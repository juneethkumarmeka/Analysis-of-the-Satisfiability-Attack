module basic_2000_20000_2500_40_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_509,In_1105);
or U1 (N_1,In_649,In_1338);
and U2 (N_2,In_1422,In_1896);
nand U3 (N_3,In_79,In_1394);
xnor U4 (N_4,In_592,In_351);
nand U5 (N_5,In_447,In_975);
and U6 (N_6,In_157,In_1525);
nand U7 (N_7,In_184,In_449);
nand U8 (N_8,In_1724,In_1624);
nand U9 (N_9,In_225,In_1985);
xnor U10 (N_10,In_810,In_1712);
nor U11 (N_11,In_947,In_913);
nand U12 (N_12,In_1894,In_1725);
xnor U13 (N_13,In_390,In_1520);
nor U14 (N_14,In_338,In_152);
or U15 (N_15,In_1884,In_937);
xnor U16 (N_16,In_1445,In_1325);
xnor U17 (N_17,In_915,In_412);
or U18 (N_18,In_1022,In_1799);
xnor U19 (N_19,In_1978,In_1284);
nor U20 (N_20,In_324,In_13);
nor U21 (N_21,In_1947,In_1072);
or U22 (N_22,In_50,In_618);
or U23 (N_23,In_1107,In_1223);
nor U24 (N_24,In_1347,In_1056);
or U25 (N_25,In_53,In_652);
nor U26 (N_26,In_678,In_172);
or U27 (N_27,In_175,In_1086);
or U28 (N_28,In_1459,In_1147);
nand U29 (N_29,In_1722,In_733);
nor U30 (N_30,In_1841,In_722);
and U31 (N_31,In_415,In_1573);
or U32 (N_32,In_1319,In_1200);
nand U33 (N_33,In_1449,In_97);
nand U34 (N_34,In_1414,In_1995);
and U35 (N_35,In_1278,In_1382);
xnor U36 (N_36,In_1388,In_740);
and U37 (N_37,In_728,In_408);
and U38 (N_38,In_761,In_307);
xor U39 (N_39,In_1025,In_567);
and U40 (N_40,In_1271,In_1345);
and U41 (N_41,In_296,In_1829);
or U42 (N_42,In_1585,In_642);
and U43 (N_43,In_1301,In_221);
and U44 (N_44,In_1914,In_884);
nor U45 (N_45,In_297,In_1583);
and U46 (N_46,In_1671,In_442);
and U47 (N_47,In_1023,In_495);
and U48 (N_48,In_630,In_811);
nor U49 (N_49,In_1146,In_207);
or U50 (N_50,In_675,In_524);
and U51 (N_51,In_1487,In_448);
and U52 (N_52,In_1685,In_1742);
xnor U53 (N_53,In_709,In_622);
or U54 (N_54,In_1792,In_1043);
or U55 (N_55,In_1352,In_1892);
or U56 (N_56,In_303,In_206);
and U57 (N_57,In_1670,In_95);
xnor U58 (N_58,In_1848,In_203);
and U59 (N_59,In_1409,In_517);
or U60 (N_60,In_1491,In_1863);
nor U61 (N_61,In_784,In_428);
and U62 (N_62,In_1898,In_596);
xnor U63 (N_63,In_269,In_1554);
nand U64 (N_64,In_1895,In_917);
and U65 (N_65,In_373,In_1603);
and U66 (N_66,In_1512,In_1996);
and U67 (N_67,In_602,In_265);
xor U68 (N_68,In_891,In_281);
nor U69 (N_69,In_781,In_289);
nor U70 (N_70,In_360,In_1210);
nand U71 (N_71,In_795,In_201);
nor U72 (N_72,In_1397,In_1622);
nor U73 (N_73,In_766,In_1256);
or U74 (N_74,In_1680,In_1068);
nor U75 (N_75,In_601,In_358);
xnor U76 (N_76,In_1510,In_1201);
or U77 (N_77,In_280,In_1618);
xor U78 (N_78,In_1953,In_1090);
or U79 (N_79,In_738,In_1251);
nor U80 (N_80,In_327,In_1366);
xnor U81 (N_81,In_1316,In_436);
xor U82 (N_82,In_1079,In_1315);
nand U83 (N_83,In_1974,In_1675);
and U84 (N_84,In_989,In_645);
or U85 (N_85,In_780,In_1800);
nor U86 (N_86,In_1137,In_1272);
or U87 (N_87,In_1760,In_1900);
nor U88 (N_88,In_246,In_1653);
nand U89 (N_89,In_1413,In_1519);
nor U90 (N_90,In_1357,In_1955);
nor U91 (N_91,In_1381,In_1172);
xor U92 (N_92,In_271,In_2);
xor U93 (N_93,In_155,In_1796);
nor U94 (N_94,In_1013,In_626);
and U95 (N_95,In_304,In_1981);
nor U96 (N_96,In_1648,In_1883);
nor U97 (N_97,In_476,In_1073);
nand U98 (N_98,In_1763,In_404);
and U99 (N_99,In_779,In_28);
nor U100 (N_100,In_341,In_1709);
or U101 (N_101,In_1836,In_1501);
nand U102 (N_102,In_123,In_922);
or U103 (N_103,In_380,In_1377);
and U104 (N_104,In_1873,In_608);
nor U105 (N_105,In_1092,In_753);
nor U106 (N_106,In_1881,In_1673);
xnor U107 (N_107,In_1493,In_229);
nand U108 (N_108,In_1007,In_597);
xor U109 (N_109,In_844,In_1729);
nand U110 (N_110,In_422,In_726);
and U111 (N_111,In_1240,In_952);
xnor U112 (N_112,In_577,In_1150);
xor U113 (N_113,In_47,In_209);
nor U114 (N_114,In_243,In_1945);
and U115 (N_115,In_1123,In_1508);
nor U116 (N_116,In_407,In_1994);
nand U117 (N_117,In_1158,In_411);
nand U118 (N_118,In_1273,In_617);
xor U119 (N_119,In_1267,In_1522);
and U120 (N_120,In_918,In_1461);
and U121 (N_121,In_39,In_1893);
or U122 (N_122,In_589,In_967);
nor U123 (N_123,In_813,In_1975);
or U124 (N_124,In_919,In_432);
and U125 (N_125,In_362,In_266);
and U126 (N_126,In_1507,In_274);
and U127 (N_127,In_1174,In_1956);
nand U128 (N_128,In_1110,In_920);
nor U129 (N_129,In_194,In_824);
xor U130 (N_130,In_1686,In_1657);
nand U131 (N_131,In_789,In_1851);
or U132 (N_132,In_1533,In_941);
xor U133 (N_133,In_1296,In_1277);
and U134 (N_134,In_292,In_790);
nor U135 (N_135,In_1921,In_174);
nand U136 (N_136,In_1918,In_1646);
nor U137 (N_137,In_1372,In_690);
xnor U138 (N_138,In_129,In_1927);
xor U139 (N_139,In_560,In_1542);
nor U140 (N_140,In_1615,In_403);
xnor U141 (N_141,In_90,In_979);
nor U142 (N_142,In_1678,In_499);
nor U143 (N_143,In_433,In_222);
nor U144 (N_144,In_725,In_775);
xnor U145 (N_145,In_89,In_809);
nor U146 (N_146,In_518,In_418);
and U147 (N_147,In_914,In_792);
nand U148 (N_148,In_664,In_859);
xor U149 (N_149,In_1517,In_992);
nand U150 (N_150,In_1323,In_1421);
nor U151 (N_151,In_1403,In_928);
or U152 (N_152,In_1604,In_333);
nand U153 (N_153,In_158,In_125);
xnor U154 (N_154,In_138,In_900);
xnor U155 (N_155,In_1327,In_1082);
and U156 (N_156,In_1489,In_530);
or U157 (N_157,In_648,In_440);
and U158 (N_158,In_774,In_854);
xnor U159 (N_159,In_425,In_434);
nand U160 (N_160,In_423,In_1130);
nand U161 (N_161,In_295,In_720);
xnor U162 (N_162,In_970,In_1784);
and U163 (N_163,In_1152,In_956);
or U164 (N_164,In_659,In_508);
nor U165 (N_165,In_1810,In_139);
xor U166 (N_166,In_549,In_1718);
or U167 (N_167,In_905,In_1039);
nor U168 (N_168,In_1915,In_1714);
xnor U169 (N_169,In_1120,In_950);
and U170 (N_170,In_1170,In_52);
nor U171 (N_171,In_598,In_1970);
and U172 (N_172,In_1085,In_543);
and U173 (N_173,In_1081,In_1231);
xnor U174 (N_174,In_1084,In_1764);
nor U175 (N_175,In_771,In_119);
nand U176 (N_176,In_1116,In_730);
xor U177 (N_177,In_1302,In_672);
or U178 (N_178,In_233,In_1404);
and U179 (N_179,In_1802,In_1237);
and U180 (N_180,In_406,In_1834);
nor U181 (N_181,In_216,In_1897);
nor U182 (N_182,In_1122,In_1570);
xnor U183 (N_183,In_122,In_1472);
nor U184 (N_184,In_1055,In_334);
nor U185 (N_185,In_1417,In_1968);
or U186 (N_186,In_1420,In_1386);
or U187 (N_187,In_977,In_888);
xor U188 (N_188,In_1650,In_200);
and U189 (N_189,In_930,In_1179);
nand U190 (N_190,In_1478,In_253);
xor U191 (N_191,In_1700,In_1854);
nand U192 (N_192,In_377,In_1053);
xor U193 (N_193,In_398,In_1629);
and U194 (N_194,In_1992,In_1496);
nand U195 (N_195,In_1463,In_1531);
or U196 (N_196,In_1115,In_706);
xnor U197 (N_197,In_1870,In_374);
nand U198 (N_198,In_646,In_1567);
nand U199 (N_199,In_1730,In_1447);
nand U200 (N_200,In_42,In_802);
xnor U201 (N_201,In_1820,In_182);
or U202 (N_202,In_1561,In_1195);
nand U203 (N_203,In_657,In_290);
nor U204 (N_204,In_1776,In_925);
xor U205 (N_205,In_559,In_1486);
or U206 (N_206,In_198,In_1581);
nor U207 (N_207,In_48,In_1415);
nor U208 (N_208,In_3,In_677);
xnor U209 (N_209,In_493,In_1088);
nand U210 (N_210,In_1750,In_1757);
or U211 (N_211,In_1346,In_1505);
or U212 (N_212,In_625,In_1249);
nor U213 (N_213,In_87,In_247);
nand U214 (N_214,In_882,In_1003);
and U215 (N_215,In_1083,In_600);
or U216 (N_216,In_1959,In_186);
or U217 (N_217,In_1363,In_825);
and U218 (N_218,In_1563,In_1100);
or U219 (N_219,In_1103,In_1441);
nand U220 (N_220,In_1954,In_1697);
or U221 (N_221,In_1126,In_556);
and U222 (N_222,In_513,In_1495);
xor U223 (N_223,In_1232,In_108);
and U224 (N_224,In_72,In_1254);
or U225 (N_225,In_1125,In_177);
or U226 (N_226,In_1479,In_1589);
xnor U227 (N_227,In_1868,In_986);
or U228 (N_228,In_1426,In_372);
xor U229 (N_229,In_1400,In_1860);
and U230 (N_230,In_263,In_1998);
xnor U231 (N_231,In_502,In_1128);
or U232 (N_232,In_1106,In_1911);
and U233 (N_233,In_1465,In_7);
and U234 (N_234,In_1824,In_717);
nand U235 (N_235,In_565,In_399);
and U236 (N_236,In_910,In_193);
or U237 (N_237,In_381,In_1818);
xnor U238 (N_238,In_591,In_829);
nand U239 (N_239,In_150,In_909);
xor U240 (N_240,In_156,In_1108);
xor U241 (N_241,In_955,In_1785);
nand U242 (N_242,In_1821,In_1932);
nand U243 (N_243,In_1234,In_583);
nand U244 (N_244,In_1687,In_1205);
xnor U245 (N_245,In_976,In_933);
nand U246 (N_246,In_1229,In_1017);
nor U247 (N_247,In_1752,In_456);
xnor U248 (N_248,In_29,In_1853);
or U249 (N_249,In_1578,In_767);
xnor U250 (N_250,In_1588,In_841);
xor U251 (N_251,In_1221,In_1934);
and U252 (N_252,In_980,In_1736);
or U253 (N_253,In_366,In_865);
xor U254 (N_254,In_587,In_1018);
nand U255 (N_255,In_356,In_18);
or U256 (N_256,In_1024,In_1064);
and U257 (N_257,In_1188,In_1194);
and U258 (N_258,In_106,In_760);
nand U259 (N_259,In_1973,In_1333);
and U260 (N_260,In_309,In_1813);
xor U261 (N_261,In_1161,In_113);
nand U262 (N_262,In_552,In_1983);
nor U263 (N_263,In_593,In_41);
and U264 (N_264,In_663,In_566);
nand U265 (N_265,In_741,In_1560);
nand U266 (N_266,In_929,In_118);
xor U267 (N_267,In_1075,In_797);
nand U268 (N_268,In_1546,In_1002);
xor U269 (N_269,In_1530,In_395);
nor U270 (N_270,In_10,In_778);
and U271 (N_271,In_91,In_1102);
or U272 (N_272,In_575,In_1539);
xor U273 (N_273,In_77,In_1300);
or U274 (N_274,In_1155,In_1708);
and U275 (N_275,In_1935,In_651);
nand U276 (N_276,In_564,In_562);
and U277 (N_277,In_852,In_335);
nor U278 (N_278,In_945,In_1384);
nand U279 (N_279,In_1861,In_1011);
nand U280 (N_280,In_671,In_429);
nor U281 (N_281,In_287,In_638);
nor U282 (N_282,In_727,In_25);
or U283 (N_283,In_1074,In_109);
xor U284 (N_284,In_595,In_1541);
or U285 (N_285,In_1497,In_1034);
and U286 (N_286,In_1875,In_629);
xor U287 (N_287,In_1839,In_1211);
xnor U288 (N_288,In_1242,In_143);
and U289 (N_289,In_951,In_528);
xor U290 (N_290,In_365,In_1795);
nand U291 (N_291,In_1250,In_537);
nand U292 (N_292,In_1966,In_161);
and U293 (N_293,In_1564,In_1499);
nor U294 (N_294,In_49,In_101);
nor U295 (N_295,In_314,In_1040);
nand U296 (N_296,In_444,In_734);
nor U297 (N_297,In_1266,In_259);
nand U298 (N_298,In_299,In_1396);
or U299 (N_299,In_1227,In_1524);
nand U300 (N_300,In_801,In_1312);
xor U301 (N_301,In_1832,In_890);
nor U302 (N_302,In_1662,In_264);
or U303 (N_303,In_704,In_896);
and U304 (N_304,In_620,In_1723);
nor U305 (N_305,In_1635,In_1288);
and U306 (N_306,In_1367,In_847);
or U307 (N_307,In_1586,In_1590);
nand U308 (N_308,In_1941,In_427);
nor U309 (N_309,In_1481,In_1735);
or U310 (N_310,In_1610,In_1297);
or U311 (N_311,In_111,In_1798);
nand U312 (N_312,In_1765,In_228);
nor U313 (N_313,In_223,In_1644);
xnor U314 (N_314,In_765,In_886);
nor U315 (N_315,In_1852,In_301);
and U316 (N_316,In_827,In_1833);
and U317 (N_317,In_1429,In_777);
and U318 (N_318,In_1702,In_1913);
nand U319 (N_319,In_145,In_1408);
and U320 (N_320,In_506,In_416);
or U321 (N_321,In_1719,In_1609);
xor U322 (N_322,In_454,In_417);
nor U323 (N_323,In_1387,In_1584);
nor U324 (N_324,In_1295,In_1807);
and U325 (N_325,In_1245,In_1849);
nor U326 (N_326,In_1940,In_1744);
or U327 (N_327,In_1690,In_1236);
or U328 (N_328,In_1926,In_1880);
nand U329 (N_329,In_1577,In_504);
and U330 (N_330,In_644,In_687);
xor U331 (N_331,In_57,In_38);
nor U332 (N_332,In_908,In_1427);
nor U333 (N_333,In_1544,In_1933);
or U334 (N_334,In_655,In_85);
nand U335 (N_335,In_1743,In_911);
and U336 (N_336,In_1480,In_545);
nor U337 (N_337,In_1777,In_569);
and U338 (N_338,In_453,In_1412);
and U339 (N_339,In_1326,In_1356);
nor U340 (N_340,In_368,In_1208);
and U341 (N_341,In_26,In_1937);
xor U342 (N_342,In_1255,In_808);
nand U343 (N_343,In_838,In_1494);
or U344 (N_344,In_514,In_519);
nor U345 (N_345,In_1141,In_1630);
or U346 (N_346,In_788,In_885);
xor U347 (N_347,In_496,In_195);
nor U348 (N_348,In_1337,In_940);
xor U349 (N_349,In_117,In_1228);
xor U350 (N_350,In_204,In_1207);
xnor U351 (N_351,In_527,In_468);
and U352 (N_352,In_1647,In_349);
nand U353 (N_353,In_165,In_308);
xnor U354 (N_354,In_192,In_1672);
or U355 (N_355,In_1734,In_58);
nand U356 (N_356,In_1938,In_189);
nand U357 (N_357,In_1238,In_60);
nor U358 (N_358,In_68,In_1485);
xnor U359 (N_359,In_1840,In_234);
nand U360 (N_360,In_379,In_1287);
and U361 (N_361,In_1909,In_1149);
and U362 (N_362,In_1104,In_628);
nand U363 (N_363,In_458,In_1948);
and U364 (N_364,In_1329,In_1314);
nand U365 (N_365,In_1607,In_751);
or U366 (N_366,In_1264,In_1661);
xnor U367 (N_367,In_872,In_553);
or U368 (N_368,In_1925,In_1021);
or U369 (N_369,In_685,In_831);
or U370 (N_370,In_1176,In_1303);
nor U371 (N_371,In_1318,In_1260);
or U372 (N_372,In_612,In_1643);
or U373 (N_373,In_1674,In_1655);
xor U374 (N_374,In_782,In_1593);
and U375 (N_375,In_1457,In_798);
nor U376 (N_376,In_1634,In_898);
nor U377 (N_377,In_864,In_742);
nand U378 (N_378,In_401,In_1866);
nor U379 (N_379,In_550,In_1339);
nand U380 (N_380,In_46,In_1929);
and U381 (N_381,In_669,In_492);
xnor U382 (N_382,In_547,In_936);
and U383 (N_383,In_1376,In_1551);
nor U384 (N_384,In_267,In_22);
nand U385 (N_385,In_213,In_1660);
or U386 (N_386,In_397,In_1317);
and U387 (N_387,In_1733,In_1825);
and U388 (N_388,In_1026,In_754);
nor U389 (N_389,In_1523,In_185);
xor U390 (N_390,In_1789,In_1191);
and U391 (N_391,In_1354,In_1448);
xnor U392 (N_392,In_1136,In_1450);
xnor U393 (N_393,In_791,In_631);
nand U394 (N_394,In_1378,In_1964);
or U395 (N_395,In_1095,In_949);
nor U396 (N_396,In_44,In_837);
and U397 (N_397,In_1716,In_1094);
and U398 (N_398,In_1342,In_1132);
nor U399 (N_399,In_953,In_1484);
and U400 (N_400,In_1117,In_1154);
nor U401 (N_401,In_993,In_100);
and U402 (N_402,In_343,In_64);
or U403 (N_403,In_1566,In_604);
xor U404 (N_404,In_1683,In_160);
or U405 (N_405,In_1721,In_1157);
nand U406 (N_406,In_1640,In_220);
or U407 (N_407,In_1035,In_1248);
and U408 (N_408,In_959,In_277);
or U409 (N_409,In_1877,In_1008);
xor U410 (N_410,In_772,In_387);
and U411 (N_411,In_839,In_261);
nor U412 (N_412,In_619,In_1440);
or U413 (N_413,In_93,In_1727);
or U414 (N_414,In_1555,In_557);
xnor U415 (N_415,In_1855,In_1202);
and U416 (N_416,In_1419,In_27);
or U417 (N_417,In_1401,In_806);
or U418 (N_418,In_1061,In_20);
or U419 (N_419,In_1768,In_1862);
or U420 (N_420,In_962,In_446);
nor U421 (N_421,In_59,In_1268);
nor U422 (N_422,In_1431,In_969);
nor U423 (N_423,In_1748,In_660);
or U424 (N_424,In_318,In_235);
nor U425 (N_425,In_1455,In_1812);
nor U426 (N_426,In_1028,In_1946);
or U427 (N_427,In_1599,In_1737);
and U428 (N_428,In_1691,In_921);
and U429 (N_429,In_1428,In_1783);
and U430 (N_430,In_1951,In_586);
xor U431 (N_431,In_450,In_36);
or U432 (N_432,In_142,In_31);
or U433 (N_433,In_1699,In_1726);
nand U434 (N_434,In_822,In_439);
or U435 (N_435,In_1867,In_357);
and U436 (N_436,In_291,In_666);
and U437 (N_437,In_252,In_1279);
nor U438 (N_438,In_1842,In_1753);
xor U439 (N_439,In_643,In_298);
nand U440 (N_440,In_856,In_799);
and U441 (N_441,In_972,In_441);
xnor U442 (N_442,In_1679,In_982);
xor U443 (N_443,In_1532,In_1121);
and U444 (N_444,In_1012,In_1321);
nor U445 (N_445,In_302,In_1416);
nand U446 (N_446,In_1649,In_83);
xor U447 (N_447,In_1580,In_997);
nand U448 (N_448,In_347,In_133);
nand U449 (N_449,In_1163,In_239);
or U450 (N_450,In_467,In_424);
and U451 (N_451,In_226,In_712);
nand U452 (N_452,In_1960,In_1451);
nand U453 (N_453,In_1715,In_1304);
nor U454 (N_454,In_98,In_762);
nand U455 (N_455,In_1475,In_1667);
or U456 (N_456,In_457,In_1059);
and U457 (N_457,In_1516,In_1626);
nand U458 (N_458,In_1473,In_1399);
nor U459 (N_459,In_743,In_1299);
xnor U460 (N_460,In_1612,In_1991);
xnor U461 (N_461,In_1693,In_1731);
nand U462 (N_462,In_964,In_1659);
xor U463 (N_463,In_238,In_1222);
xor U464 (N_464,In_103,In_756);
and U465 (N_465,In_1823,In_419);
nor U466 (N_466,In_1910,In_710);
nor U467 (N_467,In_1253,In_1889);
or U468 (N_468,In_14,In_1374);
nor U469 (N_469,In_199,In_497);
and U470 (N_470,In_627,In_361);
and U471 (N_471,In_823,In_805);
or U472 (N_472,In_74,In_578);
nand U473 (N_473,In_330,In_1771);
nor U474 (N_474,In_214,In_1182);
nand U475 (N_475,In_1280,In_1196);
nor U476 (N_476,In_178,In_948);
nor U477 (N_477,In_1423,In_1804);
nand U478 (N_478,In_1769,In_8);
nor U479 (N_479,In_535,In_1019);
and U480 (N_480,In_1052,In_1037);
or U481 (N_481,In_1676,In_662);
or U482 (N_482,In_276,In_1057);
nand U483 (N_483,In_211,In_1504);
nor U484 (N_484,In_1442,In_485);
xor U485 (N_485,In_286,In_1171);
xor U486 (N_486,In_1905,In_1952);
xnor U487 (N_487,In_1114,In_1632);
nand U488 (N_488,In_1605,In_279);
and U489 (N_489,In_674,In_255);
and U490 (N_490,In_1907,In_1269);
nand U491 (N_491,In_245,In_676);
nor U492 (N_492,In_479,In_701);
and U493 (N_493,In_1097,In_258);
nor U494 (N_494,In_268,In_1886);
nor U495 (N_495,In_376,In_606);
xor U496 (N_496,In_1193,In_1917);
and U497 (N_497,In_594,In_804);
or U498 (N_498,In_491,In_1289);
nor U499 (N_499,In_317,In_1000);
nand U500 (N_500,N_244,In_465);
and U501 (N_501,In_927,In_708);
and U502 (N_502,N_159,N_219);
or U503 (N_503,In_688,N_118);
xnor U504 (N_504,In_680,N_419);
xnor U505 (N_505,N_161,In_1212);
nor U506 (N_506,In_484,In_392);
nand U507 (N_507,In_1432,In_1741);
or U508 (N_508,N_382,In_723);
nor U509 (N_509,In_1434,In_1217);
nand U510 (N_510,N_56,N_2);
or U511 (N_511,In_1692,In_1282);
nor U512 (N_512,N_192,In_1864);
and U513 (N_513,N_110,N_234);
xnor U514 (N_514,N_367,In_906);
nor U515 (N_515,In_1131,In_1048);
xnor U516 (N_516,N_439,N_453);
and U517 (N_517,In_1828,In_869);
nand U518 (N_518,N_74,In_540);
xor U519 (N_519,N_495,In_293);
nand U520 (N_520,In_1984,N_227);
nand U521 (N_521,In_1838,N_251);
nand U522 (N_522,In_187,In_19);
nor U523 (N_523,In_1410,In_926);
or U524 (N_524,In_1856,In_1666);
nor U525 (N_525,In_78,In_1592);
or U526 (N_526,In_776,In_1540);
xor U527 (N_527,In_1930,In_582);
and U528 (N_528,In_210,N_129);
nor U529 (N_529,In_821,In_1587);
xnor U530 (N_530,N_246,In_421);
nand U531 (N_531,In_350,N_148);
and U532 (N_532,N_43,In_1305);
xor U533 (N_533,In_1270,N_135);
or U534 (N_534,In_515,In_1890);
and U535 (N_535,In_1882,In_531);
or U536 (N_536,In_320,In_636);
nor U537 (N_537,N_39,In_1140);
or U538 (N_538,In_490,In_1454);
xor U539 (N_539,In_1701,In_516);
and U540 (N_540,In_1916,In_1135);
xor U541 (N_541,In_463,In_1831);
nor U542 (N_542,In_431,N_272);
nor U543 (N_543,In_402,N_152);
nor U544 (N_544,N_353,In_1703);
or U545 (N_545,In_1383,N_311);
xnor U546 (N_546,In_147,N_40);
nand U547 (N_547,N_177,In_176);
xor U548 (N_548,In_1470,In_1569);
nand U549 (N_549,N_273,In_739);
and U550 (N_550,N_408,N_320);
and U551 (N_551,In_1936,N_326);
or U552 (N_552,In_1225,In_1732);
and U553 (N_553,N_105,In_849);
and U554 (N_554,In_1774,In_1464);
and U555 (N_555,N_405,In_24);
nor U556 (N_556,In_683,In_249);
and U557 (N_557,In_932,In_1698);
nand U558 (N_558,N_262,In_533);
nand U559 (N_559,In_1617,In_579);
and U560 (N_560,In_1625,In_637);
xor U561 (N_561,In_546,In_800);
nand U562 (N_562,In_1358,In_414);
and U563 (N_563,In_461,In_1281);
and U564 (N_564,In_1446,In_866);
nand U565 (N_565,In_632,In_1772);
nor U566 (N_566,In_1320,In_873);
nand U567 (N_567,N_21,In_1005);
nand U568 (N_568,N_255,N_238);
or U569 (N_569,In_1694,In_173);
and U570 (N_570,In_1341,In_934);
nor U571 (N_571,In_624,N_68);
nor U572 (N_572,In_251,In_105);
and U573 (N_573,In_1187,N_113);
nand U574 (N_574,In_721,N_71);
nor U575 (N_575,In_737,In_494);
or U576 (N_576,In_1198,In_700);
nor U577 (N_577,N_25,N_346);
nor U578 (N_578,N_266,N_204);
and U579 (N_579,In_505,In_1924);
or U580 (N_580,In_783,N_7);
nand U581 (N_581,In_1060,In_256);
and U582 (N_582,In_316,In_332);
xnor U583 (N_583,In_1335,In_1294);
nor U584 (N_584,In_994,In_1558);
xnor U585 (N_585,In_1355,N_137);
and U586 (N_586,In_183,In_215);
or U587 (N_587,In_1751,In_40);
and U588 (N_588,In_1596,In_1192);
nand U589 (N_589,In_724,In_435);
and U590 (N_590,In_1139,In_1990);
nor U591 (N_591,N_35,In_1247);
nor U592 (N_592,In_1490,In_466);
xor U593 (N_593,In_285,N_387);
nor U594 (N_594,In_745,N_224);
and U595 (N_595,In_682,In_999);
nor U596 (N_596,N_37,In_1901);
xnor U597 (N_597,In_471,In_1298);
xnor U598 (N_598,In_382,In_694);
nor U599 (N_599,In_1243,In_1259);
xor U600 (N_600,N_257,N_93);
nand U601 (N_601,In_375,In_590);
xor U602 (N_602,In_998,N_478);
nor U603 (N_603,In_1109,In_196);
xor U604 (N_604,In_1160,N_443);
xnor U605 (N_605,N_165,N_225);
and U606 (N_606,In_1521,In_1572);
nor U607 (N_607,N_28,In_1156);
xnor U608 (N_608,In_1579,N_190);
and U609 (N_609,In_715,N_452);
xnor U610 (N_610,In_1565,In_1912);
xnor U611 (N_611,In_654,N_446);
nand U612 (N_612,In_1613,In_814);
and U613 (N_613,N_15,In_534);
and U614 (N_614,N_427,In_75);
and U615 (N_615,In_294,N_26);
and U616 (N_616,In_526,N_116);
and U617 (N_617,In_1600,N_141);
and U618 (N_618,In_353,N_352);
nor U619 (N_619,N_0,In_803);
nand U620 (N_620,N_53,In_1185);
and U621 (N_621,In_1159,In_88);
and U622 (N_622,N_302,N_107);
or U623 (N_623,In_1393,In_1215);
nand U624 (N_624,In_963,N_319);
xor U625 (N_625,In_1226,In_481);
or U626 (N_626,In_580,In_770);
xor U627 (N_627,N_388,In_1283);
nand U628 (N_628,N_348,In_1928);
and U629 (N_629,In_1099,In_786);
and U630 (N_630,N_167,In_470);
nor U631 (N_631,N_441,In_1276);
nand U632 (N_632,In_899,In_1595);
nor U633 (N_633,In_1274,In_1636);
xnor U634 (N_634,In_984,N_8);
or U635 (N_635,N_111,In_393);
and U636 (N_636,In_988,N_145);
nand U637 (N_637,N_76,N_403);
nor U638 (N_638,In_1001,N_416);
and U639 (N_639,In_853,In_1781);
and U640 (N_640,In_958,In_1706);
xor U641 (N_641,In_1816,N_97);
or U642 (N_642,In_383,N_45);
nand U643 (N_643,N_378,In_1309);
nand U644 (N_644,In_120,N_444);
nand U645 (N_645,N_41,N_456);
and U646 (N_646,In_1754,N_98);
nand U647 (N_647,N_306,In_140);
and U648 (N_648,N_343,In_136);
xnor U649 (N_649,In_1756,N_125);
and U650 (N_650,N_373,In_313);
nand U651 (N_651,In_1656,In_1826);
or U652 (N_652,In_1373,N_278);
xnor U653 (N_653,In_1098,In_1835);
and U654 (N_654,N_428,N_289);
nor U655 (N_655,N_109,In_218);
and U656 (N_656,N_140,N_330);
or U657 (N_657,N_384,In_1214);
and U658 (N_658,In_716,N_412);
or U659 (N_659,In_149,N_150);
nor U660 (N_660,N_187,In_746);
nor U661 (N_661,N_48,In_1353);
xnor U662 (N_662,In_1552,In_1197);
xor U663 (N_663,In_56,In_1545);
nor U664 (N_664,In_699,N_166);
and U665 (N_665,In_735,In_1747);
nand U666 (N_666,N_130,In_1371);
xnor U667 (N_667,In_581,In_863);
or U668 (N_668,In_231,In_355);
nand U669 (N_669,In_840,N_312);
nand U670 (N_670,In_713,In_208);
nand U671 (N_671,In_1819,N_108);
xor U672 (N_672,In_639,In_1257);
nor U673 (N_673,N_12,In_1608);
and U674 (N_674,In_278,In_1999);
and U675 (N_675,In_34,N_196);
nand U676 (N_676,N_241,In_438);
nor U677 (N_677,In_1220,In_1285);
nor U678 (N_678,In_273,In_1350);
or U679 (N_679,In_1704,N_214);
and U680 (N_680,N_31,N_437);
nand U681 (N_681,In_469,In_1165);
or U682 (N_682,In_1045,N_142);
and U683 (N_683,N_149,N_341);
and U684 (N_684,N_497,In_154);
nand U685 (N_685,In_23,N_182);
nor U686 (N_686,N_295,N_211);
xnor U687 (N_687,In_472,In_1628);
xor U688 (N_688,N_30,N_459);
and U689 (N_689,In_1652,In_462);
or U690 (N_690,In_1637,N_83);
nor U691 (N_691,N_480,In_112);
or U692 (N_692,In_1888,In_389);
and U693 (N_693,In_1988,In_1641);
nor U694 (N_694,In_875,N_496);
and U695 (N_695,N_79,In_523);
or U696 (N_696,In_116,In_938);
and U697 (N_697,N_379,N_285);
nor U698 (N_698,N_414,In_939);
or U699 (N_699,In_310,N_163);
nand U700 (N_700,N_88,In_1986);
xnor U701 (N_701,In_1963,In_883);
nor U702 (N_702,In_61,N_374);
xor U703 (N_703,N_304,N_136);
nand U704 (N_704,In_260,N_410);
nor U705 (N_705,N_261,N_174);
nand U706 (N_706,In_661,N_6);
nor U707 (N_707,In_1456,N_393);
nand U708 (N_708,N_347,N_77);
nand U709 (N_709,N_117,N_314);
and U710 (N_710,In_148,In_284);
nand U711 (N_711,N_205,N_92);
or U712 (N_712,In_1014,In_924);
nand U713 (N_713,In_1129,In_1717);
nor U714 (N_714,N_69,In_520);
xnor U715 (N_715,In_1786,N_466);
or U716 (N_716,In_1307,N_89);
and U717 (N_717,In_443,N_194);
nor U718 (N_718,N_184,N_217);
nor U719 (N_719,In_828,N_334);
nor U720 (N_720,In_270,In_1293);
xnor U721 (N_721,In_599,In_1186);
and U722 (N_722,In_615,N_332);
nor U723 (N_723,In_966,In_1965);
or U724 (N_724,In_190,N_336);
xor U725 (N_725,N_286,In_81);
or U726 (N_726,In_1950,N_440);
or U727 (N_727,In_871,N_49);
and U728 (N_728,In_1793,N_175);
and U729 (N_729,In_1076,N_133);
or U730 (N_730,N_421,In_1275);
or U731 (N_731,N_323,N_366);
nand U732 (N_732,In_257,In_32);
and U733 (N_733,In_614,N_270);
and U734 (N_734,In_45,N_297);
xnor U735 (N_735,N_147,In_71);
nand U736 (N_736,In_227,In_410);
and U737 (N_737,In_237,In_1391);
and U738 (N_738,In_1111,N_247);
xnor U739 (N_739,N_164,N_260);
nor U740 (N_740,In_254,In_1536);
or U741 (N_741,In_1474,N_60);
nor U742 (N_742,In_1920,In_1844);
and U743 (N_743,N_402,N_123);
nor U744 (N_744,N_423,In_1906);
nor U745 (N_745,N_18,In_1550);
and U746 (N_746,N_328,In_501);
and U747 (N_747,N_114,N_181);
nand U748 (N_748,In_971,In_1462);
and U749 (N_749,In_1958,N_256);
and U750 (N_750,N_386,In_110);
nor U751 (N_751,N_377,In_692);
and U752 (N_752,N_360,In_1483);
nand U753 (N_753,In_1181,In_1601);
or U754 (N_754,In_1746,In_968);
nand U755 (N_755,In_785,In_1993);
or U756 (N_756,N_58,In_1395);
xnor U757 (N_757,N_209,In_1817);
nand U758 (N_758,In_0,N_121);
or U759 (N_759,N_33,In_473);
or U760 (N_760,N_356,In_224);
nor U761 (N_761,In_92,In_641);
nor U762 (N_762,In_17,In_1885);
and U763 (N_763,In_188,In_1939);
or U764 (N_764,In_1364,N_212);
and U765 (N_765,In_344,In_1847);
nand U766 (N_766,In_1639,In_37);
nor U767 (N_767,N_14,In_1113);
nand U768 (N_768,In_329,N_34);
nor U769 (N_769,In_80,In_342);
and U770 (N_770,In_127,In_1096);
nor U771 (N_771,In_115,N_27);
or U772 (N_772,In_1290,In_719);
and U773 (N_773,N_442,In_820);
nor U774 (N_774,N_363,In_340);
nand U775 (N_775,In_987,In_1582);
and U776 (N_776,In_1411,N_216);
or U777 (N_777,In_1989,In_300);
xnor U778 (N_778,N_430,In_1511);
nor U779 (N_779,In_146,In_679);
and U780 (N_780,In_748,In_529);
or U781 (N_781,In_850,In_345);
nand U782 (N_782,N_265,In_1077);
nand U783 (N_783,N_372,In_191);
xnor U784 (N_784,In_525,In_1070);
and U785 (N_785,In_76,In_607);
nor U786 (N_786,In_1611,In_460);
nand U787 (N_787,N_447,N_395);
and U788 (N_788,In_1943,In_1620);
or U789 (N_789,In_1534,In_1328);
nor U790 (N_790,In_1859,N_154);
and U791 (N_791,In_554,N_19);
and U792 (N_792,N_51,In_1801);
nor U793 (N_793,N_476,In_539);
nor U794 (N_794,In_1169,In_833);
and U795 (N_795,In_510,N_55);
or U796 (N_796,N_344,In_507);
xnor U797 (N_797,In_1931,In_1425);
or U798 (N_798,N_417,N_84);
and U799 (N_799,N_299,In_319);
and U800 (N_800,In_879,In_1553);
xnor U801 (N_801,N_325,In_1961);
xnor U802 (N_802,N_385,N_127);
and U803 (N_803,N_94,In_749);
and U804 (N_804,In_1591,In_1846);
nand U805 (N_805,In_1224,In_695);
nand U806 (N_806,In_1684,In_1173);
and U807 (N_807,N_86,In_1324);
nand U808 (N_808,N_337,N_482);
and U809 (N_809,N_349,In_634);
nor U810 (N_810,N_143,In_1468);
or U811 (N_811,N_90,In_306);
and U812 (N_812,In_1788,N_342);
or U813 (N_813,In_1665,In_1642);
or U814 (N_814,N_1,In_475);
xor U815 (N_815,In_1261,In_1502);
or U816 (N_816,In_1518,In_1619);
nand U817 (N_817,In_478,In_1044);
xor U818 (N_818,In_114,In_862);
or U819 (N_819,In_1368,N_100);
nand U820 (N_820,In_54,In_1969);
nor U821 (N_821,N_425,In_130);
and U822 (N_822,In_315,In_1526);
nor U823 (N_823,In_877,In_1677);
nor U824 (N_824,N_406,In_826);
xnor U825 (N_825,In_703,N_485);
nand U826 (N_826,In_1923,In_647);
nor U827 (N_827,N_243,In_354);
nand U828 (N_828,In_1015,N_193);
and U829 (N_829,N_433,In_684);
and U830 (N_830,In_1543,In_1392);
and U831 (N_831,In_1987,In_1230);
and U832 (N_832,N_345,N_280);
and U833 (N_833,In_558,In_1244);
nor U834 (N_834,In_1087,N_106);
or U835 (N_835,N_279,In_352);
or U836 (N_836,N_274,In_691);
and U837 (N_837,N_358,In_794);
or U838 (N_838,N_350,In_755);
and U839 (N_839,In_1047,N_488);
or U840 (N_840,In_990,N_245);
nor U841 (N_841,In_1379,In_1791);
and U842 (N_842,In_1433,N_321);
or U843 (N_843,N_375,In_1738);
and U844 (N_844,N_80,In_1492);
or U845 (N_845,In_1405,N_22);
nor U846 (N_846,In_141,In_1488);
or U847 (N_847,In_1498,N_200);
xnor U848 (N_848,N_239,In_1334);
nand U849 (N_849,In_1979,In_665);
nand U850 (N_850,In_656,N_486);
xnor U851 (N_851,N_73,In_860);
xnor U852 (N_852,In_282,In_30);
nand U853 (N_853,In_1203,In_452);
or U854 (N_854,N_47,N_310);
or U855 (N_855,In_1857,In_322);
xnor U856 (N_856,In_170,In_217);
or U857 (N_857,In_576,N_481);
nor U858 (N_858,In_732,N_383);
nand U859 (N_859,In_983,In_1209);
or U860 (N_860,In_616,N_70);
xnor U861 (N_861,In_1904,N_368);
and U862 (N_862,In_1407,N_242);
nor U863 (N_863,In_1042,In_769);
xor U864 (N_864,In_121,In_548);
nor U865 (N_865,In_1658,N_198);
or U866 (N_866,In_288,In_9);
or U867 (N_867,In_511,In_1361);
nand U868 (N_868,N_369,N_138);
nand U869 (N_869,In_1980,In_1899);
nand U870 (N_870,In_1453,In_845);
and U871 (N_871,In_1571,N_499);
and U872 (N_872,In_610,In_1503);
or U873 (N_873,In_339,In_336);
nor U874 (N_874,In_1041,In_1547);
nand U875 (N_875,In_241,In_151);
nand U876 (N_876,N_120,N_23);
or U877 (N_877,In_892,N_426);
xor U878 (N_878,N_315,N_489);
nand U879 (N_879,In_521,In_1779);
and U880 (N_880,N_288,N_355);
and U881 (N_881,In_916,N_78);
nand U882 (N_882,In_1168,N_54);
nand U883 (N_883,N_240,In_1471);
nor U884 (N_884,N_458,N_20);
and U885 (N_885,In_584,In_1054);
and U886 (N_886,N_479,In_759);
nor U887 (N_887,In_1286,In_1167);
nor U888 (N_888,In_1443,In_1606);
nand U889 (N_889,In_1466,In_1755);
and U890 (N_890,N_407,In_1476);
nor U891 (N_891,N_206,In_1614);
and U892 (N_892,In_1009,N_188);
or U893 (N_893,N_221,In_830);
and U894 (N_894,N_253,N_418);
nand U895 (N_895,In_1770,N_170);
xnor U896 (N_896,In_1668,N_329);
and U897 (N_897,In_1038,In_1576);
nor U898 (N_898,N_61,N_85);
nor U899 (N_899,N_483,In_1124);
nand U900 (N_900,N_354,N_264);
xnor U901 (N_901,In_1809,N_237);
or U902 (N_902,In_1438,In_698);
or U903 (N_903,In_104,In_1696);
or U904 (N_904,In_551,In_1664);
nand U905 (N_905,In_832,In_1233);
nor U906 (N_906,In_1942,In_1362);
or U907 (N_907,In_1291,In_1265);
nor U908 (N_908,In_1344,In_1878);
and U909 (N_909,In_359,In_846);
nor U910 (N_910,In_420,N_131);
and U911 (N_911,N_228,In_673);
and U912 (N_912,In_394,In_1811);
nand U913 (N_913,N_498,In_1380);
nand U914 (N_914,In_1199,In_834);
or U915 (N_915,In_328,N_308);
nor U916 (N_916,In_1213,In_1982);
or U917 (N_917,In_1654,N_226);
or U918 (N_918,In_391,In_1313);
nand U919 (N_919,N_210,N_411);
nor U920 (N_920,In_902,In_1621);
xor U921 (N_921,N_208,In_1252);
xor U922 (N_922,In_1069,In_69);
nor U923 (N_923,In_1967,In_995);
nand U924 (N_924,N_119,N_450);
xnor U925 (N_925,N_335,In_35);
and U926 (N_926,In_1051,In_135);
xnor U927 (N_927,In_144,N_178);
nor U928 (N_928,In_1365,In_681);
nand U929 (N_929,In_1311,N_477);
and U930 (N_930,N_317,In_1976);
and U931 (N_931,N_156,N_461);
nand U932 (N_932,In_126,N_397);
nor U933 (N_933,N_268,N_296);
nand U934 (N_934,In_842,In_965);
nand U935 (N_935,In_179,N_236);
and U936 (N_936,In_1216,N_454);
nand U937 (N_937,N_294,In_1134);
and U938 (N_938,In_1308,N_422);
xnor U939 (N_939,N_235,In_1127);
nand U940 (N_940,N_112,In_66);
and U941 (N_941,In_1067,In_131);
nand U942 (N_942,In_67,In_793);
xor U943 (N_943,In_1370,In_538);
or U944 (N_944,N_487,In_413);
nor U945 (N_945,N_464,N_364);
nor U946 (N_946,N_173,N_11);
or U947 (N_947,In_1340,In_689);
nor U948 (N_948,N_168,In_1437);
and U949 (N_949,N_316,In_693);
nor U950 (N_950,N_313,N_465);
xnor U951 (N_951,In_752,In_312);
nand U952 (N_952,In_1118,N_176);
nand U953 (N_953,In_1235,In_1027);
or U954 (N_954,In_244,N_468);
nor U955 (N_955,In_1616,In_1598);
nor U956 (N_956,N_5,In_1310);
or U957 (N_957,In_166,In_1469);
or U958 (N_958,In_996,N_132);
or U959 (N_959,N_438,In_63);
nand U960 (N_960,In_65,In_62);
xor U961 (N_961,In_262,In_500);
or U962 (N_962,N_104,N_259);
or U963 (N_963,In_1062,In_718);
nor U964 (N_964,In_1369,In_1871);
or U965 (N_965,In_82,In_1359);
xnor U966 (N_966,In_757,In_532);
xor U967 (N_967,In_1548,In_981);
nand U968 (N_968,In_1773,In_571);
xor U969 (N_969,N_415,In_1375);
and U970 (N_970,In_137,N_380);
nand U971 (N_971,In_961,N_409);
nor U972 (N_972,In_1594,N_394);
nor U973 (N_973,N_24,In_1360);
and U974 (N_974,In_219,In_807);
nand U975 (N_975,N_122,In_1033);
or U976 (N_976,N_186,In_897);
or U977 (N_977,In_1239,In_653);
nor U978 (N_978,In_482,N_324);
nor U979 (N_979,In_1049,N_81);
and U980 (N_980,In_1145,N_162);
xor U981 (N_981,N_371,In_1740);
or U982 (N_982,In_1262,In_385);
nand U983 (N_983,In_498,In_55);
nor U984 (N_984,N_263,In_1138);
or U985 (N_985,In_1500,N_115);
and U986 (N_986,In_667,N_213);
xor U987 (N_987,N_460,In_1790);
nor U988 (N_988,N_404,N_36);
nor U989 (N_989,In_574,In_773);
and U990 (N_990,In_640,N_359);
nand U991 (N_991,In_1477,In_1759);
xor U992 (N_992,N_381,N_473);
or U993 (N_993,In_1997,In_702);
nand U994 (N_994,N_215,In_205);
nor U995 (N_995,In_1631,N_431);
and U996 (N_996,In_605,In_1803);
and U997 (N_997,In_459,In_409);
nor U998 (N_998,N_435,In_1663);
or U999 (N_999,In_1874,In_163);
or U1000 (N_1000,N_538,N_50);
xor U1001 (N_1001,In_1066,N_955);
and U1002 (N_1002,N_782,In_1460);
nor U1003 (N_1003,N_362,N_815);
nand U1004 (N_1004,In_168,N_508);
xor U1005 (N_1005,In_1713,N_637);
and U1006 (N_1006,N_868,In_696);
nand U1007 (N_1007,In_974,N_757);
xnor U1008 (N_1008,N_980,In_1903);
xnor U1009 (N_1009,N_233,N_462);
nor U1010 (N_1010,In_1183,In_86);
nand U1011 (N_1011,In_668,N_770);
nor U1012 (N_1012,N_704,N_391);
nor U1013 (N_1013,N_959,N_972);
and U1014 (N_1014,In_369,In_812);
and U1015 (N_1015,N_976,N_854);
and U1016 (N_1016,N_886,N_604);
nand U1017 (N_1017,N_715,In_796);
nand U1018 (N_1018,N_936,In_386);
nand U1019 (N_1019,In_1843,In_1681);
and U1020 (N_1020,N_361,In_881);
nand U1021 (N_1021,N_928,In_613);
nor U1022 (N_1022,In_396,N_605);
nand U1023 (N_1023,N_678,N_768);
nor U1024 (N_1024,N_275,In_1827);
or U1025 (N_1025,N_911,In_1845);
nand U1026 (N_1026,N_57,N_277);
xnor U1027 (N_1027,In_1010,In_1922);
and U1028 (N_1028,N_822,In_1837);
and U1029 (N_1029,N_682,N_941);
nor U1030 (N_1030,N_666,In_585);
or U1031 (N_1031,N_207,In_1876);
and U1032 (N_1032,N_4,In_1142);
xor U1033 (N_1033,N_281,N_449);
nand U1034 (N_1034,N_847,N_101);
nand U1035 (N_1035,N_844,N_721);
or U1036 (N_1036,In_51,N_624);
nor U1037 (N_1037,N_665,N_744);
nand U1038 (N_1038,In_991,In_1306);
nor U1039 (N_1039,N_622,In_946);
or U1040 (N_1040,N_613,N_523);
nor U1041 (N_1041,In_363,N_396);
nor U1042 (N_1042,In_16,In_1241);
or U1043 (N_1043,In_1908,In_1292);
and U1044 (N_1044,N_659,N_837);
or U1045 (N_1045,N_572,N_983);
nor U1046 (N_1046,In_1112,N_559);
nand U1047 (N_1047,N_191,N_484);
nor U1048 (N_1048,N_796,N_231);
xnor U1049 (N_1049,N_520,In_1151);
xnor U1050 (N_1050,N_158,N_725);
nand U1051 (N_1051,N_964,N_755);
nor U1052 (N_1052,In_1538,N_608);
xor U1053 (N_1053,In_405,N_694);
or U1054 (N_1054,In_563,In_1865);
xor U1055 (N_1055,N_917,In_73);
nand U1056 (N_1056,N_580,In_570);
nand U1057 (N_1057,N_989,N_541);
or U1058 (N_1058,N_745,N_685);
nor U1059 (N_1059,In_1078,In_236);
and U1060 (N_1060,In_1148,In_711);
xor U1061 (N_1061,In_70,In_895);
or U1062 (N_1062,N_970,N_649);
or U1063 (N_1063,N_290,In_1418);
xor U1064 (N_1064,N_988,N_436);
nand U1065 (N_1065,N_893,N_820);
or U1066 (N_1066,N_399,N_775);
nor U1067 (N_1067,In_544,In_107);
or U1068 (N_1068,N_871,In_21);
nor U1069 (N_1069,N_612,N_772);
nor U1070 (N_1070,N_303,In_388);
and U1071 (N_1071,In_483,N_690);
or U1072 (N_1072,N_500,N_203);
xnor U1073 (N_1073,N_590,N_891);
xnor U1074 (N_1074,N_475,In_705);
and U1075 (N_1075,N_327,N_581);
and U1076 (N_1076,In_973,In_1030);
nand U1077 (N_1077,N_522,In_1556);
or U1078 (N_1078,N_810,In_819);
and U1079 (N_1079,N_639,N_492);
xor U1080 (N_1080,N_863,N_783);
xnor U1081 (N_1081,In_1004,In_1549);
or U1082 (N_1082,N_573,In_474);
nor U1083 (N_1083,N_888,In_954);
nor U1084 (N_1084,N_636,In_488);
nand U1085 (N_1085,N_987,In_1080);
nor U1086 (N_1086,N_67,N_986);
and U1087 (N_1087,In_1815,N_931);
or U1088 (N_1088,In_164,N_708);
or U1089 (N_1089,N_786,N_900);
and U1090 (N_1090,In_96,N_897);
and U1091 (N_1091,N_699,In_128);
nor U1092 (N_1092,N_218,In_1133);
and U1093 (N_1093,N_128,In_371);
or U1094 (N_1094,In_1190,N_518);
xor U1095 (N_1095,N_940,N_753);
and U1096 (N_1096,N_773,N_562);
nor U1097 (N_1097,In_1535,In_1602);
nor U1098 (N_1098,N_766,N_776);
or U1099 (N_1099,In_1218,In_1206);
or U1100 (N_1100,In_1872,N_656);
nand U1101 (N_1101,N_514,In_250);
and U1102 (N_1102,In_1575,N_826);
xnor U1103 (N_1103,N_183,N_630);
nor U1104 (N_1104,In_848,In_758);
nor U1105 (N_1105,N_827,N_392);
xnor U1106 (N_1106,N_287,N_781);
nand U1107 (N_1107,In_1514,N_66);
or U1108 (N_1108,In_763,N_709);
xor U1109 (N_1109,In_1063,N_856);
xor U1110 (N_1110,In_1794,N_223);
and U1111 (N_1111,N_716,In_768);
or U1112 (N_1112,In_1006,N_924);
xor U1113 (N_1113,N_977,N_501);
nand U1114 (N_1114,N_582,In_868);
or U1115 (N_1115,N_723,In_124);
or U1116 (N_1116,N_915,N_851);
and U1117 (N_1117,In_348,N_575);
nor U1118 (N_1118,N_926,In_818);
xor U1119 (N_1119,N_880,N_777);
nand U1120 (N_1120,N_293,In_1020);
nand U1121 (N_1121,N_904,N_29);
xnor U1122 (N_1122,N_735,In_815);
xor U1123 (N_1123,N_17,N_700);
and U1124 (N_1124,N_677,N_724);
xnor U1125 (N_1125,N_623,N_13);
xnor U1126 (N_1126,N_706,N_617);
nand U1127 (N_1127,N_401,In_985);
nor U1128 (N_1128,N_146,N_890);
xnor U1129 (N_1129,N_606,N_570);
and U1130 (N_1130,In_744,N_512);
nor U1131 (N_1131,N_560,In_326);
xnor U1132 (N_1132,In_202,N_788);
nor U1133 (N_1133,N_370,In_904);
and U1134 (N_1134,N_919,N_833);
nor U1135 (N_1135,N_874,N_519);
xor U1136 (N_1136,N_865,N_730);
xnor U1137 (N_1137,N_843,In_1153);
nand U1138 (N_1138,In_1879,N_771);
and U1139 (N_1139,In_750,N_944);
nand U1140 (N_1140,In_1482,N_791);
nor U1141 (N_1141,N_920,N_197);
nor U1142 (N_1142,N_185,N_935);
nor U1143 (N_1143,N_722,N_797);
nand U1144 (N_1144,N_599,In_1390);
and U1145 (N_1145,N_269,N_248);
or U1146 (N_1146,N_832,N_276);
and U1147 (N_1147,In_171,N_565);
xnor U1148 (N_1148,N_503,N_583);
nand U1149 (N_1149,N_713,In_907);
nand U1150 (N_1150,N_710,N_870);
nor U1151 (N_1151,N_884,N_852);
and U1152 (N_1152,N_841,N_591);
or U1153 (N_1153,N_738,N_739);
nor U1154 (N_1154,In_729,In_650);
nor U1155 (N_1155,N_63,N_764);
or U1156 (N_1156,N_938,In_230);
or U1157 (N_1157,N_793,N_648);
and U1158 (N_1158,N_829,N_937);
and U1159 (N_1159,In_1184,N_697);
nand U1160 (N_1160,In_1031,N_711);
nor U1161 (N_1161,In_1430,N_760);
nand U1162 (N_1162,N_653,In_1089);
or U1163 (N_1163,In_1246,N_676);
and U1164 (N_1164,N_470,In_1204);
nor U1165 (N_1165,N_905,In_686);
nand U1166 (N_1166,N_635,N_814);
and U1167 (N_1167,N_547,In_240);
nor U1168 (N_1168,N_860,N_284);
and U1169 (N_1169,N_762,N_990);
xor U1170 (N_1170,N_953,N_620);
nand U1171 (N_1171,N_967,In_169);
nand U1172 (N_1172,In_861,N_201);
or U1173 (N_1173,In_855,N_564);
or U1174 (N_1174,N_758,In_181);
and U1175 (N_1175,N_340,N_979);
nor U1176 (N_1176,In_33,In_878);
nand U1177 (N_1177,N_601,N_567);
or U1178 (N_1178,In_1119,N_550);
or U1179 (N_1179,N_835,N_463);
xnor U1180 (N_1180,N_655,N_712);
and U1181 (N_1181,N_72,N_579);
or U1182 (N_1182,N_526,In_1633);
nand U1183 (N_1183,N_309,N_333);
and U1184 (N_1184,In_912,N_513);
or U1185 (N_1185,In_1452,N_803);
or U1186 (N_1186,N_647,N_658);
xor U1187 (N_1187,In_1651,N_997);
or U1188 (N_1188,N_999,N_740);
xor U1189 (N_1189,N_864,N_857);
or U1190 (N_1190,N_792,N_491);
nor U1191 (N_1191,N_530,N_292);
nor U1192 (N_1192,N_674,In_1745);
and U1193 (N_1193,In_903,N_602);
xor U1194 (N_1194,N_763,In_132);
xor U1195 (N_1195,N_151,In_1189);
xor U1196 (N_1196,N_966,N_515);
or U1197 (N_1197,N_831,N_958);
and U1198 (N_1198,N_534,N_918);
and U1199 (N_1199,In_935,N_254);
xor U1200 (N_1200,N_848,N_896);
and U1201 (N_1201,In_1762,N_688);
and U1202 (N_1202,In_489,N_413);
xnor U1203 (N_1203,N_646,N_734);
xor U1204 (N_1204,In_1949,In_1797);
or U1205 (N_1205,N_774,N_322);
xnor U1206 (N_1206,N_10,N_853);
xnor U1207 (N_1207,N_859,N_202);
nand U1208 (N_1208,In_1623,N_532);
nand U1209 (N_1209,In_487,N_574);
nor U1210 (N_1210,In_889,N_737);
nor U1211 (N_1211,N_875,In_1780);
and U1212 (N_1212,In_1065,N_616);
nor U1213 (N_1213,In_747,N_651);
nor U1214 (N_1214,N_943,In_1219);
or U1215 (N_1215,In_787,In_858);
xor U1216 (N_1216,N_907,N_765);
nand U1217 (N_1217,N_895,N_785);
nand U1218 (N_1218,In_43,In_816);
or U1219 (N_1219,N_806,In_817);
nand U1220 (N_1220,In_364,N_873);
or U1221 (N_1221,N_729,N_642);
and U1222 (N_1222,In_1091,N_157);
xnor U1223 (N_1223,N_555,N_930);
xor U1224 (N_1224,In_923,N_759);
or U1225 (N_1225,N_179,N_539);
and U1226 (N_1226,In_503,N_593);
xnor U1227 (N_1227,N_645,N_301);
xnor U1228 (N_1228,N_736,In_542);
nand U1229 (N_1229,N_102,In_180);
xor U1230 (N_1230,N_790,In_1330);
or U1231 (N_1231,In_437,In_1406);
nor U1232 (N_1232,N_691,N_511);
nor U1233 (N_1233,N_921,In_6);
and U1234 (N_1234,In_311,N_641);
nand U1235 (N_1235,In_880,In_572);
nand U1236 (N_1236,N_922,In_573);
xnor U1237 (N_1237,N_657,N_742);
nor U1238 (N_1238,In_1180,N_586);
xnor U1239 (N_1239,N_733,N_628);
and U1240 (N_1240,N_172,In_1778);
or U1241 (N_1241,In_1739,In_1775);
nor U1242 (N_1242,N_684,N_732);
nor U1243 (N_1243,In_1143,N_846);
and U1244 (N_1244,N_300,In_455);
and U1245 (N_1245,N_885,N_821);
xnor U1246 (N_1246,N_795,In_1711);
or U1247 (N_1247,N_950,In_1);
xnor U1248 (N_1248,In_960,In_94);
nor U1249 (N_1249,N_878,In_876);
or U1250 (N_1250,N_189,In_367);
and U1251 (N_1251,In_1814,N_751);
or U1252 (N_1252,N_934,In_1175);
or U1253 (N_1253,N_91,N_801);
and U1254 (N_1254,In_1971,In_835);
nor U1255 (N_1255,N_524,N_981);
and U1256 (N_1256,N_720,N_991);
nor U1257 (N_1257,In_159,N_982);
nand U1258 (N_1258,In_1162,N_726);
nand U1259 (N_1259,N_536,N_675);
xor U1260 (N_1260,N_872,N_563);
or U1261 (N_1261,N_747,N_861);
or U1262 (N_1262,In_1919,N_610);
xor U1263 (N_1263,N_927,In_764);
xor U1264 (N_1264,N_794,N_472);
nor U1265 (N_1265,In_867,N_728);
nor U1266 (N_1266,N_467,N_933);
nor U1267 (N_1267,N_42,N_968);
nor U1268 (N_1268,N_546,In_400);
xor U1269 (N_1269,N_901,N_561);
xnor U1270 (N_1270,In_1050,In_843);
or U1271 (N_1271,N_578,In_321);
nor U1272 (N_1272,In_1568,N_683);
xor U1273 (N_1273,In_1164,N_879);
xor U1274 (N_1274,N_834,In_870);
or U1275 (N_1275,N_705,In_1444);
and U1276 (N_1276,N_680,In_283);
nor U1277 (N_1277,N_898,N_855);
xnor U1278 (N_1278,In_212,In_305);
nand U1279 (N_1279,In_931,N_695);
nand U1280 (N_1280,N_965,N_974);
nor U1281 (N_1281,N_65,In_1758);
nand U1282 (N_1282,N_818,N_502);
or U1283 (N_1283,N_3,In_480);
xnor U1284 (N_1284,N_544,N_625);
and U1285 (N_1285,N_681,In_874);
and U1286 (N_1286,N_126,In_1032);
nor U1287 (N_1287,In_1962,N_634);
or U1288 (N_1288,In_248,In_1029);
nor U1289 (N_1289,N_761,In_603);
and U1290 (N_1290,N_894,N_445);
xor U1291 (N_1291,In_1336,N_619);
xnor U1292 (N_1292,N_957,N_517);
nand U1293 (N_1293,N_881,In_1389);
xnor U1294 (N_1294,In_541,N_542);
xnor U1295 (N_1295,N_96,In_242);
or U1296 (N_1296,N_588,N_836);
nor U1297 (N_1297,In_731,N_516);
xnor U1298 (N_1298,N_670,N_660);
and U1299 (N_1299,N_587,N_800);
xor U1300 (N_1300,N_731,In_153);
xor U1301 (N_1301,In_1343,In_736);
xnor U1302 (N_1302,N_995,N_823);
nand U1303 (N_1303,N_535,N_845);
or U1304 (N_1304,N_808,N_714);
nand U1305 (N_1305,In_944,N_64);
or U1306 (N_1306,N_903,In_1529);
nand U1307 (N_1307,N_929,In_1705);
nand U1308 (N_1308,N_945,In_1806);
xnor U1309 (N_1309,N_95,N_99);
or U1310 (N_1310,N_932,N_153);
and U1311 (N_1311,In_1178,N_631);
nand U1312 (N_1312,In_12,N_789);
and U1313 (N_1313,N_38,N_671);
nor U1314 (N_1314,N_663,N_828);
and U1315 (N_1315,In_555,In_197);
nand U1316 (N_1316,N_595,N_271);
nor U1317 (N_1317,N_862,N_975);
or U1318 (N_1318,N_994,N_305);
and U1319 (N_1319,In_658,In_325);
or U1320 (N_1320,In_1627,N_925);
xor U1321 (N_1321,In_588,N_180);
nor U1322 (N_1322,N_858,N_672);
or U1323 (N_1323,N_16,N_597);
nand U1324 (N_1324,N_804,N_52);
or U1325 (N_1325,In_697,In_1822);
nand U1326 (N_1326,In_1557,N_780);
and U1327 (N_1327,In_346,N_553);
xor U1328 (N_1328,N_521,N_510);
or U1329 (N_1329,N_155,In_370);
nand U1330 (N_1330,N_252,In_11);
xor U1331 (N_1331,N_509,N_199);
or U1332 (N_1332,In_1850,In_384);
xor U1333 (N_1333,N_506,N_883);
nor U1334 (N_1334,N_557,In_901);
nor U1335 (N_1335,N_457,N_973);
and U1336 (N_1336,N_961,N_842);
and U1337 (N_1337,N_830,In_1805);
and U1338 (N_1338,N_229,In_1527);
xnor U1339 (N_1339,N_719,N_916);
nor U1340 (N_1340,N_906,N_993);
or U1341 (N_1341,N_171,N_626);
xnor U1342 (N_1342,N_82,N_507);
nand U1343 (N_1343,N_494,N_638);
or U1344 (N_1344,In_4,In_512);
or U1345 (N_1345,In_1902,In_1351);
and U1346 (N_1346,N_490,N_839);
and U1347 (N_1347,In_714,N_331);
or U1348 (N_1348,N_661,N_779);
nand U1349 (N_1349,In_1513,In_1036);
xor U1350 (N_1350,N_551,In_1385);
nor U1351 (N_1351,In_84,N_752);
nor U1352 (N_1352,In_1537,In_1695);
or U1353 (N_1353,N_568,N_451);
xnor U1354 (N_1354,N_669,N_954);
or U1355 (N_1355,In_943,N_432);
xor U1356 (N_1356,N_840,N_869);
nand U1357 (N_1357,N_769,N_650);
or U1358 (N_1358,In_430,In_331);
xor U1359 (N_1359,N_679,N_813);
nand U1360 (N_1360,In_337,N_338);
nor U1361 (N_1361,In_894,In_1515);
nand U1362 (N_1362,N_914,In_1638);
xnor U1363 (N_1363,N_689,N_420);
or U1364 (N_1364,N_632,N_250);
or U1365 (N_1365,In_1263,N_942);
or U1366 (N_1366,N_767,In_1559);
xor U1367 (N_1367,N_799,N_46);
nand U1368 (N_1368,N_139,In_836);
nand U1369 (N_1369,In_1348,In_1689);
nor U1370 (N_1370,In_477,N_577);
nor U1371 (N_1371,N_662,N_640);
nand U1372 (N_1372,N_947,N_543);
nand U1373 (N_1373,N_529,In_1957);
nor U1374 (N_1374,N_971,N_998);
nand U1375 (N_1375,In_15,N_717);
xor U1376 (N_1376,N_504,N_748);
and U1377 (N_1377,N_889,In_451);
nor U1378 (N_1378,In_1177,In_1766);
or U1379 (N_1379,N_819,N_448);
or U1380 (N_1380,N_908,N_62);
nand U1381 (N_1381,N_727,N_357);
nand U1382 (N_1382,In_1562,N_609);
and U1383 (N_1383,N_592,In_1688);
and U1384 (N_1384,N_817,N_692);
and U1385 (N_1385,N_32,N_554);
or U1386 (N_1386,N_960,N_985);
or U1387 (N_1387,N_627,In_232);
or U1388 (N_1388,N_87,N_812);
nand U1389 (N_1389,N_258,N_389);
or U1390 (N_1390,N_603,N_594);
or U1391 (N_1391,In_851,In_464);
or U1392 (N_1392,N_741,In_1787);
nand U1393 (N_1393,In_1891,N_558);
nor U1394 (N_1394,N_667,In_167);
xor U1395 (N_1395,N_144,N_615);
and U1396 (N_1396,N_505,N_249);
and U1397 (N_1397,In_1322,In_1093);
and U1398 (N_1398,In_609,N_339);
nand U1399 (N_1399,In_1645,N_291);
xnor U1400 (N_1400,N_802,In_1869);
nand U1401 (N_1401,N_984,In_162);
xor U1402 (N_1402,N_298,N_307);
nor U1403 (N_1403,In_1720,In_1682);
nand U1404 (N_1404,In_536,In_1071);
nor U1405 (N_1405,N_702,In_1506);
xnor U1406 (N_1406,In_568,N_811);
nor U1407 (N_1407,In_522,N_556);
and U1408 (N_1408,N_754,In_272);
xor U1409 (N_1409,N_525,N_548);
xor U1410 (N_1410,In_1398,N_493);
xnor U1411 (N_1411,In_445,N_805);
xnor U1412 (N_1412,N_824,N_816);
and U1413 (N_1413,N_687,N_571);
xor U1414 (N_1414,N_912,N_825);
nor U1415 (N_1415,N_877,N_232);
nor U1416 (N_1416,N_698,N_696);
or U1417 (N_1417,N_267,N_282);
or U1418 (N_1418,In_1402,In_486);
or U1419 (N_1419,N_549,N_621);
nor U1420 (N_1420,N_633,N_756);
and U1421 (N_1421,N_283,N_629);
and U1422 (N_1422,In_1101,In_1858);
nand U1423 (N_1423,N_607,N_913);
and U1424 (N_1424,N_952,N_614);
and U1425 (N_1425,N_44,N_956);
xnor U1426 (N_1426,In_1830,N_222);
nand U1427 (N_1427,N_784,In_1728);
nor U1428 (N_1428,N_9,N_531);
or U1429 (N_1429,N_618,In_635);
xnor U1430 (N_1430,In_1887,N_668);
nand U1431 (N_1431,In_942,N_598);
or U1432 (N_1432,N_566,N_134);
nor U1433 (N_1433,In_1574,In_5);
nand U1434 (N_1434,In_1016,N_537);
nand U1435 (N_1435,N_807,N_400);
nand U1436 (N_1436,In_1258,N_923);
xor U1437 (N_1437,In_1331,N_643);
nor U1438 (N_1438,N_746,N_743);
xor U1439 (N_1439,N_398,In_1767);
nand U1440 (N_1440,N_429,N_750);
and U1441 (N_1441,N_701,In_134);
xnor U1442 (N_1442,In_1424,N_474);
xnor U1443 (N_1443,In_1332,N_527);
nand U1444 (N_1444,N_946,N_169);
xor U1445 (N_1445,In_1597,N_652);
or U1446 (N_1446,In_623,In_99);
nand U1447 (N_1447,In_887,In_707);
nand U1448 (N_1448,In_323,N_948);
and U1449 (N_1449,In_1435,N_902);
nor U1450 (N_1450,N_992,In_102);
xor U1451 (N_1451,In_1782,N_664);
or U1452 (N_1452,In_378,N_469);
nand U1453 (N_1453,N_318,In_1749);
and U1454 (N_1454,N_351,N_160);
nor U1455 (N_1455,In_1349,N_195);
nor U1456 (N_1456,N_978,In_1046);
or U1457 (N_1457,In_1972,N_600);
nand U1458 (N_1458,N_939,In_633);
nor U1459 (N_1459,N_673,In_1058);
and U1460 (N_1460,In_426,N_585);
and U1461 (N_1461,In_1528,N_124);
nor U1462 (N_1462,N_644,In_1436);
nor U1463 (N_1463,N_533,In_957);
nand U1464 (N_1464,N_540,N_75);
or U1465 (N_1465,N_230,In_611);
or U1466 (N_1466,N_809,N_390);
nand U1467 (N_1467,N_552,N_866);
xnor U1468 (N_1468,N_798,N_596);
and U1469 (N_1469,N_59,In_1944);
nor U1470 (N_1470,N_892,N_996);
xor U1471 (N_1471,In_1710,In_1439);
and U1472 (N_1472,In_275,In_1707);
nor U1473 (N_1473,N_528,N_849);
or U1474 (N_1474,N_103,N_365);
nand U1475 (N_1475,N_876,In_857);
xnor U1476 (N_1476,In_1977,N_963);
nand U1477 (N_1477,N_589,N_867);
nand U1478 (N_1478,N_576,In_621);
and U1479 (N_1479,N_584,N_693);
nand U1480 (N_1480,N_951,N_882);
or U1481 (N_1481,N_838,N_910);
nand U1482 (N_1482,N_899,In_1166);
and U1483 (N_1483,N_434,N_569);
and U1484 (N_1484,In_1669,N_455);
and U1485 (N_1485,N_654,N_686);
and U1486 (N_1486,In_893,N_778);
and U1487 (N_1487,In_1144,N_707);
nand U1488 (N_1488,In_1458,N_969);
nand U1489 (N_1489,N_850,N_703);
nor U1490 (N_1490,N_376,In_1467);
or U1491 (N_1491,In_1808,N_962);
xor U1492 (N_1492,N_545,N_718);
xor U1493 (N_1493,N_220,N_949);
nor U1494 (N_1494,In_1761,N_909);
nand U1495 (N_1495,In_978,N_424);
xor U1496 (N_1496,In_670,N_471);
or U1497 (N_1497,In_1509,N_887);
or U1498 (N_1498,In_561,N_749);
and U1499 (N_1499,N_611,N_787);
nor U1500 (N_1500,N_1437,N_1496);
or U1501 (N_1501,N_1036,N_1206);
and U1502 (N_1502,N_1458,N_1377);
nand U1503 (N_1503,N_1100,N_1389);
and U1504 (N_1504,N_1204,N_1148);
or U1505 (N_1505,N_1007,N_1258);
nand U1506 (N_1506,N_1121,N_1275);
or U1507 (N_1507,N_1215,N_1338);
nand U1508 (N_1508,N_1308,N_1305);
and U1509 (N_1509,N_1037,N_1281);
or U1510 (N_1510,N_1440,N_1114);
nor U1511 (N_1511,N_1091,N_1015);
nor U1512 (N_1512,N_1196,N_1236);
xor U1513 (N_1513,N_1263,N_1311);
nor U1514 (N_1514,N_1240,N_1133);
nand U1515 (N_1515,N_1097,N_1428);
and U1516 (N_1516,N_1270,N_1390);
nand U1517 (N_1517,N_1083,N_1464);
or U1518 (N_1518,N_1029,N_1071);
or U1519 (N_1519,N_1024,N_1408);
nand U1520 (N_1520,N_1156,N_1465);
nor U1521 (N_1521,N_1213,N_1127);
nor U1522 (N_1522,N_1191,N_1339);
and U1523 (N_1523,N_1495,N_1126);
nor U1524 (N_1524,N_1313,N_1144);
xnor U1525 (N_1525,N_1084,N_1259);
nand U1526 (N_1526,N_1216,N_1486);
nand U1527 (N_1527,N_1019,N_1177);
and U1528 (N_1528,N_1287,N_1406);
xnor U1529 (N_1529,N_1260,N_1005);
and U1530 (N_1530,N_1488,N_1183);
xnor U1531 (N_1531,N_1018,N_1143);
and U1532 (N_1532,N_1055,N_1025);
nand U1533 (N_1533,N_1374,N_1310);
nand U1534 (N_1534,N_1164,N_1209);
nand U1535 (N_1535,N_1052,N_1239);
or U1536 (N_1536,N_1494,N_1237);
nor U1537 (N_1537,N_1448,N_1343);
or U1538 (N_1538,N_1132,N_1423);
or U1539 (N_1539,N_1013,N_1011);
or U1540 (N_1540,N_1393,N_1466);
and U1541 (N_1541,N_1452,N_1009);
and U1542 (N_1542,N_1131,N_1353);
or U1543 (N_1543,N_1101,N_1093);
xnor U1544 (N_1544,N_1075,N_1397);
xnor U1545 (N_1545,N_1090,N_1199);
xor U1546 (N_1546,N_1219,N_1170);
or U1547 (N_1547,N_1264,N_1290);
or U1548 (N_1548,N_1327,N_1003);
nand U1549 (N_1549,N_1181,N_1016);
nor U1550 (N_1550,N_1252,N_1441);
and U1551 (N_1551,N_1340,N_1032);
nor U1552 (N_1552,N_1140,N_1421);
xor U1553 (N_1553,N_1360,N_1073);
xnor U1554 (N_1554,N_1256,N_1438);
xnor U1555 (N_1555,N_1253,N_1443);
nor U1556 (N_1556,N_1254,N_1155);
or U1557 (N_1557,N_1372,N_1094);
and U1558 (N_1558,N_1371,N_1321);
nand U1559 (N_1559,N_1493,N_1300);
nor U1560 (N_1560,N_1195,N_1161);
nor U1561 (N_1561,N_1328,N_1033);
or U1562 (N_1562,N_1298,N_1113);
nand U1563 (N_1563,N_1008,N_1173);
nand U1564 (N_1564,N_1370,N_1030);
nand U1565 (N_1565,N_1230,N_1307);
nand U1566 (N_1566,N_1192,N_1415);
nand U1567 (N_1567,N_1401,N_1068);
or U1568 (N_1568,N_1431,N_1469);
xor U1569 (N_1569,N_1391,N_1381);
or U1570 (N_1570,N_1282,N_1346);
xnor U1571 (N_1571,N_1329,N_1444);
nand U1572 (N_1572,N_1320,N_1233);
or U1573 (N_1573,N_1153,N_1373);
xnor U1574 (N_1574,N_1169,N_1108);
and U1575 (N_1575,N_1442,N_1330);
xnor U1576 (N_1576,N_1026,N_1424);
and U1577 (N_1577,N_1242,N_1301);
nand U1578 (N_1578,N_1061,N_1483);
xnor U1579 (N_1579,N_1355,N_1398);
nand U1580 (N_1580,N_1194,N_1349);
or U1581 (N_1581,N_1103,N_1080);
or U1582 (N_1582,N_1277,N_1366);
nand U1583 (N_1583,N_1064,N_1269);
xor U1584 (N_1584,N_1189,N_1210);
nor U1585 (N_1585,N_1102,N_1250);
xnor U1586 (N_1586,N_1375,N_1010);
and U1587 (N_1587,N_1367,N_1413);
and U1588 (N_1588,N_1070,N_1382);
nand U1589 (N_1589,N_1356,N_1337);
xnor U1590 (N_1590,N_1481,N_1165);
and U1591 (N_1591,N_1176,N_1089);
nand U1592 (N_1592,N_1067,N_1455);
nand U1593 (N_1593,N_1409,N_1333);
nor U1594 (N_1594,N_1014,N_1081);
nor U1595 (N_1595,N_1106,N_1490);
nor U1596 (N_1596,N_1023,N_1386);
nor U1597 (N_1597,N_1359,N_1352);
nor U1598 (N_1598,N_1396,N_1418);
nor U1599 (N_1599,N_1474,N_1150);
xor U1600 (N_1600,N_1147,N_1178);
nor U1601 (N_1601,N_1420,N_1416);
and U1602 (N_1602,N_1109,N_1472);
xnor U1603 (N_1603,N_1066,N_1475);
xor U1604 (N_1604,N_1317,N_1280);
and U1605 (N_1605,N_1208,N_1456);
nor U1606 (N_1606,N_1085,N_1268);
xnor U1607 (N_1607,N_1119,N_1471);
nand U1608 (N_1608,N_1395,N_1491);
xnor U1609 (N_1609,N_1202,N_1358);
xnor U1610 (N_1610,N_1246,N_1146);
nor U1611 (N_1611,N_1099,N_1046);
xor U1612 (N_1612,N_1405,N_1043);
nand U1613 (N_1613,N_1244,N_1225);
nor U1614 (N_1614,N_1168,N_1412);
and U1615 (N_1615,N_1453,N_1040);
and U1616 (N_1616,N_1257,N_1478);
or U1617 (N_1617,N_1378,N_1457);
nor U1618 (N_1618,N_1086,N_1198);
and U1619 (N_1619,N_1088,N_1283);
and U1620 (N_1620,N_1384,N_1432);
and U1621 (N_1621,N_1053,N_1439);
and U1622 (N_1622,N_1492,N_1187);
or U1623 (N_1623,N_1312,N_1057);
nand U1624 (N_1624,N_1115,N_1163);
and U1625 (N_1625,N_1228,N_1351);
or U1626 (N_1626,N_1429,N_1303);
or U1627 (N_1627,N_1309,N_1104);
and U1628 (N_1628,N_1231,N_1159);
nor U1629 (N_1629,N_1188,N_1141);
nor U1630 (N_1630,N_1235,N_1142);
or U1631 (N_1631,N_1223,N_1262);
or U1632 (N_1632,N_1482,N_1368);
and U1633 (N_1633,N_1266,N_1069);
or U1634 (N_1634,N_1054,N_1123);
nor U1635 (N_1635,N_1294,N_1417);
or U1636 (N_1636,N_1020,N_1274);
or U1637 (N_1637,N_1332,N_1051);
nand U1638 (N_1638,N_1357,N_1145);
nand U1639 (N_1639,N_1049,N_1179);
nor U1640 (N_1640,N_1203,N_1473);
or U1641 (N_1641,N_1468,N_1182);
nor U1642 (N_1642,N_1082,N_1403);
or U1643 (N_1643,N_1092,N_1460);
nand U1644 (N_1644,N_1407,N_1385);
nor U1645 (N_1645,N_1222,N_1136);
nand U1646 (N_1646,N_1433,N_1434);
and U1647 (N_1647,N_1285,N_1076);
xor U1648 (N_1648,N_1447,N_1134);
nand U1649 (N_1649,N_1463,N_1489);
nand U1650 (N_1650,N_1435,N_1487);
nor U1651 (N_1651,N_1111,N_1427);
nor U1652 (N_1652,N_1324,N_1251);
nor U1653 (N_1653,N_1291,N_1331);
xor U1654 (N_1654,N_1039,N_1002);
and U1655 (N_1655,N_1342,N_1289);
xnor U1656 (N_1656,N_1034,N_1379);
and U1657 (N_1657,N_1214,N_1380);
nand U1658 (N_1658,N_1001,N_1157);
nor U1659 (N_1659,N_1265,N_1387);
and U1660 (N_1660,N_1217,N_1334);
xor U1661 (N_1661,N_1392,N_1035);
xnor U1662 (N_1662,N_1234,N_1363);
and U1663 (N_1663,N_1162,N_1446);
and U1664 (N_1664,N_1063,N_1220);
or U1665 (N_1665,N_1062,N_1158);
or U1666 (N_1666,N_1326,N_1038);
nand U1667 (N_1667,N_1430,N_1139);
nand U1668 (N_1668,N_1449,N_1243);
or U1669 (N_1669,N_1175,N_1295);
nor U1670 (N_1670,N_1369,N_1459);
nand U1671 (N_1671,N_1314,N_1167);
or U1672 (N_1672,N_1364,N_1171);
xor U1673 (N_1673,N_1484,N_1462);
nor U1674 (N_1674,N_1044,N_1322);
nand U1675 (N_1675,N_1226,N_1318);
nor U1676 (N_1676,N_1273,N_1004);
nand U1677 (N_1677,N_1047,N_1229);
nor U1678 (N_1678,N_1212,N_1184);
and U1679 (N_1679,N_1293,N_1344);
nor U1680 (N_1680,N_1031,N_1261);
or U1681 (N_1681,N_1211,N_1404);
or U1682 (N_1682,N_1249,N_1152);
xor U1683 (N_1683,N_1479,N_1095);
xnor U1684 (N_1684,N_1028,N_1297);
and U1685 (N_1685,N_1477,N_1302);
and U1686 (N_1686,N_1027,N_1135);
nor U1687 (N_1687,N_1323,N_1450);
or U1688 (N_1688,N_1410,N_1299);
xnor U1689 (N_1689,N_1096,N_1050);
and U1690 (N_1690,N_1445,N_1006);
or U1691 (N_1691,N_1247,N_1306);
or U1692 (N_1692,N_1098,N_1394);
nor U1693 (N_1693,N_1454,N_1154);
xnor U1694 (N_1694,N_1172,N_1335);
and U1695 (N_1695,N_1315,N_1400);
or U1696 (N_1696,N_1078,N_1436);
nor U1697 (N_1697,N_1174,N_1221);
nand U1698 (N_1698,N_1151,N_1079);
nor U1699 (N_1699,N_1354,N_1185);
or U1700 (N_1700,N_1218,N_1124);
or U1701 (N_1701,N_1021,N_1497);
or U1702 (N_1702,N_1227,N_1402);
nor U1703 (N_1703,N_1341,N_1325);
xor U1704 (N_1704,N_1267,N_1205);
xor U1705 (N_1705,N_1319,N_1058);
and U1706 (N_1706,N_1348,N_1045);
xor U1707 (N_1707,N_1012,N_1110);
nand U1708 (N_1708,N_1105,N_1350);
nand U1709 (N_1709,N_1074,N_1248);
xnor U1710 (N_1710,N_1180,N_1383);
xnor U1711 (N_1711,N_1480,N_1365);
and U1712 (N_1712,N_1336,N_1042);
nor U1713 (N_1713,N_1232,N_1041);
or U1714 (N_1714,N_1426,N_1361);
nor U1715 (N_1715,N_1276,N_1166);
and U1716 (N_1716,N_1138,N_1451);
and U1717 (N_1717,N_1316,N_1065);
and U1718 (N_1718,N_1160,N_1238);
or U1719 (N_1719,N_1255,N_1304);
and U1720 (N_1720,N_1284,N_1499);
xnor U1721 (N_1721,N_1129,N_1241);
nor U1722 (N_1722,N_1059,N_1118);
nor U1723 (N_1723,N_1286,N_1122);
xnor U1724 (N_1724,N_1422,N_1117);
nor U1725 (N_1725,N_1072,N_1467);
or U1726 (N_1726,N_1087,N_1470);
nand U1727 (N_1727,N_1278,N_1279);
and U1728 (N_1728,N_1272,N_1120);
xnor U1729 (N_1729,N_1461,N_1388);
or U1730 (N_1730,N_1137,N_1190);
xnor U1731 (N_1731,N_1498,N_1207);
nand U1732 (N_1732,N_1077,N_1200);
nand U1733 (N_1733,N_1125,N_1476);
or U1734 (N_1734,N_1271,N_1414);
xor U1735 (N_1735,N_1296,N_1347);
nand U1736 (N_1736,N_1000,N_1022);
xnor U1737 (N_1737,N_1411,N_1197);
or U1738 (N_1738,N_1345,N_1376);
nor U1739 (N_1739,N_1186,N_1017);
or U1740 (N_1740,N_1116,N_1048);
nand U1741 (N_1741,N_1288,N_1130);
nor U1742 (N_1742,N_1485,N_1193);
and U1743 (N_1743,N_1245,N_1128);
or U1744 (N_1744,N_1362,N_1060);
nor U1745 (N_1745,N_1224,N_1056);
and U1746 (N_1746,N_1112,N_1201);
xor U1747 (N_1747,N_1292,N_1419);
nand U1748 (N_1748,N_1425,N_1107);
xnor U1749 (N_1749,N_1149,N_1399);
nand U1750 (N_1750,N_1029,N_1086);
xor U1751 (N_1751,N_1286,N_1480);
or U1752 (N_1752,N_1227,N_1029);
nor U1753 (N_1753,N_1121,N_1134);
or U1754 (N_1754,N_1045,N_1174);
or U1755 (N_1755,N_1495,N_1032);
nand U1756 (N_1756,N_1445,N_1399);
and U1757 (N_1757,N_1422,N_1002);
nand U1758 (N_1758,N_1066,N_1496);
and U1759 (N_1759,N_1228,N_1365);
nand U1760 (N_1760,N_1468,N_1216);
nand U1761 (N_1761,N_1239,N_1389);
xnor U1762 (N_1762,N_1241,N_1392);
nor U1763 (N_1763,N_1269,N_1344);
and U1764 (N_1764,N_1126,N_1101);
xor U1765 (N_1765,N_1116,N_1235);
and U1766 (N_1766,N_1106,N_1129);
nor U1767 (N_1767,N_1024,N_1003);
or U1768 (N_1768,N_1212,N_1078);
nand U1769 (N_1769,N_1367,N_1432);
nor U1770 (N_1770,N_1388,N_1474);
nor U1771 (N_1771,N_1123,N_1338);
or U1772 (N_1772,N_1080,N_1481);
and U1773 (N_1773,N_1335,N_1398);
and U1774 (N_1774,N_1207,N_1495);
and U1775 (N_1775,N_1456,N_1486);
or U1776 (N_1776,N_1024,N_1224);
and U1777 (N_1777,N_1280,N_1366);
nand U1778 (N_1778,N_1277,N_1302);
or U1779 (N_1779,N_1270,N_1052);
nand U1780 (N_1780,N_1286,N_1430);
xnor U1781 (N_1781,N_1063,N_1378);
nand U1782 (N_1782,N_1472,N_1490);
and U1783 (N_1783,N_1479,N_1351);
nand U1784 (N_1784,N_1047,N_1084);
nand U1785 (N_1785,N_1264,N_1144);
nand U1786 (N_1786,N_1476,N_1042);
or U1787 (N_1787,N_1429,N_1467);
and U1788 (N_1788,N_1019,N_1499);
or U1789 (N_1789,N_1350,N_1404);
nor U1790 (N_1790,N_1021,N_1391);
and U1791 (N_1791,N_1015,N_1165);
and U1792 (N_1792,N_1130,N_1080);
nand U1793 (N_1793,N_1429,N_1127);
nor U1794 (N_1794,N_1382,N_1061);
xor U1795 (N_1795,N_1080,N_1040);
xnor U1796 (N_1796,N_1152,N_1138);
xnor U1797 (N_1797,N_1087,N_1267);
nand U1798 (N_1798,N_1012,N_1447);
or U1799 (N_1799,N_1339,N_1093);
xor U1800 (N_1800,N_1193,N_1116);
or U1801 (N_1801,N_1173,N_1432);
nor U1802 (N_1802,N_1164,N_1376);
and U1803 (N_1803,N_1152,N_1253);
nor U1804 (N_1804,N_1422,N_1436);
or U1805 (N_1805,N_1238,N_1032);
xor U1806 (N_1806,N_1081,N_1290);
nand U1807 (N_1807,N_1381,N_1372);
or U1808 (N_1808,N_1374,N_1154);
and U1809 (N_1809,N_1170,N_1074);
and U1810 (N_1810,N_1198,N_1106);
or U1811 (N_1811,N_1053,N_1321);
and U1812 (N_1812,N_1192,N_1446);
and U1813 (N_1813,N_1358,N_1448);
or U1814 (N_1814,N_1349,N_1386);
or U1815 (N_1815,N_1064,N_1132);
or U1816 (N_1816,N_1221,N_1423);
and U1817 (N_1817,N_1099,N_1110);
and U1818 (N_1818,N_1212,N_1196);
and U1819 (N_1819,N_1109,N_1447);
nor U1820 (N_1820,N_1060,N_1023);
and U1821 (N_1821,N_1054,N_1458);
nor U1822 (N_1822,N_1098,N_1489);
nor U1823 (N_1823,N_1007,N_1289);
xnor U1824 (N_1824,N_1033,N_1096);
nand U1825 (N_1825,N_1069,N_1221);
nand U1826 (N_1826,N_1129,N_1310);
or U1827 (N_1827,N_1136,N_1104);
and U1828 (N_1828,N_1347,N_1196);
or U1829 (N_1829,N_1082,N_1349);
xor U1830 (N_1830,N_1418,N_1241);
or U1831 (N_1831,N_1290,N_1478);
and U1832 (N_1832,N_1232,N_1384);
nor U1833 (N_1833,N_1269,N_1067);
and U1834 (N_1834,N_1237,N_1362);
nor U1835 (N_1835,N_1363,N_1401);
nand U1836 (N_1836,N_1432,N_1182);
and U1837 (N_1837,N_1326,N_1390);
xnor U1838 (N_1838,N_1389,N_1155);
or U1839 (N_1839,N_1419,N_1114);
nor U1840 (N_1840,N_1029,N_1464);
nor U1841 (N_1841,N_1132,N_1282);
nand U1842 (N_1842,N_1336,N_1088);
and U1843 (N_1843,N_1442,N_1376);
or U1844 (N_1844,N_1074,N_1037);
or U1845 (N_1845,N_1072,N_1395);
or U1846 (N_1846,N_1426,N_1244);
or U1847 (N_1847,N_1329,N_1037);
xor U1848 (N_1848,N_1223,N_1065);
nand U1849 (N_1849,N_1357,N_1117);
nor U1850 (N_1850,N_1440,N_1041);
and U1851 (N_1851,N_1007,N_1090);
nor U1852 (N_1852,N_1274,N_1277);
nand U1853 (N_1853,N_1490,N_1298);
nand U1854 (N_1854,N_1118,N_1297);
or U1855 (N_1855,N_1378,N_1118);
nor U1856 (N_1856,N_1233,N_1436);
and U1857 (N_1857,N_1465,N_1110);
nand U1858 (N_1858,N_1170,N_1089);
and U1859 (N_1859,N_1218,N_1248);
nor U1860 (N_1860,N_1467,N_1289);
xnor U1861 (N_1861,N_1026,N_1440);
or U1862 (N_1862,N_1285,N_1455);
xnor U1863 (N_1863,N_1257,N_1189);
nand U1864 (N_1864,N_1079,N_1386);
xor U1865 (N_1865,N_1179,N_1183);
and U1866 (N_1866,N_1303,N_1398);
nand U1867 (N_1867,N_1420,N_1188);
or U1868 (N_1868,N_1328,N_1179);
xor U1869 (N_1869,N_1335,N_1348);
or U1870 (N_1870,N_1131,N_1396);
and U1871 (N_1871,N_1120,N_1012);
and U1872 (N_1872,N_1247,N_1442);
or U1873 (N_1873,N_1075,N_1280);
nor U1874 (N_1874,N_1449,N_1204);
and U1875 (N_1875,N_1035,N_1150);
xor U1876 (N_1876,N_1050,N_1352);
or U1877 (N_1877,N_1345,N_1486);
nor U1878 (N_1878,N_1037,N_1298);
and U1879 (N_1879,N_1115,N_1202);
or U1880 (N_1880,N_1499,N_1052);
xor U1881 (N_1881,N_1112,N_1088);
and U1882 (N_1882,N_1074,N_1254);
or U1883 (N_1883,N_1205,N_1284);
or U1884 (N_1884,N_1076,N_1249);
and U1885 (N_1885,N_1143,N_1292);
or U1886 (N_1886,N_1457,N_1334);
xnor U1887 (N_1887,N_1440,N_1363);
and U1888 (N_1888,N_1100,N_1385);
and U1889 (N_1889,N_1432,N_1215);
xnor U1890 (N_1890,N_1300,N_1156);
nand U1891 (N_1891,N_1491,N_1307);
nor U1892 (N_1892,N_1419,N_1232);
nand U1893 (N_1893,N_1401,N_1427);
nor U1894 (N_1894,N_1333,N_1299);
xnor U1895 (N_1895,N_1386,N_1149);
and U1896 (N_1896,N_1271,N_1418);
or U1897 (N_1897,N_1262,N_1098);
xnor U1898 (N_1898,N_1065,N_1442);
nor U1899 (N_1899,N_1430,N_1002);
and U1900 (N_1900,N_1021,N_1181);
nor U1901 (N_1901,N_1165,N_1074);
nor U1902 (N_1902,N_1440,N_1491);
or U1903 (N_1903,N_1007,N_1059);
nand U1904 (N_1904,N_1421,N_1253);
and U1905 (N_1905,N_1144,N_1166);
nand U1906 (N_1906,N_1226,N_1372);
nor U1907 (N_1907,N_1492,N_1419);
nand U1908 (N_1908,N_1391,N_1025);
nand U1909 (N_1909,N_1129,N_1059);
xnor U1910 (N_1910,N_1280,N_1231);
nand U1911 (N_1911,N_1096,N_1426);
nor U1912 (N_1912,N_1486,N_1252);
xor U1913 (N_1913,N_1368,N_1481);
nand U1914 (N_1914,N_1172,N_1468);
and U1915 (N_1915,N_1240,N_1293);
xor U1916 (N_1916,N_1156,N_1431);
or U1917 (N_1917,N_1100,N_1091);
and U1918 (N_1918,N_1315,N_1471);
nor U1919 (N_1919,N_1172,N_1074);
and U1920 (N_1920,N_1007,N_1390);
nand U1921 (N_1921,N_1070,N_1408);
or U1922 (N_1922,N_1313,N_1307);
xor U1923 (N_1923,N_1450,N_1404);
nand U1924 (N_1924,N_1124,N_1060);
nand U1925 (N_1925,N_1096,N_1456);
nand U1926 (N_1926,N_1321,N_1445);
xor U1927 (N_1927,N_1067,N_1200);
xor U1928 (N_1928,N_1359,N_1271);
xor U1929 (N_1929,N_1286,N_1426);
nand U1930 (N_1930,N_1089,N_1432);
nor U1931 (N_1931,N_1269,N_1235);
and U1932 (N_1932,N_1067,N_1466);
xnor U1933 (N_1933,N_1202,N_1310);
nand U1934 (N_1934,N_1396,N_1282);
and U1935 (N_1935,N_1004,N_1354);
or U1936 (N_1936,N_1173,N_1284);
nand U1937 (N_1937,N_1390,N_1275);
or U1938 (N_1938,N_1371,N_1393);
nand U1939 (N_1939,N_1385,N_1436);
or U1940 (N_1940,N_1198,N_1010);
nand U1941 (N_1941,N_1446,N_1306);
xnor U1942 (N_1942,N_1261,N_1386);
nand U1943 (N_1943,N_1269,N_1246);
xor U1944 (N_1944,N_1044,N_1212);
nand U1945 (N_1945,N_1163,N_1370);
nand U1946 (N_1946,N_1253,N_1326);
nand U1947 (N_1947,N_1399,N_1092);
nand U1948 (N_1948,N_1018,N_1264);
or U1949 (N_1949,N_1428,N_1217);
nand U1950 (N_1950,N_1185,N_1086);
nor U1951 (N_1951,N_1063,N_1432);
nand U1952 (N_1952,N_1041,N_1478);
nand U1953 (N_1953,N_1308,N_1409);
or U1954 (N_1954,N_1457,N_1055);
nand U1955 (N_1955,N_1276,N_1021);
nor U1956 (N_1956,N_1361,N_1372);
nor U1957 (N_1957,N_1486,N_1093);
nand U1958 (N_1958,N_1292,N_1393);
nand U1959 (N_1959,N_1021,N_1265);
or U1960 (N_1960,N_1448,N_1415);
or U1961 (N_1961,N_1183,N_1207);
xnor U1962 (N_1962,N_1098,N_1371);
and U1963 (N_1963,N_1146,N_1274);
nor U1964 (N_1964,N_1131,N_1292);
nor U1965 (N_1965,N_1154,N_1150);
or U1966 (N_1966,N_1005,N_1338);
or U1967 (N_1967,N_1178,N_1402);
nand U1968 (N_1968,N_1426,N_1391);
and U1969 (N_1969,N_1321,N_1062);
nand U1970 (N_1970,N_1198,N_1075);
nor U1971 (N_1971,N_1087,N_1393);
and U1972 (N_1972,N_1467,N_1113);
nor U1973 (N_1973,N_1246,N_1334);
or U1974 (N_1974,N_1282,N_1340);
nor U1975 (N_1975,N_1394,N_1074);
xor U1976 (N_1976,N_1184,N_1233);
nand U1977 (N_1977,N_1420,N_1297);
nand U1978 (N_1978,N_1350,N_1358);
nand U1979 (N_1979,N_1321,N_1452);
nor U1980 (N_1980,N_1408,N_1206);
and U1981 (N_1981,N_1180,N_1171);
nor U1982 (N_1982,N_1388,N_1203);
nor U1983 (N_1983,N_1136,N_1436);
or U1984 (N_1984,N_1073,N_1029);
xnor U1985 (N_1985,N_1257,N_1008);
nor U1986 (N_1986,N_1392,N_1157);
xnor U1987 (N_1987,N_1135,N_1383);
and U1988 (N_1988,N_1111,N_1188);
nand U1989 (N_1989,N_1185,N_1317);
nand U1990 (N_1990,N_1183,N_1023);
or U1991 (N_1991,N_1384,N_1311);
or U1992 (N_1992,N_1376,N_1411);
nor U1993 (N_1993,N_1006,N_1416);
nand U1994 (N_1994,N_1384,N_1067);
xor U1995 (N_1995,N_1411,N_1059);
and U1996 (N_1996,N_1245,N_1378);
xor U1997 (N_1997,N_1456,N_1011);
xnor U1998 (N_1998,N_1422,N_1418);
or U1999 (N_1999,N_1484,N_1306);
and U2000 (N_2000,N_1703,N_1779);
xnor U2001 (N_2001,N_1933,N_1626);
nor U2002 (N_2002,N_1745,N_1609);
nor U2003 (N_2003,N_1602,N_1675);
xnor U2004 (N_2004,N_1606,N_1920);
xor U2005 (N_2005,N_1564,N_1708);
or U2006 (N_2006,N_1665,N_1692);
nand U2007 (N_2007,N_1818,N_1760);
xor U2008 (N_2008,N_1529,N_1746);
nor U2009 (N_2009,N_1770,N_1991);
and U2010 (N_2010,N_1721,N_1573);
or U2011 (N_2011,N_1637,N_1852);
and U2012 (N_2012,N_1872,N_1542);
or U2013 (N_2013,N_1955,N_1739);
or U2014 (N_2014,N_1887,N_1571);
or U2015 (N_2015,N_1572,N_1923);
and U2016 (N_2016,N_1695,N_1783);
nor U2017 (N_2017,N_1881,N_1617);
xnor U2018 (N_2018,N_1752,N_1592);
xnor U2019 (N_2019,N_1577,N_1851);
xnor U2020 (N_2020,N_1987,N_1913);
xor U2021 (N_2021,N_1669,N_1605);
nand U2022 (N_2022,N_1788,N_1869);
xnor U2023 (N_2023,N_1828,N_1724);
nor U2024 (N_2024,N_1927,N_1984);
and U2025 (N_2025,N_1641,N_1960);
nor U2026 (N_2026,N_1799,N_1751);
or U2027 (N_2027,N_1849,N_1627);
or U2028 (N_2028,N_1514,N_1956);
nand U2029 (N_2029,N_1599,N_1722);
or U2030 (N_2030,N_1657,N_1836);
nand U2031 (N_2031,N_1509,N_1890);
nor U2032 (N_2032,N_1670,N_1524);
xor U2033 (N_2033,N_1750,N_1638);
nand U2034 (N_2034,N_1698,N_1504);
and U2035 (N_2035,N_1996,N_1723);
xor U2036 (N_2036,N_1846,N_1541);
xnor U2037 (N_2037,N_1674,N_1747);
nor U2038 (N_2038,N_1965,N_1676);
xnor U2039 (N_2039,N_1531,N_1903);
or U2040 (N_2040,N_1550,N_1651);
nor U2041 (N_2041,N_1500,N_1748);
xor U2042 (N_2042,N_1953,N_1850);
and U2043 (N_2043,N_1888,N_1644);
and U2044 (N_2044,N_1696,N_1734);
and U2045 (N_2045,N_1757,N_1900);
and U2046 (N_2046,N_1697,N_1883);
nor U2047 (N_2047,N_1772,N_1523);
nor U2048 (N_2048,N_1587,N_1691);
nand U2049 (N_2049,N_1507,N_1689);
xnor U2050 (N_2050,N_1798,N_1568);
nor U2051 (N_2051,N_1875,N_1969);
nand U2052 (N_2052,N_1536,N_1777);
or U2053 (N_2053,N_1904,N_1865);
nand U2054 (N_2054,N_1966,N_1906);
or U2055 (N_2055,N_1639,N_1655);
nor U2056 (N_2056,N_1807,N_1744);
nor U2057 (N_2057,N_1824,N_1800);
nor U2058 (N_2058,N_1805,N_1552);
xor U2059 (N_2059,N_1539,N_1905);
or U2060 (N_2060,N_1738,N_1535);
nand U2061 (N_2061,N_1650,N_1700);
xnor U2062 (N_2062,N_1827,N_1837);
or U2063 (N_2063,N_1997,N_1974);
nand U2064 (N_2064,N_1726,N_1516);
or U2065 (N_2065,N_1988,N_1601);
nor U2066 (N_2066,N_1716,N_1947);
xnor U2067 (N_2067,N_1634,N_1753);
nor U2068 (N_2068,N_1928,N_1505);
nand U2069 (N_2069,N_1917,N_1860);
or U2070 (N_2070,N_1645,N_1719);
xnor U2071 (N_2071,N_1709,N_1635);
nor U2072 (N_2072,N_1527,N_1553);
or U2073 (N_2073,N_1858,N_1512);
and U2074 (N_2074,N_1999,N_1876);
nand U2075 (N_2075,N_1714,N_1658);
xnor U2076 (N_2076,N_1802,N_1902);
nand U2077 (N_2077,N_1936,N_1791);
nand U2078 (N_2078,N_1793,N_1604);
or U2079 (N_2079,N_1831,N_1593);
or U2080 (N_2080,N_1702,N_1688);
or U2081 (N_2081,N_1782,N_1896);
nand U2082 (N_2082,N_1582,N_1652);
xor U2083 (N_2083,N_1768,N_1502);
nor U2084 (N_2084,N_1813,N_1742);
and U2085 (N_2085,N_1855,N_1707);
and U2086 (N_2086,N_1518,N_1563);
nand U2087 (N_2087,N_1659,N_1623);
xor U2088 (N_2088,N_1642,N_1620);
xnor U2089 (N_2089,N_1909,N_1621);
nand U2090 (N_2090,N_1961,N_1771);
and U2091 (N_2091,N_1545,N_1957);
or U2092 (N_2092,N_1986,N_1784);
and U2093 (N_2093,N_1806,N_1671);
nand U2094 (N_2094,N_1559,N_1517);
nor U2095 (N_2095,N_1832,N_1546);
xnor U2096 (N_2096,N_1977,N_1954);
nand U2097 (N_2097,N_1787,N_1854);
or U2098 (N_2098,N_1715,N_1610);
nor U2099 (N_2099,N_1893,N_1501);
or U2100 (N_2100,N_1942,N_1841);
nor U2101 (N_2101,N_1581,N_1543);
nand U2102 (N_2102,N_1725,N_1838);
nor U2103 (N_2103,N_1950,N_1861);
and U2104 (N_2104,N_1801,N_1873);
nand U2105 (N_2105,N_1878,N_1548);
nor U2106 (N_2106,N_1976,N_1882);
nand U2107 (N_2107,N_1911,N_1561);
nor U2108 (N_2108,N_1737,N_1754);
nand U2109 (N_2109,N_1576,N_1557);
xnor U2110 (N_2110,N_1778,N_1534);
nor U2111 (N_2111,N_1661,N_1835);
or U2112 (N_2112,N_1975,N_1774);
xnor U2113 (N_2113,N_1503,N_1560);
and U2114 (N_2114,N_1990,N_1985);
nor U2115 (N_2115,N_1677,N_1736);
or U2116 (N_2116,N_1590,N_1720);
nand U2117 (N_2117,N_1575,N_1622);
and U2118 (N_2118,N_1515,N_1919);
or U2119 (N_2119,N_1845,N_1643);
xnor U2120 (N_2120,N_1664,N_1585);
nor U2121 (N_2121,N_1992,N_1810);
nor U2122 (N_2122,N_1717,N_1843);
nand U2123 (N_2123,N_1816,N_1673);
nand U2124 (N_2124,N_1558,N_1863);
and U2125 (N_2125,N_1765,N_1764);
or U2126 (N_2126,N_1648,N_1769);
or U2127 (N_2127,N_1598,N_1815);
nand U2128 (N_2128,N_1857,N_1615);
xnor U2129 (N_2129,N_1756,N_1898);
or U2130 (N_2130,N_1944,N_1897);
nor U2131 (N_2131,N_1762,N_1660);
nand U2132 (N_2132,N_1781,N_1958);
nand U2133 (N_2133,N_1586,N_1684);
nand U2134 (N_2134,N_1629,N_1994);
nor U2135 (N_2135,N_1600,N_1856);
nor U2136 (N_2136,N_1993,N_1834);
nand U2137 (N_2137,N_1759,N_1740);
nand U2138 (N_2138,N_1755,N_1879);
and U2139 (N_2139,N_1767,N_1662);
xor U2140 (N_2140,N_1729,N_1711);
xor U2141 (N_2141,N_1780,N_1825);
nand U2142 (N_2142,N_1940,N_1580);
or U2143 (N_2143,N_1728,N_1654);
or U2144 (N_2144,N_1538,N_1519);
nor U2145 (N_2145,N_1636,N_1595);
nand U2146 (N_2146,N_1973,N_1924);
nand U2147 (N_2147,N_1663,N_1926);
nor U2148 (N_2148,N_1792,N_1971);
nand U2149 (N_2149,N_1591,N_1667);
and U2150 (N_2150,N_1706,N_1693);
xor U2151 (N_2151,N_1916,N_1574);
and U2152 (N_2152,N_1946,N_1611);
nand U2153 (N_2153,N_1649,N_1628);
nor U2154 (N_2154,N_1797,N_1943);
nor U2155 (N_2155,N_1945,N_1565);
nand U2156 (N_2156,N_1690,N_1833);
and U2157 (N_2157,N_1533,N_1932);
xnor U2158 (N_2158,N_1980,N_1814);
nor U2159 (N_2159,N_1619,N_1867);
nand U2160 (N_2160,N_1795,N_1853);
or U2161 (N_2161,N_1579,N_1921);
or U2162 (N_2162,N_1597,N_1525);
or U2163 (N_2163,N_1699,N_1732);
and U2164 (N_2164,N_1683,N_1866);
nand U2165 (N_2165,N_1521,N_1907);
and U2166 (N_2166,N_1870,N_1511);
and U2167 (N_2167,N_1938,N_1889);
nand U2168 (N_2168,N_1613,N_1967);
or U2169 (N_2169,N_1998,N_1794);
and U2170 (N_2170,N_1914,N_1625);
xor U2171 (N_2171,N_1808,N_1868);
and U2172 (N_2172,N_1848,N_1951);
nor U2173 (N_2173,N_1761,N_1989);
nand U2174 (N_2174,N_1567,N_1970);
and U2175 (N_2175,N_1922,N_1821);
nand U2176 (N_2176,N_1891,N_1895);
or U2177 (N_2177,N_1981,N_1948);
nor U2178 (N_2178,N_1631,N_1962);
xnor U2179 (N_2179,N_1547,N_1822);
nor U2180 (N_2180,N_1679,N_1937);
or U2181 (N_2181,N_1830,N_1829);
nand U2182 (N_2182,N_1880,N_1812);
nand U2183 (N_2183,N_1862,N_1584);
nor U2184 (N_2184,N_1624,N_1847);
nand U2185 (N_2185,N_1508,N_1666);
nor U2186 (N_2186,N_1551,N_1978);
or U2187 (N_2187,N_1840,N_1710);
and U2188 (N_2188,N_1647,N_1859);
and U2189 (N_2189,N_1886,N_1968);
xnor U2190 (N_2190,N_1823,N_1885);
nor U2191 (N_2191,N_1930,N_1935);
nor U2192 (N_2192,N_1532,N_1963);
and U2193 (N_2193,N_1758,N_1730);
nor U2194 (N_2194,N_1520,N_1983);
xor U2195 (N_2195,N_1803,N_1939);
nor U2196 (N_2196,N_1570,N_1712);
and U2197 (N_2197,N_1653,N_1526);
nor U2198 (N_2198,N_1607,N_1894);
and U2199 (N_2199,N_1640,N_1809);
or U2200 (N_2200,N_1646,N_1632);
xnor U2201 (N_2201,N_1817,N_1934);
nor U2202 (N_2202,N_1733,N_1680);
and U2203 (N_2203,N_1510,N_1796);
xnor U2204 (N_2204,N_1773,N_1979);
or U2205 (N_2205,N_1931,N_1844);
nand U2206 (N_2206,N_1910,N_1952);
xor U2207 (N_2207,N_1589,N_1608);
and U2208 (N_2208,N_1704,N_1537);
and U2209 (N_2209,N_1735,N_1705);
xnor U2210 (N_2210,N_1915,N_1995);
xor U2211 (N_2211,N_1901,N_1618);
or U2212 (N_2212,N_1694,N_1776);
nand U2213 (N_2213,N_1826,N_1775);
nor U2214 (N_2214,N_1701,N_1682);
nand U2215 (N_2215,N_1596,N_1842);
nand U2216 (N_2216,N_1540,N_1630);
and U2217 (N_2217,N_1566,N_1763);
nand U2218 (N_2218,N_1982,N_1549);
nand U2219 (N_2219,N_1614,N_1672);
nor U2220 (N_2220,N_1633,N_1685);
nor U2221 (N_2221,N_1569,N_1941);
nand U2222 (N_2222,N_1949,N_1686);
nor U2223 (N_2223,N_1959,N_1713);
nand U2224 (N_2224,N_1743,N_1544);
nor U2225 (N_2225,N_1528,N_1656);
xnor U2226 (N_2226,N_1603,N_1877);
or U2227 (N_2227,N_1790,N_1731);
nor U2228 (N_2228,N_1554,N_1668);
nor U2229 (N_2229,N_1506,N_1804);
and U2230 (N_2230,N_1786,N_1749);
and U2231 (N_2231,N_1892,N_1874);
and U2232 (N_2232,N_1819,N_1718);
or U2233 (N_2233,N_1918,N_1964);
nor U2234 (N_2234,N_1530,N_1678);
and U2235 (N_2235,N_1583,N_1594);
and U2236 (N_2236,N_1899,N_1766);
nor U2237 (N_2237,N_1912,N_1871);
nor U2238 (N_2238,N_1612,N_1789);
nand U2239 (N_2239,N_1925,N_1556);
and U2240 (N_2240,N_1727,N_1588);
nand U2241 (N_2241,N_1522,N_1578);
nand U2242 (N_2242,N_1687,N_1864);
xor U2243 (N_2243,N_1741,N_1555);
xnor U2244 (N_2244,N_1562,N_1884);
and U2245 (N_2245,N_1908,N_1929);
nor U2246 (N_2246,N_1513,N_1839);
xnor U2247 (N_2247,N_1616,N_1820);
xor U2248 (N_2248,N_1811,N_1681);
xor U2249 (N_2249,N_1972,N_1785);
or U2250 (N_2250,N_1526,N_1736);
or U2251 (N_2251,N_1605,N_1702);
or U2252 (N_2252,N_1732,N_1987);
and U2253 (N_2253,N_1855,N_1964);
and U2254 (N_2254,N_1785,N_1960);
or U2255 (N_2255,N_1948,N_1943);
nor U2256 (N_2256,N_1527,N_1862);
and U2257 (N_2257,N_1536,N_1943);
nor U2258 (N_2258,N_1808,N_1703);
nand U2259 (N_2259,N_1562,N_1958);
nor U2260 (N_2260,N_1628,N_1508);
nor U2261 (N_2261,N_1927,N_1706);
nand U2262 (N_2262,N_1621,N_1517);
or U2263 (N_2263,N_1600,N_1562);
and U2264 (N_2264,N_1973,N_1661);
nand U2265 (N_2265,N_1847,N_1933);
nand U2266 (N_2266,N_1881,N_1522);
xor U2267 (N_2267,N_1593,N_1816);
xnor U2268 (N_2268,N_1923,N_1740);
nor U2269 (N_2269,N_1975,N_1557);
and U2270 (N_2270,N_1547,N_1742);
and U2271 (N_2271,N_1950,N_1520);
nor U2272 (N_2272,N_1875,N_1581);
and U2273 (N_2273,N_1502,N_1943);
nor U2274 (N_2274,N_1670,N_1616);
nand U2275 (N_2275,N_1563,N_1647);
and U2276 (N_2276,N_1933,N_1862);
xor U2277 (N_2277,N_1848,N_1544);
and U2278 (N_2278,N_1980,N_1913);
or U2279 (N_2279,N_1764,N_1509);
nand U2280 (N_2280,N_1597,N_1654);
nand U2281 (N_2281,N_1744,N_1543);
nand U2282 (N_2282,N_1601,N_1804);
xor U2283 (N_2283,N_1971,N_1516);
nand U2284 (N_2284,N_1661,N_1589);
and U2285 (N_2285,N_1645,N_1774);
nand U2286 (N_2286,N_1775,N_1847);
nand U2287 (N_2287,N_1643,N_1556);
nor U2288 (N_2288,N_1678,N_1872);
nand U2289 (N_2289,N_1792,N_1898);
and U2290 (N_2290,N_1680,N_1827);
xnor U2291 (N_2291,N_1860,N_1659);
or U2292 (N_2292,N_1949,N_1919);
or U2293 (N_2293,N_1536,N_1576);
or U2294 (N_2294,N_1626,N_1902);
or U2295 (N_2295,N_1714,N_1558);
xnor U2296 (N_2296,N_1815,N_1717);
xor U2297 (N_2297,N_1935,N_1826);
and U2298 (N_2298,N_1754,N_1620);
and U2299 (N_2299,N_1785,N_1708);
and U2300 (N_2300,N_1819,N_1991);
nand U2301 (N_2301,N_1981,N_1529);
nand U2302 (N_2302,N_1851,N_1595);
nor U2303 (N_2303,N_1811,N_1804);
xnor U2304 (N_2304,N_1564,N_1914);
or U2305 (N_2305,N_1614,N_1707);
and U2306 (N_2306,N_1639,N_1596);
or U2307 (N_2307,N_1558,N_1915);
nor U2308 (N_2308,N_1947,N_1724);
nor U2309 (N_2309,N_1763,N_1526);
and U2310 (N_2310,N_1614,N_1891);
or U2311 (N_2311,N_1573,N_1536);
nor U2312 (N_2312,N_1653,N_1520);
xor U2313 (N_2313,N_1651,N_1749);
and U2314 (N_2314,N_1780,N_1680);
nor U2315 (N_2315,N_1979,N_1598);
or U2316 (N_2316,N_1965,N_1770);
nand U2317 (N_2317,N_1767,N_1587);
and U2318 (N_2318,N_1500,N_1844);
nand U2319 (N_2319,N_1898,N_1641);
nor U2320 (N_2320,N_1962,N_1584);
or U2321 (N_2321,N_1908,N_1745);
and U2322 (N_2322,N_1633,N_1985);
or U2323 (N_2323,N_1785,N_1558);
nor U2324 (N_2324,N_1873,N_1655);
and U2325 (N_2325,N_1900,N_1917);
and U2326 (N_2326,N_1720,N_1600);
xor U2327 (N_2327,N_1783,N_1981);
and U2328 (N_2328,N_1962,N_1723);
xnor U2329 (N_2329,N_1894,N_1819);
nand U2330 (N_2330,N_1690,N_1727);
or U2331 (N_2331,N_1565,N_1616);
or U2332 (N_2332,N_1833,N_1660);
nand U2333 (N_2333,N_1736,N_1849);
and U2334 (N_2334,N_1745,N_1762);
or U2335 (N_2335,N_1747,N_1741);
and U2336 (N_2336,N_1690,N_1778);
and U2337 (N_2337,N_1639,N_1721);
and U2338 (N_2338,N_1836,N_1541);
or U2339 (N_2339,N_1746,N_1519);
nand U2340 (N_2340,N_1567,N_1746);
or U2341 (N_2341,N_1936,N_1526);
or U2342 (N_2342,N_1899,N_1706);
xor U2343 (N_2343,N_1733,N_1937);
xor U2344 (N_2344,N_1991,N_1578);
xnor U2345 (N_2345,N_1624,N_1564);
xnor U2346 (N_2346,N_1703,N_1768);
or U2347 (N_2347,N_1813,N_1689);
nand U2348 (N_2348,N_1602,N_1992);
and U2349 (N_2349,N_1615,N_1902);
nand U2350 (N_2350,N_1876,N_1894);
or U2351 (N_2351,N_1846,N_1810);
xor U2352 (N_2352,N_1937,N_1863);
and U2353 (N_2353,N_1793,N_1557);
xnor U2354 (N_2354,N_1638,N_1606);
xnor U2355 (N_2355,N_1622,N_1943);
nor U2356 (N_2356,N_1795,N_1725);
and U2357 (N_2357,N_1523,N_1966);
nor U2358 (N_2358,N_1503,N_1747);
or U2359 (N_2359,N_1726,N_1566);
or U2360 (N_2360,N_1999,N_1530);
and U2361 (N_2361,N_1572,N_1860);
nand U2362 (N_2362,N_1755,N_1815);
and U2363 (N_2363,N_1863,N_1857);
xor U2364 (N_2364,N_1828,N_1537);
xnor U2365 (N_2365,N_1819,N_1540);
xor U2366 (N_2366,N_1615,N_1907);
or U2367 (N_2367,N_1809,N_1788);
and U2368 (N_2368,N_1760,N_1544);
nand U2369 (N_2369,N_1659,N_1613);
nand U2370 (N_2370,N_1655,N_1523);
and U2371 (N_2371,N_1892,N_1724);
nand U2372 (N_2372,N_1975,N_1693);
nor U2373 (N_2373,N_1939,N_1513);
or U2374 (N_2374,N_1773,N_1638);
and U2375 (N_2375,N_1790,N_1607);
nor U2376 (N_2376,N_1514,N_1507);
nand U2377 (N_2377,N_1772,N_1750);
nand U2378 (N_2378,N_1799,N_1691);
or U2379 (N_2379,N_1789,N_1984);
xnor U2380 (N_2380,N_1988,N_1728);
nor U2381 (N_2381,N_1626,N_1536);
nand U2382 (N_2382,N_1672,N_1731);
nand U2383 (N_2383,N_1860,N_1539);
nand U2384 (N_2384,N_1627,N_1640);
nand U2385 (N_2385,N_1942,N_1894);
and U2386 (N_2386,N_1910,N_1747);
and U2387 (N_2387,N_1686,N_1650);
or U2388 (N_2388,N_1536,N_1565);
nor U2389 (N_2389,N_1950,N_1542);
nor U2390 (N_2390,N_1799,N_1551);
nor U2391 (N_2391,N_1590,N_1849);
or U2392 (N_2392,N_1809,N_1976);
nand U2393 (N_2393,N_1955,N_1970);
and U2394 (N_2394,N_1744,N_1600);
nand U2395 (N_2395,N_1938,N_1669);
or U2396 (N_2396,N_1868,N_1881);
and U2397 (N_2397,N_1772,N_1719);
or U2398 (N_2398,N_1940,N_1870);
nor U2399 (N_2399,N_1810,N_1776);
nor U2400 (N_2400,N_1746,N_1808);
or U2401 (N_2401,N_1551,N_1795);
nor U2402 (N_2402,N_1600,N_1939);
nor U2403 (N_2403,N_1592,N_1767);
or U2404 (N_2404,N_1979,N_1527);
or U2405 (N_2405,N_1721,N_1729);
or U2406 (N_2406,N_1554,N_1632);
xor U2407 (N_2407,N_1604,N_1689);
or U2408 (N_2408,N_1500,N_1618);
and U2409 (N_2409,N_1529,N_1654);
or U2410 (N_2410,N_1834,N_1691);
xor U2411 (N_2411,N_1569,N_1800);
and U2412 (N_2412,N_1935,N_1881);
nor U2413 (N_2413,N_1856,N_1930);
xor U2414 (N_2414,N_1713,N_1920);
xnor U2415 (N_2415,N_1880,N_1938);
nor U2416 (N_2416,N_1972,N_1554);
nor U2417 (N_2417,N_1650,N_1933);
or U2418 (N_2418,N_1996,N_1679);
nand U2419 (N_2419,N_1914,N_1661);
nor U2420 (N_2420,N_1672,N_1907);
nand U2421 (N_2421,N_1725,N_1903);
xor U2422 (N_2422,N_1694,N_1766);
or U2423 (N_2423,N_1827,N_1655);
and U2424 (N_2424,N_1998,N_1566);
and U2425 (N_2425,N_1957,N_1616);
and U2426 (N_2426,N_1874,N_1884);
nand U2427 (N_2427,N_1672,N_1551);
xnor U2428 (N_2428,N_1941,N_1511);
nor U2429 (N_2429,N_1897,N_1723);
and U2430 (N_2430,N_1572,N_1559);
nand U2431 (N_2431,N_1773,N_1947);
and U2432 (N_2432,N_1804,N_1624);
or U2433 (N_2433,N_1597,N_1684);
or U2434 (N_2434,N_1750,N_1888);
xor U2435 (N_2435,N_1890,N_1533);
and U2436 (N_2436,N_1844,N_1970);
xnor U2437 (N_2437,N_1779,N_1921);
nand U2438 (N_2438,N_1522,N_1955);
and U2439 (N_2439,N_1810,N_1677);
and U2440 (N_2440,N_1940,N_1710);
xnor U2441 (N_2441,N_1936,N_1580);
xor U2442 (N_2442,N_1842,N_1646);
xor U2443 (N_2443,N_1965,N_1856);
and U2444 (N_2444,N_1638,N_1962);
or U2445 (N_2445,N_1639,N_1569);
nand U2446 (N_2446,N_1877,N_1559);
and U2447 (N_2447,N_1556,N_1954);
nor U2448 (N_2448,N_1608,N_1530);
and U2449 (N_2449,N_1512,N_1862);
or U2450 (N_2450,N_1594,N_1926);
or U2451 (N_2451,N_1733,N_1629);
and U2452 (N_2452,N_1847,N_1649);
and U2453 (N_2453,N_1919,N_1664);
nor U2454 (N_2454,N_1655,N_1695);
or U2455 (N_2455,N_1858,N_1557);
nor U2456 (N_2456,N_1751,N_1654);
nand U2457 (N_2457,N_1977,N_1846);
nand U2458 (N_2458,N_1567,N_1701);
nand U2459 (N_2459,N_1696,N_1864);
and U2460 (N_2460,N_1732,N_1772);
and U2461 (N_2461,N_1641,N_1722);
and U2462 (N_2462,N_1985,N_1813);
and U2463 (N_2463,N_1718,N_1815);
and U2464 (N_2464,N_1630,N_1784);
nand U2465 (N_2465,N_1604,N_1610);
nand U2466 (N_2466,N_1670,N_1988);
nand U2467 (N_2467,N_1618,N_1555);
or U2468 (N_2468,N_1613,N_1948);
nand U2469 (N_2469,N_1857,N_1623);
and U2470 (N_2470,N_1700,N_1736);
and U2471 (N_2471,N_1758,N_1894);
nand U2472 (N_2472,N_1883,N_1924);
and U2473 (N_2473,N_1759,N_1544);
xor U2474 (N_2474,N_1621,N_1697);
xnor U2475 (N_2475,N_1887,N_1836);
xor U2476 (N_2476,N_1527,N_1731);
nand U2477 (N_2477,N_1670,N_1727);
and U2478 (N_2478,N_1619,N_1578);
or U2479 (N_2479,N_1560,N_1737);
and U2480 (N_2480,N_1689,N_1952);
or U2481 (N_2481,N_1975,N_1846);
nand U2482 (N_2482,N_1866,N_1693);
and U2483 (N_2483,N_1785,N_1634);
or U2484 (N_2484,N_1530,N_1513);
nor U2485 (N_2485,N_1681,N_1882);
nor U2486 (N_2486,N_1982,N_1999);
and U2487 (N_2487,N_1512,N_1735);
or U2488 (N_2488,N_1820,N_1809);
xnor U2489 (N_2489,N_1724,N_1996);
nor U2490 (N_2490,N_1955,N_1931);
nor U2491 (N_2491,N_1679,N_1668);
xnor U2492 (N_2492,N_1890,N_1841);
xor U2493 (N_2493,N_1845,N_1518);
nor U2494 (N_2494,N_1873,N_1832);
or U2495 (N_2495,N_1844,N_1678);
nor U2496 (N_2496,N_1658,N_1972);
or U2497 (N_2497,N_1522,N_1788);
xnor U2498 (N_2498,N_1952,N_1938);
and U2499 (N_2499,N_1640,N_1984);
xor U2500 (N_2500,N_2341,N_2173);
xnor U2501 (N_2501,N_2412,N_2118);
and U2502 (N_2502,N_2382,N_2486);
nor U2503 (N_2503,N_2241,N_2469);
nor U2504 (N_2504,N_2286,N_2218);
nor U2505 (N_2505,N_2493,N_2162);
nand U2506 (N_2506,N_2045,N_2062);
nor U2507 (N_2507,N_2312,N_2001);
nor U2508 (N_2508,N_2338,N_2110);
nor U2509 (N_2509,N_2109,N_2029);
or U2510 (N_2510,N_2200,N_2405);
and U2511 (N_2511,N_2255,N_2306);
nor U2512 (N_2512,N_2335,N_2316);
xor U2513 (N_2513,N_2258,N_2104);
xor U2514 (N_2514,N_2346,N_2215);
xor U2515 (N_2515,N_2299,N_2055);
nor U2516 (N_2516,N_2112,N_2424);
or U2517 (N_2517,N_2330,N_2024);
and U2518 (N_2518,N_2047,N_2008);
or U2519 (N_2519,N_2261,N_2383);
nor U2520 (N_2520,N_2453,N_2149);
and U2521 (N_2521,N_2157,N_2441);
or U2522 (N_2522,N_2189,N_2248);
or U2523 (N_2523,N_2030,N_2042);
or U2524 (N_2524,N_2334,N_2415);
xor U2525 (N_2525,N_2426,N_2259);
or U2526 (N_2526,N_2183,N_2379);
xor U2527 (N_2527,N_2434,N_2016);
nand U2528 (N_2528,N_2211,N_2343);
or U2529 (N_2529,N_2369,N_2127);
xnor U2530 (N_2530,N_2221,N_2375);
and U2531 (N_2531,N_2284,N_2454);
nor U2532 (N_2532,N_2365,N_2397);
nor U2533 (N_2533,N_2219,N_2410);
and U2534 (N_2534,N_2317,N_2195);
and U2535 (N_2535,N_2083,N_2311);
and U2536 (N_2536,N_2264,N_2000);
xor U2537 (N_2537,N_2082,N_2452);
nand U2538 (N_2538,N_2425,N_2021);
and U2539 (N_2539,N_2287,N_2011);
xor U2540 (N_2540,N_2491,N_2433);
xnor U2541 (N_2541,N_2194,N_2488);
xor U2542 (N_2542,N_2033,N_2467);
or U2543 (N_2543,N_2065,N_2459);
or U2544 (N_2544,N_2440,N_2117);
nand U2545 (N_2545,N_2006,N_2435);
nor U2546 (N_2546,N_2199,N_2014);
nand U2547 (N_2547,N_2172,N_2290);
or U2548 (N_2548,N_2253,N_2096);
and U2549 (N_2549,N_2374,N_2023);
or U2550 (N_2550,N_2318,N_2304);
xor U2551 (N_2551,N_2308,N_2244);
nor U2552 (N_2552,N_2420,N_2164);
xor U2553 (N_2553,N_2305,N_2446);
nand U2554 (N_2554,N_2007,N_2429);
or U2555 (N_2555,N_2396,N_2430);
nor U2556 (N_2556,N_2128,N_2310);
and U2557 (N_2557,N_2391,N_2087);
xnor U2558 (N_2558,N_2296,N_2091);
or U2559 (N_2559,N_2050,N_2009);
or U2560 (N_2560,N_2034,N_2140);
and U2561 (N_2561,N_2465,N_2487);
or U2562 (N_2562,N_2276,N_2394);
and U2563 (N_2563,N_2484,N_2285);
or U2564 (N_2564,N_2460,N_2404);
nor U2565 (N_2565,N_2378,N_2462);
nor U2566 (N_2566,N_2409,N_2278);
xnor U2567 (N_2567,N_2414,N_2086);
nor U2568 (N_2568,N_2483,N_2456);
nor U2569 (N_2569,N_2431,N_2307);
nand U2570 (N_2570,N_2191,N_2471);
nand U2571 (N_2571,N_2282,N_2300);
and U2572 (N_2572,N_2231,N_2399);
nand U2573 (N_2573,N_2324,N_2075);
xnor U2574 (N_2574,N_2090,N_2381);
xor U2575 (N_2575,N_2158,N_2130);
xnor U2576 (N_2576,N_2068,N_2201);
nand U2577 (N_2577,N_2245,N_2099);
nor U2578 (N_2578,N_2057,N_2327);
and U2579 (N_2579,N_2035,N_2040);
nand U2580 (N_2580,N_2283,N_2210);
or U2581 (N_2581,N_2060,N_2468);
or U2582 (N_2582,N_2407,N_2344);
nand U2583 (N_2583,N_2279,N_2103);
nor U2584 (N_2584,N_2406,N_2223);
xnor U2585 (N_2585,N_2249,N_2386);
nor U2586 (N_2586,N_2037,N_2098);
nor U2587 (N_2587,N_2333,N_2178);
or U2588 (N_2588,N_2170,N_2018);
nor U2589 (N_2589,N_2227,N_2234);
nor U2590 (N_2590,N_2085,N_2228);
nand U2591 (N_2591,N_2095,N_2137);
nor U2592 (N_2592,N_2078,N_2266);
nor U2593 (N_2593,N_2202,N_2289);
xnor U2594 (N_2594,N_2072,N_2256);
xnor U2595 (N_2595,N_2461,N_2269);
or U2596 (N_2596,N_2108,N_2036);
nand U2597 (N_2597,N_2364,N_2362);
or U2598 (N_2598,N_2247,N_2153);
nor U2599 (N_2599,N_2438,N_2163);
nand U2600 (N_2600,N_2190,N_2226);
nand U2601 (N_2601,N_2133,N_2229);
or U2602 (N_2602,N_2076,N_2161);
and U2603 (N_2603,N_2455,N_2268);
or U2604 (N_2604,N_2193,N_2233);
nand U2605 (N_2605,N_2031,N_2359);
nand U2606 (N_2606,N_2063,N_2361);
xor U2607 (N_2607,N_2336,N_2353);
or U2608 (N_2608,N_2373,N_2054);
xnor U2609 (N_2609,N_2070,N_2146);
and U2610 (N_2610,N_2222,N_2134);
xor U2611 (N_2611,N_2175,N_2303);
or U2612 (N_2612,N_2052,N_2182);
or U2613 (N_2613,N_2297,N_2225);
xor U2614 (N_2614,N_2220,N_2114);
and U2615 (N_2615,N_2489,N_2351);
nor U2616 (N_2616,N_2402,N_2411);
nand U2617 (N_2617,N_2464,N_2155);
and U2618 (N_2618,N_2192,N_2432);
nand U2619 (N_2619,N_2315,N_2025);
nor U2620 (N_2620,N_2003,N_2092);
xnor U2621 (N_2621,N_2165,N_2478);
xnor U2622 (N_2622,N_2358,N_2198);
nand U2623 (N_2623,N_2337,N_2094);
or U2624 (N_2624,N_2398,N_2214);
xor U2625 (N_2625,N_2458,N_2026);
nand U2626 (N_2626,N_2295,N_2450);
and U2627 (N_2627,N_2292,N_2348);
nor U2628 (N_2628,N_2445,N_2498);
xnor U2629 (N_2629,N_2122,N_2254);
or U2630 (N_2630,N_2345,N_2235);
or U2631 (N_2631,N_2027,N_2107);
and U2632 (N_2632,N_2013,N_2265);
and U2633 (N_2633,N_2101,N_2332);
nor U2634 (N_2634,N_2143,N_2106);
or U2635 (N_2635,N_2097,N_2288);
nor U2636 (N_2636,N_2370,N_2230);
nor U2637 (N_2637,N_2367,N_2120);
or U2638 (N_2638,N_2197,N_2105);
or U2639 (N_2639,N_2102,N_2490);
or U2640 (N_2640,N_2419,N_2262);
nand U2641 (N_2641,N_2319,N_2115);
nand U2642 (N_2642,N_2320,N_2022);
nand U2643 (N_2643,N_2472,N_2213);
xnor U2644 (N_2644,N_2499,N_2387);
nand U2645 (N_2645,N_2015,N_2160);
or U2646 (N_2646,N_2205,N_2119);
and U2647 (N_2647,N_2251,N_2475);
and U2648 (N_2648,N_2041,N_2185);
and U2649 (N_2649,N_2028,N_2147);
xnor U2650 (N_2650,N_2314,N_2084);
nor U2651 (N_2651,N_2238,N_2243);
nand U2652 (N_2652,N_2340,N_2207);
nand U2653 (N_2653,N_2196,N_2088);
xor U2654 (N_2654,N_2270,N_2372);
and U2655 (N_2655,N_2321,N_2174);
and U2656 (N_2656,N_2368,N_2302);
and U2657 (N_2657,N_2236,N_2326);
or U2658 (N_2658,N_2171,N_2043);
nor U2659 (N_2659,N_2049,N_2492);
nor U2660 (N_2660,N_2141,N_2208);
nor U2661 (N_2661,N_2093,N_2217);
xor U2662 (N_2662,N_2377,N_2322);
and U2663 (N_2663,N_2131,N_2145);
nor U2664 (N_2664,N_2357,N_2389);
or U2665 (N_2665,N_2017,N_2395);
or U2666 (N_2666,N_2126,N_2277);
or U2667 (N_2667,N_2239,N_2350);
xnor U2668 (N_2668,N_2044,N_2002);
and U2669 (N_2669,N_2129,N_2206);
xnor U2670 (N_2670,N_2476,N_2156);
nand U2671 (N_2671,N_2242,N_2298);
and U2672 (N_2672,N_2355,N_2176);
nand U2673 (N_2673,N_2212,N_2442);
nor U2674 (N_2674,N_2293,N_2309);
nor U2675 (N_2675,N_2449,N_2080);
xor U2676 (N_2676,N_2051,N_2271);
or U2677 (N_2677,N_2485,N_2148);
nor U2678 (N_2678,N_2166,N_2479);
and U2679 (N_2679,N_2366,N_2418);
xor U2680 (N_2680,N_2111,N_2046);
xnor U2681 (N_2681,N_2342,N_2463);
or U2682 (N_2682,N_2413,N_2482);
or U2683 (N_2683,N_2132,N_2142);
and U2684 (N_2684,N_2301,N_2349);
xor U2685 (N_2685,N_2480,N_2474);
or U2686 (N_2686,N_2329,N_2451);
nand U2687 (N_2687,N_2186,N_2038);
or U2688 (N_2688,N_2177,N_2204);
xnor U2689 (N_2689,N_2376,N_2039);
xnor U2690 (N_2690,N_2100,N_2447);
and U2691 (N_2691,N_2073,N_2135);
xor U2692 (N_2692,N_2237,N_2352);
and U2693 (N_2693,N_2074,N_2356);
or U2694 (N_2694,N_2354,N_2089);
xnor U2695 (N_2695,N_2392,N_2181);
nand U2696 (N_2696,N_2184,N_2058);
xnor U2697 (N_2697,N_2281,N_2403);
and U2698 (N_2698,N_2187,N_2466);
xor U2699 (N_2699,N_2116,N_2152);
xnor U2700 (N_2700,N_2053,N_2064);
or U2701 (N_2701,N_2470,N_2019);
or U2702 (N_2702,N_2428,N_2457);
and U2703 (N_2703,N_2067,N_2380);
xnor U2704 (N_2704,N_2439,N_2497);
xnor U2705 (N_2705,N_2159,N_2401);
xnor U2706 (N_2706,N_2246,N_2209);
nand U2707 (N_2707,N_2384,N_2416);
nand U2708 (N_2708,N_2180,N_2390);
or U2709 (N_2709,N_2151,N_2275);
nand U2710 (N_2710,N_2291,N_2313);
nor U2711 (N_2711,N_2077,N_2144);
nand U2712 (N_2712,N_2121,N_2331);
nor U2713 (N_2713,N_2168,N_2477);
xor U2714 (N_2714,N_2494,N_2079);
xnor U2715 (N_2715,N_2444,N_2005);
or U2716 (N_2716,N_2150,N_2056);
nor U2717 (N_2717,N_2123,N_2136);
nor U2718 (N_2718,N_2360,N_2436);
xor U2719 (N_2719,N_2260,N_2169);
nand U2720 (N_2720,N_2417,N_2385);
nand U2721 (N_2721,N_2481,N_2280);
nand U2722 (N_2722,N_2179,N_2393);
xnor U2723 (N_2723,N_2495,N_2294);
xnor U2724 (N_2724,N_2216,N_2081);
or U2725 (N_2725,N_2257,N_2421);
nor U2726 (N_2726,N_2422,N_2347);
nor U2727 (N_2727,N_2113,N_2363);
or U2728 (N_2728,N_2203,N_2124);
nor U2729 (N_2729,N_2061,N_2125);
or U2730 (N_2730,N_2423,N_2020);
or U2731 (N_2731,N_2267,N_2069);
and U2732 (N_2732,N_2328,N_2188);
nor U2733 (N_2733,N_2273,N_2012);
xnor U2734 (N_2734,N_2010,N_2388);
nand U2735 (N_2735,N_2437,N_2071);
and U2736 (N_2736,N_2448,N_2443);
and U2737 (N_2737,N_2272,N_2496);
or U2738 (N_2738,N_2263,N_2004);
and U2739 (N_2739,N_2154,N_2224);
xnor U2740 (N_2740,N_2473,N_2408);
and U2741 (N_2741,N_2167,N_2325);
or U2742 (N_2742,N_2323,N_2059);
nor U2743 (N_2743,N_2250,N_2252);
nand U2744 (N_2744,N_2371,N_2427);
and U2745 (N_2745,N_2139,N_2048);
or U2746 (N_2746,N_2032,N_2232);
nand U2747 (N_2747,N_2066,N_2274);
or U2748 (N_2748,N_2138,N_2339);
and U2749 (N_2749,N_2240,N_2400);
nand U2750 (N_2750,N_2494,N_2356);
nor U2751 (N_2751,N_2022,N_2480);
nand U2752 (N_2752,N_2484,N_2392);
nor U2753 (N_2753,N_2259,N_2465);
nor U2754 (N_2754,N_2210,N_2088);
xnor U2755 (N_2755,N_2445,N_2084);
nor U2756 (N_2756,N_2225,N_2074);
nor U2757 (N_2757,N_2131,N_2086);
nor U2758 (N_2758,N_2312,N_2384);
or U2759 (N_2759,N_2488,N_2051);
nor U2760 (N_2760,N_2369,N_2411);
or U2761 (N_2761,N_2499,N_2267);
nor U2762 (N_2762,N_2366,N_2326);
nand U2763 (N_2763,N_2067,N_2476);
xor U2764 (N_2764,N_2251,N_2366);
and U2765 (N_2765,N_2358,N_2159);
nand U2766 (N_2766,N_2217,N_2053);
and U2767 (N_2767,N_2310,N_2359);
and U2768 (N_2768,N_2125,N_2349);
nor U2769 (N_2769,N_2211,N_2436);
xnor U2770 (N_2770,N_2364,N_2487);
and U2771 (N_2771,N_2007,N_2004);
nand U2772 (N_2772,N_2162,N_2426);
nor U2773 (N_2773,N_2250,N_2353);
nor U2774 (N_2774,N_2217,N_2224);
or U2775 (N_2775,N_2497,N_2389);
xor U2776 (N_2776,N_2444,N_2352);
nand U2777 (N_2777,N_2189,N_2015);
nand U2778 (N_2778,N_2344,N_2259);
nor U2779 (N_2779,N_2248,N_2439);
xor U2780 (N_2780,N_2229,N_2136);
or U2781 (N_2781,N_2107,N_2053);
nand U2782 (N_2782,N_2106,N_2035);
nand U2783 (N_2783,N_2459,N_2238);
and U2784 (N_2784,N_2479,N_2491);
nand U2785 (N_2785,N_2249,N_2100);
or U2786 (N_2786,N_2197,N_2145);
or U2787 (N_2787,N_2206,N_2056);
nor U2788 (N_2788,N_2465,N_2448);
nor U2789 (N_2789,N_2272,N_2248);
and U2790 (N_2790,N_2050,N_2349);
xnor U2791 (N_2791,N_2047,N_2451);
xnor U2792 (N_2792,N_2182,N_2372);
nor U2793 (N_2793,N_2033,N_2474);
nand U2794 (N_2794,N_2210,N_2029);
and U2795 (N_2795,N_2298,N_2439);
or U2796 (N_2796,N_2043,N_2210);
and U2797 (N_2797,N_2395,N_2066);
or U2798 (N_2798,N_2008,N_2041);
nor U2799 (N_2799,N_2127,N_2149);
xnor U2800 (N_2800,N_2092,N_2312);
xor U2801 (N_2801,N_2017,N_2300);
xor U2802 (N_2802,N_2307,N_2226);
nor U2803 (N_2803,N_2079,N_2003);
xor U2804 (N_2804,N_2015,N_2087);
and U2805 (N_2805,N_2389,N_2491);
xor U2806 (N_2806,N_2222,N_2238);
or U2807 (N_2807,N_2056,N_2398);
or U2808 (N_2808,N_2473,N_2229);
and U2809 (N_2809,N_2256,N_2109);
xor U2810 (N_2810,N_2112,N_2080);
nand U2811 (N_2811,N_2178,N_2001);
nor U2812 (N_2812,N_2091,N_2174);
xnor U2813 (N_2813,N_2461,N_2173);
and U2814 (N_2814,N_2142,N_2105);
or U2815 (N_2815,N_2340,N_2499);
nand U2816 (N_2816,N_2318,N_2034);
xnor U2817 (N_2817,N_2088,N_2316);
and U2818 (N_2818,N_2322,N_2374);
xor U2819 (N_2819,N_2035,N_2085);
nor U2820 (N_2820,N_2195,N_2133);
and U2821 (N_2821,N_2364,N_2427);
nand U2822 (N_2822,N_2186,N_2031);
or U2823 (N_2823,N_2189,N_2110);
or U2824 (N_2824,N_2029,N_2384);
or U2825 (N_2825,N_2451,N_2353);
nand U2826 (N_2826,N_2491,N_2131);
nor U2827 (N_2827,N_2343,N_2078);
or U2828 (N_2828,N_2316,N_2455);
or U2829 (N_2829,N_2033,N_2294);
xnor U2830 (N_2830,N_2041,N_2383);
and U2831 (N_2831,N_2095,N_2032);
xnor U2832 (N_2832,N_2187,N_2082);
nand U2833 (N_2833,N_2440,N_2065);
nor U2834 (N_2834,N_2089,N_2455);
and U2835 (N_2835,N_2098,N_2187);
or U2836 (N_2836,N_2146,N_2385);
nor U2837 (N_2837,N_2170,N_2132);
and U2838 (N_2838,N_2056,N_2055);
or U2839 (N_2839,N_2459,N_2099);
or U2840 (N_2840,N_2423,N_2480);
nor U2841 (N_2841,N_2489,N_2004);
nor U2842 (N_2842,N_2084,N_2473);
and U2843 (N_2843,N_2039,N_2368);
nand U2844 (N_2844,N_2130,N_2392);
nor U2845 (N_2845,N_2077,N_2114);
or U2846 (N_2846,N_2077,N_2461);
and U2847 (N_2847,N_2365,N_2334);
nand U2848 (N_2848,N_2298,N_2151);
nor U2849 (N_2849,N_2153,N_2481);
and U2850 (N_2850,N_2344,N_2377);
xor U2851 (N_2851,N_2203,N_2465);
or U2852 (N_2852,N_2139,N_2430);
nor U2853 (N_2853,N_2373,N_2169);
nor U2854 (N_2854,N_2399,N_2361);
nor U2855 (N_2855,N_2446,N_2225);
xor U2856 (N_2856,N_2337,N_2031);
nor U2857 (N_2857,N_2470,N_2164);
nand U2858 (N_2858,N_2406,N_2453);
xnor U2859 (N_2859,N_2065,N_2380);
nor U2860 (N_2860,N_2485,N_2373);
or U2861 (N_2861,N_2311,N_2255);
or U2862 (N_2862,N_2069,N_2270);
nor U2863 (N_2863,N_2235,N_2384);
xor U2864 (N_2864,N_2425,N_2206);
xnor U2865 (N_2865,N_2069,N_2391);
and U2866 (N_2866,N_2307,N_2488);
xor U2867 (N_2867,N_2067,N_2122);
nand U2868 (N_2868,N_2116,N_2094);
or U2869 (N_2869,N_2431,N_2201);
nand U2870 (N_2870,N_2457,N_2382);
and U2871 (N_2871,N_2006,N_2159);
nor U2872 (N_2872,N_2259,N_2021);
and U2873 (N_2873,N_2262,N_2093);
nand U2874 (N_2874,N_2225,N_2232);
nor U2875 (N_2875,N_2241,N_2208);
nor U2876 (N_2876,N_2068,N_2296);
nand U2877 (N_2877,N_2022,N_2170);
nor U2878 (N_2878,N_2372,N_2165);
nand U2879 (N_2879,N_2347,N_2029);
xnor U2880 (N_2880,N_2116,N_2374);
or U2881 (N_2881,N_2202,N_2037);
or U2882 (N_2882,N_2182,N_2126);
nor U2883 (N_2883,N_2266,N_2080);
xor U2884 (N_2884,N_2342,N_2169);
nand U2885 (N_2885,N_2292,N_2295);
xor U2886 (N_2886,N_2372,N_2448);
and U2887 (N_2887,N_2306,N_2373);
nor U2888 (N_2888,N_2468,N_2425);
or U2889 (N_2889,N_2168,N_2119);
or U2890 (N_2890,N_2302,N_2283);
xor U2891 (N_2891,N_2353,N_2464);
nand U2892 (N_2892,N_2212,N_2062);
and U2893 (N_2893,N_2093,N_2434);
or U2894 (N_2894,N_2051,N_2473);
nor U2895 (N_2895,N_2394,N_2493);
nor U2896 (N_2896,N_2474,N_2434);
nand U2897 (N_2897,N_2067,N_2254);
xnor U2898 (N_2898,N_2023,N_2406);
and U2899 (N_2899,N_2026,N_2125);
or U2900 (N_2900,N_2392,N_2295);
and U2901 (N_2901,N_2241,N_2152);
nand U2902 (N_2902,N_2382,N_2326);
nor U2903 (N_2903,N_2354,N_2130);
nand U2904 (N_2904,N_2497,N_2036);
nor U2905 (N_2905,N_2102,N_2406);
nor U2906 (N_2906,N_2156,N_2148);
nand U2907 (N_2907,N_2124,N_2331);
nor U2908 (N_2908,N_2453,N_2437);
nand U2909 (N_2909,N_2252,N_2106);
nand U2910 (N_2910,N_2373,N_2062);
xnor U2911 (N_2911,N_2201,N_2200);
or U2912 (N_2912,N_2282,N_2112);
nand U2913 (N_2913,N_2379,N_2496);
or U2914 (N_2914,N_2227,N_2410);
nor U2915 (N_2915,N_2136,N_2429);
nand U2916 (N_2916,N_2299,N_2291);
and U2917 (N_2917,N_2407,N_2117);
and U2918 (N_2918,N_2203,N_2441);
xor U2919 (N_2919,N_2001,N_2348);
nor U2920 (N_2920,N_2109,N_2294);
xor U2921 (N_2921,N_2163,N_2277);
nand U2922 (N_2922,N_2112,N_2362);
and U2923 (N_2923,N_2038,N_2400);
xor U2924 (N_2924,N_2482,N_2489);
xor U2925 (N_2925,N_2253,N_2021);
nand U2926 (N_2926,N_2259,N_2164);
or U2927 (N_2927,N_2238,N_2328);
xor U2928 (N_2928,N_2230,N_2128);
nor U2929 (N_2929,N_2096,N_2443);
or U2930 (N_2930,N_2416,N_2046);
xnor U2931 (N_2931,N_2392,N_2209);
and U2932 (N_2932,N_2482,N_2144);
and U2933 (N_2933,N_2022,N_2476);
nand U2934 (N_2934,N_2426,N_2034);
and U2935 (N_2935,N_2211,N_2428);
nor U2936 (N_2936,N_2054,N_2331);
or U2937 (N_2937,N_2001,N_2330);
nor U2938 (N_2938,N_2109,N_2210);
nor U2939 (N_2939,N_2212,N_2412);
and U2940 (N_2940,N_2109,N_2372);
and U2941 (N_2941,N_2163,N_2034);
nand U2942 (N_2942,N_2346,N_2246);
and U2943 (N_2943,N_2043,N_2356);
and U2944 (N_2944,N_2384,N_2220);
and U2945 (N_2945,N_2040,N_2480);
xor U2946 (N_2946,N_2486,N_2132);
or U2947 (N_2947,N_2121,N_2441);
and U2948 (N_2948,N_2031,N_2380);
or U2949 (N_2949,N_2106,N_2009);
nor U2950 (N_2950,N_2280,N_2275);
nor U2951 (N_2951,N_2386,N_2129);
or U2952 (N_2952,N_2414,N_2234);
nor U2953 (N_2953,N_2452,N_2420);
nor U2954 (N_2954,N_2498,N_2375);
nor U2955 (N_2955,N_2376,N_2058);
nor U2956 (N_2956,N_2054,N_2333);
xnor U2957 (N_2957,N_2277,N_2080);
nand U2958 (N_2958,N_2412,N_2045);
xor U2959 (N_2959,N_2201,N_2434);
or U2960 (N_2960,N_2080,N_2050);
and U2961 (N_2961,N_2324,N_2234);
nor U2962 (N_2962,N_2068,N_2209);
nand U2963 (N_2963,N_2350,N_2044);
and U2964 (N_2964,N_2398,N_2061);
xnor U2965 (N_2965,N_2108,N_2098);
or U2966 (N_2966,N_2429,N_2308);
nor U2967 (N_2967,N_2349,N_2066);
and U2968 (N_2968,N_2005,N_2300);
or U2969 (N_2969,N_2097,N_2165);
or U2970 (N_2970,N_2344,N_2411);
or U2971 (N_2971,N_2352,N_2131);
xor U2972 (N_2972,N_2258,N_2084);
or U2973 (N_2973,N_2269,N_2040);
nor U2974 (N_2974,N_2497,N_2041);
xnor U2975 (N_2975,N_2059,N_2479);
xnor U2976 (N_2976,N_2234,N_2448);
nand U2977 (N_2977,N_2360,N_2243);
nor U2978 (N_2978,N_2400,N_2029);
or U2979 (N_2979,N_2358,N_2483);
or U2980 (N_2980,N_2391,N_2456);
nand U2981 (N_2981,N_2434,N_2367);
xnor U2982 (N_2982,N_2272,N_2065);
nor U2983 (N_2983,N_2201,N_2136);
xor U2984 (N_2984,N_2143,N_2117);
nand U2985 (N_2985,N_2154,N_2213);
nor U2986 (N_2986,N_2342,N_2242);
nand U2987 (N_2987,N_2375,N_2121);
and U2988 (N_2988,N_2429,N_2281);
xnor U2989 (N_2989,N_2364,N_2005);
or U2990 (N_2990,N_2397,N_2255);
nand U2991 (N_2991,N_2190,N_2484);
nand U2992 (N_2992,N_2464,N_2146);
xnor U2993 (N_2993,N_2490,N_2035);
nand U2994 (N_2994,N_2398,N_2081);
or U2995 (N_2995,N_2372,N_2346);
and U2996 (N_2996,N_2096,N_2457);
or U2997 (N_2997,N_2404,N_2150);
and U2998 (N_2998,N_2242,N_2473);
nor U2999 (N_2999,N_2159,N_2330);
nor U3000 (N_3000,N_2644,N_2915);
nor U3001 (N_3001,N_2710,N_2734);
nand U3002 (N_3002,N_2592,N_2613);
nand U3003 (N_3003,N_2525,N_2507);
xor U3004 (N_3004,N_2810,N_2890);
nand U3005 (N_3005,N_2912,N_2696);
and U3006 (N_3006,N_2987,N_2673);
xnor U3007 (N_3007,N_2858,N_2751);
or U3008 (N_3008,N_2919,N_2582);
nand U3009 (N_3009,N_2714,N_2950);
and U3010 (N_3010,N_2889,N_2554);
or U3011 (N_3011,N_2952,N_2593);
nor U3012 (N_3012,N_2578,N_2505);
or U3013 (N_3013,N_2743,N_2579);
nand U3014 (N_3014,N_2670,N_2686);
or U3015 (N_3015,N_2532,N_2882);
and U3016 (N_3016,N_2865,N_2977);
nor U3017 (N_3017,N_2960,N_2654);
nand U3018 (N_3018,N_2756,N_2971);
or U3019 (N_3019,N_2610,N_2638);
xor U3020 (N_3020,N_2989,N_2930);
nand U3021 (N_3021,N_2556,N_2885);
nor U3022 (N_3022,N_2985,N_2551);
and U3023 (N_3023,N_2732,N_2851);
nor U3024 (N_3024,N_2716,N_2522);
xnor U3025 (N_3025,N_2776,N_2903);
nor U3026 (N_3026,N_2516,N_2720);
nand U3027 (N_3027,N_2856,N_2777);
nand U3028 (N_3028,N_2968,N_2519);
and U3029 (N_3029,N_2785,N_2596);
nor U3030 (N_3030,N_2826,N_2941);
nor U3031 (N_3031,N_2850,N_2786);
or U3032 (N_3032,N_2991,N_2605);
nor U3033 (N_3033,N_2833,N_2929);
nor U3034 (N_3034,N_2626,N_2565);
nor U3035 (N_3035,N_2778,N_2552);
nand U3036 (N_3036,N_2840,N_2923);
nor U3037 (N_3037,N_2924,N_2528);
or U3038 (N_3038,N_2747,N_2750);
or U3039 (N_3039,N_2913,N_2540);
or U3040 (N_3040,N_2719,N_2650);
xnor U3041 (N_3041,N_2633,N_2748);
or U3042 (N_3042,N_2689,N_2606);
or U3043 (N_3043,N_2945,N_2764);
xnor U3044 (N_3044,N_2741,N_2667);
nor U3045 (N_3045,N_2585,N_2555);
nand U3046 (N_3046,N_2708,N_2940);
nand U3047 (N_3047,N_2523,N_2509);
nor U3048 (N_3048,N_2944,N_2958);
xor U3049 (N_3049,N_2895,N_2946);
and U3050 (N_3050,N_2706,N_2869);
nor U3051 (N_3051,N_2517,N_2775);
nand U3052 (N_3052,N_2543,N_2934);
nand U3053 (N_3053,N_2699,N_2953);
nand U3054 (N_3054,N_2894,N_2918);
or U3055 (N_3055,N_2587,N_2811);
nand U3056 (N_3056,N_2625,N_2725);
nand U3057 (N_3057,N_2692,N_2653);
nand U3058 (N_3058,N_2768,N_2938);
xor U3059 (N_3059,N_2612,N_2855);
nor U3060 (N_3060,N_2992,N_2622);
or U3061 (N_3061,N_2904,N_2683);
nand U3062 (N_3062,N_2691,N_2588);
nand U3063 (N_3063,N_2922,N_2570);
or U3064 (N_3064,N_2760,N_2624);
xnor U3065 (N_3065,N_2539,N_2986);
or U3066 (N_3066,N_2729,N_2600);
and U3067 (N_3067,N_2602,N_2640);
or U3068 (N_3068,N_2513,N_2998);
or U3069 (N_3069,N_2503,N_2726);
nand U3070 (N_3070,N_2680,N_2707);
nand U3071 (N_3071,N_2907,N_2619);
xnor U3072 (N_3072,N_2510,N_2685);
nand U3073 (N_3073,N_2550,N_2808);
or U3074 (N_3074,N_2717,N_2835);
and U3075 (N_3075,N_2701,N_2787);
and U3076 (N_3076,N_2576,N_2676);
or U3077 (N_3077,N_2979,N_2949);
or U3078 (N_3078,N_2661,N_2749);
or U3079 (N_3079,N_2766,N_2780);
nand U3080 (N_3080,N_2873,N_2901);
or U3081 (N_3081,N_2688,N_2642);
and U3082 (N_3082,N_2623,N_2893);
nor U3083 (N_3083,N_2942,N_2862);
nand U3084 (N_3084,N_2698,N_2871);
xor U3085 (N_3085,N_2713,N_2982);
xnor U3086 (N_3086,N_2620,N_2783);
or U3087 (N_3087,N_2879,N_2595);
nor U3088 (N_3088,N_2700,N_2662);
nor U3089 (N_3089,N_2796,N_2860);
or U3090 (N_3090,N_2562,N_2527);
xor U3091 (N_3091,N_2993,N_2621);
or U3092 (N_3092,N_2542,N_2534);
and U3093 (N_3093,N_2872,N_2891);
or U3094 (N_3094,N_2997,N_2731);
xor U3095 (N_3095,N_2880,N_2791);
nor U3096 (N_3096,N_2788,N_2607);
nand U3097 (N_3097,N_2917,N_2800);
xor U3098 (N_3098,N_2859,N_2802);
and U3099 (N_3099,N_2837,N_2843);
nand U3100 (N_3100,N_2886,N_2765);
xor U3101 (N_3101,N_2666,N_2948);
nor U3102 (N_3102,N_2795,N_2844);
and U3103 (N_3103,N_2853,N_2704);
xnor U3104 (N_3104,N_2951,N_2921);
and U3105 (N_3105,N_2656,N_2966);
xnor U3106 (N_3106,N_2736,N_2687);
and U3107 (N_3107,N_2599,N_2658);
or U3108 (N_3108,N_2645,N_2611);
or U3109 (N_3109,N_2506,N_2641);
or U3110 (N_3110,N_2639,N_2976);
nor U3111 (N_3111,N_2967,N_2573);
nor U3112 (N_3112,N_2936,N_2723);
nand U3113 (N_3113,N_2758,N_2836);
or U3114 (N_3114,N_2888,N_2730);
or U3115 (N_3115,N_2630,N_2695);
and U3116 (N_3116,N_2518,N_2501);
nand U3117 (N_3117,N_2580,N_2793);
or U3118 (N_3118,N_2694,N_2744);
or U3119 (N_3119,N_2931,N_2779);
or U3120 (N_3120,N_2804,N_2569);
and U3121 (N_3121,N_2679,N_2927);
nor U3122 (N_3122,N_2549,N_2925);
nand U3123 (N_3123,N_2712,N_2847);
nor U3124 (N_3124,N_2845,N_2737);
nand U3125 (N_3125,N_2868,N_2502);
nand U3126 (N_3126,N_2660,N_2589);
nand U3127 (N_3127,N_2838,N_2545);
xor U3128 (N_3128,N_2628,N_2636);
nand U3129 (N_3129,N_2863,N_2957);
nand U3130 (N_3130,N_2892,N_2818);
nand U3131 (N_3131,N_2995,N_2659);
and U3132 (N_3132,N_2875,N_2947);
nand U3133 (N_3133,N_2914,N_2801);
or U3134 (N_3134,N_2575,N_2740);
xnor U3135 (N_3135,N_2981,N_2728);
xor U3136 (N_3136,N_2854,N_2754);
nor U3137 (N_3137,N_2646,N_2813);
nand U3138 (N_3138,N_2684,N_2681);
nand U3139 (N_3139,N_2905,N_2789);
and U3140 (N_3140,N_2559,N_2512);
xor U3141 (N_3141,N_2671,N_2781);
and U3142 (N_3142,N_2965,N_2933);
or U3143 (N_3143,N_2887,N_2537);
or U3144 (N_3144,N_2896,N_2735);
and U3145 (N_3145,N_2900,N_2797);
or U3146 (N_3146,N_2648,N_2842);
and U3147 (N_3147,N_2757,N_2561);
or U3148 (N_3148,N_2530,N_2964);
nand U3149 (N_3149,N_2830,N_2742);
xor U3150 (N_3150,N_2746,N_2665);
or U3151 (N_3151,N_2805,N_2832);
nor U3152 (N_3152,N_2798,N_2821);
or U3153 (N_3153,N_2822,N_2643);
and U3154 (N_3154,N_2697,N_2583);
xnor U3155 (N_3155,N_2738,N_2655);
or U3156 (N_3156,N_2515,N_2771);
or U3157 (N_3157,N_2883,N_2548);
xnor U3158 (N_3158,N_2682,N_2755);
xnor U3159 (N_3159,N_2935,N_2975);
nand U3160 (N_3160,N_2718,N_2500);
nor U3161 (N_3161,N_2572,N_2631);
and U3162 (N_3162,N_2910,N_2649);
and U3163 (N_3163,N_2647,N_2829);
nand U3164 (N_3164,N_2560,N_2897);
and U3165 (N_3165,N_2721,N_2669);
nor U3166 (N_3166,N_2615,N_2999);
and U3167 (N_3167,N_2807,N_2564);
xor U3168 (N_3168,N_2908,N_2547);
nand U3169 (N_3169,N_2663,N_2841);
nor U3170 (N_3170,N_2831,N_2806);
nor U3171 (N_3171,N_2514,N_2752);
nand U3172 (N_3172,N_2531,N_2943);
nand U3173 (N_3173,N_2774,N_2815);
xnor U3174 (N_3174,N_2745,N_2814);
nand U3175 (N_3175,N_2767,N_2651);
nor U3176 (N_3176,N_2970,N_2614);
xor U3177 (N_3177,N_2809,N_2703);
nand U3178 (N_3178,N_2533,N_2857);
xor U3179 (N_3179,N_2616,N_2784);
nor U3180 (N_3180,N_2727,N_2792);
xnor U3181 (N_3181,N_2761,N_2693);
xnor U3182 (N_3182,N_2586,N_2541);
or U3183 (N_3183,N_2911,N_2773);
nand U3184 (N_3184,N_2823,N_2916);
nor U3185 (N_3185,N_2820,N_2790);
and U3186 (N_3186,N_2920,N_2584);
xor U3187 (N_3187,N_2996,N_2972);
nand U3188 (N_3188,N_2978,N_2902);
xor U3189 (N_3189,N_2508,N_2603);
xnor U3190 (N_3190,N_2724,N_2980);
and U3191 (N_3191,N_2963,N_2668);
or U3192 (N_3192,N_2772,N_2617);
xnor U3193 (N_3193,N_2794,N_2799);
nor U3194 (N_3194,N_2812,N_2544);
xnor U3195 (N_3195,N_2594,N_2962);
nand U3196 (N_3196,N_2878,N_2990);
xor U3197 (N_3197,N_2711,N_2898);
nand U3198 (N_3198,N_2637,N_2803);
and U3199 (N_3199,N_2598,N_2909);
or U3200 (N_3200,N_2846,N_2526);
nand U3201 (N_3201,N_2675,N_2816);
nand U3202 (N_3202,N_2881,N_2994);
nor U3203 (N_3203,N_2827,N_2866);
nor U3204 (N_3204,N_2674,N_2874);
nor U3205 (N_3205,N_2652,N_2877);
nor U3206 (N_3206,N_2954,N_2702);
nand U3207 (N_3207,N_2635,N_2769);
and U3208 (N_3208,N_2715,N_2961);
xor U3209 (N_3209,N_2690,N_2884);
and U3210 (N_3210,N_2535,N_2571);
xnor U3211 (N_3211,N_2627,N_2536);
xor U3212 (N_3212,N_2566,N_2739);
and U3213 (N_3213,N_2973,N_2817);
xor U3214 (N_3214,N_2988,N_2664);
nor U3215 (N_3215,N_2849,N_2591);
nor U3216 (N_3216,N_2770,N_2733);
xor U3217 (N_3217,N_2722,N_2618);
and U3218 (N_3218,N_2601,N_2557);
xor U3219 (N_3219,N_2538,N_2906);
nor U3220 (N_3220,N_2870,N_2529);
nor U3221 (N_3221,N_2546,N_2705);
nand U3222 (N_3222,N_2558,N_2932);
xor U3223 (N_3223,N_2763,N_2782);
or U3224 (N_3224,N_2937,N_2928);
xnor U3225 (N_3225,N_2959,N_2597);
xor U3226 (N_3226,N_2955,N_2864);
or U3227 (N_3227,N_2520,N_2553);
nand U3228 (N_3228,N_2574,N_2672);
nor U3229 (N_3229,N_2629,N_2511);
nor U3230 (N_3230,N_2521,N_2825);
and U3231 (N_3231,N_2969,N_2608);
xnor U3232 (N_3232,N_2867,N_2848);
xor U3233 (N_3233,N_2568,N_2590);
or U3234 (N_3234,N_2876,N_2604);
xor U3235 (N_3235,N_2899,N_2828);
nor U3236 (N_3236,N_2834,N_2504);
and U3237 (N_3237,N_2956,N_2567);
or U3238 (N_3238,N_2984,N_2759);
xor U3239 (N_3239,N_2753,N_2819);
xnor U3240 (N_3240,N_2657,N_2824);
xor U3241 (N_3241,N_2632,N_2634);
and U3242 (N_3242,N_2709,N_2852);
nand U3243 (N_3243,N_2524,N_2762);
nand U3244 (N_3244,N_2577,N_2974);
xor U3245 (N_3245,N_2939,N_2983);
or U3246 (N_3246,N_2677,N_2926);
xor U3247 (N_3247,N_2563,N_2581);
nand U3248 (N_3248,N_2609,N_2861);
nor U3249 (N_3249,N_2678,N_2839);
or U3250 (N_3250,N_2552,N_2836);
and U3251 (N_3251,N_2750,N_2731);
and U3252 (N_3252,N_2737,N_2785);
and U3253 (N_3253,N_2953,N_2693);
and U3254 (N_3254,N_2584,N_2664);
or U3255 (N_3255,N_2572,N_2525);
nand U3256 (N_3256,N_2684,N_2926);
and U3257 (N_3257,N_2883,N_2880);
and U3258 (N_3258,N_2598,N_2505);
nand U3259 (N_3259,N_2686,N_2538);
or U3260 (N_3260,N_2736,N_2982);
nand U3261 (N_3261,N_2718,N_2599);
or U3262 (N_3262,N_2922,N_2695);
nor U3263 (N_3263,N_2507,N_2600);
or U3264 (N_3264,N_2619,N_2753);
or U3265 (N_3265,N_2836,N_2676);
and U3266 (N_3266,N_2525,N_2562);
or U3267 (N_3267,N_2654,N_2752);
or U3268 (N_3268,N_2828,N_2736);
xor U3269 (N_3269,N_2892,N_2522);
xor U3270 (N_3270,N_2784,N_2773);
xnor U3271 (N_3271,N_2710,N_2850);
xnor U3272 (N_3272,N_2925,N_2783);
or U3273 (N_3273,N_2619,N_2774);
or U3274 (N_3274,N_2857,N_2619);
and U3275 (N_3275,N_2597,N_2650);
or U3276 (N_3276,N_2905,N_2904);
and U3277 (N_3277,N_2627,N_2525);
and U3278 (N_3278,N_2859,N_2723);
nor U3279 (N_3279,N_2534,N_2858);
or U3280 (N_3280,N_2720,N_2941);
nor U3281 (N_3281,N_2881,N_2604);
nor U3282 (N_3282,N_2941,N_2943);
nor U3283 (N_3283,N_2909,N_2946);
xor U3284 (N_3284,N_2992,N_2572);
or U3285 (N_3285,N_2599,N_2900);
and U3286 (N_3286,N_2891,N_2517);
and U3287 (N_3287,N_2673,N_2830);
xor U3288 (N_3288,N_2775,N_2818);
nand U3289 (N_3289,N_2614,N_2755);
and U3290 (N_3290,N_2621,N_2628);
nor U3291 (N_3291,N_2989,N_2983);
nand U3292 (N_3292,N_2552,N_2969);
nand U3293 (N_3293,N_2836,N_2619);
nor U3294 (N_3294,N_2506,N_2693);
nand U3295 (N_3295,N_2695,N_2665);
nor U3296 (N_3296,N_2926,N_2954);
or U3297 (N_3297,N_2525,N_2818);
and U3298 (N_3298,N_2625,N_2803);
or U3299 (N_3299,N_2779,N_2957);
nand U3300 (N_3300,N_2854,N_2882);
nor U3301 (N_3301,N_2859,N_2676);
or U3302 (N_3302,N_2777,N_2974);
and U3303 (N_3303,N_2751,N_2638);
nand U3304 (N_3304,N_2697,N_2503);
nand U3305 (N_3305,N_2721,N_2798);
or U3306 (N_3306,N_2971,N_2999);
nor U3307 (N_3307,N_2614,N_2540);
nand U3308 (N_3308,N_2645,N_2520);
nor U3309 (N_3309,N_2830,N_2653);
xor U3310 (N_3310,N_2629,N_2851);
or U3311 (N_3311,N_2871,N_2696);
xor U3312 (N_3312,N_2969,N_2907);
and U3313 (N_3313,N_2759,N_2831);
xnor U3314 (N_3314,N_2937,N_2664);
nor U3315 (N_3315,N_2558,N_2984);
xnor U3316 (N_3316,N_2998,N_2520);
nand U3317 (N_3317,N_2996,N_2512);
xnor U3318 (N_3318,N_2714,N_2906);
and U3319 (N_3319,N_2826,N_2830);
nor U3320 (N_3320,N_2925,N_2959);
or U3321 (N_3321,N_2756,N_2976);
nor U3322 (N_3322,N_2591,N_2995);
nand U3323 (N_3323,N_2555,N_2680);
and U3324 (N_3324,N_2804,N_2633);
or U3325 (N_3325,N_2767,N_2670);
or U3326 (N_3326,N_2776,N_2603);
or U3327 (N_3327,N_2724,N_2749);
nor U3328 (N_3328,N_2515,N_2655);
and U3329 (N_3329,N_2612,N_2992);
and U3330 (N_3330,N_2845,N_2637);
xor U3331 (N_3331,N_2674,N_2786);
or U3332 (N_3332,N_2621,N_2933);
nor U3333 (N_3333,N_2827,N_2821);
nand U3334 (N_3334,N_2965,N_2724);
and U3335 (N_3335,N_2745,N_2586);
xor U3336 (N_3336,N_2906,N_2705);
nand U3337 (N_3337,N_2974,N_2763);
and U3338 (N_3338,N_2647,N_2717);
xnor U3339 (N_3339,N_2703,N_2678);
nor U3340 (N_3340,N_2535,N_2550);
xnor U3341 (N_3341,N_2679,N_2974);
and U3342 (N_3342,N_2850,N_2597);
or U3343 (N_3343,N_2857,N_2515);
or U3344 (N_3344,N_2537,N_2522);
nand U3345 (N_3345,N_2874,N_2878);
xnor U3346 (N_3346,N_2916,N_2773);
nand U3347 (N_3347,N_2512,N_2871);
and U3348 (N_3348,N_2899,N_2908);
nand U3349 (N_3349,N_2554,N_2801);
nor U3350 (N_3350,N_2519,N_2695);
nor U3351 (N_3351,N_2681,N_2687);
nand U3352 (N_3352,N_2506,N_2930);
xnor U3353 (N_3353,N_2736,N_2881);
xnor U3354 (N_3354,N_2746,N_2507);
and U3355 (N_3355,N_2544,N_2590);
nor U3356 (N_3356,N_2965,N_2817);
xnor U3357 (N_3357,N_2982,N_2587);
and U3358 (N_3358,N_2983,N_2527);
and U3359 (N_3359,N_2730,N_2788);
and U3360 (N_3360,N_2662,N_2728);
xnor U3361 (N_3361,N_2695,N_2820);
nand U3362 (N_3362,N_2831,N_2967);
and U3363 (N_3363,N_2772,N_2917);
xor U3364 (N_3364,N_2724,N_2624);
nand U3365 (N_3365,N_2862,N_2644);
nor U3366 (N_3366,N_2614,N_2570);
or U3367 (N_3367,N_2578,N_2721);
nand U3368 (N_3368,N_2966,N_2888);
nand U3369 (N_3369,N_2535,N_2988);
xor U3370 (N_3370,N_2888,N_2995);
or U3371 (N_3371,N_2953,N_2904);
nor U3372 (N_3372,N_2991,N_2983);
or U3373 (N_3373,N_2990,N_2577);
nand U3374 (N_3374,N_2674,N_2730);
nand U3375 (N_3375,N_2949,N_2894);
xor U3376 (N_3376,N_2577,N_2636);
or U3377 (N_3377,N_2927,N_2529);
xnor U3378 (N_3378,N_2801,N_2930);
nor U3379 (N_3379,N_2967,N_2572);
or U3380 (N_3380,N_2946,N_2710);
nand U3381 (N_3381,N_2771,N_2586);
xor U3382 (N_3382,N_2590,N_2814);
xor U3383 (N_3383,N_2902,N_2941);
xor U3384 (N_3384,N_2681,N_2963);
nor U3385 (N_3385,N_2531,N_2927);
or U3386 (N_3386,N_2728,N_2671);
nand U3387 (N_3387,N_2766,N_2967);
nor U3388 (N_3388,N_2786,N_2621);
nor U3389 (N_3389,N_2927,N_2665);
nand U3390 (N_3390,N_2561,N_2629);
or U3391 (N_3391,N_2783,N_2767);
and U3392 (N_3392,N_2971,N_2617);
or U3393 (N_3393,N_2849,N_2507);
nor U3394 (N_3394,N_2641,N_2801);
or U3395 (N_3395,N_2898,N_2708);
xnor U3396 (N_3396,N_2821,N_2833);
nor U3397 (N_3397,N_2753,N_2515);
and U3398 (N_3398,N_2893,N_2630);
xnor U3399 (N_3399,N_2773,N_2544);
nor U3400 (N_3400,N_2893,N_2597);
xor U3401 (N_3401,N_2859,N_2819);
and U3402 (N_3402,N_2662,N_2773);
or U3403 (N_3403,N_2675,N_2952);
xnor U3404 (N_3404,N_2572,N_2938);
or U3405 (N_3405,N_2986,N_2899);
nand U3406 (N_3406,N_2715,N_2676);
xnor U3407 (N_3407,N_2966,N_2989);
xor U3408 (N_3408,N_2712,N_2522);
or U3409 (N_3409,N_2625,N_2783);
xnor U3410 (N_3410,N_2838,N_2754);
nor U3411 (N_3411,N_2865,N_2515);
nand U3412 (N_3412,N_2512,N_2777);
nand U3413 (N_3413,N_2907,N_2518);
nor U3414 (N_3414,N_2513,N_2879);
nand U3415 (N_3415,N_2811,N_2987);
xor U3416 (N_3416,N_2873,N_2913);
or U3417 (N_3417,N_2701,N_2537);
xnor U3418 (N_3418,N_2981,N_2985);
nand U3419 (N_3419,N_2744,N_2909);
nor U3420 (N_3420,N_2948,N_2736);
or U3421 (N_3421,N_2786,N_2854);
nand U3422 (N_3422,N_2911,N_2712);
nor U3423 (N_3423,N_2997,N_2689);
nand U3424 (N_3424,N_2855,N_2700);
nand U3425 (N_3425,N_2639,N_2637);
xor U3426 (N_3426,N_2997,N_2633);
and U3427 (N_3427,N_2533,N_2869);
xor U3428 (N_3428,N_2765,N_2903);
xor U3429 (N_3429,N_2981,N_2649);
or U3430 (N_3430,N_2667,N_2526);
and U3431 (N_3431,N_2877,N_2992);
and U3432 (N_3432,N_2764,N_2563);
xnor U3433 (N_3433,N_2832,N_2942);
or U3434 (N_3434,N_2643,N_2896);
nand U3435 (N_3435,N_2664,N_2538);
and U3436 (N_3436,N_2840,N_2755);
nor U3437 (N_3437,N_2968,N_2567);
or U3438 (N_3438,N_2604,N_2865);
and U3439 (N_3439,N_2824,N_2949);
xnor U3440 (N_3440,N_2670,N_2863);
xnor U3441 (N_3441,N_2915,N_2849);
or U3442 (N_3442,N_2576,N_2668);
nand U3443 (N_3443,N_2835,N_2844);
or U3444 (N_3444,N_2609,N_2875);
and U3445 (N_3445,N_2666,N_2518);
or U3446 (N_3446,N_2525,N_2553);
or U3447 (N_3447,N_2972,N_2641);
xnor U3448 (N_3448,N_2935,N_2599);
and U3449 (N_3449,N_2696,N_2532);
or U3450 (N_3450,N_2905,N_2791);
and U3451 (N_3451,N_2802,N_2683);
and U3452 (N_3452,N_2753,N_2587);
or U3453 (N_3453,N_2996,N_2541);
nand U3454 (N_3454,N_2874,N_2986);
nor U3455 (N_3455,N_2699,N_2702);
or U3456 (N_3456,N_2835,N_2649);
and U3457 (N_3457,N_2506,N_2640);
or U3458 (N_3458,N_2908,N_2764);
nor U3459 (N_3459,N_2701,N_2611);
nand U3460 (N_3460,N_2720,N_2676);
or U3461 (N_3461,N_2612,N_2509);
or U3462 (N_3462,N_2830,N_2713);
and U3463 (N_3463,N_2830,N_2567);
xor U3464 (N_3464,N_2674,N_2618);
and U3465 (N_3465,N_2926,N_2671);
nand U3466 (N_3466,N_2504,N_2599);
and U3467 (N_3467,N_2886,N_2525);
nor U3468 (N_3468,N_2574,N_2730);
or U3469 (N_3469,N_2522,N_2619);
or U3470 (N_3470,N_2610,N_2731);
and U3471 (N_3471,N_2527,N_2702);
or U3472 (N_3472,N_2836,N_2614);
nor U3473 (N_3473,N_2523,N_2732);
nand U3474 (N_3474,N_2965,N_2610);
nand U3475 (N_3475,N_2909,N_2922);
xor U3476 (N_3476,N_2625,N_2881);
nand U3477 (N_3477,N_2614,N_2799);
xnor U3478 (N_3478,N_2988,N_2738);
nor U3479 (N_3479,N_2677,N_2551);
xnor U3480 (N_3480,N_2774,N_2996);
xor U3481 (N_3481,N_2681,N_2561);
or U3482 (N_3482,N_2820,N_2642);
or U3483 (N_3483,N_2752,N_2911);
nor U3484 (N_3484,N_2590,N_2531);
xor U3485 (N_3485,N_2927,N_2548);
nand U3486 (N_3486,N_2827,N_2783);
and U3487 (N_3487,N_2846,N_2765);
xor U3488 (N_3488,N_2589,N_2953);
nand U3489 (N_3489,N_2921,N_2538);
xor U3490 (N_3490,N_2789,N_2569);
or U3491 (N_3491,N_2647,N_2837);
xnor U3492 (N_3492,N_2928,N_2860);
nor U3493 (N_3493,N_2851,N_2707);
nand U3494 (N_3494,N_2916,N_2584);
xor U3495 (N_3495,N_2776,N_2535);
nor U3496 (N_3496,N_2815,N_2716);
nand U3497 (N_3497,N_2852,N_2522);
or U3498 (N_3498,N_2710,N_2910);
nor U3499 (N_3499,N_2884,N_2789);
or U3500 (N_3500,N_3213,N_3276);
and U3501 (N_3501,N_3383,N_3287);
or U3502 (N_3502,N_3490,N_3084);
and U3503 (N_3503,N_3325,N_3046);
nand U3504 (N_3504,N_3464,N_3482);
xor U3505 (N_3505,N_3074,N_3223);
or U3506 (N_3506,N_3251,N_3060);
xor U3507 (N_3507,N_3115,N_3127);
nor U3508 (N_3508,N_3369,N_3378);
xor U3509 (N_3509,N_3112,N_3049);
nand U3510 (N_3510,N_3061,N_3089);
and U3511 (N_3511,N_3456,N_3004);
or U3512 (N_3512,N_3437,N_3097);
or U3513 (N_3513,N_3452,N_3343);
nand U3514 (N_3514,N_3023,N_3182);
nor U3515 (N_3515,N_3096,N_3289);
xor U3516 (N_3516,N_3384,N_3457);
and U3517 (N_3517,N_3387,N_3044);
and U3518 (N_3518,N_3405,N_3245);
or U3519 (N_3519,N_3226,N_3022);
xor U3520 (N_3520,N_3390,N_3282);
nor U3521 (N_3521,N_3497,N_3180);
nor U3522 (N_3522,N_3431,N_3400);
nor U3523 (N_3523,N_3170,N_3380);
nor U3524 (N_3524,N_3110,N_3359);
and U3525 (N_3525,N_3140,N_3016);
and U3526 (N_3526,N_3391,N_3056);
or U3527 (N_3527,N_3485,N_3346);
nor U3528 (N_3528,N_3007,N_3135);
and U3529 (N_3529,N_3263,N_3364);
xnor U3530 (N_3530,N_3072,N_3026);
and U3531 (N_3531,N_3093,N_3336);
nand U3532 (N_3532,N_3206,N_3261);
xnor U3533 (N_3533,N_3113,N_3069);
nand U3534 (N_3534,N_3045,N_3453);
or U3535 (N_3535,N_3329,N_3114);
and U3536 (N_3536,N_3001,N_3487);
xor U3537 (N_3537,N_3429,N_3296);
or U3538 (N_3538,N_3129,N_3143);
nor U3539 (N_3539,N_3273,N_3350);
or U3540 (N_3540,N_3164,N_3165);
nor U3541 (N_3541,N_3322,N_3011);
nor U3542 (N_3542,N_3407,N_3435);
or U3543 (N_3543,N_3411,N_3377);
nor U3544 (N_3544,N_3462,N_3106);
xnor U3545 (N_3545,N_3416,N_3412);
xnor U3546 (N_3546,N_3393,N_3076);
nand U3547 (N_3547,N_3066,N_3250);
nand U3548 (N_3548,N_3493,N_3181);
or U3549 (N_3549,N_3150,N_3098);
and U3550 (N_3550,N_3006,N_3328);
nor U3551 (N_3551,N_3057,N_3190);
and U3552 (N_3552,N_3302,N_3363);
or U3553 (N_3553,N_3252,N_3237);
or U3554 (N_3554,N_3185,N_3025);
or U3555 (N_3555,N_3036,N_3428);
nor U3556 (N_3556,N_3399,N_3275);
xnor U3557 (N_3557,N_3100,N_3173);
xnor U3558 (N_3558,N_3238,N_3065);
nor U3559 (N_3559,N_3230,N_3027);
xnor U3560 (N_3560,N_3099,N_3055);
or U3561 (N_3561,N_3280,N_3402);
nand U3562 (N_3562,N_3316,N_3395);
and U3563 (N_3563,N_3345,N_3332);
nand U3564 (N_3564,N_3196,N_3444);
xnor U3565 (N_3565,N_3175,N_3422);
xnor U3566 (N_3566,N_3063,N_3342);
and U3567 (N_3567,N_3019,N_3310);
and U3568 (N_3568,N_3448,N_3126);
or U3569 (N_3569,N_3147,N_3078);
xor U3570 (N_3570,N_3153,N_3091);
nor U3571 (N_3571,N_3246,N_3494);
nand U3572 (N_3572,N_3235,N_3403);
or U3573 (N_3573,N_3291,N_3201);
or U3574 (N_3574,N_3161,N_3268);
and U3575 (N_3575,N_3174,N_3212);
and U3576 (N_3576,N_3272,N_3210);
nor U3577 (N_3577,N_3458,N_3151);
nor U3578 (N_3578,N_3095,N_3389);
or U3579 (N_3579,N_3087,N_3463);
and U3580 (N_3580,N_3119,N_3320);
xnor U3581 (N_3581,N_3205,N_3303);
or U3582 (N_3582,N_3495,N_3498);
xor U3583 (N_3583,N_3123,N_3202);
xnor U3584 (N_3584,N_3171,N_3081);
and U3585 (N_3585,N_3312,N_3481);
xnor U3586 (N_3586,N_3461,N_3187);
and U3587 (N_3587,N_3484,N_3349);
nor U3588 (N_3588,N_3160,N_3128);
and U3589 (N_3589,N_3386,N_3301);
nor U3590 (N_3590,N_3353,N_3366);
and U3591 (N_3591,N_3020,N_3274);
and U3592 (N_3592,N_3396,N_3042);
nor U3593 (N_3593,N_3483,N_3382);
nor U3594 (N_3594,N_3440,N_3469);
nand U3595 (N_3595,N_3133,N_3433);
xor U3596 (N_3596,N_3374,N_3092);
and U3597 (N_3597,N_3136,N_3079);
or U3598 (N_3598,N_3459,N_3334);
nand U3599 (N_3599,N_3008,N_3077);
or U3600 (N_3600,N_3284,N_3002);
nor U3601 (N_3601,N_3313,N_3466);
nand U3602 (N_3602,N_3293,N_3299);
nand U3603 (N_3603,N_3264,N_3169);
or U3604 (N_3604,N_3130,N_3064);
nor U3605 (N_3605,N_3050,N_3294);
xnor U3606 (N_3606,N_3124,N_3253);
nand U3607 (N_3607,N_3224,N_3362);
nand U3608 (N_3608,N_3259,N_3376);
nand U3609 (N_3609,N_3474,N_3239);
xor U3610 (N_3610,N_3271,N_3247);
and U3611 (N_3611,N_3297,N_3028);
xor U3612 (N_3612,N_3300,N_3473);
nor U3613 (N_3613,N_3214,N_3496);
nor U3614 (N_3614,N_3138,N_3357);
xnor U3615 (N_3615,N_3356,N_3218);
or U3616 (N_3616,N_3015,N_3305);
nand U3617 (N_3617,N_3471,N_3186);
and U3618 (N_3618,N_3162,N_3075);
nor U3619 (N_3619,N_3267,N_3118);
xnor U3620 (N_3620,N_3281,N_3441);
and U3621 (N_3621,N_3286,N_3260);
and U3622 (N_3622,N_3470,N_3032);
or U3623 (N_3623,N_3101,N_3005);
xnor U3624 (N_3624,N_3054,N_3472);
and U3625 (N_3625,N_3053,N_3047);
nor U3626 (N_3626,N_3070,N_3331);
or U3627 (N_3627,N_3195,N_3090);
and U3628 (N_3628,N_3365,N_3241);
xnor U3629 (N_3629,N_3058,N_3339);
or U3630 (N_3630,N_3012,N_3154);
nand U3631 (N_3631,N_3211,N_3168);
xor U3632 (N_3632,N_3425,N_3255);
xnor U3633 (N_3633,N_3492,N_3447);
and U3634 (N_3634,N_3499,N_3258);
or U3635 (N_3635,N_3385,N_3232);
or U3636 (N_3636,N_3432,N_3240);
or U3637 (N_3637,N_3103,N_3073);
xnor U3638 (N_3638,N_3468,N_3475);
xor U3639 (N_3639,N_3326,N_3409);
nand U3640 (N_3640,N_3315,N_3419);
or U3641 (N_3641,N_3397,N_3330);
and U3642 (N_3642,N_3478,N_3159);
xor U3643 (N_3643,N_3242,N_3455);
nor U3644 (N_3644,N_3145,N_3269);
nor U3645 (N_3645,N_3406,N_3184);
nand U3646 (N_3646,N_3489,N_3010);
and U3647 (N_3647,N_3318,N_3003);
nor U3648 (N_3648,N_3183,N_3144);
nor U3649 (N_3649,N_3141,N_3401);
nor U3650 (N_3650,N_3051,N_3423);
xnor U3651 (N_3651,N_3107,N_3236);
xnor U3652 (N_3652,N_3220,N_3225);
and U3653 (N_3653,N_3415,N_3085);
nor U3654 (N_3654,N_3352,N_3337);
or U3655 (N_3655,N_3449,N_3229);
nand U3656 (N_3656,N_3338,N_3347);
nor U3657 (N_3657,N_3341,N_3348);
or U3658 (N_3658,N_3013,N_3217);
or U3659 (N_3659,N_3094,N_3413);
and U3660 (N_3660,N_3361,N_3249);
nor U3661 (N_3661,N_3421,N_3108);
nor U3662 (N_3662,N_3228,N_3248);
nor U3663 (N_3663,N_3277,N_3270);
xnor U3664 (N_3664,N_3031,N_3373);
nor U3665 (N_3665,N_3424,N_3434);
or U3666 (N_3666,N_3290,N_3368);
or U3667 (N_3667,N_3367,N_3048);
or U3668 (N_3668,N_3059,N_3445);
or U3669 (N_3669,N_3436,N_3351);
or U3670 (N_3670,N_3360,N_3176);
or U3671 (N_3671,N_3120,N_3139);
nand U3672 (N_3672,N_3354,N_3163);
or U3673 (N_3673,N_3319,N_3102);
nor U3674 (N_3674,N_3278,N_3324);
and U3675 (N_3675,N_3134,N_3039);
and U3676 (N_3676,N_3388,N_3137);
nand U3677 (N_3677,N_3306,N_3035);
nor U3678 (N_3678,N_3283,N_3323);
nand U3679 (N_3679,N_3000,N_3465);
nor U3680 (N_3680,N_3193,N_3179);
and U3681 (N_3681,N_3111,N_3146);
xnor U3682 (N_3682,N_3430,N_3295);
nand U3683 (N_3683,N_3370,N_3109);
or U3684 (N_3684,N_3189,N_3062);
and U3685 (N_3685,N_3067,N_3321);
nand U3686 (N_3686,N_3132,N_3344);
or U3687 (N_3687,N_3335,N_3298);
nand U3688 (N_3688,N_3256,N_3398);
and U3689 (N_3689,N_3191,N_3037);
or U3690 (N_3690,N_3410,N_3142);
nor U3691 (N_3691,N_3254,N_3450);
nor U3692 (N_3692,N_3314,N_3041);
and U3693 (N_3693,N_3265,N_3488);
and U3694 (N_3694,N_3199,N_3317);
or U3695 (N_3695,N_3204,N_3426);
and U3696 (N_3696,N_3408,N_3418);
xor U3697 (N_3697,N_3486,N_3038);
and U3698 (N_3698,N_3443,N_3192);
or U3699 (N_3699,N_3355,N_3207);
nor U3700 (N_3700,N_3309,N_3197);
nor U3701 (N_3701,N_3491,N_3172);
and U3702 (N_3702,N_3071,N_3231);
nand U3703 (N_3703,N_3243,N_3446);
nor U3704 (N_3704,N_3024,N_3279);
nor U3705 (N_3705,N_3311,N_3188);
nor U3706 (N_3706,N_3379,N_3477);
and U3707 (N_3707,N_3121,N_3266);
nor U3708 (N_3708,N_3149,N_3308);
nand U3709 (N_3709,N_3104,N_3476);
xor U3710 (N_3710,N_3009,N_3417);
nor U3711 (N_3711,N_3014,N_3152);
nand U3712 (N_3712,N_3375,N_3304);
and U3713 (N_3713,N_3414,N_3030);
nor U3714 (N_3714,N_3166,N_3033);
and U3715 (N_3715,N_3451,N_3381);
and U3716 (N_3716,N_3125,N_3285);
nand U3717 (N_3717,N_3262,N_3167);
xor U3718 (N_3718,N_3017,N_3480);
nand U3719 (N_3719,N_3333,N_3178);
xnor U3720 (N_3720,N_3122,N_3083);
xor U3721 (N_3721,N_3467,N_3340);
nand U3722 (N_3722,N_3244,N_3157);
nand U3723 (N_3723,N_3392,N_3068);
or U3724 (N_3724,N_3216,N_3439);
nor U3725 (N_3725,N_3233,N_3292);
nor U3726 (N_3726,N_3257,N_3288);
or U3727 (N_3727,N_3221,N_3194);
nand U3728 (N_3728,N_3394,N_3209);
xor U3729 (N_3729,N_3442,N_3080);
nand U3730 (N_3730,N_3043,N_3372);
xor U3731 (N_3731,N_3040,N_3117);
and U3732 (N_3732,N_3454,N_3029);
nor U3733 (N_3733,N_3427,N_3158);
xor U3734 (N_3734,N_3307,N_3021);
xnor U3735 (N_3735,N_3219,N_3198);
and U3736 (N_3736,N_3148,N_3034);
xnor U3737 (N_3737,N_3327,N_3131);
xor U3738 (N_3738,N_3088,N_3438);
nor U3739 (N_3739,N_3203,N_3222);
nor U3740 (N_3740,N_3105,N_3116);
or U3741 (N_3741,N_3155,N_3215);
xnor U3742 (N_3742,N_3052,N_3156);
xor U3743 (N_3743,N_3018,N_3177);
and U3744 (N_3744,N_3082,N_3479);
nor U3745 (N_3745,N_3086,N_3208);
nand U3746 (N_3746,N_3200,N_3234);
nor U3747 (N_3747,N_3371,N_3404);
or U3748 (N_3748,N_3227,N_3460);
xor U3749 (N_3749,N_3420,N_3358);
nand U3750 (N_3750,N_3476,N_3206);
nor U3751 (N_3751,N_3015,N_3002);
or U3752 (N_3752,N_3476,N_3011);
nand U3753 (N_3753,N_3247,N_3265);
nor U3754 (N_3754,N_3183,N_3019);
or U3755 (N_3755,N_3056,N_3446);
or U3756 (N_3756,N_3054,N_3201);
xnor U3757 (N_3757,N_3453,N_3278);
and U3758 (N_3758,N_3305,N_3440);
and U3759 (N_3759,N_3216,N_3428);
and U3760 (N_3760,N_3269,N_3322);
or U3761 (N_3761,N_3351,N_3231);
xor U3762 (N_3762,N_3293,N_3294);
and U3763 (N_3763,N_3142,N_3205);
or U3764 (N_3764,N_3490,N_3112);
and U3765 (N_3765,N_3082,N_3402);
xnor U3766 (N_3766,N_3033,N_3435);
or U3767 (N_3767,N_3126,N_3259);
nor U3768 (N_3768,N_3358,N_3129);
or U3769 (N_3769,N_3008,N_3131);
xor U3770 (N_3770,N_3078,N_3204);
nand U3771 (N_3771,N_3241,N_3416);
nand U3772 (N_3772,N_3217,N_3443);
xnor U3773 (N_3773,N_3377,N_3073);
and U3774 (N_3774,N_3087,N_3044);
or U3775 (N_3775,N_3442,N_3397);
nor U3776 (N_3776,N_3346,N_3337);
and U3777 (N_3777,N_3302,N_3170);
nor U3778 (N_3778,N_3067,N_3359);
nand U3779 (N_3779,N_3258,N_3374);
nand U3780 (N_3780,N_3284,N_3445);
xor U3781 (N_3781,N_3457,N_3067);
and U3782 (N_3782,N_3275,N_3496);
xor U3783 (N_3783,N_3244,N_3367);
nor U3784 (N_3784,N_3389,N_3270);
xor U3785 (N_3785,N_3332,N_3129);
nor U3786 (N_3786,N_3101,N_3160);
nor U3787 (N_3787,N_3182,N_3365);
or U3788 (N_3788,N_3051,N_3108);
or U3789 (N_3789,N_3051,N_3029);
xnor U3790 (N_3790,N_3084,N_3352);
xor U3791 (N_3791,N_3035,N_3335);
nand U3792 (N_3792,N_3181,N_3255);
xnor U3793 (N_3793,N_3358,N_3257);
and U3794 (N_3794,N_3466,N_3337);
or U3795 (N_3795,N_3089,N_3037);
and U3796 (N_3796,N_3294,N_3135);
or U3797 (N_3797,N_3047,N_3382);
or U3798 (N_3798,N_3448,N_3193);
and U3799 (N_3799,N_3450,N_3382);
xor U3800 (N_3800,N_3069,N_3159);
nand U3801 (N_3801,N_3457,N_3450);
nor U3802 (N_3802,N_3270,N_3200);
nor U3803 (N_3803,N_3202,N_3109);
or U3804 (N_3804,N_3455,N_3207);
nand U3805 (N_3805,N_3481,N_3327);
or U3806 (N_3806,N_3144,N_3156);
nand U3807 (N_3807,N_3087,N_3162);
xor U3808 (N_3808,N_3212,N_3498);
or U3809 (N_3809,N_3261,N_3011);
or U3810 (N_3810,N_3490,N_3241);
or U3811 (N_3811,N_3376,N_3248);
xor U3812 (N_3812,N_3448,N_3256);
and U3813 (N_3813,N_3165,N_3316);
or U3814 (N_3814,N_3325,N_3073);
xnor U3815 (N_3815,N_3147,N_3399);
xor U3816 (N_3816,N_3209,N_3239);
nand U3817 (N_3817,N_3284,N_3107);
or U3818 (N_3818,N_3302,N_3333);
nor U3819 (N_3819,N_3171,N_3297);
and U3820 (N_3820,N_3226,N_3394);
xor U3821 (N_3821,N_3352,N_3046);
nand U3822 (N_3822,N_3052,N_3021);
or U3823 (N_3823,N_3304,N_3443);
nand U3824 (N_3824,N_3166,N_3098);
xor U3825 (N_3825,N_3340,N_3386);
and U3826 (N_3826,N_3471,N_3173);
nor U3827 (N_3827,N_3417,N_3470);
nand U3828 (N_3828,N_3130,N_3160);
nor U3829 (N_3829,N_3027,N_3344);
xor U3830 (N_3830,N_3184,N_3482);
xor U3831 (N_3831,N_3458,N_3363);
and U3832 (N_3832,N_3380,N_3145);
xnor U3833 (N_3833,N_3013,N_3321);
or U3834 (N_3834,N_3480,N_3059);
xnor U3835 (N_3835,N_3243,N_3221);
or U3836 (N_3836,N_3310,N_3004);
xnor U3837 (N_3837,N_3228,N_3420);
nand U3838 (N_3838,N_3131,N_3446);
nand U3839 (N_3839,N_3063,N_3312);
nor U3840 (N_3840,N_3364,N_3262);
or U3841 (N_3841,N_3204,N_3383);
xnor U3842 (N_3842,N_3237,N_3377);
xnor U3843 (N_3843,N_3410,N_3029);
nor U3844 (N_3844,N_3188,N_3193);
nand U3845 (N_3845,N_3359,N_3338);
and U3846 (N_3846,N_3217,N_3170);
xnor U3847 (N_3847,N_3305,N_3455);
nor U3848 (N_3848,N_3360,N_3071);
and U3849 (N_3849,N_3018,N_3408);
and U3850 (N_3850,N_3297,N_3436);
and U3851 (N_3851,N_3246,N_3371);
xnor U3852 (N_3852,N_3278,N_3274);
xor U3853 (N_3853,N_3495,N_3352);
nand U3854 (N_3854,N_3170,N_3375);
and U3855 (N_3855,N_3053,N_3413);
nand U3856 (N_3856,N_3466,N_3449);
and U3857 (N_3857,N_3306,N_3039);
or U3858 (N_3858,N_3348,N_3316);
nand U3859 (N_3859,N_3456,N_3010);
nor U3860 (N_3860,N_3402,N_3099);
or U3861 (N_3861,N_3431,N_3238);
and U3862 (N_3862,N_3335,N_3409);
nor U3863 (N_3863,N_3170,N_3147);
nor U3864 (N_3864,N_3218,N_3035);
nor U3865 (N_3865,N_3095,N_3378);
or U3866 (N_3866,N_3212,N_3132);
xnor U3867 (N_3867,N_3358,N_3266);
nor U3868 (N_3868,N_3387,N_3045);
nor U3869 (N_3869,N_3443,N_3245);
nand U3870 (N_3870,N_3461,N_3357);
xor U3871 (N_3871,N_3388,N_3374);
xnor U3872 (N_3872,N_3298,N_3417);
or U3873 (N_3873,N_3138,N_3378);
nor U3874 (N_3874,N_3079,N_3360);
nor U3875 (N_3875,N_3260,N_3378);
nor U3876 (N_3876,N_3170,N_3389);
nor U3877 (N_3877,N_3416,N_3099);
xnor U3878 (N_3878,N_3009,N_3162);
xor U3879 (N_3879,N_3028,N_3098);
xor U3880 (N_3880,N_3254,N_3077);
xnor U3881 (N_3881,N_3419,N_3348);
or U3882 (N_3882,N_3383,N_3443);
or U3883 (N_3883,N_3221,N_3237);
nand U3884 (N_3884,N_3206,N_3236);
xor U3885 (N_3885,N_3219,N_3120);
xnor U3886 (N_3886,N_3297,N_3220);
or U3887 (N_3887,N_3092,N_3311);
or U3888 (N_3888,N_3253,N_3095);
or U3889 (N_3889,N_3251,N_3023);
or U3890 (N_3890,N_3376,N_3382);
nor U3891 (N_3891,N_3125,N_3291);
xnor U3892 (N_3892,N_3193,N_3199);
nor U3893 (N_3893,N_3254,N_3142);
or U3894 (N_3894,N_3236,N_3375);
xnor U3895 (N_3895,N_3349,N_3132);
or U3896 (N_3896,N_3166,N_3083);
nand U3897 (N_3897,N_3072,N_3338);
and U3898 (N_3898,N_3069,N_3416);
nand U3899 (N_3899,N_3325,N_3318);
or U3900 (N_3900,N_3131,N_3194);
nor U3901 (N_3901,N_3488,N_3095);
nor U3902 (N_3902,N_3063,N_3147);
nor U3903 (N_3903,N_3295,N_3206);
nand U3904 (N_3904,N_3209,N_3469);
and U3905 (N_3905,N_3179,N_3286);
nand U3906 (N_3906,N_3143,N_3018);
nor U3907 (N_3907,N_3354,N_3423);
nand U3908 (N_3908,N_3058,N_3273);
and U3909 (N_3909,N_3488,N_3007);
and U3910 (N_3910,N_3016,N_3397);
nand U3911 (N_3911,N_3340,N_3017);
nor U3912 (N_3912,N_3078,N_3022);
nand U3913 (N_3913,N_3381,N_3077);
nand U3914 (N_3914,N_3496,N_3088);
xor U3915 (N_3915,N_3416,N_3005);
xnor U3916 (N_3916,N_3014,N_3186);
nand U3917 (N_3917,N_3161,N_3375);
and U3918 (N_3918,N_3060,N_3331);
xnor U3919 (N_3919,N_3312,N_3350);
xnor U3920 (N_3920,N_3305,N_3331);
and U3921 (N_3921,N_3319,N_3063);
or U3922 (N_3922,N_3468,N_3153);
nor U3923 (N_3923,N_3487,N_3188);
nor U3924 (N_3924,N_3491,N_3110);
nand U3925 (N_3925,N_3385,N_3118);
nor U3926 (N_3926,N_3302,N_3491);
nor U3927 (N_3927,N_3335,N_3216);
nand U3928 (N_3928,N_3257,N_3386);
nand U3929 (N_3929,N_3114,N_3036);
xnor U3930 (N_3930,N_3199,N_3450);
and U3931 (N_3931,N_3225,N_3206);
nor U3932 (N_3932,N_3142,N_3270);
or U3933 (N_3933,N_3460,N_3134);
xnor U3934 (N_3934,N_3164,N_3261);
and U3935 (N_3935,N_3495,N_3324);
or U3936 (N_3936,N_3384,N_3485);
nor U3937 (N_3937,N_3489,N_3176);
xor U3938 (N_3938,N_3096,N_3440);
nand U3939 (N_3939,N_3093,N_3458);
or U3940 (N_3940,N_3308,N_3027);
nor U3941 (N_3941,N_3031,N_3418);
or U3942 (N_3942,N_3287,N_3356);
or U3943 (N_3943,N_3072,N_3282);
or U3944 (N_3944,N_3346,N_3418);
and U3945 (N_3945,N_3381,N_3209);
nor U3946 (N_3946,N_3056,N_3123);
nor U3947 (N_3947,N_3382,N_3389);
xor U3948 (N_3948,N_3332,N_3213);
nand U3949 (N_3949,N_3291,N_3368);
nand U3950 (N_3950,N_3290,N_3049);
nand U3951 (N_3951,N_3398,N_3022);
nor U3952 (N_3952,N_3231,N_3199);
nor U3953 (N_3953,N_3045,N_3145);
or U3954 (N_3954,N_3221,N_3344);
or U3955 (N_3955,N_3474,N_3272);
nand U3956 (N_3956,N_3248,N_3491);
and U3957 (N_3957,N_3364,N_3497);
and U3958 (N_3958,N_3448,N_3359);
and U3959 (N_3959,N_3405,N_3138);
or U3960 (N_3960,N_3063,N_3202);
and U3961 (N_3961,N_3466,N_3023);
nor U3962 (N_3962,N_3107,N_3033);
nor U3963 (N_3963,N_3085,N_3454);
or U3964 (N_3964,N_3173,N_3410);
and U3965 (N_3965,N_3209,N_3341);
nand U3966 (N_3966,N_3004,N_3256);
and U3967 (N_3967,N_3240,N_3355);
nand U3968 (N_3968,N_3440,N_3310);
or U3969 (N_3969,N_3011,N_3140);
nand U3970 (N_3970,N_3155,N_3285);
nand U3971 (N_3971,N_3444,N_3016);
nand U3972 (N_3972,N_3200,N_3376);
nand U3973 (N_3973,N_3319,N_3422);
and U3974 (N_3974,N_3033,N_3410);
xnor U3975 (N_3975,N_3053,N_3140);
and U3976 (N_3976,N_3425,N_3381);
nor U3977 (N_3977,N_3091,N_3250);
or U3978 (N_3978,N_3464,N_3457);
or U3979 (N_3979,N_3010,N_3127);
xor U3980 (N_3980,N_3136,N_3035);
or U3981 (N_3981,N_3281,N_3252);
nor U3982 (N_3982,N_3236,N_3190);
and U3983 (N_3983,N_3030,N_3098);
nand U3984 (N_3984,N_3281,N_3210);
nand U3985 (N_3985,N_3268,N_3281);
nor U3986 (N_3986,N_3301,N_3241);
nor U3987 (N_3987,N_3000,N_3158);
xor U3988 (N_3988,N_3113,N_3141);
xor U3989 (N_3989,N_3216,N_3169);
nor U3990 (N_3990,N_3101,N_3077);
xnor U3991 (N_3991,N_3386,N_3078);
nand U3992 (N_3992,N_3191,N_3464);
nand U3993 (N_3993,N_3394,N_3244);
xnor U3994 (N_3994,N_3435,N_3108);
xor U3995 (N_3995,N_3140,N_3151);
nand U3996 (N_3996,N_3387,N_3119);
or U3997 (N_3997,N_3012,N_3088);
nor U3998 (N_3998,N_3494,N_3000);
and U3999 (N_3999,N_3072,N_3043);
and U4000 (N_4000,N_3666,N_3535);
nand U4001 (N_4001,N_3677,N_3854);
xor U4002 (N_4002,N_3701,N_3532);
and U4003 (N_4003,N_3849,N_3507);
nor U4004 (N_4004,N_3927,N_3841);
xor U4005 (N_4005,N_3725,N_3605);
nor U4006 (N_4006,N_3846,N_3964);
nor U4007 (N_4007,N_3604,N_3529);
xor U4008 (N_4008,N_3610,N_3731);
nor U4009 (N_4009,N_3993,N_3974);
and U4010 (N_4010,N_3903,N_3843);
and U4011 (N_4011,N_3991,N_3543);
xnor U4012 (N_4012,N_3660,N_3819);
nand U4013 (N_4013,N_3918,N_3641);
nor U4014 (N_4014,N_3675,N_3852);
and U4015 (N_4015,N_3625,N_3602);
xnor U4016 (N_4016,N_3975,N_3549);
and U4017 (N_4017,N_3788,N_3945);
and U4018 (N_4018,N_3693,N_3779);
nand U4019 (N_4019,N_3805,N_3594);
nand U4020 (N_4020,N_3899,N_3703);
or U4021 (N_4021,N_3674,N_3957);
xor U4022 (N_4022,N_3867,N_3822);
and U4023 (N_4023,N_3868,N_3729);
and U4024 (N_4024,N_3670,N_3613);
or U4025 (N_4025,N_3542,N_3934);
or U4026 (N_4026,N_3679,N_3614);
xnor U4027 (N_4027,N_3711,N_3773);
or U4028 (N_4028,N_3801,N_3950);
xnor U4029 (N_4029,N_3816,N_3592);
nor U4030 (N_4030,N_3545,N_3980);
nand U4031 (N_4031,N_3859,N_3683);
xor U4032 (N_4032,N_3560,N_3633);
nor U4033 (N_4033,N_3530,N_3659);
xnor U4034 (N_4034,N_3962,N_3664);
nor U4035 (N_4035,N_3796,N_3724);
nand U4036 (N_4036,N_3735,N_3907);
xnor U4037 (N_4037,N_3580,N_3887);
or U4038 (N_4038,N_3533,N_3622);
and U4039 (N_4039,N_3932,N_3893);
nor U4040 (N_4040,N_3989,N_3869);
and U4041 (N_4041,N_3699,N_3621);
and U4042 (N_4042,N_3896,N_3971);
nand U4043 (N_4043,N_3730,N_3866);
and U4044 (N_4044,N_3727,N_3949);
nand U4045 (N_4045,N_3515,N_3704);
xor U4046 (N_4046,N_3764,N_3810);
or U4047 (N_4047,N_3759,N_3690);
nand U4048 (N_4048,N_3995,N_3557);
and U4049 (N_4049,N_3789,N_3923);
nor U4050 (N_4050,N_3829,N_3563);
or U4051 (N_4051,N_3953,N_3818);
and U4052 (N_4052,N_3576,N_3760);
xnor U4053 (N_4053,N_3910,N_3501);
or U4054 (N_4054,N_3774,N_3908);
and U4055 (N_4055,N_3740,N_3994);
nand U4056 (N_4056,N_3909,N_3514);
nand U4057 (N_4057,N_3698,N_3981);
or U4058 (N_4058,N_3714,N_3860);
nor U4059 (N_4059,N_3966,N_3642);
or U4060 (N_4060,N_3914,N_3657);
nor U4061 (N_4061,N_3820,N_3570);
or U4062 (N_4062,N_3987,N_3551);
and U4063 (N_4063,N_3799,N_3746);
and U4064 (N_4064,N_3607,N_3894);
nor U4065 (N_4065,N_3871,N_3983);
nand U4066 (N_4066,N_3750,N_3716);
and U4067 (N_4067,N_3598,N_3900);
nand U4068 (N_4068,N_3784,N_3895);
xnor U4069 (N_4069,N_3525,N_3733);
nand U4070 (N_4070,N_3958,N_3722);
and U4071 (N_4071,N_3700,N_3952);
xnor U4072 (N_4072,N_3970,N_3692);
or U4073 (N_4073,N_3837,N_3655);
nor U4074 (N_4074,N_3567,N_3520);
or U4075 (N_4075,N_3536,N_3850);
or U4076 (N_4076,N_3857,N_3999);
xnor U4077 (N_4077,N_3654,N_3890);
or U4078 (N_4078,N_3876,N_3782);
xnor U4079 (N_4079,N_3941,N_3673);
nand U4080 (N_4080,N_3645,N_3873);
xnor U4081 (N_4081,N_3769,N_3972);
nand U4082 (N_4082,N_3806,N_3590);
and U4083 (N_4083,N_3845,N_3745);
or U4084 (N_4084,N_3628,N_3791);
and U4085 (N_4085,N_3574,N_3901);
and U4086 (N_4086,N_3526,N_3689);
nor U4087 (N_4087,N_3636,N_3646);
nand U4088 (N_4088,N_3736,N_3835);
nand U4089 (N_4089,N_3978,N_3577);
or U4090 (N_4090,N_3634,N_3765);
nor U4091 (N_4091,N_3943,N_3865);
nand U4092 (N_4092,N_3540,N_3924);
xnor U4093 (N_4093,N_3794,N_3875);
xor U4094 (N_4094,N_3640,N_3627);
xor U4095 (N_4095,N_3824,N_3737);
nand U4096 (N_4096,N_3930,N_3620);
xnor U4097 (N_4097,N_3783,N_3742);
or U4098 (N_4098,N_3798,N_3967);
or U4099 (N_4099,N_3508,N_3635);
or U4100 (N_4100,N_3591,N_3696);
and U4101 (N_4101,N_3720,N_3911);
xor U4102 (N_4102,N_3792,N_3606);
nor U4103 (N_4103,N_3874,N_3979);
xnor U4104 (N_4104,N_3548,N_3732);
or U4105 (N_4105,N_3647,N_3787);
nand U4106 (N_4106,N_3573,N_3878);
and U4107 (N_4107,N_3889,N_3648);
nand U4108 (N_4108,N_3938,N_3644);
nor U4109 (N_4109,N_3990,N_3597);
nand U4110 (N_4110,N_3763,N_3596);
nand U4111 (N_4111,N_3856,N_3800);
nor U4112 (N_4112,N_3506,N_3617);
xor U4113 (N_4113,N_3821,N_3752);
nor U4114 (N_4114,N_3955,N_3539);
nor U4115 (N_4115,N_3559,N_3504);
nand U4116 (N_4116,N_3582,N_3685);
and U4117 (N_4117,N_3906,N_3578);
and U4118 (N_4118,N_3511,N_3589);
xnor U4119 (N_4119,N_3702,N_3947);
nand U4120 (N_4120,N_3982,N_3826);
nor U4121 (N_4121,N_3919,N_3804);
xnor U4122 (N_4122,N_3917,N_3780);
xor U4123 (N_4123,N_3695,N_3968);
and U4124 (N_4124,N_3961,N_3681);
nor U4125 (N_4125,N_3808,N_3913);
and U4126 (N_4126,N_3985,N_3505);
nand U4127 (N_4127,N_3753,N_3969);
nor U4128 (N_4128,N_3743,N_3652);
xnor U4129 (N_4129,N_3925,N_3562);
xor U4130 (N_4130,N_3823,N_3584);
nand U4131 (N_4131,N_3797,N_3715);
xnor U4132 (N_4132,N_3656,N_3882);
nand U4133 (N_4133,N_3976,N_3717);
nand U4134 (N_4134,N_3768,N_3948);
nand U4135 (N_4135,N_3767,N_3687);
and U4136 (N_4136,N_3940,N_3997);
or U4137 (N_4137,N_3847,N_3738);
nand U4138 (N_4138,N_3863,N_3619);
nand U4139 (N_4139,N_3631,N_3946);
nand U4140 (N_4140,N_3802,N_3706);
nand U4141 (N_4141,N_3682,N_3726);
or U4142 (N_4142,N_3762,N_3749);
or U4143 (N_4143,N_3747,N_3877);
and U4144 (N_4144,N_3755,N_3748);
nand U4145 (N_4145,N_3830,N_3708);
xnor U4146 (N_4146,N_3684,N_3928);
nor U4147 (N_4147,N_3963,N_3612);
nor U4148 (N_4148,N_3609,N_3579);
nor U4149 (N_4149,N_3828,N_3537);
nand U4150 (N_4150,N_3944,N_3977);
nand U4151 (N_4151,N_3915,N_3521);
or U4152 (N_4152,N_3758,N_3771);
and U4153 (N_4153,N_3676,N_3757);
nor U4154 (N_4154,N_3547,N_3776);
xor U4155 (N_4155,N_3965,N_3793);
or U4156 (N_4156,N_3766,N_3888);
or U4157 (N_4157,N_3996,N_3541);
xnor U4158 (N_4158,N_3565,N_3658);
nand U4159 (N_4159,N_3569,N_3669);
and U4160 (N_4160,N_3571,N_3761);
and U4161 (N_4161,N_3500,N_3516);
or U4162 (N_4162,N_3637,N_3650);
nor U4163 (N_4163,N_3886,N_3513);
or U4164 (N_4164,N_3840,N_3709);
and U4165 (N_4165,N_3916,N_3601);
or U4166 (N_4166,N_3705,N_3951);
xnor U4167 (N_4167,N_3667,N_3528);
nand U4168 (N_4168,N_3661,N_3772);
xor U4169 (N_4169,N_3599,N_3723);
or U4170 (N_4170,N_3831,N_3524);
xnor U4171 (N_4171,N_3555,N_3686);
nand U4172 (N_4172,N_3629,N_3992);
and U4173 (N_4173,N_3575,N_3904);
or U4174 (N_4174,N_3986,N_3643);
xor U4175 (N_4175,N_3812,N_3825);
nor U4176 (N_4176,N_3833,N_3956);
nor U4177 (N_4177,N_3593,N_3939);
or U4178 (N_4178,N_3552,N_3546);
and U4179 (N_4179,N_3814,N_3785);
or U4180 (N_4180,N_3663,N_3626);
or U4181 (N_4181,N_3921,N_3756);
nand U4182 (N_4182,N_3861,N_3639);
or U4183 (N_4183,N_3827,N_3694);
xnor U4184 (N_4184,N_3572,N_3662);
or U4185 (N_4185,N_3898,N_3554);
xor U4186 (N_4186,N_3836,N_3531);
nor U4187 (N_4187,N_3936,N_3885);
nor U4188 (N_4188,N_3544,N_3853);
nand U4189 (N_4189,N_3777,N_3710);
and U4190 (N_4190,N_3608,N_3522);
xor U4191 (N_4191,N_3988,N_3671);
and U4192 (N_4192,N_3728,N_3568);
or U4193 (N_4193,N_3902,N_3998);
nand U4194 (N_4194,N_3960,N_3653);
nor U4195 (N_4195,N_3811,N_3618);
nor U4196 (N_4196,N_3973,N_3564);
and U4197 (N_4197,N_3632,N_3984);
nor U4198 (N_4198,N_3600,N_3512);
nand U4199 (N_4199,N_3510,N_3550);
xor U4200 (N_4200,N_3770,N_3834);
xnor U4201 (N_4201,N_3668,N_3807);
nand U4202 (N_4202,N_3739,N_3842);
or U4203 (N_4203,N_3795,N_3817);
nor U4204 (N_4204,N_3623,N_3844);
or U4205 (N_4205,N_3697,N_3581);
xor U4206 (N_4206,N_3931,N_3527);
nand U4207 (N_4207,N_3721,N_3680);
and U4208 (N_4208,N_3615,N_3558);
and U4209 (N_4209,N_3864,N_3855);
and U4210 (N_4210,N_3870,N_3832);
or U4211 (N_4211,N_3707,N_3616);
nand U4212 (N_4212,N_3588,N_3920);
or U4213 (N_4213,N_3790,N_3712);
xor U4214 (N_4214,N_3942,N_3651);
nand U4215 (N_4215,N_3809,N_3713);
or U4216 (N_4216,N_3638,N_3879);
and U4217 (N_4217,N_3518,N_3803);
nor U4218 (N_4218,N_3534,N_3517);
nand U4219 (N_4219,N_3611,N_3858);
xor U4220 (N_4220,N_3880,N_3935);
nand U4221 (N_4221,N_3839,N_3678);
or U4222 (N_4222,N_3905,N_3929);
and U4223 (N_4223,N_3718,N_3933);
nor U4224 (N_4224,N_3851,N_3624);
xnor U4225 (N_4225,N_3926,N_3954);
or U4226 (N_4226,N_3538,N_3922);
nand U4227 (N_4227,N_3744,N_3891);
nor U4228 (N_4228,N_3523,N_3775);
or U4229 (N_4229,N_3553,N_3665);
nor U4230 (N_4230,N_3556,N_3881);
and U4231 (N_4231,N_3741,N_3587);
nor U4232 (N_4232,N_3872,N_3786);
and U4233 (N_4233,N_3892,N_3586);
nor U4234 (N_4234,N_3519,N_3848);
nand U4235 (N_4235,N_3719,N_3630);
xor U4236 (N_4236,N_3561,N_3566);
nand U4237 (N_4237,N_3897,N_3912);
xor U4238 (N_4238,N_3734,N_3509);
nor U4239 (N_4239,N_3778,N_3754);
xor U4240 (N_4240,N_3503,N_3959);
xnor U4241 (N_4241,N_3649,N_3862);
xnor U4242 (N_4242,N_3502,N_3603);
nor U4243 (N_4243,N_3595,N_3815);
nand U4244 (N_4244,N_3688,N_3583);
nor U4245 (N_4245,N_3838,N_3813);
nor U4246 (N_4246,N_3884,N_3691);
or U4247 (N_4247,N_3937,N_3585);
nor U4248 (N_4248,N_3883,N_3751);
xnor U4249 (N_4249,N_3781,N_3672);
or U4250 (N_4250,N_3865,N_3942);
nor U4251 (N_4251,N_3839,N_3574);
or U4252 (N_4252,N_3882,N_3935);
nand U4253 (N_4253,N_3701,N_3835);
nor U4254 (N_4254,N_3599,N_3549);
nor U4255 (N_4255,N_3808,N_3575);
and U4256 (N_4256,N_3999,N_3596);
nand U4257 (N_4257,N_3879,N_3865);
or U4258 (N_4258,N_3532,N_3880);
xor U4259 (N_4259,N_3623,N_3867);
nand U4260 (N_4260,N_3839,N_3797);
or U4261 (N_4261,N_3508,N_3630);
nor U4262 (N_4262,N_3675,N_3581);
nor U4263 (N_4263,N_3941,N_3738);
xor U4264 (N_4264,N_3994,N_3620);
nor U4265 (N_4265,N_3824,N_3659);
or U4266 (N_4266,N_3547,N_3789);
nand U4267 (N_4267,N_3701,N_3703);
nor U4268 (N_4268,N_3749,N_3871);
nor U4269 (N_4269,N_3578,N_3678);
and U4270 (N_4270,N_3701,N_3558);
or U4271 (N_4271,N_3524,N_3596);
nand U4272 (N_4272,N_3949,N_3792);
nand U4273 (N_4273,N_3509,N_3686);
or U4274 (N_4274,N_3682,N_3911);
nor U4275 (N_4275,N_3653,N_3921);
and U4276 (N_4276,N_3903,N_3886);
nor U4277 (N_4277,N_3587,N_3901);
xnor U4278 (N_4278,N_3936,N_3831);
nand U4279 (N_4279,N_3657,N_3826);
or U4280 (N_4280,N_3827,N_3821);
nand U4281 (N_4281,N_3934,N_3646);
nor U4282 (N_4282,N_3859,N_3674);
nand U4283 (N_4283,N_3827,N_3829);
and U4284 (N_4284,N_3611,N_3696);
nor U4285 (N_4285,N_3915,N_3868);
nor U4286 (N_4286,N_3792,N_3675);
or U4287 (N_4287,N_3709,N_3689);
nor U4288 (N_4288,N_3607,N_3568);
nor U4289 (N_4289,N_3722,N_3751);
xor U4290 (N_4290,N_3988,N_3667);
xnor U4291 (N_4291,N_3633,N_3895);
nand U4292 (N_4292,N_3652,N_3816);
and U4293 (N_4293,N_3642,N_3683);
nor U4294 (N_4294,N_3553,N_3980);
and U4295 (N_4295,N_3653,N_3584);
or U4296 (N_4296,N_3969,N_3987);
or U4297 (N_4297,N_3944,N_3909);
xnor U4298 (N_4298,N_3571,N_3971);
and U4299 (N_4299,N_3647,N_3877);
and U4300 (N_4300,N_3832,N_3598);
or U4301 (N_4301,N_3644,N_3913);
and U4302 (N_4302,N_3804,N_3574);
or U4303 (N_4303,N_3510,N_3756);
and U4304 (N_4304,N_3970,N_3606);
nor U4305 (N_4305,N_3761,N_3567);
nor U4306 (N_4306,N_3846,N_3575);
or U4307 (N_4307,N_3926,N_3945);
xnor U4308 (N_4308,N_3665,N_3562);
and U4309 (N_4309,N_3823,N_3775);
xnor U4310 (N_4310,N_3708,N_3990);
xor U4311 (N_4311,N_3805,N_3551);
xor U4312 (N_4312,N_3652,N_3980);
or U4313 (N_4313,N_3763,N_3571);
xor U4314 (N_4314,N_3856,N_3597);
and U4315 (N_4315,N_3538,N_3801);
nand U4316 (N_4316,N_3575,N_3763);
nor U4317 (N_4317,N_3601,N_3777);
nor U4318 (N_4318,N_3727,N_3811);
xor U4319 (N_4319,N_3554,N_3891);
or U4320 (N_4320,N_3898,N_3705);
nand U4321 (N_4321,N_3631,N_3546);
nor U4322 (N_4322,N_3866,N_3843);
nor U4323 (N_4323,N_3873,N_3719);
or U4324 (N_4324,N_3650,N_3723);
and U4325 (N_4325,N_3851,N_3964);
nor U4326 (N_4326,N_3635,N_3879);
xor U4327 (N_4327,N_3957,N_3796);
nor U4328 (N_4328,N_3945,N_3546);
xnor U4329 (N_4329,N_3852,N_3979);
and U4330 (N_4330,N_3732,N_3611);
and U4331 (N_4331,N_3626,N_3886);
and U4332 (N_4332,N_3971,N_3645);
or U4333 (N_4333,N_3870,N_3532);
or U4334 (N_4334,N_3720,N_3826);
nor U4335 (N_4335,N_3559,N_3890);
xnor U4336 (N_4336,N_3853,N_3866);
xor U4337 (N_4337,N_3720,N_3533);
and U4338 (N_4338,N_3502,N_3666);
nand U4339 (N_4339,N_3723,N_3691);
xnor U4340 (N_4340,N_3944,N_3630);
xnor U4341 (N_4341,N_3704,N_3615);
nand U4342 (N_4342,N_3670,N_3811);
nor U4343 (N_4343,N_3517,N_3537);
nor U4344 (N_4344,N_3990,N_3980);
xnor U4345 (N_4345,N_3846,N_3972);
nor U4346 (N_4346,N_3820,N_3779);
and U4347 (N_4347,N_3959,N_3828);
nand U4348 (N_4348,N_3939,N_3700);
xnor U4349 (N_4349,N_3612,N_3660);
xnor U4350 (N_4350,N_3541,N_3779);
nand U4351 (N_4351,N_3726,N_3850);
nor U4352 (N_4352,N_3587,N_3564);
and U4353 (N_4353,N_3740,N_3734);
nor U4354 (N_4354,N_3978,N_3693);
xnor U4355 (N_4355,N_3514,N_3582);
nand U4356 (N_4356,N_3610,N_3679);
nor U4357 (N_4357,N_3958,N_3748);
and U4358 (N_4358,N_3585,N_3870);
or U4359 (N_4359,N_3828,N_3504);
nand U4360 (N_4360,N_3893,N_3570);
xnor U4361 (N_4361,N_3969,N_3642);
or U4362 (N_4362,N_3839,N_3635);
or U4363 (N_4363,N_3878,N_3817);
and U4364 (N_4364,N_3650,N_3552);
nor U4365 (N_4365,N_3757,N_3902);
nor U4366 (N_4366,N_3830,N_3673);
and U4367 (N_4367,N_3901,N_3854);
nor U4368 (N_4368,N_3602,N_3762);
nor U4369 (N_4369,N_3986,N_3660);
nand U4370 (N_4370,N_3798,N_3672);
xnor U4371 (N_4371,N_3839,N_3509);
xor U4372 (N_4372,N_3944,N_3842);
and U4373 (N_4373,N_3851,N_3669);
and U4374 (N_4374,N_3992,N_3789);
nor U4375 (N_4375,N_3962,N_3652);
and U4376 (N_4376,N_3723,N_3976);
and U4377 (N_4377,N_3872,N_3964);
or U4378 (N_4378,N_3549,N_3965);
nand U4379 (N_4379,N_3867,N_3965);
nand U4380 (N_4380,N_3840,N_3683);
and U4381 (N_4381,N_3810,N_3852);
nor U4382 (N_4382,N_3716,N_3541);
and U4383 (N_4383,N_3968,N_3669);
and U4384 (N_4384,N_3840,N_3520);
nor U4385 (N_4385,N_3632,N_3977);
xnor U4386 (N_4386,N_3987,N_3508);
and U4387 (N_4387,N_3967,N_3538);
or U4388 (N_4388,N_3882,N_3770);
xor U4389 (N_4389,N_3843,N_3692);
nor U4390 (N_4390,N_3862,N_3996);
nand U4391 (N_4391,N_3746,N_3823);
nand U4392 (N_4392,N_3688,N_3884);
and U4393 (N_4393,N_3751,N_3761);
nand U4394 (N_4394,N_3502,N_3599);
and U4395 (N_4395,N_3537,N_3508);
or U4396 (N_4396,N_3531,N_3912);
and U4397 (N_4397,N_3811,N_3718);
and U4398 (N_4398,N_3505,N_3772);
and U4399 (N_4399,N_3920,N_3823);
nor U4400 (N_4400,N_3759,N_3863);
nand U4401 (N_4401,N_3993,N_3682);
or U4402 (N_4402,N_3514,N_3776);
or U4403 (N_4403,N_3933,N_3628);
nand U4404 (N_4404,N_3916,N_3997);
or U4405 (N_4405,N_3983,N_3962);
and U4406 (N_4406,N_3809,N_3608);
xor U4407 (N_4407,N_3880,N_3765);
and U4408 (N_4408,N_3659,N_3575);
nor U4409 (N_4409,N_3927,N_3784);
xnor U4410 (N_4410,N_3794,N_3917);
and U4411 (N_4411,N_3793,N_3674);
xor U4412 (N_4412,N_3958,N_3569);
nand U4413 (N_4413,N_3682,N_3684);
xor U4414 (N_4414,N_3874,N_3743);
xnor U4415 (N_4415,N_3746,N_3765);
nor U4416 (N_4416,N_3818,N_3709);
and U4417 (N_4417,N_3913,N_3712);
xor U4418 (N_4418,N_3547,N_3716);
or U4419 (N_4419,N_3838,N_3523);
nand U4420 (N_4420,N_3791,N_3658);
nand U4421 (N_4421,N_3742,N_3848);
or U4422 (N_4422,N_3983,N_3591);
or U4423 (N_4423,N_3548,N_3871);
or U4424 (N_4424,N_3617,N_3939);
and U4425 (N_4425,N_3676,N_3890);
and U4426 (N_4426,N_3879,N_3613);
nand U4427 (N_4427,N_3793,N_3647);
xor U4428 (N_4428,N_3888,N_3977);
nor U4429 (N_4429,N_3765,N_3564);
nand U4430 (N_4430,N_3577,N_3818);
nor U4431 (N_4431,N_3610,N_3510);
nand U4432 (N_4432,N_3602,N_3821);
xnor U4433 (N_4433,N_3780,N_3961);
xnor U4434 (N_4434,N_3502,N_3832);
nor U4435 (N_4435,N_3802,N_3635);
nand U4436 (N_4436,N_3938,N_3717);
nand U4437 (N_4437,N_3528,N_3727);
xnor U4438 (N_4438,N_3684,N_3954);
xor U4439 (N_4439,N_3504,N_3631);
or U4440 (N_4440,N_3955,N_3965);
nand U4441 (N_4441,N_3514,N_3596);
nand U4442 (N_4442,N_3810,N_3785);
xnor U4443 (N_4443,N_3627,N_3960);
xor U4444 (N_4444,N_3920,N_3538);
and U4445 (N_4445,N_3685,N_3967);
nor U4446 (N_4446,N_3693,N_3807);
or U4447 (N_4447,N_3695,N_3898);
and U4448 (N_4448,N_3593,N_3765);
or U4449 (N_4449,N_3841,N_3918);
nand U4450 (N_4450,N_3817,N_3880);
or U4451 (N_4451,N_3758,N_3901);
nand U4452 (N_4452,N_3955,N_3609);
and U4453 (N_4453,N_3976,N_3715);
xnor U4454 (N_4454,N_3814,N_3963);
xnor U4455 (N_4455,N_3579,N_3942);
xor U4456 (N_4456,N_3574,N_3561);
or U4457 (N_4457,N_3618,N_3883);
nor U4458 (N_4458,N_3589,N_3898);
nor U4459 (N_4459,N_3565,N_3687);
nor U4460 (N_4460,N_3981,N_3884);
nor U4461 (N_4461,N_3927,N_3697);
and U4462 (N_4462,N_3901,N_3999);
and U4463 (N_4463,N_3687,N_3800);
and U4464 (N_4464,N_3695,N_3509);
and U4465 (N_4465,N_3566,N_3645);
nand U4466 (N_4466,N_3970,N_3707);
or U4467 (N_4467,N_3869,N_3888);
xnor U4468 (N_4468,N_3666,N_3902);
nor U4469 (N_4469,N_3780,N_3918);
and U4470 (N_4470,N_3588,N_3986);
and U4471 (N_4471,N_3657,N_3991);
or U4472 (N_4472,N_3699,N_3841);
nand U4473 (N_4473,N_3783,N_3735);
xnor U4474 (N_4474,N_3737,N_3580);
xnor U4475 (N_4475,N_3595,N_3631);
or U4476 (N_4476,N_3713,N_3622);
xnor U4477 (N_4477,N_3892,N_3772);
xnor U4478 (N_4478,N_3845,N_3961);
or U4479 (N_4479,N_3805,N_3509);
nand U4480 (N_4480,N_3782,N_3503);
xnor U4481 (N_4481,N_3849,N_3935);
and U4482 (N_4482,N_3687,N_3669);
xnor U4483 (N_4483,N_3618,N_3939);
nand U4484 (N_4484,N_3622,N_3573);
or U4485 (N_4485,N_3880,N_3690);
or U4486 (N_4486,N_3544,N_3724);
and U4487 (N_4487,N_3591,N_3661);
nand U4488 (N_4488,N_3843,N_3574);
and U4489 (N_4489,N_3594,N_3697);
nand U4490 (N_4490,N_3690,N_3528);
or U4491 (N_4491,N_3810,N_3986);
xnor U4492 (N_4492,N_3959,N_3965);
nor U4493 (N_4493,N_3935,N_3532);
and U4494 (N_4494,N_3521,N_3838);
nor U4495 (N_4495,N_3736,N_3975);
nand U4496 (N_4496,N_3520,N_3729);
nor U4497 (N_4497,N_3602,N_3656);
and U4498 (N_4498,N_3570,N_3813);
nor U4499 (N_4499,N_3838,N_3733);
xnor U4500 (N_4500,N_4017,N_4051);
or U4501 (N_4501,N_4206,N_4067);
xnor U4502 (N_4502,N_4012,N_4226);
nand U4503 (N_4503,N_4375,N_4100);
and U4504 (N_4504,N_4308,N_4006);
nand U4505 (N_4505,N_4269,N_4315);
or U4506 (N_4506,N_4187,N_4204);
and U4507 (N_4507,N_4013,N_4142);
nand U4508 (N_4508,N_4086,N_4075);
nor U4509 (N_4509,N_4309,N_4121);
nor U4510 (N_4510,N_4177,N_4288);
nor U4511 (N_4511,N_4411,N_4173);
or U4512 (N_4512,N_4267,N_4426);
xnor U4513 (N_4513,N_4373,N_4182);
nor U4514 (N_4514,N_4330,N_4070);
xor U4515 (N_4515,N_4245,N_4359);
nor U4516 (N_4516,N_4088,N_4366);
nor U4517 (N_4517,N_4311,N_4369);
nor U4518 (N_4518,N_4495,N_4171);
and U4519 (N_4519,N_4300,N_4314);
xor U4520 (N_4520,N_4328,N_4413);
or U4521 (N_4521,N_4188,N_4024);
nor U4522 (N_4522,N_4239,N_4072);
and U4523 (N_4523,N_4068,N_4062);
nor U4524 (N_4524,N_4263,N_4224);
nor U4525 (N_4525,N_4140,N_4454);
or U4526 (N_4526,N_4167,N_4053);
or U4527 (N_4527,N_4451,N_4305);
nor U4528 (N_4528,N_4418,N_4014);
and U4529 (N_4529,N_4238,N_4136);
or U4530 (N_4530,N_4194,N_4228);
and U4531 (N_4531,N_4069,N_4223);
and U4532 (N_4532,N_4107,N_4452);
xor U4533 (N_4533,N_4437,N_4444);
nor U4534 (N_4534,N_4307,N_4139);
or U4535 (N_4535,N_4403,N_4443);
xnor U4536 (N_4536,N_4380,N_4487);
xor U4537 (N_4537,N_4360,N_4478);
or U4538 (N_4538,N_4317,N_4496);
nand U4539 (N_4539,N_4423,N_4470);
and U4540 (N_4540,N_4337,N_4011);
or U4541 (N_4541,N_4215,N_4093);
nor U4542 (N_4542,N_4128,N_4271);
nor U4543 (N_4543,N_4483,N_4132);
nor U4544 (N_4544,N_4414,N_4479);
xnor U4545 (N_4545,N_4220,N_4207);
or U4546 (N_4546,N_4202,N_4023);
xnor U4547 (N_4547,N_4196,N_4421);
nand U4548 (N_4548,N_4394,N_4120);
nor U4549 (N_4549,N_4165,N_4218);
nor U4550 (N_4550,N_4250,N_4092);
nand U4551 (N_4551,N_4117,N_4001);
xor U4552 (N_4552,N_4382,N_4335);
nor U4553 (N_4553,N_4404,N_4018);
or U4554 (N_4554,N_4339,N_4231);
or U4555 (N_4555,N_4159,N_4105);
or U4556 (N_4556,N_4243,N_4091);
and U4557 (N_4557,N_4449,N_4417);
nand U4558 (N_4558,N_4321,N_4343);
or U4559 (N_4559,N_4374,N_4276);
nand U4560 (N_4560,N_4219,N_4054);
nor U4561 (N_4561,N_4342,N_4242);
nand U4562 (N_4562,N_4230,N_4189);
xor U4563 (N_4563,N_4032,N_4161);
nor U4564 (N_4564,N_4448,N_4212);
nor U4565 (N_4565,N_4025,N_4410);
nand U4566 (N_4566,N_4358,N_4367);
and U4567 (N_4567,N_4047,N_4131);
and U4568 (N_4568,N_4365,N_4489);
nand U4569 (N_4569,N_4210,N_4026);
xnor U4570 (N_4570,N_4148,N_4334);
nand U4571 (N_4571,N_4457,N_4261);
or U4572 (N_4572,N_4119,N_4232);
xor U4573 (N_4573,N_4313,N_4061);
nand U4574 (N_4574,N_4249,N_4424);
and U4575 (N_4575,N_4370,N_4402);
and U4576 (N_4576,N_4450,N_4278);
and U4577 (N_4577,N_4281,N_4116);
xor U4578 (N_4578,N_4327,N_4420);
nand U4579 (N_4579,N_4262,N_4270);
nor U4580 (N_4580,N_4272,N_4259);
and U4581 (N_4581,N_4453,N_4133);
and U4582 (N_4582,N_4482,N_4429);
xnor U4583 (N_4583,N_4298,N_4038);
and U4584 (N_4584,N_4235,N_4430);
nand U4585 (N_4585,N_4035,N_4466);
nand U4586 (N_4586,N_4246,N_4106);
or U4587 (N_4587,N_4217,N_4055);
nor U4588 (N_4588,N_4279,N_4101);
nand U4589 (N_4589,N_4080,N_4052);
nor U4590 (N_4590,N_4118,N_4033);
xnor U4591 (N_4591,N_4344,N_4265);
or U4592 (N_4592,N_4056,N_4324);
nand U4593 (N_4593,N_4077,N_4178);
or U4594 (N_4594,N_4166,N_4213);
nor U4595 (N_4595,N_4110,N_4493);
or U4596 (N_4596,N_4310,N_4176);
nand U4597 (N_4597,N_4058,N_4458);
or U4598 (N_4598,N_4211,N_4114);
nand U4599 (N_4599,N_4170,N_4323);
nor U4600 (N_4600,N_4233,N_4350);
nand U4601 (N_4601,N_4346,N_4497);
nor U4602 (N_4602,N_4361,N_4192);
nor U4603 (N_4603,N_4280,N_4073);
xnor U4604 (N_4604,N_4152,N_4486);
nand U4605 (N_4605,N_4274,N_4398);
xor U4606 (N_4606,N_4349,N_4000);
and U4607 (N_4607,N_4353,N_4289);
and U4608 (N_4608,N_4151,N_4150);
nand U4609 (N_4609,N_4008,N_4456);
xor U4610 (N_4610,N_4144,N_4090);
xor U4611 (N_4611,N_4010,N_4184);
or U4612 (N_4612,N_4439,N_4419);
nor U4613 (N_4613,N_4352,N_4094);
nor U4614 (N_4614,N_4368,N_4416);
and U4615 (N_4615,N_4009,N_4029);
nor U4616 (N_4616,N_4282,N_4354);
nand U4617 (N_4617,N_4180,N_4492);
xor U4618 (N_4618,N_4490,N_4376);
nand U4619 (N_4619,N_4332,N_4143);
or U4620 (N_4620,N_4391,N_4399);
or U4621 (N_4621,N_4434,N_4294);
xor U4622 (N_4622,N_4351,N_4472);
and U4623 (N_4623,N_4221,N_4147);
xnor U4624 (N_4624,N_4467,N_4113);
nand U4625 (N_4625,N_4169,N_4007);
nor U4626 (N_4626,N_4163,N_4260);
nor U4627 (N_4627,N_4301,N_4195);
and U4628 (N_4628,N_4464,N_4256);
or U4629 (N_4629,N_4155,N_4461);
and U4630 (N_4630,N_4126,N_4021);
nor U4631 (N_4631,N_4469,N_4338);
xnor U4632 (N_4632,N_4129,N_4084);
nand U4633 (N_4633,N_4293,N_4227);
and U4634 (N_4634,N_4463,N_4112);
nand U4635 (N_4635,N_4441,N_4198);
and U4636 (N_4636,N_4157,N_4388);
xnor U4637 (N_4637,N_4040,N_4442);
xnor U4638 (N_4638,N_4225,N_4074);
and U4639 (N_4639,N_4059,N_4401);
and U4640 (N_4640,N_4480,N_4162);
nor U4641 (N_4641,N_4438,N_4409);
xor U4642 (N_4642,N_4076,N_4331);
nor U4643 (N_4643,N_4273,N_4205);
or U4644 (N_4644,N_4048,N_4042);
xor U4645 (N_4645,N_4336,N_4244);
nand U4646 (N_4646,N_4002,N_4115);
or U4647 (N_4647,N_4320,N_4200);
or U4648 (N_4648,N_4499,N_4415);
nand U4649 (N_4649,N_4371,N_4340);
and U4650 (N_4650,N_4085,N_4175);
nand U4651 (N_4651,N_4381,N_4156);
nand U4652 (N_4652,N_4095,N_4099);
xnor U4653 (N_4653,N_4108,N_4494);
xor U4654 (N_4654,N_4397,N_4216);
or U4655 (N_4655,N_4179,N_4193);
nor U4656 (N_4656,N_4462,N_4248);
xor U4657 (N_4657,N_4020,N_4037);
nor U4658 (N_4658,N_4385,N_4459);
or U4659 (N_4659,N_4465,N_4283);
nor U4660 (N_4660,N_4087,N_4304);
xor U4661 (N_4661,N_4476,N_4135);
nor U4662 (N_4662,N_4043,N_4477);
nor U4663 (N_4663,N_4030,N_4446);
nand U4664 (N_4664,N_4146,N_4064);
nor U4665 (N_4665,N_4395,N_4066);
and U4666 (N_4666,N_4378,N_4015);
xor U4667 (N_4667,N_4425,N_4183);
nor U4668 (N_4668,N_4237,N_4318);
and U4669 (N_4669,N_4363,N_4407);
nor U4670 (N_4670,N_4473,N_4109);
nand U4671 (N_4671,N_4364,N_4252);
and U4672 (N_4672,N_4316,N_4333);
and U4673 (N_4673,N_4104,N_4057);
nor U4674 (N_4674,N_4362,N_4191);
xnor U4675 (N_4675,N_4474,N_4172);
or U4676 (N_4676,N_4081,N_4357);
nor U4677 (N_4677,N_4125,N_4181);
nor U4678 (N_4678,N_4266,N_4435);
or U4679 (N_4679,N_4185,N_4285);
xor U4680 (N_4680,N_4275,N_4158);
or U4681 (N_4681,N_4019,N_4297);
nor U4682 (N_4682,N_4400,N_4186);
nor U4683 (N_4683,N_4005,N_4329);
or U4684 (N_4684,N_4386,N_4284);
or U4685 (N_4685,N_4022,N_4138);
or U4686 (N_4686,N_4432,N_4460);
nor U4687 (N_4687,N_4341,N_4379);
nand U4688 (N_4688,N_4290,N_4291);
or U4689 (N_4689,N_4372,N_4050);
nand U4690 (N_4690,N_4436,N_4071);
nor U4691 (N_4691,N_4440,N_4287);
nor U4692 (N_4692,N_4326,N_4199);
nor U4693 (N_4693,N_4063,N_4445);
and U4694 (N_4694,N_4103,N_4392);
nor U4695 (N_4695,N_4471,N_4097);
or U4696 (N_4696,N_4145,N_4137);
xnor U4697 (N_4697,N_4078,N_4234);
and U4698 (N_4698,N_4236,N_4277);
nand U4699 (N_4699,N_4264,N_4447);
xnor U4700 (N_4700,N_4240,N_4154);
nor U4701 (N_4701,N_4422,N_4406);
and U4702 (N_4702,N_4168,N_4396);
xor U4703 (N_4703,N_4488,N_4312);
nor U4704 (N_4704,N_4355,N_4098);
nand U4705 (N_4705,N_4255,N_4468);
or U4706 (N_4706,N_4229,N_4433);
nor U4707 (N_4707,N_4127,N_4498);
and U4708 (N_4708,N_4122,N_4306);
and U4709 (N_4709,N_4102,N_4299);
nand U4710 (N_4710,N_4197,N_4174);
and U4711 (N_4711,N_4491,N_4083);
nand U4712 (N_4712,N_4455,N_4208);
or U4713 (N_4713,N_4079,N_4347);
nor U4714 (N_4714,N_4296,N_4253);
nand U4715 (N_4715,N_4384,N_4427);
and U4716 (N_4716,N_4004,N_4377);
xnor U4717 (N_4717,N_4153,N_4003);
nand U4718 (N_4718,N_4222,N_4412);
nor U4719 (N_4719,N_4484,N_4201);
nor U4720 (N_4720,N_4209,N_4134);
nand U4721 (N_4721,N_4065,N_4475);
nand U4722 (N_4722,N_4303,N_4041);
nand U4723 (N_4723,N_4428,N_4345);
and U4724 (N_4724,N_4481,N_4164);
xnor U4725 (N_4725,N_4258,N_4124);
and U4726 (N_4726,N_4039,N_4387);
or U4727 (N_4727,N_4044,N_4257);
nand U4728 (N_4728,N_4251,N_4348);
nor U4729 (N_4729,N_4027,N_4268);
xor U4730 (N_4730,N_4302,N_4046);
nand U4731 (N_4731,N_4254,N_4082);
and U4732 (N_4732,N_4247,N_4390);
nand U4733 (N_4733,N_4203,N_4130);
nand U4734 (N_4734,N_4319,N_4241);
nor U4735 (N_4735,N_4111,N_4393);
nor U4736 (N_4736,N_4089,N_4031);
and U4737 (N_4737,N_4034,N_4016);
nand U4738 (N_4738,N_4405,N_4160);
and U4739 (N_4739,N_4123,N_4389);
or U4740 (N_4740,N_4431,N_4286);
or U4741 (N_4741,N_4096,N_4036);
and U4742 (N_4742,N_4292,N_4028);
nand U4743 (N_4743,N_4214,N_4295);
nand U4744 (N_4744,N_4408,N_4149);
or U4745 (N_4745,N_4383,N_4356);
or U4746 (N_4746,N_4325,N_4190);
nand U4747 (N_4747,N_4485,N_4049);
or U4748 (N_4748,N_4322,N_4141);
xnor U4749 (N_4749,N_4045,N_4060);
nor U4750 (N_4750,N_4221,N_4212);
and U4751 (N_4751,N_4168,N_4199);
nor U4752 (N_4752,N_4084,N_4103);
nand U4753 (N_4753,N_4180,N_4133);
nand U4754 (N_4754,N_4404,N_4133);
nor U4755 (N_4755,N_4162,N_4096);
or U4756 (N_4756,N_4267,N_4009);
and U4757 (N_4757,N_4307,N_4427);
nand U4758 (N_4758,N_4029,N_4190);
or U4759 (N_4759,N_4022,N_4241);
or U4760 (N_4760,N_4060,N_4447);
xor U4761 (N_4761,N_4209,N_4401);
nor U4762 (N_4762,N_4070,N_4344);
nand U4763 (N_4763,N_4286,N_4002);
and U4764 (N_4764,N_4365,N_4140);
xor U4765 (N_4765,N_4379,N_4478);
xnor U4766 (N_4766,N_4008,N_4278);
nand U4767 (N_4767,N_4108,N_4175);
xor U4768 (N_4768,N_4348,N_4147);
nor U4769 (N_4769,N_4063,N_4370);
and U4770 (N_4770,N_4483,N_4164);
nand U4771 (N_4771,N_4330,N_4226);
or U4772 (N_4772,N_4439,N_4434);
and U4773 (N_4773,N_4073,N_4288);
nor U4774 (N_4774,N_4231,N_4027);
nand U4775 (N_4775,N_4263,N_4415);
nand U4776 (N_4776,N_4354,N_4230);
xor U4777 (N_4777,N_4276,N_4210);
or U4778 (N_4778,N_4229,N_4411);
or U4779 (N_4779,N_4417,N_4034);
xor U4780 (N_4780,N_4125,N_4275);
xnor U4781 (N_4781,N_4474,N_4367);
nor U4782 (N_4782,N_4460,N_4379);
or U4783 (N_4783,N_4415,N_4056);
nor U4784 (N_4784,N_4358,N_4010);
nand U4785 (N_4785,N_4316,N_4454);
or U4786 (N_4786,N_4485,N_4457);
or U4787 (N_4787,N_4103,N_4393);
xnor U4788 (N_4788,N_4466,N_4096);
or U4789 (N_4789,N_4489,N_4434);
nand U4790 (N_4790,N_4303,N_4142);
and U4791 (N_4791,N_4184,N_4498);
xor U4792 (N_4792,N_4248,N_4334);
nand U4793 (N_4793,N_4494,N_4472);
xor U4794 (N_4794,N_4010,N_4193);
and U4795 (N_4795,N_4334,N_4310);
nor U4796 (N_4796,N_4118,N_4318);
and U4797 (N_4797,N_4090,N_4377);
nand U4798 (N_4798,N_4078,N_4143);
nand U4799 (N_4799,N_4032,N_4273);
nor U4800 (N_4800,N_4123,N_4260);
nor U4801 (N_4801,N_4395,N_4389);
nor U4802 (N_4802,N_4101,N_4162);
xor U4803 (N_4803,N_4385,N_4172);
and U4804 (N_4804,N_4203,N_4317);
xnor U4805 (N_4805,N_4113,N_4361);
nor U4806 (N_4806,N_4340,N_4224);
nand U4807 (N_4807,N_4008,N_4095);
nand U4808 (N_4808,N_4044,N_4224);
nor U4809 (N_4809,N_4469,N_4104);
or U4810 (N_4810,N_4388,N_4192);
or U4811 (N_4811,N_4417,N_4153);
or U4812 (N_4812,N_4004,N_4286);
nand U4813 (N_4813,N_4173,N_4372);
and U4814 (N_4814,N_4434,N_4252);
and U4815 (N_4815,N_4119,N_4091);
and U4816 (N_4816,N_4080,N_4171);
or U4817 (N_4817,N_4446,N_4190);
and U4818 (N_4818,N_4160,N_4110);
or U4819 (N_4819,N_4012,N_4164);
and U4820 (N_4820,N_4272,N_4257);
or U4821 (N_4821,N_4268,N_4366);
nand U4822 (N_4822,N_4386,N_4090);
nor U4823 (N_4823,N_4360,N_4036);
nor U4824 (N_4824,N_4395,N_4469);
or U4825 (N_4825,N_4193,N_4178);
xor U4826 (N_4826,N_4420,N_4407);
and U4827 (N_4827,N_4457,N_4181);
nand U4828 (N_4828,N_4054,N_4327);
or U4829 (N_4829,N_4037,N_4090);
nand U4830 (N_4830,N_4366,N_4328);
xor U4831 (N_4831,N_4131,N_4472);
or U4832 (N_4832,N_4113,N_4237);
nand U4833 (N_4833,N_4162,N_4152);
nor U4834 (N_4834,N_4309,N_4352);
and U4835 (N_4835,N_4329,N_4111);
nand U4836 (N_4836,N_4008,N_4390);
nor U4837 (N_4837,N_4232,N_4252);
nor U4838 (N_4838,N_4088,N_4279);
nand U4839 (N_4839,N_4271,N_4015);
or U4840 (N_4840,N_4073,N_4158);
or U4841 (N_4841,N_4429,N_4045);
nand U4842 (N_4842,N_4120,N_4141);
nor U4843 (N_4843,N_4080,N_4346);
xnor U4844 (N_4844,N_4374,N_4444);
nand U4845 (N_4845,N_4440,N_4029);
xor U4846 (N_4846,N_4307,N_4230);
nand U4847 (N_4847,N_4247,N_4072);
nor U4848 (N_4848,N_4148,N_4300);
xor U4849 (N_4849,N_4389,N_4209);
xnor U4850 (N_4850,N_4405,N_4397);
xor U4851 (N_4851,N_4270,N_4453);
xnor U4852 (N_4852,N_4294,N_4297);
nor U4853 (N_4853,N_4302,N_4179);
nor U4854 (N_4854,N_4395,N_4219);
and U4855 (N_4855,N_4426,N_4430);
nand U4856 (N_4856,N_4406,N_4069);
nor U4857 (N_4857,N_4101,N_4377);
and U4858 (N_4858,N_4257,N_4013);
and U4859 (N_4859,N_4246,N_4019);
or U4860 (N_4860,N_4089,N_4245);
and U4861 (N_4861,N_4165,N_4041);
or U4862 (N_4862,N_4302,N_4432);
or U4863 (N_4863,N_4308,N_4485);
and U4864 (N_4864,N_4358,N_4339);
nor U4865 (N_4865,N_4255,N_4254);
nand U4866 (N_4866,N_4396,N_4472);
or U4867 (N_4867,N_4329,N_4238);
nor U4868 (N_4868,N_4256,N_4367);
and U4869 (N_4869,N_4453,N_4187);
xor U4870 (N_4870,N_4315,N_4431);
or U4871 (N_4871,N_4483,N_4155);
or U4872 (N_4872,N_4030,N_4200);
nor U4873 (N_4873,N_4225,N_4286);
and U4874 (N_4874,N_4018,N_4068);
and U4875 (N_4875,N_4374,N_4118);
or U4876 (N_4876,N_4445,N_4360);
nand U4877 (N_4877,N_4002,N_4328);
nor U4878 (N_4878,N_4409,N_4389);
and U4879 (N_4879,N_4370,N_4064);
and U4880 (N_4880,N_4140,N_4033);
xnor U4881 (N_4881,N_4418,N_4063);
nand U4882 (N_4882,N_4436,N_4488);
or U4883 (N_4883,N_4459,N_4212);
nand U4884 (N_4884,N_4443,N_4020);
nor U4885 (N_4885,N_4081,N_4184);
and U4886 (N_4886,N_4205,N_4008);
nand U4887 (N_4887,N_4489,N_4403);
nor U4888 (N_4888,N_4231,N_4260);
nand U4889 (N_4889,N_4497,N_4440);
or U4890 (N_4890,N_4280,N_4242);
nor U4891 (N_4891,N_4251,N_4097);
xnor U4892 (N_4892,N_4271,N_4277);
or U4893 (N_4893,N_4039,N_4480);
and U4894 (N_4894,N_4373,N_4068);
xnor U4895 (N_4895,N_4292,N_4096);
nand U4896 (N_4896,N_4081,N_4008);
and U4897 (N_4897,N_4112,N_4167);
or U4898 (N_4898,N_4010,N_4348);
nand U4899 (N_4899,N_4310,N_4190);
xor U4900 (N_4900,N_4294,N_4249);
nand U4901 (N_4901,N_4446,N_4047);
nand U4902 (N_4902,N_4205,N_4247);
nor U4903 (N_4903,N_4148,N_4458);
nor U4904 (N_4904,N_4127,N_4481);
and U4905 (N_4905,N_4247,N_4094);
or U4906 (N_4906,N_4310,N_4339);
or U4907 (N_4907,N_4264,N_4304);
or U4908 (N_4908,N_4484,N_4067);
or U4909 (N_4909,N_4161,N_4327);
xnor U4910 (N_4910,N_4019,N_4487);
or U4911 (N_4911,N_4052,N_4179);
or U4912 (N_4912,N_4013,N_4062);
nand U4913 (N_4913,N_4094,N_4452);
xnor U4914 (N_4914,N_4491,N_4379);
and U4915 (N_4915,N_4231,N_4457);
and U4916 (N_4916,N_4083,N_4241);
and U4917 (N_4917,N_4007,N_4025);
or U4918 (N_4918,N_4092,N_4161);
or U4919 (N_4919,N_4122,N_4031);
or U4920 (N_4920,N_4236,N_4211);
or U4921 (N_4921,N_4319,N_4238);
or U4922 (N_4922,N_4469,N_4303);
or U4923 (N_4923,N_4057,N_4000);
or U4924 (N_4924,N_4122,N_4324);
and U4925 (N_4925,N_4377,N_4485);
or U4926 (N_4926,N_4497,N_4199);
and U4927 (N_4927,N_4461,N_4315);
nand U4928 (N_4928,N_4295,N_4004);
or U4929 (N_4929,N_4301,N_4108);
nor U4930 (N_4930,N_4436,N_4252);
xnor U4931 (N_4931,N_4357,N_4175);
xnor U4932 (N_4932,N_4099,N_4474);
xnor U4933 (N_4933,N_4130,N_4122);
nand U4934 (N_4934,N_4146,N_4357);
or U4935 (N_4935,N_4441,N_4489);
or U4936 (N_4936,N_4483,N_4339);
nor U4937 (N_4937,N_4374,N_4418);
nor U4938 (N_4938,N_4013,N_4191);
and U4939 (N_4939,N_4383,N_4466);
nor U4940 (N_4940,N_4465,N_4126);
nor U4941 (N_4941,N_4140,N_4430);
xnor U4942 (N_4942,N_4053,N_4433);
nand U4943 (N_4943,N_4078,N_4474);
nor U4944 (N_4944,N_4277,N_4242);
nand U4945 (N_4945,N_4280,N_4032);
nor U4946 (N_4946,N_4231,N_4056);
or U4947 (N_4947,N_4098,N_4050);
nand U4948 (N_4948,N_4229,N_4363);
and U4949 (N_4949,N_4003,N_4330);
or U4950 (N_4950,N_4279,N_4428);
nor U4951 (N_4951,N_4331,N_4340);
or U4952 (N_4952,N_4298,N_4082);
nor U4953 (N_4953,N_4482,N_4412);
nand U4954 (N_4954,N_4479,N_4424);
and U4955 (N_4955,N_4054,N_4089);
xnor U4956 (N_4956,N_4448,N_4159);
nand U4957 (N_4957,N_4362,N_4248);
xor U4958 (N_4958,N_4054,N_4034);
and U4959 (N_4959,N_4325,N_4155);
or U4960 (N_4960,N_4037,N_4112);
nor U4961 (N_4961,N_4133,N_4245);
or U4962 (N_4962,N_4219,N_4020);
or U4963 (N_4963,N_4104,N_4298);
and U4964 (N_4964,N_4253,N_4429);
xor U4965 (N_4965,N_4354,N_4358);
xnor U4966 (N_4966,N_4436,N_4158);
and U4967 (N_4967,N_4464,N_4242);
xnor U4968 (N_4968,N_4153,N_4331);
xnor U4969 (N_4969,N_4176,N_4343);
or U4970 (N_4970,N_4272,N_4049);
nor U4971 (N_4971,N_4108,N_4249);
nand U4972 (N_4972,N_4342,N_4051);
nand U4973 (N_4973,N_4430,N_4264);
nand U4974 (N_4974,N_4296,N_4408);
or U4975 (N_4975,N_4317,N_4022);
or U4976 (N_4976,N_4187,N_4359);
or U4977 (N_4977,N_4003,N_4234);
or U4978 (N_4978,N_4499,N_4233);
or U4979 (N_4979,N_4170,N_4134);
nand U4980 (N_4980,N_4266,N_4402);
nand U4981 (N_4981,N_4222,N_4405);
nand U4982 (N_4982,N_4107,N_4058);
nand U4983 (N_4983,N_4419,N_4078);
nand U4984 (N_4984,N_4366,N_4234);
or U4985 (N_4985,N_4252,N_4353);
nor U4986 (N_4986,N_4297,N_4147);
nor U4987 (N_4987,N_4472,N_4124);
or U4988 (N_4988,N_4226,N_4178);
xor U4989 (N_4989,N_4202,N_4312);
and U4990 (N_4990,N_4118,N_4272);
nand U4991 (N_4991,N_4250,N_4144);
nor U4992 (N_4992,N_4224,N_4439);
or U4993 (N_4993,N_4014,N_4383);
nor U4994 (N_4994,N_4206,N_4313);
or U4995 (N_4995,N_4163,N_4246);
nand U4996 (N_4996,N_4212,N_4023);
and U4997 (N_4997,N_4092,N_4451);
and U4998 (N_4998,N_4151,N_4429);
and U4999 (N_4999,N_4238,N_4012);
and U5000 (N_5000,N_4640,N_4718);
or U5001 (N_5001,N_4649,N_4800);
nand U5002 (N_5002,N_4513,N_4545);
xnor U5003 (N_5003,N_4654,N_4760);
nand U5004 (N_5004,N_4607,N_4602);
and U5005 (N_5005,N_4621,N_4971);
nor U5006 (N_5006,N_4542,N_4966);
and U5007 (N_5007,N_4989,N_4773);
or U5008 (N_5008,N_4574,N_4864);
nand U5009 (N_5009,N_4777,N_4944);
nand U5010 (N_5010,N_4518,N_4772);
nand U5011 (N_5011,N_4550,N_4529);
or U5012 (N_5012,N_4844,N_4949);
and U5013 (N_5013,N_4778,N_4852);
or U5014 (N_5014,N_4657,N_4715);
or U5015 (N_5015,N_4661,N_4551);
xnor U5016 (N_5016,N_4722,N_4911);
nor U5017 (N_5017,N_4616,N_4546);
xor U5018 (N_5018,N_4538,N_4857);
xor U5019 (N_5019,N_4978,N_4660);
or U5020 (N_5020,N_4577,N_4957);
and U5021 (N_5021,N_4779,N_4558);
or U5022 (N_5022,N_4817,N_4757);
nand U5023 (N_5023,N_4974,N_4797);
nor U5024 (N_5024,N_4848,N_4633);
nand U5025 (N_5025,N_4963,N_4882);
xnor U5026 (N_5026,N_4643,N_4625);
nand U5027 (N_5027,N_4664,N_4548);
nand U5028 (N_5028,N_4587,N_4886);
or U5029 (N_5029,N_4935,N_4884);
xor U5030 (N_5030,N_4940,N_4980);
xor U5031 (N_5031,N_4680,N_4759);
xnor U5032 (N_5032,N_4557,N_4975);
nor U5033 (N_5033,N_4601,N_4766);
nor U5034 (N_5034,N_4860,N_4917);
or U5035 (N_5035,N_4690,N_4893);
and U5036 (N_5036,N_4798,N_4856);
and U5037 (N_5037,N_4736,N_4863);
nand U5038 (N_5038,N_4555,N_4571);
or U5039 (N_5039,N_4704,N_4630);
xor U5040 (N_5040,N_4977,N_4885);
or U5041 (N_5041,N_4794,N_4818);
and U5042 (N_5042,N_4527,N_4990);
nand U5043 (N_5043,N_4628,N_4849);
nand U5044 (N_5044,N_4727,N_4645);
and U5045 (N_5045,N_4941,N_4682);
xnor U5046 (N_5046,N_4994,N_4728);
nor U5047 (N_5047,N_4908,N_4522);
and U5048 (N_5048,N_4540,N_4676);
nand U5049 (N_5049,N_4827,N_4929);
or U5050 (N_5050,N_4892,N_4952);
xor U5051 (N_5051,N_4776,N_4973);
or U5052 (N_5052,N_4932,N_4739);
nand U5053 (N_5053,N_4784,N_4795);
nand U5054 (N_5054,N_4667,N_4562);
nor U5055 (N_5055,N_4655,N_4516);
nand U5056 (N_5056,N_4641,N_4585);
and U5057 (N_5057,N_4726,N_4854);
or U5058 (N_5058,N_4716,N_4679);
xor U5059 (N_5059,N_4501,N_4956);
nor U5060 (N_5060,N_4737,N_4568);
nor U5061 (N_5061,N_4702,N_4638);
and U5062 (N_5062,N_4671,N_4626);
or U5063 (N_5063,N_4830,N_4572);
xor U5064 (N_5064,N_4543,N_4821);
nor U5065 (N_5065,N_4693,N_4532);
nand U5066 (N_5066,N_4811,N_4976);
or U5067 (N_5067,N_4672,N_4711);
and U5068 (N_5068,N_4582,N_4687);
and U5069 (N_5069,N_4517,N_4662);
xor U5070 (N_5070,N_4559,N_4874);
nor U5071 (N_5071,N_4951,N_4822);
and U5072 (N_5072,N_4781,N_4719);
and U5073 (N_5073,N_4926,N_4521);
and U5074 (N_5074,N_4697,N_4890);
nor U5075 (N_5075,N_4696,N_4708);
xnor U5076 (N_5076,N_4899,N_4705);
or U5077 (N_5077,N_4820,N_4945);
nor U5078 (N_5078,N_4933,N_4510);
or U5079 (N_5079,N_4898,N_4701);
nand U5080 (N_5080,N_4507,N_4534);
nand U5081 (N_5081,N_4786,N_4775);
or U5082 (N_5082,N_4544,N_4868);
nor U5083 (N_5083,N_4912,N_4783);
nor U5084 (N_5084,N_4596,N_4919);
xor U5085 (N_5085,N_4694,N_4599);
nor U5086 (N_5086,N_4564,N_4803);
nand U5087 (N_5087,N_4888,N_4560);
nand U5088 (N_5088,N_4825,N_4724);
xnor U5089 (N_5089,N_4717,N_4823);
nand U5090 (N_5090,N_4734,N_4629);
nand U5091 (N_5091,N_4814,N_4554);
and U5092 (N_5092,N_4648,N_4593);
and U5093 (N_5093,N_4646,N_4962);
nor U5094 (N_5094,N_4598,N_4921);
and U5095 (N_5095,N_4519,N_4749);
xnor U5096 (N_5096,N_4509,N_4580);
nand U5097 (N_5097,N_4604,N_4605);
nor U5098 (N_5098,N_4878,N_4806);
nor U5099 (N_5099,N_4731,N_4525);
nor U5100 (N_5100,N_4665,N_4647);
and U5101 (N_5101,N_4829,N_4746);
nor U5102 (N_5102,N_4905,N_4793);
or U5103 (N_5103,N_4553,N_4758);
or U5104 (N_5104,N_4824,N_4922);
and U5105 (N_5105,N_4549,N_4755);
or U5106 (N_5106,N_4618,N_4901);
xnor U5107 (N_5107,N_4608,N_4653);
and U5108 (N_5108,N_4565,N_4541);
xnor U5109 (N_5109,N_4903,N_4624);
or U5110 (N_5110,N_4762,N_4658);
nand U5111 (N_5111,N_4867,N_4981);
xnor U5112 (N_5112,N_4812,N_4635);
xor U5113 (N_5113,N_4918,N_4502);
and U5114 (N_5114,N_4859,N_4740);
nor U5115 (N_5115,N_4833,N_4879);
and U5116 (N_5116,N_4907,N_4897);
nor U5117 (N_5117,N_4505,N_4865);
nand U5118 (N_5118,N_4733,N_4896);
and U5119 (N_5119,N_4927,N_4575);
or U5120 (N_5120,N_4928,N_4637);
or U5121 (N_5121,N_4620,N_4799);
xnor U5122 (N_5122,N_4858,N_4556);
and U5123 (N_5123,N_4894,N_4953);
and U5124 (N_5124,N_4531,N_4984);
xor U5125 (N_5125,N_4887,N_4998);
xor U5126 (N_5126,N_4750,N_4752);
nand U5127 (N_5127,N_4508,N_4828);
nor U5128 (N_5128,N_4906,N_4670);
nor U5129 (N_5129,N_4579,N_4881);
or U5130 (N_5130,N_4735,N_4843);
nor U5131 (N_5131,N_4997,N_4815);
xnor U5132 (N_5132,N_4732,N_4685);
or U5133 (N_5133,N_4700,N_4594);
or U5134 (N_5134,N_4652,N_4695);
and U5135 (N_5135,N_4802,N_4603);
nand U5136 (N_5136,N_4526,N_4774);
nand U5137 (N_5137,N_4769,N_4872);
nor U5138 (N_5138,N_4831,N_4677);
or U5139 (N_5139,N_4841,N_4561);
or U5140 (N_5140,N_4850,N_4925);
nor U5141 (N_5141,N_4835,N_4663);
nand U5142 (N_5142,N_4613,N_4832);
nor U5143 (N_5143,N_4668,N_4612);
and U5144 (N_5144,N_4714,N_4656);
nor U5145 (N_5145,N_4651,N_4623);
nand U5146 (N_5146,N_4983,N_4745);
nor U5147 (N_5147,N_4744,N_4987);
xnor U5148 (N_5148,N_4808,N_4581);
or U5149 (N_5149,N_4816,N_4563);
and U5150 (N_5150,N_4590,N_4909);
xnor U5151 (N_5151,N_4567,N_4875);
nor U5152 (N_5152,N_4788,N_4611);
xor U5153 (N_5153,N_4606,N_4876);
nand U5154 (N_5154,N_4790,N_4960);
xnor U5155 (N_5155,N_4834,N_4851);
nand U5156 (N_5156,N_4920,N_4782);
nand U5157 (N_5157,N_4995,N_4780);
or U5158 (N_5158,N_4871,N_4609);
xnor U5159 (N_5159,N_4877,N_4619);
xor U5160 (N_5160,N_4883,N_4725);
nor U5161 (N_5161,N_4615,N_4805);
or U5162 (N_5162,N_4855,N_4991);
and U5163 (N_5163,N_4692,N_4504);
nor U5164 (N_5164,N_4937,N_4523);
and U5165 (N_5165,N_4669,N_4709);
nor U5166 (N_5166,N_4889,N_4589);
xnor U5167 (N_5167,N_4578,N_4847);
xnor U5168 (N_5168,N_4636,N_4916);
nand U5169 (N_5169,N_4576,N_4934);
xnor U5170 (N_5170,N_4853,N_4913);
nor U5171 (N_5171,N_4979,N_4970);
or U5172 (N_5172,N_4570,N_4747);
or U5173 (N_5173,N_4533,N_4678);
nand U5174 (N_5174,N_4915,N_4684);
xor U5175 (N_5175,N_4787,N_4809);
and U5176 (N_5176,N_4699,N_4836);
and U5177 (N_5177,N_4520,N_4552);
or U5178 (N_5178,N_4535,N_4753);
nor U5179 (N_5179,N_4595,N_4845);
or U5180 (N_5180,N_4955,N_4703);
and U5181 (N_5181,N_4985,N_4767);
or U5182 (N_5182,N_4796,N_4791);
and U5183 (N_5183,N_4614,N_4583);
or U5184 (N_5184,N_4768,N_4675);
and U5185 (N_5185,N_4964,N_4710);
nand U5186 (N_5186,N_4939,N_4756);
nor U5187 (N_5187,N_4943,N_4738);
or U5188 (N_5188,N_4988,N_4807);
or U5189 (N_5189,N_4547,N_4754);
or U5190 (N_5190,N_4720,N_4634);
xnor U5191 (N_5191,N_4792,N_4958);
nor U5192 (N_5192,N_4683,N_4999);
and U5193 (N_5193,N_4511,N_4761);
nor U5194 (N_5194,N_4959,N_4610);
or U5195 (N_5195,N_4763,N_4723);
nand U5196 (N_5196,N_4537,N_4873);
and U5197 (N_5197,N_4968,N_4642);
nor U5198 (N_5198,N_4539,N_4967);
xnor U5199 (N_5199,N_4826,N_4961);
nand U5200 (N_5200,N_4942,N_4528);
and U5201 (N_5201,N_4515,N_4804);
and U5202 (N_5202,N_4617,N_4673);
or U5203 (N_5203,N_4741,N_4586);
nand U5204 (N_5204,N_4644,N_4721);
or U5205 (N_5205,N_4904,N_4712);
and U5206 (N_5206,N_4837,N_4659);
and U5207 (N_5207,N_4946,N_4992);
nor U5208 (N_5208,N_4742,N_4842);
or U5209 (N_5209,N_4713,N_4627);
or U5210 (N_5210,N_4691,N_4938);
and U5211 (N_5211,N_4530,N_4923);
nand U5212 (N_5212,N_4972,N_4764);
xnor U5213 (N_5213,N_4503,N_4506);
nand U5214 (N_5214,N_4666,N_4839);
or U5215 (N_5215,N_4982,N_4771);
nor U5216 (N_5216,N_4986,N_4914);
nand U5217 (N_5217,N_4639,N_4588);
nor U5218 (N_5218,N_4930,N_4900);
or U5219 (N_5219,N_4948,N_4765);
xnor U5220 (N_5220,N_4674,N_4631);
or U5221 (N_5221,N_4566,N_4748);
xor U5222 (N_5222,N_4751,N_4969);
nor U5223 (N_5223,N_4870,N_4632);
nor U5224 (N_5224,N_4869,N_4846);
nand U5225 (N_5225,N_4698,N_4686);
nor U5226 (N_5226,N_4838,N_4861);
xor U5227 (N_5227,N_4597,N_4895);
nand U5228 (N_5228,N_4512,N_4810);
and U5229 (N_5229,N_4785,N_4965);
nor U5230 (N_5230,N_4947,N_4743);
xor U5231 (N_5231,N_4840,N_4500);
nand U5232 (N_5232,N_4729,N_4569);
nand U5233 (N_5233,N_4592,N_4688);
nand U5234 (N_5234,N_4880,N_4689);
xnor U5235 (N_5235,N_4707,N_4891);
and U5236 (N_5236,N_4706,N_4996);
nor U5237 (N_5237,N_4524,N_4622);
and U5238 (N_5238,N_4931,N_4954);
xor U5239 (N_5239,N_4730,N_4514);
and U5240 (N_5240,N_4993,N_4573);
nor U5241 (N_5241,N_4910,N_4950);
and U5242 (N_5242,N_4902,N_4770);
nand U5243 (N_5243,N_4681,N_4600);
xnor U5244 (N_5244,N_4650,N_4819);
and U5245 (N_5245,N_4591,N_4584);
and U5246 (N_5246,N_4936,N_4789);
nor U5247 (N_5247,N_4924,N_4801);
xor U5248 (N_5248,N_4862,N_4536);
or U5249 (N_5249,N_4813,N_4866);
nand U5250 (N_5250,N_4769,N_4681);
nand U5251 (N_5251,N_4650,N_4866);
nand U5252 (N_5252,N_4566,N_4619);
nand U5253 (N_5253,N_4552,N_4835);
xor U5254 (N_5254,N_4698,N_4961);
or U5255 (N_5255,N_4540,N_4523);
nor U5256 (N_5256,N_4751,N_4578);
nand U5257 (N_5257,N_4734,N_4702);
xnor U5258 (N_5258,N_4877,N_4851);
nand U5259 (N_5259,N_4882,N_4753);
and U5260 (N_5260,N_4741,N_4585);
nor U5261 (N_5261,N_4516,N_4689);
nor U5262 (N_5262,N_4804,N_4637);
and U5263 (N_5263,N_4637,N_4650);
xor U5264 (N_5264,N_4564,N_4720);
or U5265 (N_5265,N_4971,N_4806);
nor U5266 (N_5266,N_4845,N_4763);
nor U5267 (N_5267,N_4900,N_4813);
xnor U5268 (N_5268,N_4642,N_4557);
nor U5269 (N_5269,N_4770,N_4828);
and U5270 (N_5270,N_4566,N_4768);
nand U5271 (N_5271,N_4580,N_4626);
xnor U5272 (N_5272,N_4828,N_4604);
nand U5273 (N_5273,N_4558,N_4795);
and U5274 (N_5274,N_4686,N_4970);
and U5275 (N_5275,N_4925,N_4936);
and U5276 (N_5276,N_4665,N_4538);
xnor U5277 (N_5277,N_4617,N_4905);
and U5278 (N_5278,N_4805,N_4747);
xor U5279 (N_5279,N_4960,N_4535);
or U5280 (N_5280,N_4644,N_4769);
xnor U5281 (N_5281,N_4857,N_4856);
nand U5282 (N_5282,N_4780,N_4936);
nor U5283 (N_5283,N_4708,N_4760);
and U5284 (N_5284,N_4571,N_4789);
nand U5285 (N_5285,N_4611,N_4509);
xor U5286 (N_5286,N_4747,N_4563);
and U5287 (N_5287,N_4854,N_4849);
and U5288 (N_5288,N_4613,N_4977);
nor U5289 (N_5289,N_4969,N_4706);
nor U5290 (N_5290,N_4905,N_4613);
and U5291 (N_5291,N_4911,N_4577);
nor U5292 (N_5292,N_4752,N_4961);
xor U5293 (N_5293,N_4896,N_4635);
xor U5294 (N_5294,N_4895,N_4632);
xor U5295 (N_5295,N_4746,N_4544);
nand U5296 (N_5296,N_4666,N_4750);
or U5297 (N_5297,N_4836,N_4819);
and U5298 (N_5298,N_4682,N_4912);
or U5299 (N_5299,N_4601,N_4889);
and U5300 (N_5300,N_4755,N_4655);
xor U5301 (N_5301,N_4822,N_4872);
or U5302 (N_5302,N_4861,N_4679);
nand U5303 (N_5303,N_4620,N_4889);
nand U5304 (N_5304,N_4750,N_4894);
xnor U5305 (N_5305,N_4714,N_4540);
nor U5306 (N_5306,N_4851,N_4678);
or U5307 (N_5307,N_4576,N_4584);
nand U5308 (N_5308,N_4781,N_4799);
nor U5309 (N_5309,N_4688,N_4766);
xor U5310 (N_5310,N_4516,N_4730);
and U5311 (N_5311,N_4954,N_4852);
and U5312 (N_5312,N_4621,N_4510);
and U5313 (N_5313,N_4720,N_4547);
or U5314 (N_5314,N_4825,N_4836);
nand U5315 (N_5315,N_4596,N_4850);
xnor U5316 (N_5316,N_4824,N_4690);
nor U5317 (N_5317,N_4637,N_4777);
xnor U5318 (N_5318,N_4785,N_4614);
and U5319 (N_5319,N_4769,N_4863);
nor U5320 (N_5320,N_4867,N_4962);
or U5321 (N_5321,N_4635,N_4734);
or U5322 (N_5322,N_4993,N_4844);
and U5323 (N_5323,N_4805,N_4773);
or U5324 (N_5324,N_4937,N_4588);
and U5325 (N_5325,N_4994,N_4548);
nor U5326 (N_5326,N_4777,N_4788);
xnor U5327 (N_5327,N_4503,N_4533);
and U5328 (N_5328,N_4863,N_4696);
xnor U5329 (N_5329,N_4829,N_4832);
or U5330 (N_5330,N_4913,N_4563);
nor U5331 (N_5331,N_4607,N_4686);
nand U5332 (N_5332,N_4988,N_4981);
nand U5333 (N_5333,N_4888,N_4951);
nor U5334 (N_5334,N_4878,N_4789);
xnor U5335 (N_5335,N_4795,N_4863);
or U5336 (N_5336,N_4508,N_4584);
nor U5337 (N_5337,N_4556,N_4586);
nor U5338 (N_5338,N_4647,N_4839);
and U5339 (N_5339,N_4764,N_4746);
xor U5340 (N_5340,N_4778,N_4954);
nor U5341 (N_5341,N_4847,N_4701);
xnor U5342 (N_5342,N_4672,N_4596);
nand U5343 (N_5343,N_4935,N_4803);
xnor U5344 (N_5344,N_4815,N_4673);
nor U5345 (N_5345,N_4630,N_4841);
xnor U5346 (N_5346,N_4628,N_4873);
nor U5347 (N_5347,N_4649,N_4996);
or U5348 (N_5348,N_4551,N_4973);
nor U5349 (N_5349,N_4568,N_4957);
or U5350 (N_5350,N_4974,N_4937);
and U5351 (N_5351,N_4591,N_4542);
and U5352 (N_5352,N_4594,N_4603);
nor U5353 (N_5353,N_4610,N_4504);
nand U5354 (N_5354,N_4514,N_4841);
nor U5355 (N_5355,N_4945,N_4509);
xnor U5356 (N_5356,N_4500,N_4863);
nor U5357 (N_5357,N_4500,N_4849);
or U5358 (N_5358,N_4988,N_4649);
nor U5359 (N_5359,N_4968,N_4841);
and U5360 (N_5360,N_4933,N_4582);
xnor U5361 (N_5361,N_4734,N_4536);
xor U5362 (N_5362,N_4626,N_4628);
or U5363 (N_5363,N_4881,N_4627);
or U5364 (N_5364,N_4720,N_4814);
and U5365 (N_5365,N_4880,N_4749);
xnor U5366 (N_5366,N_4593,N_4987);
and U5367 (N_5367,N_4618,N_4635);
xnor U5368 (N_5368,N_4959,N_4722);
xnor U5369 (N_5369,N_4981,N_4718);
nor U5370 (N_5370,N_4926,N_4779);
and U5371 (N_5371,N_4515,N_4855);
nand U5372 (N_5372,N_4842,N_4802);
or U5373 (N_5373,N_4615,N_4655);
and U5374 (N_5374,N_4506,N_4910);
or U5375 (N_5375,N_4619,N_4978);
or U5376 (N_5376,N_4559,N_4814);
or U5377 (N_5377,N_4679,N_4629);
nand U5378 (N_5378,N_4815,N_4545);
or U5379 (N_5379,N_4732,N_4618);
nand U5380 (N_5380,N_4596,N_4629);
nand U5381 (N_5381,N_4612,N_4911);
nor U5382 (N_5382,N_4515,N_4924);
and U5383 (N_5383,N_4505,N_4693);
xnor U5384 (N_5384,N_4851,N_4549);
and U5385 (N_5385,N_4676,N_4721);
xnor U5386 (N_5386,N_4775,N_4895);
nor U5387 (N_5387,N_4902,N_4693);
nand U5388 (N_5388,N_4682,N_4543);
nor U5389 (N_5389,N_4551,N_4731);
nand U5390 (N_5390,N_4575,N_4924);
xor U5391 (N_5391,N_4643,N_4766);
and U5392 (N_5392,N_4970,N_4539);
or U5393 (N_5393,N_4891,N_4509);
nor U5394 (N_5394,N_4881,N_4860);
or U5395 (N_5395,N_4570,N_4826);
or U5396 (N_5396,N_4993,N_4744);
and U5397 (N_5397,N_4512,N_4890);
xor U5398 (N_5398,N_4886,N_4658);
nand U5399 (N_5399,N_4625,N_4822);
nor U5400 (N_5400,N_4578,N_4716);
or U5401 (N_5401,N_4953,N_4815);
or U5402 (N_5402,N_4829,N_4721);
or U5403 (N_5403,N_4897,N_4964);
or U5404 (N_5404,N_4524,N_4787);
nor U5405 (N_5405,N_4703,N_4585);
or U5406 (N_5406,N_4816,N_4570);
nor U5407 (N_5407,N_4841,N_4823);
and U5408 (N_5408,N_4795,N_4853);
and U5409 (N_5409,N_4794,N_4858);
and U5410 (N_5410,N_4695,N_4959);
or U5411 (N_5411,N_4948,N_4516);
or U5412 (N_5412,N_4599,N_4860);
nand U5413 (N_5413,N_4908,N_4732);
or U5414 (N_5414,N_4753,N_4639);
nand U5415 (N_5415,N_4571,N_4894);
nand U5416 (N_5416,N_4678,N_4968);
xor U5417 (N_5417,N_4568,N_4501);
nand U5418 (N_5418,N_4580,N_4619);
and U5419 (N_5419,N_4693,N_4707);
and U5420 (N_5420,N_4624,N_4803);
nand U5421 (N_5421,N_4660,N_4576);
nand U5422 (N_5422,N_4539,N_4717);
nand U5423 (N_5423,N_4892,N_4578);
xor U5424 (N_5424,N_4505,N_4543);
nor U5425 (N_5425,N_4619,N_4836);
nor U5426 (N_5426,N_4713,N_4907);
nor U5427 (N_5427,N_4754,N_4511);
nand U5428 (N_5428,N_4643,N_4504);
or U5429 (N_5429,N_4818,N_4983);
nor U5430 (N_5430,N_4919,N_4871);
and U5431 (N_5431,N_4510,N_4960);
nand U5432 (N_5432,N_4630,N_4825);
or U5433 (N_5433,N_4812,N_4968);
and U5434 (N_5434,N_4825,N_4927);
or U5435 (N_5435,N_4675,N_4624);
nor U5436 (N_5436,N_4621,N_4902);
nand U5437 (N_5437,N_4569,N_4585);
nor U5438 (N_5438,N_4570,N_4922);
xnor U5439 (N_5439,N_4787,N_4870);
xor U5440 (N_5440,N_4740,N_4976);
xnor U5441 (N_5441,N_4633,N_4908);
xor U5442 (N_5442,N_4789,N_4740);
or U5443 (N_5443,N_4506,N_4695);
nor U5444 (N_5444,N_4974,N_4689);
nor U5445 (N_5445,N_4692,N_4773);
or U5446 (N_5446,N_4847,N_4947);
or U5447 (N_5447,N_4783,N_4685);
nand U5448 (N_5448,N_4800,N_4686);
xnor U5449 (N_5449,N_4772,N_4761);
nor U5450 (N_5450,N_4875,N_4677);
nand U5451 (N_5451,N_4552,N_4800);
nor U5452 (N_5452,N_4934,N_4528);
and U5453 (N_5453,N_4870,N_4651);
xor U5454 (N_5454,N_4986,N_4668);
nor U5455 (N_5455,N_4579,N_4708);
or U5456 (N_5456,N_4783,N_4617);
nor U5457 (N_5457,N_4924,N_4573);
nor U5458 (N_5458,N_4886,N_4540);
or U5459 (N_5459,N_4555,N_4797);
or U5460 (N_5460,N_4884,N_4692);
xnor U5461 (N_5461,N_4982,N_4863);
nand U5462 (N_5462,N_4756,N_4997);
or U5463 (N_5463,N_4927,N_4763);
and U5464 (N_5464,N_4612,N_4567);
nor U5465 (N_5465,N_4770,N_4803);
or U5466 (N_5466,N_4917,N_4632);
nand U5467 (N_5467,N_4754,N_4778);
xnor U5468 (N_5468,N_4583,N_4687);
nor U5469 (N_5469,N_4502,N_4781);
nand U5470 (N_5470,N_4627,N_4579);
nand U5471 (N_5471,N_4697,N_4636);
nand U5472 (N_5472,N_4895,N_4784);
or U5473 (N_5473,N_4826,N_4822);
nand U5474 (N_5474,N_4964,N_4884);
or U5475 (N_5475,N_4914,N_4577);
nand U5476 (N_5476,N_4871,N_4578);
or U5477 (N_5477,N_4966,N_4509);
or U5478 (N_5478,N_4728,N_4970);
nand U5479 (N_5479,N_4657,N_4779);
xnor U5480 (N_5480,N_4719,N_4737);
nor U5481 (N_5481,N_4655,N_4934);
nor U5482 (N_5482,N_4813,N_4780);
nand U5483 (N_5483,N_4851,N_4520);
or U5484 (N_5484,N_4875,N_4580);
nand U5485 (N_5485,N_4519,N_4954);
nor U5486 (N_5486,N_4825,N_4938);
or U5487 (N_5487,N_4973,N_4912);
nand U5488 (N_5488,N_4644,N_4861);
or U5489 (N_5489,N_4904,N_4841);
nor U5490 (N_5490,N_4549,N_4709);
nand U5491 (N_5491,N_4789,N_4518);
and U5492 (N_5492,N_4876,N_4779);
nand U5493 (N_5493,N_4984,N_4696);
nor U5494 (N_5494,N_4768,N_4600);
nand U5495 (N_5495,N_4737,N_4793);
and U5496 (N_5496,N_4920,N_4855);
and U5497 (N_5497,N_4812,N_4742);
xor U5498 (N_5498,N_4522,N_4852);
and U5499 (N_5499,N_4552,N_4955);
and U5500 (N_5500,N_5245,N_5028);
xnor U5501 (N_5501,N_5089,N_5364);
or U5502 (N_5502,N_5435,N_5149);
and U5503 (N_5503,N_5204,N_5487);
and U5504 (N_5504,N_5485,N_5313);
and U5505 (N_5505,N_5175,N_5271);
nor U5506 (N_5506,N_5244,N_5053);
or U5507 (N_5507,N_5197,N_5168);
and U5508 (N_5508,N_5125,N_5082);
xnor U5509 (N_5509,N_5280,N_5355);
nand U5510 (N_5510,N_5206,N_5387);
and U5511 (N_5511,N_5259,N_5151);
or U5512 (N_5512,N_5333,N_5339);
and U5513 (N_5513,N_5170,N_5145);
or U5514 (N_5514,N_5220,N_5296);
nor U5515 (N_5515,N_5103,N_5134);
xor U5516 (N_5516,N_5369,N_5063);
nor U5517 (N_5517,N_5320,N_5338);
nand U5518 (N_5518,N_5256,N_5236);
nand U5519 (N_5519,N_5099,N_5349);
or U5520 (N_5520,N_5463,N_5423);
xnor U5521 (N_5521,N_5161,N_5179);
xnor U5522 (N_5522,N_5061,N_5076);
xnor U5523 (N_5523,N_5428,N_5273);
nor U5524 (N_5524,N_5407,N_5167);
nor U5525 (N_5525,N_5458,N_5129);
xor U5526 (N_5526,N_5288,N_5230);
nor U5527 (N_5527,N_5238,N_5264);
nor U5528 (N_5528,N_5469,N_5345);
nand U5529 (N_5529,N_5000,N_5427);
xor U5530 (N_5530,N_5111,N_5107);
nand U5531 (N_5531,N_5295,N_5316);
and U5532 (N_5532,N_5050,N_5101);
nand U5533 (N_5533,N_5362,N_5497);
and U5534 (N_5534,N_5222,N_5065);
nor U5535 (N_5535,N_5400,N_5274);
nand U5536 (N_5536,N_5038,N_5009);
xor U5537 (N_5537,N_5377,N_5212);
or U5538 (N_5538,N_5329,N_5224);
and U5539 (N_5539,N_5301,N_5095);
nor U5540 (N_5540,N_5247,N_5409);
xnor U5541 (N_5541,N_5386,N_5043);
nor U5542 (N_5542,N_5291,N_5140);
nor U5543 (N_5543,N_5182,N_5121);
or U5544 (N_5544,N_5173,N_5371);
xor U5545 (N_5545,N_5115,N_5327);
or U5546 (N_5546,N_5039,N_5491);
nor U5547 (N_5547,N_5334,N_5356);
and U5548 (N_5548,N_5252,N_5020);
and U5549 (N_5549,N_5010,N_5122);
xor U5550 (N_5550,N_5193,N_5464);
nor U5551 (N_5551,N_5144,N_5127);
nand U5552 (N_5552,N_5051,N_5433);
xnor U5553 (N_5553,N_5462,N_5282);
nor U5554 (N_5554,N_5283,N_5277);
or U5555 (N_5555,N_5359,N_5156);
and U5556 (N_5556,N_5395,N_5120);
nor U5557 (N_5557,N_5185,N_5284);
nand U5558 (N_5558,N_5106,N_5195);
and U5559 (N_5559,N_5452,N_5304);
nor U5560 (N_5560,N_5308,N_5315);
nor U5561 (N_5561,N_5293,N_5209);
or U5562 (N_5562,N_5399,N_5331);
nand U5563 (N_5563,N_5036,N_5449);
xnor U5564 (N_5564,N_5011,N_5314);
nor U5565 (N_5565,N_5326,N_5214);
nand U5566 (N_5566,N_5133,N_5303);
or U5567 (N_5567,N_5171,N_5080);
and U5568 (N_5568,N_5437,N_5154);
and U5569 (N_5569,N_5225,N_5201);
xnor U5570 (N_5570,N_5146,N_5380);
nand U5571 (N_5571,N_5354,N_5232);
nor U5572 (N_5572,N_5059,N_5418);
nor U5573 (N_5573,N_5461,N_5309);
and U5574 (N_5574,N_5219,N_5058);
xnor U5575 (N_5575,N_5057,N_5251);
or U5576 (N_5576,N_5162,N_5396);
xor U5577 (N_5577,N_5176,N_5227);
nand U5578 (N_5578,N_5202,N_5105);
nand U5579 (N_5579,N_5071,N_5360);
nand U5580 (N_5580,N_5310,N_5451);
and U5581 (N_5581,N_5319,N_5114);
xor U5582 (N_5582,N_5445,N_5254);
nor U5583 (N_5583,N_5088,N_5441);
xnor U5584 (N_5584,N_5450,N_5215);
xnor U5585 (N_5585,N_5322,N_5004);
nand U5586 (N_5586,N_5078,N_5055);
xnor U5587 (N_5587,N_5015,N_5024);
nor U5588 (N_5588,N_5198,N_5228);
xor U5589 (N_5589,N_5279,N_5023);
xor U5590 (N_5590,N_5174,N_5079);
and U5591 (N_5591,N_5372,N_5443);
and U5592 (N_5592,N_5012,N_5148);
and U5593 (N_5593,N_5081,N_5286);
nor U5594 (N_5594,N_5052,N_5203);
or U5595 (N_5595,N_5302,N_5434);
nand U5596 (N_5596,N_5477,N_5332);
xnor U5597 (N_5597,N_5471,N_5474);
xnor U5598 (N_5598,N_5479,N_5233);
nand U5599 (N_5599,N_5022,N_5073);
nor U5600 (N_5600,N_5229,N_5067);
xnor U5601 (N_5601,N_5401,N_5292);
or U5602 (N_5602,N_5272,N_5027);
nor U5603 (N_5603,N_5131,N_5218);
xor U5604 (N_5604,N_5221,N_5457);
nand U5605 (N_5605,N_5318,N_5268);
and U5606 (N_5606,N_5448,N_5064);
nor U5607 (N_5607,N_5180,N_5460);
or U5608 (N_5608,N_5306,N_5139);
nor U5609 (N_5609,N_5152,N_5062);
and U5610 (N_5610,N_5172,N_5499);
xor U5611 (N_5611,N_5379,N_5416);
or U5612 (N_5612,N_5002,N_5070);
nor U5613 (N_5613,N_5410,N_5041);
xnor U5614 (N_5614,N_5192,N_5265);
and U5615 (N_5615,N_5368,N_5253);
xor U5616 (N_5616,N_5047,N_5142);
xnor U5617 (N_5617,N_5137,N_5424);
xor U5618 (N_5618,N_5110,N_5455);
nor U5619 (N_5619,N_5217,N_5031);
nor U5620 (N_5620,N_5431,N_5388);
and U5621 (N_5621,N_5187,N_5132);
nand U5622 (N_5622,N_5014,N_5237);
or U5623 (N_5623,N_5408,N_5459);
xor U5624 (N_5624,N_5208,N_5030);
or U5625 (N_5625,N_5261,N_5413);
xnor U5626 (N_5626,N_5382,N_5033);
and U5627 (N_5627,N_5083,N_5008);
and U5628 (N_5628,N_5323,N_5381);
nand U5629 (N_5629,N_5444,N_5376);
xnor U5630 (N_5630,N_5472,N_5034);
and U5631 (N_5631,N_5365,N_5116);
or U5632 (N_5632,N_5235,N_5164);
xor U5633 (N_5633,N_5178,N_5420);
or U5634 (N_5634,N_5398,N_5210);
nor U5635 (N_5635,N_5275,N_5231);
nor U5636 (N_5636,N_5417,N_5211);
nand U5637 (N_5637,N_5013,N_5049);
and U5638 (N_5638,N_5084,N_5397);
and U5639 (N_5639,N_5317,N_5367);
or U5640 (N_5640,N_5478,N_5335);
or U5641 (N_5641,N_5188,N_5475);
nor U5642 (N_5642,N_5340,N_5046);
or U5643 (N_5643,N_5337,N_5312);
xor U5644 (N_5644,N_5263,N_5223);
xnor U5645 (N_5645,N_5032,N_5422);
nand U5646 (N_5646,N_5299,N_5189);
or U5647 (N_5647,N_5234,N_5135);
or U5648 (N_5648,N_5138,N_5343);
and U5649 (N_5649,N_5026,N_5124);
and U5650 (N_5650,N_5037,N_5199);
and U5651 (N_5651,N_5126,N_5109);
and U5652 (N_5652,N_5141,N_5447);
nor U5653 (N_5653,N_5200,N_5196);
nor U5654 (N_5654,N_5007,N_5147);
xor U5655 (N_5655,N_5108,N_5393);
and U5656 (N_5656,N_5442,N_5130);
xor U5657 (N_5657,N_5328,N_5021);
nand U5658 (N_5658,N_5440,N_5025);
or U5659 (N_5659,N_5456,N_5091);
and U5660 (N_5660,N_5425,N_5404);
xnor U5661 (N_5661,N_5045,N_5029);
nand U5662 (N_5662,N_5163,N_5287);
nand U5663 (N_5663,N_5255,N_5392);
nand U5664 (N_5664,N_5412,N_5085);
nor U5665 (N_5665,N_5098,N_5157);
or U5666 (N_5666,N_5366,N_5240);
xor U5667 (N_5667,N_5260,N_5205);
xnor U5668 (N_5668,N_5490,N_5439);
or U5669 (N_5669,N_5239,N_5006);
and U5670 (N_5670,N_5348,N_5426);
nand U5671 (N_5671,N_5361,N_5430);
and U5672 (N_5672,N_5289,N_5415);
nor U5673 (N_5673,N_5352,N_5118);
or U5674 (N_5674,N_5429,N_5311);
nor U5675 (N_5675,N_5074,N_5281);
or U5676 (N_5676,N_5068,N_5258);
xnor U5677 (N_5677,N_5470,N_5489);
nor U5678 (N_5678,N_5066,N_5384);
xnor U5679 (N_5679,N_5480,N_5092);
nand U5680 (N_5680,N_5241,N_5072);
nor U5681 (N_5681,N_5128,N_5019);
nand U5682 (N_5682,N_5394,N_5297);
or U5683 (N_5683,N_5484,N_5042);
nor U5684 (N_5684,N_5097,N_5207);
and U5685 (N_5685,N_5096,N_5181);
or U5686 (N_5686,N_5267,N_5136);
and U5687 (N_5687,N_5153,N_5242);
xor U5688 (N_5688,N_5270,N_5001);
or U5689 (N_5689,N_5075,N_5165);
nor U5690 (N_5690,N_5307,N_5373);
nor U5691 (N_5691,N_5243,N_5159);
nor U5692 (N_5692,N_5482,N_5093);
nand U5693 (N_5693,N_5465,N_5276);
xnor U5694 (N_5694,N_5446,N_5184);
and U5695 (N_5695,N_5325,N_5411);
xnor U5696 (N_5696,N_5246,N_5090);
xnor U5697 (N_5697,N_5488,N_5285);
nand U5698 (N_5698,N_5060,N_5496);
or U5699 (N_5699,N_5190,N_5191);
and U5700 (N_5700,N_5389,N_5390);
or U5701 (N_5701,N_5467,N_5363);
nor U5702 (N_5702,N_5077,N_5017);
xor U5703 (N_5703,N_5432,N_5269);
or U5704 (N_5704,N_5391,N_5414);
nand U5705 (N_5705,N_5492,N_5005);
and U5706 (N_5706,N_5100,N_5321);
nor U5707 (N_5707,N_5018,N_5344);
xor U5708 (N_5708,N_5374,N_5421);
nand U5709 (N_5709,N_5113,N_5300);
and U5710 (N_5710,N_5419,N_5370);
or U5711 (N_5711,N_5087,N_5155);
and U5712 (N_5712,N_5406,N_5158);
nor U5713 (N_5713,N_5336,N_5104);
nand U5714 (N_5714,N_5495,N_5056);
xor U5715 (N_5715,N_5358,N_5453);
nand U5716 (N_5716,N_5177,N_5290);
or U5717 (N_5717,N_5438,N_5375);
or U5718 (N_5718,N_5346,N_5102);
or U5719 (N_5719,N_5486,N_5040);
and U5720 (N_5720,N_5117,N_5123);
and U5721 (N_5721,N_5226,N_5351);
nand U5722 (N_5722,N_5330,N_5342);
xnor U5723 (N_5723,N_5494,N_5213);
nor U5724 (N_5724,N_5216,N_5402);
nand U5725 (N_5725,N_5383,N_5454);
nand U5726 (N_5726,N_5347,N_5166);
nor U5727 (N_5727,N_5498,N_5054);
xnor U5728 (N_5728,N_5186,N_5249);
nor U5729 (N_5729,N_5385,N_5112);
xnor U5730 (N_5730,N_5086,N_5278);
xnor U5731 (N_5731,N_5341,N_5481);
nand U5732 (N_5732,N_5003,N_5350);
nor U5733 (N_5733,N_5143,N_5324);
nand U5734 (N_5734,N_5476,N_5044);
xor U5735 (N_5735,N_5248,N_5493);
nand U5736 (N_5736,N_5194,N_5183);
or U5737 (N_5737,N_5169,N_5483);
nor U5738 (N_5738,N_5035,N_5353);
xor U5739 (N_5739,N_5466,N_5150);
or U5740 (N_5740,N_5250,N_5298);
nor U5741 (N_5741,N_5294,N_5468);
or U5742 (N_5742,N_5048,N_5357);
nand U5743 (N_5743,N_5160,N_5473);
or U5744 (N_5744,N_5119,N_5094);
nand U5745 (N_5745,N_5257,N_5405);
nor U5746 (N_5746,N_5403,N_5436);
nand U5747 (N_5747,N_5069,N_5266);
or U5748 (N_5748,N_5262,N_5016);
and U5749 (N_5749,N_5378,N_5305);
nor U5750 (N_5750,N_5497,N_5191);
xnor U5751 (N_5751,N_5019,N_5081);
xor U5752 (N_5752,N_5479,N_5106);
nor U5753 (N_5753,N_5376,N_5048);
xor U5754 (N_5754,N_5057,N_5458);
nor U5755 (N_5755,N_5491,N_5231);
or U5756 (N_5756,N_5001,N_5387);
or U5757 (N_5757,N_5049,N_5174);
and U5758 (N_5758,N_5404,N_5030);
nor U5759 (N_5759,N_5242,N_5135);
xor U5760 (N_5760,N_5279,N_5280);
or U5761 (N_5761,N_5004,N_5447);
xor U5762 (N_5762,N_5455,N_5085);
nand U5763 (N_5763,N_5049,N_5211);
nor U5764 (N_5764,N_5138,N_5276);
xnor U5765 (N_5765,N_5025,N_5225);
nor U5766 (N_5766,N_5160,N_5495);
nor U5767 (N_5767,N_5098,N_5393);
or U5768 (N_5768,N_5308,N_5347);
nand U5769 (N_5769,N_5103,N_5497);
xnor U5770 (N_5770,N_5183,N_5242);
and U5771 (N_5771,N_5159,N_5253);
nor U5772 (N_5772,N_5175,N_5307);
xnor U5773 (N_5773,N_5293,N_5392);
or U5774 (N_5774,N_5391,N_5174);
xnor U5775 (N_5775,N_5222,N_5401);
and U5776 (N_5776,N_5428,N_5483);
nand U5777 (N_5777,N_5454,N_5056);
and U5778 (N_5778,N_5357,N_5300);
and U5779 (N_5779,N_5123,N_5366);
xor U5780 (N_5780,N_5341,N_5216);
xor U5781 (N_5781,N_5018,N_5072);
nor U5782 (N_5782,N_5069,N_5184);
or U5783 (N_5783,N_5373,N_5231);
xor U5784 (N_5784,N_5172,N_5394);
nand U5785 (N_5785,N_5242,N_5446);
or U5786 (N_5786,N_5222,N_5338);
and U5787 (N_5787,N_5393,N_5118);
or U5788 (N_5788,N_5228,N_5281);
nand U5789 (N_5789,N_5458,N_5164);
nand U5790 (N_5790,N_5251,N_5110);
nand U5791 (N_5791,N_5367,N_5330);
or U5792 (N_5792,N_5012,N_5442);
and U5793 (N_5793,N_5136,N_5100);
nor U5794 (N_5794,N_5404,N_5188);
nand U5795 (N_5795,N_5060,N_5103);
or U5796 (N_5796,N_5031,N_5247);
and U5797 (N_5797,N_5496,N_5055);
xnor U5798 (N_5798,N_5188,N_5305);
or U5799 (N_5799,N_5296,N_5452);
xnor U5800 (N_5800,N_5179,N_5409);
nor U5801 (N_5801,N_5160,N_5226);
xor U5802 (N_5802,N_5153,N_5478);
and U5803 (N_5803,N_5488,N_5111);
or U5804 (N_5804,N_5224,N_5430);
and U5805 (N_5805,N_5061,N_5151);
nand U5806 (N_5806,N_5356,N_5280);
and U5807 (N_5807,N_5458,N_5281);
or U5808 (N_5808,N_5478,N_5357);
and U5809 (N_5809,N_5287,N_5269);
and U5810 (N_5810,N_5037,N_5041);
xnor U5811 (N_5811,N_5372,N_5171);
or U5812 (N_5812,N_5041,N_5319);
nor U5813 (N_5813,N_5103,N_5458);
and U5814 (N_5814,N_5008,N_5158);
and U5815 (N_5815,N_5116,N_5208);
or U5816 (N_5816,N_5168,N_5018);
xnor U5817 (N_5817,N_5481,N_5185);
and U5818 (N_5818,N_5322,N_5146);
or U5819 (N_5819,N_5106,N_5259);
or U5820 (N_5820,N_5133,N_5454);
nor U5821 (N_5821,N_5060,N_5297);
and U5822 (N_5822,N_5127,N_5370);
xnor U5823 (N_5823,N_5011,N_5384);
or U5824 (N_5824,N_5352,N_5392);
nand U5825 (N_5825,N_5137,N_5061);
nand U5826 (N_5826,N_5041,N_5024);
xor U5827 (N_5827,N_5090,N_5341);
or U5828 (N_5828,N_5167,N_5385);
and U5829 (N_5829,N_5373,N_5160);
nand U5830 (N_5830,N_5490,N_5034);
and U5831 (N_5831,N_5242,N_5079);
nand U5832 (N_5832,N_5060,N_5161);
xnor U5833 (N_5833,N_5273,N_5106);
xnor U5834 (N_5834,N_5152,N_5331);
or U5835 (N_5835,N_5192,N_5151);
xnor U5836 (N_5836,N_5212,N_5262);
xor U5837 (N_5837,N_5223,N_5429);
and U5838 (N_5838,N_5091,N_5373);
xor U5839 (N_5839,N_5062,N_5083);
and U5840 (N_5840,N_5425,N_5185);
nand U5841 (N_5841,N_5454,N_5186);
or U5842 (N_5842,N_5454,N_5199);
and U5843 (N_5843,N_5479,N_5071);
nand U5844 (N_5844,N_5289,N_5131);
and U5845 (N_5845,N_5361,N_5120);
and U5846 (N_5846,N_5143,N_5115);
nor U5847 (N_5847,N_5305,N_5252);
nand U5848 (N_5848,N_5487,N_5166);
xor U5849 (N_5849,N_5159,N_5204);
nor U5850 (N_5850,N_5060,N_5053);
xor U5851 (N_5851,N_5385,N_5072);
and U5852 (N_5852,N_5392,N_5126);
or U5853 (N_5853,N_5178,N_5436);
and U5854 (N_5854,N_5426,N_5247);
nand U5855 (N_5855,N_5379,N_5310);
xnor U5856 (N_5856,N_5027,N_5404);
nand U5857 (N_5857,N_5228,N_5118);
nand U5858 (N_5858,N_5258,N_5405);
or U5859 (N_5859,N_5036,N_5219);
and U5860 (N_5860,N_5078,N_5195);
and U5861 (N_5861,N_5253,N_5324);
nor U5862 (N_5862,N_5343,N_5237);
and U5863 (N_5863,N_5295,N_5348);
and U5864 (N_5864,N_5334,N_5296);
xor U5865 (N_5865,N_5362,N_5115);
and U5866 (N_5866,N_5318,N_5375);
nor U5867 (N_5867,N_5186,N_5075);
xnor U5868 (N_5868,N_5481,N_5258);
or U5869 (N_5869,N_5128,N_5162);
and U5870 (N_5870,N_5492,N_5381);
or U5871 (N_5871,N_5450,N_5462);
nor U5872 (N_5872,N_5042,N_5028);
and U5873 (N_5873,N_5134,N_5463);
or U5874 (N_5874,N_5485,N_5037);
or U5875 (N_5875,N_5263,N_5164);
xor U5876 (N_5876,N_5152,N_5067);
and U5877 (N_5877,N_5120,N_5350);
nand U5878 (N_5878,N_5075,N_5334);
nand U5879 (N_5879,N_5481,N_5079);
or U5880 (N_5880,N_5118,N_5082);
nor U5881 (N_5881,N_5287,N_5166);
and U5882 (N_5882,N_5317,N_5351);
or U5883 (N_5883,N_5180,N_5440);
nand U5884 (N_5884,N_5361,N_5455);
nand U5885 (N_5885,N_5128,N_5215);
nor U5886 (N_5886,N_5342,N_5409);
xor U5887 (N_5887,N_5293,N_5197);
xor U5888 (N_5888,N_5045,N_5206);
xnor U5889 (N_5889,N_5027,N_5182);
xnor U5890 (N_5890,N_5074,N_5037);
and U5891 (N_5891,N_5232,N_5355);
and U5892 (N_5892,N_5256,N_5379);
xor U5893 (N_5893,N_5355,N_5294);
or U5894 (N_5894,N_5373,N_5342);
or U5895 (N_5895,N_5165,N_5214);
xnor U5896 (N_5896,N_5105,N_5187);
or U5897 (N_5897,N_5192,N_5064);
and U5898 (N_5898,N_5323,N_5397);
nand U5899 (N_5899,N_5443,N_5094);
nand U5900 (N_5900,N_5193,N_5499);
and U5901 (N_5901,N_5190,N_5073);
xor U5902 (N_5902,N_5427,N_5086);
or U5903 (N_5903,N_5135,N_5033);
and U5904 (N_5904,N_5237,N_5309);
or U5905 (N_5905,N_5080,N_5158);
and U5906 (N_5906,N_5219,N_5222);
nor U5907 (N_5907,N_5494,N_5274);
and U5908 (N_5908,N_5280,N_5288);
nand U5909 (N_5909,N_5131,N_5209);
and U5910 (N_5910,N_5209,N_5428);
xor U5911 (N_5911,N_5140,N_5043);
nor U5912 (N_5912,N_5496,N_5098);
nor U5913 (N_5913,N_5095,N_5409);
nor U5914 (N_5914,N_5332,N_5487);
or U5915 (N_5915,N_5087,N_5062);
nand U5916 (N_5916,N_5124,N_5358);
and U5917 (N_5917,N_5382,N_5236);
and U5918 (N_5918,N_5138,N_5029);
or U5919 (N_5919,N_5135,N_5355);
xnor U5920 (N_5920,N_5461,N_5044);
nand U5921 (N_5921,N_5165,N_5451);
and U5922 (N_5922,N_5315,N_5115);
nor U5923 (N_5923,N_5469,N_5269);
xnor U5924 (N_5924,N_5350,N_5240);
nand U5925 (N_5925,N_5187,N_5052);
and U5926 (N_5926,N_5472,N_5140);
nand U5927 (N_5927,N_5368,N_5243);
nor U5928 (N_5928,N_5074,N_5370);
and U5929 (N_5929,N_5208,N_5490);
nand U5930 (N_5930,N_5497,N_5233);
or U5931 (N_5931,N_5024,N_5197);
and U5932 (N_5932,N_5071,N_5455);
nand U5933 (N_5933,N_5161,N_5278);
nand U5934 (N_5934,N_5268,N_5463);
nand U5935 (N_5935,N_5195,N_5286);
and U5936 (N_5936,N_5397,N_5149);
nor U5937 (N_5937,N_5270,N_5219);
or U5938 (N_5938,N_5286,N_5347);
or U5939 (N_5939,N_5248,N_5391);
xor U5940 (N_5940,N_5158,N_5247);
or U5941 (N_5941,N_5391,N_5102);
xor U5942 (N_5942,N_5391,N_5116);
or U5943 (N_5943,N_5329,N_5051);
xor U5944 (N_5944,N_5470,N_5228);
nand U5945 (N_5945,N_5247,N_5148);
or U5946 (N_5946,N_5271,N_5051);
xnor U5947 (N_5947,N_5428,N_5453);
or U5948 (N_5948,N_5403,N_5399);
nand U5949 (N_5949,N_5455,N_5201);
nand U5950 (N_5950,N_5076,N_5073);
or U5951 (N_5951,N_5324,N_5171);
or U5952 (N_5952,N_5142,N_5058);
or U5953 (N_5953,N_5275,N_5450);
nor U5954 (N_5954,N_5323,N_5057);
and U5955 (N_5955,N_5211,N_5014);
nor U5956 (N_5956,N_5019,N_5007);
xnor U5957 (N_5957,N_5109,N_5107);
or U5958 (N_5958,N_5129,N_5337);
or U5959 (N_5959,N_5440,N_5439);
xnor U5960 (N_5960,N_5198,N_5455);
nand U5961 (N_5961,N_5300,N_5443);
and U5962 (N_5962,N_5070,N_5163);
or U5963 (N_5963,N_5469,N_5338);
or U5964 (N_5964,N_5042,N_5072);
and U5965 (N_5965,N_5088,N_5296);
and U5966 (N_5966,N_5042,N_5372);
nor U5967 (N_5967,N_5082,N_5187);
nand U5968 (N_5968,N_5183,N_5425);
or U5969 (N_5969,N_5240,N_5306);
xnor U5970 (N_5970,N_5000,N_5372);
or U5971 (N_5971,N_5001,N_5363);
and U5972 (N_5972,N_5256,N_5323);
and U5973 (N_5973,N_5154,N_5233);
nand U5974 (N_5974,N_5221,N_5056);
or U5975 (N_5975,N_5233,N_5052);
nand U5976 (N_5976,N_5466,N_5186);
nand U5977 (N_5977,N_5341,N_5306);
nor U5978 (N_5978,N_5017,N_5171);
xor U5979 (N_5979,N_5026,N_5113);
or U5980 (N_5980,N_5202,N_5493);
and U5981 (N_5981,N_5452,N_5350);
xor U5982 (N_5982,N_5246,N_5329);
xnor U5983 (N_5983,N_5406,N_5093);
xnor U5984 (N_5984,N_5144,N_5486);
nand U5985 (N_5985,N_5450,N_5029);
and U5986 (N_5986,N_5493,N_5252);
and U5987 (N_5987,N_5282,N_5038);
nand U5988 (N_5988,N_5049,N_5105);
or U5989 (N_5989,N_5039,N_5036);
or U5990 (N_5990,N_5471,N_5467);
and U5991 (N_5991,N_5248,N_5290);
nor U5992 (N_5992,N_5288,N_5135);
xnor U5993 (N_5993,N_5377,N_5338);
nor U5994 (N_5994,N_5299,N_5057);
or U5995 (N_5995,N_5451,N_5198);
nand U5996 (N_5996,N_5265,N_5151);
nand U5997 (N_5997,N_5126,N_5383);
and U5998 (N_5998,N_5411,N_5453);
xor U5999 (N_5999,N_5212,N_5210);
nand U6000 (N_6000,N_5527,N_5778);
or U6001 (N_6001,N_5980,N_5981);
and U6002 (N_6002,N_5931,N_5547);
nand U6003 (N_6003,N_5625,N_5835);
nor U6004 (N_6004,N_5824,N_5875);
nand U6005 (N_6005,N_5869,N_5630);
nand U6006 (N_6006,N_5945,N_5811);
or U6007 (N_6007,N_5592,N_5564);
nand U6008 (N_6008,N_5615,N_5871);
nor U6009 (N_6009,N_5999,N_5705);
xnor U6010 (N_6010,N_5745,N_5728);
xnor U6011 (N_6011,N_5954,N_5982);
nand U6012 (N_6012,N_5925,N_5569);
nor U6013 (N_6013,N_5635,N_5560);
nor U6014 (N_6014,N_5856,N_5932);
and U6015 (N_6015,N_5755,N_5947);
nand U6016 (N_6016,N_5566,N_5520);
nor U6017 (N_6017,N_5846,N_5666);
and U6018 (N_6018,N_5712,N_5752);
nor U6019 (N_6019,N_5791,N_5938);
xor U6020 (N_6020,N_5785,N_5961);
nor U6021 (N_6021,N_5594,N_5538);
xnor U6022 (N_6022,N_5736,N_5927);
nand U6023 (N_6023,N_5814,N_5909);
nor U6024 (N_6024,N_5895,N_5861);
and U6025 (N_6025,N_5536,N_5739);
nand U6026 (N_6026,N_5949,N_5583);
and U6027 (N_6027,N_5512,N_5985);
nand U6028 (N_6028,N_5679,N_5612);
nor U6029 (N_6029,N_5575,N_5567);
xor U6030 (N_6030,N_5986,N_5524);
and U6031 (N_6031,N_5995,N_5907);
nor U6032 (N_6032,N_5530,N_5720);
and U6033 (N_6033,N_5775,N_5650);
or U6034 (N_6034,N_5879,N_5891);
nor U6035 (N_6035,N_5936,N_5704);
xor U6036 (N_6036,N_5678,N_5796);
or U6037 (N_6037,N_5550,N_5793);
nand U6038 (N_6038,N_5661,N_5855);
xnor U6039 (N_6039,N_5733,N_5649);
or U6040 (N_6040,N_5826,N_5781);
nor U6041 (N_6041,N_5528,N_5888);
xnor U6042 (N_6042,N_5957,N_5699);
or U6043 (N_6043,N_5970,N_5800);
xnor U6044 (N_6044,N_5944,N_5554);
or U6045 (N_6045,N_5509,N_5545);
and U6046 (N_6046,N_5929,N_5677);
and U6047 (N_6047,N_5843,N_5614);
nand U6048 (N_6048,N_5882,N_5659);
nor U6049 (N_6049,N_5546,N_5588);
nor U6050 (N_6050,N_5977,N_5764);
and U6051 (N_6051,N_5953,N_5783);
or U6052 (N_6052,N_5818,N_5549);
and U6053 (N_6053,N_5806,N_5820);
or U6054 (N_6054,N_5672,N_5717);
and U6055 (N_6055,N_5997,N_5765);
xor U6056 (N_6056,N_5795,N_5578);
nor U6057 (N_6057,N_5671,N_5600);
and U6058 (N_6058,N_5517,N_5548);
xor U6059 (N_6059,N_5631,N_5725);
xor U6060 (N_6060,N_5700,N_5807);
or U6061 (N_6061,N_5817,N_5878);
and U6062 (N_6062,N_5762,N_5884);
nor U6063 (N_6063,N_5643,N_5770);
and U6064 (N_6064,N_5786,N_5663);
or U6065 (N_6065,N_5722,N_5889);
xnor U6066 (N_6066,N_5732,N_5747);
and U6067 (N_6067,N_5809,N_5577);
and U6068 (N_6068,N_5868,N_5911);
nor U6069 (N_6069,N_5711,N_5771);
nor U6070 (N_6070,N_5919,N_5816);
xnor U6071 (N_6071,N_5853,N_5767);
xnor U6072 (N_6072,N_5810,N_5697);
nand U6073 (N_6073,N_5860,N_5563);
nand U6074 (N_6074,N_5555,N_5862);
xnor U6075 (N_6075,N_5518,N_5965);
or U6076 (N_6076,N_5832,N_5611);
nand U6077 (N_6077,N_5708,N_5952);
nor U6078 (N_6078,N_5808,N_5887);
or U6079 (N_6079,N_5539,N_5974);
xnor U6080 (N_6080,N_5993,N_5780);
or U6081 (N_6081,N_5601,N_5616);
and U6082 (N_6082,N_5730,N_5664);
and U6083 (N_6083,N_5680,N_5591);
or U6084 (N_6084,N_5833,N_5948);
xor U6085 (N_6085,N_5798,N_5758);
nor U6086 (N_6086,N_5768,N_5731);
nand U6087 (N_6087,N_5589,N_5813);
nor U6088 (N_6088,N_5918,N_5676);
or U6089 (N_6089,N_5667,N_5942);
and U6090 (N_6090,N_5573,N_5684);
xnor U6091 (N_6091,N_5541,N_5941);
or U6092 (N_6092,N_5501,N_5845);
nand U6093 (N_6093,N_5557,N_5966);
nor U6094 (N_6094,N_5877,N_5960);
xor U6095 (N_6095,N_5587,N_5513);
xnor U6096 (N_6096,N_5754,N_5531);
nand U6097 (N_6097,N_5865,N_5963);
nor U6098 (N_6098,N_5831,N_5702);
or U6099 (N_6099,N_5804,N_5913);
nor U6100 (N_6100,N_5946,N_5610);
and U6101 (N_6101,N_5928,N_5850);
or U6102 (N_6102,N_5782,N_5844);
or U6103 (N_6103,N_5572,N_5522);
xnor U6104 (N_6104,N_5607,N_5701);
nand U6105 (N_6105,N_5962,N_5883);
and U6106 (N_6106,N_5924,N_5683);
nand U6107 (N_6107,N_5709,N_5551);
nor U6108 (N_6108,N_5935,N_5593);
and U6109 (N_6109,N_5787,N_5734);
nor U6110 (N_6110,N_5742,N_5606);
or U6111 (N_6111,N_5759,N_5823);
nand U6112 (N_6112,N_5933,N_5828);
nor U6113 (N_6113,N_5690,N_5639);
or U6114 (N_6114,N_5714,N_5516);
or U6115 (N_6115,N_5689,N_5802);
and U6116 (N_6116,N_5633,N_5648);
xnor U6117 (N_6117,N_5596,N_5978);
or U6118 (N_6118,N_5642,N_5898);
and U6119 (N_6119,N_5797,N_5543);
and U6120 (N_6120,N_5901,N_5653);
nor U6121 (N_6121,N_5707,N_5735);
xor U6122 (N_6122,N_5652,N_5784);
nand U6123 (N_6123,N_5638,N_5568);
xor U6124 (N_6124,N_5685,N_5529);
nor U6125 (N_6125,N_5912,N_5988);
nor U6126 (N_6126,N_5620,N_5523);
or U6127 (N_6127,N_5983,N_5696);
or U6128 (N_6128,N_5915,N_5655);
or U6129 (N_6129,N_5830,N_5632);
nor U6130 (N_6130,N_5608,N_5744);
nor U6131 (N_6131,N_5951,N_5837);
nand U6132 (N_6132,N_5729,N_5687);
and U6133 (N_6133,N_5867,N_5971);
xnor U6134 (N_6134,N_5864,N_5674);
nand U6135 (N_6135,N_5723,N_5761);
or U6136 (N_6136,N_5975,N_5506);
nor U6137 (N_6137,N_5605,N_5822);
nor U6138 (N_6138,N_5662,N_5562);
xnor U6139 (N_6139,N_5640,N_5571);
and U6140 (N_6140,N_5646,N_5604);
nor U6141 (N_6141,N_5553,N_5902);
nand U6142 (N_6142,N_5794,N_5598);
and U6143 (N_6143,N_5644,N_5922);
and U6144 (N_6144,N_5852,N_5623);
and U6145 (N_6145,N_5899,N_5738);
nor U6146 (N_6146,N_5967,N_5503);
xor U6147 (N_6147,N_5827,N_5719);
nor U6148 (N_6148,N_5920,N_5519);
nor U6149 (N_6149,N_5724,N_5552);
xor U6150 (N_6150,N_5619,N_5848);
xor U6151 (N_6151,N_5658,N_5576);
xor U6152 (N_6152,N_5741,N_5636);
nor U6153 (N_6153,N_5900,N_5657);
nor U6154 (N_6154,N_5859,N_5579);
xnor U6155 (N_6155,N_5815,N_5968);
nand U6156 (N_6156,N_5597,N_5502);
nor U6157 (N_6157,N_5556,N_5613);
xnor U6158 (N_6158,N_5984,N_5976);
xnor U6159 (N_6159,N_5609,N_5698);
nand U6160 (N_6160,N_5656,N_5626);
xnor U6161 (N_6161,N_5505,N_5989);
and U6162 (N_6162,N_5651,N_5673);
nand U6163 (N_6163,N_5670,N_5737);
xnor U6164 (N_6164,N_5621,N_5574);
xnor U6165 (N_6165,N_5972,N_5950);
nand U6166 (N_6166,N_5703,N_5637);
xor U6167 (N_6167,N_5774,N_5792);
nor U6168 (N_6168,N_5873,N_5964);
or U6169 (N_6169,N_5559,N_5668);
xor U6170 (N_6170,N_5540,N_5990);
nor U6171 (N_6171,N_5532,N_5885);
or U6172 (N_6172,N_5743,N_5544);
and U6173 (N_6173,N_5956,N_5841);
or U6174 (N_6174,N_5803,N_5746);
nand U6175 (N_6175,N_5876,N_5749);
nand U6176 (N_6176,N_5504,N_5716);
or U6177 (N_6177,N_5688,N_5838);
xnor U6178 (N_6178,N_5669,N_5525);
xnor U6179 (N_6179,N_5894,N_5776);
and U6180 (N_6180,N_5854,N_5763);
nand U6181 (N_6181,N_5533,N_5991);
and U6182 (N_6182,N_5872,N_5681);
or U6183 (N_6183,N_5940,N_5586);
and U6184 (N_6184,N_5617,N_5558);
nor U6185 (N_6185,N_5706,N_5721);
xor U6186 (N_6186,N_5590,N_5773);
xor U6187 (N_6187,N_5694,N_5727);
nor U6188 (N_6188,N_5629,N_5713);
and U6189 (N_6189,N_5602,N_5939);
and U6190 (N_6190,N_5585,N_5599);
nor U6191 (N_6191,N_5760,N_5840);
xor U6192 (N_6192,N_5923,N_5926);
or U6193 (N_6193,N_5582,N_5624);
and U6194 (N_6194,N_5847,N_5757);
nand U6195 (N_6195,N_5842,N_5996);
nand U6196 (N_6196,N_5665,N_5955);
nor U6197 (N_6197,N_5890,N_5777);
or U6198 (N_6198,N_5686,N_5937);
or U6199 (N_6199,N_5779,N_5969);
nor U6200 (N_6200,N_5819,N_5851);
nor U6201 (N_6201,N_5914,N_5691);
nand U6202 (N_6202,N_5805,N_5904);
and U6203 (N_6203,N_5751,N_5500);
nand U6204 (N_6204,N_5570,N_5866);
xor U6205 (N_6205,N_5726,N_5511);
or U6206 (N_6206,N_5881,N_5839);
or U6207 (N_6207,N_5829,N_5998);
nor U6208 (N_6208,N_5897,N_5718);
nor U6209 (N_6209,N_5910,N_5789);
and U6210 (N_6210,N_5618,N_5740);
or U6211 (N_6211,N_5535,N_5580);
and U6212 (N_6212,N_5695,N_5682);
or U6213 (N_6213,N_5748,N_5870);
xnor U6214 (N_6214,N_5788,N_5858);
or U6215 (N_6215,N_5906,N_5581);
or U6216 (N_6216,N_5959,N_5790);
or U6217 (N_6217,N_5510,N_5654);
nor U6218 (N_6218,N_5934,N_5692);
xor U6219 (N_6219,N_5534,N_5515);
and U6220 (N_6220,N_5834,N_5908);
and U6221 (N_6221,N_5756,N_5508);
nor U6222 (N_6222,N_5992,N_5892);
xnor U6223 (N_6223,N_5584,N_5622);
xnor U6224 (N_6224,N_5772,N_5863);
xnor U6225 (N_6225,N_5849,N_5514);
nand U6226 (N_6226,N_5526,N_5921);
or U6227 (N_6227,N_5521,N_5903);
nand U6228 (N_6228,N_5595,N_5542);
or U6229 (N_6229,N_5821,N_5766);
nor U6230 (N_6230,N_5627,N_5943);
nor U6231 (N_6231,N_5973,N_5930);
or U6232 (N_6232,N_5880,N_5916);
or U6233 (N_6233,N_5836,N_5507);
or U6234 (N_6234,N_5812,N_5628);
nor U6235 (N_6235,N_5994,N_5893);
or U6236 (N_6236,N_5769,N_5801);
xnor U6237 (N_6237,N_5874,N_5537);
or U6238 (N_6238,N_5886,N_5799);
nand U6239 (N_6239,N_5645,N_5979);
xor U6240 (N_6240,N_5647,N_5634);
or U6241 (N_6241,N_5917,N_5750);
xor U6242 (N_6242,N_5675,N_5715);
nand U6243 (N_6243,N_5603,N_5905);
and U6244 (N_6244,N_5565,N_5825);
xnor U6245 (N_6245,N_5641,N_5710);
xor U6246 (N_6246,N_5753,N_5987);
nand U6247 (N_6247,N_5693,N_5857);
or U6248 (N_6248,N_5958,N_5561);
xnor U6249 (N_6249,N_5660,N_5896);
and U6250 (N_6250,N_5772,N_5507);
nor U6251 (N_6251,N_5609,N_5950);
or U6252 (N_6252,N_5545,N_5528);
or U6253 (N_6253,N_5712,N_5575);
and U6254 (N_6254,N_5524,N_5846);
nand U6255 (N_6255,N_5700,N_5610);
or U6256 (N_6256,N_5509,N_5868);
and U6257 (N_6257,N_5640,N_5967);
nand U6258 (N_6258,N_5530,N_5513);
nor U6259 (N_6259,N_5524,N_5983);
nor U6260 (N_6260,N_5966,N_5579);
or U6261 (N_6261,N_5788,N_5658);
xor U6262 (N_6262,N_5812,N_5541);
nand U6263 (N_6263,N_5892,N_5953);
nand U6264 (N_6264,N_5779,N_5701);
nand U6265 (N_6265,N_5708,N_5715);
xor U6266 (N_6266,N_5734,N_5852);
or U6267 (N_6267,N_5984,N_5920);
or U6268 (N_6268,N_5823,N_5940);
and U6269 (N_6269,N_5506,N_5565);
nor U6270 (N_6270,N_5539,N_5936);
or U6271 (N_6271,N_5877,N_5700);
and U6272 (N_6272,N_5911,N_5773);
or U6273 (N_6273,N_5596,N_5970);
or U6274 (N_6274,N_5811,N_5683);
nor U6275 (N_6275,N_5736,N_5977);
xnor U6276 (N_6276,N_5731,N_5947);
nor U6277 (N_6277,N_5637,N_5761);
nor U6278 (N_6278,N_5619,N_5539);
or U6279 (N_6279,N_5737,N_5540);
or U6280 (N_6280,N_5568,N_5561);
nand U6281 (N_6281,N_5692,N_5973);
nand U6282 (N_6282,N_5926,N_5670);
nor U6283 (N_6283,N_5970,N_5948);
nand U6284 (N_6284,N_5930,N_5612);
xnor U6285 (N_6285,N_5787,N_5707);
and U6286 (N_6286,N_5932,N_5501);
nand U6287 (N_6287,N_5537,N_5710);
or U6288 (N_6288,N_5672,N_5806);
and U6289 (N_6289,N_5900,N_5956);
and U6290 (N_6290,N_5944,N_5715);
nor U6291 (N_6291,N_5652,N_5721);
or U6292 (N_6292,N_5887,N_5856);
and U6293 (N_6293,N_5960,N_5832);
or U6294 (N_6294,N_5778,N_5708);
nor U6295 (N_6295,N_5847,N_5658);
nand U6296 (N_6296,N_5689,N_5719);
and U6297 (N_6297,N_5797,N_5652);
nand U6298 (N_6298,N_5674,N_5943);
nor U6299 (N_6299,N_5888,N_5692);
xor U6300 (N_6300,N_5593,N_5517);
nor U6301 (N_6301,N_5575,N_5658);
nor U6302 (N_6302,N_5712,N_5956);
nor U6303 (N_6303,N_5698,N_5622);
nand U6304 (N_6304,N_5944,N_5522);
and U6305 (N_6305,N_5551,N_5613);
nor U6306 (N_6306,N_5747,N_5873);
and U6307 (N_6307,N_5733,N_5630);
nor U6308 (N_6308,N_5814,N_5591);
xnor U6309 (N_6309,N_5848,N_5796);
xnor U6310 (N_6310,N_5731,N_5717);
and U6311 (N_6311,N_5826,N_5520);
nor U6312 (N_6312,N_5889,N_5874);
and U6313 (N_6313,N_5579,N_5699);
and U6314 (N_6314,N_5820,N_5832);
and U6315 (N_6315,N_5750,N_5970);
nor U6316 (N_6316,N_5821,N_5990);
xnor U6317 (N_6317,N_5527,N_5909);
and U6318 (N_6318,N_5816,N_5999);
nand U6319 (N_6319,N_5548,N_5521);
or U6320 (N_6320,N_5716,N_5673);
and U6321 (N_6321,N_5954,N_5911);
or U6322 (N_6322,N_5637,N_5893);
and U6323 (N_6323,N_5624,N_5998);
nor U6324 (N_6324,N_5562,N_5977);
or U6325 (N_6325,N_5706,N_5994);
nor U6326 (N_6326,N_5585,N_5733);
or U6327 (N_6327,N_5611,N_5920);
and U6328 (N_6328,N_5613,N_5672);
nor U6329 (N_6329,N_5628,N_5847);
or U6330 (N_6330,N_5634,N_5727);
nor U6331 (N_6331,N_5962,N_5723);
xnor U6332 (N_6332,N_5746,N_5676);
and U6333 (N_6333,N_5681,N_5532);
and U6334 (N_6334,N_5849,N_5598);
and U6335 (N_6335,N_5856,N_5625);
nand U6336 (N_6336,N_5532,N_5508);
or U6337 (N_6337,N_5954,N_5693);
and U6338 (N_6338,N_5611,N_5873);
nand U6339 (N_6339,N_5507,N_5626);
nand U6340 (N_6340,N_5640,N_5573);
nor U6341 (N_6341,N_5687,N_5777);
nand U6342 (N_6342,N_5791,N_5677);
or U6343 (N_6343,N_5604,N_5855);
nand U6344 (N_6344,N_5612,N_5859);
or U6345 (N_6345,N_5797,N_5506);
xnor U6346 (N_6346,N_5891,N_5895);
nand U6347 (N_6347,N_5659,N_5517);
nand U6348 (N_6348,N_5942,N_5935);
or U6349 (N_6349,N_5506,N_5549);
xor U6350 (N_6350,N_5718,N_5810);
xnor U6351 (N_6351,N_5951,N_5741);
xnor U6352 (N_6352,N_5532,N_5706);
or U6353 (N_6353,N_5941,N_5991);
and U6354 (N_6354,N_5768,N_5848);
and U6355 (N_6355,N_5764,N_5708);
xor U6356 (N_6356,N_5505,N_5582);
and U6357 (N_6357,N_5549,N_5707);
nor U6358 (N_6358,N_5807,N_5548);
and U6359 (N_6359,N_5797,N_5534);
nor U6360 (N_6360,N_5512,N_5694);
and U6361 (N_6361,N_5812,N_5890);
nor U6362 (N_6362,N_5686,N_5778);
xor U6363 (N_6363,N_5864,N_5946);
nand U6364 (N_6364,N_5536,N_5869);
nand U6365 (N_6365,N_5999,N_5536);
and U6366 (N_6366,N_5740,N_5736);
xor U6367 (N_6367,N_5657,N_5570);
or U6368 (N_6368,N_5681,N_5885);
nor U6369 (N_6369,N_5831,N_5628);
nor U6370 (N_6370,N_5503,N_5610);
and U6371 (N_6371,N_5576,N_5571);
nand U6372 (N_6372,N_5592,N_5867);
nor U6373 (N_6373,N_5585,N_5784);
nand U6374 (N_6374,N_5887,N_5749);
xnor U6375 (N_6375,N_5707,N_5531);
xnor U6376 (N_6376,N_5899,N_5613);
nand U6377 (N_6377,N_5706,N_5899);
or U6378 (N_6378,N_5893,N_5657);
or U6379 (N_6379,N_5701,N_5753);
nand U6380 (N_6380,N_5987,N_5801);
xor U6381 (N_6381,N_5972,N_5758);
nor U6382 (N_6382,N_5807,N_5989);
nor U6383 (N_6383,N_5591,N_5586);
and U6384 (N_6384,N_5787,N_5912);
or U6385 (N_6385,N_5579,N_5536);
or U6386 (N_6386,N_5725,N_5641);
or U6387 (N_6387,N_5987,N_5797);
nor U6388 (N_6388,N_5594,N_5531);
xor U6389 (N_6389,N_5986,N_5798);
xnor U6390 (N_6390,N_5683,N_5737);
xor U6391 (N_6391,N_5962,N_5909);
and U6392 (N_6392,N_5544,N_5895);
or U6393 (N_6393,N_5914,N_5827);
nand U6394 (N_6394,N_5534,N_5766);
xor U6395 (N_6395,N_5962,N_5768);
xor U6396 (N_6396,N_5838,N_5769);
or U6397 (N_6397,N_5982,N_5994);
nor U6398 (N_6398,N_5878,N_5955);
nand U6399 (N_6399,N_5941,N_5960);
and U6400 (N_6400,N_5672,N_5635);
nor U6401 (N_6401,N_5778,N_5718);
nor U6402 (N_6402,N_5975,N_5787);
nand U6403 (N_6403,N_5900,N_5666);
nand U6404 (N_6404,N_5847,N_5948);
nor U6405 (N_6405,N_5949,N_5778);
nor U6406 (N_6406,N_5864,N_5758);
nand U6407 (N_6407,N_5986,N_5607);
nor U6408 (N_6408,N_5668,N_5821);
and U6409 (N_6409,N_5856,N_5667);
nand U6410 (N_6410,N_5881,N_5788);
xnor U6411 (N_6411,N_5670,N_5609);
nor U6412 (N_6412,N_5610,N_5591);
xnor U6413 (N_6413,N_5558,N_5711);
nor U6414 (N_6414,N_5643,N_5653);
or U6415 (N_6415,N_5933,N_5552);
and U6416 (N_6416,N_5690,N_5776);
and U6417 (N_6417,N_5919,N_5893);
xor U6418 (N_6418,N_5922,N_5824);
xnor U6419 (N_6419,N_5932,N_5773);
xnor U6420 (N_6420,N_5520,N_5845);
or U6421 (N_6421,N_5816,N_5861);
and U6422 (N_6422,N_5858,N_5903);
xor U6423 (N_6423,N_5733,N_5981);
xnor U6424 (N_6424,N_5839,N_5566);
and U6425 (N_6425,N_5844,N_5563);
nor U6426 (N_6426,N_5589,N_5683);
nand U6427 (N_6427,N_5881,N_5571);
xnor U6428 (N_6428,N_5663,N_5779);
xnor U6429 (N_6429,N_5857,N_5609);
and U6430 (N_6430,N_5816,N_5921);
nand U6431 (N_6431,N_5808,N_5784);
nor U6432 (N_6432,N_5775,N_5938);
or U6433 (N_6433,N_5770,N_5900);
and U6434 (N_6434,N_5609,N_5517);
nor U6435 (N_6435,N_5791,N_5962);
and U6436 (N_6436,N_5897,N_5938);
nand U6437 (N_6437,N_5839,N_5618);
or U6438 (N_6438,N_5883,N_5945);
or U6439 (N_6439,N_5550,N_5715);
nor U6440 (N_6440,N_5537,N_5574);
and U6441 (N_6441,N_5683,N_5988);
xnor U6442 (N_6442,N_5860,N_5692);
xor U6443 (N_6443,N_5709,N_5708);
nand U6444 (N_6444,N_5781,N_5773);
xnor U6445 (N_6445,N_5823,N_5957);
nor U6446 (N_6446,N_5946,N_5512);
and U6447 (N_6447,N_5585,N_5573);
nand U6448 (N_6448,N_5784,N_5915);
xor U6449 (N_6449,N_5706,N_5939);
and U6450 (N_6450,N_5726,N_5608);
nor U6451 (N_6451,N_5910,N_5528);
nand U6452 (N_6452,N_5600,N_5571);
and U6453 (N_6453,N_5843,N_5998);
xor U6454 (N_6454,N_5880,N_5598);
or U6455 (N_6455,N_5720,N_5941);
xnor U6456 (N_6456,N_5672,N_5831);
nor U6457 (N_6457,N_5550,N_5943);
nand U6458 (N_6458,N_5583,N_5995);
nand U6459 (N_6459,N_5633,N_5682);
and U6460 (N_6460,N_5559,N_5827);
xnor U6461 (N_6461,N_5664,N_5913);
nand U6462 (N_6462,N_5943,N_5646);
xnor U6463 (N_6463,N_5936,N_5564);
or U6464 (N_6464,N_5878,N_5526);
nand U6465 (N_6465,N_5964,N_5528);
and U6466 (N_6466,N_5845,N_5573);
or U6467 (N_6467,N_5911,N_5563);
nand U6468 (N_6468,N_5733,N_5533);
nor U6469 (N_6469,N_5683,N_5621);
nand U6470 (N_6470,N_5678,N_5520);
nor U6471 (N_6471,N_5911,N_5741);
xor U6472 (N_6472,N_5535,N_5508);
and U6473 (N_6473,N_5871,N_5702);
nor U6474 (N_6474,N_5668,N_5845);
nor U6475 (N_6475,N_5683,N_5828);
xnor U6476 (N_6476,N_5735,N_5837);
xor U6477 (N_6477,N_5725,N_5625);
nand U6478 (N_6478,N_5962,N_5732);
and U6479 (N_6479,N_5930,N_5847);
and U6480 (N_6480,N_5983,N_5999);
xor U6481 (N_6481,N_5509,N_5843);
nand U6482 (N_6482,N_5813,N_5841);
nor U6483 (N_6483,N_5781,N_5884);
nand U6484 (N_6484,N_5537,N_5797);
or U6485 (N_6485,N_5947,N_5850);
xor U6486 (N_6486,N_5851,N_5969);
and U6487 (N_6487,N_5724,N_5726);
xor U6488 (N_6488,N_5739,N_5714);
nor U6489 (N_6489,N_5918,N_5754);
xor U6490 (N_6490,N_5823,N_5616);
nor U6491 (N_6491,N_5849,N_5946);
or U6492 (N_6492,N_5787,N_5844);
xnor U6493 (N_6493,N_5684,N_5972);
or U6494 (N_6494,N_5814,N_5927);
xor U6495 (N_6495,N_5789,N_5978);
nand U6496 (N_6496,N_5690,N_5513);
nand U6497 (N_6497,N_5500,N_5903);
xnor U6498 (N_6498,N_5597,N_5580);
nand U6499 (N_6499,N_5759,N_5793);
nand U6500 (N_6500,N_6221,N_6231);
and U6501 (N_6501,N_6156,N_6095);
xor U6502 (N_6502,N_6263,N_6124);
and U6503 (N_6503,N_6477,N_6373);
xor U6504 (N_6504,N_6365,N_6229);
and U6505 (N_6505,N_6108,N_6311);
nand U6506 (N_6506,N_6326,N_6459);
or U6507 (N_6507,N_6271,N_6080);
or U6508 (N_6508,N_6481,N_6044);
nor U6509 (N_6509,N_6194,N_6069);
nand U6510 (N_6510,N_6497,N_6171);
nor U6511 (N_6511,N_6362,N_6356);
nand U6512 (N_6512,N_6342,N_6375);
or U6513 (N_6513,N_6010,N_6451);
or U6514 (N_6514,N_6205,N_6254);
xor U6515 (N_6515,N_6429,N_6439);
nand U6516 (N_6516,N_6323,N_6130);
or U6517 (N_6517,N_6336,N_6167);
nor U6518 (N_6518,N_6434,N_6187);
xnor U6519 (N_6519,N_6438,N_6480);
nand U6520 (N_6520,N_6456,N_6093);
nand U6521 (N_6521,N_6275,N_6207);
nor U6522 (N_6522,N_6354,N_6183);
nand U6523 (N_6523,N_6033,N_6049);
or U6524 (N_6524,N_6152,N_6418);
and U6525 (N_6525,N_6397,N_6128);
and U6526 (N_6526,N_6064,N_6237);
nor U6527 (N_6527,N_6057,N_6235);
xnor U6528 (N_6528,N_6161,N_6097);
nor U6529 (N_6529,N_6118,N_6313);
nor U6530 (N_6530,N_6426,N_6310);
nor U6531 (N_6531,N_6471,N_6173);
or U6532 (N_6532,N_6475,N_6169);
nor U6533 (N_6533,N_6296,N_6062);
or U6534 (N_6534,N_6148,N_6184);
nand U6535 (N_6535,N_6488,N_6320);
xor U6536 (N_6536,N_6299,N_6105);
or U6537 (N_6537,N_6153,N_6021);
and U6538 (N_6538,N_6012,N_6157);
or U6539 (N_6539,N_6404,N_6084);
or U6540 (N_6540,N_6028,N_6432);
nor U6541 (N_6541,N_6328,N_6457);
or U6542 (N_6542,N_6103,N_6106);
nor U6543 (N_6543,N_6135,N_6361);
nor U6544 (N_6544,N_6151,N_6092);
nand U6545 (N_6545,N_6000,N_6266);
nand U6546 (N_6546,N_6415,N_6176);
and U6547 (N_6547,N_6467,N_6253);
or U6548 (N_6548,N_6146,N_6154);
and U6549 (N_6549,N_6117,N_6413);
nor U6550 (N_6550,N_6129,N_6408);
or U6551 (N_6551,N_6283,N_6306);
xnor U6552 (N_6552,N_6255,N_6127);
nand U6553 (N_6553,N_6465,N_6054);
nor U6554 (N_6554,N_6216,N_6494);
or U6555 (N_6555,N_6496,N_6066);
and U6556 (N_6556,N_6293,N_6339);
nor U6557 (N_6557,N_6249,N_6450);
nor U6558 (N_6558,N_6282,N_6453);
nor U6559 (N_6559,N_6192,N_6285);
xor U6560 (N_6560,N_6363,N_6380);
xnor U6561 (N_6561,N_6047,N_6198);
nand U6562 (N_6562,N_6458,N_6368);
nor U6563 (N_6563,N_6083,N_6428);
nor U6564 (N_6564,N_6498,N_6197);
or U6565 (N_6565,N_6182,N_6330);
or U6566 (N_6566,N_6341,N_6357);
and U6567 (N_6567,N_6437,N_6369);
xnor U6568 (N_6568,N_6139,N_6226);
and U6569 (N_6569,N_6111,N_6075);
or U6570 (N_6570,N_6256,N_6405);
or U6571 (N_6571,N_6360,N_6185);
xor U6572 (N_6572,N_6468,N_6203);
nand U6573 (N_6573,N_6499,N_6273);
nor U6574 (N_6574,N_6242,N_6061);
nor U6575 (N_6575,N_6208,N_6279);
nor U6576 (N_6576,N_6337,N_6303);
nor U6577 (N_6577,N_6232,N_6179);
xnor U6578 (N_6578,N_6164,N_6199);
and U6579 (N_6579,N_6052,N_6091);
and U6580 (N_6580,N_6298,N_6019);
nand U6581 (N_6581,N_6304,N_6178);
or U6582 (N_6582,N_6442,N_6238);
nand U6583 (N_6583,N_6170,N_6406);
and U6584 (N_6584,N_6445,N_6359);
xnor U6585 (N_6585,N_6291,N_6041);
nor U6586 (N_6586,N_6074,N_6324);
or U6587 (N_6587,N_6250,N_6202);
nand U6588 (N_6588,N_6007,N_6295);
and U6589 (N_6589,N_6053,N_6201);
nand U6590 (N_6590,N_6227,N_6452);
nand U6591 (N_6591,N_6140,N_6409);
nor U6592 (N_6592,N_6267,N_6213);
or U6593 (N_6593,N_6204,N_6114);
and U6594 (N_6594,N_6329,N_6476);
or U6595 (N_6595,N_6484,N_6284);
and U6596 (N_6596,N_6034,N_6463);
xnor U6597 (N_6597,N_6101,N_6414);
and U6598 (N_6598,N_6327,N_6150);
nand U6599 (N_6599,N_6030,N_6393);
or U6600 (N_6600,N_6340,N_6050);
nor U6601 (N_6601,N_6042,N_6149);
and U6602 (N_6602,N_6272,N_6089);
xor U6603 (N_6603,N_6345,N_6319);
and U6604 (N_6604,N_6421,N_6419);
or U6605 (N_6605,N_6158,N_6215);
nand U6606 (N_6606,N_6455,N_6402);
and U6607 (N_6607,N_6046,N_6018);
xnor U6608 (N_6608,N_6196,N_6400);
nor U6609 (N_6609,N_6024,N_6314);
and U6610 (N_6610,N_6412,N_6248);
xor U6611 (N_6611,N_6073,N_6276);
or U6612 (N_6612,N_6035,N_6020);
nand U6613 (N_6613,N_6219,N_6113);
nand U6614 (N_6614,N_6444,N_6430);
or U6615 (N_6615,N_6258,N_6241);
nor U6616 (N_6616,N_6087,N_6121);
nand U6617 (N_6617,N_6200,N_6165);
nor U6618 (N_6618,N_6487,N_6260);
xor U6619 (N_6619,N_6411,N_6358);
or U6620 (N_6620,N_6206,N_6252);
nand U6621 (N_6621,N_6190,N_6220);
xor U6622 (N_6622,N_6399,N_6063);
or U6623 (N_6623,N_6144,N_6321);
or U6624 (N_6624,N_6268,N_6441);
nand U6625 (N_6625,N_6486,N_6214);
and U6626 (N_6626,N_6004,N_6056);
nor U6627 (N_6627,N_6243,N_6120);
nor U6628 (N_6628,N_6302,N_6349);
and U6629 (N_6629,N_6222,N_6239);
xor U6630 (N_6630,N_6338,N_6294);
nand U6631 (N_6631,N_6236,N_6068);
nor U6632 (N_6632,N_6223,N_6076);
nand U6633 (N_6633,N_6281,N_6446);
or U6634 (N_6634,N_6464,N_6043);
or U6635 (N_6635,N_6423,N_6265);
or U6636 (N_6636,N_6315,N_6489);
nand U6637 (N_6637,N_6479,N_6134);
nor U6638 (N_6638,N_6388,N_6462);
nand U6639 (N_6639,N_6211,N_6482);
and U6640 (N_6640,N_6013,N_6228);
nand U6641 (N_6641,N_6225,N_6096);
nor U6642 (N_6642,N_6261,N_6278);
nor U6643 (N_6643,N_6383,N_6060);
and U6644 (N_6644,N_6188,N_6259);
nor U6645 (N_6645,N_6424,N_6318);
xnor U6646 (N_6646,N_6079,N_6138);
or U6647 (N_6647,N_6448,N_6290);
or U6648 (N_6648,N_6191,N_6193);
nor U6649 (N_6649,N_6372,N_6472);
or U6650 (N_6650,N_6297,N_6377);
nor U6651 (N_6651,N_6071,N_6022);
xor U6652 (N_6652,N_6131,N_6332);
or U6653 (N_6653,N_6367,N_6309);
nor U6654 (N_6654,N_6233,N_6287);
nand U6655 (N_6655,N_6123,N_6417);
nor U6656 (N_6656,N_6343,N_6174);
xor U6657 (N_6657,N_6015,N_6029);
and U6658 (N_6658,N_6023,N_6466);
and U6659 (N_6659,N_6186,N_6147);
xor U6660 (N_6660,N_6391,N_6474);
or U6661 (N_6661,N_6422,N_6017);
xor U6662 (N_6662,N_6112,N_6346);
and U6663 (N_6663,N_6104,N_6433);
nor U6664 (N_6664,N_6011,N_6435);
or U6665 (N_6665,N_6366,N_6269);
or U6666 (N_6666,N_6085,N_6002);
nand U6667 (N_6667,N_6300,N_6172);
nand U6668 (N_6668,N_6110,N_6316);
nand U6669 (N_6669,N_6387,N_6055);
nor U6670 (N_6670,N_6051,N_6348);
nor U6671 (N_6671,N_6335,N_6122);
and U6672 (N_6672,N_6485,N_6065);
xor U6673 (N_6673,N_6257,N_6478);
nand U6674 (N_6674,N_6132,N_6246);
nand U6675 (N_6675,N_6425,N_6155);
or U6676 (N_6676,N_6159,N_6067);
xnor U6677 (N_6677,N_6385,N_6447);
and U6678 (N_6678,N_6492,N_6045);
nand U6679 (N_6679,N_6088,N_6078);
nand U6680 (N_6680,N_6027,N_6100);
or U6681 (N_6681,N_6005,N_6014);
nor U6682 (N_6682,N_6077,N_6039);
xor U6683 (N_6683,N_6251,N_6119);
and U6684 (N_6684,N_6440,N_6195);
nor U6685 (N_6685,N_6469,N_6059);
or U6686 (N_6686,N_6026,N_6379);
and U6687 (N_6687,N_6003,N_6277);
xor U6688 (N_6688,N_6137,N_6224);
nor U6689 (N_6689,N_6142,N_6431);
or U6690 (N_6690,N_6016,N_6334);
and U6691 (N_6691,N_6352,N_6410);
or U6692 (N_6692,N_6416,N_6090);
nand U6693 (N_6693,N_6280,N_6376);
and U6694 (N_6694,N_6230,N_6308);
nand U6695 (N_6695,N_6245,N_6307);
nor U6696 (N_6696,N_6333,N_6037);
or U6697 (N_6697,N_6436,N_6420);
and U6698 (N_6698,N_6160,N_6086);
nor U6699 (N_6699,N_6109,N_6389);
and U6700 (N_6700,N_6305,N_6145);
or U6701 (N_6701,N_6394,N_6036);
xor U6702 (N_6702,N_6133,N_6382);
nor U6703 (N_6703,N_6292,N_6009);
nand U6704 (N_6704,N_6331,N_6312);
xnor U6705 (N_6705,N_6180,N_6098);
and U6706 (N_6706,N_6136,N_6163);
and U6707 (N_6707,N_6364,N_6166);
and U6708 (N_6708,N_6244,N_6381);
or U6709 (N_6709,N_6371,N_6264);
nand U6710 (N_6710,N_6141,N_6384);
xnor U6711 (N_6711,N_6370,N_6168);
and U6712 (N_6712,N_6262,N_6001);
nand U6713 (N_6713,N_6353,N_6143);
nor U6714 (N_6714,N_6403,N_6470);
or U6715 (N_6715,N_6483,N_6102);
and U6716 (N_6716,N_6473,N_6407);
nand U6717 (N_6717,N_6031,N_6162);
or U6718 (N_6718,N_6490,N_6286);
nand U6719 (N_6719,N_6247,N_6181);
nor U6720 (N_6720,N_6378,N_6025);
xor U6721 (N_6721,N_6115,N_6048);
or U6722 (N_6722,N_6038,N_6374);
and U6723 (N_6723,N_6386,N_6006);
and U6724 (N_6724,N_6317,N_6107);
nand U6725 (N_6725,N_6218,N_6427);
nand U6726 (N_6726,N_6082,N_6390);
or U6727 (N_6727,N_6392,N_6288);
and U6728 (N_6728,N_6460,N_6240);
nor U6729 (N_6729,N_6212,N_6495);
and U6730 (N_6730,N_6325,N_6189);
and U6731 (N_6731,N_6289,N_6350);
nor U6732 (N_6732,N_6355,N_6322);
or U6733 (N_6733,N_6175,N_6396);
nand U6734 (N_6734,N_6209,N_6094);
and U6735 (N_6735,N_6058,N_6443);
or U6736 (N_6736,N_6449,N_6301);
or U6737 (N_6737,N_6493,N_6274);
or U6738 (N_6738,N_6401,N_6081);
and U6739 (N_6739,N_6125,N_6032);
nand U6740 (N_6740,N_6217,N_6491);
nand U6741 (N_6741,N_6461,N_6099);
nand U6742 (N_6742,N_6454,N_6072);
and U6743 (N_6743,N_6070,N_6398);
xor U6744 (N_6744,N_6040,N_6008);
or U6745 (N_6745,N_6351,N_6116);
nand U6746 (N_6746,N_6344,N_6126);
and U6747 (N_6747,N_6234,N_6177);
and U6748 (N_6748,N_6210,N_6270);
or U6749 (N_6749,N_6347,N_6395);
nand U6750 (N_6750,N_6463,N_6375);
nand U6751 (N_6751,N_6460,N_6499);
nor U6752 (N_6752,N_6441,N_6390);
nor U6753 (N_6753,N_6156,N_6430);
xnor U6754 (N_6754,N_6190,N_6490);
xor U6755 (N_6755,N_6211,N_6253);
or U6756 (N_6756,N_6474,N_6419);
and U6757 (N_6757,N_6265,N_6158);
nor U6758 (N_6758,N_6204,N_6289);
or U6759 (N_6759,N_6308,N_6311);
or U6760 (N_6760,N_6496,N_6003);
nand U6761 (N_6761,N_6130,N_6317);
nand U6762 (N_6762,N_6167,N_6292);
xor U6763 (N_6763,N_6319,N_6393);
nand U6764 (N_6764,N_6360,N_6332);
nor U6765 (N_6765,N_6073,N_6364);
xor U6766 (N_6766,N_6442,N_6211);
nand U6767 (N_6767,N_6187,N_6072);
and U6768 (N_6768,N_6237,N_6260);
and U6769 (N_6769,N_6075,N_6170);
xnor U6770 (N_6770,N_6056,N_6169);
or U6771 (N_6771,N_6104,N_6369);
or U6772 (N_6772,N_6480,N_6452);
and U6773 (N_6773,N_6284,N_6255);
xor U6774 (N_6774,N_6473,N_6046);
xnor U6775 (N_6775,N_6303,N_6284);
nand U6776 (N_6776,N_6016,N_6330);
nor U6777 (N_6777,N_6000,N_6230);
or U6778 (N_6778,N_6377,N_6407);
and U6779 (N_6779,N_6143,N_6412);
and U6780 (N_6780,N_6101,N_6061);
xor U6781 (N_6781,N_6466,N_6233);
or U6782 (N_6782,N_6372,N_6458);
nand U6783 (N_6783,N_6050,N_6473);
nand U6784 (N_6784,N_6242,N_6219);
nor U6785 (N_6785,N_6327,N_6077);
nor U6786 (N_6786,N_6227,N_6326);
or U6787 (N_6787,N_6090,N_6092);
and U6788 (N_6788,N_6371,N_6107);
xnor U6789 (N_6789,N_6439,N_6179);
xnor U6790 (N_6790,N_6420,N_6085);
xor U6791 (N_6791,N_6292,N_6365);
xor U6792 (N_6792,N_6130,N_6001);
nor U6793 (N_6793,N_6246,N_6009);
xor U6794 (N_6794,N_6069,N_6319);
or U6795 (N_6795,N_6016,N_6233);
and U6796 (N_6796,N_6464,N_6155);
nand U6797 (N_6797,N_6081,N_6410);
xor U6798 (N_6798,N_6125,N_6180);
xnor U6799 (N_6799,N_6319,N_6196);
xnor U6800 (N_6800,N_6414,N_6173);
nand U6801 (N_6801,N_6298,N_6372);
or U6802 (N_6802,N_6302,N_6402);
nand U6803 (N_6803,N_6129,N_6082);
or U6804 (N_6804,N_6005,N_6002);
nor U6805 (N_6805,N_6237,N_6224);
xor U6806 (N_6806,N_6379,N_6044);
nand U6807 (N_6807,N_6120,N_6469);
and U6808 (N_6808,N_6393,N_6196);
or U6809 (N_6809,N_6420,N_6017);
and U6810 (N_6810,N_6321,N_6293);
or U6811 (N_6811,N_6251,N_6098);
nand U6812 (N_6812,N_6333,N_6305);
nor U6813 (N_6813,N_6297,N_6304);
xor U6814 (N_6814,N_6327,N_6287);
xnor U6815 (N_6815,N_6274,N_6303);
xnor U6816 (N_6816,N_6079,N_6295);
and U6817 (N_6817,N_6298,N_6105);
and U6818 (N_6818,N_6195,N_6395);
and U6819 (N_6819,N_6341,N_6248);
nor U6820 (N_6820,N_6226,N_6411);
and U6821 (N_6821,N_6296,N_6054);
and U6822 (N_6822,N_6218,N_6071);
and U6823 (N_6823,N_6039,N_6305);
or U6824 (N_6824,N_6103,N_6240);
xnor U6825 (N_6825,N_6438,N_6491);
nor U6826 (N_6826,N_6068,N_6314);
nor U6827 (N_6827,N_6381,N_6254);
xor U6828 (N_6828,N_6435,N_6062);
xor U6829 (N_6829,N_6292,N_6123);
nand U6830 (N_6830,N_6143,N_6487);
xor U6831 (N_6831,N_6295,N_6313);
nand U6832 (N_6832,N_6117,N_6351);
nor U6833 (N_6833,N_6026,N_6279);
xnor U6834 (N_6834,N_6160,N_6022);
nand U6835 (N_6835,N_6348,N_6208);
or U6836 (N_6836,N_6247,N_6326);
nand U6837 (N_6837,N_6104,N_6405);
or U6838 (N_6838,N_6464,N_6137);
or U6839 (N_6839,N_6082,N_6224);
xor U6840 (N_6840,N_6099,N_6400);
xnor U6841 (N_6841,N_6314,N_6477);
nand U6842 (N_6842,N_6245,N_6305);
nand U6843 (N_6843,N_6222,N_6124);
nand U6844 (N_6844,N_6148,N_6440);
and U6845 (N_6845,N_6330,N_6277);
xor U6846 (N_6846,N_6305,N_6214);
nor U6847 (N_6847,N_6358,N_6362);
or U6848 (N_6848,N_6002,N_6204);
and U6849 (N_6849,N_6456,N_6360);
nand U6850 (N_6850,N_6084,N_6258);
or U6851 (N_6851,N_6266,N_6280);
xnor U6852 (N_6852,N_6221,N_6286);
and U6853 (N_6853,N_6493,N_6105);
and U6854 (N_6854,N_6394,N_6080);
or U6855 (N_6855,N_6285,N_6385);
or U6856 (N_6856,N_6388,N_6203);
nand U6857 (N_6857,N_6278,N_6007);
or U6858 (N_6858,N_6173,N_6321);
or U6859 (N_6859,N_6040,N_6444);
and U6860 (N_6860,N_6200,N_6262);
xor U6861 (N_6861,N_6052,N_6425);
and U6862 (N_6862,N_6161,N_6235);
nand U6863 (N_6863,N_6270,N_6154);
xor U6864 (N_6864,N_6488,N_6339);
xor U6865 (N_6865,N_6337,N_6442);
or U6866 (N_6866,N_6115,N_6326);
nor U6867 (N_6867,N_6025,N_6003);
and U6868 (N_6868,N_6336,N_6305);
or U6869 (N_6869,N_6252,N_6060);
xor U6870 (N_6870,N_6225,N_6280);
nand U6871 (N_6871,N_6415,N_6379);
nand U6872 (N_6872,N_6435,N_6203);
or U6873 (N_6873,N_6004,N_6028);
or U6874 (N_6874,N_6318,N_6394);
nor U6875 (N_6875,N_6199,N_6234);
and U6876 (N_6876,N_6457,N_6353);
nor U6877 (N_6877,N_6315,N_6159);
and U6878 (N_6878,N_6137,N_6182);
and U6879 (N_6879,N_6157,N_6471);
or U6880 (N_6880,N_6142,N_6008);
xnor U6881 (N_6881,N_6348,N_6489);
xnor U6882 (N_6882,N_6002,N_6206);
and U6883 (N_6883,N_6458,N_6229);
or U6884 (N_6884,N_6176,N_6163);
nor U6885 (N_6885,N_6363,N_6454);
nor U6886 (N_6886,N_6104,N_6110);
nand U6887 (N_6887,N_6274,N_6420);
and U6888 (N_6888,N_6397,N_6289);
nor U6889 (N_6889,N_6274,N_6204);
xor U6890 (N_6890,N_6356,N_6090);
nand U6891 (N_6891,N_6213,N_6114);
nor U6892 (N_6892,N_6385,N_6081);
xnor U6893 (N_6893,N_6036,N_6392);
nor U6894 (N_6894,N_6278,N_6214);
nor U6895 (N_6895,N_6434,N_6046);
or U6896 (N_6896,N_6432,N_6000);
xnor U6897 (N_6897,N_6461,N_6468);
nand U6898 (N_6898,N_6051,N_6129);
xnor U6899 (N_6899,N_6294,N_6122);
xor U6900 (N_6900,N_6082,N_6409);
nand U6901 (N_6901,N_6067,N_6483);
and U6902 (N_6902,N_6337,N_6343);
nand U6903 (N_6903,N_6107,N_6386);
nor U6904 (N_6904,N_6417,N_6297);
nand U6905 (N_6905,N_6234,N_6189);
xnor U6906 (N_6906,N_6050,N_6216);
nor U6907 (N_6907,N_6243,N_6137);
nand U6908 (N_6908,N_6205,N_6108);
nor U6909 (N_6909,N_6051,N_6058);
nor U6910 (N_6910,N_6231,N_6075);
and U6911 (N_6911,N_6486,N_6435);
nand U6912 (N_6912,N_6406,N_6360);
and U6913 (N_6913,N_6267,N_6178);
nand U6914 (N_6914,N_6182,N_6209);
or U6915 (N_6915,N_6126,N_6460);
xor U6916 (N_6916,N_6475,N_6252);
nand U6917 (N_6917,N_6329,N_6044);
xnor U6918 (N_6918,N_6019,N_6359);
xor U6919 (N_6919,N_6327,N_6465);
and U6920 (N_6920,N_6315,N_6018);
or U6921 (N_6921,N_6445,N_6173);
nor U6922 (N_6922,N_6384,N_6373);
and U6923 (N_6923,N_6272,N_6315);
xnor U6924 (N_6924,N_6472,N_6319);
nand U6925 (N_6925,N_6466,N_6170);
xnor U6926 (N_6926,N_6437,N_6040);
nand U6927 (N_6927,N_6307,N_6262);
xnor U6928 (N_6928,N_6183,N_6268);
and U6929 (N_6929,N_6080,N_6123);
nand U6930 (N_6930,N_6067,N_6184);
nor U6931 (N_6931,N_6157,N_6230);
or U6932 (N_6932,N_6317,N_6185);
and U6933 (N_6933,N_6109,N_6104);
nor U6934 (N_6934,N_6272,N_6342);
nor U6935 (N_6935,N_6053,N_6308);
or U6936 (N_6936,N_6046,N_6293);
and U6937 (N_6937,N_6003,N_6460);
or U6938 (N_6938,N_6120,N_6139);
or U6939 (N_6939,N_6151,N_6269);
and U6940 (N_6940,N_6225,N_6377);
nor U6941 (N_6941,N_6408,N_6145);
xor U6942 (N_6942,N_6184,N_6108);
xor U6943 (N_6943,N_6232,N_6145);
xor U6944 (N_6944,N_6087,N_6186);
nand U6945 (N_6945,N_6495,N_6139);
and U6946 (N_6946,N_6100,N_6417);
xnor U6947 (N_6947,N_6018,N_6173);
and U6948 (N_6948,N_6410,N_6045);
or U6949 (N_6949,N_6189,N_6448);
or U6950 (N_6950,N_6244,N_6141);
nand U6951 (N_6951,N_6493,N_6045);
and U6952 (N_6952,N_6049,N_6293);
nor U6953 (N_6953,N_6333,N_6151);
nand U6954 (N_6954,N_6044,N_6325);
nor U6955 (N_6955,N_6087,N_6170);
and U6956 (N_6956,N_6187,N_6292);
xnor U6957 (N_6957,N_6174,N_6060);
or U6958 (N_6958,N_6271,N_6236);
and U6959 (N_6959,N_6377,N_6111);
and U6960 (N_6960,N_6155,N_6184);
nand U6961 (N_6961,N_6071,N_6499);
or U6962 (N_6962,N_6076,N_6063);
nand U6963 (N_6963,N_6085,N_6076);
nor U6964 (N_6964,N_6312,N_6347);
xor U6965 (N_6965,N_6001,N_6478);
and U6966 (N_6966,N_6399,N_6152);
or U6967 (N_6967,N_6026,N_6314);
nor U6968 (N_6968,N_6400,N_6219);
xor U6969 (N_6969,N_6297,N_6076);
or U6970 (N_6970,N_6171,N_6095);
or U6971 (N_6971,N_6353,N_6198);
xnor U6972 (N_6972,N_6350,N_6305);
nor U6973 (N_6973,N_6175,N_6033);
and U6974 (N_6974,N_6456,N_6375);
nor U6975 (N_6975,N_6262,N_6395);
nor U6976 (N_6976,N_6019,N_6142);
nor U6977 (N_6977,N_6325,N_6489);
or U6978 (N_6978,N_6146,N_6430);
nand U6979 (N_6979,N_6212,N_6211);
xnor U6980 (N_6980,N_6128,N_6173);
and U6981 (N_6981,N_6166,N_6314);
xor U6982 (N_6982,N_6052,N_6272);
xor U6983 (N_6983,N_6045,N_6145);
nor U6984 (N_6984,N_6358,N_6005);
nor U6985 (N_6985,N_6305,N_6121);
and U6986 (N_6986,N_6100,N_6368);
or U6987 (N_6987,N_6353,N_6266);
xor U6988 (N_6988,N_6280,N_6432);
xor U6989 (N_6989,N_6489,N_6112);
and U6990 (N_6990,N_6045,N_6446);
or U6991 (N_6991,N_6433,N_6227);
or U6992 (N_6992,N_6234,N_6188);
or U6993 (N_6993,N_6134,N_6373);
and U6994 (N_6994,N_6157,N_6400);
and U6995 (N_6995,N_6127,N_6191);
nand U6996 (N_6996,N_6051,N_6309);
or U6997 (N_6997,N_6395,N_6035);
nor U6998 (N_6998,N_6486,N_6492);
and U6999 (N_6999,N_6321,N_6250);
xor U7000 (N_7000,N_6714,N_6572);
xor U7001 (N_7001,N_6820,N_6701);
and U7002 (N_7002,N_6595,N_6673);
nor U7003 (N_7003,N_6978,N_6733);
or U7004 (N_7004,N_6586,N_6767);
nor U7005 (N_7005,N_6950,N_6615);
and U7006 (N_7006,N_6598,N_6888);
nand U7007 (N_7007,N_6509,N_6954);
xor U7008 (N_7008,N_6651,N_6982);
and U7009 (N_7009,N_6793,N_6958);
xnor U7010 (N_7010,N_6623,N_6965);
nor U7011 (N_7011,N_6696,N_6530);
and U7012 (N_7012,N_6736,N_6527);
nand U7013 (N_7013,N_6859,N_6500);
nand U7014 (N_7014,N_6636,N_6578);
nor U7015 (N_7015,N_6554,N_6787);
xor U7016 (N_7016,N_6824,N_6577);
or U7017 (N_7017,N_6992,N_6920);
or U7018 (N_7018,N_6790,N_6924);
xor U7019 (N_7019,N_6908,N_6570);
or U7020 (N_7020,N_6981,N_6605);
or U7021 (N_7021,N_6743,N_6617);
and U7022 (N_7022,N_6597,N_6721);
nand U7023 (N_7023,N_6872,N_6682);
or U7024 (N_7024,N_6699,N_6875);
nand U7025 (N_7025,N_6629,N_6735);
or U7026 (N_7026,N_6678,N_6739);
xor U7027 (N_7027,N_6976,N_6728);
or U7028 (N_7028,N_6960,N_6776);
and U7029 (N_7029,N_6553,N_6877);
and U7030 (N_7030,N_6786,N_6513);
xnor U7031 (N_7031,N_6510,N_6825);
nand U7032 (N_7032,N_6907,N_6987);
xnor U7033 (N_7033,N_6983,N_6549);
and U7034 (N_7034,N_6706,N_6810);
or U7035 (N_7035,N_6634,N_6528);
xnor U7036 (N_7036,N_6945,N_6800);
nor U7037 (N_7037,N_6949,N_6871);
nand U7038 (N_7038,N_6564,N_6953);
and U7039 (N_7039,N_6775,N_6964);
nand U7040 (N_7040,N_6923,N_6971);
and U7041 (N_7041,N_6681,N_6690);
or U7042 (N_7042,N_6588,N_6635);
nor U7043 (N_7043,N_6555,N_6547);
nor U7044 (N_7044,N_6722,N_6688);
or U7045 (N_7045,N_6947,N_6752);
or U7046 (N_7046,N_6791,N_6637);
nor U7047 (N_7047,N_6503,N_6799);
or U7048 (N_7048,N_6813,N_6957);
and U7049 (N_7049,N_6990,N_6870);
nand U7050 (N_7050,N_6687,N_6977);
and U7051 (N_7051,N_6524,N_6677);
nor U7052 (N_7052,N_6993,N_6755);
nor U7053 (N_7053,N_6878,N_6779);
or U7054 (N_7054,N_6643,N_6780);
xnor U7055 (N_7055,N_6695,N_6667);
or U7056 (N_7056,N_6638,N_6656);
and U7057 (N_7057,N_6517,N_6552);
xnor U7058 (N_7058,N_6796,N_6589);
and U7059 (N_7059,N_6864,N_6904);
or U7060 (N_7060,N_6812,N_6873);
nand U7061 (N_7061,N_6898,N_6550);
or U7062 (N_7062,N_6819,N_6742);
nor U7063 (N_7063,N_6763,N_6934);
and U7064 (N_7064,N_6559,N_6841);
and U7065 (N_7065,N_6816,N_6557);
nand U7066 (N_7066,N_6565,N_6918);
or U7067 (N_7067,N_6794,N_6525);
or U7068 (N_7068,N_6846,N_6508);
xnor U7069 (N_7069,N_6838,N_6609);
xnor U7070 (N_7070,N_6862,N_6882);
xnor U7071 (N_7071,N_6737,N_6744);
nand U7072 (N_7072,N_6863,N_6808);
or U7073 (N_7073,N_6698,N_6713);
xor U7074 (N_7074,N_6631,N_6533);
and U7075 (N_7075,N_6540,N_6913);
nor U7076 (N_7076,N_6804,N_6649);
nand U7077 (N_7077,N_6658,N_6967);
xor U7078 (N_7078,N_6545,N_6647);
nand U7079 (N_7079,N_6785,N_6853);
nor U7080 (N_7080,N_6622,N_6959);
nand U7081 (N_7081,N_6546,N_6818);
nand U7082 (N_7082,N_6675,N_6917);
nor U7083 (N_7083,N_6968,N_6939);
or U7084 (N_7084,N_6703,N_6876);
or U7085 (N_7085,N_6778,N_6608);
and U7086 (N_7086,N_6581,N_6680);
xor U7087 (N_7087,N_6516,N_6847);
xnor U7088 (N_7088,N_6860,N_6828);
or U7089 (N_7089,N_6669,N_6887);
xnor U7090 (N_7090,N_6640,N_6946);
or U7091 (N_7091,N_6788,N_6966);
xnor U7092 (N_7092,N_6831,N_6769);
xnor U7093 (N_7093,N_6532,N_6973);
and U7094 (N_7094,N_6940,N_6972);
xnor U7095 (N_7095,N_6844,N_6732);
nand U7096 (N_7096,N_6970,N_6895);
or U7097 (N_7097,N_6580,N_6995);
nor U7098 (N_7098,N_6770,N_6576);
or U7099 (N_7099,N_6782,N_6584);
or U7100 (N_7100,N_6852,N_6627);
nand U7101 (N_7101,N_6806,N_6618);
or U7102 (N_7102,N_6760,N_6865);
or U7103 (N_7103,N_6988,N_6541);
xnor U7104 (N_7104,N_6952,N_6792);
or U7105 (N_7105,N_6817,N_6543);
nand U7106 (N_7106,N_6511,N_6684);
and U7107 (N_7107,N_6807,N_6891);
xor U7108 (N_7108,N_6653,N_6815);
nor U7109 (N_7109,N_6512,N_6544);
and U7110 (N_7110,N_6884,N_6826);
nand U7111 (N_7111,N_6539,N_6676);
nor U7112 (N_7112,N_6910,N_6975);
and U7113 (N_7113,N_6842,N_6520);
nor U7114 (N_7114,N_6652,N_6630);
nand U7115 (N_7115,N_6845,N_6628);
or U7116 (N_7116,N_6674,N_6936);
and U7117 (N_7117,N_6521,N_6625);
and U7118 (N_7118,N_6601,N_6811);
nand U7119 (N_7119,N_6648,N_6849);
or U7120 (N_7120,N_6611,N_6955);
and U7121 (N_7121,N_6592,N_6963);
xnor U7122 (N_7122,N_6603,N_6585);
and U7123 (N_7123,N_6663,N_6748);
nor U7124 (N_7124,N_6612,N_6626);
or U7125 (N_7125,N_6566,N_6919);
nand U7126 (N_7126,N_6768,N_6777);
and U7127 (N_7127,N_6890,N_6747);
xor U7128 (N_7128,N_6902,N_6996);
or U7129 (N_7129,N_6542,N_6504);
nand U7130 (N_7130,N_6602,N_6644);
nor U7131 (N_7131,N_6537,N_6929);
nor U7132 (N_7132,N_6892,N_6814);
nand U7133 (N_7133,N_6914,N_6507);
and U7134 (N_7134,N_6938,N_6518);
and U7135 (N_7135,N_6843,N_6839);
nand U7136 (N_7136,N_6702,N_6754);
and U7137 (N_7137,N_6932,N_6789);
nor U7138 (N_7138,N_6764,N_6740);
and U7139 (N_7139,N_6704,N_6762);
xor U7140 (N_7140,N_6526,N_6632);
or U7141 (N_7141,N_6725,N_6986);
xnor U7142 (N_7142,N_6874,N_6717);
and U7143 (N_7143,N_6896,N_6691);
nand U7144 (N_7144,N_6650,N_6579);
xnor U7145 (N_7145,N_6915,N_6529);
nand U7146 (N_7146,N_6997,N_6869);
and U7147 (N_7147,N_6858,N_6994);
nor U7148 (N_7148,N_6784,N_6620);
nor U7149 (N_7149,N_6671,N_6999);
nor U7150 (N_7150,N_6686,N_6519);
xor U7151 (N_7151,N_6587,N_6829);
xor U7152 (N_7152,N_6745,N_6604);
xnor U7153 (N_7153,N_6944,N_6837);
nor U7154 (N_7154,N_6948,N_6591);
nand U7155 (N_7155,N_6772,N_6607);
nand U7156 (N_7156,N_6501,N_6633);
nor U7157 (N_7157,N_6962,N_6989);
or U7158 (N_7158,N_6548,N_6880);
nand U7159 (N_7159,N_6606,N_6912);
or U7160 (N_7160,N_6646,N_6998);
or U7161 (N_7161,N_6855,N_6921);
nand U7162 (N_7162,N_6720,N_6573);
xor U7163 (N_7163,N_6942,N_6613);
and U7164 (N_7164,N_6710,N_6505);
xnor U7165 (N_7165,N_6645,N_6594);
nand U7166 (N_7166,N_6734,N_6803);
and U7167 (N_7167,N_6832,N_6502);
nand U7168 (N_7168,N_6655,N_6935);
nor U7169 (N_7169,N_6668,N_6657);
xor U7170 (N_7170,N_6905,N_6823);
and U7171 (N_7171,N_6596,N_6582);
nor U7172 (N_7172,N_6773,N_6802);
or U7173 (N_7173,N_6980,N_6761);
xor U7174 (N_7174,N_6991,N_6750);
nor U7175 (N_7175,N_6569,N_6746);
xnor U7176 (N_7176,N_6535,N_6759);
nand U7177 (N_7177,N_6883,N_6700);
xor U7178 (N_7178,N_6599,N_6719);
xor U7179 (N_7179,N_6639,N_6619);
and U7180 (N_7180,N_6903,N_6600);
xor U7181 (N_7181,N_6538,N_6900);
xnor U7182 (N_7182,N_6941,N_6834);
and U7183 (N_7183,N_6560,N_6621);
or U7184 (N_7184,N_6556,N_6765);
or U7185 (N_7185,N_6563,N_6795);
nand U7186 (N_7186,N_6689,N_6897);
or U7187 (N_7187,N_6567,N_6709);
or U7188 (N_7188,N_6575,N_6729);
or U7189 (N_7189,N_6916,N_6536);
and U7190 (N_7190,N_6672,N_6801);
nor U7191 (N_7191,N_6665,N_6984);
or U7192 (N_7192,N_6659,N_6705);
xnor U7193 (N_7193,N_6979,N_6711);
nand U7194 (N_7194,N_6766,N_6901);
xnor U7195 (N_7195,N_6835,N_6857);
nor U7196 (N_7196,N_6868,N_6783);
xnor U7197 (N_7197,N_6827,N_6753);
or U7198 (N_7198,N_6583,N_6666);
or U7199 (N_7199,N_6985,N_6757);
nor U7200 (N_7200,N_6833,N_6894);
nand U7201 (N_7201,N_6731,N_6889);
or U7202 (N_7202,N_6679,N_6642);
or U7203 (N_7203,N_6574,N_6534);
xnor U7204 (N_7204,N_6809,N_6523);
xnor U7205 (N_7205,N_6723,N_6693);
xnor U7206 (N_7206,N_6571,N_6797);
nand U7207 (N_7207,N_6562,N_6848);
nand U7208 (N_7208,N_6641,N_6692);
nor U7209 (N_7209,N_6751,N_6683);
nor U7210 (N_7210,N_6707,N_6856);
or U7211 (N_7211,N_6911,N_6593);
and U7212 (N_7212,N_6726,N_6610);
xnor U7213 (N_7213,N_6718,N_6730);
or U7214 (N_7214,N_6926,N_6738);
and U7215 (N_7215,N_6774,N_6624);
or U7216 (N_7216,N_6798,N_6616);
nor U7217 (N_7217,N_6660,N_6879);
nand U7218 (N_7218,N_6937,N_6771);
nor U7219 (N_7219,N_6531,N_6506);
xnor U7220 (N_7220,N_6727,N_6781);
nor U7221 (N_7221,N_6851,N_6861);
or U7222 (N_7222,N_6850,N_6712);
xnor U7223 (N_7223,N_6925,N_6974);
nand U7224 (N_7224,N_6956,N_6885);
nor U7225 (N_7225,N_6694,N_6933);
nor U7226 (N_7226,N_6724,N_6836);
xnor U7227 (N_7227,N_6922,N_6951);
nand U7228 (N_7228,N_6715,N_6685);
nor U7229 (N_7229,N_6822,N_6830);
and U7230 (N_7230,N_6961,N_6906);
xnor U7231 (N_7231,N_6558,N_6840);
and U7232 (N_7232,N_6662,N_6881);
xnor U7233 (N_7233,N_6930,N_6590);
and U7234 (N_7234,N_6758,N_6697);
nand U7235 (N_7235,N_6670,N_6909);
nand U7236 (N_7236,N_6514,N_6561);
nand U7237 (N_7237,N_6931,N_6821);
nand U7238 (N_7238,N_6899,N_6886);
and U7239 (N_7239,N_6568,N_6927);
and U7240 (N_7240,N_6893,N_6664);
nand U7241 (N_7241,N_6928,N_6614);
or U7242 (N_7242,N_6805,N_6708);
xnor U7243 (N_7243,N_6867,N_6654);
xor U7244 (N_7244,N_6866,N_6741);
nand U7245 (N_7245,N_6969,N_6749);
xnor U7246 (N_7246,N_6756,N_6716);
nand U7247 (N_7247,N_6854,N_6515);
nand U7248 (N_7248,N_6943,N_6551);
and U7249 (N_7249,N_6661,N_6522);
xor U7250 (N_7250,N_6518,N_6946);
nand U7251 (N_7251,N_6726,N_6557);
xnor U7252 (N_7252,N_6881,N_6549);
nor U7253 (N_7253,N_6949,N_6944);
and U7254 (N_7254,N_6729,N_6720);
and U7255 (N_7255,N_6617,N_6796);
and U7256 (N_7256,N_6883,N_6637);
nand U7257 (N_7257,N_6749,N_6663);
nor U7258 (N_7258,N_6738,N_6629);
and U7259 (N_7259,N_6814,N_6592);
xnor U7260 (N_7260,N_6510,N_6963);
or U7261 (N_7261,N_6609,N_6643);
xnor U7262 (N_7262,N_6675,N_6639);
nor U7263 (N_7263,N_6728,N_6540);
or U7264 (N_7264,N_6828,N_6554);
and U7265 (N_7265,N_6715,N_6615);
xor U7266 (N_7266,N_6909,N_6682);
and U7267 (N_7267,N_6902,N_6600);
or U7268 (N_7268,N_6968,N_6792);
and U7269 (N_7269,N_6575,N_6644);
or U7270 (N_7270,N_6980,N_6740);
and U7271 (N_7271,N_6894,N_6523);
and U7272 (N_7272,N_6828,N_6545);
nand U7273 (N_7273,N_6822,N_6939);
nand U7274 (N_7274,N_6660,N_6509);
nand U7275 (N_7275,N_6538,N_6929);
nand U7276 (N_7276,N_6985,N_6865);
nor U7277 (N_7277,N_6628,N_6876);
xnor U7278 (N_7278,N_6604,N_6946);
and U7279 (N_7279,N_6536,N_6978);
nand U7280 (N_7280,N_6834,N_6959);
xor U7281 (N_7281,N_6863,N_6750);
xor U7282 (N_7282,N_6571,N_6808);
nor U7283 (N_7283,N_6942,N_6770);
nor U7284 (N_7284,N_6686,N_6533);
nand U7285 (N_7285,N_6885,N_6753);
nand U7286 (N_7286,N_6724,N_6717);
nand U7287 (N_7287,N_6787,N_6973);
or U7288 (N_7288,N_6842,N_6704);
nor U7289 (N_7289,N_6774,N_6886);
nand U7290 (N_7290,N_6726,N_6503);
or U7291 (N_7291,N_6785,N_6838);
nor U7292 (N_7292,N_6503,N_6755);
xor U7293 (N_7293,N_6821,N_6765);
nand U7294 (N_7294,N_6546,N_6701);
nor U7295 (N_7295,N_6622,N_6879);
xnor U7296 (N_7296,N_6861,N_6676);
and U7297 (N_7297,N_6502,N_6613);
nand U7298 (N_7298,N_6544,N_6876);
or U7299 (N_7299,N_6523,N_6695);
nor U7300 (N_7300,N_6561,N_6922);
or U7301 (N_7301,N_6713,N_6610);
and U7302 (N_7302,N_6867,N_6990);
and U7303 (N_7303,N_6692,N_6856);
nand U7304 (N_7304,N_6594,N_6955);
and U7305 (N_7305,N_6514,N_6848);
nor U7306 (N_7306,N_6975,N_6713);
or U7307 (N_7307,N_6740,N_6876);
nand U7308 (N_7308,N_6539,N_6911);
nor U7309 (N_7309,N_6560,N_6654);
or U7310 (N_7310,N_6842,N_6746);
nor U7311 (N_7311,N_6679,N_6535);
nor U7312 (N_7312,N_6578,N_6781);
nor U7313 (N_7313,N_6691,N_6642);
nand U7314 (N_7314,N_6913,N_6510);
or U7315 (N_7315,N_6906,N_6874);
and U7316 (N_7316,N_6860,N_6662);
or U7317 (N_7317,N_6882,N_6815);
nand U7318 (N_7318,N_6766,N_6657);
xnor U7319 (N_7319,N_6502,N_6528);
or U7320 (N_7320,N_6601,N_6985);
nand U7321 (N_7321,N_6717,N_6981);
nand U7322 (N_7322,N_6819,N_6674);
and U7323 (N_7323,N_6623,N_6969);
or U7324 (N_7324,N_6843,N_6959);
nand U7325 (N_7325,N_6651,N_6526);
nand U7326 (N_7326,N_6858,N_6708);
xnor U7327 (N_7327,N_6508,N_6996);
nor U7328 (N_7328,N_6875,N_6818);
or U7329 (N_7329,N_6940,N_6811);
nor U7330 (N_7330,N_6661,N_6821);
and U7331 (N_7331,N_6913,N_6649);
nor U7332 (N_7332,N_6978,N_6644);
and U7333 (N_7333,N_6758,N_6946);
nand U7334 (N_7334,N_6583,N_6760);
nand U7335 (N_7335,N_6847,N_6522);
xnor U7336 (N_7336,N_6705,N_6822);
nand U7337 (N_7337,N_6545,N_6724);
or U7338 (N_7338,N_6954,N_6681);
nor U7339 (N_7339,N_6573,N_6886);
xor U7340 (N_7340,N_6507,N_6930);
nor U7341 (N_7341,N_6637,N_6806);
or U7342 (N_7342,N_6862,N_6554);
or U7343 (N_7343,N_6998,N_6805);
or U7344 (N_7344,N_6804,N_6680);
nand U7345 (N_7345,N_6594,N_6623);
nand U7346 (N_7346,N_6954,N_6890);
nor U7347 (N_7347,N_6533,N_6725);
or U7348 (N_7348,N_6926,N_6837);
nor U7349 (N_7349,N_6733,N_6972);
and U7350 (N_7350,N_6782,N_6656);
and U7351 (N_7351,N_6605,N_6789);
and U7352 (N_7352,N_6969,N_6934);
and U7353 (N_7353,N_6761,N_6748);
xor U7354 (N_7354,N_6994,N_6766);
or U7355 (N_7355,N_6940,N_6647);
xor U7356 (N_7356,N_6701,N_6609);
nor U7357 (N_7357,N_6987,N_6787);
and U7358 (N_7358,N_6967,N_6913);
nor U7359 (N_7359,N_6756,N_6667);
and U7360 (N_7360,N_6998,N_6865);
and U7361 (N_7361,N_6707,N_6512);
xnor U7362 (N_7362,N_6890,N_6591);
and U7363 (N_7363,N_6893,N_6762);
nand U7364 (N_7364,N_6572,N_6541);
or U7365 (N_7365,N_6987,N_6744);
xnor U7366 (N_7366,N_6653,N_6591);
nor U7367 (N_7367,N_6589,N_6661);
nand U7368 (N_7368,N_6726,N_6773);
or U7369 (N_7369,N_6959,N_6627);
nand U7370 (N_7370,N_6606,N_6501);
xnor U7371 (N_7371,N_6752,N_6903);
xor U7372 (N_7372,N_6607,N_6506);
nor U7373 (N_7373,N_6900,N_6848);
or U7374 (N_7374,N_6924,N_6888);
and U7375 (N_7375,N_6729,N_6524);
xnor U7376 (N_7376,N_6860,N_6973);
and U7377 (N_7377,N_6590,N_6502);
and U7378 (N_7378,N_6559,N_6684);
xnor U7379 (N_7379,N_6632,N_6633);
nand U7380 (N_7380,N_6590,N_6804);
nor U7381 (N_7381,N_6620,N_6656);
and U7382 (N_7382,N_6783,N_6799);
xnor U7383 (N_7383,N_6742,N_6585);
xnor U7384 (N_7384,N_6730,N_6875);
xor U7385 (N_7385,N_6582,N_6576);
and U7386 (N_7386,N_6521,N_6678);
nor U7387 (N_7387,N_6744,N_6640);
nand U7388 (N_7388,N_6631,N_6874);
nand U7389 (N_7389,N_6904,N_6901);
nor U7390 (N_7390,N_6509,N_6568);
nand U7391 (N_7391,N_6928,N_6981);
xnor U7392 (N_7392,N_6796,N_6713);
nand U7393 (N_7393,N_6835,N_6774);
nor U7394 (N_7394,N_6643,N_6834);
nor U7395 (N_7395,N_6571,N_6795);
or U7396 (N_7396,N_6652,N_6539);
and U7397 (N_7397,N_6954,N_6813);
nor U7398 (N_7398,N_6858,N_6976);
xor U7399 (N_7399,N_6773,N_6610);
nand U7400 (N_7400,N_6564,N_6703);
nor U7401 (N_7401,N_6521,N_6550);
xnor U7402 (N_7402,N_6691,N_6583);
nand U7403 (N_7403,N_6787,N_6663);
and U7404 (N_7404,N_6768,N_6583);
or U7405 (N_7405,N_6673,N_6828);
and U7406 (N_7406,N_6726,N_6608);
nand U7407 (N_7407,N_6892,N_6620);
xor U7408 (N_7408,N_6899,N_6624);
nand U7409 (N_7409,N_6789,N_6764);
xnor U7410 (N_7410,N_6782,N_6997);
nand U7411 (N_7411,N_6881,N_6651);
nor U7412 (N_7412,N_6636,N_6918);
nand U7413 (N_7413,N_6862,N_6679);
nand U7414 (N_7414,N_6994,N_6838);
nand U7415 (N_7415,N_6727,N_6944);
or U7416 (N_7416,N_6800,N_6898);
nor U7417 (N_7417,N_6989,N_6779);
or U7418 (N_7418,N_6995,N_6851);
or U7419 (N_7419,N_6972,N_6695);
or U7420 (N_7420,N_6920,N_6970);
nor U7421 (N_7421,N_6559,N_6820);
or U7422 (N_7422,N_6718,N_6664);
and U7423 (N_7423,N_6566,N_6771);
xor U7424 (N_7424,N_6801,N_6643);
nand U7425 (N_7425,N_6783,N_6949);
nor U7426 (N_7426,N_6871,N_6959);
and U7427 (N_7427,N_6909,N_6637);
and U7428 (N_7428,N_6870,N_6988);
or U7429 (N_7429,N_6841,N_6968);
xnor U7430 (N_7430,N_6549,N_6555);
and U7431 (N_7431,N_6507,N_6961);
nor U7432 (N_7432,N_6690,N_6612);
nor U7433 (N_7433,N_6825,N_6737);
xnor U7434 (N_7434,N_6744,N_6977);
xor U7435 (N_7435,N_6895,N_6807);
nand U7436 (N_7436,N_6724,N_6866);
or U7437 (N_7437,N_6653,N_6742);
xor U7438 (N_7438,N_6889,N_6516);
and U7439 (N_7439,N_6784,N_6779);
or U7440 (N_7440,N_6587,N_6500);
or U7441 (N_7441,N_6637,N_6932);
nor U7442 (N_7442,N_6751,N_6554);
xor U7443 (N_7443,N_6706,N_6967);
or U7444 (N_7444,N_6987,N_6888);
nand U7445 (N_7445,N_6896,N_6614);
or U7446 (N_7446,N_6988,N_6673);
or U7447 (N_7447,N_6908,N_6888);
or U7448 (N_7448,N_6808,N_6911);
or U7449 (N_7449,N_6781,N_6618);
nor U7450 (N_7450,N_6702,N_6675);
nand U7451 (N_7451,N_6852,N_6767);
nand U7452 (N_7452,N_6597,N_6912);
nand U7453 (N_7453,N_6852,N_6920);
and U7454 (N_7454,N_6782,N_6917);
nor U7455 (N_7455,N_6976,N_6793);
nand U7456 (N_7456,N_6837,N_6590);
and U7457 (N_7457,N_6628,N_6658);
and U7458 (N_7458,N_6625,N_6777);
or U7459 (N_7459,N_6692,N_6616);
nand U7460 (N_7460,N_6862,N_6888);
nor U7461 (N_7461,N_6614,N_6951);
xor U7462 (N_7462,N_6863,N_6960);
or U7463 (N_7463,N_6698,N_6756);
nand U7464 (N_7464,N_6903,N_6981);
xor U7465 (N_7465,N_6914,N_6508);
nor U7466 (N_7466,N_6962,N_6601);
xor U7467 (N_7467,N_6618,N_6940);
nor U7468 (N_7468,N_6612,N_6598);
xnor U7469 (N_7469,N_6965,N_6565);
nor U7470 (N_7470,N_6995,N_6882);
nand U7471 (N_7471,N_6772,N_6642);
xor U7472 (N_7472,N_6806,N_6697);
xor U7473 (N_7473,N_6756,N_6556);
and U7474 (N_7474,N_6594,N_6905);
nand U7475 (N_7475,N_6654,N_6752);
and U7476 (N_7476,N_6969,N_6602);
nand U7477 (N_7477,N_6959,N_6720);
xnor U7478 (N_7478,N_6706,N_6538);
or U7479 (N_7479,N_6585,N_6581);
or U7480 (N_7480,N_6871,N_6847);
nand U7481 (N_7481,N_6501,N_6934);
nor U7482 (N_7482,N_6964,N_6998);
nor U7483 (N_7483,N_6865,N_6903);
and U7484 (N_7484,N_6565,N_6661);
and U7485 (N_7485,N_6545,N_6771);
xnor U7486 (N_7486,N_6586,N_6840);
or U7487 (N_7487,N_6795,N_6741);
nand U7488 (N_7488,N_6979,N_6713);
nor U7489 (N_7489,N_6668,N_6727);
xnor U7490 (N_7490,N_6709,N_6996);
or U7491 (N_7491,N_6663,N_6693);
and U7492 (N_7492,N_6735,N_6832);
nand U7493 (N_7493,N_6695,N_6745);
or U7494 (N_7494,N_6813,N_6947);
nand U7495 (N_7495,N_6561,N_6767);
xor U7496 (N_7496,N_6966,N_6690);
and U7497 (N_7497,N_6868,N_6538);
xor U7498 (N_7498,N_6958,N_6601);
nand U7499 (N_7499,N_6954,N_6846);
nand U7500 (N_7500,N_7468,N_7090);
nor U7501 (N_7501,N_7000,N_7247);
nor U7502 (N_7502,N_7458,N_7404);
xnor U7503 (N_7503,N_7444,N_7215);
nor U7504 (N_7504,N_7153,N_7199);
nor U7505 (N_7505,N_7350,N_7167);
and U7506 (N_7506,N_7355,N_7335);
nand U7507 (N_7507,N_7193,N_7138);
nand U7508 (N_7508,N_7222,N_7329);
nor U7509 (N_7509,N_7409,N_7460);
xnor U7510 (N_7510,N_7428,N_7139);
nand U7511 (N_7511,N_7319,N_7175);
and U7512 (N_7512,N_7192,N_7146);
nor U7513 (N_7513,N_7183,N_7361);
or U7514 (N_7514,N_7011,N_7191);
or U7515 (N_7515,N_7122,N_7379);
nor U7516 (N_7516,N_7418,N_7165);
nor U7517 (N_7517,N_7328,N_7145);
xnor U7518 (N_7518,N_7053,N_7268);
or U7519 (N_7519,N_7026,N_7063);
or U7520 (N_7520,N_7180,N_7318);
nand U7521 (N_7521,N_7315,N_7030);
or U7522 (N_7522,N_7432,N_7367);
xor U7523 (N_7523,N_7473,N_7278);
nand U7524 (N_7524,N_7024,N_7203);
nand U7525 (N_7525,N_7486,N_7491);
and U7526 (N_7526,N_7250,N_7414);
nor U7527 (N_7527,N_7371,N_7225);
and U7528 (N_7528,N_7457,N_7112);
nor U7529 (N_7529,N_7287,N_7077);
nor U7530 (N_7530,N_7382,N_7127);
and U7531 (N_7531,N_7185,N_7177);
nor U7532 (N_7532,N_7440,N_7244);
nand U7533 (N_7533,N_7010,N_7277);
nor U7534 (N_7534,N_7331,N_7378);
and U7535 (N_7535,N_7014,N_7128);
nor U7536 (N_7536,N_7320,N_7370);
nor U7537 (N_7537,N_7276,N_7241);
xnor U7538 (N_7538,N_7248,N_7263);
and U7539 (N_7539,N_7495,N_7448);
and U7540 (N_7540,N_7304,N_7240);
nand U7541 (N_7541,N_7195,N_7072);
or U7542 (N_7542,N_7364,N_7303);
xor U7543 (N_7543,N_7060,N_7123);
xor U7544 (N_7544,N_7237,N_7269);
nand U7545 (N_7545,N_7197,N_7478);
or U7546 (N_7546,N_7251,N_7252);
or U7547 (N_7547,N_7305,N_7462);
and U7548 (N_7548,N_7156,N_7299);
nor U7549 (N_7549,N_7254,N_7200);
xnor U7550 (N_7550,N_7298,N_7366);
nor U7551 (N_7551,N_7217,N_7333);
nand U7552 (N_7552,N_7066,N_7451);
xnor U7553 (N_7553,N_7372,N_7330);
nand U7554 (N_7554,N_7051,N_7037);
and U7555 (N_7555,N_7293,N_7079);
nand U7556 (N_7556,N_7392,N_7282);
or U7557 (N_7557,N_7407,N_7004);
and U7558 (N_7558,N_7336,N_7463);
nor U7559 (N_7559,N_7201,N_7442);
nand U7560 (N_7560,N_7308,N_7196);
xor U7561 (N_7561,N_7226,N_7424);
nor U7562 (N_7562,N_7006,N_7106);
and U7563 (N_7563,N_7322,N_7068);
xnor U7564 (N_7564,N_7365,N_7098);
or U7565 (N_7565,N_7485,N_7403);
nor U7566 (N_7566,N_7040,N_7357);
and U7567 (N_7567,N_7398,N_7313);
and U7568 (N_7568,N_7005,N_7074);
nor U7569 (N_7569,N_7291,N_7317);
nor U7570 (N_7570,N_7290,N_7160);
nor U7571 (N_7571,N_7441,N_7162);
nor U7572 (N_7572,N_7323,N_7255);
and U7573 (N_7573,N_7274,N_7016);
xor U7574 (N_7574,N_7121,N_7373);
or U7575 (N_7575,N_7102,N_7368);
nor U7576 (N_7576,N_7129,N_7267);
xnor U7577 (N_7577,N_7389,N_7301);
and U7578 (N_7578,N_7309,N_7345);
or U7579 (N_7579,N_7342,N_7397);
nor U7580 (N_7580,N_7143,N_7114);
nor U7581 (N_7581,N_7085,N_7474);
xor U7582 (N_7582,N_7232,N_7429);
nor U7583 (N_7583,N_7209,N_7271);
xnor U7584 (N_7584,N_7411,N_7047);
and U7585 (N_7585,N_7234,N_7352);
nor U7586 (N_7586,N_7480,N_7136);
xnor U7587 (N_7587,N_7360,N_7294);
nand U7588 (N_7588,N_7246,N_7111);
nand U7589 (N_7589,N_7093,N_7369);
and U7590 (N_7590,N_7224,N_7281);
or U7591 (N_7591,N_7386,N_7339);
xnor U7592 (N_7592,N_7029,N_7038);
xor U7593 (N_7593,N_7067,N_7101);
and U7594 (N_7594,N_7083,N_7300);
nand U7595 (N_7595,N_7306,N_7097);
or U7596 (N_7596,N_7264,N_7494);
nand U7597 (N_7597,N_7384,N_7110);
and U7598 (N_7598,N_7438,N_7376);
nor U7599 (N_7599,N_7058,N_7481);
nor U7600 (N_7600,N_7338,N_7270);
and U7601 (N_7601,N_7140,N_7316);
nor U7602 (N_7602,N_7163,N_7210);
and U7603 (N_7603,N_7169,N_7283);
xnor U7604 (N_7604,N_7344,N_7184);
or U7605 (N_7605,N_7325,N_7132);
or U7606 (N_7606,N_7326,N_7166);
nor U7607 (N_7607,N_7479,N_7449);
and U7608 (N_7608,N_7099,N_7483);
and U7609 (N_7609,N_7312,N_7109);
xnor U7610 (N_7610,N_7311,N_7340);
or U7611 (N_7611,N_7158,N_7425);
and U7612 (N_7612,N_7235,N_7289);
or U7613 (N_7613,N_7141,N_7296);
xnor U7614 (N_7614,N_7455,N_7057);
and U7615 (N_7615,N_7133,N_7050);
nor U7616 (N_7616,N_7154,N_7266);
and U7617 (N_7617,N_7108,N_7170);
or U7618 (N_7618,N_7456,N_7332);
nor U7619 (N_7619,N_7280,N_7260);
and U7620 (N_7620,N_7236,N_7008);
or U7621 (N_7621,N_7159,N_7190);
nor U7622 (N_7622,N_7454,N_7238);
or U7623 (N_7623,N_7437,N_7061);
or U7624 (N_7624,N_7064,N_7374);
nand U7625 (N_7625,N_7214,N_7076);
and U7626 (N_7626,N_7489,N_7490);
or U7627 (N_7627,N_7406,N_7436);
or U7628 (N_7628,N_7233,N_7484);
nor U7629 (N_7629,N_7383,N_7487);
nor U7630 (N_7630,N_7095,N_7105);
nor U7631 (N_7631,N_7206,N_7245);
and U7632 (N_7632,N_7080,N_7034);
nor U7633 (N_7633,N_7033,N_7186);
nand U7634 (N_7634,N_7261,N_7086);
nand U7635 (N_7635,N_7262,N_7205);
nor U7636 (N_7636,N_7001,N_7243);
nand U7637 (N_7637,N_7465,N_7045);
and U7638 (N_7638,N_7116,N_7354);
and U7639 (N_7639,N_7459,N_7092);
nor U7640 (N_7640,N_7426,N_7477);
nor U7641 (N_7641,N_7071,N_7035);
xnor U7642 (N_7642,N_7015,N_7178);
or U7643 (N_7643,N_7118,N_7216);
or U7644 (N_7644,N_7211,N_7385);
nor U7645 (N_7645,N_7279,N_7272);
or U7646 (N_7646,N_7430,N_7391);
or U7647 (N_7647,N_7131,N_7130);
and U7648 (N_7648,N_7493,N_7229);
nand U7649 (N_7649,N_7288,N_7221);
and U7650 (N_7650,N_7137,N_7410);
nor U7651 (N_7651,N_7019,N_7416);
xor U7652 (N_7652,N_7189,N_7117);
nand U7653 (N_7653,N_7218,N_7075);
xnor U7654 (N_7654,N_7171,N_7452);
nand U7655 (N_7655,N_7120,N_7394);
or U7656 (N_7656,N_7073,N_7400);
xor U7657 (N_7657,N_7179,N_7334);
nor U7658 (N_7658,N_7343,N_7056);
nor U7659 (N_7659,N_7401,N_7124);
and U7660 (N_7660,N_7049,N_7087);
xnor U7661 (N_7661,N_7198,N_7230);
or U7662 (N_7662,N_7273,N_7070);
nand U7663 (N_7663,N_7302,N_7052);
nand U7664 (N_7664,N_7393,N_7027);
nand U7665 (N_7665,N_7395,N_7445);
xnor U7666 (N_7666,N_7464,N_7062);
or U7667 (N_7667,N_7249,N_7161);
nor U7668 (N_7668,N_7054,N_7482);
xnor U7669 (N_7669,N_7084,N_7018);
or U7670 (N_7670,N_7256,N_7443);
nor U7671 (N_7671,N_7172,N_7174);
and U7672 (N_7672,N_7337,N_7496);
xor U7673 (N_7673,N_7275,N_7492);
xnor U7674 (N_7674,N_7155,N_7324);
and U7675 (N_7675,N_7286,N_7469);
nor U7676 (N_7676,N_7498,N_7023);
nand U7677 (N_7677,N_7119,N_7147);
xnor U7678 (N_7678,N_7002,N_7427);
and U7679 (N_7679,N_7497,N_7041);
or U7680 (N_7680,N_7048,N_7134);
nand U7681 (N_7681,N_7349,N_7025);
nor U7682 (N_7682,N_7212,N_7013);
and U7683 (N_7683,N_7447,N_7188);
nand U7684 (N_7684,N_7433,N_7009);
xor U7685 (N_7685,N_7113,N_7055);
xnor U7686 (N_7686,N_7152,N_7021);
or U7687 (N_7687,N_7100,N_7126);
xor U7688 (N_7688,N_7078,N_7346);
xor U7689 (N_7689,N_7380,N_7341);
xor U7690 (N_7690,N_7377,N_7069);
nand U7691 (N_7691,N_7204,N_7297);
nor U7692 (N_7692,N_7417,N_7043);
nor U7693 (N_7693,N_7168,N_7164);
or U7694 (N_7694,N_7450,N_7347);
nand U7695 (N_7695,N_7042,N_7327);
or U7696 (N_7696,N_7017,N_7423);
nand U7697 (N_7697,N_7434,N_7413);
or U7698 (N_7698,N_7356,N_7007);
nand U7699 (N_7699,N_7307,N_7399);
nand U7700 (N_7700,N_7157,N_7499);
and U7701 (N_7701,N_7476,N_7292);
or U7702 (N_7702,N_7223,N_7096);
and U7703 (N_7703,N_7031,N_7470);
nand U7704 (N_7704,N_7135,N_7396);
xor U7705 (N_7705,N_7419,N_7036);
and U7706 (N_7706,N_7089,N_7351);
nand U7707 (N_7707,N_7231,N_7151);
or U7708 (N_7708,N_7412,N_7453);
xnor U7709 (N_7709,N_7358,N_7435);
and U7710 (N_7710,N_7348,N_7421);
xnor U7711 (N_7711,N_7115,N_7181);
nor U7712 (N_7712,N_7461,N_7022);
nor U7713 (N_7713,N_7020,N_7388);
nor U7714 (N_7714,N_7488,N_7295);
and U7715 (N_7715,N_7353,N_7439);
or U7716 (N_7716,N_7239,N_7142);
or U7717 (N_7717,N_7032,N_7202);
xnor U7718 (N_7718,N_7359,N_7094);
nor U7719 (N_7719,N_7472,N_7173);
and U7720 (N_7720,N_7059,N_7107);
or U7721 (N_7721,N_7242,N_7284);
xor U7722 (N_7722,N_7381,N_7467);
xnor U7723 (N_7723,N_7228,N_7375);
xnor U7724 (N_7724,N_7402,N_7253);
and U7725 (N_7725,N_7431,N_7285);
or U7726 (N_7726,N_7321,N_7471);
nor U7727 (N_7727,N_7104,N_7257);
and U7728 (N_7728,N_7422,N_7265);
xnor U7729 (N_7729,N_7028,N_7103);
and U7730 (N_7730,N_7149,N_7259);
nor U7731 (N_7731,N_7310,N_7208);
nor U7732 (N_7732,N_7082,N_7390);
and U7733 (N_7733,N_7219,N_7408);
or U7734 (N_7734,N_7446,N_7125);
xor U7735 (N_7735,N_7220,N_7387);
xor U7736 (N_7736,N_7207,N_7187);
or U7737 (N_7737,N_7213,N_7012);
and U7738 (N_7738,N_7258,N_7466);
nand U7739 (N_7739,N_7144,N_7314);
and U7740 (N_7740,N_7405,N_7182);
or U7741 (N_7741,N_7088,N_7148);
xor U7742 (N_7742,N_7046,N_7150);
xnor U7743 (N_7743,N_7363,N_7039);
nand U7744 (N_7744,N_7475,N_7362);
or U7745 (N_7745,N_7227,N_7415);
or U7746 (N_7746,N_7065,N_7081);
nand U7747 (N_7747,N_7194,N_7091);
nand U7748 (N_7748,N_7176,N_7044);
nand U7749 (N_7749,N_7003,N_7420);
nand U7750 (N_7750,N_7372,N_7002);
or U7751 (N_7751,N_7409,N_7152);
or U7752 (N_7752,N_7373,N_7140);
nand U7753 (N_7753,N_7116,N_7016);
xor U7754 (N_7754,N_7408,N_7189);
or U7755 (N_7755,N_7482,N_7151);
nor U7756 (N_7756,N_7045,N_7479);
nor U7757 (N_7757,N_7445,N_7011);
or U7758 (N_7758,N_7454,N_7445);
nor U7759 (N_7759,N_7019,N_7261);
or U7760 (N_7760,N_7361,N_7138);
xnor U7761 (N_7761,N_7169,N_7422);
and U7762 (N_7762,N_7413,N_7346);
or U7763 (N_7763,N_7454,N_7245);
nor U7764 (N_7764,N_7168,N_7128);
or U7765 (N_7765,N_7339,N_7324);
nor U7766 (N_7766,N_7267,N_7014);
nor U7767 (N_7767,N_7474,N_7357);
xor U7768 (N_7768,N_7016,N_7392);
and U7769 (N_7769,N_7178,N_7378);
nand U7770 (N_7770,N_7443,N_7249);
nand U7771 (N_7771,N_7292,N_7378);
or U7772 (N_7772,N_7010,N_7152);
nor U7773 (N_7773,N_7414,N_7266);
xnor U7774 (N_7774,N_7119,N_7273);
or U7775 (N_7775,N_7005,N_7323);
nor U7776 (N_7776,N_7293,N_7206);
and U7777 (N_7777,N_7469,N_7050);
nand U7778 (N_7778,N_7139,N_7359);
and U7779 (N_7779,N_7094,N_7413);
and U7780 (N_7780,N_7055,N_7044);
nand U7781 (N_7781,N_7061,N_7405);
and U7782 (N_7782,N_7084,N_7207);
nand U7783 (N_7783,N_7193,N_7101);
xnor U7784 (N_7784,N_7081,N_7090);
and U7785 (N_7785,N_7470,N_7033);
nor U7786 (N_7786,N_7488,N_7083);
or U7787 (N_7787,N_7016,N_7265);
nor U7788 (N_7788,N_7197,N_7429);
or U7789 (N_7789,N_7465,N_7447);
or U7790 (N_7790,N_7036,N_7155);
nand U7791 (N_7791,N_7378,N_7453);
and U7792 (N_7792,N_7167,N_7031);
nand U7793 (N_7793,N_7257,N_7175);
or U7794 (N_7794,N_7131,N_7091);
or U7795 (N_7795,N_7428,N_7303);
and U7796 (N_7796,N_7485,N_7263);
nor U7797 (N_7797,N_7072,N_7478);
nand U7798 (N_7798,N_7267,N_7490);
or U7799 (N_7799,N_7285,N_7016);
nand U7800 (N_7800,N_7180,N_7042);
nand U7801 (N_7801,N_7188,N_7428);
xor U7802 (N_7802,N_7018,N_7229);
or U7803 (N_7803,N_7204,N_7453);
xnor U7804 (N_7804,N_7228,N_7435);
xnor U7805 (N_7805,N_7302,N_7199);
nor U7806 (N_7806,N_7074,N_7476);
nor U7807 (N_7807,N_7055,N_7006);
xnor U7808 (N_7808,N_7444,N_7260);
and U7809 (N_7809,N_7290,N_7272);
nand U7810 (N_7810,N_7066,N_7282);
xor U7811 (N_7811,N_7155,N_7204);
or U7812 (N_7812,N_7298,N_7467);
nand U7813 (N_7813,N_7296,N_7255);
nor U7814 (N_7814,N_7079,N_7358);
xor U7815 (N_7815,N_7366,N_7256);
nor U7816 (N_7816,N_7086,N_7289);
nand U7817 (N_7817,N_7175,N_7429);
xor U7818 (N_7818,N_7468,N_7247);
nor U7819 (N_7819,N_7187,N_7361);
and U7820 (N_7820,N_7185,N_7441);
xor U7821 (N_7821,N_7316,N_7209);
and U7822 (N_7822,N_7306,N_7364);
nand U7823 (N_7823,N_7041,N_7308);
or U7824 (N_7824,N_7346,N_7142);
or U7825 (N_7825,N_7325,N_7012);
nand U7826 (N_7826,N_7495,N_7003);
and U7827 (N_7827,N_7479,N_7266);
xnor U7828 (N_7828,N_7438,N_7437);
and U7829 (N_7829,N_7477,N_7428);
xor U7830 (N_7830,N_7102,N_7275);
xnor U7831 (N_7831,N_7065,N_7361);
nor U7832 (N_7832,N_7157,N_7244);
nand U7833 (N_7833,N_7164,N_7468);
and U7834 (N_7834,N_7489,N_7324);
nor U7835 (N_7835,N_7365,N_7274);
nor U7836 (N_7836,N_7108,N_7056);
and U7837 (N_7837,N_7397,N_7355);
nand U7838 (N_7838,N_7045,N_7426);
or U7839 (N_7839,N_7114,N_7192);
nor U7840 (N_7840,N_7201,N_7132);
nand U7841 (N_7841,N_7192,N_7294);
or U7842 (N_7842,N_7401,N_7376);
or U7843 (N_7843,N_7280,N_7154);
xor U7844 (N_7844,N_7236,N_7210);
and U7845 (N_7845,N_7148,N_7075);
xnor U7846 (N_7846,N_7132,N_7377);
and U7847 (N_7847,N_7213,N_7300);
nor U7848 (N_7848,N_7238,N_7102);
and U7849 (N_7849,N_7499,N_7445);
or U7850 (N_7850,N_7254,N_7324);
nor U7851 (N_7851,N_7157,N_7315);
or U7852 (N_7852,N_7197,N_7328);
or U7853 (N_7853,N_7372,N_7452);
and U7854 (N_7854,N_7361,N_7490);
or U7855 (N_7855,N_7435,N_7457);
nand U7856 (N_7856,N_7444,N_7464);
nor U7857 (N_7857,N_7464,N_7314);
or U7858 (N_7858,N_7380,N_7370);
xor U7859 (N_7859,N_7360,N_7434);
or U7860 (N_7860,N_7143,N_7314);
nor U7861 (N_7861,N_7347,N_7361);
and U7862 (N_7862,N_7058,N_7328);
nor U7863 (N_7863,N_7030,N_7163);
nor U7864 (N_7864,N_7069,N_7230);
nor U7865 (N_7865,N_7450,N_7138);
and U7866 (N_7866,N_7248,N_7001);
xor U7867 (N_7867,N_7446,N_7081);
xnor U7868 (N_7868,N_7235,N_7006);
xor U7869 (N_7869,N_7129,N_7008);
or U7870 (N_7870,N_7240,N_7438);
nor U7871 (N_7871,N_7108,N_7373);
nand U7872 (N_7872,N_7429,N_7491);
and U7873 (N_7873,N_7003,N_7223);
xnor U7874 (N_7874,N_7423,N_7221);
and U7875 (N_7875,N_7367,N_7240);
xnor U7876 (N_7876,N_7213,N_7486);
nand U7877 (N_7877,N_7171,N_7011);
nor U7878 (N_7878,N_7499,N_7107);
or U7879 (N_7879,N_7079,N_7060);
and U7880 (N_7880,N_7201,N_7333);
xnor U7881 (N_7881,N_7018,N_7469);
and U7882 (N_7882,N_7188,N_7171);
xor U7883 (N_7883,N_7011,N_7351);
xor U7884 (N_7884,N_7028,N_7389);
and U7885 (N_7885,N_7102,N_7067);
and U7886 (N_7886,N_7029,N_7360);
or U7887 (N_7887,N_7085,N_7025);
and U7888 (N_7888,N_7448,N_7346);
nor U7889 (N_7889,N_7365,N_7301);
nand U7890 (N_7890,N_7291,N_7402);
nand U7891 (N_7891,N_7079,N_7099);
nor U7892 (N_7892,N_7455,N_7209);
or U7893 (N_7893,N_7267,N_7194);
nor U7894 (N_7894,N_7245,N_7255);
or U7895 (N_7895,N_7061,N_7111);
or U7896 (N_7896,N_7125,N_7322);
xnor U7897 (N_7897,N_7474,N_7330);
and U7898 (N_7898,N_7224,N_7470);
or U7899 (N_7899,N_7312,N_7105);
xor U7900 (N_7900,N_7466,N_7014);
xor U7901 (N_7901,N_7081,N_7077);
xor U7902 (N_7902,N_7201,N_7237);
or U7903 (N_7903,N_7446,N_7423);
nand U7904 (N_7904,N_7319,N_7464);
nor U7905 (N_7905,N_7338,N_7465);
nand U7906 (N_7906,N_7341,N_7045);
and U7907 (N_7907,N_7436,N_7049);
xnor U7908 (N_7908,N_7062,N_7486);
nand U7909 (N_7909,N_7064,N_7181);
nor U7910 (N_7910,N_7416,N_7037);
or U7911 (N_7911,N_7179,N_7078);
and U7912 (N_7912,N_7242,N_7486);
nand U7913 (N_7913,N_7046,N_7081);
or U7914 (N_7914,N_7015,N_7382);
or U7915 (N_7915,N_7167,N_7149);
and U7916 (N_7916,N_7351,N_7358);
nor U7917 (N_7917,N_7464,N_7338);
nand U7918 (N_7918,N_7158,N_7405);
nand U7919 (N_7919,N_7444,N_7350);
or U7920 (N_7920,N_7253,N_7373);
xor U7921 (N_7921,N_7170,N_7019);
or U7922 (N_7922,N_7317,N_7139);
and U7923 (N_7923,N_7038,N_7235);
nand U7924 (N_7924,N_7270,N_7236);
nor U7925 (N_7925,N_7483,N_7245);
or U7926 (N_7926,N_7053,N_7405);
nand U7927 (N_7927,N_7135,N_7306);
and U7928 (N_7928,N_7242,N_7347);
nand U7929 (N_7929,N_7270,N_7446);
nor U7930 (N_7930,N_7361,N_7049);
and U7931 (N_7931,N_7035,N_7085);
and U7932 (N_7932,N_7248,N_7160);
nand U7933 (N_7933,N_7292,N_7468);
xnor U7934 (N_7934,N_7242,N_7138);
nor U7935 (N_7935,N_7415,N_7222);
nor U7936 (N_7936,N_7331,N_7037);
or U7937 (N_7937,N_7133,N_7200);
and U7938 (N_7938,N_7191,N_7400);
nand U7939 (N_7939,N_7381,N_7238);
and U7940 (N_7940,N_7475,N_7375);
nand U7941 (N_7941,N_7251,N_7310);
xor U7942 (N_7942,N_7168,N_7179);
and U7943 (N_7943,N_7061,N_7320);
xnor U7944 (N_7944,N_7064,N_7199);
xnor U7945 (N_7945,N_7117,N_7176);
xor U7946 (N_7946,N_7094,N_7130);
xnor U7947 (N_7947,N_7158,N_7187);
and U7948 (N_7948,N_7230,N_7430);
nor U7949 (N_7949,N_7454,N_7184);
and U7950 (N_7950,N_7288,N_7193);
and U7951 (N_7951,N_7085,N_7128);
and U7952 (N_7952,N_7467,N_7009);
or U7953 (N_7953,N_7011,N_7166);
nor U7954 (N_7954,N_7408,N_7102);
xor U7955 (N_7955,N_7145,N_7467);
and U7956 (N_7956,N_7472,N_7105);
nand U7957 (N_7957,N_7464,N_7339);
xor U7958 (N_7958,N_7410,N_7145);
xor U7959 (N_7959,N_7494,N_7482);
and U7960 (N_7960,N_7258,N_7033);
nor U7961 (N_7961,N_7399,N_7291);
or U7962 (N_7962,N_7029,N_7485);
xor U7963 (N_7963,N_7189,N_7176);
nor U7964 (N_7964,N_7312,N_7489);
nor U7965 (N_7965,N_7406,N_7016);
nand U7966 (N_7966,N_7470,N_7430);
nand U7967 (N_7967,N_7277,N_7046);
or U7968 (N_7968,N_7201,N_7124);
xor U7969 (N_7969,N_7334,N_7181);
and U7970 (N_7970,N_7254,N_7341);
nand U7971 (N_7971,N_7069,N_7216);
and U7972 (N_7972,N_7246,N_7278);
nor U7973 (N_7973,N_7194,N_7484);
nor U7974 (N_7974,N_7243,N_7020);
xnor U7975 (N_7975,N_7157,N_7335);
or U7976 (N_7976,N_7312,N_7410);
nand U7977 (N_7977,N_7363,N_7220);
xnor U7978 (N_7978,N_7415,N_7178);
or U7979 (N_7979,N_7010,N_7413);
and U7980 (N_7980,N_7015,N_7029);
xnor U7981 (N_7981,N_7014,N_7332);
or U7982 (N_7982,N_7468,N_7238);
and U7983 (N_7983,N_7196,N_7101);
nand U7984 (N_7984,N_7307,N_7230);
xor U7985 (N_7985,N_7224,N_7043);
nand U7986 (N_7986,N_7495,N_7312);
nand U7987 (N_7987,N_7066,N_7202);
xnor U7988 (N_7988,N_7213,N_7471);
and U7989 (N_7989,N_7215,N_7398);
and U7990 (N_7990,N_7434,N_7117);
and U7991 (N_7991,N_7049,N_7183);
nand U7992 (N_7992,N_7374,N_7133);
or U7993 (N_7993,N_7198,N_7481);
and U7994 (N_7994,N_7112,N_7010);
or U7995 (N_7995,N_7326,N_7065);
nand U7996 (N_7996,N_7042,N_7222);
xnor U7997 (N_7997,N_7223,N_7125);
and U7998 (N_7998,N_7025,N_7046);
xnor U7999 (N_7999,N_7455,N_7423);
nand U8000 (N_8000,N_7932,N_7959);
and U8001 (N_8001,N_7737,N_7874);
and U8002 (N_8002,N_7502,N_7715);
nand U8003 (N_8003,N_7859,N_7803);
nor U8004 (N_8004,N_7678,N_7636);
nor U8005 (N_8005,N_7721,N_7856);
or U8006 (N_8006,N_7758,N_7894);
xnor U8007 (N_8007,N_7882,N_7848);
or U8008 (N_8008,N_7569,N_7509);
and U8009 (N_8009,N_7812,N_7699);
xor U8010 (N_8010,N_7974,N_7897);
and U8011 (N_8011,N_7814,N_7806);
xor U8012 (N_8012,N_7809,N_7765);
nor U8013 (N_8013,N_7731,N_7710);
and U8014 (N_8014,N_7876,N_7658);
xnor U8015 (N_8015,N_7837,N_7650);
nor U8016 (N_8016,N_7981,N_7573);
nor U8017 (N_8017,N_7786,N_7682);
nor U8018 (N_8018,N_7749,N_7960);
and U8019 (N_8019,N_7780,N_7553);
or U8020 (N_8020,N_7598,N_7671);
nor U8021 (N_8021,N_7823,N_7936);
or U8022 (N_8022,N_7541,N_7578);
and U8023 (N_8023,N_7795,N_7612);
and U8024 (N_8024,N_7742,N_7924);
nor U8025 (N_8025,N_7632,N_7910);
and U8026 (N_8026,N_7602,N_7638);
nand U8027 (N_8027,N_7588,N_7555);
nand U8028 (N_8028,N_7750,N_7889);
nand U8029 (N_8029,N_7655,N_7937);
nand U8030 (N_8030,N_7911,N_7623);
or U8031 (N_8031,N_7935,N_7739);
and U8032 (N_8032,N_7993,N_7982);
nor U8033 (N_8033,N_7881,N_7593);
nand U8034 (N_8034,N_7620,N_7672);
nand U8035 (N_8035,N_7648,N_7515);
nor U8036 (N_8036,N_7627,N_7985);
nand U8037 (N_8037,N_7722,N_7679);
or U8038 (N_8038,N_7585,N_7857);
and U8039 (N_8039,N_7862,N_7783);
nand U8040 (N_8040,N_7766,N_7868);
nor U8041 (N_8041,N_7759,N_7528);
and U8042 (N_8042,N_7531,N_7666);
nor U8043 (N_8043,N_7551,N_7549);
xor U8044 (N_8044,N_7810,N_7797);
nand U8045 (N_8045,N_7727,N_7827);
and U8046 (N_8046,N_7639,N_7805);
xnor U8047 (N_8047,N_7907,N_7940);
nor U8048 (N_8048,N_7559,N_7660);
and U8049 (N_8049,N_7538,N_7953);
nor U8050 (N_8050,N_7927,N_7608);
or U8051 (N_8051,N_7664,N_7979);
xor U8052 (N_8052,N_7522,N_7928);
or U8053 (N_8053,N_7550,N_7842);
nor U8054 (N_8054,N_7646,N_7500);
and U8055 (N_8055,N_7929,N_7586);
nand U8056 (N_8056,N_7668,N_7505);
nand U8057 (N_8057,N_7649,N_7820);
nor U8058 (N_8058,N_7767,N_7886);
and U8059 (N_8059,N_7733,N_7734);
and U8060 (N_8060,N_7700,N_7616);
nand U8061 (N_8061,N_7657,N_7869);
nor U8062 (N_8062,N_7770,N_7663);
or U8063 (N_8063,N_7594,N_7922);
nand U8064 (N_8064,N_7796,N_7808);
xnor U8065 (N_8065,N_7730,N_7961);
nor U8066 (N_8066,N_7512,N_7514);
xor U8067 (N_8067,N_7879,N_7614);
or U8068 (N_8068,N_7818,N_7508);
nand U8069 (N_8069,N_7893,N_7754);
xnor U8070 (N_8070,N_7871,N_7792);
or U8071 (N_8071,N_7822,N_7850);
xnor U8072 (N_8072,N_7587,N_7618);
nor U8073 (N_8073,N_7776,N_7839);
nand U8074 (N_8074,N_7788,N_7983);
or U8075 (N_8075,N_7851,N_7525);
nand U8076 (N_8076,N_7507,N_7607);
and U8077 (N_8077,N_7619,N_7916);
and U8078 (N_8078,N_7622,N_7757);
nand U8079 (N_8079,N_7908,N_7813);
nand U8080 (N_8080,N_7943,N_7728);
nor U8081 (N_8081,N_7833,N_7933);
or U8082 (N_8082,N_7977,N_7630);
nand U8083 (N_8083,N_7954,N_7694);
nor U8084 (N_8084,N_7527,N_7652);
nand U8085 (N_8085,N_7909,N_7704);
nor U8086 (N_8086,N_7884,N_7661);
and U8087 (N_8087,N_7952,N_7878);
xor U8088 (N_8088,N_7540,N_7942);
xor U8089 (N_8089,N_7624,N_7853);
nor U8090 (N_8090,N_7637,N_7504);
xnor U8091 (N_8091,N_7877,N_7501);
nor U8092 (N_8092,N_7873,N_7854);
nor U8093 (N_8093,N_7867,N_7831);
or U8094 (N_8094,N_7891,N_7965);
and U8095 (N_8095,N_7536,N_7662);
nand U8096 (N_8096,N_7740,N_7510);
or U8097 (N_8097,N_7844,N_7571);
nand U8098 (N_8098,N_7816,N_7978);
xor U8099 (N_8099,N_7611,N_7811);
and U8100 (N_8100,N_7926,N_7968);
and U8101 (N_8101,N_7885,N_7702);
or U8102 (N_8102,N_7775,N_7579);
nand U8103 (N_8103,N_7539,N_7519);
xor U8104 (N_8104,N_7785,N_7976);
nor U8105 (N_8105,N_7617,N_7986);
nand U8106 (N_8106,N_7870,N_7847);
and U8107 (N_8107,N_7606,N_7980);
and U8108 (N_8108,N_7930,N_7774);
xnor U8109 (N_8109,N_7784,N_7950);
nor U8110 (N_8110,N_7777,N_7596);
or U8111 (N_8111,N_7526,N_7503);
nor U8112 (N_8112,N_7898,N_7688);
xor U8113 (N_8113,N_7790,N_7970);
xor U8114 (N_8114,N_7957,N_7745);
and U8115 (N_8115,N_7567,N_7905);
or U8116 (N_8116,N_7934,N_7609);
and U8117 (N_8117,N_7902,N_7691);
nor U8118 (N_8118,N_7529,N_7801);
xnor U8119 (N_8119,N_7676,N_7755);
nand U8120 (N_8120,N_7925,N_7782);
xnor U8121 (N_8121,N_7904,N_7689);
xor U8122 (N_8122,N_7725,N_7709);
or U8123 (N_8123,N_7963,N_7582);
or U8124 (N_8124,N_7975,N_7656);
or U8125 (N_8125,N_7724,N_7667);
or U8126 (N_8126,N_7992,N_7561);
nor U8127 (N_8127,N_7523,N_7761);
xor U8128 (N_8128,N_7872,N_7938);
and U8129 (N_8129,N_7613,N_7695);
or U8130 (N_8130,N_7703,N_7684);
or U8131 (N_8131,N_7610,N_7717);
nor U8132 (N_8132,N_7866,N_7799);
xor U8133 (N_8133,N_7517,N_7732);
or U8134 (N_8134,N_7651,N_7696);
xor U8135 (N_8135,N_7955,N_7535);
or U8136 (N_8136,N_7800,N_7888);
and U8137 (N_8137,N_7990,N_7971);
and U8138 (N_8138,N_7941,N_7912);
or U8139 (N_8139,N_7572,N_7534);
or U8140 (N_8140,N_7537,N_7764);
nand U8141 (N_8141,N_7923,N_7746);
nor U8142 (N_8142,N_7726,N_7697);
nor U8143 (N_8143,N_7506,N_7883);
or U8144 (N_8144,N_7706,N_7583);
xor U8145 (N_8145,N_7565,N_7643);
or U8146 (N_8146,N_7964,N_7631);
xor U8147 (N_8147,N_7736,N_7798);
nand U8148 (N_8148,N_7988,N_7892);
nor U8149 (N_8149,N_7675,N_7584);
and U8150 (N_8150,N_7680,N_7832);
nand U8151 (N_8151,N_7778,N_7563);
xor U8152 (N_8152,N_7865,N_7969);
nor U8153 (N_8153,N_7793,N_7747);
or U8154 (N_8154,N_7591,N_7544);
nand U8155 (N_8155,N_7719,N_7570);
or U8156 (N_8156,N_7875,N_7580);
nand U8157 (N_8157,N_7962,N_7713);
nand U8158 (N_8158,N_7558,N_7511);
xnor U8159 (N_8159,N_7677,N_7768);
or U8160 (N_8160,N_7673,N_7966);
nand U8161 (N_8161,N_7599,N_7521);
nor U8162 (N_8162,N_7674,N_7906);
xor U8163 (N_8163,N_7789,N_7642);
or U8164 (N_8164,N_7633,N_7920);
or U8165 (N_8165,N_7686,N_7903);
or U8166 (N_8166,N_7698,N_7751);
nor U8167 (N_8167,N_7654,N_7524);
nand U8168 (N_8168,N_7665,N_7855);
and U8169 (N_8169,N_7575,N_7995);
xor U8170 (N_8170,N_7989,N_7690);
nor U8171 (N_8171,N_7645,N_7560);
nand U8172 (N_8172,N_7753,N_7804);
or U8173 (N_8173,N_7948,N_7997);
or U8174 (N_8174,N_7513,N_7821);
and U8175 (N_8175,N_7773,N_7647);
nor U8176 (N_8176,N_7826,N_7817);
or U8177 (N_8177,N_7849,N_7946);
nand U8178 (N_8178,N_7914,N_7752);
nand U8179 (N_8179,N_7951,N_7807);
nand U8180 (N_8180,N_7824,N_7835);
nor U8181 (N_8181,N_7685,N_7779);
nor U8182 (N_8182,N_7917,N_7836);
or U8183 (N_8183,N_7973,N_7748);
xor U8184 (N_8184,N_7998,N_7603);
xnor U8185 (N_8185,N_7828,N_7772);
and U8186 (N_8186,N_7597,N_7653);
or U8187 (N_8187,N_7687,N_7987);
nor U8188 (N_8188,N_7520,N_7564);
nor U8189 (N_8189,N_7838,N_7843);
nand U8190 (N_8190,N_7716,N_7845);
nand U8191 (N_8191,N_7815,N_7589);
and U8192 (N_8192,N_7944,N_7945);
or U8193 (N_8193,N_7556,N_7621);
or U8194 (N_8194,N_7840,N_7547);
or U8195 (N_8195,N_7825,N_7533);
xnor U8196 (N_8196,N_7738,N_7545);
nor U8197 (N_8197,N_7635,N_7967);
xnor U8198 (N_8198,N_7899,N_7605);
nor U8199 (N_8199,N_7600,N_7781);
or U8200 (N_8200,N_7919,N_7999);
xor U8201 (N_8201,N_7791,N_7723);
and U8202 (N_8202,N_7756,N_7846);
nand U8203 (N_8203,N_7984,N_7890);
and U8204 (N_8204,N_7729,N_7595);
or U8205 (N_8205,N_7802,N_7601);
xor U8206 (N_8206,N_7711,N_7915);
and U8207 (N_8207,N_7590,N_7626);
nor U8208 (N_8208,N_7735,N_7532);
nand U8209 (N_8209,N_7896,N_7895);
nand U8210 (N_8210,N_7939,N_7577);
and U8211 (N_8211,N_7829,N_7834);
or U8212 (N_8212,N_7760,N_7763);
or U8213 (N_8213,N_7628,N_7592);
and U8214 (N_8214,N_7629,N_7743);
and U8215 (N_8215,N_7861,N_7681);
or U8216 (N_8216,N_7542,N_7887);
and U8217 (N_8217,N_7769,N_7819);
or U8218 (N_8218,N_7956,N_7741);
xor U8219 (N_8219,N_7554,N_7996);
or U8220 (N_8220,N_7787,N_7701);
nand U8221 (N_8221,N_7659,N_7880);
or U8222 (N_8222,N_7858,N_7994);
nor U8223 (N_8223,N_7708,N_7864);
or U8224 (N_8224,N_7518,N_7991);
and U8225 (N_8225,N_7705,N_7604);
and U8226 (N_8226,N_7530,N_7640);
and U8227 (N_8227,N_7718,N_7901);
nand U8228 (N_8228,N_7949,N_7860);
and U8229 (N_8229,N_7720,N_7693);
and U8230 (N_8230,N_7947,N_7615);
xnor U8231 (N_8231,N_7744,N_7921);
or U8232 (N_8232,N_7712,N_7771);
or U8233 (N_8233,N_7576,N_7913);
and U8234 (N_8234,N_7670,N_7574);
nor U8235 (N_8235,N_7707,N_7566);
xor U8236 (N_8236,N_7634,N_7683);
nand U8237 (N_8237,N_7543,N_7863);
and U8238 (N_8238,N_7762,N_7562);
nor U8239 (N_8239,N_7714,N_7557);
and U8240 (N_8240,N_7900,N_7852);
xor U8241 (N_8241,N_7669,N_7625);
nand U8242 (N_8242,N_7641,N_7830);
nor U8243 (N_8243,N_7931,N_7552);
or U8244 (N_8244,N_7958,N_7644);
nor U8245 (N_8245,N_7581,N_7548);
or U8246 (N_8246,N_7516,N_7794);
and U8247 (N_8247,N_7692,N_7972);
xor U8248 (N_8248,N_7546,N_7841);
nand U8249 (N_8249,N_7568,N_7918);
nor U8250 (N_8250,N_7910,N_7741);
nor U8251 (N_8251,N_7653,N_7853);
and U8252 (N_8252,N_7521,N_7504);
and U8253 (N_8253,N_7838,N_7959);
or U8254 (N_8254,N_7601,N_7720);
nand U8255 (N_8255,N_7855,N_7789);
nand U8256 (N_8256,N_7594,N_7544);
nand U8257 (N_8257,N_7758,N_7681);
nor U8258 (N_8258,N_7603,N_7842);
nor U8259 (N_8259,N_7996,N_7552);
xnor U8260 (N_8260,N_7934,N_7554);
nand U8261 (N_8261,N_7552,N_7593);
nor U8262 (N_8262,N_7789,N_7660);
or U8263 (N_8263,N_7669,N_7742);
or U8264 (N_8264,N_7721,N_7607);
or U8265 (N_8265,N_7937,N_7656);
nor U8266 (N_8266,N_7593,N_7592);
nand U8267 (N_8267,N_7518,N_7531);
and U8268 (N_8268,N_7862,N_7527);
nor U8269 (N_8269,N_7879,N_7898);
and U8270 (N_8270,N_7726,N_7545);
and U8271 (N_8271,N_7544,N_7632);
nor U8272 (N_8272,N_7512,N_7968);
and U8273 (N_8273,N_7818,N_7787);
or U8274 (N_8274,N_7648,N_7641);
xnor U8275 (N_8275,N_7793,N_7507);
xor U8276 (N_8276,N_7744,N_7708);
and U8277 (N_8277,N_7921,N_7853);
nand U8278 (N_8278,N_7555,N_7605);
and U8279 (N_8279,N_7712,N_7673);
nor U8280 (N_8280,N_7517,N_7698);
and U8281 (N_8281,N_7678,N_7507);
and U8282 (N_8282,N_7806,N_7555);
and U8283 (N_8283,N_7874,N_7788);
nor U8284 (N_8284,N_7995,N_7748);
and U8285 (N_8285,N_7911,N_7503);
nor U8286 (N_8286,N_7633,N_7754);
or U8287 (N_8287,N_7916,N_7966);
nand U8288 (N_8288,N_7816,N_7880);
nand U8289 (N_8289,N_7611,N_7634);
and U8290 (N_8290,N_7952,N_7963);
nor U8291 (N_8291,N_7633,N_7500);
nand U8292 (N_8292,N_7811,N_7936);
xor U8293 (N_8293,N_7550,N_7889);
nand U8294 (N_8294,N_7531,N_7613);
nor U8295 (N_8295,N_7792,N_7902);
xor U8296 (N_8296,N_7654,N_7547);
nor U8297 (N_8297,N_7870,N_7875);
or U8298 (N_8298,N_7943,N_7555);
nor U8299 (N_8299,N_7704,N_7873);
nor U8300 (N_8300,N_7590,N_7828);
and U8301 (N_8301,N_7989,N_7601);
xor U8302 (N_8302,N_7819,N_7874);
and U8303 (N_8303,N_7727,N_7728);
nand U8304 (N_8304,N_7690,N_7706);
xnor U8305 (N_8305,N_7780,N_7760);
or U8306 (N_8306,N_7825,N_7731);
nor U8307 (N_8307,N_7748,N_7822);
and U8308 (N_8308,N_7874,N_7718);
nor U8309 (N_8309,N_7745,N_7972);
nor U8310 (N_8310,N_7627,N_7774);
nand U8311 (N_8311,N_7835,N_7851);
xnor U8312 (N_8312,N_7536,N_7647);
nand U8313 (N_8313,N_7714,N_7782);
nand U8314 (N_8314,N_7983,N_7645);
nor U8315 (N_8315,N_7853,N_7737);
nand U8316 (N_8316,N_7983,N_7690);
xnor U8317 (N_8317,N_7647,N_7791);
or U8318 (N_8318,N_7536,N_7703);
nand U8319 (N_8319,N_7931,N_7967);
nand U8320 (N_8320,N_7533,N_7652);
nand U8321 (N_8321,N_7873,N_7723);
or U8322 (N_8322,N_7518,N_7928);
nand U8323 (N_8323,N_7685,N_7843);
xor U8324 (N_8324,N_7714,N_7873);
and U8325 (N_8325,N_7540,N_7607);
nand U8326 (N_8326,N_7600,N_7719);
nand U8327 (N_8327,N_7858,N_7792);
nand U8328 (N_8328,N_7569,N_7694);
nor U8329 (N_8329,N_7602,N_7979);
nor U8330 (N_8330,N_7662,N_7799);
and U8331 (N_8331,N_7794,N_7628);
nor U8332 (N_8332,N_7578,N_7941);
and U8333 (N_8333,N_7866,N_7530);
xor U8334 (N_8334,N_7753,N_7628);
nand U8335 (N_8335,N_7852,N_7779);
xor U8336 (N_8336,N_7770,N_7582);
xor U8337 (N_8337,N_7618,N_7973);
nor U8338 (N_8338,N_7991,N_7734);
xor U8339 (N_8339,N_7964,N_7759);
xor U8340 (N_8340,N_7632,N_7651);
nor U8341 (N_8341,N_7727,N_7833);
nor U8342 (N_8342,N_7885,N_7512);
xor U8343 (N_8343,N_7585,N_7510);
or U8344 (N_8344,N_7848,N_7729);
nor U8345 (N_8345,N_7740,N_7984);
and U8346 (N_8346,N_7589,N_7673);
xnor U8347 (N_8347,N_7934,N_7930);
nand U8348 (N_8348,N_7874,N_7591);
nand U8349 (N_8349,N_7870,N_7876);
or U8350 (N_8350,N_7810,N_7920);
nor U8351 (N_8351,N_7690,N_7707);
or U8352 (N_8352,N_7928,N_7947);
nand U8353 (N_8353,N_7631,N_7744);
or U8354 (N_8354,N_7948,N_7640);
and U8355 (N_8355,N_7510,N_7929);
and U8356 (N_8356,N_7862,N_7507);
and U8357 (N_8357,N_7747,N_7805);
and U8358 (N_8358,N_7516,N_7661);
and U8359 (N_8359,N_7941,N_7750);
or U8360 (N_8360,N_7980,N_7880);
nand U8361 (N_8361,N_7628,N_7969);
nand U8362 (N_8362,N_7604,N_7811);
nand U8363 (N_8363,N_7815,N_7528);
nor U8364 (N_8364,N_7816,N_7615);
or U8365 (N_8365,N_7651,N_7745);
xnor U8366 (N_8366,N_7587,N_7563);
xnor U8367 (N_8367,N_7905,N_7645);
nor U8368 (N_8368,N_7934,N_7867);
or U8369 (N_8369,N_7956,N_7976);
or U8370 (N_8370,N_7825,N_7795);
xnor U8371 (N_8371,N_7870,N_7644);
nand U8372 (N_8372,N_7602,N_7863);
xor U8373 (N_8373,N_7790,N_7807);
xnor U8374 (N_8374,N_7547,N_7664);
or U8375 (N_8375,N_7939,N_7575);
or U8376 (N_8376,N_7676,N_7669);
and U8377 (N_8377,N_7593,N_7549);
and U8378 (N_8378,N_7808,N_7870);
and U8379 (N_8379,N_7784,N_7724);
xor U8380 (N_8380,N_7845,N_7629);
or U8381 (N_8381,N_7692,N_7870);
nand U8382 (N_8382,N_7980,N_7957);
nor U8383 (N_8383,N_7960,N_7932);
xnor U8384 (N_8384,N_7741,N_7679);
and U8385 (N_8385,N_7673,N_7633);
nor U8386 (N_8386,N_7866,N_7950);
nand U8387 (N_8387,N_7789,N_7551);
and U8388 (N_8388,N_7797,N_7973);
and U8389 (N_8389,N_7963,N_7989);
and U8390 (N_8390,N_7648,N_7815);
or U8391 (N_8391,N_7567,N_7685);
and U8392 (N_8392,N_7865,N_7555);
or U8393 (N_8393,N_7955,N_7574);
or U8394 (N_8394,N_7674,N_7737);
and U8395 (N_8395,N_7877,N_7711);
or U8396 (N_8396,N_7906,N_7854);
and U8397 (N_8397,N_7892,N_7557);
or U8398 (N_8398,N_7928,N_7917);
and U8399 (N_8399,N_7749,N_7837);
nand U8400 (N_8400,N_7964,N_7772);
nand U8401 (N_8401,N_7574,N_7993);
or U8402 (N_8402,N_7969,N_7710);
nor U8403 (N_8403,N_7882,N_7826);
or U8404 (N_8404,N_7891,N_7676);
nand U8405 (N_8405,N_7528,N_7817);
and U8406 (N_8406,N_7869,N_7640);
and U8407 (N_8407,N_7750,N_7960);
xnor U8408 (N_8408,N_7536,N_7627);
and U8409 (N_8409,N_7715,N_7619);
nor U8410 (N_8410,N_7942,N_7957);
nor U8411 (N_8411,N_7540,N_7686);
xnor U8412 (N_8412,N_7558,N_7728);
nand U8413 (N_8413,N_7839,N_7694);
nor U8414 (N_8414,N_7555,N_7743);
and U8415 (N_8415,N_7798,N_7784);
or U8416 (N_8416,N_7832,N_7578);
or U8417 (N_8417,N_7591,N_7590);
and U8418 (N_8418,N_7692,N_7596);
nor U8419 (N_8419,N_7750,N_7886);
xnor U8420 (N_8420,N_7903,N_7649);
or U8421 (N_8421,N_7607,N_7712);
nand U8422 (N_8422,N_7828,N_7953);
nor U8423 (N_8423,N_7840,N_7515);
xnor U8424 (N_8424,N_7720,N_7689);
nor U8425 (N_8425,N_7943,N_7873);
and U8426 (N_8426,N_7690,N_7926);
or U8427 (N_8427,N_7824,N_7779);
xor U8428 (N_8428,N_7865,N_7938);
nor U8429 (N_8429,N_7916,N_7882);
nand U8430 (N_8430,N_7758,N_7957);
xnor U8431 (N_8431,N_7658,N_7500);
xor U8432 (N_8432,N_7657,N_7641);
nand U8433 (N_8433,N_7939,N_7503);
nand U8434 (N_8434,N_7657,N_7748);
xor U8435 (N_8435,N_7593,N_7697);
xnor U8436 (N_8436,N_7962,N_7670);
xnor U8437 (N_8437,N_7992,N_7650);
xor U8438 (N_8438,N_7708,N_7890);
xnor U8439 (N_8439,N_7927,N_7513);
and U8440 (N_8440,N_7656,N_7856);
or U8441 (N_8441,N_7675,N_7873);
nor U8442 (N_8442,N_7929,N_7534);
nor U8443 (N_8443,N_7959,N_7736);
or U8444 (N_8444,N_7935,N_7918);
nand U8445 (N_8445,N_7764,N_7977);
or U8446 (N_8446,N_7581,N_7557);
nor U8447 (N_8447,N_7570,N_7766);
and U8448 (N_8448,N_7751,N_7671);
nand U8449 (N_8449,N_7816,N_7665);
nor U8450 (N_8450,N_7868,N_7995);
and U8451 (N_8451,N_7812,N_7899);
xnor U8452 (N_8452,N_7908,N_7597);
and U8453 (N_8453,N_7749,N_7833);
nand U8454 (N_8454,N_7855,N_7862);
or U8455 (N_8455,N_7852,N_7646);
nand U8456 (N_8456,N_7782,N_7766);
xor U8457 (N_8457,N_7716,N_7780);
or U8458 (N_8458,N_7971,N_7873);
or U8459 (N_8459,N_7820,N_7648);
and U8460 (N_8460,N_7709,N_7949);
and U8461 (N_8461,N_7675,N_7549);
or U8462 (N_8462,N_7778,N_7541);
and U8463 (N_8463,N_7806,N_7564);
nor U8464 (N_8464,N_7980,N_7691);
nor U8465 (N_8465,N_7920,N_7908);
or U8466 (N_8466,N_7668,N_7683);
and U8467 (N_8467,N_7652,N_7517);
xor U8468 (N_8468,N_7853,N_7710);
or U8469 (N_8469,N_7722,N_7936);
or U8470 (N_8470,N_7679,N_7684);
and U8471 (N_8471,N_7990,N_7750);
nor U8472 (N_8472,N_7850,N_7564);
nor U8473 (N_8473,N_7998,N_7978);
or U8474 (N_8474,N_7656,N_7744);
nor U8475 (N_8475,N_7867,N_7642);
nand U8476 (N_8476,N_7766,N_7503);
nor U8477 (N_8477,N_7634,N_7597);
xor U8478 (N_8478,N_7941,N_7740);
or U8479 (N_8479,N_7897,N_7841);
xor U8480 (N_8480,N_7884,N_7507);
xor U8481 (N_8481,N_7893,N_7638);
or U8482 (N_8482,N_7865,N_7864);
xnor U8483 (N_8483,N_7840,N_7894);
xor U8484 (N_8484,N_7867,N_7721);
xnor U8485 (N_8485,N_7684,N_7624);
nor U8486 (N_8486,N_7615,N_7951);
xnor U8487 (N_8487,N_7889,N_7866);
and U8488 (N_8488,N_7756,N_7568);
and U8489 (N_8489,N_7600,N_7605);
nor U8490 (N_8490,N_7855,N_7835);
nor U8491 (N_8491,N_7624,N_7565);
xnor U8492 (N_8492,N_7903,N_7729);
and U8493 (N_8493,N_7538,N_7984);
xnor U8494 (N_8494,N_7969,N_7740);
xor U8495 (N_8495,N_7557,N_7970);
or U8496 (N_8496,N_7959,N_7772);
and U8497 (N_8497,N_7782,N_7778);
nor U8498 (N_8498,N_7967,N_7557);
xnor U8499 (N_8499,N_7870,N_7678);
or U8500 (N_8500,N_8456,N_8103);
nor U8501 (N_8501,N_8297,N_8231);
nand U8502 (N_8502,N_8492,N_8322);
xor U8503 (N_8503,N_8155,N_8288);
nor U8504 (N_8504,N_8120,N_8212);
xor U8505 (N_8505,N_8023,N_8036);
nor U8506 (N_8506,N_8240,N_8066);
xor U8507 (N_8507,N_8087,N_8356);
or U8508 (N_8508,N_8257,N_8001);
nor U8509 (N_8509,N_8056,N_8355);
or U8510 (N_8510,N_8168,N_8274);
nor U8511 (N_8511,N_8141,N_8494);
nor U8512 (N_8512,N_8265,N_8013);
nand U8513 (N_8513,N_8064,N_8409);
nand U8514 (N_8514,N_8382,N_8326);
and U8515 (N_8515,N_8394,N_8243);
xor U8516 (N_8516,N_8200,N_8445);
xor U8517 (N_8517,N_8174,N_8453);
and U8518 (N_8518,N_8289,N_8019);
or U8519 (N_8519,N_8049,N_8061);
nor U8520 (N_8520,N_8415,N_8338);
or U8521 (N_8521,N_8258,N_8006);
nor U8522 (N_8522,N_8408,N_8316);
and U8523 (N_8523,N_8248,N_8135);
nand U8524 (N_8524,N_8365,N_8410);
and U8525 (N_8525,N_8438,N_8245);
or U8526 (N_8526,N_8011,N_8283);
xnor U8527 (N_8527,N_8392,N_8101);
or U8528 (N_8528,N_8478,N_8312);
or U8529 (N_8529,N_8221,N_8208);
or U8530 (N_8530,N_8439,N_8089);
and U8531 (N_8531,N_8018,N_8232);
and U8532 (N_8532,N_8241,N_8154);
nor U8533 (N_8533,N_8127,N_8102);
or U8534 (N_8534,N_8260,N_8470);
and U8535 (N_8535,N_8096,N_8166);
xnor U8536 (N_8536,N_8170,N_8107);
nand U8537 (N_8537,N_8163,N_8042);
or U8538 (N_8538,N_8205,N_8063);
and U8539 (N_8539,N_8395,N_8071);
xor U8540 (N_8540,N_8175,N_8372);
nor U8541 (N_8541,N_8278,N_8449);
or U8542 (N_8542,N_8165,N_8310);
and U8543 (N_8543,N_8458,N_8325);
xnor U8544 (N_8544,N_8369,N_8189);
nor U8545 (N_8545,N_8239,N_8086);
nand U8546 (N_8546,N_8176,N_8040);
xnor U8547 (N_8547,N_8424,N_8124);
or U8548 (N_8548,N_8062,N_8311);
or U8549 (N_8549,N_8129,N_8003);
nor U8550 (N_8550,N_8303,N_8268);
or U8551 (N_8551,N_8055,N_8448);
nor U8552 (N_8552,N_8052,N_8426);
nor U8553 (N_8553,N_8111,N_8463);
nand U8554 (N_8554,N_8179,N_8192);
or U8555 (N_8555,N_8053,N_8216);
or U8556 (N_8556,N_8477,N_8084);
nand U8557 (N_8557,N_8405,N_8466);
and U8558 (N_8558,N_8475,N_8304);
and U8559 (N_8559,N_8389,N_8264);
and U8560 (N_8560,N_8157,N_8381);
xnor U8561 (N_8561,N_8217,N_8237);
nor U8562 (N_8562,N_8495,N_8110);
xor U8563 (N_8563,N_8060,N_8029);
nor U8564 (N_8564,N_8413,N_8139);
xnor U8565 (N_8565,N_8423,N_8306);
and U8566 (N_8566,N_8436,N_8173);
and U8567 (N_8567,N_8204,N_8222);
nor U8568 (N_8568,N_8353,N_8030);
or U8569 (N_8569,N_8285,N_8065);
nand U8570 (N_8570,N_8333,N_8076);
nor U8571 (N_8571,N_8223,N_8476);
and U8572 (N_8572,N_8359,N_8004);
xor U8573 (N_8573,N_8295,N_8272);
nor U8574 (N_8574,N_8201,N_8469);
nor U8575 (N_8575,N_8330,N_8235);
nand U8576 (N_8576,N_8000,N_8197);
xor U8577 (N_8577,N_8002,N_8227);
and U8578 (N_8578,N_8115,N_8486);
nand U8579 (N_8579,N_8400,N_8454);
nand U8580 (N_8580,N_8387,N_8341);
nand U8581 (N_8581,N_8432,N_8468);
or U8582 (N_8582,N_8420,N_8024);
xor U8583 (N_8583,N_8350,N_8499);
xor U8584 (N_8584,N_8207,N_8090);
or U8585 (N_8585,N_8347,N_8109);
xor U8586 (N_8586,N_8277,N_8186);
nand U8587 (N_8587,N_8412,N_8203);
nand U8588 (N_8588,N_8151,N_8038);
xor U8589 (N_8589,N_8298,N_8016);
or U8590 (N_8590,N_8380,N_8128);
or U8591 (N_8591,N_8397,N_8095);
nor U8592 (N_8592,N_8122,N_8370);
or U8593 (N_8593,N_8421,N_8206);
and U8594 (N_8594,N_8150,N_8323);
or U8595 (N_8595,N_8242,N_8336);
and U8596 (N_8596,N_8075,N_8443);
nand U8597 (N_8597,N_8352,N_8185);
nand U8598 (N_8598,N_8136,N_8044);
or U8599 (N_8599,N_8181,N_8167);
and U8600 (N_8600,N_8318,N_8007);
and U8601 (N_8601,N_8043,N_8249);
xor U8602 (N_8602,N_8244,N_8028);
xnor U8603 (N_8603,N_8309,N_8403);
and U8604 (N_8604,N_8045,N_8373);
nor U8605 (N_8605,N_8198,N_8296);
nand U8606 (N_8606,N_8319,N_8273);
xnor U8607 (N_8607,N_8488,N_8396);
nand U8608 (N_8608,N_8282,N_8270);
nor U8609 (N_8609,N_8329,N_8366);
xor U8610 (N_8610,N_8098,N_8349);
or U8611 (N_8611,N_8020,N_8427);
nor U8612 (N_8612,N_8374,N_8346);
nand U8613 (N_8613,N_8378,N_8262);
and U8614 (N_8614,N_8450,N_8280);
and U8615 (N_8615,N_8251,N_8057);
and U8616 (N_8616,N_8269,N_8481);
or U8617 (N_8617,N_8491,N_8379);
or U8618 (N_8618,N_8498,N_8188);
xor U8619 (N_8619,N_8073,N_8255);
xor U8620 (N_8620,N_8119,N_8497);
nor U8621 (N_8621,N_8471,N_8401);
nand U8622 (N_8622,N_8482,N_8292);
nor U8623 (N_8623,N_8105,N_8085);
or U8624 (N_8624,N_8091,N_8404);
or U8625 (N_8625,N_8375,N_8088);
nand U8626 (N_8626,N_8254,N_8158);
xor U8627 (N_8627,N_8331,N_8035);
and U8628 (N_8628,N_8286,N_8080);
nand U8629 (N_8629,N_8225,N_8148);
xor U8630 (N_8630,N_8348,N_8146);
nor U8631 (N_8631,N_8140,N_8210);
nand U8632 (N_8632,N_8496,N_8314);
and U8633 (N_8633,N_8428,N_8339);
and U8634 (N_8634,N_8108,N_8183);
nor U8635 (N_8635,N_8259,N_8407);
or U8636 (N_8636,N_8388,N_8164);
nor U8637 (N_8637,N_8229,N_8133);
nor U8638 (N_8638,N_8162,N_8191);
xor U8639 (N_8639,N_8376,N_8039);
xnor U8640 (N_8640,N_8074,N_8440);
and U8641 (N_8641,N_8434,N_8238);
nand U8642 (N_8642,N_8072,N_8113);
and U8643 (N_8643,N_8473,N_8358);
xnor U8644 (N_8644,N_8145,N_8290);
or U8645 (N_8645,N_8327,N_8187);
and U8646 (N_8646,N_8414,N_8017);
nand U8647 (N_8647,N_8461,N_8067);
nor U8648 (N_8648,N_8256,N_8429);
nor U8649 (N_8649,N_8435,N_8377);
xor U8650 (N_8650,N_8058,N_8250);
or U8651 (N_8651,N_8411,N_8361);
nand U8652 (N_8652,N_8281,N_8209);
xnor U8653 (N_8653,N_8487,N_8144);
nand U8654 (N_8654,N_8357,N_8234);
or U8655 (N_8655,N_8368,N_8069);
nor U8656 (N_8656,N_8160,N_8332);
nand U8657 (N_8657,N_8093,N_8425);
nand U8658 (N_8658,N_8236,N_8169);
nand U8659 (N_8659,N_8483,N_8480);
nand U8660 (N_8660,N_8195,N_8048);
nand U8661 (N_8661,N_8138,N_8399);
xnor U8662 (N_8662,N_8070,N_8328);
or U8663 (N_8663,N_8125,N_8334);
and U8664 (N_8664,N_8100,N_8418);
nand U8665 (N_8665,N_8032,N_8300);
xor U8666 (N_8666,N_8081,N_8194);
nand U8667 (N_8667,N_8180,N_8253);
nand U8668 (N_8668,N_8083,N_8178);
and U8669 (N_8669,N_8267,N_8233);
xor U8670 (N_8670,N_8123,N_8159);
and U8671 (N_8671,N_8172,N_8246);
nand U8672 (N_8672,N_8031,N_8305);
or U8673 (N_8673,N_8182,N_8014);
nor U8674 (N_8674,N_8082,N_8433);
xnor U8675 (N_8675,N_8010,N_8079);
nand U8676 (N_8676,N_8193,N_8026);
xnor U8677 (N_8677,N_8112,N_8485);
or U8678 (N_8678,N_8228,N_8340);
and U8679 (N_8679,N_8266,N_8118);
nand U8680 (N_8680,N_8287,N_8479);
xor U8681 (N_8681,N_8021,N_8099);
or U8682 (N_8682,N_8293,N_8219);
or U8683 (N_8683,N_8008,N_8094);
or U8684 (N_8684,N_8291,N_8390);
nand U8685 (N_8685,N_8416,N_8371);
or U8686 (N_8686,N_8106,N_8009);
nand U8687 (N_8687,N_8360,N_8383);
or U8688 (N_8688,N_8153,N_8431);
nor U8689 (N_8689,N_8059,N_8313);
xnor U8690 (N_8690,N_8452,N_8131);
nor U8691 (N_8691,N_8230,N_8104);
nand U8692 (N_8692,N_8391,N_8302);
and U8693 (N_8693,N_8137,N_8385);
or U8694 (N_8694,N_8337,N_8493);
xnor U8695 (N_8695,N_8398,N_8051);
and U8696 (N_8696,N_8215,N_8247);
nand U8697 (N_8697,N_8263,N_8344);
nor U8698 (N_8698,N_8114,N_8417);
nand U8699 (N_8699,N_8050,N_8457);
xor U8700 (N_8700,N_8279,N_8442);
or U8701 (N_8701,N_8462,N_8046);
xnor U8702 (N_8702,N_8342,N_8022);
nor U8703 (N_8703,N_8308,N_8474);
nor U8704 (N_8704,N_8224,N_8324);
nand U8705 (N_8705,N_8132,N_8315);
and U8706 (N_8706,N_8218,N_8444);
nand U8707 (N_8707,N_8386,N_8252);
and U8708 (N_8708,N_8455,N_8393);
nor U8709 (N_8709,N_8345,N_8467);
and U8710 (N_8710,N_8092,N_8078);
and U8711 (N_8711,N_8156,N_8134);
nand U8712 (N_8712,N_8484,N_8199);
and U8713 (N_8713,N_8307,N_8275);
and U8714 (N_8714,N_8367,N_8190);
nor U8715 (N_8715,N_8402,N_8460);
nand U8716 (N_8716,N_8211,N_8294);
nand U8717 (N_8717,N_8271,N_8220);
or U8718 (N_8718,N_8130,N_8213);
or U8719 (N_8719,N_8047,N_8490);
xor U8720 (N_8720,N_8097,N_8142);
xor U8721 (N_8721,N_8116,N_8284);
and U8722 (N_8722,N_8459,N_8214);
or U8723 (N_8723,N_8430,N_8437);
xor U8724 (N_8724,N_8184,N_8041);
nor U8725 (N_8725,N_8171,N_8012);
and U8726 (N_8726,N_8447,N_8152);
xnor U8727 (N_8727,N_8465,N_8422);
and U8728 (N_8728,N_8299,N_8161);
xor U8729 (N_8729,N_8202,N_8363);
or U8730 (N_8730,N_8005,N_8384);
or U8731 (N_8731,N_8301,N_8177);
and U8732 (N_8732,N_8027,N_8321);
nor U8733 (N_8733,N_8149,N_8419);
or U8734 (N_8734,N_8364,N_8489);
and U8735 (N_8735,N_8143,N_8054);
or U8736 (N_8736,N_8261,N_8196);
xnor U8737 (N_8737,N_8451,N_8406);
nor U8738 (N_8738,N_8472,N_8464);
nand U8739 (N_8739,N_8015,N_8441);
nor U8740 (N_8740,N_8117,N_8317);
nor U8741 (N_8741,N_8121,N_8320);
nand U8742 (N_8742,N_8068,N_8362);
xor U8743 (N_8743,N_8147,N_8037);
xor U8744 (N_8744,N_8276,N_8033);
or U8745 (N_8745,N_8126,N_8077);
nor U8746 (N_8746,N_8226,N_8354);
or U8747 (N_8747,N_8034,N_8335);
or U8748 (N_8748,N_8351,N_8343);
and U8749 (N_8749,N_8025,N_8446);
or U8750 (N_8750,N_8471,N_8419);
nand U8751 (N_8751,N_8218,N_8291);
nor U8752 (N_8752,N_8197,N_8461);
or U8753 (N_8753,N_8433,N_8229);
or U8754 (N_8754,N_8008,N_8107);
and U8755 (N_8755,N_8499,N_8212);
nand U8756 (N_8756,N_8460,N_8060);
and U8757 (N_8757,N_8348,N_8349);
and U8758 (N_8758,N_8066,N_8108);
nor U8759 (N_8759,N_8291,N_8326);
or U8760 (N_8760,N_8138,N_8416);
nor U8761 (N_8761,N_8096,N_8127);
xor U8762 (N_8762,N_8060,N_8238);
nor U8763 (N_8763,N_8284,N_8151);
and U8764 (N_8764,N_8341,N_8455);
nor U8765 (N_8765,N_8472,N_8489);
nor U8766 (N_8766,N_8467,N_8157);
xnor U8767 (N_8767,N_8091,N_8432);
or U8768 (N_8768,N_8274,N_8419);
nor U8769 (N_8769,N_8018,N_8239);
nand U8770 (N_8770,N_8188,N_8098);
nand U8771 (N_8771,N_8357,N_8417);
and U8772 (N_8772,N_8324,N_8323);
nor U8773 (N_8773,N_8482,N_8248);
nand U8774 (N_8774,N_8393,N_8059);
xnor U8775 (N_8775,N_8184,N_8495);
nor U8776 (N_8776,N_8240,N_8440);
and U8777 (N_8777,N_8230,N_8238);
nand U8778 (N_8778,N_8080,N_8372);
xnor U8779 (N_8779,N_8346,N_8353);
xnor U8780 (N_8780,N_8242,N_8206);
and U8781 (N_8781,N_8005,N_8332);
nor U8782 (N_8782,N_8109,N_8462);
or U8783 (N_8783,N_8473,N_8465);
or U8784 (N_8784,N_8173,N_8147);
xor U8785 (N_8785,N_8183,N_8333);
nor U8786 (N_8786,N_8014,N_8337);
nand U8787 (N_8787,N_8083,N_8156);
xor U8788 (N_8788,N_8292,N_8446);
nand U8789 (N_8789,N_8001,N_8442);
xnor U8790 (N_8790,N_8311,N_8233);
nor U8791 (N_8791,N_8155,N_8062);
nor U8792 (N_8792,N_8217,N_8475);
or U8793 (N_8793,N_8182,N_8064);
or U8794 (N_8794,N_8304,N_8026);
and U8795 (N_8795,N_8204,N_8328);
and U8796 (N_8796,N_8117,N_8185);
xnor U8797 (N_8797,N_8169,N_8446);
nand U8798 (N_8798,N_8401,N_8148);
or U8799 (N_8799,N_8075,N_8168);
nand U8800 (N_8800,N_8188,N_8486);
and U8801 (N_8801,N_8267,N_8468);
xnor U8802 (N_8802,N_8233,N_8249);
and U8803 (N_8803,N_8341,N_8054);
nand U8804 (N_8804,N_8152,N_8475);
nand U8805 (N_8805,N_8237,N_8064);
nand U8806 (N_8806,N_8305,N_8041);
xnor U8807 (N_8807,N_8013,N_8364);
and U8808 (N_8808,N_8163,N_8421);
xnor U8809 (N_8809,N_8084,N_8176);
or U8810 (N_8810,N_8048,N_8115);
or U8811 (N_8811,N_8037,N_8297);
or U8812 (N_8812,N_8230,N_8265);
and U8813 (N_8813,N_8070,N_8392);
and U8814 (N_8814,N_8479,N_8454);
and U8815 (N_8815,N_8495,N_8166);
nor U8816 (N_8816,N_8192,N_8188);
xnor U8817 (N_8817,N_8493,N_8128);
nand U8818 (N_8818,N_8408,N_8436);
nand U8819 (N_8819,N_8386,N_8171);
nor U8820 (N_8820,N_8055,N_8325);
or U8821 (N_8821,N_8058,N_8107);
or U8822 (N_8822,N_8479,N_8455);
xor U8823 (N_8823,N_8463,N_8211);
nor U8824 (N_8824,N_8120,N_8200);
and U8825 (N_8825,N_8366,N_8462);
nand U8826 (N_8826,N_8059,N_8072);
nor U8827 (N_8827,N_8342,N_8016);
nor U8828 (N_8828,N_8096,N_8363);
or U8829 (N_8829,N_8122,N_8158);
and U8830 (N_8830,N_8379,N_8087);
or U8831 (N_8831,N_8152,N_8131);
or U8832 (N_8832,N_8472,N_8075);
nor U8833 (N_8833,N_8032,N_8074);
xor U8834 (N_8834,N_8479,N_8061);
nor U8835 (N_8835,N_8402,N_8251);
xnor U8836 (N_8836,N_8498,N_8067);
and U8837 (N_8837,N_8203,N_8321);
nand U8838 (N_8838,N_8092,N_8284);
and U8839 (N_8839,N_8475,N_8073);
nand U8840 (N_8840,N_8277,N_8179);
nand U8841 (N_8841,N_8090,N_8203);
nand U8842 (N_8842,N_8044,N_8175);
nand U8843 (N_8843,N_8018,N_8370);
nor U8844 (N_8844,N_8244,N_8228);
nor U8845 (N_8845,N_8270,N_8045);
or U8846 (N_8846,N_8054,N_8466);
nand U8847 (N_8847,N_8405,N_8217);
xor U8848 (N_8848,N_8120,N_8227);
nor U8849 (N_8849,N_8417,N_8067);
nand U8850 (N_8850,N_8422,N_8288);
or U8851 (N_8851,N_8377,N_8131);
and U8852 (N_8852,N_8205,N_8359);
or U8853 (N_8853,N_8242,N_8371);
nand U8854 (N_8854,N_8010,N_8294);
and U8855 (N_8855,N_8302,N_8064);
nor U8856 (N_8856,N_8042,N_8077);
and U8857 (N_8857,N_8012,N_8052);
or U8858 (N_8858,N_8365,N_8250);
nor U8859 (N_8859,N_8102,N_8438);
or U8860 (N_8860,N_8001,N_8338);
xnor U8861 (N_8861,N_8298,N_8072);
xnor U8862 (N_8862,N_8351,N_8087);
nand U8863 (N_8863,N_8230,N_8323);
or U8864 (N_8864,N_8276,N_8429);
or U8865 (N_8865,N_8153,N_8449);
nor U8866 (N_8866,N_8494,N_8093);
xor U8867 (N_8867,N_8330,N_8447);
nor U8868 (N_8868,N_8255,N_8123);
and U8869 (N_8869,N_8042,N_8496);
xor U8870 (N_8870,N_8040,N_8095);
or U8871 (N_8871,N_8322,N_8002);
nand U8872 (N_8872,N_8210,N_8083);
or U8873 (N_8873,N_8145,N_8100);
nand U8874 (N_8874,N_8179,N_8359);
and U8875 (N_8875,N_8224,N_8403);
and U8876 (N_8876,N_8331,N_8157);
nand U8877 (N_8877,N_8324,N_8036);
and U8878 (N_8878,N_8478,N_8154);
nor U8879 (N_8879,N_8033,N_8248);
nor U8880 (N_8880,N_8032,N_8332);
nand U8881 (N_8881,N_8311,N_8293);
nor U8882 (N_8882,N_8235,N_8138);
nor U8883 (N_8883,N_8432,N_8280);
or U8884 (N_8884,N_8031,N_8453);
nand U8885 (N_8885,N_8060,N_8139);
nor U8886 (N_8886,N_8449,N_8429);
xor U8887 (N_8887,N_8123,N_8378);
and U8888 (N_8888,N_8401,N_8047);
or U8889 (N_8889,N_8430,N_8266);
nand U8890 (N_8890,N_8391,N_8055);
and U8891 (N_8891,N_8025,N_8294);
xor U8892 (N_8892,N_8040,N_8154);
or U8893 (N_8893,N_8376,N_8253);
and U8894 (N_8894,N_8299,N_8229);
and U8895 (N_8895,N_8238,N_8463);
nand U8896 (N_8896,N_8055,N_8174);
or U8897 (N_8897,N_8280,N_8238);
nor U8898 (N_8898,N_8131,N_8133);
or U8899 (N_8899,N_8106,N_8192);
or U8900 (N_8900,N_8144,N_8363);
nor U8901 (N_8901,N_8193,N_8104);
nand U8902 (N_8902,N_8400,N_8417);
nor U8903 (N_8903,N_8414,N_8072);
nand U8904 (N_8904,N_8322,N_8427);
or U8905 (N_8905,N_8012,N_8006);
or U8906 (N_8906,N_8126,N_8399);
nand U8907 (N_8907,N_8034,N_8321);
nand U8908 (N_8908,N_8134,N_8266);
or U8909 (N_8909,N_8124,N_8104);
or U8910 (N_8910,N_8338,N_8208);
nand U8911 (N_8911,N_8165,N_8440);
xnor U8912 (N_8912,N_8028,N_8224);
xor U8913 (N_8913,N_8475,N_8453);
xnor U8914 (N_8914,N_8462,N_8086);
nand U8915 (N_8915,N_8386,N_8259);
nand U8916 (N_8916,N_8115,N_8107);
nor U8917 (N_8917,N_8262,N_8037);
xnor U8918 (N_8918,N_8050,N_8344);
or U8919 (N_8919,N_8124,N_8464);
nand U8920 (N_8920,N_8046,N_8279);
xor U8921 (N_8921,N_8427,N_8074);
nand U8922 (N_8922,N_8441,N_8251);
nor U8923 (N_8923,N_8487,N_8440);
xor U8924 (N_8924,N_8185,N_8402);
and U8925 (N_8925,N_8077,N_8057);
nand U8926 (N_8926,N_8283,N_8326);
xor U8927 (N_8927,N_8174,N_8268);
xnor U8928 (N_8928,N_8489,N_8152);
or U8929 (N_8929,N_8364,N_8376);
xnor U8930 (N_8930,N_8394,N_8315);
nand U8931 (N_8931,N_8064,N_8345);
or U8932 (N_8932,N_8185,N_8060);
or U8933 (N_8933,N_8011,N_8401);
or U8934 (N_8934,N_8039,N_8371);
or U8935 (N_8935,N_8139,N_8070);
and U8936 (N_8936,N_8075,N_8192);
and U8937 (N_8937,N_8430,N_8476);
nor U8938 (N_8938,N_8428,N_8088);
xnor U8939 (N_8939,N_8309,N_8297);
xnor U8940 (N_8940,N_8090,N_8001);
and U8941 (N_8941,N_8453,N_8231);
and U8942 (N_8942,N_8169,N_8099);
nor U8943 (N_8943,N_8364,N_8057);
or U8944 (N_8944,N_8293,N_8079);
nor U8945 (N_8945,N_8454,N_8006);
and U8946 (N_8946,N_8499,N_8020);
xnor U8947 (N_8947,N_8320,N_8018);
nand U8948 (N_8948,N_8378,N_8027);
or U8949 (N_8949,N_8360,N_8100);
xor U8950 (N_8950,N_8372,N_8066);
nand U8951 (N_8951,N_8099,N_8398);
nor U8952 (N_8952,N_8219,N_8123);
or U8953 (N_8953,N_8196,N_8385);
nand U8954 (N_8954,N_8097,N_8386);
nand U8955 (N_8955,N_8378,N_8275);
or U8956 (N_8956,N_8090,N_8066);
nor U8957 (N_8957,N_8063,N_8058);
xor U8958 (N_8958,N_8440,N_8226);
nand U8959 (N_8959,N_8226,N_8322);
nand U8960 (N_8960,N_8009,N_8383);
xnor U8961 (N_8961,N_8167,N_8161);
nor U8962 (N_8962,N_8389,N_8244);
and U8963 (N_8963,N_8469,N_8350);
and U8964 (N_8964,N_8042,N_8432);
and U8965 (N_8965,N_8013,N_8410);
or U8966 (N_8966,N_8130,N_8344);
xor U8967 (N_8967,N_8494,N_8053);
nor U8968 (N_8968,N_8257,N_8369);
xor U8969 (N_8969,N_8448,N_8484);
or U8970 (N_8970,N_8352,N_8314);
nand U8971 (N_8971,N_8088,N_8315);
or U8972 (N_8972,N_8199,N_8170);
xor U8973 (N_8973,N_8210,N_8327);
and U8974 (N_8974,N_8137,N_8414);
nor U8975 (N_8975,N_8356,N_8284);
nand U8976 (N_8976,N_8146,N_8181);
nor U8977 (N_8977,N_8182,N_8346);
or U8978 (N_8978,N_8424,N_8056);
nand U8979 (N_8979,N_8239,N_8192);
nand U8980 (N_8980,N_8089,N_8125);
nor U8981 (N_8981,N_8224,N_8095);
and U8982 (N_8982,N_8105,N_8259);
or U8983 (N_8983,N_8155,N_8267);
nor U8984 (N_8984,N_8175,N_8261);
and U8985 (N_8985,N_8212,N_8003);
or U8986 (N_8986,N_8378,N_8130);
nor U8987 (N_8987,N_8323,N_8241);
nand U8988 (N_8988,N_8223,N_8197);
or U8989 (N_8989,N_8172,N_8391);
xor U8990 (N_8990,N_8451,N_8184);
xor U8991 (N_8991,N_8080,N_8303);
and U8992 (N_8992,N_8482,N_8412);
and U8993 (N_8993,N_8117,N_8284);
xnor U8994 (N_8994,N_8238,N_8445);
and U8995 (N_8995,N_8335,N_8047);
nand U8996 (N_8996,N_8077,N_8113);
xnor U8997 (N_8997,N_8378,N_8186);
and U8998 (N_8998,N_8062,N_8052);
nor U8999 (N_8999,N_8220,N_8496);
nand U9000 (N_9000,N_8862,N_8614);
xnor U9001 (N_9001,N_8979,N_8528);
nand U9002 (N_9002,N_8651,N_8589);
and U9003 (N_9003,N_8695,N_8908);
and U9004 (N_9004,N_8945,N_8629);
xor U9005 (N_9005,N_8621,N_8636);
and U9006 (N_9006,N_8673,N_8775);
and U9007 (N_9007,N_8592,N_8573);
and U9008 (N_9008,N_8677,N_8674);
nor U9009 (N_9009,N_8955,N_8782);
nand U9010 (N_9010,N_8502,N_8851);
nor U9011 (N_9011,N_8856,N_8549);
nor U9012 (N_9012,N_8902,N_8607);
or U9013 (N_9013,N_8662,N_8526);
and U9014 (N_9014,N_8951,N_8828);
and U9015 (N_9015,N_8714,N_8801);
or U9016 (N_9016,N_8918,N_8761);
and U9017 (N_9017,N_8909,N_8732);
nand U9018 (N_9018,N_8789,N_8539);
or U9019 (N_9019,N_8817,N_8799);
xnor U9020 (N_9020,N_8527,N_8833);
xnor U9021 (N_9021,N_8579,N_8750);
nor U9022 (N_9022,N_8944,N_8810);
or U9023 (N_9023,N_8722,N_8938);
xor U9024 (N_9024,N_8886,N_8755);
nand U9025 (N_9025,N_8564,N_8509);
and U9026 (N_9026,N_8720,N_8889);
or U9027 (N_9027,N_8942,N_8839);
nand U9028 (N_9028,N_8622,N_8800);
xnor U9029 (N_9029,N_8552,N_8704);
nand U9030 (N_9030,N_8758,N_8748);
xnor U9031 (N_9031,N_8587,N_8570);
xnor U9032 (N_9032,N_8688,N_8683);
nor U9033 (N_9033,N_8668,N_8956);
nand U9034 (N_9034,N_8531,N_8814);
xnor U9035 (N_9035,N_8515,N_8980);
nor U9036 (N_9036,N_8615,N_8725);
nor U9037 (N_9037,N_8734,N_8964);
nor U9038 (N_9038,N_8591,N_8791);
xor U9039 (N_9039,N_8792,N_8554);
nor U9040 (N_9040,N_8779,N_8565);
nor U9041 (N_9041,N_8705,N_8927);
xor U9042 (N_9042,N_8895,N_8678);
or U9043 (N_9043,N_8894,N_8638);
xor U9044 (N_9044,N_8920,N_8768);
and U9045 (N_9045,N_8596,N_8763);
or U9046 (N_9046,N_8572,N_8780);
xnor U9047 (N_9047,N_8597,N_8633);
nor U9048 (N_9048,N_8628,N_8530);
nor U9049 (N_9049,N_8544,N_8861);
or U9050 (N_9050,N_8546,N_8957);
or U9051 (N_9051,N_8643,N_8648);
and U9052 (N_9052,N_8906,N_8512);
xnor U9053 (N_9053,N_8609,N_8642);
nor U9054 (N_9054,N_8696,N_8612);
xnor U9055 (N_9055,N_8649,N_8953);
nand U9056 (N_9056,N_8690,N_8872);
and U9057 (N_9057,N_8762,N_8736);
nand U9058 (N_9058,N_8699,N_8910);
nor U9059 (N_9059,N_8666,N_8965);
nand U9060 (N_9060,N_8984,N_8553);
xnor U9061 (N_9061,N_8706,N_8811);
nor U9062 (N_9062,N_8555,N_8912);
xnor U9063 (N_9063,N_8901,N_8557);
and U9064 (N_9064,N_8876,N_8790);
and U9065 (N_9065,N_8771,N_8961);
or U9066 (N_9066,N_8610,N_8516);
or U9067 (N_9067,N_8796,N_8988);
or U9068 (N_9068,N_8939,N_8647);
nor U9069 (N_9069,N_8737,N_8693);
or U9070 (N_9070,N_8517,N_8905);
and U9071 (N_9071,N_8744,N_8657);
nor U9072 (N_9072,N_8653,N_8826);
nor U9073 (N_9073,N_8702,N_8936);
xnor U9074 (N_9074,N_8679,N_8583);
xor U9075 (N_9075,N_8694,N_8904);
xor U9076 (N_9076,N_8576,N_8729);
nand U9077 (N_9077,N_8585,N_8680);
or U9078 (N_9078,N_8562,N_8989);
or U9079 (N_9079,N_8926,N_8917);
nor U9080 (N_9080,N_8978,N_8928);
nor U9081 (N_9081,N_8787,N_8716);
nor U9082 (N_9082,N_8740,N_8924);
and U9083 (N_9083,N_8578,N_8805);
and U9084 (N_9084,N_8522,N_8825);
xor U9085 (N_9085,N_8880,N_8981);
or U9086 (N_9086,N_8563,N_8869);
or U9087 (N_9087,N_8560,N_8850);
xor U9088 (N_9088,N_8903,N_8946);
nor U9089 (N_9089,N_8923,N_8631);
or U9090 (N_9090,N_8671,N_8672);
and U9091 (N_9091,N_8646,N_8540);
nand U9092 (N_9092,N_8745,N_8593);
nor U9093 (N_9093,N_8871,N_8670);
or U9094 (N_9094,N_8602,N_8599);
nor U9095 (N_9095,N_8764,N_8739);
xnor U9096 (N_9096,N_8533,N_8626);
nor U9097 (N_9097,N_8959,N_8824);
and U9098 (N_9098,N_8529,N_8934);
or U9099 (N_9099,N_8543,N_8689);
or U9100 (N_9100,N_8568,N_8849);
and U9101 (N_9101,N_8523,N_8885);
and U9102 (N_9102,N_8566,N_8759);
nand U9103 (N_9103,N_8827,N_8507);
nand U9104 (N_9104,N_8542,N_8658);
xnor U9105 (N_9105,N_8977,N_8534);
or U9106 (N_9106,N_8518,N_8687);
and U9107 (N_9107,N_8931,N_8947);
and U9108 (N_9108,N_8753,N_8855);
and U9109 (N_9109,N_8835,N_8752);
or U9110 (N_9110,N_8558,N_8656);
nand U9111 (N_9111,N_8586,N_8832);
nor U9112 (N_9112,N_8630,N_8685);
xnor U9113 (N_9113,N_8611,N_8550);
xnor U9114 (N_9114,N_8575,N_8911);
nand U9115 (N_9115,N_8858,N_8857);
nor U9116 (N_9116,N_8632,N_8510);
xor U9117 (N_9117,N_8898,N_8907);
xnor U9118 (N_9118,N_8940,N_8669);
nand U9119 (N_9119,N_8803,N_8937);
nand U9120 (N_9120,N_8598,N_8506);
xnor U9121 (N_9121,N_8691,N_8974);
or U9122 (N_9122,N_8588,N_8710);
and U9123 (N_9123,N_8618,N_8818);
xor U9124 (N_9124,N_8503,N_8584);
or U9125 (N_9125,N_8783,N_8726);
nand U9126 (N_9126,N_8508,N_8514);
xnor U9127 (N_9127,N_8891,N_8532);
xor U9128 (N_9128,N_8865,N_8500);
nand U9129 (N_9129,N_8859,N_8949);
and U9130 (N_9130,N_8541,N_8738);
nand U9131 (N_9131,N_8843,N_8773);
or U9132 (N_9132,N_8742,N_8641);
xnor U9133 (N_9133,N_8661,N_8713);
nand U9134 (N_9134,N_8548,N_8590);
and U9135 (N_9135,N_8838,N_8774);
or U9136 (N_9136,N_8581,N_8829);
or U9137 (N_9137,N_8561,N_8650);
xor U9138 (N_9138,N_8802,N_8770);
nor U9139 (N_9139,N_8766,N_8660);
xnor U9140 (N_9140,N_8958,N_8921);
nand U9141 (N_9141,N_8966,N_8987);
xor U9142 (N_9142,N_8606,N_8983);
and U9143 (N_9143,N_8675,N_8997);
or U9144 (N_9144,N_8892,N_8837);
or U9145 (N_9145,N_8950,N_8930);
and U9146 (N_9146,N_8777,N_8878);
xor U9147 (N_9147,N_8623,N_8747);
and U9148 (N_9148,N_8804,N_8913);
xor U9149 (N_9149,N_8972,N_8812);
or U9150 (N_9150,N_8976,N_8664);
and U9151 (N_9151,N_8899,N_8929);
and U9152 (N_9152,N_8816,N_8767);
and U9153 (N_9153,N_8698,N_8733);
xnor U9154 (N_9154,N_8807,N_8735);
nand U9155 (N_9155,N_8990,N_8854);
xnor U9156 (N_9156,N_8501,N_8605);
and U9157 (N_9157,N_8709,N_8846);
or U9158 (N_9158,N_8969,N_8708);
xor U9159 (N_9159,N_8724,N_8985);
xnor U9160 (N_9160,N_8692,N_8915);
nand U9161 (N_9161,N_8707,N_8995);
nor U9162 (N_9162,N_8538,N_8654);
xnor U9163 (N_9163,N_8844,N_8577);
and U9164 (N_9164,N_8848,N_8967);
nand U9165 (N_9165,N_8952,N_8613);
nand U9166 (N_9166,N_8922,N_8754);
nor U9167 (N_9167,N_8809,N_8556);
nor U9168 (N_9168,N_8594,N_8819);
nor U9169 (N_9169,N_8867,N_8667);
nor U9170 (N_9170,N_8935,N_8941);
nand U9171 (N_9171,N_8703,N_8619);
and U9172 (N_9172,N_8896,N_8731);
nand U9173 (N_9173,N_8875,N_8793);
nor U9174 (N_9174,N_8652,N_8511);
xor U9175 (N_9175,N_8879,N_8993);
or U9176 (N_9176,N_8537,N_8884);
nor U9177 (N_9177,N_8840,N_8676);
and U9178 (N_9178,N_8962,N_8645);
nor U9179 (N_9179,N_8883,N_8973);
or U9180 (N_9180,N_8785,N_8971);
nand U9181 (N_9181,N_8841,N_8788);
nand U9182 (N_9182,N_8808,N_8644);
xor U9183 (N_9183,N_8784,N_8608);
xnor U9184 (N_9184,N_8757,N_8525);
xnor U9185 (N_9185,N_8914,N_8786);
nor U9186 (N_9186,N_8756,N_8975);
and U9187 (N_9187,N_8524,N_8797);
and U9188 (N_9188,N_8635,N_8868);
xnor U9189 (N_9189,N_8870,N_8682);
nand U9190 (N_9190,N_8842,N_8919);
nand U9191 (N_9191,N_8877,N_8681);
and U9192 (N_9192,N_8864,N_8998);
or U9193 (N_9193,N_8806,N_8637);
nor U9194 (N_9194,N_8603,N_8863);
or U9195 (N_9195,N_8519,N_8569);
xor U9196 (N_9196,N_8600,N_8847);
nor U9197 (N_9197,N_8772,N_8640);
nand U9198 (N_9198,N_8749,N_8994);
xor U9199 (N_9199,N_8730,N_8711);
and U9200 (N_9200,N_8574,N_8624);
nor U9201 (N_9201,N_8992,N_8659);
or U9202 (N_9202,N_8625,N_8996);
or U9203 (N_9203,N_8852,N_8547);
or U9204 (N_9204,N_8513,N_8727);
nand U9205 (N_9205,N_8617,N_8684);
or U9206 (N_9206,N_8604,N_8504);
nand U9207 (N_9207,N_8821,N_8697);
and U9208 (N_9208,N_8890,N_8582);
nor U9209 (N_9209,N_8834,N_8535);
and U9210 (N_9210,N_8776,N_8822);
and U9211 (N_9211,N_8545,N_8663);
nor U9212 (N_9212,N_8897,N_8986);
nand U9213 (N_9213,N_8751,N_8700);
xor U9214 (N_9214,N_8743,N_8968);
or U9215 (N_9215,N_8970,N_8718);
and U9216 (N_9216,N_8798,N_8823);
or U9217 (N_9217,N_8571,N_8845);
nor U9218 (N_9218,N_8815,N_8712);
nor U9219 (N_9219,N_8620,N_8916);
xor U9220 (N_9220,N_8595,N_8580);
and U9221 (N_9221,N_8874,N_8888);
and U9222 (N_9222,N_8634,N_8616);
and U9223 (N_9223,N_8794,N_8887);
or U9224 (N_9224,N_8536,N_8723);
xnor U9225 (N_9225,N_8741,N_8963);
or U9226 (N_9226,N_8701,N_8567);
nand U9227 (N_9227,N_8639,N_8719);
nor U9228 (N_9228,N_8601,N_8520);
nand U9229 (N_9229,N_8830,N_8900);
nor U9230 (N_9230,N_8925,N_8948);
or U9231 (N_9231,N_8881,N_8760);
nor U9232 (N_9232,N_8778,N_8866);
nor U9233 (N_9233,N_8893,N_8686);
xor U9234 (N_9234,N_8860,N_8559);
xnor U9235 (N_9235,N_8717,N_8715);
xor U9236 (N_9236,N_8943,N_8627);
and U9237 (N_9237,N_8769,N_8932);
nor U9238 (N_9238,N_8765,N_8960);
nor U9239 (N_9239,N_8933,N_8873);
or U9240 (N_9240,N_8820,N_8954);
or U9241 (N_9241,N_8991,N_8521);
xor U9242 (N_9242,N_8781,N_8982);
xnor U9243 (N_9243,N_8836,N_8505);
nand U9244 (N_9244,N_8882,N_8795);
and U9245 (N_9245,N_8746,N_8813);
and U9246 (N_9246,N_8853,N_8721);
xnor U9247 (N_9247,N_8665,N_8831);
xnor U9248 (N_9248,N_8551,N_8999);
and U9249 (N_9249,N_8728,N_8655);
xor U9250 (N_9250,N_8695,N_8768);
xor U9251 (N_9251,N_8612,N_8970);
and U9252 (N_9252,N_8924,N_8937);
nor U9253 (N_9253,N_8742,N_8650);
xnor U9254 (N_9254,N_8530,N_8549);
or U9255 (N_9255,N_8656,N_8647);
and U9256 (N_9256,N_8996,N_8995);
and U9257 (N_9257,N_8808,N_8826);
xnor U9258 (N_9258,N_8887,N_8668);
and U9259 (N_9259,N_8723,N_8728);
nor U9260 (N_9260,N_8568,N_8873);
and U9261 (N_9261,N_8816,N_8963);
and U9262 (N_9262,N_8989,N_8819);
and U9263 (N_9263,N_8993,N_8830);
or U9264 (N_9264,N_8526,N_8845);
xor U9265 (N_9265,N_8502,N_8569);
nor U9266 (N_9266,N_8704,N_8526);
nor U9267 (N_9267,N_8774,N_8754);
nor U9268 (N_9268,N_8724,N_8606);
or U9269 (N_9269,N_8880,N_8754);
nand U9270 (N_9270,N_8839,N_8577);
nand U9271 (N_9271,N_8864,N_8569);
and U9272 (N_9272,N_8571,N_8559);
nor U9273 (N_9273,N_8636,N_8507);
or U9274 (N_9274,N_8836,N_8835);
xnor U9275 (N_9275,N_8715,N_8630);
nor U9276 (N_9276,N_8798,N_8880);
xor U9277 (N_9277,N_8873,N_8643);
xnor U9278 (N_9278,N_8760,N_8555);
or U9279 (N_9279,N_8925,N_8531);
nand U9280 (N_9280,N_8576,N_8552);
nand U9281 (N_9281,N_8848,N_8925);
and U9282 (N_9282,N_8691,N_8940);
xnor U9283 (N_9283,N_8589,N_8690);
nor U9284 (N_9284,N_8520,N_8674);
or U9285 (N_9285,N_8932,N_8839);
nor U9286 (N_9286,N_8730,N_8562);
nor U9287 (N_9287,N_8802,N_8749);
and U9288 (N_9288,N_8810,N_8581);
xnor U9289 (N_9289,N_8716,N_8544);
and U9290 (N_9290,N_8712,N_8652);
nand U9291 (N_9291,N_8703,N_8655);
or U9292 (N_9292,N_8933,N_8724);
nand U9293 (N_9293,N_8928,N_8878);
nor U9294 (N_9294,N_8984,N_8925);
nand U9295 (N_9295,N_8949,N_8576);
or U9296 (N_9296,N_8674,N_8968);
nor U9297 (N_9297,N_8778,N_8543);
or U9298 (N_9298,N_8760,N_8736);
nor U9299 (N_9299,N_8829,N_8927);
nand U9300 (N_9300,N_8975,N_8733);
nand U9301 (N_9301,N_8624,N_8554);
nand U9302 (N_9302,N_8525,N_8733);
nor U9303 (N_9303,N_8783,N_8931);
nor U9304 (N_9304,N_8592,N_8699);
or U9305 (N_9305,N_8899,N_8569);
nand U9306 (N_9306,N_8780,N_8662);
and U9307 (N_9307,N_8988,N_8856);
nand U9308 (N_9308,N_8522,N_8939);
nand U9309 (N_9309,N_8658,N_8510);
or U9310 (N_9310,N_8677,N_8859);
xnor U9311 (N_9311,N_8959,N_8618);
nor U9312 (N_9312,N_8864,N_8891);
or U9313 (N_9313,N_8694,N_8639);
xnor U9314 (N_9314,N_8704,N_8514);
or U9315 (N_9315,N_8542,N_8780);
and U9316 (N_9316,N_8967,N_8907);
nor U9317 (N_9317,N_8571,N_8765);
xor U9318 (N_9318,N_8803,N_8735);
or U9319 (N_9319,N_8834,N_8784);
or U9320 (N_9320,N_8622,N_8974);
and U9321 (N_9321,N_8970,N_8631);
and U9322 (N_9322,N_8831,N_8532);
or U9323 (N_9323,N_8596,N_8654);
or U9324 (N_9324,N_8622,N_8593);
xnor U9325 (N_9325,N_8851,N_8867);
xor U9326 (N_9326,N_8914,N_8823);
xor U9327 (N_9327,N_8531,N_8894);
xnor U9328 (N_9328,N_8841,N_8533);
and U9329 (N_9329,N_8840,N_8856);
nor U9330 (N_9330,N_8574,N_8908);
nor U9331 (N_9331,N_8766,N_8585);
and U9332 (N_9332,N_8953,N_8801);
xnor U9333 (N_9333,N_8599,N_8837);
nand U9334 (N_9334,N_8501,N_8877);
nor U9335 (N_9335,N_8588,N_8787);
or U9336 (N_9336,N_8684,N_8960);
nand U9337 (N_9337,N_8510,N_8589);
or U9338 (N_9338,N_8840,N_8950);
and U9339 (N_9339,N_8603,N_8763);
nand U9340 (N_9340,N_8634,N_8958);
nand U9341 (N_9341,N_8767,N_8650);
and U9342 (N_9342,N_8765,N_8827);
and U9343 (N_9343,N_8737,N_8878);
or U9344 (N_9344,N_8895,N_8970);
nor U9345 (N_9345,N_8984,N_8700);
and U9346 (N_9346,N_8541,N_8636);
nand U9347 (N_9347,N_8582,N_8608);
and U9348 (N_9348,N_8848,N_8895);
and U9349 (N_9349,N_8947,N_8511);
and U9350 (N_9350,N_8943,N_8855);
nand U9351 (N_9351,N_8734,N_8847);
nor U9352 (N_9352,N_8526,N_8838);
xor U9353 (N_9353,N_8529,N_8515);
nor U9354 (N_9354,N_8560,N_8857);
or U9355 (N_9355,N_8569,N_8983);
nor U9356 (N_9356,N_8800,N_8634);
and U9357 (N_9357,N_8647,N_8774);
xor U9358 (N_9358,N_8879,N_8899);
nand U9359 (N_9359,N_8743,N_8708);
nor U9360 (N_9360,N_8540,N_8614);
or U9361 (N_9361,N_8812,N_8566);
or U9362 (N_9362,N_8859,N_8766);
and U9363 (N_9363,N_8856,N_8500);
or U9364 (N_9364,N_8922,N_8877);
xor U9365 (N_9365,N_8743,N_8876);
or U9366 (N_9366,N_8635,N_8611);
xor U9367 (N_9367,N_8521,N_8712);
or U9368 (N_9368,N_8690,N_8819);
nor U9369 (N_9369,N_8510,N_8546);
nand U9370 (N_9370,N_8622,N_8535);
nand U9371 (N_9371,N_8734,N_8536);
nand U9372 (N_9372,N_8599,N_8703);
nor U9373 (N_9373,N_8668,N_8670);
nand U9374 (N_9374,N_8510,N_8985);
xor U9375 (N_9375,N_8864,N_8742);
or U9376 (N_9376,N_8567,N_8815);
nand U9377 (N_9377,N_8918,N_8535);
nor U9378 (N_9378,N_8703,N_8500);
nand U9379 (N_9379,N_8812,N_8510);
xnor U9380 (N_9380,N_8621,N_8526);
or U9381 (N_9381,N_8747,N_8706);
xnor U9382 (N_9382,N_8945,N_8748);
nand U9383 (N_9383,N_8617,N_8699);
or U9384 (N_9384,N_8853,N_8650);
and U9385 (N_9385,N_8694,N_8743);
nand U9386 (N_9386,N_8865,N_8984);
xor U9387 (N_9387,N_8870,N_8627);
or U9388 (N_9388,N_8715,N_8786);
and U9389 (N_9389,N_8769,N_8697);
or U9390 (N_9390,N_8780,N_8589);
or U9391 (N_9391,N_8825,N_8973);
nand U9392 (N_9392,N_8574,N_8769);
xnor U9393 (N_9393,N_8917,N_8628);
nand U9394 (N_9394,N_8669,N_8702);
and U9395 (N_9395,N_8798,N_8996);
nor U9396 (N_9396,N_8602,N_8987);
or U9397 (N_9397,N_8612,N_8746);
nor U9398 (N_9398,N_8791,N_8583);
xnor U9399 (N_9399,N_8654,N_8723);
or U9400 (N_9400,N_8564,N_8759);
xnor U9401 (N_9401,N_8885,N_8621);
xor U9402 (N_9402,N_8743,N_8830);
nand U9403 (N_9403,N_8715,N_8535);
nand U9404 (N_9404,N_8961,N_8615);
and U9405 (N_9405,N_8580,N_8703);
nor U9406 (N_9406,N_8572,N_8536);
nand U9407 (N_9407,N_8974,N_8979);
or U9408 (N_9408,N_8835,N_8677);
and U9409 (N_9409,N_8619,N_8628);
xor U9410 (N_9410,N_8763,N_8910);
xnor U9411 (N_9411,N_8948,N_8953);
and U9412 (N_9412,N_8621,N_8518);
and U9413 (N_9413,N_8722,N_8881);
xor U9414 (N_9414,N_8595,N_8743);
nor U9415 (N_9415,N_8875,N_8971);
and U9416 (N_9416,N_8761,N_8860);
or U9417 (N_9417,N_8815,N_8696);
xnor U9418 (N_9418,N_8650,N_8913);
nand U9419 (N_9419,N_8841,N_8601);
nand U9420 (N_9420,N_8872,N_8774);
and U9421 (N_9421,N_8737,N_8976);
and U9422 (N_9422,N_8712,N_8922);
xor U9423 (N_9423,N_8852,N_8893);
or U9424 (N_9424,N_8724,N_8950);
and U9425 (N_9425,N_8929,N_8872);
or U9426 (N_9426,N_8931,N_8944);
nand U9427 (N_9427,N_8982,N_8924);
xnor U9428 (N_9428,N_8997,N_8577);
xor U9429 (N_9429,N_8783,N_8523);
xor U9430 (N_9430,N_8561,N_8842);
nand U9431 (N_9431,N_8716,N_8949);
and U9432 (N_9432,N_8710,N_8687);
or U9433 (N_9433,N_8807,N_8768);
nor U9434 (N_9434,N_8816,N_8765);
nand U9435 (N_9435,N_8946,N_8525);
and U9436 (N_9436,N_8567,N_8644);
and U9437 (N_9437,N_8635,N_8686);
nand U9438 (N_9438,N_8511,N_8827);
and U9439 (N_9439,N_8741,N_8994);
nor U9440 (N_9440,N_8941,N_8806);
xor U9441 (N_9441,N_8872,N_8653);
and U9442 (N_9442,N_8519,N_8520);
or U9443 (N_9443,N_8865,N_8744);
xnor U9444 (N_9444,N_8680,N_8807);
xnor U9445 (N_9445,N_8568,N_8857);
nand U9446 (N_9446,N_8728,N_8967);
and U9447 (N_9447,N_8667,N_8967);
nor U9448 (N_9448,N_8530,N_8842);
xor U9449 (N_9449,N_8596,N_8747);
xnor U9450 (N_9450,N_8975,N_8597);
nor U9451 (N_9451,N_8899,N_8837);
xnor U9452 (N_9452,N_8675,N_8676);
or U9453 (N_9453,N_8860,N_8964);
nand U9454 (N_9454,N_8837,N_8989);
nor U9455 (N_9455,N_8540,N_8558);
nand U9456 (N_9456,N_8866,N_8537);
or U9457 (N_9457,N_8570,N_8877);
nor U9458 (N_9458,N_8659,N_8687);
nand U9459 (N_9459,N_8738,N_8669);
nor U9460 (N_9460,N_8567,N_8593);
nor U9461 (N_9461,N_8799,N_8792);
nand U9462 (N_9462,N_8858,N_8664);
nor U9463 (N_9463,N_8950,N_8800);
nor U9464 (N_9464,N_8761,N_8954);
and U9465 (N_9465,N_8724,N_8673);
nor U9466 (N_9466,N_8691,N_8966);
or U9467 (N_9467,N_8755,N_8579);
or U9468 (N_9468,N_8639,N_8814);
nor U9469 (N_9469,N_8784,N_8962);
xnor U9470 (N_9470,N_8646,N_8932);
nand U9471 (N_9471,N_8881,N_8867);
nor U9472 (N_9472,N_8812,N_8855);
nor U9473 (N_9473,N_8617,N_8730);
nor U9474 (N_9474,N_8669,N_8980);
xor U9475 (N_9475,N_8943,N_8813);
or U9476 (N_9476,N_8805,N_8843);
nor U9477 (N_9477,N_8923,N_8596);
nand U9478 (N_9478,N_8934,N_8809);
xnor U9479 (N_9479,N_8827,N_8992);
xor U9480 (N_9480,N_8873,N_8652);
and U9481 (N_9481,N_8878,N_8590);
nand U9482 (N_9482,N_8755,N_8945);
nor U9483 (N_9483,N_8756,N_8606);
nor U9484 (N_9484,N_8513,N_8768);
or U9485 (N_9485,N_8568,N_8972);
xor U9486 (N_9486,N_8644,N_8834);
nor U9487 (N_9487,N_8574,N_8601);
nand U9488 (N_9488,N_8510,N_8872);
nand U9489 (N_9489,N_8552,N_8658);
and U9490 (N_9490,N_8876,N_8694);
nor U9491 (N_9491,N_8938,N_8715);
or U9492 (N_9492,N_8995,N_8606);
and U9493 (N_9493,N_8925,N_8577);
nand U9494 (N_9494,N_8820,N_8673);
nand U9495 (N_9495,N_8890,N_8518);
nor U9496 (N_9496,N_8969,N_8761);
xnor U9497 (N_9497,N_8749,N_8785);
nor U9498 (N_9498,N_8976,N_8993);
nor U9499 (N_9499,N_8743,N_8671);
nor U9500 (N_9500,N_9201,N_9015);
nor U9501 (N_9501,N_9188,N_9086);
xor U9502 (N_9502,N_9359,N_9435);
xnor U9503 (N_9503,N_9319,N_9455);
xor U9504 (N_9504,N_9356,N_9093);
and U9505 (N_9505,N_9495,N_9223);
nor U9506 (N_9506,N_9183,N_9151);
nand U9507 (N_9507,N_9074,N_9083);
and U9508 (N_9508,N_9384,N_9366);
or U9509 (N_9509,N_9382,N_9293);
xor U9510 (N_9510,N_9374,N_9002);
nand U9511 (N_9511,N_9161,N_9367);
or U9512 (N_9512,N_9088,N_9462);
and U9513 (N_9513,N_9019,N_9412);
nor U9514 (N_9514,N_9163,N_9392);
nor U9515 (N_9515,N_9368,N_9059);
or U9516 (N_9516,N_9242,N_9136);
and U9517 (N_9517,N_9140,N_9459);
nor U9518 (N_9518,N_9383,N_9021);
and U9519 (N_9519,N_9341,N_9207);
nor U9520 (N_9520,N_9113,N_9193);
nor U9521 (N_9521,N_9471,N_9029);
and U9522 (N_9522,N_9234,N_9154);
xnor U9523 (N_9523,N_9477,N_9038);
or U9524 (N_9524,N_9022,N_9164);
xnor U9525 (N_9525,N_9122,N_9134);
and U9526 (N_9526,N_9402,N_9291);
nand U9527 (N_9527,N_9473,N_9011);
or U9528 (N_9528,N_9103,N_9185);
xor U9529 (N_9529,N_9347,N_9407);
nand U9530 (N_9530,N_9449,N_9492);
xnor U9531 (N_9531,N_9419,N_9309);
xor U9532 (N_9532,N_9068,N_9283);
xor U9533 (N_9533,N_9245,N_9428);
nor U9534 (N_9534,N_9219,N_9155);
or U9535 (N_9535,N_9150,N_9067);
xor U9536 (N_9536,N_9296,N_9196);
xnor U9537 (N_9537,N_9012,N_9376);
nor U9538 (N_9538,N_9078,N_9194);
and U9539 (N_9539,N_9127,N_9226);
xnor U9540 (N_9540,N_9486,N_9298);
nand U9541 (N_9541,N_9079,N_9446);
nor U9542 (N_9542,N_9414,N_9209);
nand U9543 (N_9543,N_9350,N_9043);
nor U9544 (N_9544,N_9186,N_9457);
and U9545 (N_9545,N_9409,N_9430);
nor U9546 (N_9546,N_9072,N_9048);
nand U9547 (N_9547,N_9420,N_9332);
or U9548 (N_9548,N_9301,N_9290);
xor U9549 (N_9549,N_9469,N_9047);
or U9550 (N_9550,N_9144,N_9070);
nand U9551 (N_9551,N_9218,N_9334);
and U9552 (N_9552,N_9212,N_9431);
nand U9553 (N_9553,N_9271,N_9046);
nand U9554 (N_9554,N_9465,N_9354);
nor U9555 (N_9555,N_9468,N_9237);
and U9556 (N_9556,N_9087,N_9413);
nor U9557 (N_9557,N_9142,N_9461);
nand U9558 (N_9558,N_9187,N_9249);
xnor U9559 (N_9559,N_9027,N_9120);
nor U9560 (N_9560,N_9128,N_9101);
and U9561 (N_9561,N_9395,N_9358);
and U9562 (N_9562,N_9126,N_9174);
and U9563 (N_9563,N_9018,N_9115);
xor U9564 (N_9564,N_9024,N_9400);
xor U9565 (N_9565,N_9317,N_9464);
or U9566 (N_9566,N_9167,N_9470);
and U9567 (N_9567,N_9479,N_9246);
xnor U9568 (N_9568,N_9270,N_9238);
xnor U9569 (N_9569,N_9233,N_9240);
or U9570 (N_9570,N_9119,N_9364);
xnor U9571 (N_9571,N_9145,N_9192);
or U9572 (N_9572,N_9453,N_9227);
xor U9573 (N_9573,N_9399,N_9482);
or U9574 (N_9574,N_9253,N_9092);
and U9575 (N_9575,N_9248,N_9125);
and U9576 (N_9576,N_9397,N_9045);
or U9577 (N_9577,N_9182,N_9321);
or U9578 (N_9578,N_9080,N_9489);
nor U9579 (N_9579,N_9386,N_9438);
nor U9580 (N_9580,N_9037,N_9104);
and U9581 (N_9581,N_9282,N_9493);
nor U9582 (N_9582,N_9342,N_9422);
nor U9583 (N_9583,N_9272,N_9236);
nand U9584 (N_9584,N_9370,N_9208);
and U9585 (N_9585,N_9322,N_9107);
xor U9586 (N_9586,N_9199,N_9143);
nor U9587 (N_9587,N_9352,N_9421);
nand U9588 (N_9588,N_9444,N_9394);
xor U9589 (N_9589,N_9443,N_9418);
xor U9590 (N_9590,N_9179,N_9456);
and U9591 (N_9591,N_9353,N_9007);
nor U9592 (N_9592,N_9472,N_9008);
xnor U9593 (N_9593,N_9427,N_9206);
xnor U9594 (N_9594,N_9138,N_9135);
xnor U9595 (N_9595,N_9279,N_9096);
or U9596 (N_9596,N_9057,N_9228);
nor U9597 (N_9597,N_9349,N_9327);
nor U9598 (N_9598,N_9035,N_9484);
or U9599 (N_9599,N_9146,N_9458);
nor U9600 (N_9600,N_9447,N_9213);
and U9601 (N_9601,N_9028,N_9255);
or U9602 (N_9602,N_9351,N_9082);
or U9603 (N_9603,N_9224,N_9222);
or U9604 (N_9604,N_9040,N_9176);
xnor U9605 (N_9605,N_9266,N_9429);
and U9606 (N_9606,N_9286,N_9445);
nor U9607 (N_9607,N_9097,N_9261);
or U9608 (N_9608,N_9280,N_9437);
or U9609 (N_9609,N_9016,N_9230);
xor U9610 (N_9610,N_9189,N_9181);
nand U9611 (N_9611,N_9066,N_9123);
xnor U9612 (N_9612,N_9110,N_9305);
nor U9613 (N_9613,N_9294,N_9162);
xor U9614 (N_9614,N_9442,N_9056);
xnor U9615 (N_9615,N_9481,N_9393);
nor U9616 (N_9616,N_9487,N_9454);
or U9617 (N_9617,N_9313,N_9398);
xor U9618 (N_9618,N_9118,N_9000);
and U9619 (N_9619,N_9090,N_9339);
nand U9620 (N_9620,N_9297,N_9203);
or U9621 (N_9621,N_9156,N_9075);
xnor U9622 (N_9622,N_9257,N_9221);
or U9623 (N_9623,N_9379,N_9378);
or U9624 (N_9624,N_9498,N_9204);
xor U9625 (N_9625,N_9084,N_9299);
and U9626 (N_9626,N_9241,N_9034);
xor U9627 (N_9627,N_9130,N_9276);
nor U9628 (N_9628,N_9404,N_9094);
nand U9629 (N_9629,N_9361,N_9335);
and U9630 (N_9630,N_9440,N_9490);
nor U9631 (N_9631,N_9244,N_9415);
xor U9632 (N_9632,N_9076,N_9129);
nand U9633 (N_9633,N_9111,N_9089);
nor U9634 (N_9634,N_9149,N_9065);
xor U9635 (N_9635,N_9106,N_9077);
nand U9636 (N_9636,N_9036,N_9256);
nand U9637 (N_9637,N_9153,N_9050);
nor U9638 (N_9638,N_9483,N_9039);
and U9639 (N_9639,N_9348,N_9258);
xor U9640 (N_9640,N_9306,N_9325);
or U9641 (N_9641,N_9160,N_9168);
or U9642 (N_9642,N_9485,N_9239);
xor U9643 (N_9643,N_9121,N_9344);
nand U9644 (N_9644,N_9346,N_9025);
xnor U9645 (N_9645,N_9217,N_9497);
nand U9646 (N_9646,N_9403,N_9439);
xor U9647 (N_9647,N_9289,N_9488);
and U9648 (N_9648,N_9053,N_9434);
nor U9649 (N_9649,N_9231,N_9265);
nor U9650 (N_9650,N_9424,N_9329);
xor U9651 (N_9651,N_9416,N_9330);
and U9652 (N_9652,N_9494,N_9051);
nand U9653 (N_9653,N_9373,N_9191);
or U9654 (N_9654,N_9085,N_9112);
nor U9655 (N_9655,N_9100,N_9463);
or U9656 (N_9656,N_9324,N_9328);
nor U9657 (N_9657,N_9452,N_9363);
and U9658 (N_9658,N_9273,N_9173);
or U9659 (N_9659,N_9172,N_9124);
nor U9660 (N_9660,N_9274,N_9190);
or U9661 (N_9661,N_9071,N_9308);
or U9662 (N_9662,N_9451,N_9433);
xor U9663 (N_9663,N_9260,N_9360);
nand U9664 (N_9664,N_9003,N_9277);
xnor U9665 (N_9665,N_9372,N_9137);
xor U9666 (N_9666,N_9158,N_9357);
nand U9667 (N_9667,N_9380,N_9425);
nor U9668 (N_9668,N_9312,N_9263);
nand U9669 (N_9669,N_9478,N_9052);
and U9670 (N_9670,N_9269,N_9252);
xor U9671 (N_9671,N_9254,N_9098);
or U9672 (N_9672,N_9017,N_9042);
nor U9673 (N_9673,N_9333,N_9281);
nor U9674 (N_9674,N_9108,N_9406);
nor U9675 (N_9675,N_9389,N_9448);
nand U9676 (N_9676,N_9307,N_9165);
nor U9677 (N_9677,N_9450,N_9300);
and U9678 (N_9678,N_9216,N_9058);
nand U9679 (N_9679,N_9030,N_9214);
xor U9680 (N_9680,N_9315,N_9320);
nand U9681 (N_9681,N_9061,N_9475);
nand U9682 (N_9682,N_9054,N_9417);
nor U9683 (N_9683,N_9365,N_9235);
and U9684 (N_9684,N_9411,N_9225);
and U9685 (N_9685,N_9467,N_9345);
or U9686 (N_9686,N_9063,N_9331);
nand U9687 (N_9687,N_9081,N_9031);
nor U9688 (N_9688,N_9006,N_9362);
xnor U9689 (N_9689,N_9041,N_9476);
or U9690 (N_9690,N_9390,N_9229);
and U9691 (N_9691,N_9278,N_9496);
nand U9692 (N_9692,N_9033,N_9243);
and U9693 (N_9693,N_9152,N_9426);
nor U9694 (N_9694,N_9436,N_9267);
and U9695 (N_9695,N_9292,N_9432);
and U9696 (N_9696,N_9009,N_9184);
xor U9697 (N_9697,N_9060,N_9287);
xor U9698 (N_9698,N_9401,N_9388);
xnor U9699 (N_9699,N_9131,N_9091);
and U9700 (N_9700,N_9026,N_9410);
and U9701 (N_9701,N_9180,N_9460);
xor U9702 (N_9702,N_9264,N_9169);
xnor U9703 (N_9703,N_9285,N_9326);
or U9704 (N_9704,N_9211,N_9371);
nor U9705 (N_9705,N_9338,N_9148);
nand U9706 (N_9706,N_9268,N_9259);
nor U9707 (N_9707,N_9064,N_9215);
xor U9708 (N_9708,N_9377,N_9369);
nor U9709 (N_9709,N_9175,N_9441);
and U9710 (N_9710,N_9004,N_9375);
and U9711 (N_9711,N_9408,N_9423);
nor U9712 (N_9712,N_9014,N_9355);
nand U9713 (N_9713,N_9251,N_9310);
nand U9714 (N_9714,N_9010,N_9069);
xor U9715 (N_9715,N_9337,N_9262);
and U9716 (N_9716,N_9117,N_9405);
and U9717 (N_9717,N_9381,N_9304);
or U9718 (N_9718,N_9099,N_9391);
or U9719 (N_9719,N_9303,N_9316);
nor U9720 (N_9720,N_9311,N_9247);
nand U9721 (N_9721,N_9020,N_9318);
nor U9722 (N_9722,N_9105,N_9499);
and U9723 (N_9723,N_9385,N_9340);
nor U9724 (N_9724,N_9197,N_9157);
or U9725 (N_9725,N_9284,N_9474);
or U9726 (N_9726,N_9055,N_9139);
xor U9727 (N_9727,N_9032,N_9178);
and U9728 (N_9728,N_9062,N_9232);
or U9729 (N_9729,N_9133,N_9200);
and U9730 (N_9730,N_9049,N_9314);
or U9731 (N_9731,N_9336,N_9396);
and U9732 (N_9732,N_9001,N_9387);
nand U9733 (N_9733,N_9210,N_9466);
xor U9734 (N_9734,N_9171,N_9170);
and U9735 (N_9735,N_9288,N_9275);
and U9736 (N_9736,N_9480,N_9177);
xnor U9737 (N_9737,N_9073,N_9295);
xnor U9738 (N_9738,N_9109,N_9202);
xnor U9739 (N_9739,N_9166,N_9491);
or U9740 (N_9740,N_9044,N_9302);
or U9741 (N_9741,N_9116,N_9005);
and U9742 (N_9742,N_9220,N_9023);
nor U9743 (N_9743,N_9095,N_9159);
nand U9744 (N_9744,N_9195,N_9013);
nand U9745 (N_9745,N_9141,N_9102);
nor U9746 (N_9746,N_9323,N_9250);
and U9747 (N_9747,N_9147,N_9132);
xnor U9748 (N_9748,N_9343,N_9114);
or U9749 (N_9749,N_9205,N_9198);
nand U9750 (N_9750,N_9245,N_9312);
nand U9751 (N_9751,N_9323,N_9056);
and U9752 (N_9752,N_9441,N_9310);
nand U9753 (N_9753,N_9047,N_9454);
nor U9754 (N_9754,N_9412,N_9119);
xnor U9755 (N_9755,N_9480,N_9353);
and U9756 (N_9756,N_9331,N_9474);
or U9757 (N_9757,N_9143,N_9347);
nand U9758 (N_9758,N_9168,N_9006);
or U9759 (N_9759,N_9119,N_9018);
nor U9760 (N_9760,N_9300,N_9031);
nor U9761 (N_9761,N_9138,N_9112);
xor U9762 (N_9762,N_9002,N_9421);
and U9763 (N_9763,N_9388,N_9072);
and U9764 (N_9764,N_9447,N_9211);
nor U9765 (N_9765,N_9342,N_9202);
nor U9766 (N_9766,N_9302,N_9258);
nand U9767 (N_9767,N_9434,N_9478);
and U9768 (N_9768,N_9229,N_9470);
or U9769 (N_9769,N_9081,N_9308);
xnor U9770 (N_9770,N_9241,N_9011);
and U9771 (N_9771,N_9088,N_9131);
nor U9772 (N_9772,N_9239,N_9086);
and U9773 (N_9773,N_9090,N_9213);
xor U9774 (N_9774,N_9255,N_9257);
xor U9775 (N_9775,N_9413,N_9055);
nor U9776 (N_9776,N_9457,N_9142);
nand U9777 (N_9777,N_9165,N_9387);
and U9778 (N_9778,N_9287,N_9122);
and U9779 (N_9779,N_9237,N_9212);
or U9780 (N_9780,N_9307,N_9274);
nor U9781 (N_9781,N_9463,N_9019);
or U9782 (N_9782,N_9289,N_9261);
nand U9783 (N_9783,N_9465,N_9444);
xor U9784 (N_9784,N_9390,N_9337);
or U9785 (N_9785,N_9454,N_9173);
and U9786 (N_9786,N_9075,N_9037);
xor U9787 (N_9787,N_9282,N_9071);
and U9788 (N_9788,N_9440,N_9080);
or U9789 (N_9789,N_9287,N_9423);
nand U9790 (N_9790,N_9269,N_9141);
and U9791 (N_9791,N_9109,N_9196);
or U9792 (N_9792,N_9165,N_9390);
and U9793 (N_9793,N_9031,N_9087);
and U9794 (N_9794,N_9418,N_9024);
nor U9795 (N_9795,N_9393,N_9198);
xor U9796 (N_9796,N_9426,N_9206);
nor U9797 (N_9797,N_9359,N_9005);
or U9798 (N_9798,N_9084,N_9376);
or U9799 (N_9799,N_9126,N_9200);
xnor U9800 (N_9800,N_9469,N_9021);
or U9801 (N_9801,N_9362,N_9375);
xnor U9802 (N_9802,N_9154,N_9096);
or U9803 (N_9803,N_9152,N_9325);
and U9804 (N_9804,N_9318,N_9098);
and U9805 (N_9805,N_9239,N_9272);
xor U9806 (N_9806,N_9467,N_9196);
nor U9807 (N_9807,N_9264,N_9286);
nand U9808 (N_9808,N_9129,N_9237);
or U9809 (N_9809,N_9362,N_9067);
or U9810 (N_9810,N_9406,N_9459);
nor U9811 (N_9811,N_9290,N_9332);
xor U9812 (N_9812,N_9346,N_9055);
and U9813 (N_9813,N_9235,N_9408);
and U9814 (N_9814,N_9287,N_9229);
xnor U9815 (N_9815,N_9220,N_9033);
or U9816 (N_9816,N_9487,N_9442);
or U9817 (N_9817,N_9393,N_9243);
nand U9818 (N_9818,N_9063,N_9198);
xor U9819 (N_9819,N_9222,N_9212);
or U9820 (N_9820,N_9057,N_9035);
nand U9821 (N_9821,N_9254,N_9388);
xnor U9822 (N_9822,N_9307,N_9083);
or U9823 (N_9823,N_9420,N_9296);
nand U9824 (N_9824,N_9026,N_9207);
nand U9825 (N_9825,N_9238,N_9142);
nor U9826 (N_9826,N_9382,N_9187);
or U9827 (N_9827,N_9477,N_9420);
xor U9828 (N_9828,N_9209,N_9420);
xor U9829 (N_9829,N_9313,N_9036);
nor U9830 (N_9830,N_9487,N_9450);
nor U9831 (N_9831,N_9025,N_9409);
xnor U9832 (N_9832,N_9385,N_9370);
nand U9833 (N_9833,N_9164,N_9174);
or U9834 (N_9834,N_9441,N_9297);
nand U9835 (N_9835,N_9180,N_9165);
nor U9836 (N_9836,N_9350,N_9483);
nor U9837 (N_9837,N_9249,N_9453);
or U9838 (N_9838,N_9381,N_9017);
nor U9839 (N_9839,N_9002,N_9217);
and U9840 (N_9840,N_9117,N_9385);
nand U9841 (N_9841,N_9325,N_9298);
nand U9842 (N_9842,N_9265,N_9390);
nor U9843 (N_9843,N_9217,N_9411);
and U9844 (N_9844,N_9483,N_9231);
xnor U9845 (N_9845,N_9222,N_9281);
and U9846 (N_9846,N_9108,N_9471);
or U9847 (N_9847,N_9125,N_9265);
and U9848 (N_9848,N_9058,N_9375);
nor U9849 (N_9849,N_9313,N_9401);
xnor U9850 (N_9850,N_9060,N_9036);
xor U9851 (N_9851,N_9470,N_9087);
and U9852 (N_9852,N_9468,N_9476);
xnor U9853 (N_9853,N_9389,N_9273);
nor U9854 (N_9854,N_9094,N_9348);
xnor U9855 (N_9855,N_9367,N_9067);
nand U9856 (N_9856,N_9498,N_9262);
xor U9857 (N_9857,N_9287,N_9432);
nor U9858 (N_9858,N_9321,N_9411);
nand U9859 (N_9859,N_9122,N_9181);
xor U9860 (N_9860,N_9159,N_9228);
xor U9861 (N_9861,N_9443,N_9456);
and U9862 (N_9862,N_9495,N_9119);
nand U9863 (N_9863,N_9407,N_9004);
nand U9864 (N_9864,N_9035,N_9024);
nor U9865 (N_9865,N_9320,N_9349);
and U9866 (N_9866,N_9359,N_9037);
xor U9867 (N_9867,N_9139,N_9173);
and U9868 (N_9868,N_9196,N_9263);
nand U9869 (N_9869,N_9070,N_9474);
and U9870 (N_9870,N_9050,N_9462);
nor U9871 (N_9871,N_9162,N_9207);
nor U9872 (N_9872,N_9182,N_9056);
xnor U9873 (N_9873,N_9371,N_9299);
or U9874 (N_9874,N_9305,N_9083);
nor U9875 (N_9875,N_9361,N_9067);
and U9876 (N_9876,N_9230,N_9272);
nand U9877 (N_9877,N_9167,N_9481);
or U9878 (N_9878,N_9314,N_9375);
or U9879 (N_9879,N_9013,N_9319);
nor U9880 (N_9880,N_9273,N_9149);
or U9881 (N_9881,N_9259,N_9091);
nand U9882 (N_9882,N_9215,N_9383);
nor U9883 (N_9883,N_9240,N_9369);
nor U9884 (N_9884,N_9242,N_9148);
or U9885 (N_9885,N_9130,N_9488);
and U9886 (N_9886,N_9483,N_9102);
or U9887 (N_9887,N_9390,N_9445);
and U9888 (N_9888,N_9135,N_9054);
nand U9889 (N_9889,N_9406,N_9444);
nand U9890 (N_9890,N_9133,N_9215);
nand U9891 (N_9891,N_9371,N_9100);
nand U9892 (N_9892,N_9034,N_9100);
xnor U9893 (N_9893,N_9221,N_9238);
xor U9894 (N_9894,N_9454,N_9470);
nand U9895 (N_9895,N_9482,N_9023);
nand U9896 (N_9896,N_9451,N_9396);
and U9897 (N_9897,N_9175,N_9116);
or U9898 (N_9898,N_9290,N_9083);
and U9899 (N_9899,N_9421,N_9310);
xor U9900 (N_9900,N_9041,N_9365);
nand U9901 (N_9901,N_9453,N_9283);
nor U9902 (N_9902,N_9038,N_9368);
or U9903 (N_9903,N_9063,N_9050);
and U9904 (N_9904,N_9098,N_9019);
xor U9905 (N_9905,N_9056,N_9259);
and U9906 (N_9906,N_9440,N_9448);
or U9907 (N_9907,N_9378,N_9073);
or U9908 (N_9908,N_9039,N_9339);
xor U9909 (N_9909,N_9256,N_9146);
nand U9910 (N_9910,N_9216,N_9425);
nand U9911 (N_9911,N_9357,N_9356);
or U9912 (N_9912,N_9496,N_9384);
nor U9913 (N_9913,N_9116,N_9115);
nor U9914 (N_9914,N_9220,N_9107);
xor U9915 (N_9915,N_9324,N_9304);
or U9916 (N_9916,N_9010,N_9386);
and U9917 (N_9917,N_9381,N_9021);
nand U9918 (N_9918,N_9465,N_9249);
xnor U9919 (N_9919,N_9422,N_9443);
nor U9920 (N_9920,N_9021,N_9426);
and U9921 (N_9921,N_9099,N_9423);
nor U9922 (N_9922,N_9121,N_9251);
nor U9923 (N_9923,N_9444,N_9146);
nand U9924 (N_9924,N_9418,N_9405);
nor U9925 (N_9925,N_9358,N_9448);
and U9926 (N_9926,N_9199,N_9279);
nor U9927 (N_9927,N_9016,N_9245);
xnor U9928 (N_9928,N_9362,N_9127);
xor U9929 (N_9929,N_9209,N_9155);
nor U9930 (N_9930,N_9385,N_9278);
and U9931 (N_9931,N_9289,N_9105);
or U9932 (N_9932,N_9464,N_9013);
and U9933 (N_9933,N_9140,N_9411);
or U9934 (N_9934,N_9022,N_9005);
nor U9935 (N_9935,N_9160,N_9385);
and U9936 (N_9936,N_9082,N_9295);
nor U9937 (N_9937,N_9334,N_9289);
xor U9938 (N_9938,N_9318,N_9301);
xnor U9939 (N_9939,N_9093,N_9027);
nand U9940 (N_9940,N_9165,N_9371);
nor U9941 (N_9941,N_9160,N_9460);
nand U9942 (N_9942,N_9373,N_9398);
nor U9943 (N_9943,N_9471,N_9416);
xor U9944 (N_9944,N_9313,N_9470);
nor U9945 (N_9945,N_9446,N_9231);
and U9946 (N_9946,N_9113,N_9140);
nor U9947 (N_9947,N_9356,N_9159);
xnor U9948 (N_9948,N_9226,N_9144);
nand U9949 (N_9949,N_9106,N_9004);
and U9950 (N_9950,N_9319,N_9374);
nor U9951 (N_9951,N_9440,N_9350);
or U9952 (N_9952,N_9239,N_9479);
nor U9953 (N_9953,N_9301,N_9355);
xnor U9954 (N_9954,N_9086,N_9141);
or U9955 (N_9955,N_9444,N_9483);
nand U9956 (N_9956,N_9173,N_9195);
nand U9957 (N_9957,N_9497,N_9373);
and U9958 (N_9958,N_9039,N_9092);
or U9959 (N_9959,N_9443,N_9032);
xnor U9960 (N_9960,N_9311,N_9054);
nand U9961 (N_9961,N_9247,N_9099);
xnor U9962 (N_9962,N_9253,N_9386);
nor U9963 (N_9963,N_9409,N_9165);
xnor U9964 (N_9964,N_9328,N_9374);
xnor U9965 (N_9965,N_9149,N_9016);
and U9966 (N_9966,N_9260,N_9499);
xnor U9967 (N_9967,N_9173,N_9375);
nand U9968 (N_9968,N_9257,N_9116);
xor U9969 (N_9969,N_9215,N_9123);
nor U9970 (N_9970,N_9254,N_9284);
nand U9971 (N_9971,N_9092,N_9376);
xor U9972 (N_9972,N_9278,N_9472);
or U9973 (N_9973,N_9444,N_9110);
and U9974 (N_9974,N_9285,N_9136);
nor U9975 (N_9975,N_9242,N_9061);
nor U9976 (N_9976,N_9264,N_9426);
and U9977 (N_9977,N_9386,N_9162);
xnor U9978 (N_9978,N_9058,N_9321);
and U9979 (N_9979,N_9107,N_9380);
nor U9980 (N_9980,N_9081,N_9337);
xnor U9981 (N_9981,N_9041,N_9426);
xnor U9982 (N_9982,N_9158,N_9348);
nor U9983 (N_9983,N_9319,N_9449);
or U9984 (N_9984,N_9045,N_9095);
and U9985 (N_9985,N_9390,N_9252);
or U9986 (N_9986,N_9126,N_9453);
xnor U9987 (N_9987,N_9279,N_9200);
nand U9988 (N_9988,N_9007,N_9343);
and U9989 (N_9989,N_9022,N_9409);
nor U9990 (N_9990,N_9256,N_9125);
xor U9991 (N_9991,N_9245,N_9366);
or U9992 (N_9992,N_9364,N_9492);
xor U9993 (N_9993,N_9150,N_9232);
nor U9994 (N_9994,N_9176,N_9296);
nor U9995 (N_9995,N_9363,N_9167);
nor U9996 (N_9996,N_9347,N_9052);
nand U9997 (N_9997,N_9471,N_9006);
nor U9998 (N_9998,N_9273,N_9201);
nor U9999 (N_9999,N_9210,N_9040);
xnor U10000 (N_10000,N_9551,N_9542);
or U10001 (N_10001,N_9722,N_9867);
or U10002 (N_10002,N_9794,N_9849);
xnor U10003 (N_10003,N_9653,N_9847);
nand U10004 (N_10004,N_9672,N_9550);
and U10005 (N_10005,N_9796,N_9891);
nand U10006 (N_10006,N_9533,N_9670);
xnor U10007 (N_10007,N_9868,N_9636);
or U10008 (N_10008,N_9797,N_9887);
nand U10009 (N_10009,N_9940,N_9615);
nand U10010 (N_10010,N_9709,N_9906);
nand U10011 (N_10011,N_9682,N_9634);
and U10012 (N_10012,N_9597,N_9714);
and U10013 (N_10013,N_9534,N_9875);
nor U10014 (N_10014,N_9541,N_9734);
or U10015 (N_10015,N_9503,N_9640);
nor U10016 (N_10016,N_9969,N_9739);
or U10017 (N_10017,N_9590,N_9989);
and U10018 (N_10018,N_9942,N_9724);
and U10019 (N_10019,N_9961,N_9567);
nor U10020 (N_10020,N_9740,N_9654);
nor U10021 (N_10021,N_9931,N_9744);
nand U10022 (N_10022,N_9823,N_9512);
nor U10023 (N_10023,N_9517,N_9878);
or U10024 (N_10024,N_9807,N_9844);
nand U10025 (N_10025,N_9516,N_9647);
nor U10026 (N_10026,N_9960,N_9816);
nand U10027 (N_10027,N_9588,N_9988);
nand U10028 (N_10028,N_9918,N_9933);
or U10029 (N_10029,N_9776,N_9997);
and U10030 (N_10030,N_9531,N_9999);
or U10031 (N_10031,N_9589,N_9558);
nor U10032 (N_10032,N_9635,N_9628);
xnor U10033 (N_10033,N_9718,N_9922);
and U10034 (N_10034,N_9610,N_9620);
or U10035 (N_10035,N_9958,N_9553);
nor U10036 (N_10036,N_9957,N_9659);
and U10037 (N_10037,N_9658,N_9519);
xor U10038 (N_10038,N_9853,N_9943);
nand U10039 (N_10039,N_9841,N_9914);
nand U10040 (N_10040,N_9748,N_9814);
nor U10041 (N_10041,N_9556,N_9566);
or U10042 (N_10042,N_9532,N_9982);
xnor U10043 (N_10043,N_9683,N_9890);
nand U10044 (N_10044,N_9905,N_9782);
nor U10045 (N_10045,N_9954,N_9858);
xnor U10046 (N_10046,N_9546,N_9848);
nand U10047 (N_10047,N_9562,N_9623);
nor U10048 (N_10048,N_9660,N_9761);
nor U10049 (N_10049,N_9843,N_9935);
or U10050 (N_10050,N_9694,N_9774);
and U10051 (N_10051,N_9622,N_9900);
nor U10052 (N_10052,N_9831,N_9547);
and U10053 (N_10053,N_9921,N_9926);
nor U10054 (N_10054,N_9674,N_9864);
nor U10055 (N_10055,N_9974,N_9779);
xnor U10056 (N_10056,N_9731,N_9990);
or U10057 (N_10057,N_9736,N_9504);
or U10058 (N_10058,N_9786,N_9563);
xnor U10059 (N_10059,N_9979,N_9869);
nor U10060 (N_10060,N_9633,N_9520);
xnor U10061 (N_10061,N_9632,N_9850);
xor U10062 (N_10062,N_9746,N_9627);
nand U10063 (N_10063,N_9525,N_9759);
or U10064 (N_10064,N_9577,N_9642);
or U10065 (N_10065,N_9506,N_9644);
and U10066 (N_10066,N_9830,N_9631);
xor U10067 (N_10067,N_9515,N_9664);
xnor U10068 (N_10068,N_9639,N_9679);
nor U10069 (N_10069,N_9675,N_9928);
xnor U10070 (N_10070,N_9536,N_9707);
nand U10071 (N_10071,N_9950,N_9981);
xor U10072 (N_10072,N_9603,N_9760);
and U10073 (N_10073,N_9938,N_9629);
and U10074 (N_10074,N_9650,N_9576);
or U10075 (N_10075,N_9993,N_9715);
xnor U10076 (N_10076,N_9835,N_9909);
nand U10077 (N_10077,N_9646,N_9575);
and U10078 (N_10078,N_9792,N_9966);
nand U10079 (N_10079,N_9641,N_9977);
nand U10080 (N_10080,N_9671,N_9535);
or U10081 (N_10081,N_9946,N_9877);
xnor U10082 (N_10082,N_9862,N_9888);
or U10083 (N_10083,N_9784,N_9666);
and U10084 (N_10084,N_9619,N_9651);
and U10085 (N_10085,N_9685,N_9713);
and U10086 (N_10086,N_9721,N_9555);
or U10087 (N_10087,N_9611,N_9897);
or U10088 (N_10088,N_9699,N_9587);
or U10089 (N_10089,N_9825,N_9729);
xor U10090 (N_10090,N_9805,N_9524);
or U10091 (N_10091,N_9757,N_9751);
or U10092 (N_10092,N_9703,N_9840);
xnor U10093 (N_10093,N_9581,N_9898);
nand U10094 (N_10094,N_9693,N_9560);
xnor U10095 (N_10095,N_9873,N_9578);
nand U10096 (N_10096,N_9872,N_9601);
nand U10097 (N_10097,N_9809,N_9965);
nor U10098 (N_10098,N_9608,N_9501);
nand U10099 (N_10099,N_9596,N_9708);
nor U10100 (N_10100,N_9885,N_9625);
nand U10101 (N_10101,N_9763,N_9549);
xnor U10102 (N_10102,N_9681,N_9829);
nor U10103 (N_10103,N_9984,N_9598);
nor U10104 (N_10104,N_9783,N_9767);
nor U10105 (N_10105,N_9604,N_9662);
nor U10106 (N_10106,N_9643,N_9856);
or U10107 (N_10107,N_9554,N_9720);
or U10108 (N_10108,N_9698,N_9834);
or U10109 (N_10109,N_9656,N_9808);
and U10110 (N_10110,N_9655,N_9665);
and U10111 (N_10111,N_9947,N_9725);
nand U10112 (N_10112,N_9710,N_9595);
nor U10113 (N_10113,N_9768,N_9913);
or U10114 (N_10114,N_9880,N_9539);
nand U10115 (N_10115,N_9815,N_9978);
and U10116 (N_10116,N_9540,N_9932);
or U10117 (N_10117,N_9518,N_9738);
nor U10118 (N_10118,N_9543,N_9996);
xnor U10119 (N_10119,N_9669,N_9509);
or U10120 (N_10120,N_9801,N_9855);
nand U10121 (N_10121,N_9579,N_9700);
xor U10122 (N_10122,N_9712,N_9583);
or U10123 (N_10123,N_9523,N_9530);
and U10124 (N_10124,N_9663,N_9874);
and U10125 (N_10125,N_9991,N_9980);
and U10126 (N_10126,N_9584,N_9800);
nor U10127 (N_10127,N_9649,N_9648);
nor U10128 (N_10128,N_9741,N_9507);
nand U10129 (N_10129,N_9750,N_9600);
and U10130 (N_10130,N_9591,N_9626);
xnor U10131 (N_10131,N_9522,N_9930);
nand U10132 (N_10132,N_9705,N_9500);
and U10133 (N_10133,N_9785,N_9852);
and U10134 (N_10134,N_9559,N_9617);
nor U10135 (N_10135,N_9962,N_9820);
and U10136 (N_10136,N_9948,N_9616);
or U10137 (N_10137,N_9521,N_9565);
nor U10138 (N_10138,N_9903,N_9895);
nor U10139 (N_10139,N_9599,N_9902);
nor U10140 (N_10140,N_9812,N_9676);
nand U10141 (N_10141,N_9952,N_9788);
xor U10142 (N_10142,N_9992,N_9689);
nor U10143 (N_10143,N_9845,N_9661);
and U10144 (N_10144,N_9630,N_9780);
or U10145 (N_10145,N_9688,N_9667);
or U10146 (N_10146,N_9963,N_9842);
or U10147 (N_10147,N_9837,N_9822);
nand U10148 (N_10148,N_9939,N_9621);
and U10149 (N_10149,N_9929,N_9983);
or U10150 (N_10150,N_9538,N_9614);
xor U10151 (N_10151,N_9706,N_9870);
xnor U10152 (N_10152,N_9505,N_9719);
or U10153 (N_10153,N_9508,N_9793);
and U10154 (N_10154,N_9702,N_9866);
and U10155 (N_10155,N_9791,N_9955);
or U10156 (N_10156,N_9771,N_9762);
and U10157 (N_10157,N_9959,N_9605);
xnor U10158 (N_10158,N_9799,N_9998);
or U10159 (N_10159,N_9936,N_9573);
and U10160 (N_10160,N_9502,N_9585);
and U10161 (N_10161,N_9732,N_9528);
and U10162 (N_10162,N_9586,N_9692);
nand U10163 (N_10163,N_9735,N_9968);
and U10164 (N_10164,N_9697,N_9896);
and U10165 (N_10165,N_9691,N_9684);
or U10166 (N_10166,N_9987,N_9937);
or U10167 (N_10167,N_9851,N_9907);
xnor U10168 (N_10168,N_9910,N_9510);
or U10169 (N_10169,N_9678,N_9986);
nor U10170 (N_10170,N_9695,N_9832);
nor U10171 (N_10171,N_9892,N_9690);
nand U10172 (N_10172,N_9728,N_9711);
and U10173 (N_10173,N_9821,N_9737);
and U10174 (N_10174,N_9917,N_9884);
nand U10175 (N_10175,N_9687,N_9733);
and U10176 (N_10176,N_9777,N_9863);
or U10177 (N_10177,N_9752,N_9609);
nand U10178 (N_10178,N_9657,N_9527);
or U10179 (N_10179,N_9985,N_9912);
nor U10180 (N_10180,N_9593,N_9971);
and U10181 (N_10181,N_9747,N_9606);
nand U10182 (N_10182,N_9861,N_9839);
nand U10183 (N_10183,N_9607,N_9511);
nor U10184 (N_10184,N_9871,N_9704);
nor U10185 (N_10185,N_9972,N_9795);
xnor U10186 (N_10186,N_9544,N_9745);
or U10187 (N_10187,N_9513,N_9904);
xor U10188 (N_10188,N_9727,N_9781);
and U10189 (N_10189,N_9548,N_9602);
or U10190 (N_10190,N_9717,N_9810);
nor U10191 (N_10191,N_9743,N_9876);
xnor U10192 (N_10192,N_9953,N_9561);
nor U10193 (N_10193,N_9537,N_9557);
nor U10194 (N_10194,N_9865,N_9753);
and U10195 (N_10195,N_9755,N_9967);
and U10196 (N_10196,N_9749,N_9970);
nand U10197 (N_10197,N_9854,N_9883);
and U10198 (N_10198,N_9723,N_9945);
xor U10199 (N_10199,N_9764,N_9770);
or U10200 (N_10200,N_9618,N_9696);
nor U10201 (N_10201,N_9819,N_9817);
or U10202 (N_10202,N_9826,N_9846);
and U10203 (N_10203,N_9552,N_9828);
xor U10204 (N_10204,N_9592,N_9824);
and U10205 (N_10205,N_9949,N_9803);
and U10206 (N_10206,N_9827,N_9879);
nand U10207 (N_10207,N_9574,N_9833);
xor U10208 (N_10208,N_9677,N_9899);
and U10209 (N_10209,N_9911,N_9778);
and U10210 (N_10210,N_9668,N_9923);
and U10211 (N_10211,N_9994,N_9813);
xor U10212 (N_10212,N_9886,N_9754);
or U10213 (N_10213,N_9951,N_9927);
nor U10214 (N_10214,N_9730,N_9529);
nor U10215 (N_10215,N_9857,N_9580);
nor U10216 (N_10216,N_9775,N_9765);
nor U10217 (N_10217,N_9901,N_9859);
xnor U10218 (N_10218,N_9758,N_9756);
nand U10219 (N_10219,N_9836,N_9956);
nor U10220 (N_10220,N_9818,N_9772);
and U10221 (N_10221,N_9790,N_9882);
nand U10222 (N_10222,N_9915,N_9716);
xnor U10223 (N_10223,N_9838,N_9806);
nand U10224 (N_10224,N_9637,N_9624);
nor U10225 (N_10225,N_9995,N_9908);
nor U10226 (N_10226,N_9545,N_9594);
xnor U10227 (N_10227,N_9894,N_9571);
xnor U10228 (N_10228,N_9798,N_9638);
nor U10229 (N_10229,N_9811,N_9572);
xnor U10230 (N_10230,N_9564,N_9773);
nand U10231 (N_10231,N_9769,N_9934);
nand U10232 (N_10232,N_9613,N_9680);
or U10233 (N_10233,N_9612,N_9570);
nand U10234 (N_10234,N_9686,N_9973);
or U10235 (N_10235,N_9976,N_9652);
and U10236 (N_10236,N_9893,N_9787);
and U10237 (N_10237,N_9860,N_9919);
or U10238 (N_10238,N_9645,N_9802);
and U10239 (N_10239,N_9568,N_9964);
and U10240 (N_10240,N_9766,N_9881);
and U10241 (N_10241,N_9916,N_9673);
nand U10242 (N_10242,N_9569,N_9514);
or U10243 (N_10243,N_9889,N_9742);
xor U10244 (N_10244,N_9944,N_9526);
nand U10245 (N_10245,N_9804,N_9726);
xnor U10246 (N_10246,N_9924,N_9789);
nor U10247 (N_10247,N_9701,N_9925);
nor U10248 (N_10248,N_9941,N_9920);
and U10249 (N_10249,N_9975,N_9582);
xor U10250 (N_10250,N_9942,N_9956);
xor U10251 (N_10251,N_9894,N_9973);
or U10252 (N_10252,N_9708,N_9773);
or U10253 (N_10253,N_9730,N_9873);
and U10254 (N_10254,N_9805,N_9675);
and U10255 (N_10255,N_9979,N_9884);
nand U10256 (N_10256,N_9668,N_9658);
xnor U10257 (N_10257,N_9686,N_9810);
nand U10258 (N_10258,N_9994,N_9664);
nor U10259 (N_10259,N_9857,N_9703);
xor U10260 (N_10260,N_9933,N_9919);
xnor U10261 (N_10261,N_9557,N_9944);
nor U10262 (N_10262,N_9867,N_9740);
or U10263 (N_10263,N_9999,N_9777);
nor U10264 (N_10264,N_9994,N_9766);
and U10265 (N_10265,N_9813,N_9662);
nor U10266 (N_10266,N_9758,N_9610);
nand U10267 (N_10267,N_9806,N_9975);
and U10268 (N_10268,N_9903,N_9681);
nor U10269 (N_10269,N_9764,N_9665);
nor U10270 (N_10270,N_9704,N_9952);
or U10271 (N_10271,N_9903,N_9686);
xor U10272 (N_10272,N_9934,N_9645);
and U10273 (N_10273,N_9698,N_9556);
nor U10274 (N_10274,N_9570,N_9987);
xor U10275 (N_10275,N_9988,N_9775);
or U10276 (N_10276,N_9911,N_9510);
nor U10277 (N_10277,N_9809,N_9945);
nand U10278 (N_10278,N_9712,N_9762);
nand U10279 (N_10279,N_9938,N_9593);
or U10280 (N_10280,N_9527,N_9683);
xnor U10281 (N_10281,N_9880,N_9588);
and U10282 (N_10282,N_9806,N_9872);
and U10283 (N_10283,N_9724,N_9612);
or U10284 (N_10284,N_9864,N_9751);
xor U10285 (N_10285,N_9931,N_9669);
xnor U10286 (N_10286,N_9603,N_9628);
and U10287 (N_10287,N_9634,N_9937);
nor U10288 (N_10288,N_9645,N_9783);
and U10289 (N_10289,N_9923,N_9740);
or U10290 (N_10290,N_9558,N_9762);
and U10291 (N_10291,N_9628,N_9681);
nor U10292 (N_10292,N_9582,N_9597);
nor U10293 (N_10293,N_9761,N_9607);
or U10294 (N_10294,N_9539,N_9936);
nand U10295 (N_10295,N_9956,N_9642);
nor U10296 (N_10296,N_9736,N_9541);
or U10297 (N_10297,N_9865,N_9666);
and U10298 (N_10298,N_9627,N_9831);
or U10299 (N_10299,N_9577,N_9566);
or U10300 (N_10300,N_9968,N_9552);
or U10301 (N_10301,N_9546,N_9719);
and U10302 (N_10302,N_9623,N_9593);
and U10303 (N_10303,N_9886,N_9692);
xor U10304 (N_10304,N_9867,N_9654);
xnor U10305 (N_10305,N_9728,N_9779);
or U10306 (N_10306,N_9807,N_9923);
nand U10307 (N_10307,N_9885,N_9933);
xor U10308 (N_10308,N_9645,N_9952);
xor U10309 (N_10309,N_9764,N_9619);
and U10310 (N_10310,N_9514,N_9560);
and U10311 (N_10311,N_9738,N_9540);
nand U10312 (N_10312,N_9729,N_9772);
nand U10313 (N_10313,N_9811,N_9635);
or U10314 (N_10314,N_9669,N_9757);
or U10315 (N_10315,N_9541,N_9500);
or U10316 (N_10316,N_9872,N_9987);
nor U10317 (N_10317,N_9716,N_9681);
nor U10318 (N_10318,N_9617,N_9698);
nor U10319 (N_10319,N_9892,N_9514);
or U10320 (N_10320,N_9574,N_9784);
xnor U10321 (N_10321,N_9986,N_9711);
nor U10322 (N_10322,N_9687,N_9737);
and U10323 (N_10323,N_9752,N_9531);
or U10324 (N_10324,N_9596,N_9667);
nor U10325 (N_10325,N_9664,N_9542);
nand U10326 (N_10326,N_9751,N_9679);
and U10327 (N_10327,N_9737,N_9894);
nor U10328 (N_10328,N_9993,N_9908);
or U10329 (N_10329,N_9794,N_9579);
and U10330 (N_10330,N_9894,N_9721);
xnor U10331 (N_10331,N_9854,N_9836);
nand U10332 (N_10332,N_9992,N_9866);
and U10333 (N_10333,N_9762,N_9714);
or U10334 (N_10334,N_9802,N_9839);
nor U10335 (N_10335,N_9565,N_9933);
nand U10336 (N_10336,N_9935,N_9974);
nand U10337 (N_10337,N_9790,N_9562);
or U10338 (N_10338,N_9616,N_9981);
nand U10339 (N_10339,N_9718,N_9532);
and U10340 (N_10340,N_9994,N_9819);
xnor U10341 (N_10341,N_9922,N_9684);
or U10342 (N_10342,N_9538,N_9580);
and U10343 (N_10343,N_9653,N_9681);
or U10344 (N_10344,N_9763,N_9918);
nand U10345 (N_10345,N_9754,N_9801);
or U10346 (N_10346,N_9767,N_9744);
or U10347 (N_10347,N_9508,N_9545);
nor U10348 (N_10348,N_9759,N_9658);
nand U10349 (N_10349,N_9674,N_9623);
nor U10350 (N_10350,N_9685,N_9936);
and U10351 (N_10351,N_9649,N_9556);
nand U10352 (N_10352,N_9741,N_9871);
nand U10353 (N_10353,N_9598,N_9507);
or U10354 (N_10354,N_9862,N_9744);
nand U10355 (N_10355,N_9886,N_9793);
nor U10356 (N_10356,N_9770,N_9696);
xnor U10357 (N_10357,N_9670,N_9654);
and U10358 (N_10358,N_9839,N_9590);
xor U10359 (N_10359,N_9690,N_9739);
and U10360 (N_10360,N_9723,N_9897);
nor U10361 (N_10361,N_9523,N_9844);
or U10362 (N_10362,N_9507,N_9995);
nand U10363 (N_10363,N_9687,N_9501);
and U10364 (N_10364,N_9531,N_9699);
nor U10365 (N_10365,N_9771,N_9774);
and U10366 (N_10366,N_9850,N_9530);
or U10367 (N_10367,N_9965,N_9854);
and U10368 (N_10368,N_9746,N_9668);
and U10369 (N_10369,N_9504,N_9985);
and U10370 (N_10370,N_9788,N_9523);
xnor U10371 (N_10371,N_9840,N_9924);
and U10372 (N_10372,N_9674,N_9586);
xor U10373 (N_10373,N_9944,N_9741);
or U10374 (N_10374,N_9872,N_9620);
xnor U10375 (N_10375,N_9785,N_9861);
or U10376 (N_10376,N_9552,N_9853);
nor U10377 (N_10377,N_9732,N_9515);
nor U10378 (N_10378,N_9949,N_9810);
nor U10379 (N_10379,N_9805,N_9988);
and U10380 (N_10380,N_9685,N_9602);
nand U10381 (N_10381,N_9604,N_9777);
xor U10382 (N_10382,N_9881,N_9618);
and U10383 (N_10383,N_9878,N_9600);
or U10384 (N_10384,N_9937,N_9944);
xnor U10385 (N_10385,N_9602,N_9523);
nand U10386 (N_10386,N_9539,N_9887);
and U10387 (N_10387,N_9891,N_9965);
and U10388 (N_10388,N_9650,N_9811);
and U10389 (N_10389,N_9824,N_9720);
nand U10390 (N_10390,N_9570,N_9757);
and U10391 (N_10391,N_9531,N_9859);
and U10392 (N_10392,N_9960,N_9967);
xnor U10393 (N_10393,N_9804,N_9500);
xnor U10394 (N_10394,N_9935,N_9580);
nand U10395 (N_10395,N_9538,N_9874);
and U10396 (N_10396,N_9977,N_9744);
and U10397 (N_10397,N_9819,N_9942);
nand U10398 (N_10398,N_9753,N_9934);
nand U10399 (N_10399,N_9831,N_9610);
or U10400 (N_10400,N_9883,N_9992);
or U10401 (N_10401,N_9644,N_9574);
nor U10402 (N_10402,N_9652,N_9749);
nand U10403 (N_10403,N_9714,N_9563);
nand U10404 (N_10404,N_9518,N_9796);
nor U10405 (N_10405,N_9768,N_9694);
or U10406 (N_10406,N_9599,N_9648);
or U10407 (N_10407,N_9778,N_9826);
and U10408 (N_10408,N_9843,N_9967);
nor U10409 (N_10409,N_9584,N_9667);
nand U10410 (N_10410,N_9709,N_9876);
nand U10411 (N_10411,N_9973,N_9513);
or U10412 (N_10412,N_9910,N_9672);
nor U10413 (N_10413,N_9675,N_9519);
nand U10414 (N_10414,N_9802,N_9872);
nand U10415 (N_10415,N_9757,N_9624);
nor U10416 (N_10416,N_9508,N_9682);
nand U10417 (N_10417,N_9974,N_9650);
and U10418 (N_10418,N_9947,N_9991);
nand U10419 (N_10419,N_9581,N_9579);
and U10420 (N_10420,N_9841,N_9667);
or U10421 (N_10421,N_9517,N_9776);
and U10422 (N_10422,N_9543,N_9683);
nor U10423 (N_10423,N_9911,N_9642);
xnor U10424 (N_10424,N_9791,N_9816);
or U10425 (N_10425,N_9754,N_9793);
and U10426 (N_10426,N_9562,N_9822);
or U10427 (N_10427,N_9766,N_9913);
xnor U10428 (N_10428,N_9956,N_9944);
nor U10429 (N_10429,N_9602,N_9797);
or U10430 (N_10430,N_9910,N_9645);
nor U10431 (N_10431,N_9677,N_9949);
nand U10432 (N_10432,N_9543,N_9560);
xnor U10433 (N_10433,N_9639,N_9858);
nand U10434 (N_10434,N_9785,N_9556);
nand U10435 (N_10435,N_9589,N_9530);
nand U10436 (N_10436,N_9713,N_9742);
and U10437 (N_10437,N_9506,N_9645);
and U10438 (N_10438,N_9686,N_9668);
nand U10439 (N_10439,N_9977,N_9904);
or U10440 (N_10440,N_9963,N_9731);
and U10441 (N_10441,N_9589,N_9997);
xor U10442 (N_10442,N_9969,N_9558);
or U10443 (N_10443,N_9552,N_9590);
nand U10444 (N_10444,N_9700,N_9963);
xor U10445 (N_10445,N_9676,N_9936);
or U10446 (N_10446,N_9511,N_9872);
nand U10447 (N_10447,N_9983,N_9901);
nand U10448 (N_10448,N_9505,N_9660);
nor U10449 (N_10449,N_9535,N_9828);
xnor U10450 (N_10450,N_9586,N_9990);
or U10451 (N_10451,N_9567,N_9919);
nor U10452 (N_10452,N_9723,N_9682);
or U10453 (N_10453,N_9770,N_9836);
xor U10454 (N_10454,N_9951,N_9557);
xnor U10455 (N_10455,N_9959,N_9553);
and U10456 (N_10456,N_9918,N_9916);
and U10457 (N_10457,N_9626,N_9536);
nor U10458 (N_10458,N_9866,N_9901);
or U10459 (N_10459,N_9915,N_9871);
or U10460 (N_10460,N_9718,N_9674);
nor U10461 (N_10461,N_9846,N_9644);
nand U10462 (N_10462,N_9688,N_9715);
nand U10463 (N_10463,N_9509,N_9943);
and U10464 (N_10464,N_9720,N_9899);
xor U10465 (N_10465,N_9567,N_9645);
nand U10466 (N_10466,N_9708,N_9997);
and U10467 (N_10467,N_9783,N_9878);
and U10468 (N_10468,N_9541,N_9540);
nand U10469 (N_10469,N_9967,N_9983);
and U10470 (N_10470,N_9863,N_9860);
and U10471 (N_10471,N_9761,N_9539);
xnor U10472 (N_10472,N_9796,N_9946);
or U10473 (N_10473,N_9586,N_9628);
or U10474 (N_10474,N_9981,N_9587);
or U10475 (N_10475,N_9827,N_9695);
and U10476 (N_10476,N_9983,N_9852);
xor U10477 (N_10477,N_9602,N_9667);
and U10478 (N_10478,N_9929,N_9822);
xor U10479 (N_10479,N_9536,N_9970);
xnor U10480 (N_10480,N_9670,N_9911);
or U10481 (N_10481,N_9730,N_9602);
and U10482 (N_10482,N_9629,N_9775);
xor U10483 (N_10483,N_9561,N_9668);
and U10484 (N_10484,N_9624,N_9953);
nand U10485 (N_10485,N_9849,N_9843);
nor U10486 (N_10486,N_9685,N_9927);
and U10487 (N_10487,N_9952,N_9579);
and U10488 (N_10488,N_9519,N_9624);
nand U10489 (N_10489,N_9881,N_9851);
xor U10490 (N_10490,N_9818,N_9769);
nor U10491 (N_10491,N_9952,N_9980);
and U10492 (N_10492,N_9649,N_9673);
and U10493 (N_10493,N_9908,N_9639);
xor U10494 (N_10494,N_9520,N_9797);
nor U10495 (N_10495,N_9889,N_9757);
or U10496 (N_10496,N_9547,N_9951);
and U10497 (N_10497,N_9621,N_9968);
nand U10498 (N_10498,N_9966,N_9571);
nor U10499 (N_10499,N_9586,N_9661);
nor U10500 (N_10500,N_10488,N_10199);
or U10501 (N_10501,N_10484,N_10163);
nand U10502 (N_10502,N_10364,N_10128);
xor U10503 (N_10503,N_10007,N_10231);
nor U10504 (N_10504,N_10466,N_10308);
xor U10505 (N_10505,N_10075,N_10464);
nand U10506 (N_10506,N_10437,N_10369);
xnor U10507 (N_10507,N_10181,N_10136);
nor U10508 (N_10508,N_10203,N_10458);
xnor U10509 (N_10509,N_10479,N_10173);
and U10510 (N_10510,N_10497,N_10202);
and U10511 (N_10511,N_10306,N_10017);
and U10512 (N_10512,N_10088,N_10122);
or U10513 (N_10513,N_10197,N_10030);
or U10514 (N_10514,N_10061,N_10120);
xor U10515 (N_10515,N_10441,N_10036);
xor U10516 (N_10516,N_10489,N_10328);
nor U10517 (N_10517,N_10216,N_10037);
and U10518 (N_10518,N_10327,N_10486);
or U10519 (N_10519,N_10326,N_10444);
nand U10520 (N_10520,N_10279,N_10057);
nor U10521 (N_10521,N_10431,N_10359);
and U10522 (N_10522,N_10131,N_10456);
or U10523 (N_10523,N_10217,N_10288);
and U10524 (N_10524,N_10370,N_10186);
or U10525 (N_10525,N_10277,N_10013);
xnor U10526 (N_10526,N_10092,N_10038);
xnor U10527 (N_10527,N_10302,N_10195);
nand U10528 (N_10528,N_10093,N_10407);
nor U10529 (N_10529,N_10244,N_10281);
or U10530 (N_10530,N_10457,N_10297);
nor U10531 (N_10531,N_10149,N_10276);
and U10532 (N_10532,N_10353,N_10460);
or U10533 (N_10533,N_10108,N_10106);
nand U10534 (N_10534,N_10085,N_10135);
xor U10535 (N_10535,N_10463,N_10132);
xor U10536 (N_10536,N_10494,N_10314);
and U10537 (N_10537,N_10212,N_10318);
or U10538 (N_10538,N_10361,N_10062);
nand U10539 (N_10539,N_10254,N_10041);
nor U10540 (N_10540,N_10298,N_10170);
nor U10541 (N_10541,N_10180,N_10099);
and U10542 (N_10542,N_10016,N_10011);
or U10543 (N_10543,N_10225,N_10176);
and U10544 (N_10544,N_10204,N_10090);
and U10545 (N_10545,N_10426,N_10159);
or U10546 (N_10546,N_10413,N_10393);
or U10547 (N_10547,N_10461,N_10351);
nor U10548 (N_10548,N_10223,N_10481);
nor U10549 (N_10549,N_10472,N_10236);
nor U10550 (N_10550,N_10070,N_10201);
or U10551 (N_10551,N_10336,N_10033);
xnor U10552 (N_10552,N_10433,N_10060);
nor U10553 (N_10553,N_10121,N_10076);
and U10554 (N_10554,N_10144,N_10452);
xor U10555 (N_10555,N_10210,N_10487);
xnor U10556 (N_10556,N_10271,N_10443);
xnor U10557 (N_10557,N_10145,N_10262);
or U10558 (N_10558,N_10304,N_10394);
nand U10559 (N_10559,N_10450,N_10415);
or U10560 (N_10560,N_10242,N_10348);
or U10561 (N_10561,N_10293,N_10005);
xor U10562 (N_10562,N_10250,N_10332);
nand U10563 (N_10563,N_10429,N_10403);
and U10564 (N_10564,N_10490,N_10385);
and U10565 (N_10565,N_10410,N_10357);
nand U10566 (N_10566,N_10229,N_10107);
nand U10567 (N_10567,N_10072,N_10226);
xor U10568 (N_10568,N_10171,N_10100);
nor U10569 (N_10569,N_10193,N_10148);
xor U10570 (N_10570,N_10356,N_10454);
xor U10571 (N_10571,N_10377,N_10367);
xor U10572 (N_10572,N_10268,N_10152);
nand U10573 (N_10573,N_10470,N_10014);
xor U10574 (N_10574,N_10074,N_10028);
nor U10575 (N_10575,N_10485,N_10096);
xnor U10576 (N_10576,N_10333,N_10065);
and U10577 (N_10577,N_10143,N_10315);
or U10578 (N_10578,N_10018,N_10162);
nand U10579 (N_10579,N_10004,N_10255);
or U10580 (N_10580,N_10300,N_10027);
nand U10581 (N_10581,N_10425,N_10246);
or U10582 (N_10582,N_10418,N_10267);
or U10583 (N_10583,N_10087,N_10329);
and U10584 (N_10584,N_10423,N_10139);
nor U10585 (N_10585,N_10167,N_10000);
xnor U10586 (N_10586,N_10445,N_10233);
and U10587 (N_10587,N_10051,N_10227);
nand U10588 (N_10588,N_10430,N_10408);
nand U10589 (N_10589,N_10138,N_10161);
and U10590 (N_10590,N_10307,N_10113);
xnor U10591 (N_10591,N_10183,N_10218);
nor U10592 (N_10592,N_10105,N_10346);
xor U10593 (N_10593,N_10234,N_10048);
nand U10594 (N_10594,N_10035,N_10272);
and U10595 (N_10595,N_10260,N_10256);
or U10596 (N_10596,N_10140,N_10383);
nor U10597 (N_10597,N_10240,N_10335);
and U10598 (N_10598,N_10436,N_10118);
nand U10599 (N_10599,N_10371,N_10378);
or U10600 (N_10600,N_10147,N_10134);
or U10601 (N_10601,N_10398,N_10438);
or U10602 (N_10602,N_10241,N_10182);
and U10603 (N_10603,N_10400,N_10282);
or U10604 (N_10604,N_10200,N_10311);
and U10605 (N_10605,N_10360,N_10355);
and U10606 (N_10606,N_10101,N_10372);
nor U10607 (N_10607,N_10191,N_10285);
and U10608 (N_10608,N_10015,N_10290);
nor U10609 (N_10609,N_10273,N_10362);
xnor U10610 (N_10610,N_10006,N_10402);
and U10611 (N_10611,N_10416,N_10386);
and U10612 (N_10612,N_10230,N_10341);
nor U10613 (N_10613,N_10495,N_10141);
nor U10614 (N_10614,N_10381,N_10350);
nand U10615 (N_10615,N_10067,N_10428);
or U10616 (N_10616,N_10097,N_10366);
or U10617 (N_10617,N_10373,N_10153);
nor U10618 (N_10618,N_10449,N_10387);
xnor U10619 (N_10619,N_10211,N_10059);
and U10620 (N_10620,N_10069,N_10185);
or U10621 (N_10621,N_10160,N_10330);
nor U10622 (N_10622,N_10082,N_10248);
xor U10623 (N_10623,N_10349,N_10114);
nand U10624 (N_10624,N_10239,N_10053);
and U10625 (N_10625,N_10492,N_10352);
nor U10626 (N_10626,N_10363,N_10208);
nand U10627 (N_10627,N_10468,N_10404);
xor U10628 (N_10628,N_10042,N_10280);
xor U10629 (N_10629,N_10079,N_10344);
xnor U10630 (N_10630,N_10414,N_10001);
nand U10631 (N_10631,N_10409,N_10469);
xnor U10632 (N_10632,N_10411,N_10274);
nand U10633 (N_10633,N_10104,N_10392);
or U10634 (N_10634,N_10374,N_10050);
nor U10635 (N_10635,N_10265,N_10112);
or U10636 (N_10636,N_10026,N_10179);
nor U10637 (N_10637,N_10368,N_10440);
xnor U10638 (N_10638,N_10483,N_10467);
or U10639 (N_10639,N_10146,N_10309);
xnor U10640 (N_10640,N_10261,N_10382);
xor U10641 (N_10641,N_10405,N_10220);
nor U10642 (N_10642,N_10124,N_10039);
xnor U10643 (N_10643,N_10046,N_10459);
xor U10644 (N_10644,N_10156,N_10157);
and U10645 (N_10645,N_10102,N_10083);
nor U10646 (N_10646,N_10068,N_10365);
nor U10647 (N_10647,N_10294,N_10324);
xnor U10648 (N_10648,N_10024,N_10286);
nand U10649 (N_10649,N_10435,N_10063);
and U10650 (N_10650,N_10189,N_10424);
or U10651 (N_10651,N_10040,N_10482);
nand U10652 (N_10652,N_10137,N_10275);
and U10653 (N_10653,N_10342,N_10071);
nor U10654 (N_10654,N_10119,N_10094);
or U10655 (N_10655,N_10192,N_10086);
and U10656 (N_10656,N_10080,N_10379);
nand U10657 (N_10657,N_10177,N_10129);
and U10658 (N_10658,N_10009,N_10044);
nor U10659 (N_10659,N_10008,N_10187);
or U10660 (N_10660,N_10310,N_10184);
nor U10661 (N_10661,N_10178,N_10023);
or U10662 (N_10662,N_10020,N_10130);
xnor U10663 (N_10663,N_10194,N_10451);
or U10664 (N_10664,N_10209,N_10150);
xor U10665 (N_10665,N_10228,N_10391);
nand U10666 (N_10666,N_10066,N_10109);
nor U10667 (N_10667,N_10376,N_10439);
xnor U10668 (N_10668,N_10213,N_10455);
or U10669 (N_10669,N_10078,N_10316);
xnor U10670 (N_10670,N_10269,N_10343);
and U10671 (N_10671,N_10055,N_10238);
xnor U10672 (N_10672,N_10207,N_10442);
or U10673 (N_10673,N_10084,N_10476);
and U10674 (N_10674,N_10012,N_10043);
and U10675 (N_10675,N_10251,N_10299);
or U10676 (N_10676,N_10295,N_10421);
and U10677 (N_10677,N_10125,N_10224);
or U10678 (N_10678,N_10221,N_10253);
or U10679 (N_10679,N_10320,N_10338);
and U10680 (N_10680,N_10243,N_10312);
or U10681 (N_10681,N_10205,N_10258);
nand U10682 (N_10682,N_10115,N_10422);
xor U10683 (N_10683,N_10049,N_10264);
nor U10684 (N_10684,N_10358,N_10222);
nor U10685 (N_10685,N_10127,N_10245);
and U10686 (N_10686,N_10188,N_10303);
and U10687 (N_10687,N_10396,N_10175);
nand U10688 (N_10688,N_10287,N_10206);
nor U10689 (N_10689,N_10263,N_10214);
nand U10690 (N_10690,N_10462,N_10133);
nand U10691 (N_10691,N_10031,N_10165);
and U10692 (N_10692,N_10491,N_10022);
or U10693 (N_10693,N_10142,N_10103);
and U10694 (N_10694,N_10434,N_10313);
or U10695 (N_10695,N_10412,N_10252);
and U10696 (N_10696,N_10323,N_10319);
nand U10697 (N_10697,N_10052,N_10420);
xor U10698 (N_10698,N_10045,N_10389);
nand U10699 (N_10699,N_10499,N_10446);
or U10700 (N_10700,N_10453,N_10432);
xnor U10701 (N_10701,N_10278,N_10081);
nand U10702 (N_10702,N_10337,N_10475);
nor U10703 (N_10703,N_10419,N_10126);
xnor U10704 (N_10704,N_10190,N_10375);
and U10705 (N_10705,N_10219,N_10390);
nand U10706 (N_10706,N_10098,N_10388);
or U10707 (N_10707,N_10283,N_10073);
nand U10708 (N_10708,N_10003,N_10291);
xor U10709 (N_10709,N_10447,N_10091);
or U10710 (N_10710,N_10032,N_10002);
nand U10711 (N_10711,N_10010,N_10384);
xor U10712 (N_10712,N_10117,N_10448);
xnor U10713 (N_10713,N_10164,N_10334);
nand U10714 (N_10714,N_10340,N_10301);
xor U10715 (N_10715,N_10331,N_10168);
or U10716 (N_10716,N_10347,N_10465);
and U10717 (N_10717,N_10056,N_10077);
xor U10718 (N_10718,N_10284,N_10417);
or U10719 (N_10719,N_10480,N_10172);
nand U10720 (N_10720,N_10025,N_10174);
nand U10721 (N_10721,N_10166,N_10054);
and U10722 (N_10722,N_10401,N_10111);
xnor U10723 (N_10723,N_10292,N_10322);
xnor U10724 (N_10724,N_10270,N_10498);
nand U10725 (N_10725,N_10305,N_10047);
nand U10726 (N_10726,N_10493,N_10198);
nor U10727 (N_10727,N_10259,N_10395);
nor U10728 (N_10728,N_10232,N_10289);
nor U10729 (N_10729,N_10266,N_10169);
nand U10730 (N_10730,N_10123,N_10380);
and U10731 (N_10731,N_10158,N_10496);
or U10732 (N_10732,N_10317,N_10325);
nor U10733 (N_10733,N_10196,N_10215);
and U10734 (N_10734,N_10058,N_10473);
xor U10735 (N_10735,N_10406,N_10345);
or U10736 (N_10736,N_10064,N_10154);
nand U10737 (N_10737,N_10399,N_10110);
nand U10738 (N_10738,N_10034,N_10474);
nand U10739 (N_10739,N_10089,N_10249);
nor U10740 (N_10740,N_10471,N_10339);
xnor U10741 (N_10741,N_10237,N_10155);
or U10742 (N_10742,N_10247,N_10151);
nor U10743 (N_10743,N_10019,N_10095);
and U10744 (N_10744,N_10321,N_10257);
nor U10745 (N_10745,N_10477,N_10478);
nand U10746 (N_10746,N_10296,N_10116);
and U10747 (N_10747,N_10235,N_10029);
nor U10748 (N_10748,N_10397,N_10427);
xnor U10749 (N_10749,N_10354,N_10021);
xnor U10750 (N_10750,N_10263,N_10149);
nand U10751 (N_10751,N_10373,N_10441);
nand U10752 (N_10752,N_10334,N_10112);
xnor U10753 (N_10753,N_10442,N_10350);
or U10754 (N_10754,N_10392,N_10470);
and U10755 (N_10755,N_10259,N_10245);
nor U10756 (N_10756,N_10468,N_10236);
and U10757 (N_10757,N_10255,N_10077);
xnor U10758 (N_10758,N_10479,N_10249);
nand U10759 (N_10759,N_10302,N_10278);
nor U10760 (N_10760,N_10438,N_10402);
xor U10761 (N_10761,N_10435,N_10213);
or U10762 (N_10762,N_10203,N_10160);
nor U10763 (N_10763,N_10414,N_10491);
xor U10764 (N_10764,N_10313,N_10394);
nand U10765 (N_10765,N_10127,N_10181);
and U10766 (N_10766,N_10498,N_10047);
or U10767 (N_10767,N_10441,N_10444);
and U10768 (N_10768,N_10406,N_10076);
xor U10769 (N_10769,N_10091,N_10058);
or U10770 (N_10770,N_10385,N_10006);
xnor U10771 (N_10771,N_10263,N_10318);
xnor U10772 (N_10772,N_10096,N_10172);
nand U10773 (N_10773,N_10469,N_10281);
nor U10774 (N_10774,N_10349,N_10411);
nor U10775 (N_10775,N_10157,N_10025);
or U10776 (N_10776,N_10455,N_10423);
and U10777 (N_10777,N_10038,N_10440);
nand U10778 (N_10778,N_10226,N_10097);
and U10779 (N_10779,N_10423,N_10060);
nand U10780 (N_10780,N_10007,N_10038);
and U10781 (N_10781,N_10085,N_10411);
and U10782 (N_10782,N_10026,N_10224);
or U10783 (N_10783,N_10223,N_10365);
nor U10784 (N_10784,N_10243,N_10095);
and U10785 (N_10785,N_10275,N_10439);
nor U10786 (N_10786,N_10383,N_10134);
xor U10787 (N_10787,N_10081,N_10415);
or U10788 (N_10788,N_10388,N_10077);
xor U10789 (N_10789,N_10312,N_10198);
and U10790 (N_10790,N_10004,N_10113);
nand U10791 (N_10791,N_10336,N_10407);
nand U10792 (N_10792,N_10483,N_10098);
nor U10793 (N_10793,N_10149,N_10063);
and U10794 (N_10794,N_10206,N_10148);
xnor U10795 (N_10795,N_10060,N_10026);
xor U10796 (N_10796,N_10170,N_10141);
and U10797 (N_10797,N_10272,N_10016);
or U10798 (N_10798,N_10333,N_10097);
and U10799 (N_10799,N_10096,N_10351);
nand U10800 (N_10800,N_10303,N_10278);
nand U10801 (N_10801,N_10411,N_10374);
nand U10802 (N_10802,N_10471,N_10468);
or U10803 (N_10803,N_10222,N_10438);
or U10804 (N_10804,N_10062,N_10301);
nor U10805 (N_10805,N_10332,N_10100);
xnor U10806 (N_10806,N_10135,N_10118);
nor U10807 (N_10807,N_10024,N_10421);
nor U10808 (N_10808,N_10053,N_10219);
nor U10809 (N_10809,N_10393,N_10444);
nand U10810 (N_10810,N_10343,N_10028);
nand U10811 (N_10811,N_10155,N_10261);
xnor U10812 (N_10812,N_10388,N_10169);
or U10813 (N_10813,N_10390,N_10366);
xnor U10814 (N_10814,N_10223,N_10272);
nor U10815 (N_10815,N_10413,N_10323);
nor U10816 (N_10816,N_10123,N_10289);
nand U10817 (N_10817,N_10191,N_10224);
nor U10818 (N_10818,N_10366,N_10011);
xor U10819 (N_10819,N_10228,N_10496);
nand U10820 (N_10820,N_10189,N_10305);
nand U10821 (N_10821,N_10406,N_10209);
nand U10822 (N_10822,N_10412,N_10229);
or U10823 (N_10823,N_10259,N_10313);
or U10824 (N_10824,N_10272,N_10080);
and U10825 (N_10825,N_10282,N_10008);
nand U10826 (N_10826,N_10044,N_10095);
nand U10827 (N_10827,N_10160,N_10097);
or U10828 (N_10828,N_10367,N_10204);
nor U10829 (N_10829,N_10452,N_10451);
nor U10830 (N_10830,N_10066,N_10264);
and U10831 (N_10831,N_10250,N_10197);
xor U10832 (N_10832,N_10119,N_10226);
nor U10833 (N_10833,N_10154,N_10061);
and U10834 (N_10834,N_10334,N_10499);
xnor U10835 (N_10835,N_10359,N_10435);
xor U10836 (N_10836,N_10292,N_10297);
or U10837 (N_10837,N_10277,N_10068);
xor U10838 (N_10838,N_10118,N_10056);
nand U10839 (N_10839,N_10019,N_10157);
or U10840 (N_10840,N_10022,N_10490);
xor U10841 (N_10841,N_10238,N_10394);
nand U10842 (N_10842,N_10012,N_10325);
and U10843 (N_10843,N_10420,N_10262);
xor U10844 (N_10844,N_10342,N_10471);
nand U10845 (N_10845,N_10479,N_10320);
and U10846 (N_10846,N_10408,N_10208);
nor U10847 (N_10847,N_10017,N_10429);
xor U10848 (N_10848,N_10285,N_10124);
nor U10849 (N_10849,N_10025,N_10101);
xor U10850 (N_10850,N_10185,N_10147);
xor U10851 (N_10851,N_10321,N_10199);
and U10852 (N_10852,N_10067,N_10020);
xnor U10853 (N_10853,N_10203,N_10074);
nand U10854 (N_10854,N_10366,N_10063);
or U10855 (N_10855,N_10039,N_10474);
or U10856 (N_10856,N_10454,N_10005);
nor U10857 (N_10857,N_10190,N_10459);
and U10858 (N_10858,N_10351,N_10496);
xnor U10859 (N_10859,N_10199,N_10208);
or U10860 (N_10860,N_10043,N_10041);
xor U10861 (N_10861,N_10272,N_10398);
nor U10862 (N_10862,N_10410,N_10133);
and U10863 (N_10863,N_10395,N_10381);
or U10864 (N_10864,N_10458,N_10335);
or U10865 (N_10865,N_10496,N_10155);
and U10866 (N_10866,N_10033,N_10416);
nor U10867 (N_10867,N_10468,N_10141);
xnor U10868 (N_10868,N_10219,N_10214);
nor U10869 (N_10869,N_10002,N_10013);
xnor U10870 (N_10870,N_10348,N_10269);
nor U10871 (N_10871,N_10434,N_10307);
xnor U10872 (N_10872,N_10474,N_10392);
nand U10873 (N_10873,N_10420,N_10088);
nand U10874 (N_10874,N_10495,N_10267);
or U10875 (N_10875,N_10039,N_10309);
and U10876 (N_10876,N_10040,N_10483);
nand U10877 (N_10877,N_10146,N_10072);
nor U10878 (N_10878,N_10196,N_10396);
and U10879 (N_10879,N_10313,N_10113);
or U10880 (N_10880,N_10065,N_10387);
nor U10881 (N_10881,N_10361,N_10085);
and U10882 (N_10882,N_10198,N_10340);
xnor U10883 (N_10883,N_10363,N_10290);
or U10884 (N_10884,N_10129,N_10423);
nor U10885 (N_10885,N_10428,N_10269);
nand U10886 (N_10886,N_10224,N_10307);
nand U10887 (N_10887,N_10414,N_10154);
and U10888 (N_10888,N_10103,N_10061);
and U10889 (N_10889,N_10152,N_10326);
nand U10890 (N_10890,N_10402,N_10442);
xnor U10891 (N_10891,N_10000,N_10280);
nor U10892 (N_10892,N_10186,N_10492);
nand U10893 (N_10893,N_10005,N_10234);
and U10894 (N_10894,N_10208,N_10177);
or U10895 (N_10895,N_10110,N_10375);
nor U10896 (N_10896,N_10057,N_10141);
nand U10897 (N_10897,N_10089,N_10466);
and U10898 (N_10898,N_10049,N_10180);
nand U10899 (N_10899,N_10237,N_10063);
nand U10900 (N_10900,N_10311,N_10108);
and U10901 (N_10901,N_10236,N_10160);
nand U10902 (N_10902,N_10320,N_10046);
and U10903 (N_10903,N_10028,N_10247);
xnor U10904 (N_10904,N_10385,N_10451);
and U10905 (N_10905,N_10156,N_10278);
nor U10906 (N_10906,N_10448,N_10461);
or U10907 (N_10907,N_10495,N_10065);
and U10908 (N_10908,N_10410,N_10359);
and U10909 (N_10909,N_10115,N_10143);
nor U10910 (N_10910,N_10136,N_10219);
nor U10911 (N_10911,N_10349,N_10056);
nand U10912 (N_10912,N_10431,N_10111);
nor U10913 (N_10913,N_10295,N_10067);
xnor U10914 (N_10914,N_10209,N_10444);
nor U10915 (N_10915,N_10319,N_10145);
xor U10916 (N_10916,N_10299,N_10436);
xnor U10917 (N_10917,N_10096,N_10099);
nand U10918 (N_10918,N_10183,N_10165);
or U10919 (N_10919,N_10456,N_10222);
or U10920 (N_10920,N_10079,N_10413);
nand U10921 (N_10921,N_10413,N_10463);
or U10922 (N_10922,N_10451,N_10141);
xor U10923 (N_10923,N_10471,N_10168);
nor U10924 (N_10924,N_10382,N_10138);
nand U10925 (N_10925,N_10344,N_10125);
and U10926 (N_10926,N_10340,N_10224);
nor U10927 (N_10927,N_10283,N_10259);
and U10928 (N_10928,N_10450,N_10391);
nand U10929 (N_10929,N_10494,N_10273);
xnor U10930 (N_10930,N_10357,N_10463);
nand U10931 (N_10931,N_10361,N_10286);
and U10932 (N_10932,N_10269,N_10337);
nor U10933 (N_10933,N_10228,N_10168);
nand U10934 (N_10934,N_10371,N_10353);
xnor U10935 (N_10935,N_10462,N_10157);
nand U10936 (N_10936,N_10144,N_10124);
xor U10937 (N_10937,N_10031,N_10142);
and U10938 (N_10938,N_10140,N_10139);
xnor U10939 (N_10939,N_10389,N_10150);
nor U10940 (N_10940,N_10378,N_10057);
xnor U10941 (N_10941,N_10272,N_10122);
nor U10942 (N_10942,N_10171,N_10456);
nor U10943 (N_10943,N_10170,N_10080);
and U10944 (N_10944,N_10063,N_10358);
nand U10945 (N_10945,N_10046,N_10463);
nor U10946 (N_10946,N_10452,N_10460);
and U10947 (N_10947,N_10005,N_10021);
and U10948 (N_10948,N_10098,N_10468);
nand U10949 (N_10949,N_10475,N_10230);
nand U10950 (N_10950,N_10456,N_10467);
nor U10951 (N_10951,N_10088,N_10143);
xor U10952 (N_10952,N_10301,N_10465);
and U10953 (N_10953,N_10393,N_10143);
and U10954 (N_10954,N_10496,N_10326);
nand U10955 (N_10955,N_10486,N_10456);
nor U10956 (N_10956,N_10309,N_10233);
nand U10957 (N_10957,N_10055,N_10375);
and U10958 (N_10958,N_10120,N_10068);
nand U10959 (N_10959,N_10092,N_10376);
nand U10960 (N_10960,N_10450,N_10003);
and U10961 (N_10961,N_10423,N_10030);
nor U10962 (N_10962,N_10174,N_10076);
and U10963 (N_10963,N_10335,N_10088);
nand U10964 (N_10964,N_10467,N_10209);
nand U10965 (N_10965,N_10292,N_10095);
nand U10966 (N_10966,N_10096,N_10388);
xor U10967 (N_10967,N_10196,N_10399);
xor U10968 (N_10968,N_10185,N_10276);
xnor U10969 (N_10969,N_10107,N_10157);
or U10970 (N_10970,N_10346,N_10309);
nand U10971 (N_10971,N_10434,N_10364);
nor U10972 (N_10972,N_10478,N_10399);
xor U10973 (N_10973,N_10196,N_10392);
and U10974 (N_10974,N_10043,N_10011);
xor U10975 (N_10975,N_10454,N_10420);
or U10976 (N_10976,N_10011,N_10435);
nor U10977 (N_10977,N_10287,N_10305);
xnor U10978 (N_10978,N_10353,N_10015);
xnor U10979 (N_10979,N_10246,N_10402);
nand U10980 (N_10980,N_10055,N_10479);
or U10981 (N_10981,N_10129,N_10351);
nand U10982 (N_10982,N_10377,N_10169);
and U10983 (N_10983,N_10327,N_10374);
or U10984 (N_10984,N_10271,N_10496);
nor U10985 (N_10985,N_10201,N_10222);
and U10986 (N_10986,N_10433,N_10447);
nand U10987 (N_10987,N_10243,N_10205);
xor U10988 (N_10988,N_10126,N_10077);
nor U10989 (N_10989,N_10448,N_10280);
and U10990 (N_10990,N_10361,N_10379);
nand U10991 (N_10991,N_10117,N_10335);
or U10992 (N_10992,N_10072,N_10191);
nand U10993 (N_10993,N_10499,N_10247);
and U10994 (N_10994,N_10287,N_10304);
nor U10995 (N_10995,N_10111,N_10272);
and U10996 (N_10996,N_10233,N_10411);
nor U10997 (N_10997,N_10391,N_10384);
xnor U10998 (N_10998,N_10155,N_10466);
and U10999 (N_10999,N_10498,N_10273);
xnor U11000 (N_11000,N_10754,N_10605);
and U11001 (N_11001,N_10867,N_10748);
and U11002 (N_11002,N_10523,N_10686);
or U11003 (N_11003,N_10584,N_10769);
or U11004 (N_11004,N_10690,N_10619);
xnor U11005 (N_11005,N_10931,N_10961);
and U11006 (N_11006,N_10892,N_10580);
and U11007 (N_11007,N_10646,N_10777);
xor U11008 (N_11008,N_10661,N_10723);
and U11009 (N_11009,N_10551,N_10796);
nand U11010 (N_11010,N_10744,N_10573);
nand U11011 (N_11011,N_10572,N_10697);
nand U11012 (N_11012,N_10878,N_10921);
xor U11013 (N_11013,N_10631,N_10770);
nand U11014 (N_11014,N_10505,N_10622);
and U11015 (N_11015,N_10630,N_10677);
nor U11016 (N_11016,N_10706,N_10984);
xor U11017 (N_11017,N_10797,N_10521);
and U11018 (N_11018,N_10950,N_10876);
nand U11019 (N_11019,N_10731,N_10774);
nand U11020 (N_11020,N_10919,N_10541);
nor U11021 (N_11021,N_10801,N_10575);
and U11022 (N_11022,N_10717,N_10740);
nor U11023 (N_11023,N_10645,N_10910);
and U11024 (N_11024,N_10592,N_10597);
xor U11025 (N_11025,N_10904,N_10850);
and U11026 (N_11026,N_10888,N_10675);
or U11027 (N_11027,N_10739,N_10752);
and U11028 (N_11028,N_10606,N_10940);
or U11029 (N_11029,N_10725,N_10745);
xor U11030 (N_11030,N_10847,N_10542);
nor U11031 (N_11031,N_10989,N_10762);
nand U11032 (N_11032,N_10596,N_10798);
nor U11033 (N_11033,N_10555,N_10900);
or U11034 (N_11034,N_10535,N_10872);
nand U11035 (N_11035,N_10817,N_10917);
or U11036 (N_11036,N_10969,N_10670);
or U11037 (N_11037,N_10648,N_10810);
or U11038 (N_11038,N_10789,N_10966);
or U11039 (N_11039,N_10826,N_10565);
xor U11040 (N_11040,N_10906,N_10928);
nand U11041 (N_11041,N_10559,N_10895);
and U11042 (N_11042,N_10621,N_10517);
nor U11043 (N_11043,N_10953,N_10612);
or U11044 (N_11044,N_10977,N_10979);
nand U11045 (N_11045,N_10530,N_10948);
or U11046 (N_11046,N_10845,N_10874);
nand U11047 (N_11047,N_10511,N_10807);
and U11048 (N_11048,N_10837,N_10776);
or U11049 (N_11049,N_10624,N_10784);
nand U11050 (N_11050,N_10960,N_10662);
nor U11051 (N_11051,N_10885,N_10768);
or U11052 (N_11052,N_10506,N_10897);
and U11053 (N_11053,N_10985,N_10841);
nand U11054 (N_11054,N_10813,N_10663);
nor U11055 (N_11055,N_10997,N_10665);
and U11056 (N_11056,N_10652,N_10905);
nor U11057 (N_11057,N_10839,N_10974);
nand U11058 (N_11058,N_10554,N_10773);
xor U11059 (N_11059,N_10550,N_10537);
xor U11060 (N_11060,N_10628,N_10812);
xor U11061 (N_11061,N_10684,N_10791);
nor U11062 (N_11062,N_10964,N_10608);
nor U11063 (N_11063,N_10669,N_10693);
and U11064 (N_11064,N_10560,N_10660);
xnor U11065 (N_11065,N_10503,N_10879);
or U11066 (N_11066,N_10688,N_10852);
and U11067 (N_11067,N_10519,N_10558);
and U11068 (N_11068,N_10702,N_10911);
nor U11069 (N_11069,N_10793,N_10716);
or U11070 (N_11070,N_10994,N_10935);
or U11071 (N_11071,N_10603,N_10644);
nand U11072 (N_11072,N_10576,N_10593);
nor U11073 (N_11073,N_10894,N_10790);
or U11074 (N_11074,N_10933,N_10712);
xnor U11075 (N_11075,N_10830,N_10949);
nor U11076 (N_11076,N_10861,N_10756);
or U11077 (N_11077,N_10705,N_10779);
and U11078 (N_11078,N_10722,N_10549);
nor U11079 (N_11079,N_10868,N_10912);
xor U11080 (N_11080,N_10816,N_10833);
xor U11081 (N_11081,N_10863,N_10650);
xor U11082 (N_11082,N_10751,N_10577);
nand U11083 (N_11083,N_10678,N_10540);
or U11084 (N_11084,N_10522,N_10823);
or U11085 (N_11085,N_10988,N_10618);
and U11086 (N_11086,N_10999,N_10610);
nor U11087 (N_11087,N_10729,N_10512);
nand U11088 (N_11088,N_10855,N_10902);
and U11089 (N_11089,N_10673,N_10724);
nand U11090 (N_11090,N_10591,N_10923);
nand U11091 (N_11091,N_10991,N_10736);
nand U11092 (N_11092,N_10757,N_10681);
or U11093 (N_11093,N_10636,N_10938);
or U11094 (N_11094,N_10571,N_10766);
nor U11095 (N_11095,N_10835,N_10708);
nor U11096 (N_11096,N_10915,N_10500);
nand U11097 (N_11097,N_10553,N_10598);
and U11098 (N_11098,N_10860,N_10844);
nor U11099 (N_11099,N_10590,N_10909);
xor U11100 (N_11100,N_10761,N_10747);
or U11101 (N_11101,N_10891,N_10694);
or U11102 (N_11102,N_10941,N_10846);
nor U11103 (N_11103,N_10834,N_10604);
nand U11104 (N_11104,N_10875,N_10795);
nand U11105 (N_11105,N_10857,N_10959);
or U11106 (N_11106,N_10674,N_10973);
and U11107 (N_11107,N_10581,N_10849);
xor U11108 (N_11108,N_10585,N_10651);
xnor U11109 (N_11109,N_10514,N_10516);
or U11110 (N_11110,N_10914,N_10924);
or U11111 (N_11111,N_10682,N_10574);
or U11112 (N_11112,N_10962,N_10561);
xnor U11113 (N_11113,N_10643,N_10714);
nor U11114 (N_11114,N_10548,N_10567);
nand U11115 (N_11115,N_10956,N_10582);
or U11116 (N_11116,N_10704,N_10562);
or U11117 (N_11117,N_10840,N_10749);
nor U11118 (N_11118,N_10710,N_10726);
nor U11119 (N_11119,N_10800,N_10901);
or U11120 (N_11120,N_10713,N_10502);
nand U11121 (N_11121,N_10806,N_10727);
nor U11122 (N_11122,N_10890,N_10822);
and U11123 (N_11123,N_10864,N_10711);
nand U11124 (N_11124,N_10544,N_10952);
nand U11125 (N_11125,N_10570,N_10926);
and U11126 (N_11126,N_10738,N_10589);
xor U11127 (N_11127,N_10680,N_10831);
xor U11128 (N_11128,N_10613,N_10629);
xor U11129 (N_11129,N_10944,N_10758);
nor U11130 (N_11130,N_10653,N_10578);
nand U11131 (N_11131,N_10918,N_10657);
nor U11132 (N_11132,N_10664,N_10579);
nor U11133 (N_11133,N_10683,N_10907);
or U11134 (N_11134,N_10980,N_10818);
xor U11135 (N_11135,N_10943,N_10764);
xnor U11136 (N_11136,N_10615,N_10767);
nand U11137 (N_11137,N_10987,N_10750);
nor U11138 (N_11138,N_10536,N_10529);
xor U11139 (N_11139,N_10692,N_10937);
or U11140 (N_11140,N_10945,N_10785);
nand U11141 (N_11141,N_10946,N_10720);
or U11142 (N_11142,N_10689,N_10698);
and U11143 (N_11143,N_10707,N_10869);
xor U11144 (N_11144,N_10709,N_10531);
nand U11145 (N_11145,N_10734,N_10982);
xnor U11146 (N_11146,N_10998,N_10760);
and U11147 (N_11147,N_10534,N_10996);
xor U11148 (N_11148,N_10504,N_10882);
xnor U11149 (N_11149,N_10922,N_10715);
and U11150 (N_11150,N_10967,N_10899);
nand U11151 (N_11151,N_10975,N_10859);
nor U11152 (N_11152,N_10815,N_10913);
or U11153 (N_11153,N_10583,N_10616);
nand U11154 (N_11154,N_10676,N_10925);
and U11155 (N_11155,N_10866,N_10611);
and U11156 (N_11156,N_10695,N_10699);
and U11157 (N_11157,N_10543,N_10625);
nor U11158 (N_11158,N_10970,N_10955);
nor U11159 (N_11159,N_10641,N_10501);
xor U11160 (N_11160,N_10799,N_10829);
xnor U11161 (N_11161,N_10755,N_10654);
or U11162 (N_11162,N_10658,N_10626);
xnor U11163 (N_11163,N_10842,N_10851);
and U11164 (N_11164,N_10557,N_10701);
and U11165 (N_11165,N_10667,N_10545);
xor U11166 (N_11166,N_10746,N_10633);
xor U11167 (N_11167,N_10507,N_10775);
xor U11168 (N_11168,N_10871,N_10836);
nor U11169 (N_11169,N_10634,N_10930);
nand U11170 (N_11170,N_10958,N_10820);
nand U11171 (N_11171,N_10508,N_10929);
or U11172 (N_11172,N_10513,N_10787);
and U11173 (N_11173,N_10995,N_10771);
and U11174 (N_11174,N_10916,N_10656);
or U11175 (N_11175,N_10783,N_10765);
and U11176 (N_11176,N_10951,N_10968);
or U11177 (N_11177,N_10642,N_10903);
or U11178 (N_11178,N_10732,N_10632);
nor U11179 (N_11179,N_10599,N_10600);
or U11180 (N_11180,N_10649,N_10635);
xor U11181 (N_11181,N_10533,N_10886);
nand U11182 (N_11182,N_10623,N_10957);
nand U11183 (N_11183,N_10547,N_10898);
and U11184 (N_11184,N_10990,N_10788);
nor U11185 (N_11185,N_10883,N_10856);
nor U11186 (N_11186,N_10602,N_10965);
xnor U11187 (N_11187,N_10936,N_10908);
nand U11188 (N_11188,N_10881,N_10568);
nor U11189 (N_11189,N_10672,N_10753);
or U11190 (N_11190,N_10601,N_10696);
or U11191 (N_11191,N_10587,N_10614);
nor U11192 (N_11192,N_10728,N_10877);
nand U11193 (N_11193,N_10978,N_10742);
or U11194 (N_11194,N_10538,N_10927);
nor U11195 (N_11195,N_10743,N_10862);
or U11196 (N_11196,N_10920,N_10700);
nand U11197 (N_11197,N_10832,N_10853);
nor U11198 (N_11198,N_10887,N_10719);
nand U11199 (N_11199,N_10792,N_10526);
nand U11200 (N_11200,N_10821,N_10735);
and U11201 (N_11201,N_10983,N_10786);
xnor U11202 (N_11202,N_10976,N_10532);
and U11203 (N_11203,N_10647,N_10620);
xor U11204 (N_11204,N_10594,N_10848);
nor U11205 (N_11205,N_10963,N_10563);
xor U11206 (N_11206,N_10564,N_10528);
xnor U11207 (N_11207,N_10981,N_10638);
nand U11208 (N_11208,N_10838,N_10781);
or U11209 (N_11209,N_10679,N_10527);
xnor U11210 (N_11210,N_10763,N_10827);
and U11211 (N_11211,N_10947,N_10971);
nor U11212 (N_11212,N_10640,N_10873);
or U11213 (N_11213,N_10659,N_10896);
xor U11214 (N_11214,N_10992,N_10730);
nand U11215 (N_11215,N_10782,N_10627);
nor U11216 (N_11216,N_10939,N_10655);
xor U11217 (N_11217,N_10954,N_10804);
and U11218 (N_11218,N_10607,N_10510);
nand U11219 (N_11219,N_10880,N_10552);
xor U11220 (N_11220,N_10802,N_10586);
xor U11221 (N_11221,N_10721,N_10778);
and U11222 (N_11222,N_10794,N_10843);
xnor U11223 (N_11223,N_10825,N_10805);
nand U11224 (N_11224,N_10685,N_10870);
xor U11225 (N_11225,N_10703,N_10518);
and U11226 (N_11226,N_10525,N_10828);
xnor U11227 (N_11227,N_10737,N_10520);
xor U11228 (N_11228,N_10854,N_10824);
and U11229 (N_11229,N_10671,N_10556);
nor U11230 (N_11230,N_10865,N_10637);
nand U11231 (N_11231,N_10609,N_10539);
nor U11232 (N_11232,N_10741,N_10819);
xor U11233 (N_11233,N_10889,N_10759);
and U11234 (N_11234,N_10666,N_10566);
or U11235 (N_11235,N_10809,N_10546);
nand U11236 (N_11236,N_10808,N_10858);
and U11237 (N_11237,N_10617,N_10588);
or U11238 (N_11238,N_10509,N_10814);
and U11239 (N_11239,N_10780,N_10668);
and U11240 (N_11240,N_10595,N_10772);
or U11241 (N_11241,N_10893,N_10687);
and U11242 (N_11242,N_10972,N_10733);
or U11243 (N_11243,N_10932,N_10986);
or U11244 (N_11244,N_10639,N_10811);
and U11245 (N_11245,N_10934,N_10942);
nand U11246 (N_11246,N_10803,N_10718);
and U11247 (N_11247,N_10569,N_10515);
or U11248 (N_11248,N_10524,N_10691);
nor U11249 (N_11249,N_10884,N_10993);
and U11250 (N_11250,N_10975,N_10510);
nand U11251 (N_11251,N_10873,N_10551);
nor U11252 (N_11252,N_10583,N_10708);
xnor U11253 (N_11253,N_10744,N_10797);
xnor U11254 (N_11254,N_10738,N_10542);
nand U11255 (N_11255,N_10939,N_10745);
nor U11256 (N_11256,N_10716,N_10858);
nand U11257 (N_11257,N_10720,N_10874);
or U11258 (N_11258,N_10655,N_10594);
or U11259 (N_11259,N_10589,N_10792);
nor U11260 (N_11260,N_10873,N_10936);
or U11261 (N_11261,N_10736,N_10809);
nand U11262 (N_11262,N_10808,N_10667);
or U11263 (N_11263,N_10746,N_10822);
or U11264 (N_11264,N_10955,N_10938);
nor U11265 (N_11265,N_10901,N_10970);
or U11266 (N_11266,N_10551,N_10647);
nor U11267 (N_11267,N_10750,N_10872);
nor U11268 (N_11268,N_10886,N_10566);
and U11269 (N_11269,N_10943,N_10515);
nand U11270 (N_11270,N_10506,N_10539);
nand U11271 (N_11271,N_10979,N_10814);
and U11272 (N_11272,N_10852,N_10816);
nand U11273 (N_11273,N_10653,N_10512);
or U11274 (N_11274,N_10583,N_10711);
nand U11275 (N_11275,N_10894,N_10846);
nor U11276 (N_11276,N_10933,N_10605);
xnor U11277 (N_11277,N_10665,N_10657);
nor U11278 (N_11278,N_10901,N_10703);
nor U11279 (N_11279,N_10877,N_10924);
nor U11280 (N_11280,N_10999,N_10697);
nand U11281 (N_11281,N_10514,N_10623);
xnor U11282 (N_11282,N_10877,N_10544);
nand U11283 (N_11283,N_10772,N_10814);
and U11284 (N_11284,N_10867,N_10928);
nor U11285 (N_11285,N_10976,N_10900);
xnor U11286 (N_11286,N_10623,N_10691);
nor U11287 (N_11287,N_10862,N_10551);
nand U11288 (N_11288,N_10815,N_10988);
nand U11289 (N_11289,N_10510,N_10799);
or U11290 (N_11290,N_10538,N_10941);
nand U11291 (N_11291,N_10611,N_10671);
or U11292 (N_11292,N_10772,N_10831);
nand U11293 (N_11293,N_10564,N_10888);
nor U11294 (N_11294,N_10928,N_10640);
or U11295 (N_11295,N_10501,N_10795);
nor U11296 (N_11296,N_10732,N_10926);
xnor U11297 (N_11297,N_10956,N_10623);
xnor U11298 (N_11298,N_10621,N_10725);
nand U11299 (N_11299,N_10614,N_10786);
nand U11300 (N_11300,N_10761,N_10568);
nor U11301 (N_11301,N_10633,N_10661);
nor U11302 (N_11302,N_10538,N_10604);
nor U11303 (N_11303,N_10952,N_10666);
and U11304 (N_11304,N_10975,N_10845);
nor U11305 (N_11305,N_10717,N_10919);
nor U11306 (N_11306,N_10814,N_10532);
or U11307 (N_11307,N_10691,N_10784);
nor U11308 (N_11308,N_10840,N_10991);
or U11309 (N_11309,N_10737,N_10771);
nor U11310 (N_11310,N_10835,N_10678);
nand U11311 (N_11311,N_10518,N_10722);
xor U11312 (N_11312,N_10618,N_10600);
nand U11313 (N_11313,N_10604,N_10526);
xor U11314 (N_11314,N_10894,N_10508);
nor U11315 (N_11315,N_10832,N_10761);
and U11316 (N_11316,N_10585,N_10719);
nand U11317 (N_11317,N_10505,N_10833);
nor U11318 (N_11318,N_10799,N_10934);
nand U11319 (N_11319,N_10919,N_10808);
nand U11320 (N_11320,N_10725,N_10692);
and U11321 (N_11321,N_10808,N_10854);
nor U11322 (N_11322,N_10996,N_10770);
nor U11323 (N_11323,N_10835,N_10816);
xor U11324 (N_11324,N_10558,N_10882);
and U11325 (N_11325,N_10695,N_10827);
nor U11326 (N_11326,N_10657,N_10566);
nand U11327 (N_11327,N_10599,N_10578);
and U11328 (N_11328,N_10543,N_10510);
xor U11329 (N_11329,N_10984,N_10516);
xor U11330 (N_11330,N_10857,N_10794);
nor U11331 (N_11331,N_10739,N_10947);
or U11332 (N_11332,N_10712,N_10640);
nand U11333 (N_11333,N_10552,N_10805);
xnor U11334 (N_11334,N_10746,N_10581);
and U11335 (N_11335,N_10638,N_10716);
or U11336 (N_11336,N_10885,N_10671);
nor U11337 (N_11337,N_10934,N_10653);
xor U11338 (N_11338,N_10766,N_10623);
nand U11339 (N_11339,N_10722,N_10836);
xor U11340 (N_11340,N_10617,N_10959);
nor U11341 (N_11341,N_10866,N_10895);
and U11342 (N_11342,N_10695,N_10583);
or U11343 (N_11343,N_10986,N_10776);
nor U11344 (N_11344,N_10892,N_10965);
nor U11345 (N_11345,N_10910,N_10771);
xor U11346 (N_11346,N_10708,N_10532);
nand U11347 (N_11347,N_10591,N_10956);
nand U11348 (N_11348,N_10696,N_10500);
and U11349 (N_11349,N_10847,N_10945);
xnor U11350 (N_11350,N_10548,N_10651);
or U11351 (N_11351,N_10633,N_10853);
nand U11352 (N_11352,N_10799,N_10566);
and U11353 (N_11353,N_10899,N_10841);
nor U11354 (N_11354,N_10647,N_10583);
nor U11355 (N_11355,N_10968,N_10572);
and U11356 (N_11356,N_10858,N_10578);
and U11357 (N_11357,N_10765,N_10742);
nand U11358 (N_11358,N_10552,N_10563);
and U11359 (N_11359,N_10871,N_10559);
xor U11360 (N_11360,N_10543,N_10679);
and U11361 (N_11361,N_10532,N_10954);
nand U11362 (N_11362,N_10869,N_10993);
and U11363 (N_11363,N_10863,N_10587);
nand U11364 (N_11364,N_10966,N_10761);
and U11365 (N_11365,N_10553,N_10787);
or U11366 (N_11366,N_10741,N_10988);
nand U11367 (N_11367,N_10782,N_10557);
and U11368 (N_11368,N_10955,N_10937);
xnor U11369 (N_11369,N_10636,N_10946);
and U11370 (N_11370,N_10996,N_10984);
and U11371 (N_11371,N_10606,N_10620);
nor U11372 (N_11372,N_10854,N_10583);
or U11373 (N_11373,N_10711,N_10661);
or U11374 (N_11374,N_10568,N_10514);
and U11375 (N_11375,N_10673,N_10601);
nand U11376 (N_11376,N_10508,N_10871);
nor U11377 (N_11377,N_10661,N_10957);
and U11378 (N_11378,N_10912,N_10750);
xnor U11379 (N_11379,N_10597,N_10678);
nor U11380 (N_11380,N_10816,N_10558);
or U11381 (N_11381,N_10919,N_10502);
nand U11382 (N_11382,N_10901,N_10678);
nand U11383 (N_11383,N_10935,N_10845);
or U11384 (N_11384,N_10765,N_10594);
xnor U11385 (N_11385,N_10525,N_10677);
and U11386 (N_11386,N_10875,N_10622);
and U11387 (N_11387,N_10768,N_10876);
nand U11388 (N_11388,N_10979,N_10850);
and U11389 (N_11389,N_10558,N_10679);
nor U11390 (N_11390,N_10851,N_10840);
xnor U11391 (N_11391,N_10565,N_10716);
and U11392 (N_11392,N_10908,N_10599);
nor U11393 (N_11393,N_10867,N_10558);
xnor U11394 (N_11394,N_10786,N_10598);
or U11395 (N_11395,N_10518,N_10548);
nor U11396 (N_11396,N_10969,N_10589);
nand U11397 (N_11397,N_10663,N_10661);
nor U11398 (N_11398,N_10564,N_10905);
xnor U11399 (N_11399,N_10982,N_10992);
nor U11400 (N_11400,N_10642,N_10849);
nor U11401 (N_11401,N_10547,N_10877);
or U11402 (N_11402,N_10608,N_10873);
or U11403 (N_11403,N_10736,N_10608);
nor U11404 (N_11404,N_10610,N_10594);
or U11405 (N_11405,N_10750,N_10714);
and U11406 (N_11406,N_10534,N_10552);
nor U11407 (N_11407,N_10871,N_10665);
nand U11408 (N_11408,N_10984,N_10681);
xnor U11409 (N_11409,N_10694,N_10758);
or U11410 (N_11410,N_10914,N_10965);
xor U11411 (N_11411,N_10731,N_10601);
nand U11412 (N_11412,N_10663,N_10923);
nor U11413 (N_11413,N_10696,N_10631);
or U11414 (N_11414,N_10771,N_10871);
or U11415 (N_11415,N_10814,N_10768);
nor U11416 (N_11416,N_10991,N_10605);
and U11417 (N_11417,N_10584,N_10849);
and U11418 (N_11418,N_10574,N_10702);
and U11419 (N_11419,N_10601,N_10711);
xnor U11420 (N_11420,N_10644,N_10670);
or U11421 (N_11421,N_10752,N_10578);
xnor U11422 (N_11422,N_10625,N_10528);
xnor U11423 (N_11423,N_10552,N_10783);
and U11424 (N_11424,N_10622,N_10819);
xor U11425 (N_11425,N_10683,N_10586);
xnor U11426 (N_11426,N_10707,N_10973);
and U11427 (N_11427,N_10825,N_10868);
and U11428 (N_11428,N_10578,N_10934);
and U11429 (N_11429,N_10901,N_10702);
or U11430 (N_11430,N_10502,N_10530);
or U11431 (N_11431,N_10944,N_10507);
or U11432 (N_11432,N_10956,N_10756);
and U11433 (N_11433,N_10800,N_10723);
and U11434 (N_11434,N_10575,N_10664);
nand U11435 (N_11435,N_10542,N_10926);
or U11436 (N_11436,N_10559,N_10770);
and U11437 (N_11437,N_10883,N_10901);
nand U11438 (N_11438,N_10784,N_10924);
or U11439 (N_11439,N_10717,N_10727);
nor U11440 (N_11440,N_10716,N_10765);
or U11441 (N_11441,N_10533,N_10961);
xnor U11442 (N_11442,N_10755,N_10520);
and U11443 (N_11443,N_10800,N_10853);
or U11444 (N_11444,N_10759,N_10585);
or U11445 (N_11445,N_10914,N_10698);
nor U11446 (N_11446,N_10759,N_10907);
xor U11447 (N_11447,N_10963,N_10950);
or U11448 (N_11448,N_10595,N_10812);
or U11449 (N_11449,N_10660,N_10915);
xnor U11450 (N_11450,N_10956,N_10755);
xor U11451 (N_11451,N_10606,N_10963);
and U11452 (N_11452,N_10514,N_10866);
nand U11453 (N_11453,N_10953,N_10835);
or U11454 (N_11454,N_10808,N_10587);
nand U11455 (N_11455,N_10653,N_10978);
and U11456 (N_11456,N_10726,N_10501);
nand U11457 (N_11457,N_10855,N_10835);
nand U11458 (N_11458,N_10679,N_10882);
and U11459 (N_11459,N_10621,N_10654);
and U11460 (N_11460,N_10933,N_10774);
nand U11461 (N_11461,N_10880,N_10733);
nand U11462 (N_11462,N_10524,N_10891);
xor U11463 (N_11463,N_10577,N_10598);
nand U11464 (N_11464,N_10531,N_10991);
xor U11465 (N_11465,N_10535,N_10971);
nor U11466 (N_11466,N_10516,N_10939);
nor U11467 (N_11467,N_10766,N_10933);
and U11468 (N_11468,N_10854,N_10544);
or U11469 (N_11469,N_10648,N_10504);
nand U11470 (N_11470,N_10787,N_10654);
or U11471 (N_11471,N_10818,N_10580);
xnor U11472 (N_11472,N_10673,N_10565);
xnor U11473 (N_11473,N_10932,N_10982);
and U11474 (N_11474,N_10862,N_10674);
nor U11475 (N_11475,N_10709,N_10876);
or U11476 (N_11476,N_10681,N_10658);
nand U11477 (N_11477,N_10713,N_10515);
xnor U11478 (N_11478,N_10667,N_10646);
and U11479 (N_11479,N_10897,N_10984);
or U11480 (N_11480,N_10874,N_10593);
xor U11481 (N_11481,N_10609,N_10961);
nand U11482 (N_11482,N_10513,N_10748);
or U11483 (N_11483,N_10500,N_10856);
nand U11484 (N_11484,N_10767,N_10998);
nand U11485 (N_11485,N_10552,N_10818);
nor U11486 (N_11486,N_10724,N_10711);
and U11487 (N_11487,N_10936,N_10851);
xor U11488 (N_11488,N_10695,N_10692);
or U11489 (N_11489,N_10617,N_10762);
nand U11490 (N_11490,N_10690,N_10856);
xnor U11491 (N_11491,N_10748,N_10832);
and U11492 (N_11492,N_10764,N_10558);
xnor U11493 (N_11493,N_10619,N_10880);
xor U11494 (N_11494,N_10989,N_10672);
and U11495 (N_11495,N_10834,N_10759);
nand U11496 (N_11496,N_10551,N_10574);
xnor U11497 (N_11497,N_10752,N_10591);
nand U11498 (N_11498,N_10611,N_10954);
or U11499 (N_11499,N_10961,N_10708);
xnor U11500 (N_11500,N_11406,N_11413);
xnor U11501 (N_11501,N_11063,N_11030);
and U11502 (N_11502,N_11131,N_11258);
and U11503 (N_11503,N_11224,N_11174);
nor U11504 (N_11504,N_11033,N_11023);
or U11505 (N_11505,N_11261,N_11394);
or U11506 (N_11506,N_11075,N_11450);
xnor U11507 (N_11507,N_11299,N_11071);
xor U11508 (N_11508,N_11113,N_11485);
xor U11509 (N_11509,N_11247,N_11456);
nor U11510 (N_11510,N_11264,N_11214);
or U11511 (N_11511,N_11269,N_11370);
xnor U11512 (N_11512,N_11260,N_11137);
or U11513 (N_11513,N_11365,N_11418);
nand U11514 (N_11514,N_11132,N_11341);
nand U11515 (N_11515,N_11211,N_11375);
and U11516 (N_11516,N_11035,N_11128);
nand U11517 (N_11517,N_11164,N_11244);
nand U11518 (N_11518,N_11161,N_11354);
or U11519 (N_11519,N_11480,N_11422);
xnor U11520 (N_11520,N_11424,N_11009);
or U11521 (N_11521,N_11191,N_11398);
xor U11522 (N_11522,N_11109,N_11275);
nor U11523 (N_11523,N_11289,N_11445);
nor U11524 (N_11524,N_11078,N_11120);
nor U11525 (N_11525,N_11389,N_11439);
and U11526 (N_11526,N_11202,N_11136);
xnor U11527 (N_11527,N_11157,N_11265);
xnor U11528 (N_11528,N_11251,N_11072);
or U11529 (N_11529,N_11068,N_11471);
nor U11530 (N_11530,N_11163,N_11177);
xor U11531 (N_11531,N_11073,N_11401);
nand U11532 (N_11532,N_11205,N_11266);
and U11533 (N_11533,N_11383,N_11477);
nand U11534 (N_11534,N_11372,N_11219);
xnor U11535 (N_11535,N_11150,N_11476);
and U11536 (N_11536,N_11312,N_11399);
nand U11537 (N_11537,N_11494,N_11179);
nor U11538 (N_11538,N_11281,N_11434);
nand U11539 (N_11539,N_11192,N_11397);
or U11540 (N_11540,N_11454,N_11210);
and U11541 (N_11541,N_11180,N_11327);
nor U11542 (N_11542,N_11472,N_11149);
xnor U11543 (N_11543,N_11252,N_11029);
xnor U11544 (N_11544,N_11402,N_11085);
or U11545 (N_11545,N_11465,N_11081);
xnor U11546 (N_11546,N_11070,N_11390);
xor U11547 (N_11547,N_11377,N_11475);
or U11548 (N_11548,N_11012,N_11206);
nand U11549 (N_11549,N_11011,N_11355);
nand U11550 (N_11550,N_11395,N_11067);
nand U11551 (N_11551,N_11125,N_11162);
xnor U11552 (N_11552,N_11057,N_11301);
nor U11553 (N_11553,N_11404,N_11169);
or U11554 (N_11554,N_11133,N_11259);
xor U11555 (N_11555,N_11138,N_11117);
xnor U11556 (N_11556,N_11099,N_11015);
nor U11557 (N_11557,N_11140,N_11385);
xor U11558 (N_11558,N_11311,N_11044);
and U11559 (N_11559,N_11280,N_11022);
nand U11560 (N_11560,N_11444,N_11055);
or U11561 (N_11561,N_11061,N_11184);
xor U11562 (N_11562,N_11178,N_11342);
xor U11563 (N_11563,N_11426,N_11145);
and U11564 (N_11564,N_11076,N_11353);
xnor U11565 (N_11565,N_11089,N_11487);
and U11566 (N_11566,N_11446,N_11302);
nand U11567 (N_11567,N_11499,N_11348);
or U11568 (N_11568,N_11069,N_11026);
xnor U11569 (N_11569,N_11002,N_11285);
nand U11570 (N_11570,N_11440,N_11196);
nor U11571 (N_11571,N_11245,N_11159);
and U11572 (N_11572,N_11139,N_11378);
xor U11573 (N_11573,N_11351,N_11154);
nand U11574 (N_11574,N_11229,N_11241);
or U11575 (N_11575,N_11168,N_11306);
nor U11576 (N_11576,N_11239,N_11336);
and U11577 (N_11577,N_11482,N_11451);
and U11578 (N_11578,N_11103,N_11056);
or U11579 (N_11579,N_11237,N_11236);
nor U11580 (N_11580,N_11101,N_11277);
and U11581 (N_11581,N_11282,N_11432);
xnor U11582 (N_11582,N_11193,N_11200);
xnor U11583 (N_11583,N_11134,N_11121);
and U11584 (N_11584,N_11442,N_11144);
nor U11585 (N_11585,N_11469,N_11235);
nor U11586 (N_11586,N_11151,N_11318);
nor U11587 (N_11587,N_11189,N_11340);
xor U11588 (N_11588,N_11291,N_11333);
nand U11589 (N_11589,N_11024,N_11160);
nor U11590 (N_11590,N_11123,N_11077);
nor U11591 (N_11591,N_11428,N_11010);
nand U11592 (N_11592,N_11152,N_11489);
xnor U11593 (N_11593,N_11062,N_11111);
xnor U11594 (N_11594,N_11021,N_11335);
or U11595 (N_11595,N_11004,N_11367);
nand U11596 (N_11596,N_11104,N_11127);
nand U11597 (N_11597,N_11126,N_11091);
nor U11598 (N_11598,N_11276,N_11330);
xnor U11599 (N_11599,N_11158,N_11000);
nand U11600 (N_11600,N_11412,N_11212);
and U11601 (N_11601,N_11182,N_11305);
nand U11602 (N_11602,N_11461,N_11097);
nor U11603 (N_11603,N_11334,N_11052);
and U11604 (N_11604,N_11246,N_11037);
or U11605 (N_11605,N_11018,N_11014);
nor U11606 (N_11606,N_11243,N_11118);
xnor U11607 (N_11607,N_11059,N_11387);
nand U11608 (N_11608,N_11005,N_11453);
nor U11609 (N_11609,N_11356,N_11462);
and U11610 (N_11610,N_11034,N_11408);
nor U11611 (N_11611,N_11230,N_11329);
nand U11612 (N_11612,N_11352,N_11017);
xor U11613 (N_11613,N_11087,N_11204);
nor U11614 (N_11614,N_11359,N_11064);
and U11615 (N_11615,N_11298,N_11316);
nand U11616 (N_11616,N_11382,N_11092);
nand U11617 (N_11617,N_11185,N_11242);
nor U11618 (N_11618,N_11488,N_11106);
nor U11619 (N_11619,N_11484,N_11297);
and U11620 (N_11620,N_11031,N_11095);
xor U11621 (N_11621,N_11107,N_11082);
xor U11622 (N_11622,N_11054,N_11415);
xor U11623 (N_11623,N_11218,N_11373);
and U11624 (N_11624,N_11114,N_11047);
nor U11625 (N_11625,N_11094,N_11400);
nor U11626 (N_11626,N_11008,N_11195);
or U11627 (N_11627,N_11417,N_11319);
or U11628 (N_11628,N_11098,N_11284);
nor U11629 (N_11629,N_11328,N_11437);
or U11630 (N_11630,N_11310,N_11255);
nor U11631 (N_11631,N_11083,N_11048);
nand U11632 (N_11632,N_11040,N_11001);
nand U11633 (N_11633,N_11074,N_11429);
and U11634 (N_11634,N_11420,N_11080);
xnor U11635 (N_11635,N_11197,N_11391);
nor U11636 (N_11636,N_11436,N_11096);
and U11637 (N_11637,N_11240,N_11231);
nor U11638 (N_11638,N_11248,N_11115);
nor U11639 (N_11639,N_11238,N_11172);
and U11640 (N_11640,N_11303,N_11495);
or U11641 (N_11641,N_11452,N_11129);
nand U11642 (N_11642,N_11227,N_11038);
and U11643 (N_11643,N_11286,N_11209);
and U11644 (N_11644,N_11287,N_11483);
xor U11645 (N_11645,N_11345,N_11296);
nand U11646 (N_11646,N_11143,N_11225);
and U11647 (N_11647,N_11166,N_11350);
nor U11648 (N_11648,N_11339,N_11267);
or U11649 (N_11649,N_11498,N_11376);
or U11650 (N_11650,N_11105,N_11006);
nand U11651 (N_11651,N_11213,N_11234);
nand U11652 (N_11652,N_11215,N_11226);
or U11653 (N_11653,N_11381,N_11438);
xnor U11654 (N_11654,N_11308,N_11183);
nor U11655 (N_11655,N_11388,N_11043);
xnor U11656 (N_11656,N_11254,N_11490);
or U11657 (N_11657,N_11407,N_11186);
xnor U11658 (N_11658,N_11263,N_11039);
xor U11659 (N_11659,N_11250,N_11171);
nor U11660 (N_11660,N_11141,N_11188);
and U11661 (N_11661,N_11435,N_11481);
or U11662 (N_11662,N_11416,N_11496);
or U11663 (N_11663,N_11216,N_11156);
nor U11664 (N_11664,N_11042,N_11016);
and U11665 (N_11665,N_11320,N_11199);
or U11666 (N_11666,N_11307,N_11368);
xor U11667 (N_11667,N_11463,N_11155);
nor U11668 (N_11668,N_11020,N_11116);
xor U11669 (N_11669,N_11201,N_11363);
or U11670 (N_11670,N_11272,N_11173);
nand U11671 (N_11671,N_11338,N_11380);
nor U11672 (N_11672,N_11403,N_11142);
or U11673 (N_11673,N_11146,N_11025);
or U11674 (N_11674,N_11423,N_11223);
or U11675 (N_11675,N_11324,N_11474);
and U11676 (N_11676,N_11203,N_11271);
nand U11677 (N_11677,N_11364,N_11460);
xnor U11678 (N_11678,N_11135,N_11253);
nand U11679 (N_11679,N_11392,N_11222);
nand U11680 (N_11680,N_11433,N_11396);
and U11681 (N_11681,N_11467,N_11362);
or U11682 (N_11682,N_11295,N_11148);
nor U11683 (N_11683,N_11466,N_11332);
nor U11684 (N_11684,N_11233,N_11268);
or U11685 (N_11685,N_11110,N_11053);
nand U11686 (N_11686,N_11283,N_11405);
and U11687 (N_11687,N_11491,N_11130);
nand U11688 (N_11688,N_11321,N_11292);
or U11689 (N_11689,N_11019,N_11084);
nor U11690 (N_11690,N_11100,N_11322);
nand U11691 (N_11691,N_11419,N_11288);
nor U11692 (N_11692,N_11293,N_11486);
and U11693 (N_11693,N_11430,N_11331);
or U11694 (N_11694,N_11256,N_11358);
nand U11695 (N_11695,N_11273,N_11167);
and U11696 (N_11696,N_11366,N_11190);
and U11697 (N_11697,N_11041,N_11431);
nand U11698 (N_11698,N_11361,N_11479);
and U11699 (N_11699,N_11176,N_11379);
xor U11700 (N_11700,N_11497,N_11217);
nand U11701 (N_11701,N_11360,N_11347);
or U11702 (N_11702,N_11349,N_11386);
and U11703 (N_11703,N_11410,N_11045);
xor U11704 (N_11704,N_11220,N_11198);
and U11705 (N_11705,N_11300,N_11175);
xor U11706 (N_11706,N_11313,N_11086);
and U11707 (N_11707,N_11343,N_11257);
xor U11708 (N_11708,N_11421,N_11443);
nand U11709 (N_11709,N_11208,N_11065);
nor U11710 (N_11710,N_11270,N_11409);
nor U11711 (N_11711,N_11414,N_11007);
nor U11712 (N_11712,N_11032,N_11337);
or U11713 (N_11713,N_11393,N_11051);
nand U11714 (N_11714,N_11459,N_11278);
or U11715 (N_11715,N_11108,N_11262);
nor U11716 (N_11716,N_11448,N_11228);
nand U11717 (N_11717,N_11124,N_11207);
xnor U11718 (N_11718,N_11425,N_11112);
or U11719 (N_11719,N_11036,N_11027);
nor U11720 (N_11720,N_11493,N_11279);
and U11721 (N_11721,N_11165,N_11079);
nor U11722 (N_11722,N_11384,N_11003);
nor U11723 (N_11723,N_11468,N_11411);
or U11724 (N_11724,N_11427,N_11371);
nor U11725 (N_11725,N_11447,N_11317);
nand U11726 (N_11726,N_11464,N_11357);
nand U11727 (N_11727,N_11323,N_11441);
xor U11728 (N_11728,N_11315,N_11093);
nor U11729 (N_11729,N_11232,N_11374);
nand U11730 (N_11730,N_11290,N_11013);
and U11731 (N_11731,N_11049,N_11470);
or U11732 (N_11732,N_11325,N_11119);
nand U11733 (N_11733,N_11478,N_11457);
or U11734 (N_11734,N_11088,N_11187);
nor U11735 (N_11735,N_11102,N_11050);
xor U11736 (N_11736,N_11181,N_11309);
xor U11737 (N_11737,N_11060,N_11028);
xor U11738 (N_11738,N_11046,N_11066);
or U11739 (N_11739,N_11294,N_11249);
nor U11740 (N_11740,N_11458,N_11369);
or U11741 (N_11741,N_11170,N_11326);
and U11742 (N_11742,N_11147,N_11221);
or U11743 (N_11743,N_11346,N_11473);
nand U11744 (N_11744,N_11449,N_11492);
or U11745 (N_11745,N_11274,N_11194);
nor U11746 (N_11746,N_11304,N_11344);
or U11747 (N_11747,N_11058,N_11314);
nor U11748 (N_11748,N_11153,N_11122);
or U11749 (N_11749,N_11090,N_11455);
xor U11750 (N_11750,N_11391,N_11215);
or U11751 (N_11751,N_11327,N_11427);
and U11752 (N_11752,N_11016,N_11256);
xnor U11753 (N_11753,N_11412,N_11441);
nand U11754 (N_11754,N_11024,N_11000);
nor U11755 (N_11755,N_11218,N_11264);
nor U11756 (N_11756,N_11351,N_11482);
nand U11757 (N_11757,N_11134,N_11323);
or U11758 (N_11758,N_11152,N_11132);
nor U11759 (N_11759,N_11279,N_11312);
xnor U11760 (N_11760,N_11120,N_11071);
nor U11761 (N_11761,N_11122,N_11405);
nor U11762 (N_11762,N_11457,N_11191);
nand U11763 (N_11763,N_11322,N_11159);
nand U11764 (N_11764,N_11365,N_11170);
xnor U11765 (N_11765,N_11109,N_11128);
xor U11766 (N_11766,N_11265,N_11481);
and U11767 (N_11767,N_11115,N_11010);
xnor U11768 (N_11768,N_11185,N_11356);
xor U11769 (N_11769,N_11241,N_11201);
xor U11770 (N_11770,N_11306,N_11330);
or U11771 (N_11771,N_11079,N_11058);
xor U11772 (N_11772,N_11192,N_11070);
nand U11773 (N_11773,N_11085,N_11229);
and U11774 (N_11774,N_11470,N_11246);
or U11775 (N_11775,N_11176,N_11340);
nor U11776 (N_11776,N_11063,N_11276);
and U11777 (N_11777,N_11487,N_11366);
nor U11778 (N_11778,N_11471,N_11320);
nor U11779 (N_11779,N_11195,N_11060);
and U11780 (N_11780,N_11199,N_11009);
and U11781 (N_11781,N_11124,N_11487);
nor U11782 (N_11782,N_11068,N_11322);
nor U11783 (N_11783,N_11082,N_11025);
nand U11784 (N_11784,N_11144,N_11170);
nand U11785 (N_11785,N_11409,N_11284);
xnor U11786 (N_11786,N_11158,N_11269);
nor U11787 (N_11787,N_11193,N_11272);
and U11788 (N_11788,N_11030,N_11311);
xnor U11789 (N_11789,N_11270,N_11016);
xnor U11790 (N_11790,N_11440,N_11122);
nand U11791 (N_11791,N_11012,N_11128);
xor U11792 (N_11792,N_11458,N_11257);
or U11793 (N_11793,N_11475,N_11421);
xnor U11794 (N_11794,N_11346,N_11077);
xor U11795 (N_11795,N_11065,N_11075);
or U11796 (N_11796,N_11469,N_11312);
xnor U11797 (N_11797,N_11277,N_11170);
xnor U11798 (N_11798,N_11451,N_11155);
nor U11799 (N_11799,N_11226,N_11403);
and U11800 (N_11800,N_11147,N_11367);
nor U11801 (N_11801,N_11035,N_11152);
or U11802 (N_11802,N_11079,N_11222);
nor U11803 (N_11803,N_11256,N_11219);
nor U11804 (N_11804,N_11018,N_11348);
nand U11805 (N_11805,N_11054,N_11475);
and U11806 (N_11806,N_11013,N_11037);
nand U11807 (N_11807,N_11347,N_11416);
xor U11808 (N_11808,N_11105,N_11157);
nor U11809 (N_11809,N_11112,N_11198);
nor U11810 (N_11810,N_11266,N_11420);
and U11811 (N_11811,N_11456,N_11237);
xor U11812 (N_11812,N_11230,N_11007);
or U11813 (N_11813,N_11053,N_11075);
and U11814 (N_11814,N_11153,N_11037);
xnor U11815 (N_11815,N_11178,N_11072);
xor U11816 (N_11816,N_11255,N_11279);
xor U11817 (N_11817,N_11363,N_11487);
or U11818 (N_11818,N_11058,N_11383);
nor U11819 (N_11819,N_11002,N_11008);
or U11820 (N_11820,N_11329,N_11104);
nor U11821 (N_11821,N_11496,N_11183);
nor U11822 (N_11822,N_11084,N_11201);
xnor U11823 (N_11823,N_11191,N_11166);
nand U11824 (N_11824,N_11342,N_11096);
nand U11825 (N_11825,N_11141,N_11366);
xor U11826 (N_11826,N_11428,N_11435);
and U11827 (N_11827,N_11344,N_11162);
and U11828 (N_11828,N_11248,N_11313);
nor U11829 (N_11829,N_11016,N_11332);
xor U11830 (N_11830,N_11165,N_11376);
and U11831 (N_11831,N_11477,N_11158);
and U11832 (N_11832,N_11437,N_11333);
xor U11833 (N_11833,N_11210,N_11354);
or U11834 (N_11834,N_11327,N_11489);
xor U11835 (N_11835,N_11362,N_11444);
nor U11836 (N_11836,N_11321,N_11367);
nor U11837 (N_11837,N_11425,N_11474);
or U11838 (N_11838,N_11239,N_11287);
xnor U11839 (N_11839,N_11234,N_11340);
or U11840 (N_11840,N_11425,N_11091);
nor U11841 (N_11841,N_11354,N_11076);
nor U11842 (N_11842,N_11363,N_11465);
xor U11843 (N_11843,N_11454,N_11353);
xnor U11844 (N_11844,N_11248,N_11369);
or U11845 (N_11845,N_11265,N_11053);
xnor U11846 (N_11846,N_11017,N_11307);
nor U11847 (N_11847,N_11369,N_11487);
nor U11848 (N_11848,N_11057,N_11239);
nand U11849 (N_11849,N_11264,N_11186);
nand U11850 (N_11850,N_11304,N_11155);
and U11851 (N_11851,N_11023,N_11360);
nor U11852 (N_11852,N_11076,N_11452);
and U11853 (N_11853,N_11090,N_11279);
and U11854 (N_11854,N_11435,N_11462);
xor U11855 (N_11855,N_11284,N_11225);
nor U11856 (N_11856,N_11380,N_11337);
xor U11857 (N_11857,N_11084,N_11004);
xnor U11858 (N_11858,N_11126,N_11436);
xor U11859 (N_11859,N_11077,N_11133);
and U11860 (N_11860,N_11238,N_11071);
nor U11861 (N_11861,N_11186,N_11193);
nand U11862 (N_11862,N_11354,N_11245);
nand U11863 (N_11863,N_11319,N_11001);
xor U11864 (N_11864,N_11153,N_11291);
or U11865 (N_11865,N_11161,N_11134);
or U11866 (N_11866,N_11233,N_11440);
nand U11867 (N_11867,N_11445,N_11185);
or U11868 (N_11868,N_11118,N_11100);
and U11869 (N_11869,N_11168,N_11305);
xor U11870 (N_11870,N_11233,N_11460);
nand U11871 (N_11871,N_11092,N_11492);
xnor U11872 (N_11872,N_11011,N_11064);
and U11873 (N_11873,N_11050,N_11052);
or U11874 (N_11874,N_11159,N_11081);
nand U11875 (N_11875,N_11157,N_11099);
or U11876 (N_11876,N_11414,N_11221);
and U11877 (N_11877,N_11341,N_11328);
or U11878 (N_11878,N_11386,N_11088);
or U11879 (N_11879,N_11157,N_11236);
nand U11880 (N_11880,N_11331,N_11151);
nor U11881 (N_11881,N_11495,N_11186);
nor U11882 (N_11882,N_11219,N_11375);
nand U11883 (N_11883,N_11015,N_11043);
nand U11884 (N_11884,N_11143,N_11042);
nand U11885 (N_11885,N_11044,N_11411);
xor U11886 (N_11886,N_11353,N_11462);
and U11887 (N_11887,N_11171,N_11452);
and U11888 (N_11888,N_11309,N_11472);
and U11889 (N_11889,N_11030,N_11023);
xor U11890 (N_11890,N_11462,N_11184);
or U11891 (N_11891,N_11026,N_11470);
or U11892 (N_11892,N_11161,N_11206);
nand U11893 (N_11893,N_11141,N_11275);
nor U11894 (N_11894,N_11003,N_11374);
xnor U11895 (N_11895,N_11163,N_11320);
nor U11896 (N_11896,N_11441,N_11276);
nor U11897 (N_11897,N_11243,N_11205);
or U11898 (N_11898,N_11360,N_11027);
and U11899 (N_11899,N_11189,N_11265);
nor U11900 (N_11900,N_11014,N_11387);
and U11901 (N_11901,N_11056,N_11004);
and U11902 (N_11902,N_11424,N_11180);
and U11903 (N_11903,N_11317,N_11245);
xnor U11904 (N_11904,N_11166,N_11087);
nor U11905 (N_11905,N_11254,N_11466);
or U11906 (N_11906,N_11173,N_11286);
nand U11907 (N_11907,N_11392,N_11061);
or U11908 (N_11908,N_11243,N_11021);
or U11909 (N_11909,N_11197,N_11459);
and U11910 (N_11910,N_11281,N_11460);
nand U11911 (N_11911,N_11185,N_11497);
nor U11912 (N_11912,N_11490,N_11444);
nor U11913 (N_11913,N_11358,N_11363);
and U11914 (N_11914,N_11409,N_11443);
xnor U11915 (N_11915,N_11315,N_11213);
and U11916 (N_11916,N_11302,N_11058);
nor U11917 (N_11917,N_11155,N_11084);
nand U11918 (N_11918,N_11017,N_11234);
or U11919 (N_11919,N_11218,N_11121);
xor U11920 (N_11920,N_11391,N_11012);
and U11921 (N_11921,N_11429,N_11065);
or U11922 (N_11922,N_11324,N_11088);
nand U11923 (N_11923,N_11059,N_11423);
or U11924 (N_11924,N_11420,N_11460);
or U11925 (N_11925,N_11394,N_11061);
nand U11926 (N_11926,N_11144,N_11178);
nor U11927 (N_11927,N_11485,N_11323);
or U11928 (N_11928,N_11144,N_11382);
xnor U11929 (N_11929,N_11205,N_11193);
nor U11930 (N_11930,N_11141,N_11434);
and U11931 (N_11931,N_11380,N_11075);
xnor U11932 (N_11932,N_11471,N_11005);
xor U11933 (N_11933,N_11282,N_11038);
nand U11934 (N_11934,N_11232,N_11388);
xor U11935 (N_11935,N_11096,N_11071);
and U11936 (N_11936,N_11217,N_11479);
nor U11937 (N_11937,N_11124,N_11390);
or U11938 (N_11938,N_11409,N_11106);
and U11939 (N_11939,N_11371,N_11470);
or U11940 (N_11940,N_11202,N_11331);
nand U11941 (N_11941,N_11373,N_11420);
nor U11942 (N_11942,N_11142,N_11123);
xor U11943 (N_11943,N_11022,N_11431);
or U11944 (N_11944,N_11095,N_11025);
nand U11945 (N_11945,N_11404,N_11036);
and U11946 (N_11946,N_11156,N_11324);
xnor U11947 (N_11947,N_11212,N_11080);
nand U11948 (N_11948,N_11355,N_11041);
xor U11949 (N_11949,N_11312,N_11334);
nor U11950 (N_11950,N_11191,N_11306);
and U11951 (N_11951,N_11330,N_11425);
nor U11952 (N_11952,N_11045,N_11194);
nor U11953 (N_11953,N_11015,N_11228);
nor U11954 (N_11954,N_11278,N_11497);
nand U11955 (N_11955,N_11143,N_11098);
nor U11956 (N_11956,N_11175,N_11097);
or U11957 (N_11957,N_11067,N_11029);
xor U11958 (N_11958,N_11452,N_11423);
xor U11959 (N_11959,N_11091,N_11403);
nor U11960 (N_11960,N_11315,N_11096);
nand U11961 (N_11961,N_11085,N_11422);
or U11962 (N_11962,N_11438,N_11196);
and U11963 (N_11963,N_11490,N_11493);
xnor U11964 (N_11964,N_11492,N_11421);
and U11965 (N_11965,N_11238,N_11433);
and U11966 (N_11966,N_11227,N_11116);
nor U11967 (N_11967,N_11059,N_11483);
nor U11968 (N_11968,N_11430,N_11208);
nand U11969 (N_11969,N_11393,N_11364);
xor U11970 (N_11970,N_11344,N_11190);
nand U11971 (N_11971,N_11390,N_11359);
or U11972 (N_11972,N_11127,N_11453);
nand U11973 (N_11973,N_11174,N_11142);
nor U11974 (N_11974,N_11437,N_11080);
xnor U11975 (N_11975,N_11094,N_11190);
nor U11976 (N_11976,N_11052,N_11145);
xor U11977 (N_11977,N_11395,N_11446);
or U11978 (N_11978,N_11120,N_11133);
or U11979 (N_11979,N_11057,N_11326);
nor U11980 (N_11980,N_11021,N_11283);
xnor U11981 (N_11981,N_11442,N_11213);
nor U11982 (N_11982,N_11045,N_11235);
and U11983 (N_11983,N_11080,N_11126);
xnor U11984 (N_11984,N_11249,N_11361);
xnor U11985 (N_11985,N_11177,N_11076);
or U11986 (N_11986,N_11417,N_11151);
and U11987 (N_11987,N_11292,N_11166);
nor U11988 (N_11988,N_11270,N_11492);
or U11989 (N_11989,N_11494,N_11031);
and U11990 (N_11990,N_11476,N_11303);
xnor U11991 (N_11991,N_11311,N_11266);
nor U11992 (N_11992,N_11261,N_11103);
xnor U11993 (N_11993,N_11113,N_11358);
xnor U11994 (N_11994,N_11242,N_11353);
and U11995 (N_11995,N_11005,N_11223);
and U11996 (N_11996,N_11156,N_11319);
or U11997 (N_11997,N_11111,N_11298);
or U11998 (N_11998,N_11146,N_11484);
nor U11999 (N_11999,N_11188,N_11273);
nand U12000 (N_12000,N_11694,N_11989);
xnor U12001 (N_12001,N_11777,N_11759);
and U12002 (N_12002,N_11839,N_11923);
nand U12003 (N_12003,N_11802,N_11710);
nand U12004 (N_12004,N_11747,N_11665);
nor U12005 (N_12005,N_11737,N_11591);
xnor U12006 (N_12006,N_11980,N_11684);
xnor U12007 (N_12007,N_11798,N_11683);
and U12008 (N_12008,N_11557,N_11960);
or U12009 (N_12009,N_11616,N_11919);
nor U12010 (N_12010,N_11744,N_11827);
or U12011 (N_12011,N_11635,N_11644);
or U12012 (N_12012,N_11696,N_11812);
nand U12013 (N_12013,N_11536,N_11745);
nor U12014 (N_12014,N_11817,N_11664);
nand U12015 (N_12015,N_11995,N_11614);
xor U12016 (N_12016,N_11996,N_11815);
or U12017 (N_12017,N_11717,N_11908);
or U12018 (N_12018,N_11766,N_11903);
nor U12019 (N_12019,N_11695,N_11970);
nor U12020 (N_12020,N_11537,N_11951);
and U12021 (N_12021,N_11879,N_11752);
and U12022 (N_12022,N_11973,N_11599);
nand U12023 (N_12023,N_11533,N_11531);
and U12024 (N_12024,N_11921,N_11966);
xor U12025 (N_12025,N_11846,N_11841);
xnor U12026 (N_12026,N_11623,N_11539);
and U12027 (N_12027,N_11613,N_11610);
and U12028 (N_12028,N_11668,N_11965);
nand U12029 (N_12029,N_11767,N_11911);
nor U12030 (N_12030,N_11605,N_11715);
and U12031 (N_12031,N_11530,N_11809);
or U12032 (N_12032,N_11849,N_11749);
xor U12033 (N_12033,N_11576,N_11918);
and U12034 (N_12034,N_11865,N_11594);
and U12035 (N_12035,N_11667,N_11579);
nand U12036 (N_12036,N_11993,N_11905);
nor U12037 (N_12037,N_11520,N_11940);
nor U12038 (N_12038,N_11816,N_11988);
xor U12039 (N_12039,N_11932,N_11915);
xnor U12040 (N_12040,N_11731,N_11834);
xnor U12041 (N_12041,N_11638,N_11859);
nor U12042 (N_12042,N_11885,N_11856);
and U12043 (N_12043,N_11652,N_11748);
and U12044 (N_12044,N_11511,N_11897);
and U12045 (N_12045,N_11831,N_11840);
or U12046 (N_12046,N_11852,N_11850);
nand U12047 (N_12047,N_11626,N_11714);
nand U12048 (N_12048,N_11797,N_11545);
xnor U12049 (N_12049,N_11874,N_11528);
xnor U12050 (N_12050,N_11627,N_11888);
nor U12051 (N_12051,N_11880,N_11632);
and U12052 (N_12052,N_11851,N_11527);
xor U12053 (N_12053,N_11907,N_11863);
nand U12054 (N_12054,N_11822,N_11588);
or U12055 (N_12055,N_11678,N_11983);
or U12056 (N_12056,N_11976,N_11990);
and U12057 (N_12057,N_11725,N_11937);
nor U12058 (N_12058,N_11743,N_11611);
xor U12059 (N_12059,N_11758,N_11895);
nor U12060 (N_12060,N_11843,N_11524);
xor U12061 (N_12061,N_11833,N_11786);
xnor U12062 (N_12062,N_11728,N_11691);
nor U12063 (N_12063,N_11662,N_11569);
nand U12064 (N_12064,N_11942,N_11708);
xor U12065 (N_12065,N_11969,N_11826);
and U12066 (N_12066,N_11663,N_11686);
or U12067 (N_12067,N_11509,N_11986);
xor U12068 (N_12068,N_11901,N_11543);
xnor U12069 (N_12069,N_11886,N_11941);
or U12070 (N_12070,N_11582,N_11612);
and U12071 (N_12071,N_11808,N_11900);
xor U12072 (N_12072,N_11596,N_11754);
and U12073 (N_12073,N_11603,N_11974);
nand U12074 (N_12074,N_11649,N_11726);
xor U12075 (N_12075,N_11924,N_11514);
nor U12076 (N_12076,N_11971,N_11523);
nor U12077 (N_12077,N_11930,N_11598);
xnor U12078 (N_12078,N_11707,N_11950);
xnor U12079 (N_12079,N_11604,N_11813);
nor U12080 (N_12080,N_11791,N_11790);
nand U12081 (N_12081,N_11674,N_11853);
nand U12082 (N_12082,N_11732,N_11875);
or U12083 (N_12083,N_11997,N_11553);
or U12084 (N_12084,N_11929,N_11653);
nand U12085 (N_12085,N_11884,N_11904);
nand U12086 (N_12086,N_11820,N_11967);
nor U12087 (N_12087,N_11621,N_11920);
or U12088 (N_12088,N_11981,N_11586);
nor U12089 (N_12089,N_11757,N_11535);
and U12090 (N_12090,N_11890,N_11887);
nand U12091 (N_12091,N_11963,N_11525);
xor U12092 (N_12092,N_11669,N_11682);
and U12093 (N_12093,N_11538,N_11810);
nand U12094 (N_12094,N_11985,N_11595);
nand U12095 (N_12095,N_11589,N_11512);
xor U12096 (N_12096,N_11601,N_11609);
xnor U12097 (N_12097,N_11938,N_11837);
and U12098 (N_12098,N_11871,N_11736);
nand U12099 (N_12099,N_11657,N_11581);
xor U12100 (N_12100,N_11824,N_11804);
or U12101 (N_12101,N_11975,N_11584);
nor U12102 (N_12102,N_11642,N_11753);
xnor U12103 (N_12103,N_11671,N_11593);
or U12104 (N_12104,N_11898,N_11585);
and U12105 (N_12105,N_11892,N_11519);
nor U12106 (N_12106,N_11639,N_11624);
nand U12107 (N_12107,N_11948,N_11724);
nor U12108 (N_12108,N_11935,N_11700);
and U12109 (N_12109,N_11855,N_11739);
nand U12110 (N_12110,N_11946,N_11910);
and U12111 (N_12111,N_11869,N_11699);
xnor U12112 (N_12112,N_11751,N_11836);
or U12113 (N_12113,N_11704,N_11858);
xor U12114 (N_12114,N_11636,N_11505);
nor U12115 (N_12115,N_11517,N_11829);
nor U12116 (N_12116,N_11814,N_11733);
and U12117 (N_12117,N_11574,N_11881);
nor U12118 (N_12118,N_11701,N_11998);
xnor U12119 (N_12119,N_11568,N_11977);
xnor U12120 (N_12120,N_11648,N_11830);
xnor U12121 (N_12121,N_11825,N_11508);
nor U12122 (N_12122,N_11534,N_11796);
nor U12123 (N_12123,N_11987,N_11925);
and U12124 (N_12124,N_11868,N_11779);
and U12125 (N_12125,N_11718,N_11952);
nand U12126 (N_12126,N_11793,N_11775);
or U12127 (N_12127,N_11558,N_11672);
nand U12128 (N_12128,N_11711,N_11773);
xnor U12129 (N_12129,N_11556,N_11734);
nor U12130 (N_12130,N_11522,N_11552);
or U12131 (N_12131,N_11889,N_11572);
and U12132 (N_12132,N_11761,N_11764);
xnor U12133 (N_12133,N_11961,N_11554);
xnor U12134 (N_12134,N_11955,N_11646);
or U12135 (N_12135,N_11742,N_11746);
nor U12136 (N_12136,N_11618,N_11762);
nor U12137 (N_12137,N_11573,N_11620);
xor U12138 (N_12138,N_11789,N_11550);
nor U12139 (N_12139,N_11785,N_11735);
or U12140 (N_12140,N_11803,N_11756);
and U12141 (N_12141,N_11953,N_11799);
nand U12142 (N_12142,N_11872,N_11811);
or U12143 (N_12143,N_11931,N_11782);
or U12144 (N_12144,N_11540,N_11592);
nor U12145 (N_12145,N_11565,N_11992);
nor U12146 (N_12146,N_11567,N_11962);
nor U12147 (N_12147,N_11628,N_11654);
nand U12148 (N_12148,N_11821,N_11548);
and U12149 (N_12149,N_11771,N_11544);
xor U12150 (N_12150,N_11689,N_11763);
and U12151 (N_12151,N_11956,N_11641);
nand U12152 (N_12152,N_11882,N_11702);
nand U12153 (N_12153,N_11549,N_11651);
or U12154 (N_12154,N_11954,N_11631);
nor U12155 (N_12155,N_11619,N_11894);
nor U12156 (N_12156,N_11560,N_11828);
xor U12157 (N_12157,N_11891,N_11949);
or U12158 (N_12158,N_11916,N_11561);
and U12159 (N_12159,N_11706,N_11640);
or U12160 (N_12160,N_11500,N_11661);
nand U12161 (N_12161,N_11692,N_11806);
and U12162 (N_12162,N_11541,N_11778);
and U12163 (N_12163,N_11917,N_11577);
nand U12164 (N_12164,N_11656,N_11842);
nand U12165 (N_12165,N_11801,N_11555);
nand U12166 (N_12166,N_11794,N_11795);
or U12167 (N_12167,N_11617,N_11713);
nor U12168 (N_12168,N_11502,N_11835);
or U12169 (N_12169,N_11964,N_11741);
or U12170 (N_12170,N_11784,N_11673);
nor U12171 (N_12171,N_11501,N_11647);
or U12172 (N_12172,N_11906,N_11518);
nand U12173 (N_12173,N_11503,N_11625);
nor U12174 (N_12174,N_11608,N_11727);
or U12175 (N_12175,N_11755,N_11781);
and U12176 (N_12176,N_11650,N_11685);
nand U12177 (N_12177,N_11721,N_11629);
nor U12178 (N_12178,N_11877,N_11902);
nand U12179 (N_12179,N_11847,N_11670);
and U12180 (N_12180,N_11690,N_11587);
nand U12181 (N_12181,N_11959,N_11972);
nand U12182 (N_12182,N_11909,N_11774);
nor U12183 (N_12183,N_11838,N_11848);
nand U12184 (N_12184,N_11760,N_11854);
nor U12185 (N_12185,N_11712,N_11643);
nor U12186 (N_12186,N_11860,N_11776);
nor U12187 (N_12187,N_11723,N_11697);
nor U12188 (N_12188,N_11547,N_11730);
and U12189 (N_12189,N_11866,N_11693);
nor U12190 (N_12190,N_11819,N_11947);
nor U12191 (N_12191,N_11677,N_11832);
xor U12192 (N_12192,N_11709,N_11637);
nand U12193 (N_12193,N_11958,N_11883);
nand U12194 (N_12194,N_11551,N_11783);
and U12195 (N_12195,N_11607,N_11633);
xnor U12196 (N_12196,N_11719,N_11676);
or U12197 (N_12197,N_11991,N_11562);
xor U12198 (N_12198,N_11563,N_11780);
xnor U12199 (N_12199,N_11893,N_11927);
or U12200 (N_12200,N_11590,N_11606);
or U12201 (N_12201,N_11688,N_11630);
nor U12202 (N_12202,N_11580,N_11666);
nand U12203 (N_12203,N_11729,N_11876);
nor U12204 (N_12204,N_11818,N_11716);
or U12205 (N_12205,N_11510,N_11571);
or U12206 (N_12206,N_11602,N_11957);
and U12207 (N_12207,N_11934,N_11750);
nand U12208 (N_12208,N_11945,N_11658);
and U12209 (N_12209,N_11979,N_11705);
and U12210 (N_12210,N_11765,N_11622);
and U12211 (N_12211,N_11655,N_11922);
xor U12212 (N_12212,N_11982,N_11660);
nand U12213 (N_12213,N_11870,N_11805);
xnor U12214 (N_12214,N_11800,N_11844);
nand U12215 (N_12215,N_11873,N_11994);
nand U12216 (N_12216,N_11845,N_11645);
xor U12217 (N_12217,N_11862,N_11740);
nand U12218 (N_12218,N_11615,N_11864);
xor U12219 (N_12219,N_11861,N_11529);
nor U12220 (N_12220,N_11807,N_11867);
and U12221 (N_12221,N_11738,N_11681);
nor U12222 (N_12222,N_11578,N_11526);
xor U12223 (N_12223,N_11720,N_11857);
nor U12224 (N_12224,N_11899,N_11597);
nor U12225 (N_12225,N_11772,N_11679);
nand U12226 (N_12226,N_11504,N_11698);
and U12227 (N_12227,N_11770,N_11566);
or U12228 (N_12228,N_11507,N_11546);
or U12229 (N_12229,N_11928,N_11943);
and U12230 (N_12230,N_11575,N_11926);
xor U12231 (N_12231,N_11687,N_11570);
or U12232 (N_12232,N_11680,N_11703);
nor U12233 (N_12233,N_11787,N_11978);
nor U12234 (N_12234,N_11914,N_11913);
nand U12235 (N_12235,N_11521,N_11999);
nand U12236 (N_12236,N_11722,N_11823);
and U12237 (N_12237,N_11600,N_11532);
and U12238 (N_12238,N_11769,N_11936);
or U12239 (N_12239,N_11792,N_11513);
xor U12240 (N_12240,N_11878,N_11768);
or U12241 (N_12241,N_11516,N_11944);
and U12242 (N_12242,N_11939,N_11968);
nand U12243 (N_12243,N_11788,N_11659);
nand U12244 (N_12244,N_11634,N_11559);
and U12245 (N_12245,N_11984,N_11583);
nand U12246 (N_12246,N_11896,N_11564);
or U12247 (N_12247,N_11506,N_11912);
nand U12248 (N_12248,N_11933,N_11542);
xnor U12249 (N_12249,N_11675,N_11515);
and U12250 (N_12250,N_11561,N_11641);
and U12251 (N_12251,N_11615,N_11598);
xor U12252 (N_12252,N_11763,N_11951);
and U12253 (N_12253,N_11786,N_11678);
nand U12254 (N_12254,N_11655,N_11617);
nor U12255 (N_12255,N_11862,N_11611);
and U12256 (N_12256,N_11898,N_11833);
or U12257 (N_12257,N_11825,N_11827);
nand U12258 (N_12258,N_11662,N_11537);
nor U12259 (N_12259,N_11578,N_11543);
or U12260 (N_12260,N_11633,N_11587);
nor U12261 (N_12261,N_11996,N_11898);
nor U12262 (N_12262,N_11808,N_11824);
or U12263 (N_12263,N_11774,N_11599);
nand U12264 (N_12264,N_11799,N_11981);
xor U12265 (N_12265,N_11775,N_11988);
xnor U12266 (N_12266,N_11765,N_11647);
nand U12267 (N_12267,N_11540,N_11607);
nor U12268 (N_12268,N_11659,N_11557);
nor U12269 (N_12269,N_11817,N_11549);
or U12270 (N_12270,N_11500,N_11640);
xor U12271 (N_12271,N_11584,N_11811);
xor U12272 (N_12272,N_11706,N_11650);
and U12273 (N_12273,N_11674,N_11511);
xnor U12274 (N_12274,N_11816,N_11863);
or U12275 (N_12275,N_11837,N_11583);
and U12276 (N_12276,N_11642,N_11802);
and U12277 (N_12277,N_11878,N_11555);
or U12278 (N_12278,N_11500,N_11783);
nand U12279 (N_12279,N_11698,N_11917);
or U12280 (N_12280,N_11655,N_11569);
or U12281 (N_12281,N_11556,N_11795);
or U12282 (N_12282,N_11702,N_11889);
nor U12283 (N_12283,N_11940,N_11606);
nand U12284 (N_12284,N_11749,N_11577);
nor U12285 (N_12285,N_11726,N_11601);
and U12286 (N_12286,N_11833,N_11820);
nand U12287 (N_12287,N_11926,N_11710);
xor U12288 (N_12288,N_11751,N_11970);
nand U12289 (N_12289,N_11657,N_11769);
and U12290 (N_12290,N_11614,N_11929);
xnor U12291 (N_12291,N_11626,N_11621);
and U12292 (N_12292,N_11889,N_11991);
nand U12293 (N_12293,N_11509,N_11669);
or U12294 (N_12294,N_11830,N_11517);
xnor U12295 (N_12295,N_11605,N_11657);
nor U12296 (N_12296,N_11804,N_11699);
nor U12297 (N_12297,N_11846,N_11691);
or U12298 (N_12298,N_11870,N_11551);
nand U12299 (N_12299,N_11733,N_11776);
and U12300 (N_12300,N_11882,N_11756);
and U12301 (N_12301,N_11630,N_11662);
xor U12302 (N_12302,N_11620,N_11585);
xnor U12303 (N_12303,N_11702,N_11660);
and U12304 (N_12304,N_11702,N_11760);
nand U12305 (N_12305,N_11959,N_11850);
and U12306 (N_12306,N_11971,N_11656);
and U12307 (N_12307,N_11597,N_11958);
nor U12308 (N_12308,N_11940,N_11808);
xnor U12309 (N_12309,N_11919,N_11501);
nor U12310 (N_12310,N_11697,N_11831);
nand U12311 (N_12311,N_11891,N_11579);
or U12312 (N_12312,N_11827,N_11838);
or U12313 (N_12313,N_11961,N_11800);
nand U12314 (N_12314,N_11770,N_11820);
and U12315 (N_12315,N_11947,N_11797);
xor U12316 (N_12316,N_11520,N_11938);
xor U12317 (N_12317,N_11581,N_11650);
or U12318 (N_12318,N_11649,N_11850);
nand U12319 (N_12319,N_11932,N_11606);
nand U12320 (N_12320,N_11610,N_11988);
and U12321 (N_12321,N_11543,N_11959);
or U12322 (N_12322,N_11773,N_11915);
nor U12323 (N_12323,N_11711,N_11826);
nor U12324 (N_12324,N_11500,N_11799);
nand U12325 (N_12325,N_11801,N_11837);
nor U12326 (N_12326,N_11931,N_11852);
xor U12327 (N_12327,N_11576,N_11833);
nor U12328 (N_12328,N_11916,N_11784);
nand U12329 (N_12329,N_11547,N_11686);
xor U12330 (N_12330,N_11999,N_11824);
or U12331 (N_12331,N_11637,N_11898);
xor U12332 (N_12332,N_11891,N_11875);
and U12333 (N_12333,N_11628,N_11680);
xor U12334 (N_12334,N_11910,N_11842);
xnor U12335 (N_12335,N_11942,N_11958);
nor U12336 (N_12336,N_11871,N_11986);
or U12337 (N_12337,N_11938,N_11642);
or U12338 (N_12338,N_11801,N_11963);
nor U12339 (N_12339,N_11727,N_11660);
and U12340 (N_12340,N_11795,N_11588);
or U12341 (N_12341,N_11545,N_11988);
or U12342 (N_12342,N_11712,N_11792);
xnor U12343 (N_12343,N_11802,N_11707);
xor U12344 (N_12344,N_11630,N_11883);
nand U12345 (N_12345,N_11660,N_11776);
nor U12346 (N_12346,N_11857,N_11587);
xnor U12347 (N_12347,N_11600,N_11870);
nor U12348 (N_12348,N_11570,N_11836);
and U12349 (N_12349,N_11778,N_11646);
or U12350 (N_12350,N_11955,N_11714);
xor U12351 (N_12351,N_11725,N_11749);
nor U12352 (N_12352,N_11853,N_11843);
or U12353 (N_12353,N_11907,N_11640);
or U12354 (N_12354,N_11563,N_11661);
or U12355 (N_12355,N_11858,N_11555);
nor U12356 (N_12356,N_11760,N_11560);
xnor U12357 (N_12357,N_11543,N_11936);
and U12358 (N_12358,N_11642,N_11652);
and U12359 (N_12359,N_11771,N_11890);
nand U12360 (N_12360,N_11909,N_11514);
or U12361 (N_12361,N_11608,N_11851);
nor U12362 (N_12362,N_11588,N_11949);
or U12363 (N_12363,N_11769,N_11885);
nor U12364 (N_12364,N_11621,N_11859);
nor U12365 (N_12365,N_11929,N_11766);
and U12366 (N_12366,N_11765,N_11763);
and U12367 (N_12367,N_11941,N_11966);
nor U12368 (N_12368,N_11814,N_11548);
nor U12369 (N_12369,N_11756,N_11593);
and U12370 (N_12370,N_11808,N_11556);
nand U12371 (N_12371,N_11599,N_11836);
xor U12372 (N_12372,N_11847,N_11787);
xnor U12373 (N_12373,N_11837,N_11626);
and U12374 (N_12374,N_11735,N_11564);
or U12375 (N_12375,N_11633,N_11584);
nor U12376 (N_12376,N_11822,N_11969);
or U12377 (N_12377,N_11955,N_11548);
and U12378 (N_12378,N_11744,N_11969);
nor U12379 (N_12379,N_11533,N_11973);
nand U12380 (N_12380,N_11621,N_11940);
and U12381 (N_12381,N_11771,N_11913);
and U12382 (N_12382,N_11655,N_11566);
xor U12383 (N_12383,N_11690,N_11683);
nor U12384 (N_12384,N_11726,N_11719);
or U12385 (N_12385,N_11892,N_11710);
nor U12386 (N_12386,N_11742,N_11796);
nand U12387 (N_12387,N_11804,N_11576);
or U12388 (N_12388,N_11849,N_11534);
nor U12389 (N_12389,N_11795,N_11893);
nand U12390 (N_12390,N_11972,N_11573);
nand U12391 (N_12391,N_11637,N_11604);
nand U12392 (N_12392,N_11977,N_11831);
nand U12393 (N_12393,N_11839,N_11507);
nor U12394 (N_12394,N_11875,N_11923);
xor U12395 (N_12395,N_11963,N_11572);
xor U12396 (N_12396,N_11953,N_11685);
and U12397 (N_12397,N_11733,N_11764);
nor U12398 (N_12398,N_11883,N_11507);
nor U12399 (N_12399,N_11569,N_11538);
and U12400 (N_12400,N_11662,N_11891);
or U12401 (N_12401,N_11646,N_11926);
and U12402 (N_12402,N_11618,N_11983);
or U12403 (N_12403,N_11982,N_11551);
or U12404 (N_12404,N_11981,N_11853);
nand U12405 (N_12405,N_11780,N_11830);
or U12406 (N_12406,N_11966,N_11893);
nand U12407 (N_12407,N_11914,N_11510);
nand U12408 (N_12408,N_11798,N_11522);
and U12409 (N_12409,N_11725,N_11744);
nor U12410 (N_12410,N_11955,N_11926);
nand U12411 (N_12411,N_11926,N_11977);
nand U12412 (N_12412,N_11522,N_11775);
or U12413 (N_12413,N_11511,N_11679);
and U12414 (N_12414,N_11652,N_11615);
and U12415 (N_12415,N_11803,N_11890);
and U12416 (N_12416,N_11924,N_11649);
and U12417 (N_12417,N_11883,N_11559);
and U12418 (N_12418,N_11923,N_11558);
nand U12419 (N_12419,N_11890,N_11783);
nor U12420 (N_12420,N_11566,N_11595);
or U12421 (N_12421,N_11948,N_11684);
and U12422 (N_12422,N_11518,N_11825);
and U12423 (N_12423,N_11811,N_11637);
nor U12424 (N_12424,N_11788,N_11829);
nand U12425 (N_12425,N_11971,N_11815);
nor U12426 (N_12426,N_11787,N_11639);
xor U12427 (N_12427,N_11685,N_11986);
nand U12428 (N_12428,N_11994,N_11893);
xor U12429 (N_12429,N_11785,N_11866);
nand U12430 (N_12430,N_11705,N_11936);
nand U12431 (N_12431,N_11746,N_11970);
nor U12432 (N_12432,N_11949,N_11945);
nand U12433 (N_12433,N_11855,N_11673);
nand U12434 (N_12434,N_11564,N_11955);
nor U12435 (N_12435,N_11783,N_11568);
xnor U12436 (N_12436,N_11978,N_11711);
xor U12437 (N_12437,N_11825,N_11923);
xnor U12438 (N_12438,N_11966,N_11880);
and U12439 (N_12439,N_11608,N_11656);
and U12440 (N_12440,N_11766,N_11667);
or U12441 (N_12441,N_11652,N_11937);
nand U12442 (N_12442,N_11565,N_11653);
nand U12443 (N_12443,N_11501,N_11784);
and U12444 (N_12444,N_11869,N_11668);
or U12445 (N_12445,N_11521,N_11576);
or U12446 (N_12446,N_11908,N_11935);
or U12447 (N_12447,N_11989,N_11658);
nor U12448 (N_12448,N_11891,N_11844);
nand U12449 (N_12449,N_11677,N_11623);
nand U12450 (N_12450,N_11638,N_11772);
or U12451 (N_12451,N_11681,N_11652);
and U12452 (N_12452,N_11929,N_11911);
nor U12453 (N_12453,N_11955,N_11678);
and U12454 (N_12454,N_11799,N_11825);
nor U12455 (N_12455,N_11938,N_11501);
nor U12456 (N_12456,N_11500,N_11544);
xor U12457 (N_12457,N_11997,N_11563);
xor U12458 (N_12458,N_11724,N_11937);
nand U12459 (N_12459,N_11951,N_11918);
nand U12460 (N_12460,N_11931,N_11716);
nor U12461 (N_12461,N_11780,N_11909);
nor U12462 (N_12462,N_11630,N_11904);
xnor U12463 (N_12463,N_11924,N_11588);
nand U12464 (N_12464,N_11563,N_11762);
nand U12465 (N_12465,N_11783,N_11728);
xor U12466 (N_12466,N_11748,N_11870);
xor U12467 (N_12467,N_11652,N_11968);
nand U12468 (N_12468,N_11588,N_11629);
and U12469 (N_12469,N_11850,N_11548);
nand U12470 (N_12470,N_11680,N_11581);
or U12471 (N_12471,N_11959,N_11779);
nor U12472 (N_12472,N_11958,N_11677);
nand U12473 (N_12473,N_11796,N_11902);
xnor U12474 (N_12474,N_11631,N_11821);
and U12475 (N_12475,N_11571,N_11881);
nand U12476 (N_12476,N_11796,N_11665);
nand U12477 (N_12477,N_11556,N_11626);
and U12478 (N_12478,N_11591,N_11636);
and U12479 (N_12479,N_11515,N_11892);
nor U12480 (N_12480,N_11809,N_11983);
and U12481 (N_12481,N_11859,N_11515);
nor U12482 (N_12482,N_11844,N_11553);
nor U12483 (N_12483,N_11601,N_11571);
and U12484 (N_12484,N_11612,N_11871);
or U12485 (N_12485,N_11986,N_11925);
or U12486 (N_12486,N_11721,N_11924);
nor U12487 (N_12487,N_11666,N_11765);
nor U12488 (N_12488,N_11693,N_11709);
nor U12489 (N_12489,N_11905,N_11977);
nand U12490 (N_12490,N_11615,N_11889);
nand U12491 (N_12491,N_11580,N_11836);
xnor U12492 (N_12492,N_11830,N_11886);
xnor U12493 (N_12493,N_11605,N_11833);
and U12494 (N_12494,N_11866,N_11573);
and U12495 (N_12495,N_11557,N_11778);
and U12496 (N_12496,N_11875,N_11863);
or U12497 (N_12497,N_11956,N_11813);
and U12498 (N_12498,N_11618,N_11979);
xor U12499 (N_12499,N_11943,N_11956);
and U12500 (N_12500,N_12037,N_12142);
xnor U12501 (N_12501,N_12379,N_12116);
nor U12502 (N_12502,N_12030,N_12102);
or U12503 (N_12503,N_12363,N_12454);
xnor U12504 (N_12504,N_12382,N_12295);
and U12505 (N_12505,N_12265,N_12251);
nor U12506 (N_12506,N_12232,N_12334);
xor U12507 (N_12507,N_12390,N_12151);
and U12508 (N_12508,N_12492,N_12278);
xor U12509 (N_12509,N_12496,N_12064);
nand U12510 (N_12510,N_12197,N_12369);
xnor U12511 (N_12511,N_12283,N_12261);
xnor U12512 (N_12512,N_12318,N_12017);
xor U12513 (N_12513,N_12333,N_12412);
or U12514 (N_12514,N_12019,N_12273);
or U12515 (N_12515,N_12188,N_12343);
and U12516 (N_12516,N_12158,N_12250);
or U12517 (N_12517,N_12422,N_12279);
nor U12518 (N_12518,N_12375,N_12244);
and U12519 (N_12519,N_12005,N_12353);
nor U12520 (N_12520,N_12374,N_12415);
nand U12521 (N_12521,N_12491,N_12267);
nand U12522 (N_12522,N_12264,N_12451);
or U12523 (N_12523,N_12266,N_12444);
nand U12524 (N_12524,N_12442,N_12337);
or U12525 (N_12525,N_12118,N_12323);
xnor U12526 (N_12526,N_12368,N_12354);
nand U12527 (N_12527,N_12080,N_12276);
and U12528 (N_12528,N_12238,N_12089);
or U12529 (N_12529,N_12067,N_12268);
and U12530 (N_12530,N_12270,N_12362);
xnor U12531 (N_12531,N_12289,N_12207);
xnor U12532 (N_12532,N_12129,N_12404);
or U12533 (N_12533,N_12445,N_12433);
or U12534 (N_12534,N_12311,N_12069);
nor U12535 (N_12535,N_12499,N_12438);
or U12536 (N_12536,N_12177,N_12044);
or U12537 (N_12537,N_12463,N_12312);
xor U12538 (N_12538,N_12141,N_12052);
and U12539 (N_12539,N_12274,N_12001);
or U12540 (N_12540,N_12408,N_12101);
nand U12541 (N_12541,N_12296,N_12436);
and U12542 (N_12542,N_12427,N_12477);
or U12543 (N_12543,N_12358,N_12332);
nand U12544 (N_12544,N_12034,N_12297);
and U12545 (N_12545,N_12465,N_12437);
nand U12546 (N_12546,N_12325,N_12128);
nor U12547 (N_12547,N_12046,N_12220);
xor U12548 (N_12548,N_12065,N_12347);
xnor U12549 (N_12549,N_12109,N_12075);
xnor U12550 (N_12550,N_12194,N_12204);
or U12551 (N_12551,N_12085,N_12348);
nand U12552 (N_12552,N_12399,N_12457);
nor U12553 (N_12553,N_12403,N_12309);
or U12554 (N_12554,N_12098,N_12303);
or U12555 (N_12555,N_12400,N_12271);
xor U12556 (N_12556,N_12466,N_12229);
nand U12557 (N_12557,N_12462,N_12235);
and U12558 (N_12558,N_12335,N_12164);
nor U12559 (N_12559,N_12062,N_12341);
and U12560 (N_12560,N_12282,N_12068);
nor U12561 (N_12561,N_12178,N_12394);
or U12562 (N_12562,N_12346,N_12191);
xor U12563 (N_12563,N_12166,N_12461);
nand U12564 (N_12564,N_12329,N_12099);
xnor U12565 (N_12565,N_12383,N_12114);
xor U12566 (N_12566,N_12136,N_12039);
or U12567 (N_12567,N_12317,N_12223);
and U12568 (N_12568,N_12228,N_12040);
xor U12569 (N_12569,N_12304,N_12010);
nor U12570 (N_12570,N_12074,N_12051);
nand U12571 (N_12571,N_12467,N_12377);
nand U12572 (N_12572,N_12108,N_12205);
xor U12573 (N_12573,N_12352,N_12149);
nor U12574 (N_12574,N_12262,N_12484);
nor U12575 (N_12575,N_12146,N_12410);
nand U12576 (N_12576,N_12219,N_12160);
and U12577 (N_12577,N_12119,N_12284);
xnor U12578 (N_12578,N_12066,N_12003);
or U12579 (N_12579,N_12198,N_12452);
or U12580 (N_12580,N_12315,N_12123);
nor U12581 (N_12581,N_12246,N_12389);
nor U12582 (N_12582,N_12104,N_12431);
and U12583 (N_12583,N_12218,N_12277);
xnor U12584 (N_12584,N_12256,N_12053);
xnor U12585 (N_12585,N_12336,N_12168);
and U12586 (N_12586,N_12161,N_12418);
and U12587 (N_12587,N_12455,N_12169);
nor U12588 (N_12588,N_12327,N_12092);
or U12589 (N_12589,N_12137,N_12090);
xnor U12590 (N_12590,N_12206,N_12260);
nand U12591 (N_12591,N_12392,N_12018);
and U12592 (N_12592,N_12026,N_12187);
nor U12593 (N_12593,N_12148,N_12294);
or U12594 (N_12594,N_12185,N_12319);
nor U12595 (N_12595,N_12331,N_12322);
nand U12596 (N_12596,N_12082,N_12456);
nor U12597 (N_12597,N_12468,N_12378);
nor U12598 (N_12598,N_12339,N_12350);
nand U12599 (N_12599,N_12401,N_12120);
nor U12600 (N_12600,N_12047,N_12371);
xnor U12601 (N_12601,N_12201,N_12012);
nor U12602 (N_12602,N_12131,N_12022);
nand U12603 (N_12603,N_12248,N_12421);
or U12604 (N_12604,N_12285,N_12395);
and U12605 (N_12605,N_12231,N_12426);
nand U12606 (N_12606,N_12416,N_12310);
nand U12607 (N_12607,N_12088,N_12439);
or U12608 (N_12608,N_12269,N_12298);
nand U12609 (N_12609,N_12073,N_12417);
xnor U12610 (N_12610,N_12247,N_12060);
nor U12611 (N_12611,N_12076,N_12095);
xnor U12612 (N_12612,N_12174,N_12487);
nand U12613 (N_12613,N_12464,N_12111);
or U12614 (N_12614,N_12171,N_12008);
xor U12615 (N_12615,N_12405,N_12113);
nor U12616 (N_12616,N_12221,N_12316);
nor U12617 (N_12617,N_12117,N_12447);
or U12618 (N_12618,N_12242,N_12470);
or U12619 (N_12619,N_12059,N_12132);
or U12620 (N_12620,N_12411,N_12497);
xnor U12621 (N_12621,N_12083,N_12225);
nand U12622 (N_12622,N_12255,N_12483);
xnor U12623 (N_12623,N_12291,N_12459);
and U12624 (N_12624,N_12173,N_12002);
and U12625 (N_12625,N_12321,N_12328);
and U12626 (N_12626,N_12428,N_12391);
nor U12627 (N_12627,N_12097,N_12349);
or U12628 (N_12628,N_12366,N_12139);
nor U12629 (N_12629,N_12100,N_12406);
nor U12630 (N_12630,N_12373,N_12007);
nand U12631 (N_12631,N_12424,N_12004);
or U12632 (N_12632,N_12121,N_12308);
xor U12633 (N_12633,N_12193,N_12125);
xor U12634 (N_12634,N_12430,N_12230);
or U12635 (N_12635,N_12480,N_12380);
xnor U12636 (N_12636,N_12450,N_12181);
and U12637 (N_12637,N_12079,N_12393);
nor U12638 (N_12638,N_12443,N_12199);
xnor U12639 (N_12639,N_12478,N_12023);
and U12640 (N_12640,N_12063,N_12184);
xnor U12641 (N_12641,N_12413,N_12195);
or U12642 (N_12642,N_12376,N_12448);
and U12643 (N_12643,N_12388,N_12330);
nor U12644 (N_12644,N_12453,N_12227);
xor U12645 (N_12645,N_12179,N_12152);
xor U12646 (N_12646,N_12140,N_12435);
xnor U12647 (N_12647,N_12275,N_12127);
and U12648 (N_12648,N_12154,N_12021);
or U12649 (N_12649,N_12014,N_12359);
nand U12650 (N_12650,N_12106,N_12407);
nand U12651 (N_12651,N_12498,N_12287);
nor U12652 (N_12652,N_12049,N_12036);
xnor U12653 (N_12653,N_12344,N_12084);
nand U12654 (N_12654,N_12471,N_12292);
nor U12655 (N_12655,N_12057,N_12087);
nor U12656 (N_12656,N_12200,N_12299);
nand U12657 (N_12657,N_12240,N_12054);
or U12658 (N_12658,N_12211,N_12110);
nor U12659 (N_12659,N_12093,N_12288);
nand U12660 (N_12660,N_12351,N_12257);
nand U12661 (N_12661,N_12214,N_12203);
and U12662 (N_12662,N_12409,N_12081);
xor U12663 (N_12663,N_12425,N_12009);
xnor U12664 (N_12664,N_12420,N_12028);
or U12665 (N_12665,N_12441,N_12027);
and U12666 (N_12666,N_12155,N_12326);
xor U12667 (N_12667,N_12045,N_12361);
or U12668 (N_12668,N_12280,N_12086);
and U12669 (N_12669,N_12189,N_12212);
and U12670 (N_12670,N_12272,N_12217);
nor U12671 (N_12671,N_12342,N_12167);
nor U12672 (N_12672,N_12135,N_12112);
nand U12673 (N_12673,N_12449,N_12460);
or U12674 (N_12674,N_12387,N_12091);
or U12675 (N_12675,N_12486,N_12286);
xnor U12676 (N_12676,N_12365,N_12489);
or U12677 (N_12677,N_12186,N_12226);
nand U12678 (N_12678,N_12048,N_12340);
or U12679 (N_12679,N_12143,N_12432);
xor U12680 (N_12680,N_12245,N_12025);
nand U12681 (N_12681,N_12234,N_12077);
nor U12682 (N_12682,N_12338,N_12306);
xor U12683 (N_12683,N_12243,N_12041);
nor U12684 (N_12684,N_12124,N_12153);
nor U12685 (N_12685,N_12020,N_12429);
xor U12686 (N_12686,N_12305,N_12133);
nor U12687 (N_12687,N_12482,N_12222);
nand U12688 (N_12688,N_12182,N_12290);
xnor U12689 (N_12689,N_12042,N_12031);
and U12690 (N_12690,N_12458,N_12381);
nand U12691 (N_12691,N_12355,N_12367);
or U12692 (N_12692,N_12253,N_12038);
nor U12693 (N_12693,N_12215,N_12006);
xor U12694 (N_12694,N_12474,N_12015);
or U12695 (N_12695,N_12050,N_12029);
and U12696 (N_12696,N_12372,N_12162);
and U12697 (N_12697,N_12150,N_12414);
nor U12698 (N_12698,N_12175,N_12024);
nor U12699 (N_12699,N_12176,N_12071);
and U12700 (N_12700,N_12145,N_12300);
nor U12701 (N_12701,N_12370,N_12016);
or U12702 (N_12702,N_12386,N_12473);
or U12703 (N_12703,N_12055,N_12281);
xor U12704 (N_12704,N_12130,N_12170);
xnor U12705 (N_12705,N_12043,N_12384);
or U12706 (N_12706,N_12239,N_12397);
xor U12707 (N_12707,N_12313,N_12192);
or U12708 (N_12708,N_12385,N_12423);
nand U12709 (N_12709,N_12476,N_12263);
nor U12710 (N_12710,N_12490,N_12398);
nor U12711 (N_12711,N_12237,N_12208);
xor U12712 (N_12712,N_12180,N_12147);
and U12713 (N_12713,N_12360,N_12494);
nand U12714 (N_12714,N_12183,N_12241);
and U12715 (N_12715,N_12488,N_12402);
and U12716 (N_12716,N_12446,N_12224);
xnor U12717 (N_12717,N_12485,N_12061);
nor U12718 (N_12718,N_12011,N_12165);
nor U12719 (N_12719,N_12254,N_12302);
or U12720 (N_12720,N_12163,N_12493);
nor U12721 (N_12721,N_12013,N_12210);
and U12722 (N_12722,N_12202,N_12236);
nand U12723 (N_12723,N_12115,N_12213);
xor U12724 (N_12724,N_12320,N_12307);
nand U12725 (N_12725,N_12209,N_12035);
or U12726 (N_12726,N_12356,N_12032);
xor U12727 (N_12727,N_12078,N_12159);
nand U12728 (N_12728,N_12472,N_12107);
and U12729 (N_12729,N_12434,N_12126);
nor U12730 (N_12730,N_12233,N_12440);
nand U12731 (N_12731,N_12479,N_12190);
xor U12732 (N_12732,N_12301,N_12475);
xnor U12733 (N_12733,N_12156,N_12396);
nor U12734 (N_12734,N_12495,N_12216);
xor U12735 (N_12735,N_12324,N_12258);
and U12736 (N_12736,N_12105,N_12293);
xnor U12737 (N_12737,N_12094,N_12252);
or U12738 (N_12738,N_12419,N_12157);
xnor U12739 (N_12739,N_12357,N_12314);
nor U12740 (N_12740,N_12103,N_12345);
or U12741 (N_12741,N_12196,N_12469);
or U12742 (N_12742,N_12138,N_12364);
nand U12743 (N_12743,N_12134,N_12070);
and U12744 (N_12744,N_12249,N_12058);
and U12745 (N_12745,N_12481,N_12144);
and U12746 (N_12746,N_12096,N_12072);
and U12747 (N_12747,N_12172,N_12056);
or U12748 (N_12748,N_12000,N_12122);
nor U12749 (N_12749,N_12259,N_12033);
or U12750 (N_12750,N_12294,N_12250);
nand U12751 (N_12751,N_12171,N_12121);
nand U12752 (N_12752,N_12009,N_12045);
xor U12753 (N_12753,N_12190,N_12404);
and U12754 (N_12754,N_12292,N_12108);
or U12755 (N_12755,N_12148,N_12153);
and U12756 (N_12756,N_12093,N_12325);
xor U12757 (N_12757,N_12336,N_12329);
xnor U12758 (N_12758,N_12128,N_12288);
xnor U12759 (N_12759,N_12346,N_12172);
or U12760 (N_12760,N_12197,N_12145);
nand U12761 (N_12761,N_12005,N_12322);
xor U12762 (N_12762,N_12102,N_12247);
nand U12763 (N_12763,N_12139,N_12447);
nand U12764 (N_12764,N_12438,N_12471);
nand U12765 (N_12765,N_12269,N_12490);
nand U12766 (N_12766,N_12184,N_12302);
or U12767 (N_12767,N_12409,N_12235);
nor U12768 (N_12768,N_12112,N_12306);
nand U12769 (N_12769,N_12128,N_12048);
nand U12770 (N_12770,N_12370,N_12090);
or U12771 (N_12771,N_12352,N_12293);
and U12772 (N_12772,N_12209,N_12181);
and U12773 (N_12773,N_12070,N_12131);
xor U12774 (N_12774,N_12367,N_12321);
or U12775 (N_12775,N_12388,N_12380);
nand U12776 (N_12776,N_12007,N_12148);
or U12777 (N_12777,N_12192,N_12195);
or U12778 (N_12778,N_12484,N_12152);
xnor U12779 (N_12779,N_12165,N_12047);
or U12780 (N_12780,N_12061,N_12258);
xor U12781 (N_12781,N_12325,N_12480);
nand U12782 (N_12782,N_12063,N_12315);
xor U12783 (N_12783,N_12446,N_12355);
and U12784 (N_12784,N_12231,N_12168);
nand U12785 (N_12785,N_12474,N_12260);
and U12786 (N_12786,N_12138,N_12304);
and U12787 (N_12787,N_12052,N_12437);
xor U12788 (N_12788,N_12015,N_12346);
xor U12789 (N_12789,N_12187,N_12483);
and U12790 (N_12790,N_12115,N_12461);
and U12791 (N_12791,N_12466,N_12100);
nor U12792 (N_12792,N_12471,N_12418);
nor U12793 (N_12793,N_12336,N_12186);
or U12794 (N_12794,N_12100,N_12474);
nor U12795 (N_12795,N_12275,N_12082);
xor U12796 (N_12796,N_12336,N_12420);
and U12797 (N_12797,N_12435,N_12014);
and U12798 (N_12798,N_12215,N_12212);
nand U12799 (N_12799,N_12139,N_12397);
xnor U12800 (N_12800,N_12470,N_12268);
xor U12801 (N_12801,N_12136,N_12235);
or U12802 (N_12802,N_12409,N_12256);
xnor U12803 (N_12803,N_12357,N_12412);
nand U12804 (N_12804,N_12077,N_12311);
xnor U12805 (N_12805,N_12490,N_12458);
or U12806 (N_12806,N_12245,N_12202);
xnor U12807 (N_12807,N_12037,N_12065);
or U12808 (N_12808,N_12163,N_12167);
xor U12809 (N_12809,N_12067,N_12290);
nand U12810 (N_12810,N_12165,N_12180);
and U12811 (N_12811,N_12004,N_12431);
xnor U12812 (N_12812,N_12082,N_12048);
or U12813 (N_12813,N_12271,N_12414);
nor U12814 (N_12814,N_12335,N_12142);
or U12815 (N_12815,N_12112,N_12397);
nor U12816 (N_12816,N_12260,N_12165);
nand U12817 (N_12817,N_12220,N_12318);
nor U12818 (N_12818,N_12263,N_12288);
or U12819 (N_12819,N_12144,N_12300);
nand U12820 (N_12820,N_12151,N_12251);
nor U12821 (N_12821,N_12358,N_12324);
and U12822 (N_12822,N_12083,N_12169);
nor U12823 (N_12823,N_12364,N_12187);
or U12824 (N_12824,N_12476,N_12353);
nor U12825 (N_12825,N_12017,N_12069);
or U12826 (N_12826,N_12042,N_12140);
xnor U12827 (N_12827,N_12348,N_12079);
xnor U12828 (N_12828,N_12110,N_12155);
nor U12829 (N_12829,N_12266,N_12142);
nor U12830 (N_12830,N_12246,N_12298);
xnor U12831 (N_12831,N_12274,N_12430);
or U12832 (N_12832,N_12351,N_12355);
or U12833 (N_12833,N_12498,N_12111);
nor U12834 (N_12834,N_12355,N_12448);
nor U12835 (N_12835,N_12137,N_12070);
nand U12836 (N_12836,N_12243,N_12258);
or U12837 (N_12837,N_12039,N_12295);
or U12838 (N_12838,N_12320,N_12129);
and U12839 (N_12839,N_12483,N_12336);
nor U12840 (N_12840,N_12356,N_12056);
nor U12841 (N_12841,N_12285,N_12070);
xor U12842 (N_12842,N_12434,N_12029);
nor U12843 (N_12843,N_12395,N_12275);
nor U12844 (N_12844,N_12066,N_12290);
nor U12845 (N_12845,N_12363,N_12420);
or U12846 (N_12846,N_12416,N_12075);
or U12847 (N_12847,N_12004,N_12259);
or U12848 (N_12848,N_12328,N_12198);
nor U12849 (N_12849,N_12113,N_12345);
or U12850 (N_12850,N_12228,N_12086);
nor U12851 (N_12851,N_12278,N_12364);
or U12852 (N_12852,N_12142,N_12263);
nor U12853 (N_12853,N_12449,N_12100);
nor U12854 (N_12854,N_12135,N_12159);
nor U12855 (N_12855,N_12269,N_12085);
or U12856 (N_12856,N_12282,N_12260);
or U12857 (N_12857,N_12358,N_12048);
or U12858 (N_12858,N_12257,N_12371);
nand U12859 (N_12859,N_12095,N_12206);
nand U12860 (N_12860,N_12466,N_12426);
nor U12861 (N_12861,N_12150,N_12145);
xnor U12862 (N_12862,N_12141,N_12110);
and U12863 (N_12863,N_12234,N_12423);
nor U12864 (N_12864,N_12099,N_12105);
nand U12865 (N_12865,N_12011,N_12473);
and U12866 (N_12866,N_12001,N_12426);
and U12867 (N_12867,N_12412,N_12163);
and U12868 (N_12868,N_12196,N_12142);
xnor U12869 (N_12869,N_12473,N_12289);
nor U12870 (N_12870,N_12458,N_12234);
and U12871 (N_12871,N_12149,N_12232);
or U12872 (N_12872,N_12078,N_12281);
nor U12873 (N_12873,N_12417,N_12355);
xor U12874 (N_12874,N_12039,N_12140);
and U12875 (N_12875,N_12250,N_12395);
nor U12876 (N_12876,N_12239,N_12450);
xor U12877 (N_12877,N_12418,N_12154);
nor U12878 (N_12878,N_12033,N_12456);
and U12879 (N_12879,N_12435,N_12459);
and U12880 (N_12880,N_12353,N_12151);
and U12881 (N_12881,N_12060,N_12166);
nor U12882 (N_12882,N_12392,N_12452);
nand U12883 (N_12883,N_12490,N_12483);
nand U12884 (N_12884,N_12003,N_12191);
and U12885 (N_12885,N_12039,N_12387);
and U12886 (N_12886,N_12202,N_12392);
and U12887 (N_12887,N_12409,N_12326);
nor U12888 (N_12888,N_12359,N_12032);
xnor U12889 (N_12889,N_12227,N_12326);
nor U12890 (N_12890,N_12039,N_12415);
xnor U12891 (N_12891,N_12493,N_12378);
or U12892 (N_12892,N_12399,N_12177);
nand U12893 (N_12893,N_12169,N_12432);
xor U12894 (N_12894,N_12129,N_12312);
xnor U12895 (N_12895,N_12048,N_12267);
nor U12896 (N_12896,N_12004,N_12142);
nor U12897 (N_12897,N_12336,N_12367);
nand U12898 (N_12898,N_12345,N_12210);
or U12899 (N_12899,N_12019,N_12101);
or U12900 (N_12900,N_12082,N_12398);
xnor U12901 (N_12901,N_12341,N_12494);
xnor U12902 (N_12902,N_12090,N_12154);
nand U12903 (N_12903,N_12200,N_12232);
nand U12904 (N_12904,N_12248,N_12120);
nand U12905 (N_12905,N_12232,N_12341);
nand U12906 (N_12906,N_12486,N_12147);
xor U12907 (N_12907,N_12292,N_12269);
or U12908 (N_12908,N_12395,N_12184);
and U12909 (N_12909,N_12289,N_12019);
nand U12910 (N_12910,N_12474,N_12087);
xnor U12911 (N_12911,N_12471,N_12218);
nand U12912 (N_12912,N_12422,N_12105);
or U12913 (N_12913,N_12211,N_12098);
and U12914 (N_12914,N_12241,N_12132);
nor U12915 (N_12915,N_12208,N_12210);
nor U12916 (N_12916,N_12383,N_12199);
nand U12917 (N_12917,N_12468,N_12379);
and U12918 (N_12918,N_12391,N_12150);
nand U12919 (N_12919,N_12115,N_12172);
nor U12920 (N_12920,N_12229,N_12448);
xor U12921 (N_12921,N_12287,N_12250);
or U12922 (N_12922,N_12016,N_12046);
and U12923 (N_12923,N_12258,N_12361);
nand U12924 (N_12924,N_12433,N_12203);
and U12925 (N_12925,N_12438,N_12114);
nor U12926 (N_12926,N_12361,N_12091);
and U12927 (N_12927,N_12253,N_12202);
nand U12928 (N_12928,N_12156,N_12340);
or U12929 (N_12929,N_12342,N_12104);
nor U12930 (N_12930,N_12460,N_12140);
nor U12931 (N_12931,N_12164,N_12046);
nor U12932 (N_12932,N_12092,N_12086);
xnor U12933 (N_12933,N_12155,N_12303);
nor U12934 (N_12934,N_12129,N_12126);
or U12935 (N_12935,N_12154,N_12263);
nor U12936 (N_12936,N_12151,N_12147);
and U12937 (N_12937,N_12191,N_12337);
nor U12938 (N_12938,N_12139,N_12145);
or U12939 (N_12939,N_12261,N_12034);
and U12940 (N_12940,N_12342,N_12263);
nand U12941 (N_12941,N_12179,N_12083);
or U12942 (N_12942,N_12370,N_12468);
xor U12943 (N_12943,N_12423,N_12468);
nor U12944 (N_12944,N_12277,N_12388);
nand U12945 (N_12945,N_12308,N_12237);
xnor U12946 (N_12946,N_12050,N_12300);
and U12947 (N_12947,N_12060,N_12093);
and U12948 (N_12948,N_12034,N_12492);
or U12949 (N_12949,N_12157,N_12063);
xnor U12950 (N_12950,N_12033,N_12349);
or U12951 (N_12951,N_12317,N_12481);
nor U12952 (N_12952,N_12447,N_12253);
nor U12953 (N_12953,N_12105,N_12490);
and U12954 (N_12954,N_12118,N_12408);
and U12955 (N_12955,N_12083,N_12170);
nand U12956 (N_12956,N_12080,N_12176);
xnor U12957 (N_12957,N_12443,N_12075);
and U12958 (N_12958,N_12205,N_12137);
xor U12959 (N_12959,N_12454,N_12484);
nand U12960 (N_12960,N_12238,N_12447);
nand U12961 (N_12961,N_12130,N_12460);
and U12962 (N_12962,N_12293,N_12469);
or U12963 (N_12963,N_12236,N_12114);
nand U12964 (N_12964,N_12082,N_12238);
and U12965 (N_12965,N_12156,N_12157);
and U12966 (N_12966,N_12202,N_12386);
and U12967 (N_12967,N_12058,N_12454);
nand U12968 (N_12968,N_12071,N_12150);
nor U12969 (N_12969,N_12040,N_12398);
nand U12970 (N_12970,N_12334,N_12063);
and U12971 (N_12971,N_12161,N_12060);
and U12972 (N_12972,N_12131,N_12163);
nand U12973 (N_12973,N_12025,N_12356);
xor U12974 (N_12974,N_12320,N_12225);
nand U12975 (N_12975,N_12295,N_12261);
or U12976 (N_12976,N_12371,N_12076);
nor U12977 (N_12977,N_12281,N_12107);
or U12978 (N_12978,N_12069,N_12338);
nor U12979 (N_12979,N_12107,N_12263);
and U12980 (N_12980,N_12067,N_12051);
or U12981 (N_12981,N_12111,N_12060);
or U12982 (N_12982,N_12253,N_12052);
nand U12983 (N_12983,N_12003,N_12069);
xor U12984 (N_12984,N_12033,N_12139);
and U12985 (N_12985,N_12104,N_12450);
nor U12986 (N_12986,N_12377,N_12341);
nor U12987 (N_12987,N_12143,N_12021);
xnor U12988 (N_12988,N_12405,N_12153);
and U12989 (N_12989,N_12102,N_12052);
xor U12990 (N_12990,N_12065,N_12094);
xnor U12991 (N_12991,N_12047,N_12309);
xnor U12992 (N_12992,N_12196,N_12149);
or U12993 (N_12993,N_12185,N_12115);
and U12994 (N_12994,N_12172,N_12069);
xnor U12995 (N_12995,N_12065,N_12286);
nand U12996 (N_12996,N_12205,N_12434);
nor U12997 (N_12997,N_12287,N_12006);
or U12998 (N_12998,N_12381,N_12315);
or U12999 (N_12999,N_12003,N_12082);
xor U13000 (N_13000,N_12910,N_12601);
nand U13001 (N_13001,N_12623,N_12664);
xor U13002 (N_13002,N_12905,N_12709);
nand U13003 (N_13003,N_12551,N_12695);
and U13004 (N_13004,N_12805,N_12611);
and U13005 (N_13005,N_12827,N_12503);
or U13006 (N_13006,N_12795,N_12908);
and U13007 (N_13007,N_12912,N_12570);
xor U13008 (N_13008,N_12927,N_12763);
or U13009 (N_13009,N_12775,N_12850);
nand U13010 (N_13010,N_12972,N_12918);
and U13011 (N_13011,N_12757,N_12577);
xor U13012 (N_13012,N_12802,N_12739);
or U13013 (N_13013,N_12837,N_12629);
nand U13014 (N_13014,N_12564,N_12703);
nand U13015 (N_13015,N_12816,N_12792);
nor U13016 (N_13016,N_12771,N_12834);
nand U13017 (N_13017,N_12929,N_12530);
or U13018 (N_13018,N_12576,N_12890);
xnor U13019 (N_13019,N_12839,N_12637);
xnor U13020 (N_13020,N_12549,N_12661);
nor U13021 (N_13021,N_12624,N_12870);
and U13022 (N_13022,N_12589,N_12559);
nor U13023 (N_13023,N_12980,N_12963);
or U13024 (N_13024,N_12959,N_12788);
xor U13025 (N_13025,N_12883,N_12854);
and U13026 (N_13026,N_12884,N_12732);
nor U13027 (N_13027,N_12777,N_12666);
xor U13028 (N_13028,N_12600,N_12644);
and U13029 (N_13029,N_12701,N_12774);
nand U13030 (N_13030,N_12627,N_12713);
nor U13031 (N_13031,N_12736,N_12741);
nor U13032 (N_13032,N_12799,N_12652);
or U13033 (N_13033,N_12533,N_12902);
nor U13034 (N_13034,N_12532,N_12989);
nand U13035 (N_13035,N_12800,N_12588);
and U13036 (N_13036,N_12614,N_12747);
and U13037 (N_13037,N_12853,N_12649);
xor U13038 (N_13038,N_12783,N_12668);
and U13039 (N_13039,N_12937,N_12803);
xnor U13040 (N_13040,N_12517,N_12746);
xor U13041 (N_13041,N_12761,N_12721);
nor U13042 (N_13042,N_12596,N_12597);
and U13043 (N_13043,N_12509,N_12572);
nor U13044 (N_13044,N_12913,N_12969);
nor U13045 (N_13045,N_12770,N_12983);
nor U13046 (N_13046,N_12906,N_12907);
nand U13047 (N_13047,N_12851,N_12791);
or U13048 (N_13048,N_12798,N_12866);
nand U13049 (N_13049,N_12840,N_12698);
and U13050 (N_13050,N_12557,N_12892);
and U13051 (N_13051,N_12943,N_12808);
nand U13052 (N_13052,N_12678,N_12960);
and U13053 (N_13053,N_12690,N_12848);
and U13054 (N_13054,N_12651,N_12582);
and U13055 (N_13055,N_12782,N_12897);
or U13056 (N_13056,N_12751,N_12683);
nand U13057 (N_13057,N_12821,N_12830);
nand U13058 (N_13058,N_12780,N_12928);
or U13059 (N_13059,N_12618,N_12710);
or U13060 (N_13060,N_12944,N_12714);
nand U13061 (N_13061,N_12767,N_12794);
nand U13062 (N_13062,N_12919,N_12645);
and U13063 (N_13063,N_12749,N_12764);
nor U13064 (N_13064,N_12641,N_12738);
nand U13065 (N_13065,N_12935,N_12612);
xor U13066 (N_13066,N_12542,N_12901);
nor U13067 (N_13067,N_12529,N_12545);
nor U13068 (N_13068,N_12541,N_12986);
or U13069 (N_13069,N_12752,N_12676);
nor U13070 (N_13070,N_12544,N_12687);
xnor U13071 (N_13071,N_12514,N_12697);
and U13072 (N_13072,N_12864,N_12616);
xnor U13073 (N_13073,N_12587,N_12941);
and U13074 (N_13074,N_12519,N_12583);
and U13075 (N_13075,N_12524,N_12622);
nor U13076 (N_13076,N_12942,N_12691);
xnor U13077 (N_13077,N_12828,N_12825);
and U13078 (N_13078,N_12797,N_12726);
or U13079 (N_13079,N_12914,N_12855);
or U13080 (N_13080,N_12565,N_12586);
nand U13081 (N_13081,N_12847,N_12879);
nor U13082 (N_13082,N_12987,N_12953);
nor U13083 (N_13083,N_12688,N_12553);
xor U13084 (N_13084,N_12638,N_12733);
or U13085 (N_13085,N_12886,N_12501);
nand U13086 (N_13086,N_12956,N_12599);
nor U13087 (N_13087,N_12820,N_12663);
nand U13088 (N_13088,N_12702,N_12671);
and U13089 (N_13089,N_12885,N_12590);
nand U13090 (N_13090,N_12762,N_12955);
or U13091 (N_13091,N_12547,N_12674);
nor U13092 (N_13092,N_12540,N_12608);
and U13093 (N_13093,N_12526,N_12900);
nor U13094 (N_13094,N_12613,N_12998);
xnor U13095 (N_13095,N_12766,N_12558);
or U13096 (N_13096,N_12996,N_12872);
nor U13097 (N_13097,N_12521,N_12745);
and U13098 (N_13098,N_12887,N_12716);
nand U13099 (N_13099,N_12968,N_12835);
nand U13100 (N_13100,N_12786,N_12575);
and U13101 (N_13101,N_12659,N_12724);
and U13102 (N_13102,N_12658,N_12573);
and U13103 (N_13103,N_12880,N_12593);
nand U13104 (N_13104,N_12778,N_12723);
or U13105 (N_13105,N_12842,N_12977);
nor U13106 (N_13106,N_12743,N_12539);
nand U13107 (N_13107,N_12954,N_12528);
or U13108 (N_13108,N_12603,N_12858);
nor U13109 (N_13109,N_12952,N_12862);
or U13110 (N_13110,N_12995,N_12833);
or U13111 (N_13111,N_12997,N_12932);
nand U13112 (N_13112,N_12926,N_12888);
and U13113 (N_13113,N_12689,N_12568);
nand U13114 (N_13114,N_12563,N_12680);
nor U13115 (N_13115,N_12648,N_12605);
and U13116 (N_13116,N_12964,N_12643);
nand U13117 (N_13117,N_12988,N_12505);
nor U13118 (N_13118,N_12734,N_12807);
or U13119 (N_13119,N_12957,N_12554);
nand U13120 (N_13120,N_12704,N_12898);
and U13121 (N_13121,N_12515,N_12699);
nor U13122 (N_13122,N_12522,N_12773);
nor U13123 (N_13123,N_12894,N_12657);
nand U13124 (N_13124,N_12779,N_12809);
nor U13125 (N_13125,N_12585,N_12580);
nor U13126 (N_13126,N_12920,N_12958);
and U13127 (N_13127,N_12868,N_12844);
nand U13128 (N_13128,N_12976,N_12843);
nand U13129 (N_13129,N_12740,N_12817);
and U13130 (N_13130,N_12630,N_12717);
nand U13131 (N_13131,N_12925,N_12889);
nand U13132 (N_13132,N_12841,N_12708);
nand U13133 (N_13133,N_12631,N_12822);
or U13134 (N_13134,N_12684,N_12707);
or U13135 (N_13135,N_12975,N_12633);
nand U13136 (N_13136,N_12653,N_12634);
or U13137 (N_13137,N_12720,N_12978);
or U13138 (N_13138,N_12829,N_12518);
nor U13139 (N_13139,N_12815,N_12536);
nand U13140 (N_13140,N_12974,N_12917);
and U13141 (N_13141,N_12660,N_12617);
xor U13142 (N_13142,N_12538,N_12874);
nand U13143 (N_13143,N_12502,N_12811);
nor U13144 (N_13144,N_12903,N_12607);
xnor U13145 (N_13145,N_12730,N_12647);
or U13146 (N_13146,N_12620,N_12504);
nand U13147 (N_13147,N_12625,N_12606);
xor U13148 (N_13148,N_12863,N_12748);
nor U13149 (N_13149,N_12686,N_12804);
nand U13150 (N_13150,N_12857,N_12673);
nand U13151 (N_13151,N_12574,N_12985);
xor U13152 (N_13152,N_12961,N_12856);
and U13153 (N_13153,N_12527,N_12970);
or U13154 (N_13154,N_12507,N_12896);
nand U13155 (N_13155,N_12694,N_12569);
nor U13156 (N_13156,N_12556,N_12621);
or U13157 (N_13157,N_12911,N_12523);
nor U13158 (N_13158,N_12966,N_12685);
and U13159 (N_13159,N_12768,N_12632);
nand U13160 (N_13160,N_12669,N_12508);
nand U13161 (N_13161,N_12846,N_12849);
nand U13162 (N_13162,N_12591,N_12873);
nand U13163 (N_13163,N_12722,N_12810);
nand U13164 (N_13164,N_12836,N_12965);
xnor U13165 (N_13165,N_12604,N_12594);
nor U13166 (N_13166,N_12772,N_12930);
and U13167 (N_13167,N_12578,N_12973);
nand U13168 (N_13168,N_12650,N_12759);
xnor U13169 (N_13169,N_12619,N_12693);
xor U13170 (N_13170,N_12560,N_12531);
or U13171 (N_13171,N_12784,N_12548);
and U13172 (N_13172,N_12512,N_12656);
xor U13173 (N_13173,N_12546,N_12991);
nor U13174 (N_13174,N_12994,N_12670);
nor U13175 (N_13175,N_12729,N_12584);
xor U13176 (N_13176,N_12737,N_12785);
nor U13177 (N_13177,N_12769,N_12877);
xor U13178 (N_13178,N_12881,N_12818);
xnor U13179 (N_13179,N_12566,N_12758);
xor U13180 (N_13180,N_12790,N_12706);
nor U13181 (N_13181,N_12990,N_12639);
xnor U13182 (N_13182,N_12999,N_12513);
nand U13183 (N_13183,N_12951,N_12940);
nand U13184 (N_13184,N_12552,N_12719);
and U13185 (N_13185,N_12787,N_12789);
and U13186 (N_13186,N_12859,N_12636);
nor U13187 (N_13187,N_12826,N_12993);
xnor U13188 (N_13188,N_12646,N_12579);
or U13189 (N_13189,N_12592,N_12510);
nand U13190 (N_13190,N_12750,N_12878);
or U13191 (N_13191,N_12852,N_12700);
nor U13192 (N_13192,N_12967,N_12675);
xor U13193 (N_13193,N_12626,N_12814);
or U13194 (N_13194,N_12715,N_12893);
nor U13195 (N_13195,N_12712,N_12662);
or U13196 (N_13196,N_12711,N_12555);
nand U13197 (N_13197,N_12754,N_12760);
and U13198 (N_13198,N_12550,N_12665);
xnor U13199 (N_13199,N_12735,N_12642);
nor U13200 (N_13200,N_12945,N_12946);
and U13201 (N_13201,N_12742,N_12876);
or U13202 (N_13202,N_12933,N_12981);
and U13203 (N_13203,N_12875,N_12755);
or U13204 (N_13204,N_12796,N_12895);
xor U13205 (N_13205,N_12654,N_12667);
and U13206 (N_13206,N_12947,N_12819);
nand U13207 (N_13207,N_12831,N_12979);
or U13208 (N_13208,N_12534,N_12725);
nand U13209 (N_13209,N_12506,N_12682);
xnor U13210 (N_13210,N_12971,N_12609);
nor U13211 (N_13211,N_12571,N_12562);
or U13212 (N_13212,N_12860,N_12635);
nand U13213 (N_13213,N_12869,N_12537);
or U13214 (N_13214,N_12561,N_12921);
nand U13215 (N_13215,N_12832,N_12744);
or U13216 (N_13216,N_12882,N_12992);
nor U13217 (N_13217,N_12610,N_12909);
or U13218 (N_13218,N_12598,N_12679);
or U13219 (N_13219,N_12602,N_12812);
or U13220 (N_13220,N_12867,N_12904);
or U13221 (N_13221,N_12776,N_12628);
nand U13222 (N_13222,N_12891,N_12899);
and U13223 (N_13223,N_12934,N_12535);
xor U13224 (N_13224,N_12681,N_12806);
xor U13225 (N_13225,N_12781,N_12939);
nand U13226 (N_13226,N_12718,N_12728);
nand U13227 (N_13227,N_12924,N_12984);
xnor U13228 (N_13228,N_12793,N_12543);
or U13229 (N_13229,N_12865,N_12936);
nand U13230 (N_13230,N_12823,N_12916);
nand U13231 (N_13231,N_12962,N_12861);
xnor U13232 (N_13232,N_12567,N_12692);
xor U13233 (N_13233,N_12677,N_12949);
nor U13234 (N_13234,N_12922,N_12520);
and U13235 (N_13235,N_12696,N_12931);
nor U13236 (N_13236,N_12871,N_12615);
or U13237 (N_13237,N_12948,N_12655);
and U13238 (N_13238,N_12672,N_12511);
nand U13239 (N_13239,N_12845,N_12516);
nand U13240 (N_13240,N_12938,N_12982);
and U13241 (N_13241,N_12765,N_12950);
nand U13242 (N_13242,N_12500,N_12731);
xnor U13243 (N_13243,N_12595,N_12525);
nand U13244 (N_13244,N_12581,N_12923);
or U13245 (N_13245,N_12756,N_12915);
nand U13246 (N_13246,N_12838,N_12824);
and U13247 (N_13247,N_12753,N_12801);
xor U13248 (N_13248,N_12813,N_12640);
nor U13249 (N_13249,N_12705,N_12727);
nand U13250 (N_13250,N_12758,N_12852);
xor U13251 (N_13251,N_12580,N_12773);
nor U13252 (N_13252,N_12967,N_12694);
and U13253 (N_13253,N_12654,N_12925);
xnor U13254 (N_13254,N_12517,N_12710);
xnor U13255 (N_13255,N_12958,N_12755);
nand U13256 (N_13256,N_12885,N_12766);
xor U13257 (N_13257,N_12687,N_12847);
xor U13258 (N_13258,N_12811,N_12812);
xnor U13259 (N_13259,N_12865,N_12517);
or U13260 (N_13260,N_12756,N_12659);
nand U13261 (N_13261,N_12929,N_12524);
nand U13262 (N_13262,N_12745,N_12838);
and U13263 (N_13263,N_12937,N_12737);
xor U13264 (N_13264,N_12847,N_12866);
nand U13265 (N_13265,N_12804,N_12548);
and U13266 (N_13266,N_12854,N_12745);
nor U13267 (N_13267,N_12586,N_12868);
nand U13268 (N_13268,N_12654,N_12693);
xor U13269 (N_13269,N_12618,N_12542);
nor U13270 (N_13270,N_12990,N_12856);
nand U13271 (N_13271,N_12711,N_12969);
or U13272 (N_13272,N_12930,N_12590);
and U13273 (N_13273,N_12731,N_12667);
nor U13274 (N_13274,N_12980,N_12552);
or U13275 (N_13275,N_12577,N_12811);
nand U13276 (N_13276,N_12654,N_12790);
nand U13277 (N_13277,N_12828,N_12569);
xor U13278 (N_13278,N_12889,N_12679);
nand U13279 (N_13279,N_12911,N_12921);
and U13280 (N_13280,N_12688,N_12580);
or U13281 (N_13281,N_12869,N_12699);
xnor U13282 (N_13282,N_12622,N_12910);
xnor U13283 (N_13283,N_12890,N_12782);
xor U13284 (N_13284,N_12783,N_12983);
nor U13285 (N_13285,N_12967,N_12514);
or U13286 (N_13286,N_12830,N_12743);
nor U13287 (N_13287,N_12606,N_12570);
xor U13288 (N_13288,N_12664,N_12732);
nand U13289 (N_13289,N_12667,N_12729);
nor U13290 (N_13290,N_12602,N_12607);
and U13291 (N_13291,N_12816,N_12701);
nor U13292 (N_13292,N_12951,N_12891);
nand U13293 (N_13293,N_12633,N_12745);
nor U13294 (N_13294,N_12647,N_12948);
and U13295 (N_13295,N_12948,N_12898);
nor U13296 (N_13296,N_12634,N_12537);
nor U13297 (N_13297,N_12707,N_12971);
or U13298 (N_13298,N_12627,N_12832);
and U13299 (N_13299,N_12633,N_12763);
and U13300 (N_13300,N_12508,N_12914);
xnor U13301 (N_13301,N_12905,N_12605);
xnor U13302 (N_13302,N_12686,N_12977);
nor U13303 (N_13303,N_12670,N_12834);
or U13304 (N_13304,N_12540,N_12782);
or U13305 (N_13305,N_12623,N_12756);
nor U13306 (N_13306,N_12962,N_12559);
nand U13307 (N_13307,N_12721,N_12504);
and U13308 (N_13308,N_12758,N_12523);
or U13309 (N_13309,N_12840,N_12841);
nand U13310 (N_13310,N_12674,N_12518);
nand U13311 (N_13311,N_12755,N_12909);
or U13312 (N_13312,N_12708,N_12728);
xnor U13313 (N_13313,N_12630,N_12955);
xnor U13314 (N_13314,N_12525,N_12861);
or U13315 (N_13315,N_12596,N_12725);
or U13316 (N_13316,N_12506,N_12724);
nand U13317 (N_13317,N_12823,N_12654);
xor U13318 (N_13318,N_12519,N_12891);
nor U13319 (N_13319,N_12691,N_12802);
nand U13320 (N_13320,N_12941,N_12905);
or U13321 (N_13321,N_12927,N_12998);
and U13322 (N_13322,N_12571,N_12891);
xor U13323 (N_13323,N_12952,N_12567);
or U13324 (N_13324,N_12857,N_12670);
xnor U13325 (N_13325,N_12837,N_12624);
or U13326 (N_13326,N_12963,N_12761);
nand U13327 (N_13327,N_12997,N_12600);
nor U13328 (N_13328,N_12579,N_12649);
and U13329 (N_13329,N_12771,N_12953);
or U13330 (N_13330,N_12580,N_12796);
and U13331 (N_13331,N_12889,N_12774);
and U13332 (N_13332,N_12877,N_12605);
nor U13333 (N_13333,N_12666,N_12940);
xnor U13334 (N_13334,N_12647,N_12779);
or U13335 (N_13335,N_12706,N_12973);
nand U13336 (N_13336,N_12815,N_12626);
nand U13337 (N_13337,N_12752,N_12651);
and U13338 (N_13338,N_12664,N_12809);
and U13339 (N_13339,N_12526,N_12791);
nand U13340 (N_13340,N_12702,N_12845);
nand U13341 (N_13341,N_12934,N_12831);
nor U13342 (N_13342,N_12933,N_12951);
or U13343 (N_13343,N_12594,N_12579);
or U13344 (N_13344,N_12813,N_12730);
nor U13345 (N_13345,N_12633,N_12657);
nand U13346 (N_13346,N_12649,N_12767);
and U13347 (N_13347,N_12890,N_12536);
or U13348 (N_13348,N_12680,N_12816);
xnor U13349 (N_13349,N_12554,N_12594);
xor U13350 (N_13350,N_12852,N_12896);
nand U13351 (N_13351,N_12622,N_12788);
and U13352 (N_13352,N_12732,N_12752);
nor U13353 (N_13353,N_12879,N_12636);
xnor U13354 (N_13354,N_12917,N_12928);
nand U13355 (N_13355,N_12503,N_12868);
or U13356 (N_13356,N_12979,N_12688);
nor U13357 (N_13357,N_12851,N_12853);
nor U13358 (N_13358,N_12747,N_12920);
and U13359 (N_13359,N_12826,N_12996);
nor U13360 (N_13360,N_12669,N_12771);
and U13361 (N_13361,N_12667,N_12876);
nor U13362 (N_13362,N_12850,N_12640);
xor U13363 (N_13363,N_12675,N_12922);
nand U13364 (N_13364,N_12829,N_12634);
and U13365 (N_13365,N_12916,N_12812);
and U13366 (N_13366,N_12538,N_12748);
nor U13367 (N_13367,N_12876,N_12598);
xor U13368 (N_13368,N_12722,N_12529);
or U13369 (N_13369,N_12843,N_12635);
xnor U13370 (N_13370,N_12864,N_12506);
or U13371 (N_13371,N_12727,N_12526);
and U13372 (N_13372,N_12989,N_12901);
or U13373 (N_13373,N_12803,N_12762);
and U13374 (N_13374,N_12921,N_12761);
xor U13375 (N_13375,N_12755,N_12650);
or U13376 (N_13376,N_12880,N_12652);
or U13377 (N_13377,N_12659,N_12905);
and U13378 (N_13378,N_12875,N_12546);
nand U13379 (N_13379,N_12923,N_12701);
xnor U13380 (N_13380,N_12725,N_12877);
nor U13381 (N_13381,N_12914,N_12883);
nand U13382 (N_13382,N_12585,N_12747);
nand U13383 (N_13383,N_12781,N_12714);
nor U13384 (N_13384,N_12624,N_12664);
nand U13385 (N_13385,N_12753,N_12654);
nor U13386 (N_13386,N_12752,N_12904);
and U13387 (N_13387,N_12705,N_12668);
and U13388 (N_13388,N_12631,N_12630);
nor U13389 (N_13389,N_12633,N_12917);
and U13390 (N_13390,N_12778,N_12903);
nand U13391 (N_13391,N_12988,N_12960);
xnor U13392 (N_13392,N_12750,N_12799);
and U13393 (N_13393,N_12501,N_12828);
or U13394 (N_13394,N_12740,N_12884);
nand U13395 (N_13395,N_12876,N_12811);
and U13396 (N_13396,N_12630,N_12829);
xor U13397 (N_13397,N_12750,N_12733);
or U13398 (N_13398,N_12998,N_12598);
or U13399 (N_13399,N_12773,N_12636);
xor U13400 (N_13400,N_12655,N_12819);
xor U13401 (N_13401,N_12546,N_12644);
or U13402 (N_13402,N_12821,N_12861);
xor U13403 (N_13403,N_12588,N_12548);
nand U13404 (N_13404,N_12753,N_12560);
and U13405 (N_13405,N_12977,N_12773);
and U13406 (N_13406,N_12567,N_12673);
nor U13407 (N_13407,N_12534,N_12604);
xnor U13408 (N_13408,N_12851,N_12798);
nand U13409 (N_13409,N_12969,N_12551);
nor U13410 (N_13410,N_12980,N_12984);
or U13411 (N_13411,N_12556,N_12819);
xnor U13412 (N_13412,N_12663,N_12608);
or U13413 (N_13413,N_12787,N_12866);
and U13414 (N_13414,N_12731,N_12952);
xnor U13415 (N_13415,N_12976,N_12528);
xor U13416 (N_13416,N_12570,N_12500);
nor U13417 (N_13417,N_12897,N_12659);
or U13418 (N_13418,N_12895,N_12622);
nor U13419 (N_13419,N_12509,N_12598);
and U13420 (N_13420,N_12918,N_12800);
or U13421 (N_13421,N_12737,N_12757);
nand U13422 (N_13422,N_12977,N_12946);
nand U13423 (N_13423,N_12714,N_12937);
xor U13424 (N_13424,N_12969,N_12810);
nand U13425 (N_13425,N_12939,N_12592);
nand U13426 (N_13426,N_12921,N_12746);
or U13427 (N_13427,N_12709,N_12699);
nand U13428 (N_13428,N_12540,N_12967);
and U13429 (N_13429,N_12539,N_12989);
or U13430 (N_13430,N_12560,N_12562);
or U13431 (N_13431,N_12610,N_12899);
nand U13432 (N_13432,N_12631,N_12549);
nand U13433 (N_13433,N_12554,N_12879);
nor U13434 (N_13434,N_12935,N_12608);
or U13435 (N_13435,N_12667,N_12742);
nand U13436 (N_13436,N_12804,N_12906);
nand U13437 (N_13437,N_12808,N_12572);
nand U13438 (N_13438,N_12797,N_12659);
and U13439 (N_13439,N_12923,N_12669);
and U13440 (N_13440,N_12539,N_12803);
nand U13441 (N_13441,N_12746,N_12803);
nand U13442 (N_13442,N_12914,N_12706);
and U13443 (N_13443,N_12639,N_12914);
nand U13444 (N_13444,N_12552,N_12716);
or U13445 (N_13445,N_12707,N_12800);
xor U13446 (N_13446,N_12902,N_12863);
xnor U13447 (N_13447,N_12727,N_12557);
nand U13448 (N_13448,N_12585,N_12730);
or U13449 (N_13449,N_12975,N_12941);
and U13450 (N_13450,N_12589,N_12852);
and U13451 (N_13451,N_12859,N_12880);
or U13452 (N_13452,N_12832,N_12883);
xor U13453 (N_13453,N_12655,N_12710);
and U13454 (N_13454,N_12887,N_12757);
or U13455 (N_13455,N_12825,N_12512);
and U13456 (N_13456,N_12759,N_12724);
xnor U13457 (N_13457,N_12531,N_12906);
xor U13458 (N_13458,N_12566,N_12929);
or U13459 (N_13459,N_12724,N_12899);
nand U13460 (N_13460,N_12800,N_12566);
and U13461 (N_13461,N_12779,N_12762);
xor U13462 (N_13462,N_12870,N_12813);
and U13463 (N_13463,N_12969,N_12895);
and U13464 (N_13464,N_12759,N_12653);
and U13465 (N_13465,N_12699,N_12570);
xnor U13466 (N_13466,N_12973,N_12940);
nand U13467 (N_13467,N_12709,N_12509);
nand U13468 (N_13468,N_12682,N_12753);
nor U13469 (N_13469,N_12547,N_12960);
and U13470 (N_13470,N_12510,N_12724);
nand U13471 (N_13471,N_12978,N_12922);
and U13472 (N_13472,N_12966,N_12900);
nor U13473 (N_13473,N_12513,N_12634);
and U13474 (N_13474,N_12724,N_12733);
nand U13475 (N_13475,N_12631,N_12917);
xor U13476 (N_13476,N_12675,N_12696);
and U13477 (N_13477,N_12901,N_12624);
or U13478 (N_13478,N_12547,N_12986);
and U13479 (N_13479,N_12570,N_12931);
xnor U13480 (N_13480,N_12831,N_12729);
xor U13481 (N_13481,N_12869,N_12794);
nor U13482 (N_13482,N_12841,N_12664);
xor U13483 (N_13483,N_12668,N_12617);
xnor U13484 (N_13484,N_12848,N_12713);
xor U13485 (N_13485,N_12747,N_12863);
nor U13486 (N_13486,N_12557,N_12835);
nor U13487 (N_13487,N_12945,N_12528);
xor U13488 (N_13488,N_12782,N_12918);
xor U13489 (N_13489,N_12865,N_12653);
or U13490 (N_13490,N_12546,N_12533);
xor U13491 (N_13491,N_12699,N_12820);
or U13492 (N_13492,N_12746,N_12876);
nand U13493 (N_13493,N_12851,N_12608);
and U13494 (N_13494,N_12759,N_12560);
nor U13495 (N_13495,N_12831,N_12639);
nor U13496 (N_13496,N_12923,N_12823);
nand U13497 (N_13497,N_12539,N_12740);
or U13498 (N_13498,N_12896,N_12967);
xor U13499 (N_13499,N_12698,N_12502);
xnor U13500 (N_13500,N_13016,N_13073);
nand U13501 (N_13501,N_13114,N_13394);
and U13502 (N_13502,N_13353,N_13191);
or U13503 (N_13503,N_13198,N_13406);
xor U13504 (N_13504,N_13455,N_13041);
nand U13505 (N_13505,N_13169,N_13117);
or U13506 (N_13506,N_13089,N_13452);
and U13507 (N_13507,N_13399,N_13082);
nor U13508 (N_13508,N_13499,N_13358);
or U13509 (N_13509,N_13087,N_13387);
nor U13510 (N_13510,N_13433,N_13485);
nand U13511 (N_13511,N_13088,N_13175);
or U13512 (N_13512,N_13483,N_13246);
and U13513 (N_13513,N_13419,N_13252);
or U13514 (N_13514,N_13446,N_13423);
nand U13515 (N_13515,N_13472,N_13075);
nand U13516 (N_13516,N_13030,N_13035);
or U13517 (N_13517,N_13385,N_13445);
nor U13518 (N_13518,N_13068,N_13340);
xor U13519 (N_13519,N_13069,N_13158);
or U13520 (N_13520,N_13378,N_13171);
nor U13521 (N_13521,N_13355,N_13392);
xnor U13522 (N_13522,N_13102,N_13360);
nand U13523 (N_13523,N_13427,N_13498);
or U13524 (N_13524,N_13202,N_13197);
and U13525 (N_13525,N_13457,N_13221);
and U13526 (N_13526,N_13413,N_13245);
xor U13527 (N_13527,N_13217,N_13255);
nand U13528 (N_13528,N_13134,N_13265);
nor U13529 (N_13529,N_13418,N_13441);
xnor U13530 (N_13530,N_13228,N_13361);
nor U13531 (N_13531,N_13193,N_13173);
nor U13532 (N_13532,N_13282,N_13319);
nand U13533 (N_13533,N_13379,N_13357);
and U13534 (N_13534,N_13318,N_13047);
nand U13535 (N_13535,N_13150,N_13425);
nand U13536 (N_13536,N_13291,N_13298);
nand U13537 (N_13537,N_13074,N_13183);
xor U13538 (N_13538,N_13060,N_13464);
nand U13539 (N_13539,N_13129,N_13316);
xor U13540 (N_13540,N_13206,N_13231);
and U13541 (N_13541,N_13421,N_13218);
or U13542 (N_13542,N_13454,N_13147);
nand U13543 (N_13543,N_13048,N_13222);
nand U13544 (N_13544,N_13177,N_13466);
and U13545 (N_13545,N_13244,N_13366);
nand U13546 (N_13546,N_13465,N_13410);
xor U13547 (N_13547,N_13431,N_13056);
nor U13548 (N_13548,N_13157,N_13142);
and U13549 (N_13549,N_13474,N_13404);
or U13550 (N_13550,N_13420,N_13154);
nand U13551 (N_13551,N_13438,N_13343);
nor U13552 (N_13552,N_13072,N_13451);
or U13553 (N_13553,N_13091,N_13223);
nand U13554 (N_13554,N_13032,N_13288);
nand U13555 (N_13555,N_13324,N_13015);
or U13556 (N_13556,N_13260,N_13444);
xor U13557 (N_13557,N_13309,N_13388);
nor U13558 (N_13558,N_13494,N_13403);
nand U13559 (N_13559,N_13144,N_13257);
xnor U13560 (N_13560,N_13335,N_13416);
and U13561 (N_13561,N_13492,N_13149);
or U13562 (N_13562,N_13266,N_13262);
and U13563 (N_13563,N_13407,N_13098);
or U13564 (N_13564,N_13373,N_13128);
nor U13565 (N_13565,N_13365,N_13468);
or U13566 (N_13566,N_13043,N_13185);
nor U13567 (N_13567,N_13151,N_13188);
and U13568 (N_13568,N_13342,N_13462);
xnor U13569 (N_13569,N_13473,N_13167);
nor U13570 (N_13570,N_13141,N_13215);
nor U13571 (N_13571,N_13352,N_13139);
nand U13572 (N_13572,N_13058,N_13414);
and U13573 (N_13573,N_13107,N_13417);
and U13574 (N_13574,N_13000,N_13349);
or U13575 (N_13575,N_13010,N_13160);
or U13576 (N_13576,N_13004,N_13039);
xor U13577 (N_13577,N_13009,N_13350);
or U13578 (N_13578,N_13315,N_13268);
nand U13579 (N_13579,N_13205,N_13290);
or U13580 (N_13580,N_13234,N_13354);
or U13581 (N_13581,N_13249,N_13334);
xnor U13582 (N_13582,N_13259,N_13370);
nor U13583 (N_13583,N_13179,N_13371);
nor U13584 (N_13584,N_13061,N_13121);
nand U13585 (N_13585,N_13375,N_13051);
nor U13586 (N_13586,N_13220,N_13148);
nor U13587 (N_13587,N_13180,N_13037);
xnor U13588 (N_13588,N_13022,N_13155);
or U13589 (N_13589,N_13424,N_13094);
or U13590 (N_13590,N_13428,N_13463);
nor U13591 (N_13591,N_13241,N_13118);
xnor U13592 (N_13592,N_13376,N_13402);
nand U13593 (N_13593,N_13186,N_13277);
nor U13594 (N_13594,N_13001,N_13014);
or U13595 (N_13595,N_13430,N_13070);
or U13596 (N_13596,N_13442,N_13256);
xor U13597 (N_13597,N_13124,N_13081);
nor U13598 (N_13598,N_13484,N_13274);
xor U13599 (N_13599,N_13284,N_13026);
and U13600 (N_13600,N_13329,N_13338);
nand U13601 (N_13601,N_13239,N_13278);
nor U13602 (N_13602,N_13398,N_13034);
or U13603 (N_13603,N_13495,N_13201);
or U13604 (N_13604,N_13140,N_13331);
xor U13605 (N_13605,N_13242,N_13025);
or U13606 (N_13606,N_13367,N_13018);
nor U13607 (N_13607,N_13199,N_13136);
or U13608 (N_13608,N_13095,N_13369);
nor U13609 (N_13609,N_13103,N_13076);
nand U13610 (N_13610,N_13168,N_13122);
or U13611 (N_13611,N_13165,N_13384);
and U13612 (N_13612,N_13045,N_13449);
and U13613 (N_13613,N_13253,N_13490);
nor U13614 (N_13614,N_13006,N_13044);
xnor U13615 (N_13615,N_13194,N_13382);
xnor U13616 (N_13616,N_13408,N_13286);
nand U13617 (N_13617,N_13381,N_13055);
and U13618 (N_13618,N_13182,N_13327);
nor U13619 (N_13619,N_13111,N_13207);
and U13620 (N_13620,N_13469,N_13448);
xnor U13621 (N_13621,N_13372,N_13187);
xor U13622 (N_13622,N_13012,N_13063);
nand U13623 (N_13623,N_13023,N_13115);
and U13624 (N_13624,N_13303,N_13166);
nand U13625 (N_13625,N_13325,N_13459);
or U13626 (N_13626,N_13059,N_13235);
or U13627 (N_13627,N_13078,N_13040);
nand U13628 (N_13628,N_13323,N_13196);
nor U13629 (N_13629,N_13250,N_13003);
xnor U13630 (N_13630,N_13028,N_13109);
nor U13631 (N_13631,N_13271,N_13108);
nand U13632 (N_13632,N_13152,N_13321);
or U13633 (N_13633,N_13460,N_13204);
xnor U13634 (N_13634,N_13304,N_13377);
nand U13635 (N_13635,N_13176,N_13052);
or U13636 (N_13636,N_13174,N_13208);
xor U13637 (N_13637,N_13230,N_13079);
xor U13638 (N_13638,N_13224,N_13393);
nand U13639 (N_13639,N_13293,N_13251);
and U13640 (N_13640,N_13153,N_13347);
nor U13641 (N_13641,N_13337,N_13137);
xor U13642 (N_13642,N_13192,N_13471);
nor U13643 (N_13643,N_13247,N_13062);
and U13644 (N_13644,N_13272,N_13054);
nand U13645 (N_13645,N_13294,N_13363);
or U13646 (N_13646,N_13049,N_13437);
xor U13647 (N_13647,N_13359,N_13119);
or U13648 (N_13648,N_13033,N_13066);
nand U13649 (N_13649,N_13046,N_13164);
nand U13650 (N_13650,N_13042,N_13105);
or U13651 (N_13651,N_13031,N_13064);
xor U13652 (N_13652,N_13050,N_13211);
and U13653 (N_13653,N_13306,N_13456);
nor U13654 (N_13654,N_13374,N_13415);
nor U13655 (N_13655,N_13112,N_13090);
nand U13656 (N_13656,N_13322,N_13085);
nor U13657 (N_13657,N_13328,N_13496);
xor U13658 (N_13658,N_13497,N_13440);
nor U13659 (N_13659,N_13178,N_13226);
xnor U13660 (N_13660,N_13096,N_13383);
or U13661 (N_13661,N_13219,N_13493);
xnor U13662 (N_13662,N_13362,N_13132);
or U13663 (N_13663,N_13084,N_13283);
or U13664 (N_13664,N_13432,N_13131);
or U13665 (N_13665,N_13475,N_13116);
xor U13666 (N_13666,N_13138,N_13299);
or U13667 (N_13667,N_13297,N_13320);
nand U13668 (N_13668,N_13332,N_13080);
or U13669 (N_13669,N_13229,N_13212);
xnor U13670 (N_13670,N_13238,N_13341);
or U13671 (N_13671,N_13214,N_13233);
and U13672 (N_13672,N_13317,N_13227);
and U13673 (N_13673,N_13021,N_13281);
and U13674 (N_13674,N_13163,N_13287);
and U13675 (N_13675,N_13036,N_13435);
or U13676 (N_13676,N_13296,N_13289);
xor U13677 (N_13677,N_13336,N_13110);
xor U13678 (N_13678,N_13491,N_13275);
xnor U13679 (N_13679,N_13305,N_13077);
and U13680 (N_13680,N_13237,N_13225);
or U13681 (N_13681,N_13184,N_13086);
nand U13682 (N_13682,N_13308,N_13434);
or U13683 (N_13683,N_13017,N_13400);
or U13684 (N_13684,N_13190,N_13461);
and U13685 (N_13685,N_13130,N_13389);
or U13686 (N_13686,N_13146,N_13487);
and U13687 (N_13687,N_13189,N_13172);
xor U13688 (N_13688,N_13326,N_13007);
xnor U13689 (N_13689,N_13307,N_13002);
nor U13690 (N_13690,N_13312,N_13258);
nand U13691 (N_13691,N_13436,N_13248);
and U13692 (N_13692,N_13203,N_13450);
xnor U13693 (N_13693,N_13093,N_13467);
nor U13694 (N_13694,N_13135,N_13264);
nand U13695 (N_13695,N_13008,N_13005);
or U13696 (N_13696,N_13270,N_13019);
xnor U13697 (N_13697,N_13443,N_13422);
xnor U13698 (N_13698,N_13453,N_13020);
or U13699 (N_13699,N_13458,N_13314);
and U13700 (N_13700,N_13162,N_13330);
or U13701 (N_13701,N_13083,N_13477);
nand U13702 (N_13702,N_13292,N_13344);
nand U13703 (N_13703,N_13395,N_13209);
and U13704 (N_13704,N_13267,N_13127);
or U13705 (N_13705,N_13302,N_13156);
nand U13706 (N_13706,N_13478,N_13261);
and U13707 (N_13707,N_13368,N_13333);
nand U13708 (N_13708,N_13024,N_13311);
xnor U13709 (N_13709,N_13067,N_13126);
nand U13710 (N_13710,N_13280,N_13489);
and U13711 (N_13711,N_13101,N_13285);
xor U13712 (N_13712,N_13488,N_13345);
or U13713 (N_13713,N_13300,N_13439);
xnor U13714 (N_13714,N_13348,N_13429);
nand U13715 (N_13715,N_13346,N_13411);
or U13716 (N_13716,N_13351,N_13479);
or U13717 (N_13717,N_13390,N_13380);
nor U13718 (N_13718,N_13027,N_13313);
nor U13719 (N_13719,N_13481,N_13013);
or U13720 (N_13720,N_13254,N_13210);
or U13721 (N_13721,N_13071,N_13405);
nor U13722 (N_13722,N_13123,N_13470);
or U13723 (N_13723,N_13486,N_13447);
or U13724 (N_13724,N_13143,N_13029);
nand U13725 (N_13725,N_13181,N_13243);
nand U13726 (N_13726,N_13240,N_13113);
nand U13727 (N_13727,N_13480,N_13263);
or U13728 (N_13728,N_13145,N_13161);
and U13729 (N_13729,N_13310,N_13213);
and U13730 (N_13730,N_13396,N_13159);
or U13731 (N_13731,N_13279,N_13100);
xor U13732 (N_13732,N_13301,N_13391);
nand U13733 (N_13733,N_13106,N_13397);
nor U13734 (N_13734,N_13038,N_13133);
or U13735 (N_13735,N_13057,N_13065);
nor U13736 (N_13736,N_13386,N_13236);
nand U13737 (N_13737,N_13273,N_13276);
xor U13738 (N_13738,N_13092,N_13232);
and U13739 (N_13739,N_13295,N_13482);
nand U13740 (N_13740,N_13195,N_13120);
nand U13741 (N_13741,N_13125,N_13104);
or U13742 (N_13742,N_13200,N_13412);
nor U13743 (N_13743,N_13170,N_13476);
xor U13744 (N_13744,N_13401,N_13216);
and U13745 (N_13745,N_13269,N_13053);
nand U13746 (N_13746,N_13364,N_13011);
and U13747 (N_13747,N_13426,N_13339);
and U13748 (N_13748,N_13097,N_13356);
and U13749 (N_13749,N_13099,N_13409);
and U13750 (N_13750,N_13194,N_13460);
nand U13751 (N_13751,N_13179,N_13301);
nand U13752 (N_13752,N_13117,N_13192);
and U13753 (N_13753,N_13297,N_13015);
and U13754 (N_13754,N_13205,N_13071);
xnor U13755 (N_13755,N_13484,N_13198);
or U13756 (N_13756,N_13406,N_13019);
xor U13757 (N_13757,N_13446,N_13286);
nand U13758 (N_13758,N_13300,N_13111);
xnor U13759 (N_13759,N_13238,N_13047);
or U13760 (N_13760,N_13264,N_13123);
nor U13761 (N_13761,N_13151,N_13460);
xnor U13762 (N_13762,N_13114,N_13463);
and U13763 (N_13763,N_13427,N_13181);
and U13764 (N_13764,N_13274,N_13423);
xnor U13765 (N_13765,N_13131,N_13319);
nand U13766 (N_13766,N_13184,N_13072);
or U13767 (N_13767,N_13193,N_13055);
and U13768 (N_13768,N_13492,N_13243);
or U13769 (N_13769,N_13021,N_13209);
or U13770 (N_13770,N_13477,N_13496);
or U13771 (N_13771,N_13120,N_13077);
or U13772 (N_13772,N_13227,N_13331);
and U13773 (N_13773,N_13478,N_13321);
or U13774 (N_13774,N_13458,N_13496);
and U13775 (N_13775,N_13220,N_13375);
or U13776 (N_13776,N_13050,N_13269);
and U13777 (N_13777,N_13237,N_13050);
xor U13778 (N_13778,N_13019,N_13152);
and U13779 (N_13779,N_13279,N_13019);
and U13780 (N_13780,N_13434,N_13278);
or U13781 (N_13781,N_13151,N_13377);
xor U13782 (N_13782,N_13412,N_13112);
nand U13783 (N_13783,N_13238,N_13070);
nand U13784 (N_13784,N_13316,N_13119);
xnor U13785 (N_13785,N_13108,N_13015);
or U13786 (N_13786,N_13292,N_13418);
xor U13787 (N_13787,N_13403,N_13247);
or U13788 (N_13788,N_13414,N_13230);
nor U13789 (N_13789,N_13132,N_13268);
nor U13790 (N_13790,N_13215,N_13241);
or U13791 (N_13791,N_13291,N_13470);
nand U13792 (N_13792,N_13202,N_13478);
nand U13793 (N_13793,N_13430,N_13476);
nand U13794 (N_13794,N_13094,N_13152);
nand U13795 (N_13795,N_13197,N_13315);
xnor U13796 (N_13796,N_13319,N_13022);
xnor U13797 (N_13797,N_13449,N_13122);
or U13798 (N_13798,N_13404,N_13145);
or U13799 (N_13799,N_13331,N_13124);
nand U13800 (N_13800,N_13251,N_13245);
nand U13801 (N_13801,N_13363,N_13454);
and U13802 (N_13802,N_13301,N_13127);
nor U13803 (N_13803,N_13077,N_13045);
nand U13804 (N_13804,N_13105,N_13220);
nand U13805 (N_13805,N_13422,N_13276);
or U13806 (N_13806,N_13112,N_13464);
xnor U13807 (N_13807,N_13432,N_13247);
or U13808 (N_13808,N_13133,N_13149);
nand U13809 (N_13809,N_13358,N_13050);
nand U13810 (N_13810,N_13043,N_13318);
or U13811 (N_13811,N_13255,N_13154);
and U13812 (N_13812,N_13044,N_13026);
nand U13813 (N_13813,N_13262,N_13109);
nor U13814 (N_13814,N_13282,N_13111);
or U13815 (N_13815,N_13298,N_13168);
and U13816 (N_13816,N_13238,N_13073);
xnor U13817 (N_13817,N_13382,N_13258);
xnor U13818 (N_13818,N_13250,N_13359);
and U13819 (N_13819,N_13483,N_13288);
nand U13820 (N_13820,N_13166,N_13049);
nand U13821 (N_13821,N_13436,N_13192);
or U13822 (N_13822,N_13295,N_13281);
or U13823 (N_13823,N_13069,N_13042);
and U13824 (N_13824,N_13178,N_13317);
xnor U13825 (N_13825,N_13206,N_13021);
and U13826 (N_13826,N_13156,N_13317);
nor U13827 (N_13827,N_13308,N_13028);
or U13828 (N_13828,N_13057,N_13372);
nor U13829 (N_13829,N_13338,N_13317);
or U13830 (N_13830,N_13315,N_13139);
or U13831 (N_13831,N_13212,N_13088);
and U13832 (N_13832,N_13490,N_13120);
or U13833 (N_13833,N_13280,N_13072);
or U13834 (N_13834,N_13423,N_13235);
nor U13835 (N_13835,N_13098,N_13232);
xnor U13836 (N_13836,N_13115,N_13241);
nand U13837 (N_13837,N_13430,N_13356);
or U13838 (N_13838,N_13374,N_13237);
nor U13839 (N_13839,N_13119,N_13389);
and U13840 (N_13840,N_13073,N_13497);
nor U13841 (N_13841,N_13207,N_13412);
xnor U13842 (N_13842,N_13146,N_13295);
xnor U13843 (N_13843,N_13156,N_13350);
or U13844 (N_13844,N_13164,N_13179);
and U13845 (N_13845,N_13091,N_13089);
xnor U13846 (N_13846,N_13127,N_13114);
nand U13847 (N_13847,N_13238,N_13264);
nand U13848 (N_13848,N_13170,N_13482);
nor U13849 (N_13849,N_13446,N_13065);
nor U13850 (N_13850,N_13373,N_13349);
nor U13851 (N_13851,N_13000,N_13085);
nor U13852 (N_13852,N_13352,N_13279);
and U13853 (N_13853,N_13338,N_13091);
xnor U13854 (N_13854,N_13067,N_13121);
or U13855 (N_13855,N_13310,N_13016);
nor U13856 (N_13856,N_13367,N_13219);
nand U13857 (N_13857,N_13121,N_13080);
and U13858 (N_13858,N_13448,N_13106);
xor U13859 (N_13859,N_13440,N_13080);
and U13860 (N_13860,N_13049,N_13310);
nor U13861 (N_13861,N_13236,N_13273);
or U13862 (N_13862,N_13474,N_13350);
and U13863 (N_13863,N_13446,N_13233);
nor U13864 (N_13864,N_13185,N_13268);
nor U13865 (N_13865,N_13453,N_13176);
nor U13866 (N_13866,N_13299,N_13482);
and U13867 (N_13867,N_13295,N_13110);
nand U13868 (N_13868,N_13099,N_13407);
or U13869 (N_13869,N_13257,N_13209);
xor U13870 (N_13870,N_13293,N_13360);
or U13871 (N_13871,N_13109,N_13048);
nand U13872 (N_13872,N_13009,N_13357);
nand U13873 (N_13873,N_13273,N_13440);
xnor U13874 (N_13874,N_13354,N_13108);
nand U13875 (N_13875,N_13423,N_13382);
or U13876 (N_13876,N_13459,N_13202);
nor U13877 (N_13877,N_13001,N_13191);
nor U13878 (N_13878,N_13017,N_13482);
or U13879 (N_13879,N_13034,N_13061);
nand U13880 (N_13880,N_13099,N_13274);
or U13881 (N_13881,N_13032,N_13151);
and U13882 (N_13882,N_13260,N_13418);
and U13883 (N_13883,N_13130,N_13018);
xnor U13884 (N_13884,N_13317,N_13305);
nor U13885 (N_13885,N_13116,N_13349);
xor U13886 (N_13886,N_13366,N_13266);
or U13887 (N_13887,N_13069,N_13084);
and U13888 (N_13888,N_13175,N_13372);
and U13889 (N_13889,N_13334,N_13022);
nor U13890 (N_13890,N_13304,N_13477);
xor U13891 (N_13891,N_13292,N_13346);
and U13892 (N_13892,N_13257,N_13022);
nand U13893 (N_13893,N_13097,N_13016);
and U13894 (N_13894,N_13438,N_13117);
xnor U13895 (N_13895,N_13400,N_13166);
nand U13896 (N_13896,N_13272,N_13299);
xnor U13897 (N_13897,N_13055,N_13076);
nand U13898 (N_13898,N_13053,N_13411);
xor U13899 (N_13899,N_13113,N_13042);
or U13900 (N_13900,N_13178,N_13314);
or U13901 (N_13901,N_13173,N_13103);
xnor U13902 (N_13902,N_13353,N_13141);
xnor U13903 (N_13903,N_13300,N_13061);
xnor U13904 (N_13904,N_13485,N_13157);
nor U13905 (N_13905,N_13468,N_13324);
or U13906 (N_13906,N_13227,N_13026);
or U13907 (N_13907,N_13483,N_13195);
xor U13908 (N_13908,N_13209,N_13172);
xor U13909 (N_13909,N_13191,N_13204);
or U13910 (N_13910,N_13317,N_13208);
xor U13911 (N_13911,N_13149,N_13314);
nor U13912 (N_13912,N_13136,N_13279);
or U13913 (N_13913,N_13098,N_13287);
xor U13914 (N_13914,N_13438,N_13460);
nor U13915 (N_13915,N_13231,N_13075);
and U13916 (N_13916,N_13165,N_13275);
nor U13917 (N_13917,N_13286,N_13299);
or U13918 (N_13918,N_13396,N_13161);
nor U13919 (N_13919,N_13189,N_13471);
nand U13920 (N_13920,N_13450,N_13151);
nor U13921 (N_13921,N_13463,N_13287);
xnor U13922 (N_13922,N_13214,N_13380);
nand U13923 (N_13923,N_13145,N_13413);
xor U13924 (N_13924,N_13368,N_13307);
xor U13925 (N_13925,N_13376,N_13156);
xor U13926 (N_13926,N_13312,N_13494);
and U13927 (N_13927,N_13252,N_13161);
nor U13928 (N_13928,N_13127,N_13247);
or U13929 (N_13929,N_13182,N_13413);
xor U13930 (N_13930,N_13292,N_13017);
or U13931 (N_13931,N_13236,N_13086);
and U13932 (N_13932,N_13332,N_13437);
xor U13933 (N_13933,N_13164,N_13420);
nand U13934 (N_13934,N_13417,N_13385);
nand U13935 (N_13935,N_13264,N_13362);
and U13936 (N_13936,N_13343,N_13464);
nor U13937 (N_13937,N_13361,N_13486);
and U13938 (N_13938,N_13278,N_13007);
and U13939 (N_13939,N_13373,N_13027);
nor U13940 (N_13940,N_13029,N_13349);
nor U13941 (N_13941,N_13483,N_13373);
or U13942 (N_13942,N_13160,N_13056);
and U13943 (N_13943,N_13180,N_13111);
and U13944 (N_13944,N_13483,N_13181);
nand U13945 (N_13945,N_13304,N_13329);
and U13946 (N_13946,N_13120,N_13420);
nor U13947 (N_13947,N_13373,N_13196);
nor U13948 (N_13948,N_13367,N_13180);
nand U13949 (N_13949,N_13150,N_13448);
or U13950 (N_13950,N_13235,N_13334);
and U13951 (N_13951,N_13213,N_13332);
nand U13952 (N_13952,N_13463,N_13124);
nor U13953 (N_13953,N_13112,N_13056);
and U13954 (N_13954,N_13007,N_13180);
or U13955 (N_13955,N_13378,N_13106);
xnor U13956 (N_13956,N_13422,N_13231);
nor U13957 (N_13957,N_13095,N_13460);
nand U13958 (N_13958,N_13115,N_13110);
and U13959 (N_13959,N_13316,N_13130);
and U13960 (N_13960,N_13185,N_13322);
xnor U13961 (N_13961,N_13360,N_13139);
nor U13962 (N_13962,N_13366,N_13378);
nand U13963 (N_13963,N_13278,N_13368);
xnor U13964 (N_13964,N_13365,N_13067);
xnor U13965 (N_13965,N_13496,N_13224);
or U13966 (N_13966,N_13299,N_13362);
and U13967 (N_13967,N_13234,N_13128);
nand U13968 (N_13968,N_13078,N_13373);
nor U13969 (N_13969,N_13489,N_13251);
xor U13970 (N_13970,N_13123,N_13466);
xnor U13971 (N_13971,N_13076,N_13116);
and U13972 (N_13972,N_13186,N_13077);
nand U13973 (N_13973,N_13009,N_13417);
or U13974 (N_13974,N_13491,N_13054);
nor U13975 (N_13975,N_13036,N_13284);
nor U13976 (N_13976,N_13340,N_13151);
nor U13977 (N_13977,N_13057,N_13040);
nand U13978 (N_13978,N_13333,N_13331);
nand U13979 (N_13979,N_13335,N_13433);
and U13980 (N_13980,N_13211,N_13392);
nand U13981 (N_13981,N_13026,N_13041);
nor U13982 (N_13982,N_13121,N_13431);
or U13983 (N_13983,N_13411,N_13297);
xor U13984 (N_13984,N_13498,N_13318);
or U13985 (N_13985,N_13122,N_13084);
and U13986 (N_13986,N_13036,N_13341);
or U13987 (N_13987,N_13471,N_13154);
and U13988 (N_13988,N_13001,N_13349);
xor U13989 (N_13989,N_13235,N_13149);
and U13990 (N_13990,N_13488,N_13499);
or U13991 (N_13991,N_13355,N_13229);
and U13992 (N_13992,N_13204,N_13228);
nor U13993 (N_13993,N_13347,N_13115);
nand U13994 (N_13994,N_13423,N_13091);
or U13995 (N_13995,N_13128,N_13482);
nand U13996 (N_13996,N_13461,N_13033);
or U13997 (N_13997,N_13165,N_13140);
and U13998 (N_13998,N_13318,N_13402);
xnor U13999 (N_13999,N_13062,N_13488);
and U14000 (N_14000,N_13862,N_13563);
and U14001 (N_14001,N_13799,N_13820);
and U14002 (N_14002,N_13510,N_13802);
nand U14003 (N_14003,N_13516,N_13785);
or U14004 (N_14004,N_13595,N_13894);
xor U14005 (N_14005,N_13755,N_13776);
and U14006 (N_14006,N_13653,N_13693);
or U14007 (N_14007,N_13819,N_13959);
xor U14008 (N_14008,N_13854,N_13912);
nand U14009 (N_14009,N_13640,N_13853);
or U14010 (N_14010,N_13977,N_13788);
xnor U14011 (N_14011,N_13791,N_13800);
or U14012 (N_14012,N_13938,N_13848);
or U14013 (N_14013,N_13571,N_13649);
or U14014 (N_14014,N_13890,N_13674);
nor U14015 (N_14015,N_13750,N_13937);
xor U14016 (N_14016,N_13960,N_13614);
nand U14017 (N_14017,N_13515,N_13817);
nand U14018 (N_14018,N_13587,N_13527);
xnor U14019 (N_14019,N_13648,N_13541);
nand U14020 (N_14020,N_13883,N_13503);
nand U14021 (N_14021,N_13903,N_13831);
and U14022 (N_14022,N_13813,N_13897);
nand U14023 (N_14023,N_13578,N_13728);
and U14024 (N_14024,N_13920,N_13878);
xor U14025 (N_14025,N_13551,N_13832);
xor U14026 (N_14026,N_13689,N_13885);
nand U14027 (N_14027,N_13526,N_13955);
and U14028 (N_14028,N_13625,N_13962);
and U14029 (N_14029,N_13624,N_13569);
nand U14030 (N_14030,N_13988,N_13880);
and U14031 (N_14031,N_13583,N_13941);
nor U14032 (N_14032,N_13661,N_13901);
xor U14033 (N_14033,N_13596,N_13570);
and U14034 (N_14034,N_13914,N_13623);
xor U14035 (N_14035,N_13740,N_13687);
and U14036 (N_14036,N_13796,N_13658);
xnor U14037 (N_14037,N_13926,N_13836);
xor U14038 (N_14038,N_13999,N_13919);
and U14039 (N_14039,N_13681,N_13718);
nand U14040 (N_14040,N_13644,N_13576);
nand U14041 (N_14041,N_13877,N_13904);
nand U14042 (N_14042,N_13879,N_13922);
xor U14043 (N_14043,N_13605,N_13752);
nand U14044 (N_14044,N_13706,N_13828);
and U14045 (N_14045,N_13609,N_13851);
nor U14046 (N_14046,N_13533,N_13845);
nand U14047 (N_14047,N_13936,N_13532);
nor U14048 (N_14048,N_13767,N_13824);
nor U14049 (N_14049,N_13835,N_13995);
nand U14050 (N_14050,N_13873,N_13782);
xnor U14051 (N_14051,N_13968,N_13697);
nand U14052 (N_14052,N_13757,N_13775);
xnor U14053 (N_14053,N_13899,N_13666);
or U14054 (N_14054,N_13603,N_13792);
nand U14055 (N_14055,N_13822,N_13908);
nor U14056 (N_14056,N_13859,N_13809);
nand U14057 (N_14057,N_13652,N_13940);
nand U14058 (N_14058,N_13865,N_13615);
or U14059 (N_14059,N_13781,N_13794);
xnor U14060 (N_14060,N_13725,N_13893);
nand U14061 (N_14061,N_13748,N_13797);
nor U14062 (N_14062,N_13506,N_13784);
xnor U14063 (N_14063,N_13778,N_13590);
nand U14064 (N_14064,N_13699,N_13954);
and U14065 (N_14065,N_13655,N_13586);
nand U14066 (N_14066,N_13882,N_13841);
or U14067 (N_14067,N_13694,N_13867);
nor U14068 (N_14068,N_13852,N_13654);
and U14069 (N_14069,N_13742,N_13975);
xor U14070 (N_14070,N_13630,N_13762);
nand U14071 (N_14071,N_13734,N_13735);
or U14072 (N_14072,N_13948,N_13850);
nand U14073 (N_14073,N_13747,N_13700);
nand U14074 (N_14074,N_13584,N_13925);
and U14075 (N_14075,N_13801,N_13994);
and U14076 (N_14076,N_13513,N_13534);
or U14077 (N_14077,N_13956,N_13556);
nor U14078 (N_14078,N_13635,N_13896);
xnor U14079 (N_14079,N_13622,N_13714);
xor U14080 (N_14080,N_13965,N_13679);
or U14081 (N_14081,N_13509,N_13729);
xnor U14082 (N_14082,N_13918,N_13834);
or U14083 (N_14083,N_13567,N_13540);
xor U14084 (N_14084,N_13838,N_13807);
xor U14085 (N_14085,N_13548,N_13927);
nor U14086 (N_14086,N_13844,N_13521);
nor U14087 (N_14087,N_13617,N_13727);
nor U14088 (N_14088,N_13857,N_13537);
xnor U14089 (N_14089,N_13935,N_13958);
and U14090 (N_14090,N_13731,N_13830);
nor U14091 (N_14091,N_13637,N_13629);
nand U14092 (N_14092,N_13712,N_13864);
or U14093 (N_14093,N_13721,N_13564);
and U14094 (N_14094,N_13626,N_13581);
nand U14095 (N_14095,N_13573,N_13677);
nor U14096 (N_14096,N_13680,N_13608);
or U14097 (N_14097,N_13501,N_13702);
nor U14098 (N_14098,N_13546,N_13972);
nor U14099 (N_14099,N_13708,N_13872);
or U14100 (N_14100,N_13783,N_13547);
xor U14101 (N_14101,N_13979,N_13722);
xor U14102 (N_14102,N_13633,N_13726);
nor U14103 (N_14103,N_13870,N_13868);
nand U14104 (N_14104,N_13939,N_13577);
nand U14105 (N_14105,N_13826,N_13924);
xor U14106 (N_14106,N_13860,N_13987);
nor U14107 (N_14107,N_13508,N_13618);
nor U14108 (N_14108,N_13665,N_13847);
xor U14109 (N_14109,N_13930,N_13507);
or U14110 (N_14110,N_13662,N_13871);
and U14111 (N_14111,N_13818,N_13620);
or U14112 (N_14112,N_13953,N_13610);
xor U14113 (N_14113,N_13759,N_13989);
xor U14114 (N_14114,N_13973,N_13898);
or U14115 (N_14115,N_13594,N_13602);
or U14116 (N_14116,N_13886,N_13566);
xor U14117 (N_14117,N_13932,N_13803);
nand U14118 (N_14118,N_13579,N_13568);
or U14119 (N_14119,N_13642,N_13631);
nand U14120 (N_14120,N_13634,N_13984);
and U14121 (N_14121,N_13849,N_13518);
or U14122 (N_14122,N_13723,N_13942);
and U14123 (N_14123,N_13833,N_13787);
and U14124 (N_14124,N_13963,N_13686);
or U14125 (N_14125,N_13713,N_13676);
xor U14126 (N_14126,N_13692,N_13542);
nand U14127 (N_14127,N_13780,N_13671);
or U14128 (N_14128,N_13812,N_13810);
xor U14129 (N_14129,N_13601,N_13668);
nand U14130 (N_14130,N_13717,N_13691);
and U14131 (N_14131,N_13651,N_13743);
or U14132 (N_14132,N_13970,N_13528);
nand U14133 (N_14133,N_13753,N_13768);
xor U14134 (N_14134,N_13565,N_13656);
nand U14135 (N_14135,N_13522,N_13805);
nor U14136 (N_14136,N_13888,N_13544);
or U14137 (N_14137,N_13967,N_13500);
nand U14138 (N_14138,N_13682,N_13843);
and U14139 (N_14139,N_13980,N_13646);
and U14140 (N_14140,N_13761,N_13993);
xnor U14141 (N_14141,N_13598,N_13763);
nand U14142 (N_14142,N_13530,N_13588);
or U14143 (N_14143,N_13952,N_13957);
nand U14144 (N_14144,N_13892,N_13823);
xnor U14145 (N_14145,N_13517,N_13933);
nand U14146 (N_14146,N_13664,N_13730);
xor U14147 (N_14147,N_13554,N_13552);
and U14148 (N_14148,N_13982,N_13811);
xnor U14149 (N_14149,N_13923,N_13690);
nand U14150 (N_14150,N_13675,N_13525);
nor U14151 (N_14151,N_13943,N_13964);
nor U14152 (N_14152,N_13876,N_13770);
or U14153 (N_14153,N_13793,N_13944);
or U14154 (N_14154,N_13531,N_13769);
xor U14155 (N_14155,N_13790,N_13705);
or U14156 (N_14156,N_13669,N_13683);
or U14157 (N_14157,N_13560,N_13981);
nor U14158 (N_14158,N_13504,N_13561);
or U14159 (N_14159,N_13558,N_13580);
or U14160 (N_14160,N_13754,N_13815);
or U14161 (N_14161,N_13766,N_13641);
or U14162 (N_14162,N_13737,N_13703);
xor U14163 (N_14163,N_13756,N_13639);
or U14164 (N_14164,N_13945,N_13921);
xnor U14165 (N_14165,N_13619,N_13971);
xnor U14166 (N_14166,N_13808,N_13745);
and U14167 (N_14167,N_13946,N_13643);
xor U14168 (N_14168,N_13719,N_13621);
and U14169 (N_14169,N_13758,N_13696);
nor U14170 (N_14170,N_13869,N_13931);
xor U14171 (N_14171,N_13724,N_13774);
and U14172 (N_14172,N_13986,N_13861);
xnor U14173 (N_14173,N_13647,N_13825);
and U14174 (N_14174,N_13779,N_13934);
or U14175 (N_14175,N_13738,N_13974);
or U14176 (N_14176,N_13559,N_13816);
nand U14177 (N_14177,N_13983,N_13604);
nor U14178 (N_14178,N_13961,N_13523);
or U14179 (N_14179,N_13519,N_13947);
or U14180 (N_14180,N_13910,N_13667);
and U14181 (N_14181,N_13911,N_13613);
nor U14182 (N_14182,N_13884,N_13688);
nor U14183 (N_14183,N_13746,N_13916);
nor U14184 (N_14184,N_13711,N_13628);
nor U14185 (N_14185,N_13996,N_13990);
nand U14186 (N_14186,N_13827,N_13804);
and U14187 (N_14187,N_13949,N_13582);
xor U14188 (N_14188,N_13593,N_13659);
nor U14189 (N_14189,N_13660,N_13611);
nand U14190 (N_14190,N_13814,N_13606);
xnor U14191 (N_14191,N_13928,N_13716);
nand U14192 (N_14192,N_13550,N_13795);
nor U14193 (N_14193,N_13751,N_13915);
or U14194 (N_14194,N_13891,N_13585);
xor U14195 (N_14195,N_13562,N_13512);
nor U14196 (N_14196,N_13900,N_13998);
nor U14197 (N_14197,N_13502,N_13991);
and U14198 (N_14198,N_13597,N_13524);
xnor U14199 (N_14199,N_13645,N_13997);
xnor U14200 (N_14200,N_13543,N_13553);
xor U14201 (N_14201,N_13839,N_13895);
nor U14202 (N_14202,N_13917,N_13875);
or U14203 (N_14203,N_13650,N_13535);
nand U14204 (N_14204,N_13858,N_13720);
nor U14205 (N_14205,N_13978,N_13549);
or U14206 (N_14206,N_13575,N_13985);
xor U14207 (N_14207,N_13663,N_13874);
nand U14208 (N_14208,N_13673,N_13710);
and U14209 (N_14209,N_13771,N_13657);
and U14210 (N_14210,N_13749,N_13889);
or U14211 (N_14211,N_13966,N_13684);
nor U14212 (N_14212,N_13765,N_13976);
nand U14213 (N_14213,N_13505,N_13760);
nand U14214 (N_14214,N_13600,N_13842);
and U14215 (N_14215,N_13950,N_13913);
nand U14216 (N_14216,N_13545,N_13638);
nor U14217 (N_14217,N_13627,N_13591);
nand U14218 (N_14218,N_13672,N_13741);
nand U14219 (N_14219,N_13529,N_13520);
nor U14220 (N_14220,N_13715,N_13840);
xor U14221 (N_14221,N_13732,N_13589);
nor U14222 (N_14222,N_13821,N_13555);
xor U14223 (N_14223,N_13902,N_13907);
or U14224 (N_14224,N_13773,N_13698);
nand U14225 (N_14225,N_13881,N_13969);
nor U14226 (N_14226,N_13670,N_13744);
xnor U14227 (N_14227,N_13736,N_13786);
xnor U14228 (N_14228,N_13704,N_13829);
and U14229 (N_14229,N_13607,N_13887);
xor U14230 (N_14230,N_13538,N_13777);
or U14231 (N_14231,N_13539,N_13709);
or U14232 (N_14232,N_13536,N_13557);
nor U14233 (N_14233,N_13511,N_13798);
nor U14234 (N_14234,N_13856,N_13906);
nor U14235 (N_14235,N_13592,N_13806);
xnor U14236 (N_14236,N_13764,N_13863);
nand U14237 (N_14237,N_13739,N_13632);
and U14238 (N_14238,N_13929,N_13572);
nand U14239 (N_14239,N_13514,N_13616);
nand U14240 (N_14240,N_13574,N_13695);
nand U14241 (N_14241,N_13789,N_13701);
and U14242 (N_14242,N_13707,N_13678);
nor U14243 (N_14243,N_13846,N_13837);
or U14244 (N_14244,N_13992,N_13599);
or U14245 (N_14245,N_13772,N_13612);
nand U14246 (N_14246,N_13636,N_13905);
nand U14247 (N_14247,N_13951,N_13733);
nor U14248 (N_14248,N_13909,N_13866);
xor U14249 (N_14249,N_13685,N_13855);
or U14250 (N_14250,N_13577,N_13594);
or U14251 (N_14251,N_13675,N_13631);
nor U14252 (N_14252,N_13509,N_13698);
nor U14253 (N_14253,N_13875,N_13989);
or U14254 (N_14254,N_13844,N_13773);
nand U14255 (N_14255,N_13799,N_13643);
nor U14256 (N_14256,N_13624,N_13613);
nand U14257 (N_14257,N_13800,N_13914);
or U14258 (N_14258,N_13938,N_13534);
nor U14259 (N_14259,N_13907,N_13812);
or U14260 (N_14260,N_13767,N_13686);
nor U14261 (N_14261,N_13758,N_13716);
nor U14262 (N_14262,N_13868,N_13613);
nand U14263 (N_14263,N_13978,N_13961);
and U14264 (N_14264,N_13609,N_13604);
nor U14265 (N_14265,N_13872,N_13512);
and U14266 (N_14266,N_13953,N_13898);
and U14267 (N_14267,N_13635,N_13786);
and U14268 (N_14268,N_13546,N_13908);
nor U14269 (N_14269,N_13923,N_13844);
and U14270 (N_14270,N_13561,N_13666);
xor U14271 (N_14271,N_13875,N_13707);
or U14272 (N_14272,N_13639,N_13540);
nor U14273 (N_14273,N_13677,N_13674);
nand U14274 (N_14274,N_13723,N_13820);
or U14275 (N_14275,N_13878,N_13951);
xor U14276 (N_14276,N_13660,N_13618);
or U14277 (N_14277,N_13577,N_13507);
and U14278 (N_14278,N_13505,N_13519);
or U14279 (N_14279,N_13848,N_13763);
nand U14280 (N_14280,N_13876,N_13582);
and U14281 (N_14281,N_13661,N_13876);
and U14282 (N_14282,N_13916,N_13651);
xor U14283 (N_14283,N_13913,N_13842);
and U14284 (N_14284,N_13615,N_13799);
or U14285 (N_14285,N_13752,N_13809);
and U14286 (N_14286,N_13717,N_13619);
nor U14287 (N_14287,N_13672,N_13810);
nand U14288 (N_14288,N_13794,N_13659);
and U14289 (N_14289,N_13789,N_13743);
and U14290 (N_14290,N_13934,N_13860);
nor U14291 (N_14291,N_13827,N_13877);
xnor U14292 (N_14292,N_13706,N_13987);
or U14293 (N_14293,N_13886,N_13884);
nand U14294 (N_14294,N_13784,N_13914);
xnor U14295 (N_14295,N_13767,N_13957);
or U14296 (N_14296,N_13966,N_13658);
and U14297 (N_14297,N_13867,N_13774);
xor U14298 (N_14298,N_13537,N_13860);
or U14299 (N_14299,N_13811,N_13517);
or U14300 (N_14300,N_13592,N_13624);
nand U14301 (N_14301,N_13653,N_13968);
xnor U14302 (N_14302,N_13633,N_13632);
nor U14303 (N_14303,N_13968,N_13798);
xor U14304 (N_14304,N_13794,N_13804);
nand U14305 (N_14305,N_13808,N_13716);
or U14306 (N_14306,N_13669,N_13648);
nor U14307 (N_14307,N_13534,N_13525);
and U14308 (N_14308,N_13791,N_13515);
nand U14309 (N_14309,N_13728,N_13773);
and U14310 (N_14310,N_13561,N_13586);
nand U14311 (N_14311,N_13976,N_13925);
and U14312 (N_14312,N_13922,N_13604);
and U14313 (N_14313,N_13708,N_13761);
xor U14314 (N_14314,N_13938,N_13897);
nor U14315 (N_14315,N_13700,N_13535);
or U14316 (N_14316,N_13871,N_13511);
nor U14317 (N_14317,N_13977,N_13557);
xor U14318 (N_14318,N_13847,N_13555);
xnor U14319 (N_14319,N_13722,N_13532);
xnor U14320 (N_14320,N_13763,N_13833);
nor U14321 (N_14321,N_13529,N_13936);
nor U14322 (N_14322,N_13809,N_13668);
nand U14323 (N_14323,N_13891,N_13858);
or U14324 (N_14324,N_13599,N_13807);
nand U14325 (N_14325,N_13773,N_13678);
or U14326 (N_14326,N_13598,N_13907);
nor U14327 (N_14327,N_13513,N_13797);
nor U14328 (N_14328,N_13895,N_13716);
and U14329 (N_14329,N_13975,N_13602);
nand U14330 (N_14330,N_13543,N_13687);
nor U14331 (N_14331,N_13738,N_13935);
xnor U14332 (N_14332,N_13539,N_13525);
and U14333 (N_14333,N_13529,N_13663);
nor U14334 (N_14334,N_13841,N_13786);
nor U14335 (N_14335,N_13718,N_13868);
and U14336 (N_14336,N_13723,N_13694);
or U14337 (N_14337,N_13940,N_13527);
nor U14338 (N_14338,N_13791,N_13631);
and U14339 (N_14339,N_13818,N_13898);
nor U14340 (N_14340,N_13550,N_13629);
or U14341 (N_14341,N_13755,N_13500);
and U14342 (N_14342,N_13630,N_13561);
xnor U14343 (N_14343,N_13590,N_13900);
nor U14344 (N_14344,N_13763,N_13750);
nor U14345 (N_14345,N_13522,N_13734);
xnor U14346 (N_14346,N_13868,N_13618);
and U14347 (N_14347,N_13792,N_13689);
xor U14348 (N_14348,N_13982,N_13564);
or U14349 (N_14349,N_13634,N_13501);
and U14350 (N_14350,N_13718,N_13980);
nand U14351 (N_14351,N_13823,N_13822);
nand U14352 (N_14352,N_13643,N_13678);
nand U14353 (N_14353,N_13721,N_13792);
xor U14354 (N_14354,N_13781,N_13532);
nor U14355 (N_14355,N_13904,N_13538);
or U14356 (N_14356,N_13797,N_13876);
and U14357 (N_14357,N_13933,N_13502);
or U14358 (N_14358,N_13683,N_13923);
and U14359 (N_14359,N_13783,N_13916);
and U14360 (N_14360,N_13601,N_13795);
xnor U14361 (N_14361,N_13523,N_13805);
and U14362 (N_14362,N_13817,N_13673);
or U14363 (N_14363,N_13881,N_13660);
xnor U14364 (N_14364,N_13710,N_13669);
or U14365 (N_14365,N_13825,N_13589);
xor U14366 (N_14366,N_13858,N_13745);
nand U14367 (N_14367,N_13757,N_13565);
and U14368 (N_14368,N_13595,N_13775);
nor U14369 (N_14369,N_13546,N_13758);
nor U14370 (N_14370,N_13899,N_13940);
nor U14371 (N_14371,N_13870,N_13596);
xnor U14372 (N_14372,N_13948,N_13720);
and U14373 (N_14373,N_13921,N_13733);
or U14374 (N_14374,N_13510,N_13705);
or U14375 (N_14375,N_13741,N_13542);
and U14376 (N_14376,N_13998,N_13801);
and U14377 (N_14377,N_13611,N_13887);
nor U14378 (N_14378,N_13533,N_13994);
xor U14379 (N_14379,N_13683,N_13799);
or U14380 (N_14380,N_13933,N_13794);
and U14381 (N_14381,N_13758,N_13558);
nand U14382 (N_14382,N_13685,N_13712);
nor U14383 (N_14383,N_13785,N_13804);
and U14384 (N_14384,N_13814,N_13561);
or U14385 (N_14385,N_13738,N_13529);
nor U14386 (N_14386,N_13589,N_13872);
or U14387 (N_14387,N_13798,N_13549);
xor U14388 (N_14388,N_13964,N_13527);
nand U14389 (N_14389,N_13647,N_13634);
and U14390 (N_14390,N_13994,N_13944);
nor U14391 (N_14391,N_13565,N_13704);
xnor U14392 (N_14392,N_13753,N_13611);
nand U14393 (N_14393,N_13858,N_13771);
or U14394 (N_14394,N_13536,N_13605);
nand U14395 (N_14395,N_13667,N_13877);
or U14396 (N_14396,N_13688,N_13652);
xor U14397 (N_14397,N_13509,N_13789);
or U14398 (N_14398,N_13838,N_13893);
nand U14399 (N_14399,N_13691,N_13896);
xor U14400 (N_14400,N_13582,N_13748);
nand U14401 (N_14401,N_13523,N_13615);
nand U14402 (N_14402,N_13950,N_13572);
and U14403 (N_14403,N_13734,N_13585);
and U14404 (N_14404,N_13835,N_13623);
or U14405 (N_14405,N_13596,N_13647);
or U14406 (N_14406,N_13566,N_13601);
and U14407 (N_14407,N_13765,N_13505);
nor U14408 (N_14408,N_13814,N_13709);
nand U14409 (N_14409,N_13760,N_13551);
and U14410 (N_14410,N_13628,N_13606);
or U14411 (N_14411,N_13729,N_13748);
xor U14412 (N_14412,N_13702,N_13886);
and U14413 (N_14413,N_13757,N_13672);
xnor U14414 (N_14414,N_13669,N_13976);
and U14415 (N_14415,N_13994,N_13983);
and U14416 (N_14416,N_13816,N_13934);
or U14417 (N_14417,N_13733,N_13762);
or U14418 (N_14418,N_13647,N_13627);
and U14419 (N_14419,N_13924,N_13677);
nor U14420 (N_14420,N_13574,N_13652);
nand U14421 (N_14421,N_13987,N_13945);
and U14422 (N_14422,N_13780,N_13693);
nor U14423 (N_14423,N_13915,N_13708);
nand U14424 (N_14424,N_13581,N_13718);
and U14425 (N_14425,N_13881,N_13970);
nand U14426 (N_14426,N_13561,N_13663);
xor U14427 (N_14427,N_13905,N_13608);
and U14428 (N_14428,N_13813,N_13682);
and U14429 (N_14429,N_13682,N_13998);
nand U14430 (N_14430,N_13516,N_13932);
xor U14431 (N_14431,N_13958,N_13704);
and U14432 (N_14432,N_13631,N_13709);
nor U14433 (N_14433,N_13591,N_13694);
nor U14434 (N_14434,N_13734,N_13877);
nand U14435 (N_14435,N_13664,N_13683);
nand U14436 (N_14436,N_13709,N_13590);
and U14437 (N_14437,N_13783,N_13674);
or U14438 (N_14438,N_13536,N_13645);
xor U14439 (N_14439,N_13674,N_13635);
or U14440 (N_14440,N_13893,N_13629);
nor U14441 (N_14441,N_13904,N_13520);
nor U14442 (N_14442,N_13577,N_13931);
nor U14443 (N_14443,N_13622,N_13875);
nand U14444 (N_14444,N_13780,N_13942);
nor U14445 (N_14445,N_13652,N_13525);
nand U14446 (N_14446,N_13802,N_13631);
xnor U14447 (N_14447,N_13513,N_13641);
and U14448 (N_14448,N_13745,N_13682);
nand U14449 (N_14449,N_13554,N_13559);
or U14450 (N_14450,N_13775,N_13696);
xor U14451 (N_14451,N_13504,N_13930);
nor U14452 (N_14452,N_13864,N_13778);
and U14453 (N_14453,N_13988,N_13866);
nor U14454 (N_14454,N_13715,N_13568);
and U14455 (N_14455,N_13622,N_13769);
nand U14456 (N_14456,N_13799,N_13551);
or U14457 (N_14457,N_13844,N_13872);
or U14458 (N_14458,N_13737,N_13546);
nand U14459 (N_14459,N_13633,N_13536);
xor U14460 (N_14460,N_13563,N_13752);
and U14461 (N_14461,N_13574,N_13694);
nor U14462 (N_14462,N_13654,N_13863);
nor U14463 (N_14463,N_13646,N_13985);
nand U14464 (N_14464,N_13875,N_13756);
nor U14465 (N_14465,N_13613,N_13536);
xnor U14466 (N_14466,N_13619,N_13691);
and U14467 (N_14467,N_13627,N_13989);
and U14468 (N_14468,N_13954,N_13786);
xor U14469 (N_14469,N_13841,N_13967);
or U14470 (N_14470,N_13812,N_13512);
or U14471 (N_14471,N_13765,N_13815);
xor U14472 (N_14472,N_13696,N_13648);
and U14473 (N_14473,N_13925,N_13947);
xor U14474 (N_14474,N_13699,N_13575);
xor U14475 (N_14475,N_13673,N_13611);
xor U14476 (N_14476,N_13935,N_13941);
nand U14477 (N_14477,N_13775,N_13814);
and U14478 (N_14478,N_13501,N_13572);
nand U14479 (N_14479,N_13748,N_13640);
xor U14480 (N_14480,N_13571,N_13710);
xnor U14481 (N_14481,N_13930,N_13501);
nand U14482 (N_14482,N_13594,N_13980);
xnor U14483 (N_14483,N_13814,N_13958);
nand U14484 (N_14484,N_13863,N_13650);
nor U14485 (N_14485,N_13863,N_13810);
and U14486 (N_14486,N_13544,N_13671);
nor U14487 (N_14487,N_13584,N_13856);
or U14488 (N_14488,N_13969,N_13973);
and U14489 (N_14489,N_13559,N_13648);
and U14490 (N_14490,N_13878,N_13534);
nand U14491 (N_14491,N_13823,N_13596);
and U14492 (N_14492,N_13729,N_13871);
or U14493 (N_14493,N_13951,N_13518);
nand U14494 (N_14494,N_13528,N_13586);
and U14495 (N_14495,N_13892,N_13652);
nand U14496 (N_14496,N_13946,N_13813);
nor U14497 (N_14497,N_13739,N_13919);
nor U14498 (N_14498,N_13969,N_13924);
and U14499 (N_14499,N_13686,N_13612);
or U14500 (N_14500,N_14249,N_14329);
nand U14501 (N_14501,N_14208,N_14492);
nor U14502 (N_14502,N_14290,N_14189);
nand U14503 (N_14503,N_14141,N_14424);
nor U14504 (N_14504,N_14077,N_14096);
nor U14505 (N_14505,N_14379,N_14456);
nand U14506 (N_14506,N_14025,N_14322);
and U14507 (N_14507,N_14114,N_14495);
and U14508 (N_14508,N_14388,N_14132);
xnor U14509 (N_14509,N_14272,N_14421);
or U14510 (N_14510,N_14371,N_14123);
nand U14511 (N_14511,N_14247,N_14246);
or U14512 (N_14512,N_14367,N_14281);
xor U14513 (N_14513,N_14201,N_14185);
nand U14514 (N_14514,N_14490,N_14211);
or U14515 (N_14515,N_14050,N_14494);
and U14516 (N_14516,N_14214,N_14269);
xor U14517 (N_14517,N_14469,N_14468);
nor U14518 (N_14518,N_14307,N_14274);
and U14519 (N_14519,N_14463,N_14280);
nand U14520 (N_14520,N_14145,N_14216);
nand U14521 (N_14521,N_14110,N_14333);
or U14522 (N_14522,N_14075,N_14170);
nand U14523 (N_14523,N_14295,N_14239);
and U14524 (N_14524,N_14093,N_14372);
xnor U14525 (N_14525,N_14302,N_14262);
nand U14526 (N_14526,N_14352,N_14271);
nand U14527 (N_14527,N_14163,N_14351);
nor U14528 (N_14528,N_14341,N_14160);
nand U14529 (N_14529,N_14104,N_14432);
and U14530 (N_14530,N_14192,N_14013);
xor U14531 (N_14531,N_14085,N_14207);
xnor U14532 (N_14532,N_14080,N_14314);
or U14533 (N_14533,N_14245,N_14299);
xnor U14534 (N_14534,N_14435,N_14476);
nand U14535 (N_14535,N_14078,N_14058);
nor U14536 (N_14536,N_14174,N_14015);
xor U14537 (N_14537,N_14045,N_14386);
nor U14538 (N_14538,N_14230,N_14312);
nand U14539 (N_14539,N_14173,N_14217);
or U14540 (N_14540,N_14266,N_14231);
xor U14541 (N_14541,N_14179,N_14199);
and U14542 (N_14542,N_14429,N_14076);
or U14543 (N_14543,N_14128,N_14489);
nor U14544 (N_14544,N_14483,N_14094);
and U14545 (N_14545,N_14018,N_14493);
xnor U14546 (N_14546,N_14115,N_14464);
nand U14547 (N_14547,N_14142,N_14182);
and U14548 (N_14548,N_14426,N_14089);
nor U14549 (N_14549,N_14027,N_14291);
xnor U14550 (N_14550,N_14487,N_14203);
or U14551 (N_14551,N_14153,N_14046);
nor U14552 (N_14552,N_14233,N_14324);
xnor U14553 (N_14553,N_14028,N_14311);
or U14554 (N_14554,N_14382,N_14306);
or U14555 (N_14555,N_14073,N_14397);
nand U14556 (N_14556,N_14229,N_14437);
nor U14557 (N_14557,N_14002,N_14418);
or U14558 (N_14558,N_14219,N_14393);
and U14559 (N_14559,N_14167,N_14036);
nand U14560 (N_14560,N_14331,N_14238);
or U14561 (N_14561,N_14254,N_14431);
xor U14562 (N_14562,N_14130,N_14406);
and U14563 (N_14563,N_14419,N_14082);
xor U14564 (N_14564,N_14156,N_14353);
nand U14565 (N_14565,N_14024,N_14081);
or U14566 (N_14566,N_14034,N_14155);
nor U14567 (N_14567,N_14359,N_14164);
and U14568 (N_14568,N_14042,N_14067);
xnor U14569 (N_14569,N_14317,N_14086);
or U14570 (N_14570,N_14008,N_14327);
nor U14571 (N_14571,N_14244,N_14480);
xnor U14572 (N_14572,N_14062,N_14477);
xnor U14573 (N_14573,N_14442,N_14482);
and U14574 (N_14574,N_14151,N_14136);
and U14575 (N_14575,N_14071,N_14068);
and U14576 (N_14576,N_14248,N_14412);
nand U14577 (N_14577,N_14445,N_14157);
nand U14578 (N_14578,N_14041,N_14378);
or U14579 (N_14579,N_14006,N_14448);
and U14580 (N_14580,N_14055,N_14091);
xor U14581 (N_14581,N_14095,N_14320);
xnor U14582 (N_14582,N_14010,N_14111);
and U14583 (N_14583,N_14102,N_14121);
or U14584 (N_14584,N_14323,N_14187);
nand U14585 (N_14585,N_14099,N_14223);
nand U14586 (N_14586,N_14385,N_14415);
and U14587 (N_14587,N_14275,N_14049);
and U14588 (N_14588,N_14172,N_14326);
nand U14589 (N_14589,N_14033,N_14175);
and U14590 (N_14590,N_14113,N_14001);
xnor U14591 (N_14591,N_14263,N_14410);
or U14592 (N_14592,N_14440,N_14334);
nand U14593 (N_14593,N_14000,N_14321);
or U14594 (N_14594,N_14169,N_14070);
xnor U14595 (N_14595,N_14003,N_14053);
xnor U14596 (N_14596,N_14105,N_14304);
and U14597 (N_14597,N_14190,N_14020);
nor U14598 (N_14598,N_14029,N_14162);
xor U14599 (N_14599,N_14079,N_14258);
nor U14600 (N_14600,N_14237,N_14444);
xor U14601 (N_14601,N_14069,N_14335);
or U14602 (N_14602,N_14138,N_14087);
and U14603 (N_14603,N_14318,N_14012);
nand U14604 (N_14604,N_14210,N_14150);
nand U14605 (N_14605,N_14471,N_14196);
and U14606 (N_14606,N_14491,N_14235);
nand U14607 (N_14607,N_14261,N_14109);
and U14608 (N_14608,N_14241,N_14116);
or U14609 (N_14609,N_14218,N_14016);
or U14610 (N_14610,N_14328,N_14242);
and U14611 (N_14611,N_14101,N_14198);
xnor U14612 (N_14612,N_14369,N_14428);
nor U14613 (N_14613,N_14017,N_14420);
nor U14614 (N_14614,N_14325,N_14066);
and U14615 (N_14615,N_14363,N_14383);
xnor U14616 (N_14616,N_14287,N_14195);
nand U14617 (N_14617,N_14227,N_14273);
xnor U14618 (N_14618,N_14349,N_14143);
and U14619 (N_14619,N_14253,N_14106);
xor U14620 (N_14620,N_14061,N_14060);
and U14621 (N_14621,N_14394,N_14090);
nor U14622 (N_14622,N_14498,N_14459);
nor U14623 (N_14623,N_14232,N_14485);
nand U14624 (N_14624,N_14004,N_14140);
nand U14625 (N_14625,N_14414,N_14276);
or U14626 (N_14626,N_14470,N_14316);
nor U14627 (N_14627,N_14204,N_14344);
xnor U14628 (N_14628,N_14159,N_14206);
nor U14629 (N_14629,N_14286,N_14403);
nor U14630 (N_14630,N_14446,N_14148);
nand U14631 (N_14631,N_14310,N_14122);
and U14632 (N_14632,N_14417,N_14222);
nand U14633 (N_14633,N_14413,N_14057);
nor U14634 (N_14634,N_14032,N_14339);
and U14635 (N_14635,N_14184,N_14396);
or U14636 (N_14636,N_14166,N_14390);
xor U14637 (N_14637,N_14308,N_14348);
nor U14638 (N_14638,N_14380,N_14243);
or U14639 (N_14639,N_14496,N_14289);
or U14640 (N_14640,N_14288,N_14059);
or U14641 (N_14641,N_14112,N_14197);
or U14642 (N_14642,N_14457,N_14285);
nand U14643 (N_14643,N_14319,N_14191);
nor U14644 (N_14644,N_14064,N_14236);
xnor U14645 (N_14645,N_14047,N_14309);
nor U14646 (N_14646,N_14220,N_14336);
xor U14647 (N_14647,N_14117,N_14165);
nand U14648 (N_14648,N_14452,N_14405);
or U14649 (N_14649,N_14072,N_14212);
nand U14650 (N_14650,N_14467,N_14293);
nor U14651 (N_14651,N_14375,N_14434);
xnor U14652 (N_14652,N_14268,N_14134);
and U14653 (N_14653,N_14011,N_14465);
and U14654 (N_14654,N_14144,N_14346);
and U14655 (N_14655,N_14399,N_14119);
and U14656 (N_14656,N_14332,N_14455);
or U14657 (N_14657,N_14256,N_14007);
or U14658 (N_14658,N_14026,N_14226);
nor U14659 (N_14659,N_14120,N_14458);
nor U14660 (N_14660,N_14466,N_14284);
nand U14661 (N_14661,N_14225,N_14313);
nor U14662 (N_14662,N_14146,N_14347);
xor U14663 (N_14663,N_14330,N_14499);
or U14664 (N_14664,N_14384,N_14368);
nand U14665 (N_14665,N_14441,N_14478);
nand U14666 (N_14666,N_14400,N_14181);
xnor U14667 (N_14667,N_14152,N_14462);
and U14668 (N_14668,N_14063,N_14065);
or U14669 (N_14669,N_14209,N_14021);
or U14670 (N_14670,N_14088,N_14161);
xnor U14671 (N_14671,N_14479,N_14257);
and U14672 (N_14672,N_14297,N_14205);
or U14673 (N_14673,N_14133,N_14449);
and U14674 (N_14674,N_14411,N_14279);
nor U14675 (N_14675,N_14461,N_14433);
or U14676 (N_14676,N_14083,N_14048);
nand U14677 (N_14677,N_14345,N_14124);
xnor U14678 (N_14678,N_14194,N_14350);
and U14679 (N_14679,N_14259,N_14129);
nor U14680 (N_14680,N_14391,N_14366);
or U14681 (N_14681,N_14044,N_14147);
nor U14682 (N_14682,N_14168,N_14381);
nand U14683 (N_14683,N_14423,N_14377);
and U14684 (N_14684,N_14402,N_14030);
xor U14685 (N_14685,N_14283,N_14355);
and U14686 (N_14686,N_14474,N_14100);
nor U14687 (N_14687,N_14398,N_14358);
xor U14688 (N_14688,N_14250,N_14387);
nor U14689 (N_14689,N_14131,N_14292);
nor U14690 (N_14690,N_14450,N_14425);
xnor U14691 (N_14691,N_14342,N_14186);
xnor U14692 (N_14692,N_14270,N_14180);
and U14693 (N_14693,N_14107,N_14497);
xnor U14694 (N_14694,N_14486,N_14296);
and U14695 (N_14695,N_14454,N_14023);
xor U14696 (N_14696,N_14427,N_14364);
nor U14697 (N_14697,N_14188,N_14215);
or U14698 (N_14698,N_14337,N_14056);
nor U14699 (N_14699,N_14038,N_14370);
nor U14700 (N_14700,N_14357,N_14224);
xor U14701 (N_14701,N_14202,N_14484);
or U14702 (N_14702,N_14255,N_14139);
and U14703 (N_14703,N_14338,N_14177);
nor U14704 (N_14704,N_14301,N_14416);
nor U14705 (N_14705,N_14014,N_14360);
and U14706 (N_14706,N_14473,N_14395);
nand U14707 (N_14707,N_14092,N_14221);
and U14708 (N_14708,N_14374,N_14125);
or U14709 (N_14709,N_14376,N_14213);
nor U14710 (N_14710,N_14481,N_14252);
xnor U14711 (N_14711,N_14365,N_14264);
xor U14712 (N_14712,N_14267,N_14392);
nor U14713 (N_14713,N_14265,N_14356);
and U14714 (N_14714,N_14282,N_14054);
xnor U14715 (N_14715,N_14475,N_14171);
xnor U14716 (N_14716,N_14251,N_14149);
or U14717 (N_14717,N_14040,N_14343);
and U14718 (N_14718,N_14009,N_14409);
or U14719 (N_14719,N_14298,N_14361);
xor U14720 (N_14720,N_14039,N_14200);
nand U14721 (N_14721,N_14260,N_14303);
and U14722 (N_14722,N_14315,N_14362);
or U14723 (N_14723,N_14404,N_14037);
nor U14724 (N_14724,N_14408,N_14447);
or U14725 (N_14725,N_14234,N_14472);
nand U14726 (N_14726,N_14135,N_14460);
nand U14727 (N_14727,N_14240,N_14407);
xnor U14728 (N_14728,N_14074,N_14005);
nor U14729 (N_14729,N_14118,N_14294);
nand U14730 (N_14730,N_14278,N_14439);
and U14731 (N_14731,N_14035,N_14401);
and U14732 (N_14732,N_14178,N_14019);
xnor U14733 (N_14733,N_14488,N_14022);
and U14734 (N_14734,N_14228,N_14422);
nor U14735 (N_14735,N_14137,N_14158);
and U14736 (N_14736,N_14103,N_14451);
or U14737 (N_14737,N_14436,N_14127);
xor U14738 (N_14738,N_14051,N_14154);
nand U14739 (N_14739,N_14389,N_14098);
nand U14740 (N_14740,N_14305,N_14043);
nand U14741 (N_14741,N_14340,N_14300);
and U14742 (N_14742,N_14438,N_14430);
nand U14743 (N_14743,N_14443,N_14031);
nor U14744 (N_14744,N_14193,N_14097);
nand U14745 (N_14745,N_14126,N_14453);
or U14746 (N_14746,N_14354,N_14176);
and U14747 (N_14747,N_14052,N_14183);
or U14748 (N_14748,N_14373,N_14084);
and U14749 (N_14749,N_14277,N_14108);
nor U14750 (N_14750,N_14123,N_14093);
nand U14751 (N_14751,N_14343,N_14138);
or U14752 (N_14752,N_14293,N_14229);
nor U14753 (N_14753,N_14207,N_14080);
xnor U14754 (N_14754,N_14467,N_14080);
nor U14755 (N_14755,N_14298,N_14145);
xnor U14756 (N_14756,N_14132,N_14264);
nor U14757 (N_14757,N_14250,N_14389);
xnor U14758 (N_14758,N_14032,N_14409);
xor U14759 (N_14759,N_14437,N_14382);
and U14760 (N_14760,N_14350,N_14362);
nand U14761 (N_14761,N_14264,N_14084);
nand U14762 (N_14762,N_14032,N_14053);
xor U14763 (N_14763,N_14342,N_14485);
nor U14764 (N_14764,N_14020,N_14006);
nand U14765 (N_14765,N_14272,N_14063);
or U14766 (N_14766,N_14325,N_14045);
or U14767 (N_14767,N_14273,N_14485);
or U14768 (N_14768,N_14126,N_14270);
xor U14769 (N_14769,N_14239,N_14113);
or U14770 (N_14770,N_14053,N_14041);
and U14771 (N_14771,N_14307,N_14026);
xor U14772 (N_14772,N_14394,N_14224);
nor U14773 (N_14773,N_14320,N_14170);
nor U14774 (N_14774,N_14228,N_14195);
nand U14775 (N_14775,N_14312,N_14182);
and U14776 (N_14776,N_14110,N_14286);
xor U14777 (N_14777,N_14319,N_14204);
or U14778 (N_14778,N_14272,N_14138);
or U14779 (N_14779,N_14465,N_14340);
xnor U14780 (N_14780,N_14346,N_14229);
nand U14781 (N_14781,N_14209,N_14376);
nand U14782 (N_14782,N_14322,N_14438);
nor U14783 (N_14783,N_14248,N_14366);
nand U14784 (N_14784,N_14350,N_14285);
nor U14785 (N_14785,N_14329,N_14477);
nand U14786 (N_14786,N_14475,N_14442);
nand U14787 (N_14787,N_14171,N_14244);
xor U14788 (N_14788,N_14089,N_14365);
or U14789 (N_14789,N_14245,N_14001);
nor U14790 (N_14790,N_14003,N_14371);
or U14791 (N_14791,N_14092,N_14377);
and U14792 (N_14792,N_14086,N_14461);
xnor U14793 (N_14793,N_14119,N_14357);
nand U14794 (N_14794,N_14211,N_14117);
nand U14795 (N_14795,N_14091,N_14015);
or U14796 (N_14796,N_14443,N_14298);
nor U14797 (N_14797,N_14220,N_14388);
nor U14798 (N_14798,N_14432,N_14142);
nand U14799 (N_14799,N_14061,N_14441);
or U14800 (N_14800,N_14375,N_14310);
or U14801 (N_14801,N_14339,N_14482);
xor U14802 (N_14802,N_14053,N_14374);
and U14803 (N_14803,N_14410,N_14075);
xnor U14804 (N_14804,N_14432,N_14120);
xor U14805 (N_14805,N_14283,N_14276);
and U14806 (N_14806,N_14365,N_14316);
and U14807 (N_14807,N_14006,N_14155);
and U14808 (N_14808,N_14466,N_14188);
nor U14809 (N_14809,N_14169,N_14142);
nor U14810 (N_14810,N_14488,N_14133);
nand U14811 (N_14811,N_14421,N_14354);
or U14812 (N_14812,N_14456,N_14293);
or U14813 (N_14813,N_14175,N_14386);
nand U14814 (N_14814,N_14154,N_14391);
and U14815 (N_14815,N_14394,N_14025);
nand U14816 (N_14816,N_14394,N_14297);
xnor U14817 (N_14817,N_14294,N_14385);
nor U14818 (N_14818,N_14473,N_14255);
xor U14819 (N_14819,N_14372,N_14305);
nand U14820 (N_14820,N_14062,N_14464);
and U14821 (N_14821,N_14285,N_14067);
xnor U14822 (N_14822,N_14136,N_14427);
or U14823 (N_14823,N_14118,N_14272);
xor U14824 (N_14824,N_14492,N_14078);
xor U14825 (N_14825,N_14050,N_14134);
nand U14826 (N_14826,N_14042,N_14401);
nor U14827 (N_14827,N_14114,N_14138);
and U14828 (N_14828,N_14190,N_14425);
nor U14829 (N_14829,N_14268,N_14496);
and U14830 (N_14830,N_14122,N_14169);
nor U14831 (N_14831,N_14467,N_14074);
xnor U14832 (N_14832,N_14208,N_14418);
and U14833 (N_14833,N_14151,N_14013);
xor U14834 (N_14834,N_14118,N_14254);
xor U14835 (N_14835,N_14415,N_14231);
xnor U14836 (N_14836,N_14041,N_14276);
or U14837 (N_14837,N_14410,N_14030);
nor U14838 (N_14838,N_14323,N_14344);
and U14839 (N_14839,N_14104,N_14281);
or U14840 (N_14840,N_14176,N_14021);
xor U14841 (N_14841,N_14338,N_14408);
and U14842 (N_14842,N_14445,N_14367);
nand U14843 (N_14843,N_14270,N_14141);
nor U14844 (N_14844,N_14199,N_14068);
xor U14845 (N_14845,N_14154,N_14143);
nand U14846 (N_14846,N_14464,N_14180);
or U14847 (N_14847,N_14274,N_14171);
and U14848 (N_14848,N_14051,N_14149);
or U14849 (N_14849,N_14382,N_14371);
nand U14850 (N_14850,N_14236,N_14156);
nor U14851 (N_14851,N_14223,N_14321);
or U14852 (N_14852,N_14229,N_14164);
nand U14853 (N_14853,N_14253,N_14043);
nand U14854 (N_14854,N_14173,N_14102);
xnor U14855 (N_14855,N_14331,N_14102);
nand U14856 (N_14856,N_14381,N_14477);
nor U14857 (N_14857,N_14082,N_14356);
nand U14858 (N_14858,N_14458,N_14360);
nor U14859 (N_14859,N_14401,N_14110);
xnor U14860 (N_14860,N_14389,N_14263);
nor U14861 (N_14861,N_14085,N_14080);
nor U14862 (N_14862,N_14083,N_14358);
nand U14863 (N_14863,N_14204,N_14469);
or U14864 (N_14864,N_14246,N_14222);
nand U14865 (N_14865,N_14091,N_14059);
xnor U14866 (N_14866,N_14016,N_14185);
and U14867 (N_14867,N_14047,N_14138);
nor U14868 (N_14868,N_14434,N_14229);
or U14869 (N_14869,N_14337,N_14204);
nand U14870 (N_14870,N_14033,N_14156);
or U14871 (N_14871,N_14251,N_14327);
nor U14872 (N_14872,N_14057,N_14366);
nor U14873 (N_14873,N_14187,N_14408);
and U14874 (N_14874,N_14045,N_14225);
nor U14875 (N_14875,N_14180,N_14418);
and U14876 (N_14876,N_14000,N_14163);
nand U14877 (N_14877,N_14405,N_14095);
and U14878 (N_14878,N_14246,N_14452);
nand U14879 (N_14879,N_14292,N_14170);
nand U14880 (N_14880,N_14377,N_14227);
nor U14881 (N_14881,N_14472,N_14448);
and U14882 (N_14882,N_14348,N_14301);
xor U14883 (N_14883,N_14087,N_14275);
nand U14884 (N_14884,N_14287,N_14021);
and U14885 (N_14885,N_14447,N_14295);
nand U14886 (N_14886,N_14184,N_14399);
nor U14887 (N_14887,N_14094,N_14116);
xor U14888 (N_14888,N_14187,N_14381);
nand U14889 (N_14889,N_14366,N_14415);
nor U14890 (N_14890,N_14434,N_14472);
xnor U14891 (N_14891,N_14224,N_14393);
nand U14892 (N_14892,N_14184,N_14480);
or U14893 (N_14893,N_14290,N_14053);
xnor U14894 (N_14894,N_14374,N_14127);
nand U14895 (N_14895,N_14000,N_14186);
nor U14896 (N_14896,N_14038,N_14158);
nand U14897 (N_14897,N_14193,N_14191);
nor U14898 (N_14898,N_14323,N_14085);
nand U14899 (N_14899,N_14037,N_14093);
xor U14900 (N_14900,N_14494,N_14102);
and U14901 (N_14901,N_14328,N_14220);
xor U14902 (N_14902,N_14241,N_14354);
nand U14903 (N_14903,N_14225,N_14345);
and U14904 (N_14904,N_14068,N_14076);
xnor U14905 (N_14905,N_14310,N_14266);
xor U14906 (N_14906,N_14414,N_14487);
xnor U14907 (N_14907,N_14070,N_14115);
nor U14908 (N_14908,N_14003,N_14020);
xnor U14909 (N_14909,N_14429,N_14374);
xnor U14910 (N_14910,N_14419,N_14279);
or U14911 (N_14911,N_14260,N_14461);
xnor U14912 (N_14912,N_14252,N_14388);
and U14913 (N_14913,N_14289,N_14099);
or U14914 (N_14914,N_14349,N_14351);
or U14915 (N_14915,N_14278,N_14110);
or U14916 (N_14916,N_14064,N_14214);
nor U14917 (N_14917,N_14438,N_14293);
nor U14918 (N_14918,N_14126,N_14065);
nor U14919 (N_14919,N_14065,N_14184);
nor U14920 (N_14920,N_14198,N_14072);
xor U14921 (N_14921,N_14445,N_14186);
nor U14922 (N_14922,N_14079,N_14048);
nor U14923 (N_14923,N_14163,N_14264);
or U14924 (N_14924,N_14344,N_14185);
nor U14925 (N_14925,N_14107,N_14219);
or U14926 (N_14926,N_14088,N_14159);
nor U14927 (N_14927,N_14329,N_14387);
nor U14928 (N_14928,N_14417,N_14335);
and U14929 (N_14929,N_14265,N_14036);
or U14930 (N_14930,N_14291,N_14020);
and U14931 (N_14931,N_14231,N_14249);
xor U14932 (N_14932,N_14249,N_14111);
xnor U14933 (N_14933,N_14303,N_14249);
nor U14934 (N_14934,N_14485,N_14265);
or U14935 (N_14935,N_14479,N_14398);
and U14936 (N_14936,N_14256,N_14081);
and U14937 (N_14937,N_14083,N_14266);
nor U14938 (N_14938,N_14095,N_14468);
xnor U14939 (N_14939,N_14133,N_14374);
xnor U14940 (N_14940,N_14291,N_14312);
nor U14941 (N_14941,N_14191,N_14330);
nand U14942 (N_14942,N_14279,N_14448);
or U14943 (N_14943,N_14185,N_14102);
or U14944 (N_14944,N_14204,N_14242);
xor U14945 (N_14945,N_14076,N_14457);
or U14946 (N_14946,N_14365,N_14325);
and U14947 (N_14947,N_14062,N_14117);
or U14948 (N_14948,N_14430,N_14185);
or U14949 (N_14949,N_14218,N_14466);
nand U14950 (N_14950,N_14379,N_14071);
and U14951 (N_14951,N_14455,N_14165);
xor U14952 (N_14952,N_14229,N_14252);
or U14953 (N_14953,N_14129,N_14195);
xnor U14954 (N_14954,N_14474,N_14352);
nor U14955 (N_14955,N_14132,N_14435);
nor U14956 (N_14956,N_14292,N_14328);
and U14957 (N_14957,N_14417,N_14366);
and U14958 (N_14958,N_14442,N_14135);
or U14959 (N_14959,N_14111,N_14489);
nor U14960 (N_14960,N_14197,N_14142);
xor U14961 (N_14961,N_14021,N_14174);
nand U14962 (N_14962,N_14360,N_14371);
nor U14963 (N_14963,N_14137,N_14218);
xnor U14964 (N_14964,N_14044,N_14432);
or U14965 (N_14965,N_14084,N_14088);
nand U14966 (N_14966,N_14365,N_14160);
and U14967 (N_14967,N_14360,N_14331);
nand U14968 (N_14968,N_14206,N_14105);
or U14969 (N_14969,N_14002,N_14171);
xnor U14970 (N_14970,N_14054,N_14484);
and U14971 (N_14971,N_14034,N_14230);
or U14972 (N_14972,N_14164,N_14176);
or U14973 (N_14973,N_14424,N_14225);
nor U14974 (N_14974,N_14171,N_14059);
and U14975 (N_14975,N_14189,N_14181);
nand U14976 (N_14976,N_14281,N_14031);
nor U14977 (N_14977,N_14317,N_14044);
nand U14978 (N_14978,N_14093,N_14162);
or U14979 (N_14979,N_14331,N_14070);
and U14980 (N_14980,N_14433,N_14454);
and U14981 (N_14981,N_14494,N_14417);
nor U14982 (N_14982,N_14214,N_14224);
and U14983 (N_14983,N_14139,N_14107);
nand U14984 (N_14984,N_14398,N_14282);
and U14985 (N_14985,N_14296,N_14297);
or U14986 (N_14986,N_14368,N_14202);
xor U14987 (N_14987,N_14229,N_14291);
xor U14988 (N_14988,N_14186,N_14057);
nor U14989 (N_14989,N_14248,N_14121);
xnor U14990 (N_14990,N_14000,N_14112);
and U14991 (N_14991,N_14341,N_14009);
and U14992 (N_14992,N_14417,N_14469);
or U14993 (N_14993,N_14366,N_14338);
xor U14994 (N_14994,N_14252,N_14139);
or U14995 (N_14995,N_14026,N_14347);
or U14996 (N_14996,N_14498,N_14374);
xnor U14997 (N_14997,N_14486,N_14314);
and U14998 (N_14998,N_14017,N_14204);
nand U14999 (N_14999,N_14371,N_14183);
nor U15000 (N_15000,N_14981,N_14904);
nor U15001 (N_15001,N_14745,N_14688);
nand U15002 (N_15002,N_14986,N_14830);
nor U15003 (N_15003,N_14679,N_14621);
and U15004 (N_15004,N_14984,N_14847);
or U15005 (N_15005,N_14531,N_14812);
nor U15006 (N_15006,N_14942,N_14881);
and U15007 (N_15007,N_14795,N_14558);
nor U15008 (N_15008,N_14713,N_14910);
nand U15009 (N_15009,N_14577,N_14726);
or U15010 (N_15010,N_14890,N_14537);
and U15011 (N_15011,N_14896,N_14870);
nand U15012 (N_15012,N_14846,N_14868);
nor U15013 (N_15013,N_14746,N_14978);
or U15014 (N_15014,N_14883,N_14584);
nand U15015 (N_15015,N_14946,N_14778);
and U15016 (N_15016,N_14667,N_14856);
or U15017 (N_15017,N_14902,N_14564);
nor U15018 (N_15018,N_14853,N_14855);
or U15019 (N_15019,N_14808,N_14570);
nor U15020 (N_15020,N_14832,N_14598);
xor U15021 (N_15021,N_14791,N_14801);
nor U15022 (N_15022,N_14879,N_14604);
or U15023 (N_15023,N_14661,N_14843);
or U15024 (N_15024,N_14916,N_14572);
nand U15025 (N_15025,N_14543,N_14692);
and U15026 (N_15026,N_14612,N_14716);
and U15027 (N_15027,N_14642,N_14618);
nor U15028 (N_15028,N_14687,N_14546);
nor U15029 (N_15029,N_14770,N_14614);
or U15030 (N_15030,N_14752,N_14833);
or U15031 (N_15031,N_14566,N_14857);
nor U15032 (N_15032,N_14559,N_14960);
nand U15033 (N_15033,N_14913,N_14571);
and U15034 (N_15034,N_14660,N_14605);
nand U15035 (N_15035,N_14888,N_14625);
xor U15036 (N_15036,N_14500,N_14641);
or U15037 (N_15037,N_14880,N_14554);
nand U15038 (N_15038,N_14810,N_14644);
xnor U15039 (N_15039,N_14908,N_14794);
xnor U15040 (N_15040,N_14875,N_14809);
and U15041 (N_15041,N_14934,N_14529);
and U15042 (N_15042,N_14979,N_14668);
nand U15043 (N_15043,N_14924,N_14517);
and U15044 (N_15044,N_14758,N_14547);
nor U15045 (N_15045,N_14613,N_14734);
nor U15046 (N_15046,N_14903,N_14686);
nand U15047 (N_15047,N_14754,N_14820);
xnor U15048 (N_15048,N_14760,N_14623);
nor U15049 (N_15049,N_14825,N_14602);
xor U15050 (N_15050,N_14741,N_14672);
and U15051 (N_15051,N_14740,N_14608);
and U15052 (N_15052,N_14592,N_14819);
xnor U15053 (N_15053,N_14957,N_14884);
nand U15054 (N_15054,N_14907,N_14528);
nor U15055 (N_15055,N_14973,N_14961);
xor U15056 (N_15056,N_14938,N_14548);
and U15057 (N_15057,N_14575,N_14863);
or U15058 (N_15058,N_14627,N_14501);
and U15059 (N_15059,N_14985,N_14899);
xor U15060 (N_15060,N_14982,N_14639);
xor U15061 (N_15061,N_14536,N_14640);
nor U15062 (N_15062,N_14698,N_14690);
nand U15063 (N_15063,N_14510,N_14802);
and U15064 (N_15064,N_14553,N_14783);
or U15065 (N_15065,N_14542,N_14527);
xor U15066 (N_15066,N_14603,N_14675);
and U15067 (N_15067,N_14892,N_14790);
nor U15068 (N_15068,N_14658,N_14622);
xor U15069 (N_15069,N_14538,N_14911);
nor U15070 (N_15070,N_14711,N_14583);
nand U15071 (N_15071,N_14872,N_14862);
and U15072 (N_15072,N_14798,N_14694);
xnor U15073 (N_15073,N_14504,N_14624);
or U15074 (N_15074,N_14834,N_14750);
nand U15075 (N_15075,N_14703,N_14997);
or U15076 (N_15076,N_14940,N_14764);
or U15077 (N_15077,N_14839,N_14681);
nor U15078 (N_15078,N_14851,N_14920);
or U15079 (N_15079,N_14817,N_14917);
nand U15080 (N_15080,N_14912,N_14569);
nand U15081 (N_15081,N_14905,N_14785);
and U15082 (N_15082,N_14789,N_14539);
nand U15083 (N_15083,N_14959,N_14534);
or U15084 (N_15084,N_14777,N_14988);
and U15085 (N_15085,N_14962,N_14873);
xnor U15086 (N_15086,N_14967,N_14898);
and U15087 (N_15087,N_14599,N_14926);
xor U15088 (N_15088,N_14742,N_14663);
and U15089 (N_15089,N_14669,N_14666);
xor U15090 (N_15090,N_14532,N_14611);
nand U15091 (N_15091,N_14943,N_14844);
xor U15092 (N_15092,N_14803,N_14933);
and U15093 (N_15093,N_14751,N_14989);
and U15094 (N_15094,N_14677,N_14582);
nor U15095 (N_15095,N_14909,N_14953);
nor U15096 (N_15096,N_14710,N_14866);
and U15097 (N_15097,N_14673,N_14956);
xnor U15098 (N_15098,N_14871,N_14990);
nor U15099 (N_15099,N_14594,N_14719);
xor U15100 (N_15100,N_14755,N_14861);
nor U15101 (N_15101,N_14561,N_14607);
nor U15102 (N_15102,N_14523,N_14771);
or U15103 (N_15103,N_14776,N_14586);
nor U15104 (N_15104,N_14796,N_14519);
or U15105 (N_15105,N_14815,N_14779);
nand U15106 (N_15106,N_14511,N_14993);
and U15107 (N_15107,N_14983,N_14712);
xor U15108 (N_15108,N_14650,N_14665);
and U15109 (N_15109,N_14972,N_14772);
xor U15110 (N_15110,N_14767,N_14593);
nand U15111 (N_15111,N_14514,N_14709);
nand U15112 (N_15112,N_14601,N_14645);
nor U15113 (N_15113,N_14841,N_14784);
xnor U15114 (N_15114,N_14701,N_14968);
and U15115 (N_15115,N_14590,N_14509);
xnor U15116 (N_15116,N_14724,N_14674);
and U15117 (N_15117,N_14632,N_14574);
nand U15118 (N_15118,N_14678,N_14797);
nand U15119 (N_15119,N_14518,N_14876);
and U15120 (N_15120,N_14971,N_14963);
xnor U15121 (N_15121,N_14524,N_14922);
nand U15122 (N_15122,N_14634,N_14630);
or U15123 (N_15123,N_14991,N_14704);
xnor U15124 (N_15124,N_14705,N_14515);
nor U15125 (N_15125,N_14721,N_14860);
xor U15126 (N_15126,N_14878,N_14588);
xnor U15127 (N_15127,N_14762,N_14620);
xnor U15128 (N_15128,N_14761,N_14889);
nor U15129 (N_15129,N_14929,N_14685);
nand U15130 (N_15130,N_14657,N_14521);
nor U15131 (N_15131,N_14507,N_14567);
xor U15132 (N_15132,N_14749,N_14702);
nand U15133 (N_15133,N_14782,N_14522);
and U15134 (N_15134,N_14949,N_14900);
and U15135 (N_15135,N_14662,N_14693);
xor U15136 (N_15136,N_14508,N_14680);
nor U15137 (N_15137,N_14718,N_14581);
nand U15138 (N_15138,N_14768,N_14747);
nor U15139 (N_15139,N_14941,N_14823);
or U15140 (N_15140,N_14565,N_14813);
nand U15141 (N_15141,N_14576,N_14787);
or U15142 (N_15142,N_14733,N_14696);
nor U15143 (N_15143,N_14732,N_14748);
xor U15144 (N_15144,N_14540,N_14597);
nor U15145 (N_15145,N_14720,N_14763);
or U15146 (N_15146,N_14589,N_14901);
nor U15147 (N_15147,N_14928,N_14579);
or U15148 (N_15148,N_14649,N_14864);
or U15149 (N_15149,N_14897,N_14974);
or U15150 (N_15150,N_14757,N_14894);
nand U15151 (N_15151,N_14513,N_14895);
nand U15152 (N_15152,N_14970,N_14730);
nor U15153 (N_15153,N_14637,N_14914);
or U15154 (N_15154,N_14775,N_14932);
or U15155 (N_15155,N_14887,N_14882);
or U15156 (N_15156,N_14617,N_14502);
nand U15157 (N_15157,N_14648,N_14838);
nand U15158 (N_15158,N_14786,N_14891);
and U15159 (N_15159,N_14654,N_14948);
nand U15160 (N_15160,N_14780,N_14950);
xnor U15161 (N_15161,N_14944,N_14736);
xnor U15162 (N_15162,N_14512,N_14999);
nor U15163 (N_15163,N_14852,N_14969);
xnor U15164 (N_15164,N_14549,N_14845);
xnor U15165 (N_15165,N_14918,N_14715);
or U15166 (N_15166,N_14708,N_14939);
and U15167 (N_15167,N_14792,N_14552);
nor U15168 (N_15168,N_14506,N_14628);
nor U15169 (N_15169,N_14615,N_14850);
nor U15170 (N_15170,N_14655,N_14869);
and U15171 (N_15171,N_14842,N_14927);
xor U15172 (N_15172,N_14865,N_14563);
or U15173 (N_15173,N_14631,N_14725);
or U15174 (N_15174,N_14930,N_14947);
or U15175 (N_15175,N_14952,N_14753);
and U15176 (N_15176,N_14859,N_14619);
nor U15177 (N_15177,N_14773,N_14626);
or U15178 (N_15178,N_14544,N_14699);
xnor U15179 (N_15179,N_14555,N_14729);
xnor U15180 (N_15180,N_14965,N_14723);
or U15181 (N_15181,N_14633,N_14530);
nor U15182 (N_15182,N_14580,N_14854);
and U15183 (N_15183,N_14828,N_14849);
and U15184 (N_15184,N_14585,N_14664);
nand U15185 (N_15185,N_14684,N_14717);
and U15186 (N_15186,N_14966,N_14811);
nand U15187 (N_15187,N_14659,N_14822);
or U15188 (N_15188,N_14526,N_14831);
nor U15189 (N_15189,N_14714,N_14996);
or U15190 (N_15190,N_14893,N_14638);
nand U15191 (N_15191,N_14806,N_14995);
nor U15192 (N_15192,N_14635,N_14818);
and U15193 (N_15193,N_14551,N_14573);
xnor U15194 (N_15194,N_14652,N_14606);
nor U15195 (N_15195,N_14520,N_14562);
nor U15196 (N_15196,N_14931,N_14925);
and U15197 (N_15197,N_14799,N_14557);
nand U15198 (N_15198,N_14656,N_14837);
xor U15199 (N_15199,N_14814,N_14816);
nor U15200 (N_15200,N_14700,N_14840);
or U15201 (N_15201,N_14835,N_14505);
or U15202 (N_15202,N_14731,N_14919);
xor U15203 (N_15203,N_14695,N_14756);
nor U15204 (N_15204,N_14568,N_14738);
nor U15205 (N_15205,N_14743,N_14643);
nand U15206 (N_15206,N_14682,N_14964);
or U15207 (N_15207,N_14578,N_14765);
nor U15208 (N_15208,N_14980,N_14937);
xor U15209 (N_15209,N_14616,N_14992);
nand U15210 (N_15210,N_14722,N_14885);
nand U15211 (N_15211,N_14535,N_14936);
or U15212 (N_15212,N_14556,N_14824);
and U15213 (N_15213,N_14848,N_14646);
and U15214 (N_15214,N_14503,N_14759);
xor U15215 (N_15215,N_14706,N_14671);
nand U15216 (N_15216,N_14945,N_14976);
and U15217 (N_15217,N_14977,N_14766);
nand U15218 (N_15218,N_14821,N_14629);
nand U15219 (N_15219,N_14739,N_14954);
or U15220 (N_15220,N_14951,N_14525);
or U15221 (N_15221,N_14923,N_14805);
xor U15222 (N_15222,N_14600,N_14827);
and U15223 (N_15223,N_14735,N_14781);
nor U15224 (N_15224,N_14533,N_14915);
nand U15225 (N_15225,N_14728,N_14935);
nand U15226 (N_15226,N_14550,N_14877);
or U15227 (N_15227,N_14800,N_14595);
nor U15228 (N_15228,N_14829,N_14921);
xnor U15229 (N_15229,N_14591,N_14636);
and U15230 (N_15230,N_14958,N_14998);
nor U15231 (N_15231,N_14804,N_14545);
nor U15232 (N_15232,N_14737,N_14867);
xnor U15233 (N_15233,N_14807,N_14874);
xnor U15234 (N_15234,N_14858,N_14955);
nand U15235 (N_15235,N_14609,N_14769);
and U15236 (N_15236,N_14653,N_14691);
xor U15237 (N_15237,N_14516,N_14676);
and U15238 (N_15238,N_14670,N_14994);
nand U15239 (N_15239,N_14689,N_14697);
and U15240 (N_15240,N_14906,N_14727);
xor U15241 (N_15241,N_14788,N_14541);
xor U15242 (N_15242,N_14975,N_14683);
xnor U15243 (N_15243,N_14826,N_14774);
xor U15244 (N_15244,N_14707,N_14744);
nor U15245 (N_15245,N_14560,N_14793);
and U15246 (N_15246,N_14886,N_14587);
xnor U15247 (N_15247,N_14651,N_14596);
or U15248 (N_15248,N_14647,N_14987);
nand U15249 (N_15249,N_14610,N_14836);
nand U15250 (N_15250,N_14850,N_14526);
or U15251 (N_15251,N_14768,N_14962);
nand U15252 (N_15252,N_14639,N_14689);
nor U15253 (N_15253,N_14532,N_14936);
and U15254 (N_15254,N_14749,N_14617);
nand U15255 (N_15255,N_14790,N_14978);
and U15256 (N_15256,N_14867,N_14994);
nor U15257 (N_15257,N_14723,N_14787);
nor U15258 (N_15258,N_14875,N_14562);
xnor U15259 (N_15259,N_14857,N_14773);
nor U15260 (N_15260,N_14809,N_14946);
or U15261 (N_15261,N_14747,N_14921);
and U15262 (N_15262,N_14686,N_14605);
and U15263 (N_15263,N_14514,N_14950);
nor U15264 (N_15264,N_14904,N_14521);
and U15265 (N_15265,N_14839,N_14952);
nor U15266 (N_15266,N_14957,N_14791);
and U15267 (N_15267,N_14625,N_14736);
and U15268 (N_15268,N_14995,N_14880);
nand U15269 (N_15269,N_14504,N_14678);
nor U15270 (N_15270,N_14709,N_14598);
xnor U15271 (N_15271,N_14741,N_14605);
and U15272 (N_15272,N_14513,N_14748);
nor U15273 (N_15273,N_14512,N_14594);
nand U15274 (N_15274,N_14816,N_14995);
nor U15275 (N_15275,N_14750,N_14998);
xnor U15276 (N_15276,N_14992,N_14679);
xnor U15277 (N_15277,N_14873,N_14831);
or U15278 (N_15278,N_14536,N_14780);
nand U15279 (N_15279,N_14934,N_14587);
or U15280 (N_15280,N_14591,N_14725);
nand U15281 (N_15281,N_14709,N_14922);
and U15282 (N_15282,N_14822,N_14912);
or U15283 (N_15283,N_14674,N_14777);
or U15284 (N_15284,N_14905,N_14997);
or U15285 (N_15285,N_14549,N_14852);
nand U15286 (N_15286,N_14611,N_14941);
and U15287 (N_15287,N_14845,N_14611);
nor U15288 (N_15288,N_14951,N_14615);
and U15289 (N_15289,N_14792,N_14892);
or U15290 (N_15290,N_14895,N_14607);
nor U15291 (N_15291,N_14875,N_14842);
xnor U15292 (N_15292,N_14741,N_14535);
and U15293 (N_15293,N_14504,N_14805);
or U15294 (N_15294,N_14522,N_14847);
or U15295 (N_15295,N_14717,N_14760);
or U15296 (N_15296,N_14932,N_14952);
or U15297 (N_15297,N_14753,N_14554);
nand U15298 (N_15298,N_14731,N_14866);
nand U15299 (N_15299,N_14786,N_14544);
or U15300 (N_15300,N_14913,N_14756);
or U15301 (N_15301,N_14585,N_14599);
nand U15302 (N_15302,N_14731,N_14938);
nor U15303 (N_15303,N_14953,N_14677);
and U15304 (N_15304,N_14952,N_14945);
nand U15305 (N_15305,N_14884,N_14801);
nor U15306 (N_15306,N_14794,N_14976);
xnor U15307 (N_15307,N_14690,N_14531);
xnor U15308 (N_15308,N_14984,N_14870);
xnor U15309 (N_15309,N_14857,N_14996);
and U15310 (N_15310,N_14908,N_14930);
or U15311 (N_15311,N_14680,N_14627);
nor U15312 (N_15312,N_14522,N_14824);
or U15313 (N_15313,N_14772,N_14829);
nor U15314 (N_15314,N_14968,N_14891);
xnor U15315 (N_15315,N_14703,N_14561);
nand U15316 (N_15316,N_14811,N_14784);
nor U15317 (N_15317,N_14924,N_14795);
nor U15318 (N_15318,N_14859,N_14934);
nor U15319 (N_15319,N_14893,N_14826);
or U15320 (N_15320,N_14636,N_14533);
and U15321 (N_15321,N_14949,N_14789);
and U15322 (N_15322,N_14512,N_14733);
and U15323 (N_15323,N_14693,N_14721);
nor U15324 (N_15324,N_14782,N_14692);
nor U15325 (N_15325,N_14979,N_14614);
and U15326 (N_15326,N_14755,N_14772);
nor U15327 (N_15327,N_14795,N_14745);
nand U15328 (N_15328,N_14683,N_14674);
nand U15329 (N_15329,N_14613,N_14693);
and U15330 (N_15330,N_14737,N_14966);
nor U15331 (N_15331,N_14943,N_14640);
xor U15332 (N_15332,N_14877,N_14635);
nand U15333 (N_15333,N_14687,N_14915);
nand U15334 (N_15334,N_14734,N_14576);
or U15335 (N_15335,N_14587,N_14593);
nand U15336 (N_15336,N_14964,N_14768);
xor U15337 (N_15337,N_14669,N_14671);
and U15338 (N_15338,N_14824,N_14636);
xnor U15339 (N_15339,N_14967,N_14506);
nor U15340 (N_15340,N_14751,N_14754);
nor U15341 (N_15341,N_14543,N_14634);
nor U15342 (N_15342,N_14816,N_14620);
nor U15343 (N_15343,N_14986,N_14539);
nor U15344 (N_15344,N_14876,N_14587);
and U15345 (N_15345,N_14514,N_14920);
and U15346 (N_15346,N_14696,N_14833);
or U15347 (N_15347,N_14719,N_14604);
and U15348 (N_15348,N_14785,N_14976);
and U15349 (N_15349,N_14661,N_14539);
or U15350 (N_15350,N_14606,N_14540);
xnor U15351 (N_15351,N_14583,N_14616);
and U15352 (N_15352,N_14794,N_14796);
xnor U15353 (N_15353,N_14790,N_14688);
nor U15354 (N_15354,N_14761,N_14940);
nand U15355 (N_15355,N_14716,N_14770);
nor U15356 (N_15356,N_14867,N_14522);
or U15357 (N_15357,N_14787,N_14910);
or U15358 (N_15358,N_14713,N_14846);
or U15359 (N_15359,N_14745,N_14579);
or U15360 (N_15360,N_14844,N_14848);
and U15361 (N_15361,N_14784,N_14518);
nand U15362 (N_15362,N_14700,N_14503);
nand U15363 (N_15363,N_14966,N_14526);
xnor U15364 (N_15364,N_14638,N_14846);
or U15365 (N_15365,N_14610,N_14587);
and U15366 (N_15366,N_14761,N_14514);
or U15367 (N_15367,N_14713,N_14518);
nor U15368 (N_15368,N_14519,N_14960);
nor U15369 (N_15369,N_14801,N_14581);
or U15370 (N_15370,N_14636,N_14891);
and U15371 (N_15371,N_14556,N_14806);
and U15372 (N_15372,N_14903,N_14716);
xor U15373 (N_15373,N_14978,N_14970);
and U15374 (N_15374,N_14870,N_14531);
xor U15375 (N_15375,N_14875,N_14920);
nor U15376 (N_15376,N_14822,N_14850);
and U15377 (N_15377,N_14968,N_14916);
and U15378 (N_15378,N_14550,N_14588);
and U15379 (N_15379,N_14816,N_14662);
or U15380 (N_15380,N_14613,N_14574);
nor U15381 (N_15381,N_14753,N_14883);
or U15382 (N_15382,N_14727,N_14794);
xnor U15383 (N_15383,N_14592,N_14931);
or U15384 (N_15384,N_14638,N_14783);
and U15385 (N_15385,N_14831,N_14960);
and U15386 (N_15386,N_14751,N_14738);
or U15387 (N_15387,N_14602,N_14555);
and U15388 (N_15388,N_14724,N_14523);
xor U15389 (N_15389,N_14997,N_14951);
or U15390 (N_15390,N_14739,N_14544);
and U15391 (N_15391,N_14665,N_14764);
nor U15392 (N_15392,N_14937,N_14565);
or U15393 (N_15393,N_14627,N_14628);
and U15394 (N_15394,N_14926,N_14921);
nand U15395 (N_15395,N_14924,N_14603);
or U15396 (N_15396,N_14777,N_14854);
xnor U15397 (N_15397,N_14510,N_14806);
or U15398 (N_15398,N_14953,N_14519);
nor U15399 (N_15399,N_14504,N_14884);
xor U15400 (N_15400,N_14613,N_14560);
nor U15401 (N_15401,N_14596,N_14616);
and U15402 (N_15402,N_14509,N_14828);
nor U15403 (N_15403,N_14625,N_14920);
and U15404 (N_15404,N_14776,N_14564);
or U15405 (N_15405,N_14997,N_14777);
or U15406 (N_15406,N_14929,N_14510);
and U15407 (N_15407,N_14659,N_14515);
nor U15408 (N_15408,N_14956,N_14751);
xnor U15409 (N_15409,N_14795,N_14589);
and U15410 (N_15410,N_14543,N_14912);
and U15411 (N_15411,N_14830,N_14589);
xor U15412 (N_15412,N_14553,N_14807);
nor U15413 (N_15413,N_14552,N_14581);
nor U15414 (N_15414,N_14935,N_14867);
nor U15415 (N_15415,N_14591,N_14650);
nor U15416 (N_15416,N_14651,N_14698);
and U15417 (N_15417,N_14901,N_14505);
or U15418 (N_15418,N_14716,N_14956);
xor U15419 (N_15419,N_14778,N_14918);
nand U15420 (N_15420,N_14980,N_14710);
and U15421 (N_15421,N_14633,N_14832);
xnor U15422 (N_15422,N_14537,N_14780);
xnor U15423 (N_15423,N_14658,N_14603);
nor U15424 (N_15424,N_14825,N_14948);
nor U15425 (N_15425,N_14919,N_14629);
or U15426 (N_15426,N_14517,N_14636);
and U15427 (N_15427,N_14530,N_14860);
xor U15428 (N_15428,N_14555,N_14553);
xor U15429 (N_15429,N_14892,N_14975);
nor U15430 (N_15430,N_14801,N_14993);
nor U15431 (N_15431,N_14500,N_14540);
xor U15432 (N_15432,N_14785,N_14772);
xor U15433 (N_15433,N_14566,N_14924);
nand U15434 (N_15434,N_14659,N_14681);
xor U15435 (N_15435,N_14656,N_14713);
xor U15436 (N_15436,N_14598,N_14503);
and U15437 (N_15437,N_14648,N_14912);
nor U15438 (N_15438,N_14799,N_14941);
and U15439 (N_15439,N_14788,N_14855);
xnor U15440 (N_15440,N_14677,N_14586);
or U15441 (N_15441,N_14970,N_14590);
or U15442 (N_15442,N_14674,N_14648);
and U15443 (N_15443,N_14951,N_14988);
nand U15444 (N_15444,N_14766,N_14584);
and U15445 (N_15445,N_14528,N_14987);
xor U15446 (N_15446,N_14827,N_14741);
nand U15447 (N_15447,N_14628,N_14526);
or U15448 (N_15448,N_14515,N_14885);
nor U15449 (N_15449,N_14941,N_14645);
nor U15450 (N_15450,N_14897,N_14971);
nor U15451 (N_15451,N_14605,N_14672);
nor U15452 (N_15452,N_14996,N_14870);
nand U15453 (N_15453,N_14781,N_14533);
xnor U15454 (N_15454,N_14775,N_14616);
nor U15455 (N_15455,N_14647,N_14554);
nor U15456 (N_15456,N_14616,N_14700);
xnor U15457 (N_15457,N_14968,N_14704);
or U15458 (N_15458,N_14766,N_14753);
nand U15459 (N_15459,N_14581,N_14608);
or U15460 (N_15460,N_14677,N_14769);
nand U15461 (N_15461,N_14574,N_14791);
and U15462 (N_15462,N_14575,N_14616);
and U15463 (N_15463,N_14854,N_14932);
nand U15464 (N_15464,N_14539,N_14527);
xnor U15465 (N_15465,N_14674,N_14948);
and U15466 (N_15466,N_14815,N_14777);
nand U15467 (N_15467,N_14942,N_14751);
xor U15468 (N_15468,N_14942,N_14759);
nand U15469 (N_15469,N_14781,N_14952);
xnor U15470 (N_15470,N_14801,N_14935);
or U15471 (N_15471,N_14895,N_14867);
and U15472 (N_15472,N_14852,N_14888);
nand U15473 (N_15473,N_14766,N_14855);
nor U15474 (N_15474,N_14677,N_14843);
and U15475 (N_15475,N_14650,N_14851);
nor U15476 (N_15476,N_14542,N_14686);
nand U15477 (N_15477,N_14717,N_14843);
or U15478 (N_15478,N_14546,N_14827);
nand U15479 (N_15479,N_14659,N_14812);
nand U15480 (N_15480,N_14828,N_14646);
xnor U15481 (N_15481,N_14767,N_14777);
xnor U15482 (N_15482,N_14785,N_14862);
nand U15483 (N_15483,N_14977,N_14826);
nand U15484 (N_15484,N_14658,N_14962);
xor U15485 (N_15485,N_14622,N_14540);
or U15486 (N_15486,N_14655,N_14932);
nand U15487 (N_15487,N_14518,N_14874);
nand U15488 (N_15488,N_14606,N_14942);
nand U15489 (N_15489,N_14929,N_14704);
and U15490 (N_15490,N_14531,N_14811);
nand U15491 (N_15491,N_14811,N_14915);
and U15492 (N_15492,N_14854,N_14563);
and U15493 (N_15493,N_14556,N_14533);
nor U15494 (N_15494,N_14963,N_14669);
xor U15495 (N_15495,N_14558,N_14500);
and U15496 (N_15496,N_14967,N_14918);
and U15497 (N_15497,N_14520,N_14522);
xor U15498 (N_15498,N_14592,N_14986);
nand U15499 (N_15499,N_14887,N_14696);
or U15500 (N_15500,N_15038,N_15119);
nand U15501 (N_15501,N_15199,N_15372);
xor U15502 (N_15502,N_15302,N_15023);
nand U15503 (N_15503,N_15024,N_15290);
xnor U15504 (N_15504,N_15462,N_15423);
xor U15505 (N_15505,N_15022,N_15483);
and U15506 (N_15506,N_15354,N_15205);
and U15507 (N_15507,N_15308,N_15149);
or U15508 (N_15508,N_15275,N_15028);
and U15509 (N_15509,N_15360,N_15318);
nor U15510 (N_15510,N_15327,N_15007);
and U15511 (N_15511,N_15320,N_15397);
or U15512 (N_15512,N_15228,N_15027);
xor U15513 (N_15513,N_15217,N_15150);
nand U15514 (N_15514,N_15341,N_15267);
nand U15515 (N_15515,N_15235,N_15059);
or U15516 (N_15516,N_15179,N_15128);
nor U15517 (N_15517,N_15435,N_15427);
xnor U15518 (N_15518,N_15090,N_15230);
nand U15519 (N_15519,N_15388,N_15417);
nand U15520 (N_15520,N_15123,N_15366);
nand U15521 (N_15521,N_15394,N_15133);
and U15522 (N_15522,N_15400,N_15041);
nor U15523 (N_15523,N_15374,N_15345);
and U15524 (N_15524,N_15499,N_15262);
nor U15525 (N_15525,N_15073,N_15068);
and U15526 (N_15526,N_15103,N_15307);
and U15527 (N_15527,N_15032,N_15373);
nor U15528 (N_15528,N_15326,N_15376);
xor U15529 (N_15529,N_15000,N_15305);
and U15530 (N_15530,N_15380,N_15110);
or U15531 (N_15531,N_15138,N_15258);
xnor U15532 (N_15532,N_15132,N_15014);
or U15533 (N_15533,N_15348,N_15448);
or U15534 (N_15534,N_15310,N_15288);
or U15535 (N_15535,N_15282,N_15003);
nor U15536 (N_15536,N_15182,N_15045);
nand U15537 (N_15537,N_15211,N_15050);
nor U15538 (N_15538,N_15304,N_15424);
nor U15539 (N_15539,N_15441,N_15410);
or U15540 (N_15540,N_15192,N_15056);
xnor U15541 (N_15541,N_15364,N_15085);
nand U15542 (N_15542,N_15418,N_15107);
or U15543 (N_15543,N_15171,N_15256);
nor U15544 (N_15544,N_15291,N_15076);
nor U15545 (N_15545,N_15449,N_15033);
nor U15546 (N_15546,N_15472,N_15488);
and U15547 (N_15547,N_15127,N_15439);
xor U15548 (N_15548,N_15195,N_15034);
nor U15549 (N_15549,N_15458,N_15347);
or U15550 (N_15550,N_15100,N_15284);
xnor U15551 (N_15551,N_15289,N_15193);
or U15552 (N_15552,N_15338,N_15158);
xor U15553 (N_15553,N_15203,N_15063);
nor U15554 (N_15554,N_15383,N_15098);
nand U15555 (N_15555,N_15329,N_15316);
nand U15556 (N_15556,N_15286,N_15479);
nor U15557 (N_15557,N_15167,N_15002);
and U15558 (N_15558,N_15361,N_15156);
and U15559 (N_15559,N_15005,N_15241);
nor U15560 (N_15560,N_15493,N_15089);
xnor U15561 (N_15561,N_15096,N_15245);
or U15562 (N_15562,N_15200,N_15064);
and U15563 (N_15563,N_15392,N_15044);
or U15564 (N_15564,N_15274,N_15224);
or U15565 (N_15565,N_15169,N_15359);
nand U15566 (N_15566,N_15476,N_15247);
nor U15567 (N_15567,N_15332,N_15145);
xor U15568 (N_15568,N_15446,N_15351);
and U15569 (N_15569,N_15140,N_15054);
or U15570 (N_15570,N_15060,N_15419);
and U15571 (N_15571,N_15378,N_15434);
or U15572 (N_15572,N_15337,N_15215);
nand U15573 (N_15573,N_15468,N_15066);
nor U15574 (N_15574,N_15019,N_15379);
or U15575 (N_15575,N_15157,N_15188);
or U15576 (N_15576,N_15450,N_15463);
xnor U15577 (N_15577,N_15384,N_15252);
xor U15578 (N_15578,N_15177,N_15105);
nor U15579 (N_15579,N_15148,N_15207);
and U15580 (N_15580,N_15191,N_15092);
xor U15581 (N_15581,N_15020,N_15480);
xnor U15582 (N_15582,N_15225,N_15136);
nor U15583 (N_15583,N_15226,N_15454);
nand U15584 (N_15584,N_15238,N_15111);
nor U15585 (N_15585,N_15264,N_15047);
nand U15586 (N_15586,N_15467,N_15081);
and U15587 (N_15587,N_15248,N_15189);
xor U15588 (N_15588,N_15294,N_15031);
or U15589 (N_15589,N_15381,N_15249);
xnor U15590 (N_15590,N_15117,N_15357);
or U15591 (N_15591,N_15037,N_15026);
nand U15592 (N_15592,N_15018,N_15387);
xnor U15593 (N_15593,N_15349,N_15404);
xor U15594 (N_15594,N_15498,N_15353);
xnor U15595 (N_15595,N_15223,N_15398);
or U15596 (N_15596,N_15058,N_15154);
xnor U15597 (N_15597,N_15227,N_15180);
nor U15598 (N_15598,N_15396,N_15315);
and U15599 (N_15599,N_15280,N_15393);
and U15600 (N_15600,N_15260,N_15429);
xnor U15601 (N_15601,N_15051,N_15276);
xor U15602 (N_15602,N_15287,N_15239);
xor U15603 (N_15603,N_15102,N_15325);
nand U15604 (N_15604,N_15155,N_15414);
nor U15605 (N_15605,N_15080,N_15303);
nor U15606 (N_15606,N_15250,N_15208);
and U15607 (N_15607,N_15415,N_15152);
nand U15608 (N_15608,N_15012,N_15421);
or U15609 (N_15609,N_15244,N_15492);
nor U15610 (N_15610,N_15432,N_15017);
nand U15611 (N_15611,N_15346,N_15481);
xnor U15612 (N_15612,N_15416,N_15444);
xnor U15613 (N_15613,N_15431,N_15229);
xor U15614 (N_15614,N_15144,N_15040);
and U15615 (N_15615,N_15457,N_15162);
or U15616 (N_15616,N_15259,N_15370);
xor U15617 (N_15617,N_15436,N_15489);
or U15618 (N_15618,N_15216,N_15163);
nand U15619 (N_15619,N_15470,N_15395);
or U15620 (N_15620,N_15322,N_15253);
or U15621 (N_15621,N_15413,N_15430);
and U15622 (N_15622,N_15328,N_15030);
nor U15623 (N_15623,N_15084,N_15214);
nor U15624 (N_15624,N_15043,N_15036);
xor U15625 (N_15625,N_15165,N_15135);
or U15626 (N_15626,N_15465,N_15442);
or U15627 (N_15627,N_15283,N_15460);
nor U15628 (N_15628,N_15118,N_15466);
nor U15629 (N_15629,N_15391,N_15129);
or U15630 (N_15630,N_15306,N_15197);
or U15631 (N_15631,N_15382,N_15069);
nand U15632 (N_15632,N_15363,N_15271);
nor U15633 (N_15633,N_15482,N_15173);
and U15634 (N_15634,N_15113,N_15025);
or U15635 (N_15635,N_15496,N_15008);
xnor U15636 (N_15636,N_15447,N_15484);
or U15637 (N_15637,N_15114,N_15141);
nand U15638 (N_15638,N_15281,N_15001);
nand U15639 (N_15639,N_15170,N_15083);
nor U15640 (N_15640,N_15137,N_15049);
nor U15641 (N_15641,N_15340,N_15052);
and U15642 (N_15642,N_15405,N_15218);
or U15643 (N_15643,N_15074,N_15240);
xnor U15644 (N_15644,N_15321,N_15433);
and U15645 (N_15645,N_15234,N_15297);
xor U15646 (N_15646,N_15086,N_15344);
xnor U15647 (N_15647,N_15131,N_15408);
or U15648 (N_15648,N_15082,N_15407);
and U15649 (N_15649,N_15355,N_15469);
or U15650 (N_15650,N_15161,N_15185);
nand U15651 (N_15651,N_15147,N_15194);
nor U15652 (N_15652,N_15166,N_15278);
xor U15653 (N_15653,N_15010,N_15006);
xor U15654 (N_15654,N_15377,N_15295);
and U15655 (N_15655,N_15046,N_15279);
nor U15656 (N_15656,N_15184,N_15485);
xor U15657 (N_15657,N_15257,N_15088);
nor U15658 (N_15658,N_15198,N_15339);
xnor U15659 (N_15659,N_15124,N_15455);
nand U15660 (N_15660,N_15473,N_15143);
xnor U15661 (N_15661,N_15425,N_15079);
xor U15662 (N_15662,N_15070,N_15263);
xnor U15663 (N_15663,N_15285,N_15159);
nand U15664 (N_15664,N_15491,N_15411);
xor U15665 (N_15665,N_15270,N_15266);
xor U15666 (N_15666,N_15035,N_15009);
or U15667 (N_15667,N_15317,N_15209);
and U15668 (N_15668,N_15204,N_15219);
nor U15669 (N_15669,N_15324,N_15101);
xnor U15670 (N_15670,N_15201,N_15115);
and U15671 (N_15671,N_15494,N_15061);
nand U15672 (N_15672,N_15309,N_15269);
xor U15673 (N_15673,N_15330,N_15072);
nor U15674 (N_15674,N_15453,N_15176);
or U15675 (N_15675,N_15146,N_15261);
xnor U15676 (N_15676,N_15222,N_15343);
or U15677 (N_15677,N_15334,N_15236);
or U15678 (N_15678,N_15233,N_15071);
nor U15679 (N_15679,N_15021,N_15095);
or U15680 (N_15680,N_15368,N_15232);
or U15681 (N_15681,N_15385,N_15104);
nor U15682 (N_15682,N_15443,N_15375);
nand U15683 (N_15683,N_15126,N_15186);
and U15684 (N_15684,N_15495,N_15451);
or U15685 (N_15685,N_15471,N_15456);
nor U15686 (N_15686,N_15153,N_15212);
xnor U15687 (N_15687,N_15093,N_15196);
or U15688 (N_15688,N_15277,N_15231);
xnor U15689 (N_15689,N_15190,N_15242);
xnor U15690 (N_15690,N_15273,N_15402);
and U15691 (N_15691,N_15369,N_15172);
xnor U15692 (N_15692,N_15174,N_15301);
nor U15693 (N_15693,N_15160,N_15265);
or U15694 (N_15694,N_15350,N_15464);
xnor U15695 (N_15695,N_15181,N_15210);
or U15696 (N_15696,N_15300,N_15412);
and U15697 (N_15697,N_15087,N_15106);
xnor U15698 (N_15698,N_15142,N_15039);
or U15699 (N_15699,N_15445,N_15125);
or U15700 (N_15700,N_15108,N_15202);
and U15701 (N_15701,N_15178,N_15251);
and U15702 (N_15702,N_15055,N_15004);
nand U15703 (N_15703,N_15389,N_15386);
or U15704 (N_15704,N_15367,N_15246);
nor U15705 (N_15705,N_15116,N_15094);
nand U15706 (N_15706,N_15091,N_15139);
nand U15707 (N_15707,N_15314,N_15065);
nor U15708 (N_15708,N_15099,N_15365);
nor U15709 (N_15709,N_15220,N_15352);
xor U15710 (N_15710,N_15187,N_15356);
or U15711 (N_15711,N_15122,N_15296);
xnor U15712 (N_15712,N_15490,N_15335);
nand U15713 (N_15713,N_15438,N_15168);
xor U15714 (N_15714,N_15486,N_15062);
and U15715 (N_15715,N_15243,N_15475);
xnor U15716 (N_15716,N_15120,N_15406);
nor U15717 (N_15717,N_15075,N_15053);
and U15718 (N_15718,N_15461,N_15097);
nor U15719 (N_15719,N_15323,N_15134);
xnor U15720 (N_15720,N_15311,N_15057);
and U15721 (N_15721,N_15221,N_15077);
xnor U15722 (N_15722,N_15151,N_15362);
xor U15723 (N_15723,N_15440,N_15497);
and U15724 (N_15724,N_15409,N_15130);
or U15725 (N_15725,N_15254,N_15015);
xor U15726 (N_15726,N_15371,N_15298);
nand U15727 (N_15727,N_15428,N_15401);
nand U15728 (N_15728,N_15067,N_15478);
nand U15729 (N_15729,N_15477,N_15164);
nand U15730 (N_15730,N_15206,N_15422);
or U15731 (N_15731,N_15333,N_15319);
nor U15732 (N_15732,N_15312,N_15013);
xor U15733 (N_15733,N_15358,N_15313);
xnor U15734 (N_15734,N_15272,N_15299);
and U15735 (N_15735,N_15078,N_15331);
nand U15736 (N_15736,N_15342,N_15011);
nor U15737 (N_15737,N_15293,N_15255);
xor U15738 (N_15738,N_15426,N_15390);
or U15739 (N_15739,N_15459,N_15403);
xor U15740 (N_15740,N_15048,N_15183);
nand U15741 (N_15741,N_15292,N_15175);
nor U15742 (N_15742,N_15016,N_15237);
nand U15743 (N_15743,N_15399,N_15437);
nor U15744 (N_15744,N_15487,N_15452);
or U15745 (N_15745,N_15420,N_15109);
xor U15746 (N_15746,N_15121,N_15112);
nand U15747 (N_15747,N_15213,N_15268);
xor U15748 (N_15748,N_15474,N_15042);
nand U15749 (N_15749,N_15336,N_15029);
and U15750 (N_15750,N_15105,N_15146);
nand U15751 (N_15751,N_15306,N_15205);
nand U15752 (N_15752,N_15380,N_15330);
nand U15753 (N_15753,N_15417,N_15336);
or U15754 (N_15754,N_15426,N_15183);
and U15755 (N_15755,N_15223,N_15376);
and U15756 (N_15756,N_15224,N_15144);
xor U15757 (N_15757,N_15395,N_15198);
nor U15758 (N_15758,N_15393,N_15126);
and U15759 (N_15759,N_15219,N_15472);
and U15760 (N_15760,N_15120,N_15205);
and U15761 (N_15761,N_15276,N_15480);
nand U15762 (N_15762,N_15000,N_15306);
xnor U15763 (N_15763,N_15233,N_15127);
xnor U15764 (N_15764,N_15118,N_15062);
and U15765 (N_15765,N_15396,N_15198);
nor U15766 (N_15766,N_15320,N_15403);
xnor U15767 (N_15767,N_15414,N_15298);
or U15768 (N_15768,N_15262,N_15306);
xnor U15769 (N_15769,N_15354,N_15039);
and U15770 (N_15770,N_15055,N_15398);
nand U15771 (N_15771,N_15378,N_15212);
and U15772 (N_15772,N_15260,N_15062);
or U15773 (N_15773,N_15398,N_15375);
xor U15774 (N_15774,N_15175,N_15219);
nand U15775 (N_15775,N_15321,N_15492);
or U15776 (N_15776,N_15162,N_15352);
nor U15777 (N_15777,N_15181,N_15324);
xnor U15778 (N_15778,N_15348,N_15053);
nor U15779 (N_15779,N_15276,N_15086);
xnor U15780 (N_15780,N_15438,N_15468);
nor U15781 (N_15781,N_15085,N_15187);
or U15782 (N_15782,N_15110,N_15164);
and U15783 (N_15783,N_15049,N_15077);
nand U15784 (N_15784,N_15465,N_15435);
or U15785 (N_15785,N_15036,N_15250);
or U15786 (N_15786,N_15095,N_15138);
and U15787 (N_15787,N_15145,N_15124);
nand U15788 (N_15788,N_15484,N_15370);
nand U15789 (N_15789,N_15085,N_15083);
and U15790 (N_15790,N_15087,N_15182);
nor U15791 (N_15791,N_15306,N_15461);
xor U15792 (N_15792,N_15076,N_15130);
xor U15793 (N_15793,N_15068,N_15312);
xor U15794 (N_15794,N_15396,N_15065);
and U15795 (N_15795,N_15181,N_15446);
and U15796 (N_15796,N_15068,N_15122);
and U15797 (N_15797,N_15183,N_15211);
or U15798 (N_15798,N_15140,N_15112);
nand U15799 (N_15799,N_15127,N_15486);
and U15800 (N_15800,N_15449,N_15066);
nand U15801 (N_15801,N_15494,N_15012);
xor U15802 (N_15802,N_15347,N_15046);
or U15803 (N_15803,N_15155,N_15340);
and U15804 (N_15804,N_15293,N_15188);
and U15805 (N_15805,N_15025,N_15135);
nor U15806 (N_15806,N_15446,N_15071);
or U15807 (N_15807,N_15045,N_15017);
and U15808 (N_15808,N_15337,N_15396);
xor U15809 (N_15809,N_15298,N_15238);
nand U15810 (N_15810,N_15446,N_15093);
and U15811 (N_15811,N_15250,N_15163);
nand U15812 (N_15812,N_15413,N_15359);
nor U15813 (N_15813,N_15122,N_15471);
or U15814 (N_15814,N_15499,N_15271);
or U15815 (N_15815,N_15200,N_15342);
nand U15816 (N_15816,N_15109,N_15113);
nor U15817 (N_15817,N_15328,N_15246);
nand U15818 (N_15818,N_15286,N_15454);
or U15819 (N_15819,N_15262,N_15003);
nand U15820 (N_15820,N_15230,N_15144);
nor U15821 (N_15821,N_15148,N_15050);
nand U15822 (N_15822,N_15164,N_15499);
nor U15823 (N_15823,N_15355,N_15210);
and U15824 (N_15824,N_15079,N_15138);
xnor U15825 (N_15825,N_15433,N_15199);
nand U15826 (N_15826,N_15258,N_15178);
nand U15827 (N_15827,N_15253,N_15401);
nand U15828 (N_15828,N_15039,N_15226);
and U15829 (N_15829,N_15357,N_15104);
and U15830 (N_15830,N_15205,N_15258);
xnor U15831 (N_15831,N_15335,N_15200);
nor U15832 (N_15832,N_15421,N_15380);
or U15833 (N_15833,N_15454,N_15271);
xnor U15834 (N_15834,N_15099,N_15361);
nand U15835 (N_15835,N_15400,N_15212);
nor U15836 (N_15836,N_15337,N_15053);
nand U15837 (N_15837,N_15280,N_15383);
nand U15838 (N_15838,N_15233,N_15017);
xor U15839 (N_15839,N_15156,N_15427);
nor U15840 (N_15840,N_15183,N_15242);
nand U15841 (N_15841,N_15437,N_15051);
nor U15842 (N_15842,N_15171,N_15138);
and U15843 (N_15843,N_15443,N_15330);
nand U15844 (N_15844,N_15040,N_15156);
xnor U15845 (N_15845,N_15071,N_15124);
and U15846 (N_15846,N_15343,N_15394);
nor U15847 (N_15847,N_15028,N_15003);
xnor U15848 (N_15848,N_15286,N_15164);
nand U15849 (N_15849,N_15478,N_15471);
or U15850 (N_15850,N_15051,N_15196);
xor U15851 (N_15851,N_15409,N_15070);
and U15852 (N_15852,N_15454,N_15456);
or U15853 (N_15853,N_15093,N_15473);
xor U15854 (N_15854,N_15353,N_15008);
or U15855 (N_15855,N_15066,N_15069);
or U15856 (N_15856,N_15012,N_15241);
nand U15857 (N_15857,N_15305,N_15092);
and U15858 (N_15858,N_15262,N_15330);
and U15859 (N_15859,N_15431,N_15090);
nand U15860 (N_15860,N_15344,N_15006);
or U15861 (N_15861,N_15207,N_15320);
or U15862 (N_15862,N_15054,N_15129);
nand U15863 (N_15863,N_15429,N_15322);
nand U15864 (N_15864,N_15212,N_15376);
nand U15865 (N_15865,N_15053,N_15264);
nor U15866 (N_15866,N_15371,N_15011);
xnor U15867 (N_15867,N_15371,N_15407);
nor U15868 (N_15868,N_15108,N_15225);
or U15869 (N_15869,N_15360,N_15492);
nand U15870 (N_15870,N_15064,N_15021);
xnor U15871 (N_15871,N_15173,N_15155);
or U15872 (N_15872,N_15243,N_15350);
and U15873 (N_15873,N_15423,N_15146);
or U15874 (N_15874,N_15058,N_15185);
nor U15875 (N_15875,N_15451,N_15051);
nor U15876 (N_15876,N_15131,N_15082);
nand U15877 (N_15877,N_15242,N_15294);
nand U15878 (N_15878,N_15157,N_15088);
nor U15879 (N_15879,N_15085,N_15218);
and U15880 (N_15880,N_15054,N_15485);
or U15881 (N_15881,N_15308,N_15243);
nand U15882 (N_15882,N_15348,N_15145);
nand U15883 (N_15883,N_15052,N_15010);
nor U15884 (N_15884,N_15118,N_15149);
and U15885 (N_15885,N_15052,N_15216);
nand U15886 (N_15886,N_15271,N_15340);
nand U15887 (N_15887,N_15161,N_15397);
xor U15888 (N_15888,N_15135,N_15092);
nand U15889 (N_15889,N_15371,N_15045);
and U15890 (N_15890,N_15081,N_15163);
nor U15891 (N_15891,N_15400,N_15250);
nor U15892 (N_15892,N_15138,N_15461);
and U15893 (N_15893,N_15201,N_15178);
and U15894 (N_15894,N_15303,N_15156);
xnor U15895 (N_15895,N_15195,N_15491);
xor U15896 (N_15896,N_15436,N_15143);
nand U15897 (N_15897,N_15360,N_15049);
nand U15898 (N_15898,N_15183,N_15060);
nor U15899 (N_15899,N_15100,N_15031);
nand U15900 (N_15900,N_15004,N_15014);
nand U15901 (N_15901,N_15324,N_15409);
xnor U15902 (N_15902,N_15243,N_15177);
nor U15903 (N_15903,N_15496,N_15312);
nand U15904 (N_15904,N_15231,N_15247);
and U15905 (N_15905,N_15454,N_15427);
and U15906 (N_15906,N_15391,N_15387);
nor U15907 (N_15907,N_15221,N_15268);
nand U15908 (N_15908,N_15122,N_15142);
and U15909 (N_15909,N_15108,N_15126);
or U15910 (N_15910,N_15138,N_15380);
nand U15911 (N_15911,N_15351,N_15488);
nand U15912 (N_15912,N_15046,N_15012);
nor U15913 (N_15913,N_15496,N_15464);
nand U15914 (N_15914,N_15109,N_15440);
nor U15915 (N_15915,N_15020,N_15037);
nor U15916 (N_15916,N_15288,N_15080);
or U15917 (N_15917,N_15098,N_15464);
nor U15918 (N_15918,N_15348,N_15420);
and U15919 (N_15919,N_15021,N_15191);
xnor U15920 (N_15920,N_15307,N_15096);
or U15921 (N_15921,N_15039,N_15476);
or U15922 (N_15922,N_15294,N_15350);
xor U15923 (N_15923,N_15356,N_15294);
nand U15924 (N_15924,N_15086,N_15104);
and U15925 (N_15925,N_15117,N_15046);
nor U15926 (N_15926,N_15406,N_15148);
or U15927 (N_15927,N_15292,N_15362);
xor U15928 (N_15928,N_15245,N_15284);
nand U15929 (N_15929,N_15029,N_15267);
nand U15930 (N_15930,N_15123,N_15268);
or U15931 (N_15931,N_15290,N_15171);
or U15932 (N_15932,N_15471,N_15183);
nand U15933 (N_15933,N_15438,N_15097);
or U15934 (N_15934,N_15217,N_15029);
nand U15935 (N_15935,N_15327,N_15207);
or U15936 (N_15936,N_15351,N_15038);
xor U15937 (N_15937,N_15244,N_15391);
nor U15938 (N_15938,N_15258,N_15496);
or U15939 (N_15939,N_15499,N_15351);
nor U15940 (N_15940,N_15439,N_15482);
and U15941 (N_15941,N_15047,N_15118);
and U15942 (N_15942,N_15103,N_15221);
nand U15943 (N_15943,N_15301,N_15035);
and U15944 (N_15944,N_15488,N_15465);
or U15945 (N_15945,N_15158,N_15132);
or U15946 (N_15946,N_15123,N_15385);
and U15947 (N_15947,N_15049,N_15351);
and U15948 (N_15948,N_15345,N_15415);
or U15949 (N_15949,N_15222,N_15130);
xor U15950 (N_15950,N_15336,N_15378);
and U15951 (N_15951,N_15270,N_15131);
or U15952 (N_15952,N_15046,N_15020);
nor U15953 (N_15953,N_15088,N_15358);
nand U15954 (N_15954,N_15499,N_15113);
xor U15955 (N_15955,N_15237,N_15151);
nand U15956 (N_15956,N_15165,N_15225);
xnor U15957 (N_15957,N_15471,N_15139);
xnor U15958 (N_15958,N_15450,N_15243);
nand U15959 (N_15959,N_15394,N_15082);
nand U15960 (N_15960,N_15160,N_15152);
and U15961 (N_15961,N_15293,N_15163);
and U15962 (N_15962,N_15325,N_15016);
and U15963 (N_15963,N_15288,N_15213);
or U15964 (N_15964,N_15027,N_15257);
xor U15965 (N_15965,N_15217,N_15196);
or U15966 (N_15966,N_15034,N_15098);
nor U15967 (N_15967,N_15146,N_15451);
and U15968 (N_15968,N_15467,N_15251);
or U15969 (N_15969,N_15490,N_15342);
nor U15970 (N_15970,N_15309,N_15421);
or U15971 (N_15971,N_15095,N_15413);
and U15972 (N_15972,N_15248,N_15111);
and U15973 (N_15973,N_15308,N_15465);
and U15974 (N_15974,N_15346,N_15136);
and U15975 (N_15975,N_15428,N_15167);
nor U15976 (N_15976,N_15375,N_15428);
or U15977 (N_15977,N_15012,N_15135);
nand U15978 (N_15978,N_15156,N_15155);
or U15979 (N_15979,N_15196,N_15434);
nand U15980 (N_15980,N_15225,N_15114);
or U15981 (N_15981,N_15238,N_15462);
nand U15982 (N_15982,N_15174,N_15189);
nor U15983 (N_15983,N_15350,N_15009);
and U15984 (N_15984,N_15363,N_15056);
xor U15985 (N_15985,N_15253,N_15064);
nand U15986 (N_15986,N_15055,N_15208);
or U15987 (N_15987,N_15041,N_15453);
nor U15988 (N_15988,N_15343,N_15160);
nand U15989 (N_15989,N_15025,N_15142);
nand U15990 (N_15990,N_15205,N_15150);
or U15991 (N_15991,N_15388,N_15059);
or U15992 (N_15992,N_15270,N_15099);
nor U15993 (N_15993,N_15344,N_15270);
or U15994 (N_15994,N_15386,N_15180);
xnor U15995 (N_15995,N_15169,N_15187);
and U15996 (N_15996,N_15200,N_15296);
nor U15997 (N_15997,N_15328,N_15014);
or U15998 (N_15998,N_15403,N_15451);
xnor U15999 (N_15999,N_15283,N_15468);
xor U16000 (N_16000,N_15661,N_15649);
or U16001 (N_16001,N_15585,N_15544);
and U16002 (N_16002,N_15796,N_15799);
xnor U16003 (N_16003,N_15528,N_15631);
nor U16004 (N_16004,N_15640,N_15687);
xor U16005 (N_16005,N_15988,N_15579);
nand U16006 (N_16006,N_15907,N_15981);
or U16007 (N_16007,N_15668,N_15549);
or U16008 (N_16008,N_15985,N_15627);
nor U16009 (N_16009,N_15896,N_15790);
nor U16010 (N_16010,N_15626,N_15674);
nor U16011 (N_16011,N_15580,N_15503);
nand U16012 (N_16012,N_15708,N_15535);
nor U16013 (N_16013,N_15866,N_15732);
xor U16014 (N_16014,N_15846,N_15712);
or U16015 (N_16015,N_15863,N_15702);
nand U16016 (N_16016,N_15798,N_15679);
nand U16017 (N_16017,N_15760,N_15812);
nor U16018 (N_16018,N_15805,N_15758);
xor U16019 (N_16019,N_15887,N_15598);
and U16020 (N_16020,N_15736,N_15891);
and U16021 (N_16021,N_15728,N_15787);
and U16022 (N_16022,N_15641,N_15623);
nand U16023 (N_16023,N_15709,N_15939);
and U16024 (N_16024,N_15664,N_15688);
nor U16025 (N_16025,N_15883,N_15817);
nand U16026 (N_16026,N_15703,N_15856);
or U16027 (N_16027,N_15783,N_15828);
and U16028 (N_16028,N_15947,N_15734);
xor U16029 (N_16029,N_15884,N_15693);
nor U16030 (N_16030,N_15595,N_15808);
nand U16031 (N_16031,N_15786,N_15807);
and U16032 (N_16032,N_15739,N_15726);
xnor U16033 (N_16033,N_15992,N_15841);
xor U16034 (N_16034,N_15672,N_15989);
nand U16035 (N_16035,N_15830,N_15659);
xnor U16036 (N_16036,N_15605,N_15554);
xnor U16037 (N_16037,N_15754,N_15762);
nand U16038 (N_16038,N_15721,N_15978);
nand U16039 (N_16039,N_15685,N_15872);
nor U16040 (N_16040,N_15952,N_15592);
and U16041 (N_16041,N_15657,N_15510);
or U16042 (N_16042,N_15602,N_15570);
xor U16043 (N_16043,N_15636,N_15561);
and U16044 (N_16044,N_15660,N_15635);
nor U16045 (N_16045,N_15996,N_15651);
or U16046 (N_16046,N_15792,N_15761);
xor U16047 (N_16047,N_15862,N_15612);
nor U16048 (N_16048,N_15615,N_15700);
and U16049 (N_16049,N_15844,N_15673);
and U16050 (N_16050,N_15861,N_15853);
and U16051 (N_16051,N_15902,N_15848);
and U16052 (N_16052,N_15776,N_15583);
nor U16053 (N_16053,N_15670,N_15698);
nor U16054 (N_16054,N_15885,N_15669);
nand U16055 (N_16055,N_15738,N_15677);
nor U16056 (N_16056,N_15737,N_15713);
nor U16057 (N_16057,N_15578,N_15513);
and U16058 (N_16058,N_15625,N_15845);
nand U16059 (N_16059,N_15825,N_15874);
or U16060 (N_16060,N_15780,N_15928);
and U16061 (N_16061,N_15600,N_15961);
nor U16062 (N_16062,N_15611,N_15701);
or U16063 (N_16063,N_15753,N_15869);
or U16064 (N_16064,N_15847,N_15935);
nor U16065 (N_16065,N_15944,N_15691);
or U16066 (N_16066,N_15684,N_15534);
nor U16067 (N_16067,N_15973,N_15552);
nand U16068 (N_16068,N_15620,N_15781);
or U16069 (N_16069,N_15810,N_15750);
and U16070 (N_16070,N_15921,N_15678);
xnor U16071 (N_16071,N_15894,N_15840);
and U16072 (N_16072,N_15746,N_15962);
and U16073 (N_16073,N_15994,N_15924);
or U16074 (N_16074,N_15551,N_15536);
and U16075 (N_16075,N_15901,N_15507);
xnor U16076 (N_16076,N_15642,N_15873);
or U16077 (N_16077,N_15904,N_15865);
nand U16078 (N_16078,N_15643,N_15991);
nand U16079 (N_16079,N_15953,N_15692);
nand U16080 (N_16080,N_15868,N_15936);
nor U16081 (N_16081,N_15725,N_15813);
xnor U16082 (N_16082,N_15997,N_15826);
and U16083 (N_16083,N_15983,N_15929);
and U16084 (N_16084,N_15543,N_15722);
and U16085 (N_16085,N_15607,N_15878);
or U16086 (N_16086,N_15571,N_15715);
and U16087 (N_16087,N_15859,N_15882);
nand U16088 (N_16088,N_15850,N_15804);
xnor U16089 (N_16089,N_15852,N_15594);
and U16090 (N_16090,N_15770,N_15509);
xnor U16091 (N_16091,N_15638,N_15771);
nor U16092 (N_16092,N_15619,N_15654);
and U16093 (N_16093,N_15724,N_15658);
or U16094 (N_16094,N_15697,N_15656);
xnor U16095 (N_16095,N_15773,N_15779);
nor U16096 (N_16096,N_15849,N_15705);
and U16097 (N_16097,N_15562,N_15714);
nand U16098 (N_16098,N_15681,N_15979);
or U16099 (N_16099,N_15806,N_15880);
or U16100 (N_16100,N_15506,N_15795);
nor U16101 (N_16101,N_15912,N_15504);
xor U16102 (N_16102,N_15555,N_15857);
or U16103 (N_16103,N_15752,N_15957);
and U16104 (N_16104,N_15926,N_15606);
nor U16105 (N_16105,N_15662,N_15596);
xnor U16106 (N_16106,N_15557,N_15976);
and U16107 (N_16107,N_15995,N_15519);
and U16108 (N_16108,N_15964,N_15614);
or U16109 (N_16109,N_15876,N_15785);
nor U16110 (N_16110,N_15581,N_15563);
nor U16111 (N_16111,N_15788,N_15689);
xnor U16112 (N_16112,N_15778,N_15937);
or U16113 (N_16113,N_15809,N_15864);
xnor U16114 (N_16114,N_15609,N_15676);
xnor U16115 (N_16115,N_15502,N_15586);
xnor U16116 (N_16116,N_15731,N_15803);
and U16117 (N_16117,N_15816,N_15858);
nand U16118 (N_16118,N_15839,N_15624);
or U16119 (N_16119,N_15637,N_15984);
xnor U16120 (N_16120,N_15965,N_15966);
xnor U16121 (N_16121,N_15815,N_15980);
nand U16122 (N_16122,N_15634,N_15843);
and U16123 (N_16123,N_15515,N_15608);
or U16124 (N_16124,N_15717,N_15801);
or U16125 (N_16125,N_15742,N_15524);
xor U16126 (N_16126,N_15572,N_15851);
nand U16127 (N_16127,N_15889,N_15834);
or U16128 (N_16128,N_15512,N_15900);
nor U16129 (N_16129,N_15967,N_15617);
nand U16130 (N_16130,N_15899,N_15516);
nand U16131 (N_16131,N_15910,N_15764);
and U16132 (N_16132,N_15974,N_15759);
nor U16133 (N_16133,N_15919,N_15821);
and U16134 (N_16134,N_15639,N_15956);
or U16135 (N_16135,N_15730,N_15559);
nor U16136 (N_16136,N_15610,N_15719);
and U16137 (N_16137,N_15975,N_15946);
nor U16138 (N_16138,N_15768,N_15723);
xor U16139 (N_16139,N_15720,N_15727);
and U16140 (N_16140,N_15569,N_15632);
and U16141 (N_16141,N_15749,N_15584);
or U16142 (N_16142,N_15818,N_15916);
and U16143 (N_16143,N_15767,N_15782);
or U16144 (N_16144,N_15622,N_15751);
and U16145 (N_16145,N_15597,N_15526);
nand U16146 (N_16146,N_15576,N_15802);
nand U16147 (N_16147,N_15893,N_15542);
and U16148 (N_16148,N_15895,N_15913);
xor U16149 (N_16149,N_15567,N_15824);
nand U16150 (N_16150,N_15890,N_15518);
and U16151 (N_16151,N_15917,N_15932);
or U16152 (N_16152,N_15970,N_15838);
xor U16153 (N_16153,N_15525,N_15682);
xnor U16154 (N_16154,N_15582,N_15558);
and U16155 (N_16155,N_15998,N_15833);
nor U16156 (N_16156,N_15699,N_15565);
nor U16157 (N_16157,N_15941,N_15925);
or U16158 (N_16158,N_15500,N_15982);
nand U16159 (N_16159,N_15945,N_15690);
nor U16160 (N_16160,N_15575,N_15948);
xnor U16161 (N_16161,N_15886,N_15573);
or U16162 (N_16162,N_15867,N_15747);
nand U16163 (N_16163,N_15560,N_15905);
or U16164 (N_16164,N_15735,N_15621);
or U16165 (N_16165,N_15832,N_15514);
or U16166 (N_16166,N_15538,N_15694);
nor U16167 (N_16167,N_15718,N_15879);
nor U16168 (N_16168,N_15971,N_15539);
nand U16169 (N_16169,N_15743,N_15791);
xnor U16170 (N_16170,N_15537,N_15505);
and U16171 (N_16171,N_15603,N_15613);
and U16172 (N_16172,N_15556,N_15855);
nand U16173 (N_16173,N_15784,N_15836);
and U16174 (N_16174,N_15666,N_15501);
nor U16175 (N_16175,N_15529,N_15593);
nor U16176 (N_16176,N_15875,N_15909);
nand U16177 (N_16177,N_15523,N_15986);
nand U16178 (N_16178,N_15527,N_15577);
nor U16179 (N_16179,N_15508,N_15811);
nor U16180 (N_16180,N_15566,N_15881);
nand U16181 (N_16181,N_15871,N_15548);
nand U16182 (N_16182,N_15568,N_15530);
and U16183 (N_16183,N_15820,N_15740);
nor U16184 (N_16184,N_15765,N_15616);
nand U16185 (N_16185,N_15633,N_15757);
or U16186 (N_16186,N_15564,N_15835);
xnor U16187 (N_16187,N_15628,N_15915);
nor U16188 (N_16188,N_15860,N_15533);
nor U16189 (N_16189,N_15958,N_15706);
or U16190 (N_16190,N_15521,N_15541);
or U16191 (N_16191,N_15733,N_15774);
nand U16192 (N_16192,N_15831,N_15763);
xnor U16193 (N_16193,N_15903,N_15748);
or U16194 (N_16194,N_15898,N_15938);
nand U16195 (N_16195,N_15959,N_15954);
xnor U16196 (N_16196,N_15990,N_15653);
xnor U16197 (N_16197,N_15794,N_15553);
and U16198 (N_16198,N_15827,N_15604);
or U16199 (N_16199,N_15854,N_15711);
or U16200 (N_16200,N_15644,N_15511);
or U16201 (N_16201,N_15665,N_15745);
nor U16202 (N_16202,N_15829,N_15531);
nor U16203 (N_16203,N_15842,N_15695);
nor U16204 (N_16204,N_15630,N_15987);
or U16205 (N_16205,N_15977,N_15772);
nor U16206 (N_16206,N_15671,N_15675);
and U16207 (N_16207,N_15645,N_15897);
or U16208 (N_16208,N_15601,N_15696);
or U16209 (N_16209,N_15972,N_15766);
and U16210 (N_16210,N_15927,N_15546);
xor U16211 (N_16211,N_15940,N_15650);
nand U16212 (N_16212,N_15591,N_15968);
nor U16213 (N_16213,N_15655,N_15933);
and U16214 (N_16214,N_15920,N_15589);
or U16215 (N_16215,N_15793,N_15943);
and U16216 (N_16216,N_15520,N_15822);
and U16217 (N_16217,N_15629,N_15663);
and U16218 (N_16218,N_15906,N_15908);
and U16219 (N_16219,N_15618,N_15814);
nand U16220 (N_16220,N_15888,N_15707);
nand U16221 (N_16221,N_15797,N_15532);
nand U16222 (N_16222,N_15969,N_15789);
xor U16223 (N_16223,N_15686,N_15942);
and U16224 (N_16224,N_15545,N_15769);
nor U16225 (N_16225,N_15777,N_15547);
or U16226 (N_16226,N_15930,N_15574);
nand U16227 (N_16227,N_15680,N_15934);
nor U16228 (N_16228,N_15652,N_15923);
xnor U16229 (N_16229,N_15540,N_15522);
nor U16230 (N_16230,N_15918,N_15710);
or U16231 (N_16231,N_15667,N_15588);
and U16232 (N_16232,N_15922,N_15951);
nand U16233 (N_16233,N_15716,N_15955);
or U16234 (N_16234,N_15999,N_15755);
or U16235 (N_16235,N_15590,N_15800);
xor U16236 (N_16236,N_15931,N_15744);
xor U16237 (N_16237,N_15517,N_15683);
nor U16238 (N_16238,N_15911,N_15819);
or U16239 (N_16239,N_15775,N_15993);
xnor U16240 (N_16240,N_15960,N_15892);
and U16241 (N_16241,N_15648,N_15646);
or U16242 (N_16242,N_15756,N_15950);
and U16243 (N_16243,N_15877,N_15949);
or U16244 (N_16244,N_15704,N_15729);
nand U16245 (N_16245,N_15647,N_15837);
xnor U16246 (N_16246,N_15963,N_15587);
and U16247 (N_16247,N_15870,N_15599);
nand U16248 (N_16248,N_15823,N_15914);
xnor U16249 (N_16249,N_15550,N_15741);
nand U16250 (N_16250,N_15928,N_15982);
nor U16251 (N_16251,N_15720,N_15760);
nand U16252 (N_16252,N_15819,N_15539);
xor U16253 (N_16253,N_15704,N_15608);
nor U16254 (N_16254,N_15670,N_15699);
nor U16255 (N_16255,N_15926,N_15756);
and U16256 (N_16256,N_15964,N_15914);
xor U16257 (N_16257,N_15566,N_15875);
or U16258 (N_16258,N_15573,N_15670);
or U16259 (N_16259,N_15814,N_15753);
or U16260 (N_16260,N_15915,N_15525);
nor U16261 (N_16261,N_15780,N_15927);
nor U16262 (N_16262,N_15755,N_15976);
nor U16263 (N_16263,N_15692,N_15689);
xnor U16264 (N_16264,N_15760,N_15620);
xnor U16265 (N_16265,N_15869,N_15953);
nor U16266 (N_16266,N_15504,N_15769);
nor U16267 (N_16267,N_15579,N_15676);
and U16268 (N_16268,N_15850,N_15743);
nand U16269 (N_16269,N_15844,N_15768);
nor U16270 (N_16270,N_15876,N_15660);
nand U16271 (N_16271,N_15865,N_15614);
and U16272 (N_16272,N_15574,N_15887);
and U16273 (N_16273,N_15922,N_15515);
and U16274 (N_16274,N_15631,N_15541);
or U16275 (N_16275,N_15926,N_15636);
and U16276 (N_16276,N_15894,N_15668);
nor U16277 (N_16277,N_15603,N_15609);
or U16278 (N_16278,N_15751,N_15573);
or U16279 (N_16279,N_15988,N_15838);
xor U16280 (N_16280,N_15593,N_15821);
or U16281 (N_16281,N_15551,N_15682);
nand U16282 (N_16282,N_15763,N_15870);
or U16283 (N_16283,N_15998,N_15617);
and U16284 (N_16284,N_15507,N_15744);
and U16285 (N_16285,N_15602,N_15751);
or U16286 (N_16286,N_15515,N_15647);
and U16287 (N_16287,N_15576,N_15700);
xor U16288 (N_16288,N_15856,N_15610);
or U16289 (N_16289,N_15557,N_15970);
and U16290 (N_16290,N_15911,N_15775);
nor U16291 (N_16291,N_15627,N_15802);
xor U16292 (N_16292,N_15751,N_15516);
or U16293 (N_16293,N_15650,N_15956);
nor U16294 (N_16294,N_15886,N_15640);
and U16295 (N_16295,N_15512,N_15923);
nor U16296 (N_16296,N_15708,N_15537);
nand U16297 (N_16297,N_15750,N_15531);
nand U16298 (N_16298,N_15522,N_15880);
nand U16299 (N_16299,N_15900,N_15668);
nand U16300 (N_16300,N_15678,N_15688);
nor U16301 (N_16301,N_15918,N_15507);
and U16302 (N_16302,N_15766,N_15715);
and U16303 (N_16303,N_15860,N_15648);
nor U16304 (N_16304,N_15691,N_15618);
and U16305 (N_16305,N_15597,N_15605);
xor U16306 (N_16306,N_15914,N_15954);
and U16307 (N_16307,N_15880,N_15505);
nand U16308 (N_16308,N_15583,N_15591);
or U16309 (N_16309,N_15857,N_15888);
nor U16310 (N_16310,N_15564,N_15775);
nor U16311 (N_16311,N_15527,N_15692);
nand U16312 (N_16312,N_15599,N_15572);
nand U16313 (N_16313,N_15877,N_15982);
and U16314 (N_16314,N_15903,N_15873);
xnor U16315 (N_16315,N_15874,N_15898);
nand U16316 (N_16316,N_15696,N_15653);
and U16317 (N_16317,N_15632,N_15617);
and U16318 (N_16318,N_15925,N_15835);
or U16319 (N_16319,N_15641,N_15826);
nand U16320 (N_16320,N_15945,N_15597);
nor U16321 (N_16321,N_15773,N_15555);
or U16322 (N_16322,N_15587,N_15710);
and U16323 (N_16323,N_15622,N_15911);
nor U16324 (N_16324,N_15590,N_15931);
and U16325 (N_16325,N_15530,N_15838);
and U16326 (N_16326,N_15898,N_15522);
xor U16327 (N_16327,N_15867,N_15977);
nand U16328 (N_16328,N_15743,N_15762);
or U16329 (N_16329,N_15573,N_15728);
or U16330 (N_16330,N_15546,N_15636);
and U16331 (N_16331,N_15765,N_15653);
nor U16332 (N_16332,N_15945,N_15599);
xnor U16333 (N_16333,N_15950,N_15792);
and U16334 (N_16334,N_15856,N_15953);
nand U16335 (N_16335,N_15798,N_15542);
xor U16336 (N_16336,N_15835,N_15516);
xnor U16337 (N_16337,N_15801,N_15917);
nand U16338 (N_16338,N_15920,N_15929);
xor U16339 (N_16339,N_15850,N_15916);
and U16340 (N_16340,N_15537,N_15927);
or U16341 (N_16341,N_15503,N_15541);
xor U16342 (N_16342,N_15546,N_15749);
xor U16343 (N_16343,N_15640,N_15834);
nor U16344 (N_16344,N_15749,N_15854);
and U16345 (N_16345,N_15522,N_15628);
or U16346 (N_16346,N_15890,N_15859);
and U16347 (N_16347,N_15959,N_15723);
and U16348 (N_16348,N_15974,N_15647);
xor U16349 (N_16349,N_15987,N_15596);
xnor U16350 (N_16350,N_15507,N_15877);
and U16351 (N_16351,N_15573,N_15615);
or U16352 (N_16352,N_15586,N_15688);
xor U16353 (N_16353,N_15646,N_15823);
nand U16354 (N_16354,N_15999,N_15938);
nand U16355 (N_16355,N_15670,N_15564);
xor U16356 (N_16356,N_15943,N_15665);
or U16357 (N_16357,N_15857,N_15612);
or U16358 (N_16358,N_15672,N_15594);
xnor U16359 (N_16359,N_15754,N_15963);
and U16360 (N_16360,N_15506,N_15893);
and U16361 (N_16361,N_15980,N_15966);
nand U16362 (N_16362,N_15989,N_15805);
xnor U16363 (N_16363,N_15751,N_15790);
or U16364 (N_16364,N_15988,N_15858);
xor U16365 (N_16365,N_15520,N_15714);
xnor U16366 (N_16366,N_15870,N_15734);
xnor U16367 (N_16367,N_15787,N_15601);
and U16368 (N_16368,N_15508,N_15768);
nor U16369 (N_16369,N_15726,N_15620);
xnor U16370 (N_16370,N_15903,N_15740);
nand U16371 (N_16371,N_15924,N_15683);
nor U16372 (N_16372,N_15925,N_15768);
nand U16373 (N_16373,N_15890,N_15936);
and U16374 (N_16374,N_15903,N_15719);
xnor U16375 (N_16375,N_15621,N_15672);
and U16376 (N_16376,N_15642,N_15581);
nor U16377 (N_16377,N_15819,N_15551);
or U16378 (N_16378,N_15557,N_15939);
and U16379 (N_16379,N_15672,N_15840);
nor U16380 (N_16380,N_15599,N_15778);
xnor U16381 (N_16381,N_15808,N_15787);
nand U16382 (N_16382,N_15967,N_15570);
and U16383 (N_16383,N_15722,N_15705);
and U16384 (N_16384,N_15725,N_15584);
nand U16385 (N_16385,N_15677,N_15910);
nand U16386 (N_16386,N_15980,N_15592);
xnor U16387 (N_16387,N_15902,N_15661);
nor U16388 (N_16388,N_15985,N_15640);
nor U16389 (N_16389,N_15886,N_15938);
nor U16390 (N_16390,N_15719,N_15590);
nand U16391 (N_16391,N_15599,N_15529);
xor U16392 (N_16392,N_15501,N_15792);
nor U16393 (N_16393,N_15626,N_15990);
and U16394 (N_16394,N_15553,N_15893);
and U16395 (N_16395,N_15658,N_15523);
nor U16396 (N_16396,N_15552,N_15860);
nor U16397 (N_16397,N_15706,N_15613);
xnor U16398 (N_16398,N_15604,N_15884);
or U16399 (N_16399,N_15662,N_15693);
or U16400 (N_16400,N_15798,N_15574);
or U16401 (N_16401,N_15765,N_15612);
and U16402 (N_16402,N_15576,N_15608);
nand U16403 (N_16403,N_15885,N_15638);
xor U16404 (N_16404,N_15749,N_15599);
or U16405 (N_16405,N_15726,N_15744);
or U16406 (N_16406,N_15508,N_15576);
or U16407 (N_16407,N_15561,N_15935);
and U16408 (N_16408,N_15876,N_15746);
xor U16409 (N_16409,N_15647,N_15582);
xor U16410 (N_16410,N_15643,N_15768);
and U16411 (N_16411,N_15837,N_15537);
and U16412 (N_16412,N_15565,N_15678);
nor U16413 (N_16413,N_15842,N_15863);
or U16414 (N_16414,N_15616,N_15768);
xnor U16415 (N_16415,N_15905,N_15769);
nor U16416 (N_16416,N_15794,N_15863);
nor U16417 (N_16417,N_15689,N_15570);
nand U16418 (N_16418,N_15889,N_15976);
nand U16419 (N_16419,N_15696,N_15568);
and U16420 (N_16420,N_15725,N_15520);
and U16421 (N_16421,N_15885,N_15927);
xor U16422 (N_16422,N_15573,N_15796);
or U16423 (N_16423,N_15988,N_15997);
and U16424 (N_16424,N_15876,N_15815);
xor U16425 (N_16425,N_15556,N_15644);
nand U16426 (N_16426,N_15963,N_15525);
or U16427 (N_16427,N_15524,N_15993);
or U16428 (N_16428,N_15676,N_15779);
nand U16429 (N_16429,N_15893,N_15541);
nand U16430 (N_16430,N_15518,N_15935);
nor U16431 (N_16431,N_15509,N_15730);
xor U16432 (N_16432,N_15719,N_15555);
nor U16433 (N_16433,N_15957,N_15833);
xor U16434 (N_16434,N_15947,N_15822);
nand U16435 (N_16435,N_15838,N_15895);
nand U16436 (N_16436,N_15522,N_15545);
and U16437 (N_16437,N_15689,N_15620);
xor U16438 (N_16438,N_15695,N_15871);
xnor U16439 (N_16439,N_15657,N_15752);
or U16440 (N_16440,N_15588,N_15987);
nand U16441 (N_16441,N_15885,N_15936);
and U16442 (N_16442,N_15718,N_15848);
nor U16443 (N_16443,N_15855,N_15664);
and U16444 (N_16444,N_15880,N_15738);
and U16445 (N_16445,N_15582,N_15683);
or U16446 (N_16446,N_15835,N_15769);
and U16447 (N_16447,N_15689,N_15584);
xor U16448 (N_16448,N_15968,N_15999);
or U16449 (N_16449,N_15934,N_15842);
nor U16450 (N_16450,N_15719,N_15818);
xnor U16451 (N_16451,N_15604,N_15593);
xor U16452 (N_16452,N_15661,N_15730);
xnor U16453 (N_16453,N_15718,N_15713);
or U16454 (N_16454,N_15983,N_15979);
or U16455 (N_16455,N_15696,N_15806);
xnor U16456 (N_16456,N_15705,N_15927);
and U16457 (N_16457,N_15718,N_15731);
or U16458 (N_16458,N_15817,N_15865);
or U16459 (N_16459,N_15695,N_15970);
xor U16460 (N_16460,N_15810,N_15938);
or U16461 (N_16461,N_15793,N_15533);
xnor U16462 (N_16462,N_15500,N_15851);
nor U16463 (N_16463,N_15740,N_15608);
xor U16464 (N_16464,N_15699,N_15609);
nor U16465 (N_16465,N_15552,N_15835);
or U16466 (N_16466,N_15521,N_15749);
and U16467 (N_16467,N_15740,N_15790);
and U16468 (N_16468,N_15987,N_15644);
or U16469 (N_16469,N_15687,N_15635);
nor U16470 (N_16470,N_15932,N_15739);
nor U16471 (N_16471,N_15878,N_15666);
and U16472 (N_16472,N_15767,N_15801);
nand U16473 (N_16473,N_15887,N_15819);
nand U16474 (N_16474,N_15854,N_15941);
nor U16475 (N_16475,N_15946,N_15720);
nor U16476 (N_16476,N_15997,N_15545);
xnor U16477 (N_16477,N_15835,N_15932);
or U16478 (N_16478,N_15810,N_15763);
nor U16479 (N_16479,N_15992,N_15979);
or U16480 (N_16480,N_15772,N_15628);
nor U16481 (N_16481,N_15678,N_15895);
and U16482 (N_16482,N_15924,N_15517);
xor U16483 (N_16483,N_15715,N_15558);
or U16484 (N_16484,N_15695,N_15853);
nand U16485 (N_16485,N_15685,N_15504);
xor U16486 (N_16486,N_15908,N_15648);
nor U16487 (N_16487,N_15571,N_15745);
nand U16488 (N_16488,N_15591,N_15909);
and U16489 (N_16489,N_15731,N_15649);
nand U16490 (N_16490,N_15514,N_15985);
nor U16491 (N_16491,N_15865,N_15818);
or U16492 (N_16492,N_15666,N_15988);
nor U16493 (N_16493,N_15524,N_15656);
nor U16494 (N_16494,N_15659,N_15664);
or U16495 (N_16495,N_15830,N_15941);
nand U16496 (N_16496,N_15503,N_15913);
nand U16497 (N_16497,N_15648,N_15954);
nand U16498 (N_16498,N_15587,N_15878);
nor U16499 (N_16499,N_15982,N_15670);
and U16500 (N_16500,N_16330,N_16224);
nor U16501 (N_16501,N_16312,N_16165);
xnor U16502 (N_16502,N_16447,N_16443);
or U16503 (N_16503,N_16218,N_16429);
or U16504 (N_16504,N_16132,N_16259);
or U16505 (N_16505,N_16261,N_16221);
nand U16506 (N_16506,N_16379,N_16463);
and U16507 (N_16507,N_16018,N_16207);
nand U16508 (N_16508,N_16237,N_16313);
and U16509 (N_16509,N_16410,N_16366);
xnor U16510 (N_16510,N_16394,N_16350);
and U16511 (N_16511,N_16436,N_16371);
nand U16512 (N_16512,N_16262,N_16135);
and U16513 (N_16513,N_16401,N_16299);
or U16514 (N_16514,N_16279,N_16157);
and U16515 (N_16515,N_16404,N_16288);
nand U16516 (N_16516,N_16470,N_16171);
and U16517 (N_16517,N_16308,N_16180);
xnor U16518 (N_16518,N_16417,N_16085);
nand U16519 (N_16519,N_16396,N_16214);
nor U16520 (N_16520,N_16021,N_16238);
xnor U16521 (N_16521,N_16307,N_16026);
xnor U16522 (N_16522,N_16211,N_16268);
and U16523 (N_16523,N_16163,N_16459);
or U16524 (N_16524,N_16141,N_16055);
and U16525 (N_16525,N_16113,N_16077);
and U16526 (N_16526,N_16497,N_16185);
and U16527 (N_16527,N_16204,N_16319);
xor U16528 (N_16528,N_16071,N_16027);
and U16529 (N_16529,N_16084,N_16206);
nor U16530 (N_16530,N_16452,N_16321);
nor U16531 (N_16531,N_16305,N_16413);
nor U16532 (N_16532,N_16037,N_16315);
or U16533 (N_16533,N_16317,N_16250);
or U16534 (N_16534,N_16166,N_16442);
and U16535 (N_16535,N_16161,N_16181);
nor U16536 (N_16536,N_16083,N_16493);
or U16537 (N_16537,N_16363,N_16300);
and U16538 (N_16538,N_16179,N_16193);
or U16539 (N_16539,N_16134,N_16292);
xnor U16540 (N_16540,N_16433,N_16223);
nor U16541 (N_16541,N_16107,N_16144);
xnor U16542 (N_16542,N_16205,N_16097);
or U16543 (N_16543,N_16040,N_16190);
nor U16544 (N_16544,N_16036,N_16395);
nand U16545 (N_16545,N_16428,N_16201);
or U16546 (N_16546,N_16286,N_16334);
nor U16547 (N_16547,N_16150,N_16478);
nor U16548 (N_16548,N_16124,N_16267);
or U16549 (N_16549,N_16147,N_16052);
nor U16550 (N_16550,N_16209,N_16473);
nand U16551 (N_16551,N_16331,N_16195);
nor U16552 (N_16552,N_16393,N_16160);
nor U16553 (N_16553,N_16121,N_16137);
or U16554 (N_16554,N_16381,N_16435);
or U16555 (N_16555,N_16047,N_16405);
nand U16556 (N_16556,N_16118,N_16215);
xor U16557 (N_16557,N_16082,N_16444);
or U16558 (N_16558,N_16353,N_16309);
nand U16559 (N_16559,N_16194,N_16189);
and U16560 (N_16560,N_16072,N_16153);
nand U16561 (N_16561,N_16461,N_16348);
and U16562 (N_16562,N_16336,N_16455);
or U16563 (N_16563,N_16271,N_16496);
and U16564 (N_16564,N_16380,N_16042);
and U16565 (N_16565,N_16054,N_16412);
nand U16566 (N_16566,N_16100,N_16246);
xnor U16567 (N_16567,N_16386,N_16297);
and U16568 (N_16568,N_16140,N_16407);
or U16569 (N_16569,N_16278,N_16074);
nor U16570 (N_16570,N_16420,N_16090);
or U16571 (N_16571,N_16337,N_16310);
and U16572 (N_16572,N_16034,N_16324);
nor U16573 (N_16573,N_16311,N_16041);
nor U16574 (N_16574,N_16392,N_16362);
nor U16575 (N_16575,N_16298,N_16007);
and U16576 (N_16576,N_16446,N_16170);
and U16577 (N_16577,N_16156,N_16199);
nand U16578 (N_16578,N_16266,N_16475);
nor U16579 (N_16579,N_16089,N_16116);
and U16580 (N_16580,N_16440,N_16245);
xor U16581 (N_16581,N_16338,N_16235);
and U16582 (N_16582,N_16468,N_16127);
and U16583 (N_16583,N_16495,N_16415);
or U16584 (N_16584,N_16432,N_16152);
nand U16585 (N_16585,N_16464,N_16354);
and U16586 (N_16586,N_16139,N_16075);
nor U16587 (N_16587,N_16051,N_16106);
xnor U16588 (N_16588,N_16225,N_16291);
xnor U16589 (N_16589,N_16372,N_16035);
or U16590 (N_16590,N_16110,N_16360);
or U16591 (N_16591,N_16426,N_16011);
xor U16592 (N_16592,N_16247,N_16332);
nand U16593 (N_16593,N_16466,N_16376);
nand U16594 (N_16594,N_16486,N_16439);
nand U16595 (N_16595,N_16364,N_16028);
xor U16596 (N_16596,N_16456,N_16397);
nand U16597 (N_16597,N_16492,N_16340);
nand U16598 (N_16598,N_16104,N_16057);
xor U16599 (N_16599,N_16458,N_16158);
nand U16600 (N_16600,N_16406,N_16045);
or U16601 (N_16601,N_16142,N_16399);
nand U16602 (N_16602,N_16065,N_16483);
and U16603 (N_16603,N_16389,N_16048);
and U16604 (N_16604,N_16341,N_16188);
or U16605 (N_16605,N_16285,N_16202);
or U16606 (N_16606,N_16320,N_16384);
xnor U16607 (N_16607,N_16129,N_16454);
nor U16608 (N_16608,N_16228,N_16236);
and U16609 (N_16609,N_16069,N_16343);
xor U16610 (N_16610,N_16377,N_16277);
or U16611 (N_16611,N_16010,N_16490);
xnor U16612 (N_16612,N_16025,N_16231);
nor U16613 (N_16613,N_16213,N_16098);
nand U16614 (N_16614,N_16164,N_16359);
and U16615 (N_16615,N_16438,N_16445);
and U16616 (N_16616,N_16070,N_16472);
and U16617 (N_16617,N_16280,N_16192);
nand U16618 (N_16618,N_16431,N_16176);
nand U16619 (N_16619,N_16451,N_16108);
or U16620 (N_16620,N_16066,N_16061);
or U16621 (N_16621,N_16208,N_16254);
and U16622 (N_16622,N_16203,N_16076);
nor U16623 (N_16623,N_16008,N_16091);
or U16624 (N_16624,N_16046,N_16339);
nand U16625 (N_16625,N_16109,N_16120);
and U16626 (N_16626,N_16335,N_16031);
or U16627 (N_16627,N_16293,N_16482);
xor U16628 (N_16628,N_16423,N_16378);
xnor U16629 (N_16629,N_16058,N_16481);
xnor U16630 (N_16630,N_16467,N_16004);
and U16631 (N_16631,N_16102,N_16159);
nor U16632 (N_16632,N_16414,N_16020);
xnor U16633 (N_16633,N_16284,N_16373);
nand U16634 (N_16634,N_16251,N_16032);
and U16635 (N_16635,N_16117,N_16002);
xor U16636 (N_16636,N_16361,N_16023);
or U16637 (N_16637,N_16487,N_16434);
xnor U16638 (N_16638,N_16453,N_16273);
nand U16639 (N_16639,N_16043,N_16148);
nor U16640 (N_16640,N_16287,N_16029);
xor U16641 (N_16641,N_16358,N_16220);
nand U16642 (N_16642,N_16145,N_16119);
xnor U16643 (N_16643,N_16197,N_16425);
and U16644 (N_16644,N_16351,N_16329);
nand U16645 (N_16645,N_16138,N_16243);
or U16646 (N_16646,N_16260,N_16347);
xor U16647 (N_16647,N_16123,N_16488);
nand U16648 (N_16648,N_16086,N_16143);
and U16649 (N_16649,N_16499,N_16050);
or U16650 (N_16650,N_16000,N_16095);
nand U16651 (N_16651,N_16187,N_16130);
xor U16652 (N_16652,N_16289,N_16128);
and U16653 (N_16653,N_16056,N_16400);
or U16654 (N_16654,N_16062,N_16263);
nor U16655 (N_16655,N_16151,N_16015);
nand U16656 (N_16656,N_16172,N_16274);
xor U16657 (N_16657,N_16244,N_16240);
nand U16658 (N_16658,N_16265,N_16409);
or U16659 (N_16659,N_16005,N_16112);
xnor U16660 (N_16660,N_16294,N_16154);
and U16661 (N_16661,N_16302,N_16345);
or U16662 (N_16662,N_16421,N_16013);
nor U16663 (N_16663,N_16126,N_16484);
or U16664 (N_16664,N_16096,N_16370);
xor U16665 (N_16665,N_16191,N_16198);
or U16666 (N_16666,N_16064,N_16184);
xor U16667 (N_16667,N_16101,N_16149);
nand U16668 (N_16668,N_16059,N_16030);
or U16669 (N_16669,N_16368,N_16441);
and U16670 (N_16670,N_16474,N_16078);
xnor U16671 (N_16671,N_16167,N_16038);
xor U16672 (N_16672,N_16326,N_16450);
nand U16673 (N_16673,N_16403,N_16318);
xnor U16674 (N_16674,N_16016,N_16009);
nand U16675 (N_16675,N_16460,N_16258);
and U16676 (N_16676,N_16080,N_16374);
or U16677 (N_16677,N_16014,N_16382);
xor U16678 (N_16678,N_16387,N_16408);
xor U16679 (N_16679,N_16178,N_16402);
nand U16680 (N_16680,N_16357,N_16019);
xnor U16681 (N_16681,N_16304,N_16063);
nand U16682 (N_16682,N_16398,N_16276);
nand U16683 (N_16683,N_16241,N_16416);
and U16684 (N_16684,N_16316,N_16115);
nor U16685 (N_16685,N_16003,N_16169);
or U16686 (N_16686,N_16437,N_16111);
and U16687 (N_16687,N_16448,N_16233);
or U16688 (N_16688,N_16323,N_16498);
and U16689 (N_16689,N_16039,N_16001);
nand U16690 (N_16690,N_16230,N_16314);
or U16691 (N_16691,N_16249,N_16229);
nand U16692 (N_16692,N_16333,N_16146);
nand U16693 (N_16693,N_16168,N_16248);
nor U16694 (N_16694,N_16099,N_16264);
and U16695 (N_16695,N_16491,N_16226);
nand U16696 (N_16696,N_16081,N_16346);
nand U16697 (N_16697,N_16217,N_16471);
and U16698 (N_16698,N_16175,N_16306);
xor U16699 (N_16699,N_16012,N_16232);
xor U16700 (N_16700,N_16212,N_16325);
and U16701 (N_16701,N_16196,N_16282);
or U16702 (N_16702,N_16272,N_16087);
xor U16703 (N_16703,N_16060,N_16256);
or U16704 (N_16704,N_16162,N_16275);
nand U16705 (N_16705,N_16131,N_16103);
nor U16706 (N_16706,N_16465,N_16369);
xnor U16707 (N_16707,N_16322,N_16344);
xnor U16708 (N_16708,N_16255,N_16219);
nand U16709 (N_16709,N_16479,N_16067);
or U16710 (N_16710,N_16480,N_16295);
xnor U16711 (N_16711,N_16173,N_16068);
xnor U16712 (N_16712,N_16186,N_16006);
or U16713 (N_16713,N_16281,N_16053);
or U16714 (N_16714,N_16270,N_16182);
xnor U16715 (N_16715,N_16352,N_16390);
or U16716 (N_16716,N_16494,N_16419);
nor U16717 (N_16717,N_16383,N_16411);
nand U16718 (N_16718,N_16355,N_16449);
nand U16719 (N_16719,N_16033,N_16327);
nor U16720 (N_16720,N_16462,N_16114);
nor U16721 (N_16721,N_16049,N_16155);
and U16722 (N_16722,N_16174,N_16093);
xnor U16723 (N_16723,N_16227,N_16257);
xnor U16724 (N_16724,N_16017,N_16125);
nor U16725 (N_16725,N_16457,N_16269);
xnor U16726 (N_16726,N_16301,N_16328);
and U16727 (N_16727,N_16122,N_16092);
nor U16728 (N_16728,N_16469,N_16356);
xor U16729 (N_16729,N_16427,N_16477);
and U16730 (N_16730,N_16476,N_16234);
and U16731 (N_16731,N_16216,N_16367);
or U16732 (N_16732,N_16430,N_16418);
or U16733 (N_16733,N_16422,N_16222);
and U16734 (N_16734,N_16088,N_16424);
and U16735 (N_16735,N_16210,N_16044);
and U16736 (N_16736,N_16094,N_16375);
xor U16737 (N_16737,N_16385,N_16200);
xor U16738 (N_16738,N_16391,N_16133);
and U16739 (N_16739,N_16485,N_16105);
xnor U16740 (N_16740,N_16024,N_16136);
nand U16741 (N_16741,N_16079,N_16296);
nand U16742 (N_16742,N_16253,N_16365);
nand U16743 (N_16743,N_16388,N_16183);
and U16744 (N_16744,N_16290,N_16239);
nor U16745 (N_16745,N_16342,N_16489);
nand U16746 (N_16746,N_16252,N_16303);
nand U16747 (N_16747,N_16283,N_16073);
and U16748 (N_16748,N_16349,N_16242);
and U16749 (N_16749,N_16177,N_16022);
xor U16750 (N_16750,N_16496,N_16079);
nand U16751 (N_16751,N_16012,N_16160);
and U16752 (N_16752,N_16361,N_16365);
or U16753 (N_16753,N_16185,N_16238);
and U16754 (N_16754,N_16131,N_16353);
nand U16755 (N_16755,N_16082,N_16073);
and U16756 (N_16756,N_16352,N_16199);
nor U16757 (N_16757,N_16122,N_16066);
nand U16758 (N_16758,N_16057,N_16097);
or U16759 (N_16759,N_16429,N_16372);
or U16760 (N_16760,N_16391,N_16044);
or U16761 (N_16761,N_16445,N_16161);
nand U16762 (N_16762,N_16284,N_16041);
nand U16763 (N_16763,N_16206,N_16481);
or U16764 (N_16764,N_16455,N_16267);
or U16765 (N_16765,N_16057,N_16368);
and U16766 (N_16766,N_16388,N_16235);
nor U16767 (N_16767,N_16114,N_16116);
nor U16768 (N_16768,N_16034,N_16065);
or U16769 (N_16769,N_16187,N_16373);
xor U16770 (N_16770,N_16306,N_16192);
or U16771 (N_16771,N_16275,N_16007);
nor U16772 (N_16772,N_16190,N_16472);
xnor U16773 (N_16773,N_16163,N_16064);
nand U16774 (N_16774,N_16404,N_16422);
nor U16775 (N_16775,N_16027,N_16100);
xnor U16776 (N_16776,N_16380,N_16023);
nand U16777 (N_16777,N_16176,N_16177);
nand U16778 (N_16778,N_16059,N_16480);
nand U16779 (N_16779,N_16017,N_16012);
and U16780 (N_16780,N_16495,N_16358);
nor U16781 (N_16781,N_16403,N_16136);
or U16782 (N_16782,N_16286,N_16232);
or U16783 (N_16783,N_16101,N_16216);
or U16784 (N_16784,N_16117,N_16021);
nand U16785 (N_16785,N_16064,N_16368);
xor U16786 (N_16786,N_16027,N_16009);
xnor U16787 (N_16787,N_16075,N_16040);
xor U16788 (N_16788,N_16477,N_16032);
xor U16789 (N_16789,N_16499,N_16269);
or U16790 (N_16790,N_16161,N_16372);
and U16791 (N_16791,N_16216,N_16349);
xor U16792 (N_16792,N_16245,N_16115);
nand U16793 (N_16793,N_16139,N_16042);
nor U16794 (N_16794,N_16334,N_16203);
xnor U16795 (N_16795,N_16490,N_16015);
or U16796 (N_16796,N_16486,N_16272);
and U16797 (N_16797,N_16480,N_16429);
and U16798 (N_16798,N_16120,N_16490);
nor U16799 (N_16799,N_16462,N_16337);
and U16800 (N_16800,N_16295,N_16017);
nor U16801 (N_16801,N_16026,N_16334);
xnor U16802 (N_16802,N_16099,N_16003);
nor U16803 (N_16803,N_16380,N_16407);
xnor U16804 (N_16804,N_16113,N_16244);
or U16805 (N_16805,N_16281,N_16324);
or U16806 (N_16806,N_16447,N_16236);
nor U16807 (N_16807,N_16212,N_16290);
and U16808 (N_16808,N_16094,N_16416);
or U16809 (N_16809,N_16186,N_16079);
or U16810 (N_16810,N_16093,N_16133);
or U16811 (N_16811,N_16323,N_16442);
or U16812 (N_16812,N_16149,N_16400);
and U16813 (N_16813,N_16463,N_16142);
nor U16814 (N_16814,N_16462,N_16049);
or U16815 (N_16815,N_16054,N_16208);
or U16816 (N_16816,N_16152,N_16297);
or U16817 (N_16817,N_16285,N_16379);
or U16818 (N_16818,N_16133,N_16059);
and U16819 (N_16819,N_16122,N_16478);
nor U16820 (N_16820,N_16483,N_16309);
nand U16821 (N_16821,N_16243,N_16069);
or U16822 (N_16822,N_16362,N_16343);
nand U16823 (N_16823,N_16405,N_16196);
nand U16824 (N_16824,N_16217,N_16265);
xor U16825 (N_16825,N_16098,N_16379);
and U16826 (N_16826,N_16421,N_16424);
nand U16827 (N_16827,N_16234,N_16492);
nor U16828 (N_16828,N_16408,N_16012);
nor U16829 (N_16829,N_16019,N_16250);
nand U16830 (N_16830,N_16498,N_16274);
nor U16831 (N_16831,N_16309,N_16316);
and U16832 (N_16832,N_16070,N_16308);
nor U16833 (N_16833,N_16496,N_16082);
nand U16834 (N_16834,N_16041,N_16038);
nand U16835 (N_16835,N_16352,N_16235);
and U16836 (N_16836,N_16043,N_16149);
or U16837 (N_16837,N_16405,N_16426);
xnor U16838 (N_16838,N_16037,N_16138);
and U16839 (N_16839,N_16127,N_16156);
and U16840 (N_16840,N_16386,N_16155);
xnor U16841 (N_16841,N_16279,N_16397);
nor U16842 (N_16842,N_16147,N_16323);
xnor U16843 (N_16843,N_16065,N_16491);
nand U16844 (N_16844,N_16414,N_16434);
nand U16845 (N_16845,N_16437,N_16361);
xnor U16846 (N_16846,N_16220,N_16170);
and U16847 (N_16847,N_16218,N_16084);
and U16848 (N_16848,N_16427,N_16016);
xnor U16849 (N_16849,N_16143,N_16437);
or U16850 (N_16850,N_16093,N_16194);
nor U16851 (N_16851,N_16043,N_16237);
xnor U16852 (N_16852,N_16427,N_16295);
xor U16853 (N_16853,N_16085,N_16390);
nor U16854 (N_16854,N_16229,N_16071);
nand U16855 (N_16855,N_16150,N_16197);
and U16856 (N_16856,N_16448,N_16122);
nor U16857 (N_16857,N_16035,N_16290);
or U16858 (N_16858,N_16326,N_16019);
nor U16859 (N_16859,N_16312,N_16132);
and U16860 (N_16860,N_16296,N_16364);
or U16861 (N_16861,N_16202,N_16013);
and U16862 (N_16862,N_16455,N_16206);
xnor U16863 (N_16863,N_16105,N_16405);
xor U16864 (N_16864,N_16084,N_16192);
xor U16865 (N_16865,N_16058,N_16222);
xor U16866 (N_16866,N_16431,N_16499);
xnor U16867 (N_16867,N_16408,N_16482);
nor U16868 (N_16868,N_16141,N_16309);
and U16869 (N_16869,N_16021,N_16114);
nor U16870 (N_16870,N_16365,N_16250);
xor U16871 (N_16871,N_16015,N_16014);
and U16872 (N_16872,N_16120,N_16421);
or U16873 (N_16873,N_16192,N_16307);
or U16874 (N_16874,N_16322,N_16309);
nand U16875 (N_16875,N_16425,N_16293);
or U16876 (N_16876,N_16208,N_16474);
nand U16877 (N_16877,N_16458,N_16180);
nor U16878 (N_16878,N_16465,N_16161);
nand U16879 (N_16879,N_16136,N_16040);
nor U16880 (N_16880,N_16379,N_16091);
or U16881 (N_16881,N_16467,N_16223);
nand U16882 (N_16882,N_16190,N_16113);
or U16883 (N_16883,N_16070,N_16384);
or U16884 (N_16884,N_16036,N_16142);
nor U16885 (N_16885,N_16229,N_16292);
nor U16886 (N_16886,N_16079,N_16280);
nand U16887 (N_16887,N_16232,N_16037);
or U16888 (N_16888,N_16452,N_16431);
or U16889 (N_16889,N_16306,N_16207);
xnor U16890 (N_16890,N_16185,N_16496);
nor U16891 (N_16891,N_16466,N_16087);
and U16892 (N_16892,N_16188,N_16374);
nand U16893 (N_16893,N_16285,N_16480);
nand U16894 (N_16894,N_16109,N_16175);
nor U16895 (N_16895,N_16407,N_16233);
nor U16896 (N_16896,N_16134,N_16024);
nor U16897 (N_16897,N_16014,N_16225);
nand U16898 (N_16898,N_16384,N_16482);
and U16899 (N_16899,N_16398,N_16150);
nor U16900 (N_16900,N_16150,N_16469);
and U16901 (N_16901,N_16025,N_16118);
xnor U16902 (N_16902,N_16464,N_16103);
nand U16903 (N_16903,N_16128,N_16304);
and U16904 (N_16904,N_16249,N_16007);
xnor U16905 (N_16905,N_16192,N_16423);
or U16906 (N_16906,N_16118,N_16122);
nor U16907 (N_16907,N_16065,N_16082);
or U16908 (N_16908,N_16121,N_16132);
or U16909 (N_16909,N_16487,N_16282);
xor U16910 (N_16910,N_16004,N_16474);
and U16911 (N_16911,N_16179,N_16229);
or U16912 (N_16912,N_16493,N_16482);
nand U16913 (N_16913,N_16499,N_16331);
nand U16914 (N_16914,N_16349,N_16168);
or U16915 (N_16915,N_16079,N_16461);
and U16916 (N_16916,N_16080,N_16011);
nor U16917 (N_16917,N_16321,N_16499);
nor U16918 (N_16918,N_16320,N_16419);
xor U16919 (N_16919,N_16407,N_16045);
nand U16920 (N_16920,N_16408,N_16010);
xor U16921 (N_16921,N_16342,N_16375);
xnor U16922 (N_16922,N_16225,N_16100);
or U16923 (N_16923,N_16101,N_16355);
or U16924 (N_16924,N_16075,N_16499);
and U16925 (N_16925,N_16224,N_16077);
or U16926 (N_16926,N_16288,N_16353);
nand U16927 (N_16927,N_16327,N_16437);
nor U16928 (N_16928,N_16492,N_16384);
and U16929 (N_16929,N_16373,N_16226);
or U16930 (N_16930,N_16219,N_16455);
and U16931 (N_16931,N_16181,N_16173);
and U16932 (N_16932,N_16319,N_16419);
xor U16933 (N_16933,N_16454,N_16406);
xnor U16934 (N_16934,N_16005,N_16343);
nand U16935 (N_16935,N_16203,N_16312);
and U16936 (N_16936,N_16392,N_16248);
xnor U16937 (N_16937,N_16499,N_16042);
nor U16938 (N_16938,N_16074,N_16428);
nand U16939 (N_16939,N_16016,N_16230);
or U16940 (N_16940,N_16397,N_16399);
and U16941 (N_16941,N_16462,N_16155);
or U16942 (N_16942,N_16086,N_16091);
and U16943 (N_16943,N_16026,N_16433);
xnor U16944 (N_16944,N_16227,N_16022);
and U16945 (N_16945,N_16410,N_16015);
or U16946 (N_16946,N_16194,N_16264);
nand U16947 (N_16947,N_16172,N_16231);
xor U16948 (N_16948,N_16128,N_16071);
or U16949 (N_16949,N_16311,N_16222);
and U16950 (N_16950,N_16362,N_16425);
xnor U16951 (N_16951,N_16380,N_16345);
and U16952 (N_16952,N_16040,N_16294);
xor U16953 (N_16953,N_16246,N_16460);
or U16954 (N_16954,N_16161,N_16368);
nor U16955 (N_16955,N_16369,N_16082);
and U16956 (N_16956,N_16305,N_16175);
nor U16957 (N_16957,N_16439,N_16421);
and U16958 (N_16958,N_16301,N_16096);
xor U16959 (N_16959,N_16321,N_16268);
and U16960 (N_16960,N_16056,N_16195);
nor U16961 (N_16961,N_16400,N_16052);
xnor U16962 (N_16962,N_16275,N_16448);
nand U16963 (N_16963,N_16449,N_16335);
or U16964 (N_16964,N_16141,N_16325);
nor U16965 (N_16965,N_16063,N_16035);
xnor U16966 (N_16966,N_16253,N_16383);
or U16967 (N_16967,N_16371,N_16307);
xnor U16968 (N_16968,N_16317,N_16050);
xor U16969 (N_16969,N_16362,N_16255);
or U16970 (N_16970,N_16100,N_16402);
nand U16971 (N_16971,N_16088,N_16224);
nor U16972 (N_16972,N_16033,N_16278);
or U16973 (N_16973,N_16324,N_16388);
xor U16974 (N_16974,N_16228,N_16051);
xor U16975 (N_16975,N_16268,N_16040);
nand U16976 (N_16976,N_16497,N_16268);
nor U16977 (N_16977,N_16077,N_16425);
and U16978 (N_16978,N_16441,N_16444);
nor U16979 (N_16979,N_16244,N_16159);
nor U16980 (N_16980,N_16063,N_16199);
and U16981 (N_16981,N_16376,N_16250);
or U16982 (N_16982,N_16044,N_16087);
and U16983 (N_16983,N_16067,N_16074);
nor U16984 (N_16984,N_16416,N_16332);
and U16985 (N_16985,N_16494,N_16036);
nor U16986 (N_16986,N_16482,N_16188);
and U16987 (N_16987,N_16262,N_16218);
or U16988 (N_16988,N_16219,N_16056);
nor U16989 (N_16989,N_16143,N_16093);
xnor U16990 (N_16990,N_16452,N_16323);
or U16991 (N_16991,N_16020,N_16134);
or U16992 (N_16992,N_16092,N_16158);
xnor U16993 (N_16993,N_16378,N_16343);
nor U16994 (N_16994,N_16253,N_16348);
or U16995 (N_16995,N_16374,N_16021);
nor U16996 (N_16996,N_16362,N_16337);
xor U16997 (N_16997,N_16029,N_16272);
and U16998 (N_16998,N_16128,N_16397);
nor U16999 (N_16999,N_16054,N_16342);
or U17000 (N_17000,N_16948,N_16995);
or U17001 (N_17001,N_16856,N_16775);
xor U17002 (N_17002,N_16745,N_16711);
nor U17003 (N_17003,N_16931,N_16639);
nand U17004 (N_17004,N_16878,N_16684);
nor U17005 (N_17005,N_16875,N_16696);
and U17006 (N_17006,N_16730,N_16968);
or U17007 (N_17007,N_16516,N_16713);
xnor U17008 (N_17008,N_16520,N_16561);
xor U17009 (N_17009,N_16946,N_16603);
or U17010 (N_17010,N_16848,N_16902);
or U17011 (N_17011,N_16820,N_16951);
or U17012 (N_17012,N_16537,N_16832);
nand U17013 (N_17013,N_16814,N_16911);
nand U17014 (N_17014,N_16766,N_16927);
nand U17015 (N_17015,N_16750,N_16892);
nand U17016 (N_17016,N_16538,N_16607);
or U17017 (N_17017,N_16563,N_16886);
nor U17018 (N_17018,N_16862,N_16715);
nor U17019 (N_17019,N_16536,N_16959);
nand U17020 (N_17020,N_16816,N_16854);
nand U17021 (N_17021,N_16828,N_16544);
or U17022 (N_17022,N_16768,N_16870);
and U17023 (N_17023,N_16518,N_16799);
or U17024 (N_17024,N_16650,N_16920);
nand U17025 (N_17025,N_16867,N_16542);
nand U17026 (N_17026,N_16926,N_16749);
xnor U17027 (N_17027,N_16534,N_16971);
nor U17028 (N_17028,N_16779,N_16554);
xor U17029 (N_17029,N_16859,N_16758);
nand U17030 (N_17030,N_16569,N_16671);
nor U17031 (N_17031,N_16982,N_16769);
or U17032 (N_17032,N_16611,N_16527);
nand U17033 (N_17033,N_16793,N_16823);
and U17034 (N_17034,N_16930,N_16756);
nor U17035 (N_17035,N_16928,N_16559);
nor U17036 (N_17036,N_16541,N_16897);
and U17037 (N_17037,N_16863,N_16784);
and U17038 (N_17038,N_16853,N_16903);
nand U17039 (N_17039,N_16701,N_16526);
and U17040 (N_17040,N_16890,N_16906);
and U17041 (N_17041,N_16532,N_16663);
and U17042 (N_17042,N_16824,N_16629);
and U17043 (N_17043,N_16970,N_16618);
and U17044 (N_17044,N_16535,N_16914);
nor U17045 (N_17045,N_16725,N_16619);
and U17046 (N_17046,N_16633,N_16679);
xnor U17047 (N_17047,N_16746,N_16547);
or U17048 (N_17048,N_16644,N_16916);
nand U17049 (N_17049,N_16702,N_16934);
xor U17050 (N_17050,N_16879,N_16693);
xor U17051 (N_17051,N_16630,N_16700);
nor U17052 (N_17052,N_16785,N_16637);
or U17053 (N_17053,N_16924,N_16577);
nand U17054 (N_17054,N_16695,N_16558);
and U17055 (N_17055,N_16628,N_16839);
nand U17056 (N_17056,N_16626,N_16591);
nand U17057 (N_17057,N_16501,N_16682);
xor U17058 (N_17058,N_16643,N_16901);
and U17059 (N_17059,N_16899,N_16976);
nand U17060 (N_17060,N_16675,N_16732);
nand U17061 (N_17061,N_16590,N_16877);
nor U17062 (N_17062,N_16938,N_16571);
and U17063 (N_17063,N_16737,N_16865);
nor U17064 (N_17064,N_16575,N_16551);
nand U17065 (N_17065,N_16767,N_16837);
nor U17066 (N_17066,N_16985,N_16858);
or U17067 (N_17067,N_16815,N_16937);
or U17068 (N_17068,N_16963,N_16964);
or U17069 (N_17069,N_16909,N_16808);
nand U17070 (N_17070,N_16720,N_16581);
nand U17071 (N_17071,N_16776,N_16600);
nor U17072 (N_17072,N_16900,N_16507);
and U17073 (N_17073,N_16975,N_16578);
nor U17074 (N_17074,N_16705,N_16810);
nor U17075 (N_17075,N_16855,N_16835);
and U17076 (N_17076,N_16990,N_16989);
nor U17077 (N_17077,N_16557,N_16662);
and U17078 (N_17078,N_16893,N_16599);
xnor U17079 (N_17079,N_16685,N_16586);
nor U17080 (N_17080,N_16743,N_16807);
nor U17081 (N_17081,N_16850,N_16648);
or U17082 (N_17082,N_16716,N_16864);
xnor U17083 (N_17083,N_16589,N_16957);
or U17084 (N_17084,N_16809,N_16986);
and U17085 (N_17085,N_16838,N_16840);
or U17086 (N_17086,N_16714,N_16861);
and U17087 (N_17087,N_16584,N_16651);
nand U17088 (N_17088,N_16821,N_16510);
xnor U17089 (N_17089,N_16585,N_16764);
xor U17090 (N_17090,N_16781,N_16513);
and U17091 (N_17091,N_16625,N_16770);
or U17092 (N_17092,N_16795,N_16978);
and U17093 (N_17093,N_16640,N_16887);
nor U17094 (N_17094,N_16717,N_16983);
nand U17095 (N_17095,N_16883,N_16772);
or U17096 (N_17096,N_16522,N_16655);
nand U17097 (N_17097,N_16857,N_16981);
and U17098 (N_17098,N_16760,N_16956);
xnor U17099 (N_17099,N_16594,N_16895);
nor U17100 (N_17100,N_16907,N_16545);
nor U17101 (N_17101,N_16869,N_16852);
and U17102 (N_17102,N_16804,N_16881);
or U17103 (N_17103,N_16708,N_16866);
or U17104 (N_17104,N_16605,N_16933);
or U17105 (N_17105,N_16778,N_16974);
nor U17106 (N_17106,N_16872,N_16952);
or U17107 (N_17107,N_16574,N_16919);
nand U17108 (N_17108,N_16972,N_16996);
or U17109 (N_17109,N_16632,N_16777);
nor U17110 (N_17110,N_16517,N_16562);
nand U17111 (N_17111,N_16979,N_16898);
xor U17112 (N_17112,N_16514,N_16741);
or U17113 (N_17113,N_16598,N_16761);
nor U17114 (N_17114,N_16642,N_16706);
nor U17115 (N_17115,N_16548,N_16967);
and U17116 (N_17116,N_16800,N_16722);
or U17117 (N_17117,N_16842,N_16621);
or U17118 (N_17118,N_16595,N_16659);
or U17119 (N_17119,N_16553,N_16891);
and U17120 (N_17120,N_16845,N_16780);
or U17121 (N_17121,N_16641,N_16576);
nor U17122 (N_17122,N_16885,N_16836);
and U17123 (N_17123,N_16936,N_16593);
xnor U17124 (N_17124,N_16546,N_16733);
nor U17125 (N_17125,N_16790,N_16588);
or U17126 (N_17126,N_16921,N_16677);
or U17127 (N_17127,N_16834,N_16751);
nor U17128 (N_17128,N_16515,N_16612);
xnor U17129 (N_17129,N_16698,N_16549);
and U17130 (N_17130,N_16673,N_16688);
nor U17131 (N_17131,N_16792,N_16676);
and U17132 (N_17132,N_16529,N_16923);
nand U17133 (N_17133,N_16998,N_16992);
xnor U17134 (N_17134,N_16694,N_16843);
nand U17135 (N_17135,N_16521,N_16844);
and U17136 (N_17136,N_16721,N_16740);
xor U17137 (N_17137,N_16500,N_16680);
and U17138 (N_17138,N_16939,N_16560);
nor U17139 (N_17139,N_16503,N_16656);
xor U17140 (N_17140,N_16782,N_16699);
xor U17141 (N_17141,N_16638,N_16580);
xor U17142 (N_17142,N_16945,N_16731);
and U17143 (N_17143,N_16666,N_16606);
nor U17144 (N_17144,N_16596,N_16966);
and U17145 (N_17145,N_16724,N_16674);
xnor U17146 (N_17146,N_16565,N_16791);
and U17147 (N_17147,N_16918,N_16636);
nor U17148 (N_17148,N_16997,N_16524);
nand U17149 (N_17149,N_16627,N_16817);
and U17150 (N_17150,N_16623,N_16718);
nand U17151 (N_17151,N_16602,N_16660);
nand U17152 (N_17152,N_16787,N_16880);
nand U17153 (N_17153,N_16753,N_16683);
or U17154 (N_17154,N_16509,N_16819);
nand U17155 (N_17155,N_16794,N_16757);
xnor U17156 (N_17156,N_16830,N_16811);
and U17157 (N_17157,N_16646,N_16691);
and U17158 (N_17158,N_16601,N_16922);
and U17159 (N_17159,N_16786,N_16993);
or U17160 (N_17160,N_16678,N_16960);
nand U17161 (N_17161,N_16727,N_16752);
xnor U17162 (N_17162,N_16729,N_16613);
nor U17163 (N_17163,N_16940,N_16788);
nor U17164 (N_17164,N_16973,N_16954);
nor U17165 (N_17165,N_16658,N_16797);
nor U17166 (N_17166,N_16999,N_16635);
nor U17167 (N_17167,N_16672,N_16894);
nor U17168 (N_17168,N_16723,N_16681);
nor U17169 (N_17169,N_16943,N_16592);
or U17170 (N_17170,N_16742,N_16915);
or U17171 (N_17171,N_16765,N_16994);
or U17172 (N_17172,N_16813,N_16735);
nand U17173 (N_17173,N_16616,N_16849);
xor U17174 (N_17174,N_16991,N_16645);
xnor U17175 (N_17175,N_16944,N_16738);
nand U17176 (N_17176,N_16608,N_16667);
nand U17177 (N_17177,N_16689,N_16803);
nor U17178 (N_17178,N_16739,N_16617);
nor U17179 (N_17179,N_16508,N_16904);
nand U17180 (N_17180,N_16736,N_16818);
and U17181 (N_17181,N_16533,N_16615);
and U17182 (N_17182,N_16851,N_16917);
nand U17183 (N_17183,N_16614,N_16707);
nor U17184 (N_17184,N_16932,N_16876);
nor U17185 (N_17185,N_16969,N_16759);
and U17186 (N_17186,N_16796,N_16846);
xnor U17187 (N_17187,N_16913,N_16528);
nor U17188 (N_17188,N_16747,N_16668);
nand U17189 (N_17189,N_16512,N_16774);
xnor U17190 (N_17190,N_16942,N_16582);
or U17191 (N_17191,N_16669,N_16511);
nor U17192 (N_17192,N_16910,N_16665);
or U17193 (N_17193,N_16609,N_16831);
xnor U17194 (N_17194,N_16755,N_16988);
or U17195 (N_17195,N_16543,N_16540);
nand U17196 (N_17196,N_16556,N_16812);
and U17197 (N_17197,N_16525,N_16965);
nor U17198 (N_17198,N_16710,N_16825);
xor U17199 (N_17199,N_16962,N_16888);
xnor U17200 (N_17200,N_16947,N_16805);
nand U17201 (N_17201,N_16806,N_16798);
or U17202 (N_17202,N_16868,N_16649);
nand U17203 (N_17203,N_16977,N_16847);
and U17204 (N_17204,N_16692,N_16624);
xor U17205 (N_17205,N_16670,N_16652);
xnor U17206 (N_17206,N_16896,N_16955);
nand U17207 (N_17207,N_16925,N_16726);
xor U17208 (N_17208,N_16773,N_16568);
nor U17209 (N_17209,N_16734,N_16929);
xnor U17210 (N_17210,N_16712,N_16506);
nand U17211 (N_17211,N_16826,N_16827);
nor U17212 (N_17212,N_16555,N_16748);
xnor U17213 (N_17213,N_16610,N_16664);
or U17214 (N_17214,N_16935,N_16871);
or U17215 (N_17215,N_16572,N_16687);
or U17216 (N_17216,N_16860,N_16530);
or U17217 (N_17217,N_16941,N_16884);
and U17218 (N_17218,N_16523,N_16690);
nor U17219 (N_17219,N_16874,N_16502);
xnor U17220 (N_17220,N_16573,N_16802);
and U17221 (N_17221,N_16719,N_16703);
xnor U17222 (N_17222,N_16873,N_16587);
or U17223 (N_17223,N_16882,N_16833);
or U17224 (N_17224,N_16709,N_16958);
and U17225 (N_17225,N_16519,N_16984);
or U17226 (N_17226,N_16539,N_16531);
nor U17227 (N_17227,N_16980,N_16550);
xor U17228 (N_17228,N_16552,N_16889);
nor U17229 (N_17229,N_16829,N_16704);
nand U17230 (N_17230,N_16771,N_16505);
or U17231 (N_17231,N_16597,N_16950);
and U17232 (N_17232,N_16686,N_16661);
and U17233 (N_17233,N_16841,N_16579);
xor U17234 (N_17234,N_16567,N_16504);
and U17235 (N_17235,N_16647,N_16622);
xnor U17236 (N_17236,N_16654,N_16789);
or U17237 (N_17237,N_16570,N_16566);
xor U17238 (N_17238,N_16631,N_16754);
xor U17239 (N_17239,N_16728,N_16653);
and U17240 (N_17240,N_16912,N_16564);
xnor U17241 (N_17241,N_16783,N_16905);
nor U17242 (N_17242,N_16987,N_16949);
nand U17243 (N_17243,N_16583,N_16762);
xnor U17244 (N_17244,N_16822,N_16604);
nor U17245 (N_17245,N_16744,N_16620);
and U17246 (N_17246,N_16953,N_16908);
or U17247 (N_17247,N_16634,N_16801);
nor U17248 (N_17248,N_16697,N_16657);
or U17249 (N_17249,N_16961,N_16763);
nor U17250 (N_17250,N_16875,N_16609);
nor U17251 (N_17251,N_16956,N_16518);
and U17252 (N_17252,N_16622,N_16635);
and U17253 (N_17253,N_16609,N_16667);
nand U17254 (N_17254,N_16940,N_16995);
xor U17255 (N_17255,N_16581,N_16729);
or U17256 (N_17256,N_16588,N_16860);
xnor U17257 (N_17257,N_16958,N_16614);
and U17258 (N_17258,N_16894,N_16962);
or U17259 (N_17259,N_16930,N_16598);
nand U17260 (N_17260,N_16621,N_16973);
nand U17261 (N_17261,N_16793,N_16653);
and U17262 (N_17262,N_16622,N_16517);
xnor U17263 (N_17263,N_16525,N_16810);
nor U17264 (N_17264,N_16604,N_16706);
and U17265 (N_17265,N_16535,N_16617);
or U17266 (N_17266,N_16696,N_16606);
nand U17267 (N_17267,N_16714,N_16767);
and U17268 (N_17268,N_16558,N_16914);
or U17269 (N_17269,N_16852,N_16885);
xnor U17270 (N_17270,N_16509,N_16633);
nand U17271 (N_17271,N_16926,N_16553);
and U17272 (N_17272,N_16858,N_16838);
nand U17273 (N_17273,N_16920,N_16876);
and U17274 (N_17274,N_16665,N_16707);
nand U17275 (N_17275,N_16985,N_16592);
nand U17276 (N_17276,N_16618,N_16735);
and U17277 (N_17277,N_16793,N_16943);
xnor U17278 (N_17278,N_16709,N_16715);
and U17279 (N_17279,N_16586,N_16508);
or U17280 (N_17280,N_16985,N_16827);
nand U17281 (N_17281,N_16990,N_16733);
nand U17282 (N_17282,N_16610,N_16724);
or U17283 (N_17283,N_16506,N_16876);
xnor U17284 (N_17284,N_16602,N_16688);
nand U17285 (N_17285,N_16995,N_16652);
xnor U17286 (N_17286,N_16997,N_16749);
or U17287 (N_17287,N_16663,N_16879);
nand U17288 (N_17288,N_16848,N_16941);
and U17289 (N_17289,N_16895,N_16519);
or U17290 (N_17290,N_16783,N_16578);
nor U17291 (N_17291,N_16933,N_16939);
and U17292 (N_17292,N_16586,N_16803);
xor U17293 (N_17293,N_16532,N_16826);
or U17294 (N_17294,N_16835,N_16520);
nor U17295 (N_17295,N_16590,N_16629);
nand U17296 (N_17296,N_16715,N_16808);
nand U17297 (N_17297,N_16982,N_16944);
nor U17298 (N_17298,N_16733,N_16538);
nor U17299 (N_17299,N_16832,N_16701);
or U17300 (N_17300,N_16661,N_16570);
or U17301 (N_17301,N_16507,N_16776);
nand U17302 (N_17302,N_16835,N_16930);
and U17303 (N_17303,N_16857,N_16556);
or U17304 (N_17304,N_16744,N_16962);
xor U17305 (N_17305,N_16542,N_16933);
nor U17306 (N_17306,N_16515,N_16745);
or U17307 (N_17307,N_16804,N_16890);
and U17308 (N_17308,N_16509,N_16702);
nor U17309 (N_17309,N_16916,N_16692);
or U17310 (N_17310,N_16708,N_16542);
nand U17311 (N_17311,N_16643,N_16850);
and U17312 (N_17312,N_16706,N_16745);
or U17313 (N_17313,N_16530,N_16871);
nor U17314 (N_17314,N_16650,N_16570);
nor U17315 (N_17315,N_16720,N_16516);
nor U17316 (N_17316,N_16893,N_16973);
and U17317 (N_17317,N_16632,N_16827);
and U17318 (N_17318,N_16552,N_16697);
nand U17319 (N_17319,N_16934,N_16946);
nor U17320 (N_17320,N_16571,N_16612);
and U17321 (N_17321,N_16888,N_16844);
or U17322 (N_17322,N_16922,N_16749);
xnor U17323 (N_17323,N_16900,N_16511);
and U17324 (N_17324,N_16536,N_16794);
xor U17325 (N_17325,N_16502,N_16511);
xor U17326 (N_17326,N_16505,N_16960);
and U17327 (N_17327,N_16648,N_16873);
nand U17328 (N_17328,N_16896,N_16608);
or U17329 (N_17329,N_16871,N_16689);
nand U17330 (N_17330,N_16979,N_16608);
xnor U17331 (N_17331,N_16714,N_16642);
nor U17332 (N_17332,N_16959,N_16730);
xor U17333 (N_17333,N_16652,N_16924);
nand U17334 (N_17334,N_16571,N_16860);
or U17335 (N_17335,N_16951,N_16783);
or U17336 (N_17336,N_16628,N_16640);
or U17337 (N_17337,N_16726,N_16685);
or U17338 (N_17338,N_16692,N_16569);
xor U17339 (N_17339,N_16807,N_16574);
or U17340 (N_17340,N_16586,N_16876);
xor U17341 (N_17341,N_16785,N_16854);
xnor U17342 (N_17342,N_16791,N_16903);
and U17343 (N_17343,N_16816,N_16728);
xnor U17344 (N_17344,N_16946,N_16895);
and U17345 (N_17345,N_16962,N_16646);
xor U17346 (N_17346,N_16950,N_16664);
xnor U17347 (N_17347,N_16748,N_16585);
xnor U17348 (N_17348,N_16595,N_16843);
xnor U17349 (N_17349,N_16600,N_16591);
or U17350 (N_17350,N_16639,N_16759);
or U17351 (N_17351,N_16908,N_16867);
and U17352 (N_17352,N_16956,N_16830);
or U17353 (N_17353,N_16862,N_16900);
xor U17354 (N_17354,N_16994,N_16851);
xnor U17355 (N_17355,N_16952,N_16715);
and U17356 (N_17356,N_16539,N_16728);
xor U17357 (N_17357,N_16785,N_16660);
nand U17358 (N_17358,N_16846,N_16889);
nor U17359 (N_17359,N_16622,N_16808);
nand U17360 (N_17360,N_16507,N_16606);
and U17361 (N_17361,N_16908,N_16617);
and U17362 (N_17362,N_16669,N_16780);
nand U17363 (N_17363,N_16659,N_16809);
nor U17364 (N_17364,N_16533,N_16850);
nor U17365 (N_17365,N_16520,N_16687);
or U17366 (N_17366,N_16679,N_16939);
xor U17367 (N_17367,N_16857,N_16520);
nand U17368 (N_17368,N_16622,N_16907);
xor U17369 (N_17369,N_16715,N_16990);
and U17370 (N_17370,N_16975,N_16679);
and U17371 (N_17371,N_16538,N_16876);
and U17372 (N_17372,N_16979,N_16578);
nand U17373 (N_17373,N_16675,N_16751);
xor U17374 (N_17374,N_16899,N_16707);
nand U17375 (N_17375,N_16833,N_16605);
or U17376 (N_17376,N_16821,N_16818);
and U17377 (N_17377,N_16787,N_16548);
xnor U17378 (N_17378,N_16540,N_16858);
and U17379 (N_17379,N_16921,N_16615);
nand U17380 (N_17380,N_16679,N_16621);
nor U17381 (N_17381,N_16620,N_16555);
nand U17382 (N_17382,N_16909,N_16712);
nand U17383 (N_17383,N_16503,N_16960);
or U17384 (N_17384,N_16556,N_16982);
xnor U17385 (N_17385,N_16985,N_16502);
xnor U17386 (N_17386,N_16563,N_16552);
nor U17387 (N_17387,N_16568,N_16618);
and U17388 (N_17388,N_16828,N_16926);
or U17389 (N_17389,N_16973,N_16589);
nor U17390 (N_17390,N_16670,N_16669);
and U17391 (N_17391,N_16732,N_16796);
nand U17392 (N_17392,N_16625,N_16531);
xor U17393 (N_17393,N_16995,N_16737);
xor U17394 (N_17394,N_16971,N_16850);
or U17395 (N_17395,N_16947,N_16602);
xor U17396 (N_17396,N_16593,N_16839);
nand U17397 (N_17397,N_16951,N_16518);
or U17398 (N_17398,N_16668,N_16968);
nand U17399 (N_17399,N_16871,N_16541);
and U17400 (N_17400,N_16993,N_16904);
and U17401 (N_17401,N_16875,N_16700);
nand U17402 (N_17402,N_16902,N_16991);
xnor U17403 (N_17403,N_16619,N_16903);
xor U17404 (N_17404,N_16777,N_16932);
xor U17405 (N_17405,N_16986,N_16951);
nor U17406 (N_17406,N_16948,N_16967);
xor U17407 (N_17407,N_16788,N_16658);
nand U17408 (N_17408,N_16615,N_16910);
or U17409 (N_17409,N_16596,N_16635);
and U17410 (N_17410,N_16673,N_16800);
nand U17411 (N_17411,N_16500,N_16999);
and U17412 (N_17412,N_16602,N_16777);
nand U17413 (N_17413,N_16763,N_16583);
or U17414 (N_17414,N_16933,N_16591);
nand U17415 (N_17415,N_16959,N_16895);
nor U17416 (N_17416,N_16688,N_16907);
or U17417 (N_17417,N_16779,N_16986);
xor U17418 (N_17418,N_16918,N_16937);
nand U17419 (N_17419,N_16749,N_16878);
nor U17420 (N_17420,N_16876,N_16792);
or U17421 (N_17421,N_16721,N_16597);
and U17422 (N_17422,N_16657,N_16715);
or U17423 (N_17423,N_16595,N_16603);
nor U17424 (N_17424,N_16799,N_16927);
or U17425 (N_17425,N_16971,N_16844);
or U17426 (N_17426,N_16878,N_16645);
nand U17427 (N_17427,N_16697,N_16907);
nor U17428 (N_17428,N_16798,N_16676);
or U17429 (N_17429,N_16676,N_16869);
xor U17430 (N_17430,N_16821,N_16981);
or U17431 (N_17431,N_16622,N_16807);
or U17432 (N_17432,N_16831,N_16633);
nand U17433 (N_17433,N_16624,N_16710);
and U17434 (N_17434,N_16794,N_16535);
or U17435 (N_17435,N_16612,N_16977);
xnor U17436 (N_17436,N_16939,N_16793);
nand U17437 (N_17437,N_16762,N_16524);
xnor U17438 (N_17438,N_16785,N_16902);
nor U17439 (N_17439,N_16886,N_16556);
xor U17440 (N_17440,N_16782,N_16624);
or U17441 (N_17441,N_16916,N_16845);
nand U17442 (N_17442,N_16887,N_16934);
and U17443 (N_17443,N_16535,N_16664);
xnor U17444 (N_17444,N_16615,N_16912);
nand U17445 (N_17445,N_16783,N_16624);
nor U17446 (N_17446,N_16756,N_16840);
nor U17447 (N_17447,N_16790,N_16590);
nor U17448 (N_17448,N_16986,N_16974);
nor U17449 (N_17449,N_16558,N_16522);
and U17450 (N_17450,N_16506,N_16679);
xor U17451 (N_17451,N_16668,N_16737);
or U17452 (N_17452,N_16919,N_16606);
or U17453 (N_17453,N_16529,N_16940);
or U17454 (N_17454,N_16960,N_16774);
nand U17455 (N_17455,N_16597,N_16748);
xor U17456 (N_17456,N_16686,N_16596);
xor U17457 (N_17457,N_16572,N_16899);
and U17458 (N_17458,N_16730,N_16865);
and U17459 (N_17459,N_16766,N_16608);
or U17460 (N_17460,N_16578,N_16814);
or U17461 (N_17461,N_16505,N_16818);
xnor U17462 (N_17462,N_16571,N_16713);
nand U17463 (N_17463,N_16834,N_16964);
nor U17464 (N_17464,N_16962,N_16975);
xnor U17465 (N_17465,N_16522,N_16650);
or U17466 (N_17466,N_16580,N_16602);
nor U17467 (N_17467,N_16821,N_16501);
or U17468 (N_17468,N_16616,N_16706);
or U17469 (N_17469,N_16990,N_16620);
nand U17470 (N_17470,N_16579,N_16837);
nand U17471 (N_17471,N_16828,N_16787);
nand U17472 (N_17472,N_16916,N_16513);
nor U17473 (N_17473,N_16855,N_16558);
and U17474 (N_17474,N_16998,N_16509);
xnor U17475 (N_17475,N_16713,N_16732);
xnor U17476 (N_17476,N_16761,N_16605);
nand U17477 (N_17477,N_16618,N_16621);
nor U17478 (N_17478,N_16887,N_16673);
nor U17479 (N_17479,N_16998,N_16622);
nor U17480 (N_17480,N_16951,N_16517);
xor U17481 (N_17481,N_16694,N_16768);
xnor U17482 (N_17482,N_16696,N_16607);
nor U17483 (N_17483,N_16657,N_16687);
or U17484 (N_17484,N_16949,N_16557);
xnor U17485 (N_17485,N_16896,N_16928);
and U17486 (N_17486,N_16746,N_16761);
nand U17487 (N_17487,N_16752,N_16562);
xnor U17488 (N_17488,N_16997,N_16523);
xnor U17489 (N_17489,N_16723,N_16957);
nand U17490 (N_17490,N_16675,N_16538);
and U17491 (N_17491,N_16775,N_16949);
or U17492 (N_17492,N_16844,N_16797);
nor U17493 (N_17493,N_16669,N_16771);
or U17494 (N_17494,N_16695,N_16725);
and U17495 (N_17495,N_16649,N_16550);
and U17496 (N_17496,N_16989,N_16902);
xor U17497 (N_17497,N_16977,N_16547);
nor U17498 (N_17498,N_16773,N_16952);
or U17499 (N_17499,N_16690,N_16835);
nand U17500 (N_17500,N_17120,N_17444);
or U17501 (N_17501,N_17168,N_17144);
nand U17502 (N_17502,N_17335,N_17198);
or U17503 (N_17503,N_17462,N_17019);
and U17504 (N_17504,N_17080,N_17219);
nor U17505 (N_17505,N_17495,N_17131);
nand U17506 (N_17506,N_17014,N_17107);
xor U17507 (N_17507,N_17244,N_17121);
and U17508 (N_17508,N_17027,N_17138);
nand U17509 (N_17509,N_17378,N_17343);
nand U17510 (N_17510,N_17347,N_17481);
xnor U17511 (N_17511,N_17383,N_17025);
or U17512 (N_17512,N_17409,N_17026);
and U17513 (N_17513,N_17263,N_17268);
nor U17514 (N_17514,N_17151,N_17452);
nor U17515 (N_17515,N_17426,N_17125);
and U17516 (N_17516,N_17057,N_17483);
xor U17517 (N_17517,N_17272,N_17251);
and U17518 (N_17518,N_17232,N_17436);
nor U17519 (N_17519,N_17275,N_17130);
xnor U17520 (N_17520,N_17078,N_17371);
or U17521 (N_17521,N_17377,N_17428);
xor U17522 (N_17522,N_17424,N_17210);
nand U17523 (N_17523,N_17306,N_17147);
and U17524 (N_17524,N_17134,N_17337);
and U17525 (N_17525,N_17466,N_17065);
nor U17526 (N_17526,N_17358,N_17240);
nor U17527 (N_17527,N_17063,N_17489);
nor U17528 (N_17528,N_17396,N_17017);
xnor U17529 (N_17529,N_17292,N_17259);
and U17530 (N_17530,N_17230,N_17357);
xnor U17531 (N_17531,N_17164,N_17160);
nand U17532 (N_17532,N_17202,N_17223);
xor U17533 (N_17533,N_17498,N_17177);
nand U17534 (N_17534,N_17088,N_17470);
and U17535 (N_17535,N_17446,N_17018);
and U17536 (N_17536,N_17294,N_17056);
or U17537 (N_17537,N_17074,N_17073);
and U17538 (N_17538,N_17200,N_17010);
nor U17539 (N_17539,N_17034,N_17264);
or U17540 (N_17540,N_17064,N_17286);
nand U17541 (N_17541,N_17171,N_17344);
nor U17542 (N_17542,N_17448,N_17234);
and U17543 (N_17543,N_17423,N_17256);
xnor U17544 (N_17544,N_17228,N_17252);
nor U17545 (N_17545,N_17174,N_17382);
or U17546 (N_17546,N_17356,N_17205);
xor U17547 (N_17547,N_17270,N_17413);
and U17548 (N_17548,N_17298,N_17077);
nand U17549 (N_17549,N_17070,N_17071);
and U17550 (N_17550,N_17109,N_17055);
nand U17551 (N_17551,N_17336,N_17053);
xnor U17552 (N_17552,N_17206,N_17432);
and U17553 (N_17553,N_17345,N_17392);
xnor U17554 (N_17554,N_17083,N_17295);
or U17555 (N_17555,N_17214,N_17415);
xnor U17556 (N_17556,N_17135,N_17283);
nor U17557 (N_17557,N_17112,N_17023);
nor U17558 (N_17558,N_17241,N_17370);
nand U17559 (N_17559,N_17373,N_17096);
nor U17560 (N_17560,N_17453,N_17299);
or U17561 (N_17561,N_17348,N_17476);
xor U17562 (N_17562,N_17410,N_17233);
xor U17563 (N_17563,N_17445,N_17167);
nand U17564 (N_17564,N_17119,N_17159);
nor U17565 (N_17565,N_17307,N_17076);
xor U17566 (N_17566,N_17290,N_17278);
or U17567 (N_17567,N_17208,N_17461);
xnor U17568 (N_17568,N_17173,N_17334);
nor U17569 (N_17569,N_17227,N_17172);
nor U17570 (N_17570,N_17439,N_17101);
nand U17571 (N_17571,N_17150,N_17485);
xnor U17572 (N_17572,N_17412,N_17261);
and U17573 (N_17573,N_17250,N_17406);
xor U17574 (N_17574,N_17490,N_17225);
nor U17575 (N_17575,N_17411,N_17108);
xor U17576 (N_17576,N_17287,N_17494);
and U17577 (N_17577,N_17280,N_17266);
or U17578 (N_17578,N_17381,N_17161);
nor U17579 (N_17579,N_17366,N_17044);
nand U17580 (N_17580,N_17199,N_17450);
nor U17581 (N_17581,N_17407,N_17408);
and U17582 (N_17582,N_17196,N_17342);
xor U17583 (N_17583,N_17218,N_17105);
and U17584 (N_17584,N_17006,N_17456);
or U17585 (N_17585,N_17184,N_17464);
nand U17586 (N_17586,N_17269,N_17005);
nor U17587 (N_17587,N_17049,N_17197);
or U17588 (N_17588,N_17089,N_17273);
nor U17589 (N_17589,N_17029,N_17060);
xnor U17590 (N_17590,N_17487,N_17169);
and U17591 (N_17591,N_17421,N_17414);
nand U17592 (N_17592,N_17098,N_17110);
or U17593 (N_17593,N_17157,N_17482);
and U17594 (N_17594,N_17440,N_17468);
nand U17595 (N_17595,N_17314,N_17441);
xor U17596 (N_17596,N_17085,N_17143);
and U17597 (N_17597,N_17166,N_17193);
or U17598 (N_17598,N_17099,N_17463);
nor U17599 (N_17599,N_17435,N_17403);
and U17600 (N_17600,N_17284,N_17431);
and U17601 (N_17601,N_17258,N_17082);
or U17602 (N_17602,N_17340,N_17380);
or U17603 (N_17603,N_17341,N_17192);
or U17604 (N_17604,N_17324,N_17308);
nand U17605 (N_17605,N_17246,N_17052);
nor U17606 (N_17606,N_17102,N_17117);
nor U17607 (N_17607,N_17021,N_17043);
or U17608 (N_17608,N_17391,N_17181);
nand U17609 (N_17609,N_17368,N_17459);
nor U17610 (N_17610,N_17028,N_17104);
xor U17611 (N_17611,N_17145,N_17066);
or U17612 (N_17612,N_17209,N_17022);
nand U17613 (N_17613,N_17187,N_17216);
nand U17614 (N_17614,N_17361,N_17020);
or U17615 (N_17615,N_17309,N_17374);
xor U17616 (N_17616,N_17058,N_17036);
nor U17617 (N_17617,N_17455,N_17402);
or U17618 (N_17618,N_17433,N_17352);
nor U17619 (N_17619,N_17221,N_17480);
xnor U17620 (N_17620,N_17457,N_17111);
or U17621 (N_17621,N_17296,N_17126);
or U17622 (N_17622,N_17115,N_17061);
nand U17623 (N_17623,N_17127,N_17301);
nand U17624 (N_17624,N_17097,N_17163);
nor U17625 (N_17625,N_17116,N_17386);
xor U17626 (N_17626,N_17247,N_17474);
xor U17627 (N_17627,N_17201,N_17437);
or U17628 (N_17628,N_17238,N_17353);
nand U17629 (N_17629,N_17090,N_17372);
nand U17630 (N_17630,N_17393,N_17087);
xnor U17631 (N_17631,N_17430,N_17322);
nand U17632 (N_17632,N_17364,N_17239);
xor U17633 (N_17633,N_17467,N_17072);
xnor U17634 (N_17634,N_17385,N_17009);
and U17635 (N_17635,N_17217,N_17154);
nor U17636 (N_17636,N_17190,N_17068);
and U17637 (N_17637,N_17041,N_17140);
and U17638 (N_17638,N_17038,N_17425);
or U17639 (N_17639,N_17422,N_17229);
xnor U17640 (N_17640,N_17062,N_17042);
and U17641 (N_17641,N_17222,N_17079);
nand U17642 (N_17642,N_17069,N_17325);
and U17643 (N_17643,N_17037,N_17323);
nor U17644 (N_17644,N_17282,N_17146);
nand U17645 (N_17645,N_17400,N_17122);
nor U17646 (N_17646,N_17458,N_17046);
and U17647 (N_17647,N_17390,N_17257);
nand U17648 (N_17648,N_17191,N_17379);
nor U17649 (N_17649,N_17367,N_17158);
nand U17650 (N_17650,N_17319,N_17451);
and U17651 (N_17651,N_17183,N_17478);
nor U17652 (N_17652,N_17152,N_17106);
xor U17653 (N_17653,N_17030,N_17103);
and U17654 (N_17654,N_17213,N_17260);
and U17655 (N_17655,N_17326,N_17339);
xor U17656 (N_17656,N_17404,N_17369);
xnor U17657 (N_17657,N_17491,N_17405);
nand U17658 (N_17658,N_17387,N_17279);
or U17659 (N_17659,N_17186,N_17024);
nand U17660 (N_17660,N_17050,N_17033);
or U17661 (N_17661,N_17248,N_17059);
nand U17662 (N_17662,N_17175,N_17417);
nand U17663 (N_17663,N_17486,N_17471);
and U17664 (N_17664,N_17189,N_17047);
or U17665 (N_17665,N_17291,N_17262);
or U17666 (N_17666,N_17304,N_17276);
and U17667 (N_17667,N_17351,N_17091);
nor U17668 (N_17668,N_17312,N_17203);
or U17669 (N_17669,N_17011,N_17300);
xnor U17670 (N_17670,N_17162,N_17472);
or U17671 (N_17671,N_17013,N_17313);
xor U17672 (N_17672,N_17418,N_17320);
xnor U17673 (N_17673,N_17315,N_17363);
or U17674 (N_17674,N_17499,N_17447);
or U17675 (N_17675,N_17084,N_17086);
nand U17676 (N_17676,N_17438,N_17460);
nor U17677 (N_17677,N_17132,N_17317);
or U17678 (N_17678,N_17092,N_17093);
nand U17679 (N_17679,N_17094,N_17204);
nor U17680 (N_17680,N_17465,N_17182);
or U17681 (N_17681,N_17195,N_17429);
xor U17682 (N_17682,N_17302,N_17350);
nor U17683 (N_17683,N_17484,N_17318);
nor U17684 (N_17684,N_17002,N_17321);
xnor U17685 (N_17685,N_17442,N_17496);
and U17686 (N_17686,N_17355,N_17277);
xnor U17687 (N_17687,N_17118,N_17016);
nor U17688 (N_17688,N_17039,N_17427);
and U17689 (N_17689,N_17349,N_17267);
or U17690 (N_17690,N_17443,N_17207);
nand U17691 (N_17691,N_17149,N_17303);
and U17692 (N_17692,N_17040,N_17156);
nor U17693 (N_17693,N_17124,N_17100);
or U17694 (N_17694,N_17274,N_17012);
xnor U17695 (N_17695,N_17285,N_17170);
and U17696 (N_17696,N_17416,N_17155);
xnor U17697 (N_17697,N_17139,N_17031);
and U17698 (N_17698,N_17449,N_17137);
xor U17699 (N_17699,N_17114,N_17311);
and U17700 (N_17700,N_17305,N_17395);
nor U17701 (N_17701,N_17129,N_17123);
nor U17702 (N_17702,N_17255,N_17376);
nor U17703 (N_17703,N_17265,N_17331);
xor U17704 (N_17704,N_17067,N_17253);
or U17705 (N_17705,N_17165,N_17237);
xnor U17706 (N_17706,N_17384,N_17288);
nor U17707 (N_17707,N_17243,N_17310);
or U17708 (N_17708,N_17330,N_17113);
nor U17709 (N_17709,N_17180,N_17211);
nand U17710 (N_17710,N_17254,N_17338);
nor U17711 (N_17711,N_17015,N_17008);
nand U17712 (N_17712,N_17420,N_17316);
nor U17713 (N_17713,N_17128,N_17188);
or U17714 (N_17714,N_17136,N_17035);
or U17715 (N_17715,N_17220,N_17394);
nand U17716 (N_17716,N_17289,N_17469);
nor U17717 (N_17717,N_17245,N_17075);
and U17718 (N_17718,N_17148,N_17051);
or U17719 (N_17719,N_17133,N_17389);
nor U17720 (N_17720,N_17488,N_17194);
nand U17721 (N_17721,N_17479,N_17329);
or U17722 (N_17722,N_17001,N_17003);
or U17723 (N_17723,N_17271,N_17492);
or U17724 (N_17724,N_17419,N_17493);
nand U17725 (N_17725,N_17327,N_17360);
xnor U17726 (N_17726,N_17176,N_17231);
nand U17727 (N_17727,N_17000,N_17399);
xor U17728 (N_17728,N_17141,N_17328);
or U17729 (N_17729,N_17475,N_17293);
nor U17730 (N_17730,N_17401,N_17153);
nand U17731 (N_17731,N_17185,N_17215);
nor U17732 (N_17732,N_17359,N_17346);
or U17733 (N_17733,N_17477,N_17142);
and U17734 (N_17734,N_17397,N_17242);
xor U17735 (N_17735,N_17236,N_17045);
or U17736 (N_17736,N_17054,N_17179);
nand U17737 (N_17737,N_17454,N_17048);
nand U17738 (N_17738,N_17212,N_17434);
xnor U17739 (N_17739,N_17365,N_17224);
nor U17740 (N_17740,N_17333,N_17178);
or U17741 (N_17741,N_17226,N_17297);
xnor U17742 (N_17742,N_17473,N_17497);
xor U17743 (N_17743,N_17375,N_17007);
nor U17744 (N_17744,N_17281,N_17388);
nor U17745 (N_17745,N_17362,N_17081);
xor U17746 (N_17746,N_17235,N_17398);
nor U17747 (N_17747,N_17095,N_17004);
or U17748 (N_17748,N_17332,N_17354);
and U17749 (N_17749,N_17032,N_17249);
or U17750 (N_17750,N_17472,N_17154);
nand U17751 (N_17751,N_17177,N_17367);
and U17752 (N_17752,N_17030,N_17273);
or U17753 (N_17753,N_17103,N_17010);
or U17754 (N_17754,N_17250,N_17045);
nand U17755 (N_17755,N_17143,N_17236);
nand U17756 (N_17756,N_17323,N_17467);
and U17757 (N_17757,N_17293,N_17012);
and U17758 (N_17758,N_17129,N_17126);
nand U17759 (N_17759,N_17022,N_17237);
nor U17760 (N_17760,N_17408,N_17413);
or U17761 (N_17761,N_17183,N_17468);
nor U17762 (N_17762,N_17178,N_17182);
and U17763 (N_17763,N_17145,N_17074);
nor U17764 (N_17764,N_17335,N_17303);
nor U17765 (N_17765,N_17208,N_17276);
nor U17766 (N_17766,N_17011,N_17414);
nor U17767 (N_17767,N_17483,N_17428);
nand U17768 (N_17768,N_17473,N_17475);
or U17769 (N_17769,N_17278,N_17198);
nor U17770 (N_17770,N_17401,N_17266);
or U17771 (N_17771,N_17070,N_17425);
and U17772 (N_17772,N_17153,N_17379);
or U17773 (N_17773,N_17049,N_17349);
xnor U17774 (N_17774,N_17113,N_17050);
or U17775 (N_17775,N_17209,N_17384);
and U17776 (N_17776,N_17184,N_17004);
and U17777 (N_17777,N_17393,N_17476);
xnor U17778 (N_17778,N_17455,N_17277);
nand U17779 (N_17779,N_17160,N_17423);
or U17780 (N_17780,N_17218,N_17128);
or U17781 (N_17781,N_17100,N_17241);
xor U17782 (N_17782,N_17429,N_17309);
xnor U17783 (N_17783,N_17417,N_17086);
xor U17784 (N_17784,N_17087,N_17461);
and U17785 (N_17785,N_17081,N_17281);
xor U17786 (N_17786,N_17254,N_17307);
xor U17787 (N_17787,N_17346,N_17434);
and U17788 (N_17788,N_17159,N_17223);
nand U17789 (N_17789,N_17493,N_17394);
nand U17790 (N_17790,N_17383,N_17126);
xnor U17791 (N_17791,N_17076,N_17245);
and U17792 (N_17792,N_17028,N_17384);
and U17793 (N_17793,N_17015,N_17457);
and U17794 (N_17794,N_17149,N_17259);
nor U17795 (N_17795,N_17035,N_17431);
and U17796 (N_17796,N_17380,N_17405);
xnor U17797 (N_17797,N_17468,N_17250);
and U17798 (N_17798,N_17339,N_17042);
or U17799 (N_17799,N_17281,N_17484);
xnor U17800 (N_17800,N_17170,N_17328);
and U17801 (N_17801,N_17187,N_17202);
or U17802 (N_17802,N_17349,N_17226);
nand U17803 (N_17803,N_17129,N_17104);
xor U17804 (N_17804,N_17091,N_17257);
xnor U17805 (N_17805,N_17338,N_17363);
xnor U17806 (N_17806,N_17064,N_17440);
nor U17807 (N_17807,N_17146,N_17154);
nor U17808 (N_17808,N_17006,N_17315);
nor U17809 (N_17809,N_17456,N_17007);
xnor U17810 (N_17810,N_17192,N_17087);
or U17811 (N_17811,N_17247,N_17309);
xnor U17812 (N_17812,N_17360,N_17115);
xor U17813 (N_17813,N_17145,N_17241);
and U17814 (N_17814,N_17071,N_17293);
xnor U17815 (N_17815,N_17374,N_17016);
nand U17816 (N_17816,N_17230,N_17417);
xor U17817 (N_17817,N_17052,N_17261);
nor U17818 (N_17818,N_17445,N_17455);
nand U17819 (N_17819,N_17246,N_17397);
and U17820 (N_17820,N_17386,N_17071);
and U17821 (N_17821,N_17262,N_17468);
nand U17822 (N_17822,N_17083,N_17198);
nand U17823 (N_17823,N_17308,N_17167);
nand U17824 (N_17824,N_17144,N_17310);
xnor U17825 (N_17825,N_17205,N_17417);
and U17826 (N_17826,N_17028,N_17417);
and U17827 (N_17827,N_17206,N_17229);
xnor U17828 (N_17828,N_17057,N_17095);
nand U17829 (N_17829,N_17272,N_17467);
nand U17830 (N_17830,N_17211,N_17385);
or U17831 (N_17831,N_17261,N_17210);
or U17832 (N_17832,N_17130,N_17254);
nand U17833 (N_17833,N_17147,N_17380);
nor U17834 (N_17834,N_17126,N_17024);
xor U17835 (N_17835,N_17432,N_17190);
nor U17836 (N_17836,N_17455,N_17306);
xor U17837 (N_17837,N_17481,N_17108);
nand U17838 (N_17838,N_17126,N_17370);
nor U17839 (N_17839,N_17344,N_17455);
nand U17840 (N_17840,N_17422,N_17302);
and U17841 (N_17841,N_17320,N_17119);
or U17842 (N_17842,N_17264,N_17301);
nand U17843 (N_17843,N_17246,N_17177);
and U17844 (N_17844,N_17359,N_17086);
xnor U17845 (N_17845,N_17358,N_17195);
or U17846 (N_17846,N_17063,N_17051);
and U17847 (N_17847,N_17395,N_17110);
and U17848 (N_17848,N_17451,N_17376);
or U17849 (N_17849,N_17442,N_17403);
nor U17850 (N_17850,N_17084,N_17161);
or U17851 (N_17851,N_17090,N_17204);
xnor U17852 (N_17852,N_17220,N_17397);
nor U17853 (N_17853,N_17393,N_17016);
nand U17854 (N_17854,N_17433,N_17228);
and U17855 (N_17855,N_17030,N_17397);
or U17856 (N_17856,N_17427,N_17386);
or U17857 (N_17857,N_17031,N_17166);
nor U17858 (N_17858,N_17210,N_17041);
nand U17859 (N_17859,N_17356,N_17478);
nor U17860 (N_17860,N_17127,N_17311);
nand U17861 (N_17861,N_17252,N_17087);
nor U17862 (N_17862,N_17045,N_17156);
or U17863 (N_17863,N_17492,N_17335);
nand U17864 (N_17864,N_17253,N_17290);
xor U17865 (N_17865,N_17099,N_17029);
and U17866 (N_17866,N_17463,N_17306);
nor U17867 (N_17867,N_17222,N_17449);
and U17868 (N_17868,N_17319,N_17232);
and U17869 (N_17869,N_17457,N_17147);
xor U17870 (N_17870,N_17256,N_17086);
nor U17871 (N_17871,N_17231,N_17471);
and U17872 (N_17872,N_17230,N_17028);
and U17873 (N_17873,N_17236,N_17250);
xor U17874 (N_17874,N_17491,N_17364);
nand U17875 (N_17875,N_17313,N_17310);
xor U17876 (N_17876,N_17147,N_17311);
nand U17877 (N_17877,N_17299,N_17236);
or U17878 (N_17878,N_17013,N_17467);
or U17879 (N_17879,N_17237,N_17116);
xor U17880 (N_17880,N_17280,N_17438);
xor U17881 (N_17881,N_17292,N_17421);
xnor U17882 (N_17882,N_17067,N_17140);
and U17883 (N_17883,N_17210,N_17047);
or U17884 (N_17884,N_17104,N_17475);
or U17885 (N_17885,N_17014,N_17468);
nor U17886 (N_17886,N_17060,N_17353);
nor U17887 (N_17887,N_17038,N_17235);
or U17888 (N_17888,N_17163,N_17217);
or U17889 (N_17889,N_17118,N_17388);
xnor U17890 (N_17890,N_17266,N_17345);
nand U17891 (N_17891,N_17293,N_17145);
nor U17892 (N_17892,N_17070,N_17144);
nor U17893 (N_17893,N_17030,N_17134);
or U17894 (N_17894,N_17285,N_17333);
or U17895 (N_17895,N_17440,N_17126);
xor U17896 (N_17896,N_17142,N_17282);
nand U17897 (N_17897,N_17137,N_17037);
nand U17898 (N_17898,N_17493,N_17431);
xor U17899 (N_17899,N_17216,N_17171);
nand U17900 (N_17900,N_17259,N_17463);
nand U17901 (N_17901,N_17466,N_17154);
or U17902 (N_17902,N_17115,N_17347);
xnor U17903 (N_17903,N_17438,N_17396);
nand U17904 (N_17904,N_17019,N_17215);
nand U17905 (N_17905,N_17352,N_17408);
xnor U17906 (N_17906,N_17102,N_17042);
xnor U17907 (N_17907,N_17158,N_17102);
or U17908 (N_17908,N_17304,N_17272);
or U17909 (N_17909,N_17447,N_17151);
nand U17910 (N_17910,N_17481,N_17061);
and U17911 (N_17911,N_17284,N_17035);
nor U17912 (N_17912,N_17143,N_17358);
or U17913 (N_17913,N_17221,N_17302);
nor U17914 (N_17914,N_17322,N_17478);
nand U17915 (N_17915,N_17212,N_17295);
nand U17916 (N_17916,N_17249,N_17350);
or U17917 (N_17917,N_17052,N_17220);
nor U17918 (N_17918,N_17464,N_17363);
xor U17919 (N_17919,N_17349,N_17059);
and U17920 (N_17920,N_17026,N_17438);
or U17921 (N_17921,N_17097,N_17370);
nor U17922 (N_17922,N_17350,N_17354);
and U17923 (N_17923,N_17233,N_17096);
nor U17924 (N_17924,N_17431,N_17350);
nand U17925 (N_17925,N_17127,N_17357);
and U17926 (N_17926,N_17250,N_17394);
and U17927 (N_17927,N_17414,N_17264);
nor U17928 (N_17928,N_17128,N_17305);
nand U17929 (N_17929,N_17143,N_17176);
nand U17930 (N_17930,N_17027,N_17189);
xnor U17931 (N_17931,N_17410,N_17411);
xor U17932 (N_17932,N_17028,N_17040);
and U17933 (N_17933,N_17001,N_17395);
xnor U17934 (N_17934,N_17131,N_17444);
or U17935 (N_17935,N_17091,N_17109);
or U17936 (N_17936,N_17346,N_17389);
nor U17937 (N_17937,N_17418,N_17197);
and U17938 (N_17938,N_17398,N_17133);
nor U17939 (N_17939,N_17104,N_17447);
xor U17940 (N_17940,N_17101,N_17427);
and U17941 (N_17941,N_17319,N_17399);
nand U17942 (N_17942,N_17307,N_17389);
nand U17943 (N_17943,N_17269,N_17368);
and U17944 (N_17944,N_17311,N_17437);
or U17945 (N_17945,N_17442,N_17349);
nor U17946 (N_17946,N_17230,N_17450);
and U17947 (N_17947,N_17180,N_17014);
nor U17948 (N_17948,N_17012,N_17479);
and U17949 (N_17949,N_17144,N_17427);
nand U17950 (N_17950,N_17175,N_17101);
xnor U17951 (N_17951,N_17393,N_17396);
nor U17952 (N_17952,N_17205,N_17077);
or U17953 (N_17953,N_17173,N_17042);
nor U17954 (N_17954,N_17302,N_17444);
and U17955 (N_17955,N_17122,N_17463);
nand U17956 (N_17956,N_17052,N_17016);
xnor U17957 (N_17957,N_17403,N_17425);
and U17958 (N_17958,N_17061,N_17045);
or U17959 (N_17959,N_17299,N_17246);
or U17960 (N_17960,N_17385,N_17432);
or U17961 (N_17961,N_17240,N_17428);
and U17962 (N_17962,N_17480,N_17306);
nor U17963 (N_17963,N_17202,N_17226);
xnor U17964 (N_17964,N_17157,N_17244);
nor U17965 (N_17965,N_17296,N_17109);
nor U17966 (N_17966,N_17437,N_17208);
nand U17967 (N_17967,N_17466,N_17462);
nor U17968 (N_17968,N_17080,N_17450);
and U17969 (N_17969,N_17486,N_17058);
and U17970 (N_17970,N_17000,N_17369);
or U17971 (N_17971,N_17216,N_17221);
nor U17972 (N_17972,N_17323,N_17283);
or U17973 (N_17973,N_17203,N_17034);
nand U17974 (N_17974,N_17037,N_17018);
nor U17975 (N_17975,N_17184,N_17288);
nand U17976 (N_17976,N_17287,N_17081);
or U17977 (N_17977,N_17005,N_17419);
and U17978 (N_17978,N_17375,N_17430);
nand U17979 (N_17979,N_17475,N_17463);
nand U17980 (N_17980,N_17361,N_17128);
and U17981 (N_17981,N_17166,N_17225);
nor U17982 (N_17982,N_17472,N_17308);
nor U17983 (N_17983,N_17200,N_17324);
xor U17984 (N_17984,N_17038,N_17198);
xor U17985 (N_17985,N_17433,N_17273);
nor U17986 (N_17986,N_17263,N_17146);
or U17987 (N_17987,N_17252,N_17349);
or U17988 (N_17988,N_17395,N_17041);
nand U17989 (N_17989,N_17192,N_17351);
xnor U17990 (N_17990,N_17249,N_17096);
xnor U17991 (N_17991,N_17002,N_17092);
nor U17992 (N_17992,N_17413,N_17024);
xor U17993 (N_17993,N_17396,N_17287);
or U17994 (N_17994,N_17267,N_17023);
and U17995 (N_17995,N_17377,N_17472);
and U17996 (N_17996,N_17077,N_17352);
nand U17997 (N_17997,N_17212,N_17438);
and U17998 (N_17998,N_17052,N_17425);
or U17999 (N_17999,N_17202,N_17305);
nor U18000 (N_18000,N_17943,N_17758);
nand U18001 (N_18001,N_17530,N_17507);
nor U18002 (N_18002,N_17951,N_17551);
and U18003 (N_18003,N_17857,N_17583);
or U18004 (N_18004,N_17839,N_17827);
and U18005 (N_18005,N_17947,N_17509);
and U18006 (N_18006,N_17990,N_17954);
xor U18007 (N_18007,N_17706,N_17993);
and U18008 (N_18008,N_17878,N_17793);
nor U18009 (N_18009,N_17974,N_17569);
or U18010 (N_18010,N_17541,N_17816);
nor U18011 (N_18011,N_17899,N_17506);
and U18012 (N_18012,N_17595,N_17739);
nand U18013 (N_18013,N_17754,N_17512);
nor U18014 (N_18014,N_17538,N_17669);
nand U18015 (N_18015,N_17599,N_17623);
or U18016 (N_18016,N_17838,N_17520);
and U18017 (N_18017,N_17880,N_17535);
and U18018 (N_18018,N_17695,N_17783);
nor U18019 (N_18019,N_17784,N_17961);
and U18020 (N_18020,N_17813,N_17871);
and U18021 (N_18021,N_17720,N_17637);
or U18022 (N_18022,N_17744,N_17722);
xnor U18023 (N_18023,N_17588,N_17982);
and U18024 (N_18024,N_17630,N_17667);
xnor U18025 (N_18025,N_17946,N_17928);
or U18026 (N_18026,N_17879,N_17929);
and U18027 (N_18027,N_17658,N_17850);
nand U18028 (N_18028,N_17619,N_17934);
or U18029 (N_18029,N_17640,N_17989);
nor U18030 (N_18030,N_17792,N_17740);
nor U18031 (N_18031,N_17514,N_17851);
and U18032 (N_18032,N_17684,N_17992);
nor U18033 (N_18033,N_17962,N_17615);
or U18034 (N_18034,N_17700,N_17876);
and U18035 (N_18035,N_17767,N_17981);
nor U18036 (N_18036,N_17930,N_17516);
and U18037 (N_18037,N_17939,N_17788);
and U18038 (N_18038,N_17896,N_17560);
nand U18039 (N_18039,N_17650,N_17859);
nor U18040 (N_18040,N_17842,N_17935);
or U18041 (N_18041,N_17906,N_17780);
nor U18042 (N_18042,N_17515,N_17620);
xor U18043 (N_18043,N_17887,N_17611);
and U18044 (N_18044,N_17873,N_17733);
or U18045 (N_18045,N_17654,N_17749);
nor U18046 (N_18046,N_17821,N_17957);
nor U18047 (N_18047,N_17950,N_17971);
or U18048 (N_18048,N_17736,N_17725);
and U18049 (N_18049,N_17846,N_17634);
or U18050 (N_18050,N_17872,N_17653);
and U18051 (N_18051,N_17984,N_17673);
xnor U18052 (N_18052,N_17689,N_17796);
xor U18053 (N_18053,N_17723,N_17729);
and U18054 (N_18054,N_17964,N_17750);
nor U18055 (N_18055,N_17881,N_17766);
xor U18056 (N_18056,N_17558,N_17748);
and U18057 (N_18057,N_17730,N_17570);
nor U18058 (N_18058,N_17718,N_17622);
xor U18059 (N_18059,N_17609,N_17837);
xnor U18060 (N_18060,N_17557,N_17546);
nor U18061 (N_18061,N_17855,N_17809);
or U18062 (N_18062,N_17973,N_17843);
nor U18063 (N_18063,N_17756,N_17913);
xnor U18064 (N_18064,N_17726,N_17605);
nand U18065 (N_18065,N_17936,N_17772);
or U18066 (N_18066,N_17676,N_17548);
nor U18067 (N_18067,N_17606,N_17870);
nand U18068 (N_18068,N_17844,N_17968);
xor U18069 (N_18069,N_17806,N_17685);
xnor U18070 (N_18070,N_17578,N_17907);
and U18071 (N_18071,N_17563,N_17521);
or U18072 (N_18072,N_17678,N_17979);
xnor U18073 (N_18073,N_17602,N_17760);
or U18074 (N_18074,N_17747,N_17817);
and U18075 (N_18075,N_17511,N_17608);
and U18076 (N_18076,N_17893,N_17918);
and U18077 (N_18077,N_17901,N_17576);
nor U18078 (N_18078,N_17713,N_17504);
nor U18079 (N_18079,N_17638,N_17841);
or U18080 (N_18080,N_17709,N_17824);
and U18081 (N_18081,N_17998,N_17745);
nor U18082 (N_18082,N_17651,N_17627);
xnor U18083 (N_18083,N_17645,N_17727);
and U18084 (N_18084,N_17549,N_17617);
and U18085 (N_18085,N_17986,N_17755);
or U18086 (N_18086,N_17539,N_17526);
nor U18087 (N_18087,N_17952,N_17501);
or U18088 (N_18088,N_17815,N_17944);
nor U18089 (N_18089,N_17581,N_17693);
or U18090 (N_18090,N_17626,N_17781);
nand U18091 (N_18091,N_17942,N_17810);
nor U18092 (N_18092,N_17687,N_17579);
nor U18093 (N_18093,N_17900,N_17932);
or U18094 (N_18094,N_17925,N_17875);
or U18095 (N_18095,N_17532,N_17519);
xnor U18096 (N_18096,N_17540,N_17829);
nand U18097 (N_18097,N_17681,N_17902);
nand U18098 (N_18098,N_17959,N_17797);
or U18099 (N_18099,N_17912,N_17778);
and U18100 (N_18100,N_17811,N_17545);
nand U18101 (N_18101,N_17775,N_17625);
and U18102 (N_18102,N_17911,N_17597);
or U18103 (N_18103,N_17735,N_17831);
nand U18104 (N_18104,N_17874,N_17594);
nand U18105 (N_18105,N_17711,N_17572);
xor U18106 (N_18106,N_17920,N_17861);
xnor U18107 (N_18107,N_17891,N_17805);
or U18108 (N_18108,N_17697,N_17728);
xnor U18109 (N_18109,N_17975,N_17629);
nand U18110 (N_18110,N_17983,N_17853);
and U18111 (N_18111,N_17789,N_17704);
or U18112 (N_18112,N_17537,N_17502);
nor U18113 (N_18113,N_17826,N_17898);
or U18114 (N_18114,N_17682,N_17799);
xor U18115 (N_18115,N_17867,N_17888);
xnor U18116 (N_18116,N_17852,N_17794);
nand U18117 (N_18117,N_17845,N_17980);
and U18118 (N_18118,N_17941,N_17690);
and U18119 (N_18119,N_17644,N_17836);
nand U18120 (N_18120,N_17927,N_17802);
or U18121 (N_18121,N_17694,N_17931);
xor U18122 (N_18122,N_17656,N_17641);
nand U18123 (N_18123,N_17812,N_17624);
nor U18124 (N_18124,N_17790,N_17856);
and U18125 (N_18125,N_17833,N_17956);
nor U18126 (N_18126,N_17719,N_17593);
nand U18127 (N_18127,N_17905,N_17568);
xnor U18128 (N_18128,N_17702,N_17643);
nand U18129 (N_18129,N_17705,N_17916);
or U18130 (N_18130,N_17777,N_17807);
nor U18131 (N_18131,N_17544,N_17863);
or U18132 (N_18132,N_17721,N_17590);
or U18133 (N_18133,N_17751,N_17786);
nand U18134 (N_18134,N_17828,N_17714);
nor U18135 (N_18135,N_17573,N_17825);
xor U18136 (N_18136,N_17610,N_17771);
xor U18137 (N_18137,N_17525,N_17921);
or U18138 (N_18138,N_17948,N_17785);
xor U18139 (N_18139,N_17529,N_17661);
nand U18140 (N_18140,N_17686,N_17591);
nand U18141 (N_18141,N_17621,N_17963);
nand U18142 (N_18142,N_17782,N_17562);
nand U18143 (N_18143,N_17988,N_17612);
and U18144 (N_18144,N_17970,N_17660);
nor U18145 (N_18145,N_17655,N_17908);
nor U18146 (N_18146,N_17742,N_17890);
nor U18147 (N_18147,N_17604,N_17741);
or U18148 (N_18148,N_17769,N_17528);
nand U18149 (N_18149,N_17701,N_17692);
nor U18150 (N_18150,N_17996,N_17864);
nor U18151 (N_18151,N_17699,N_17814);
and U18152 (N_18152,N_17691,N_17734);
and U18153 (N_18153,N_17779,N_17909);
or U18154 (N_18154,N_17584,N_17757);
and U18155 (N_18155,N_17616,N_17882);
and U18156 (N_18156,N_17798,N_17999);
or U18157 (N_18157,N_17647,N_17972);
nand U18158 (N_18158,N_17803,N_17668);
nor U18159 (N_18159,N_17915,N_17587);
nand U18160 (N_18160,N_17724,N_17768);
or U18161 (N_18161,N_17601,N_17503);
nand U18162 (N_18162,N_17577,N_17834);
nor U18163 (N_18163,N_17670,N_17567);
nand U18164 (N_18164,N_17997,N_17663);
nor U18165 (N_18165,N_17924,N_17848);
xor U18166 (N_18166,N_17613,N_17830);
nand U18167 (N_18167,N_17508,N_17533);
or U18168 (N_18168,N_17642,N_17820);
and U18169 (N_18169,N_17987,N_17832);
and U18170 (N_18170,N_17865,N_17672);
nand U18171 (N_18171,N_17554,N_17543);
xnor U18172 (N_18172,N_17737,N_17743);
or U18173 (N_18173,N_17862,N_17703);
nor U18174 (N_18174,N_17522,N_17536);
nor U18175 (N_18175,N_17565,N_17715);
xor U18176 (N_18176,N_17589,N_17712);
or U18177 (N_18177,N_17835,N_17823);
nand U18178 (N_18178,N_17860,N_17732);
nor U18179 (N_18179,N_17556,N_17534);
or U18180 (N_18180,N_17618,N_17894);
xor U18181 (N_18181,N_17903,N_17523);
or U18182 (N_18182,N_17688,N_17822);
nor U18183 (N_18183,N_17991,N_17542);
or U18184 (N_18184,N_17698,N_17636);
and U18185 (N_18185,N_17889,N_17994);
and U18186 (N_18186,N_17664,N_17804);
xor U18187 (N_18187,N_17633,N_17665);
or U18188 (N_18188,N_17598,N_17763);
xor U18189 (N_18189,N_17659,N_17883);
or U18190 (N_18190,N_17513,N_17960);
nand U18191 (N_18191,N_17679,N_17919);
nor U18192 (N_18192,N_17759,N_17868);
nand U18193 (N_18193,N_17949,N_17580);
nand U18194 (N_18194,N_17564,N_17761);
and U18195 (N_18195,N_17505,N_17877);
nand U18196 (N_18196,N_17635,N_17716);
nand U18197 (N_18197,N_17800,N_17574);
or U18198 (N_18198,N_17858,N_17914);
nor U18199 (N_18199,N_17738,N_17607);
and U18200 (N_18200,N_17886,N_17897);
nand U18201 (N_18201,N_17510,N_17631);
and U18202 (N_18202,N_17801,N_17585);
or U18203 (N_18203,N_17995,N_17531);
nor U18204 (N_18204,N_17600,N_17648);
nor U18205 (N_18205,N_17976,N_17885);
nor U18206 (N_18206,N_17603,N_17985);
and U18207 (N_18207,N_17884,N_17680);
and U18208 (N_18208,N_17808,N_17707);
nor U18209 (N_18209,N_17787,N_17552);
xor U18210 (N_18210,N_17937,N_17869);
nor U18211 (N_18211,N_17500,N_17818);
and U18212 (N_18212,N_17596,N_17965);
and U18213 (N_18213,N_17776,N_17773);
nor U18214 (N_18214,N_17649,N_17847);
nand U18215 (N_18215,N_17662,N_17746);
and U18216 (N_18216,N_17555,N_17940);
xnor U18217 (N_18217,N_17866,N_17892);
or U18218 (N_18218,N_17671,N_17517);
xor U18219 (N_18219,N_17518,N_17571);
nand U18220 (N_18220,N_17628,N_17675);
xor U18221 (N_18221,N_17657,N_17917);
nor U18222 (N_18222,N_17895,N_17770);
xor U18223 (N_18223,N_17639,N_17550);
xnor U18224 (N_18224,N_17632,N_17904);
nor U18225 (N_18225,N_17708,N_17582);
nand U18226 (N_18226,N_17945,N_17566);
nor U18227 (N_18227,N_17677,N_17969);
nor U18228 (N_18228,N_17666,N_17652);
xor U18229 (N_18229,N_17774,N_17592);
nor U18230 (N_18230,N_17559,N_17731);
or U18231 (N_18231,N_17795,N_17953);
or U18232 (N_18232,N_17955,N_17753);
nor U18233 (N_18233,N_17764,N_17717);
nor U18234 (N_18234,N_17938,N_17575);
and U18235 (N_18235,N_17527,N_17854);
and U18236 (N_18236,N_17765,N_17710);
nor U18237 (N_18237,N_17762,N_17910);
or U18238 (N_18238,N_17524,N_17674);
or U18239 (N_18239,N_17840,N_17561);
nand U18240 (N_18240,N_17977,N_17614);
nand U18241 (N_18241,N_17926,N_17696);
and U18242 (N_18242,N_17967,N_17553);
and U18243 (N_18243,N_17933,N_17683);
nor U18244 (N_18244,N_17958,N_17966);
nor U18245 (N_18245,N_17547,N_17978);
nor U18246 (N_18246,N_17752,N_17819);
nand U18247 (N_18247,N_17849,N_17923);
nor U18248 (N_18248,N_17922,N_17646);
nor U18249 (N_18249,N_17791,N_17586);
nor U18250 (N_18250,N_17994,N_17857);
or U18251 (N_18251,N_17749,N_17789);
nor U18252 (N_18252,N_17856,N_17844);
xnor U18253 (N_18253,N_17633,N_17718);
xor U18254 (N_18254,N_17751,N_17942);
or U18255 (N_18255,N_17718,N_17679);
or U18256 (N_18256,N_17531,N_17874);
xor U18257 (N_18257,N_17947,N_17735);
or U18258 (N_18258,N_17799,N_17843);
and U18259 (N_18259,N_17912,N_17751);
and U18260 (N_18260,N_17945,N_17532);
nand U18261 (N_18261,N_17915,N_17929);
and U18262 (N_18262,N_17783,N_17545);
nor U18263 (N_18263,N_17728,N_17581);
and U18264 (N_18264,N_17518,N_17746);
nor U18265 (N_18265,N_17833,N_17549);
nor U18266 (N_18266,N_17973,N_17743);
nand U18267 (N_18267,N_17699,N_17905);
and U18268 (N_18268,N_17801,N_17987);
or U18269 (N_18269,N_17536,N_17977);
nand U18270 (N_18270,N_17540,N_17931);
or U18271 (N_18271,N_17561,N_17727);
or U18272 (N_18272,N_17513,N_17584);
nor U18273 (N_18273,N_17507,N_17528);
and U18274 (N_18274,N_17517,N_17885);
and U18275 (N_18275,N_17643,N_17835);
nor U18276 (N_18276,N_17638,N_17770);
nor U18277 (N_18277,N_17927,N_17546);
nor U18278 (N_18278,N_17986,N_17588);
nor U18279 (N_18279,N_17583,N_17961);
xnor U18280 (N_18280,N_17748,N_17908);
nor U18281 (N_18281,N_17659,N_17804);
xnor U18282 (N_18282,N_17806,N_17699);
nor U18283 (N_18283,N_17509,N_17746);
nor U18284 (N_18284,N_17575,N_17952);
nand U18285 (N_18285,N_17982,N_17604);
or U18286 (N_18286,N_17611,N_17840);
xor U18287 (N_18287,N_17718,N_17737);
or U18288 (N_18288,N_17853,N_17528);
nand U18289 (N_18289,N_17574,N_17888);
nand U18290 (N_18290,N_17944,N_17524);
and U18291 (N_18291,N_17631,N_17692);
nand U18292 (N_18292,N_17503,N_17541);
or U18293 (N_18293,N_17548,N_17598);
nand U18294 (N_18294,N_17778,N_17803);
and U18295 (N_18295,N_17762,N_17751);
nand U18296 (N_18296,N_17741,N_17590);
nand U18297 (N_18297,N_17800,N_17536);
or U18298 (N_18298,N_17534,N_17555);
nor U18299 (N_18299,N_17756,N_17984);
and U18300 (N_18300,N_17969,N_17508);
or U18301 (N_18301,N_17804,N_17882);
nor U18302 (N_18302,N_17828,N_17740);
xnor U18303 (N_18303,N_17675,N_17881);
xor U18304 (N_18304,N_17632,N_17839);
xnor U18305 (N_18305,N_17626,N_17895);
xnor U18306 (N_18306,N_17679,N_17706);
or U18307 (N_18307,N_17817,N_17521);
xor U18308 (N_18308,N_17919,N_17901);
and U18309 (N_18309,N_17501,N_17974);
or U18310 (N_18310,N_17514,N_17875);
and U18311 (N_18311,N_17603,N_17635);
nand U18312 (N_18312,N_17674,N_17724);
xor U18313 (N_18313,N_17625,N_17733);
nand U18314 (N_18314,N_17985,N_17624);
nand U18315 (N_18315,N_17765,N_17558);
or U18316 (N_18316,N_17855,N_17865);
nand U18317 (N_18317,N_17539,N_17848);
xnor U18318 (N_18318,N_17710,N_17885);
or U18319 (N_18319,N_17599,N_17812);
or U18320 (N_18320,N_17610,N_17736);
or U18321 (N_18321,N_17718,N_17711);
nor U18322 (N_18322,N_17807,N_17922);
nand U18323 (N_18323,N_17835,N_17648);
or U18324 (N_18324,N_17815,N_17951);
and U18325 (N_18325,N_17993,N_17819);
nand U18326 (N_18326,N_17600,N_17521);
nor U18327 (N_18327,N_17737,N_17651);
and U18328 (N_18328,N_17961,N_17792);
xnor U18329 (N_18329,N_17961,N_17936);
xnor U18330 (N_18330,N_17716,N_17906);
xnor U18331 (N_18331,N_17517,N_17876);
or U18332 (N_18332,N_17503,N_17915);
or U18333 (N_18333,N_17802,N_17678);
or U18334 (N_18334,N_17935,N_17526);
nor U18335 (N_18335,N_17573,N_17712);
nor U18336 (N_18336,N_17719,N_17653);
and U18337 (N_18337,N_17700,N_17998);
nor U18338 (N_18338,N_17553,N_17796);
nor U18339 (N_18339,N_17732,N_17621);
and U18340 (N_18340,N_17790,N_17926);
nand U18341 (N_18341,N_17935,N_17785);
xor U18342 (N_18342,N_17828,N_17534);
nor U18343 (N_18343,N_17573,N_17633);
and U18344 (N_18344,N_17746,N_17902);
or U18345 (N_18345,N_17739,N_17567);
nor U18346 (N_18346,N_17674,N_17514);
nor U18347 (N_18347,N_17547,N_17831);
or U18348 (N_18348,N_17737,N_17640);
nor U18349 (N_18349,N_17841,N_17603);
nand U18350 (N_18350,N_17836,N_17971);
or U18351 (N_18351,N_17812,N_17517);
nor U18352 (N_18352,N_17671,N_17840);
nor U18353 (N_18353,N_17780,N_17693);
and U18354 (N_18354,N_17969,N_17642);
xnor U18355 (N_18355,N_17785,N_17534);
xnor U18356 (N_18356,N_17750,N_17812);
and U18357 (N_18357,N_17699,N_17644);
xnor U18358 (N_18358,N_17831,N_17548);
nand U18359 (N_18359,N_17859,N_17523);
and U18360 (N_18360,N_17695,N_17920);
and U18361 (N_18361,N_17754,N_17846);
or U18362 (N_18362,N_17772,N_17964);
nand U18363 (N_18363,N_17552,N_17752);
nand U18364 (N_18364,N_17612,N_17531);
or U18365 (N_18365,N_17757,N_17732);
or U18366 (N_18366,N_17737,N_17709);
nand U18367 (N_18367,N_17832,N_17898);
xnor U18368 (N_18368,N_17853,N_17845);
and U18369 (N_18369,N_17585,N_17665);
and U18370 (N_18370,N_17830,N_17928);
nor U18371 (N_18371,N_17851,N_17567);
nor U18372 (N_18372,N_17720,N_17799);
or U18373 (N_18373,N_17991,N_17708);
and U18374 (N_18374,N_17864,N_17520);
and U18375 (N_18375,N_17735,N_17623);
xnor U18376 (N_18376,N_17812,N_17554);
nand U18377 (N_18377,N_17851,N_17991);
xnor U18378 (N_18378,N_17670,N_17958);
xnor U18379 (N_18379,N_17568,N_17509);
or U18380 (N_18380,N_17526,N_17774);
and U18381 (N_18381,N_17776,N_17640);
xor U18382 (N_18382,N_17870,N_17802);
xnor U18383 (N_18383,N_17735,N_17662);
nor U18384 (N_18384,N_17597,N_17845);
nand U18385 (N_18385,N_17501,N_17833);
or U18386 (N_18386,N_17855,N_17795);
nand U18387 (N_18387,N_17646,N_17960);
xnor U18388 (N_18388,N_17778,N_17826);
nor U18389 (N_18389,N_17897,N_17901);
xnor U18390 (N_18390,N_17717,N_17924);
nand U18391 (N_18391,N_17936,N_17686);
and U18392 (N_18392,N_17567,N_17531);
and U18393 (N_18393,N_17809,N_17756);
nand U18394 (N_18394,N_17550,N_17990);
nor U18395 (N_18395,N_17872,N_17935);
nand U18396 (N_18396,N_17735,N_17993);
nand U18397 (N_18397,N_17920,N_17852);
xnor U18398 (N_18398,N_17800,N_17727);
xnor U18399 (N_18399,N_17709,N_17951);
nand U18400 (N_18400,N_17900,N_17675);
and U18401 (N_18401,N_17930,N_17947);
or U18402 (N_18402,N_17781,N_17916);
nand U18403 (N_18403,N_17572,N_17993);
and U18404 (N_18404,N_17607,N_17553);
or U18405 (N_18405,N_17521,N_17554);
or U18406 (N_18406,N_17514,N_17729);
nor U18407 (N_18407,N_17681,N_17639);
or U18408 (N_18408,N_17925,N_17695);
nor U18409 (N_18409,N_17861,N_17721);
nor U18410 (N_18410,N_17665,N_17830);
nand U18411 (N_18411,N_17978,N_17891);
nand U18412 (N_18412,N_17603,N_17830);
xnor U18413 (N_18413,N_17682,N_17722);
or U18414 (N_18414,N_17906,N_17563);
and U18415 (N_18415,N_17809,N_17598);
xor U18416 (N_18416,N_17996,N_17580);
nor U18417 (N_18417,N_17534,N_17888);
and U18418 (N_18418,N_17660,N_17726);
nand U18419 (N_18419,N_17744,N_17839);
xor U18420 (N_18420,N_17762,N_17918);
nand U18421 (N_18421,N_17656,N_17688);
and U18422 (N_18422,N_17674,N_17953);
and U18423 (N_18423,N_17686,N_17636);
nand U18424 (N_18424,N_17731,N_17797);
and U18425 (N_18425,N_17906,N_17803);
xor U18426 (N_18426,N_17541,N_17824);
xnor U18427 (N_18427,N_17632,N_17561);
nand U18428 (N_18428,N_17632,N_17505);
and U18429 (N_18429,N_17644,N_17786);
xor U18430 (N_18430,N_17756,N_17629);
or U18431 (N_18431,N_17839,N_17887);
xnor U18432 (N_18432,N_17593,N_17595);
or U18433 (N_18433,N_17720,N_17915);
and U18434 (N_18434,N_17799,N_17611);
and U18435 (N_18435,N_17948,N_17782);
nand U18436 (N_18436,N_17790,N_17611);
xor U18437 (N_18437,N_17698,N_17762);
nor U18438 (N_18438,N_17864,N_17828);
nor U18439 (N_18439,N_17602,N_17932);
nor U18440 (N_18440,N_17977,N_17567);
nand U18441 (N_18441,N_17999,N_17816);
nor U18442 (N_18442,N_17815,N_17980);
or U18443 (N_18443,N_17900,N_17962);
xor U18444 (N_18444,N_17991,N_17932);
or U18445 (N_18445,N_17583,N_17677);
or U18446 (N_18446,N_17671,N_17643);
nor U18447 (N_18447,N_17529,N_17912);
or U18448 (N_18448,N_17934,N_17505);
or U18449 (N_18449,N_17845,N_17909);
or U18450 (N_18450,N_17560,N_17804);
or U18451 (N_18451,N_17862,N_17672);
nor U18452 (N_18452,N_17912,N_17574);
nor U18453 (N_18453,N_17801,N_17871);
nand U18454 (N_18454,N_17797,N_17534);
nand U18455 (N_18455,N_17793,N_17816);
xor U18456 (N_18456,N_17852,N_17524);
and U18457 (N_18457,N_17794,N_17938);
and U18458 (N_18458,N_17517,N_17819);
xor U18459 (N_18459,N_17651,N_17534);
xnor U18460 (N_18460,N_17915,N_17516);
and U18461 (N_18461,N_17767,N_17525);
and U18462 (N_18462,N_17913,N_17800);
or U18463 (N_18463,N_17630,N_17676);
or U18464 (N_18464,N_17602,N_17834);
nand U18465 (N_18465,N_17938,N_17841);
xor U18466 (N_18466,N_17613,N_17807);
or U18467 (N_18467,N_17878,N_17978);
nor U18468 (N_18468,N_17575,N_17861);
and U18469 (N_18469,N_17517,N_17803);
nand U18470 (N_18470,N_17985,N_17889);
or U18471 (N_18471,N_17960,N_17877);
xnor U18472 (N_18472,N_17691,N_17820);
nor U18473 (N_18473,N_17975,N_17786);
and U18474 (N_18474,N_17951,N_17991);
nand U18475 (N_18475,N_17656,N_17719);
xnor U18476 (N_18476,N_17555,N_17871);
and U18477 (N_18477,N_17589,N_17851);
or U18478 (N_18478,N_17931,N_17846);
nor U18479 (N_18479,N_17665,N_17599);
xnor U18480 (N_18480,N_17717,N_17500);
xnor U18481 (N_18481,N_17754,N_17648);
or U18482 (N_18482,N_17743,N_17807);
and U18483 (N_18483,N_17962,N_17743);
and U18484 (N_18484,N_17889,N_17817);
and U18485 (N_18485,N_17994,N_17690);
or U18486 (N_18486,N_17946,N_17853);
nand U18487 (N_18487,N_17832,N_17909);
xnor U18488 (N_18488,N_17928,N_17975);
xnor U18489 (N_18489,N_17920,N_17597);
nand U18490 (N_18490,N_17769,N_17974);
nor U18491 (N_18491,N_17771,N_17693);
xor U18492 (N_18492,N_17698,N_17703);
or U18493 (N_18493,N_17675,N_17581);
and U18494 (N_18494,N_17760,N_17608);
and U18495 (N_18495,N_17576,N_17954);
nand U18496 (N_18496,N_17970,N_17654);
nand U18497 (N_18497,N_17616,N_17900);
nand U18498 (N_18498,N_17773,N_17844);
xnor U18499 (N_18499,N_17640,N_17743);
nand U18500 (N_18500,N_18064,N_18012);
and U18501 (N_18501,N_18018,N_18158);
nand U18502 (N_18502,N_18395,N_18201);
and U18503 (N_18503,N_18346,N_18045);
nand U18504 (N_18504,N_18219,N_18008);
xnor U18505 (N_18505,N_18092,N_18338);
nor U18506 (N_18506,N_18388,N_18274);
nor U18507 (N_18507,N_18448,N_18104);
or U18508 (N_18508,N_18210,N_18327);
nor U18509 (N_18509,N_18399,N_18154);
or U18510 (N_18510,N_18254,N_18013);
nor U18511 (N_18511,N_18090,N_18009);
or U18512 (N_18512,N_18357,N_18417);
nor U18513 (N_18513,N_18449,N_18204);
nor U18514 (N_18514,N_18298,N_18085);
nand U18515 (N_18515,N_18451,N_18362);
nand U18516 (N_18516,N_18056,N_18324);
and U18517 (N_18517,N_18468,N_18453);
or U18518 (N_18518,N_18176,N_18003);
nand U18519 (N_18519,N_18171,N_18321);
xnor U18520 (N_18520,N_18384,N_18285);
and U18521 (N_18521,N_18134,N_18046);
and U18522 (N_18522,N_18345,N_18236);
and U18523 (N_18523,N_18063,N_18007);
nand U18524 (N_18524,N_18366,N_18398);
nor U18525 (N_18525,N_18118,N_18438);
nand U18526 (N_18526,N_18145,N_18230);
nand U18527 (N_18527,N_18169,N_18188);
xnor U18528 (N_18528,N_18223,N_18099);
and U18529 (N_18529,N_18439,N_18049);
xnor U18530 (N_18530,N_18409,N_18101);
or U18531 (N_18531,N_18253,N_18372);
or U18532 (N_18532,N_18460,N_18126);
nand U18533 (N_18533,N_18290,N_18127);
and U18534 (N_18534,N_18226,N_18100);
xor U18535 (N_18535,N_18429,N_18132);
nand U18536 (N_18536,N_18431,N_18337);
nor U18537 (N_18537,N_18463,N_18120);
xnor U18538 (N_18538,N_18222,N_18315);
xor U18539 (N_18539,N_18456,N_18237);
or U18540 (N_18540,N_18493,N_18247);
and U18541 (N_18541,N_18491,N_18263);
or U18542 (N_18542,N_18088,N_18452);
nand U18543 (N_18543,N_18148,N_18257);
and U18544 (N_18544,N_18490,N_18113);
and U18545 (N_18545,N_18306,N_18484);
nor U18546 (N_18546,N_18107,N_18352);
nor U18547 (N_18547,N_18000,N_18200);
nand U18548 (N_18548,N_18255,N_18340);
or U18549 (N_18549,N_18279,N_18144);
xnor U18550 (N_18550,N_18047,N_18386);
nand U18551 (N_18551,N_18168,N_18331);
or U18552 (N_18552,N_18270,N_18084);
nor U18553 (N_18553,N_18311,N_18062);
nand U18554 (N_18554,N_18474,N_18291);
nor U18555 (N_18555,N_18435,N_18363);
or U18556 (N_18556,N_18425,N_18173);
xor U18557 (N_18557,N_18473,N_18488);
and U18558 (N_18558,N_18241,N_18117);
nor U18559 (N_18559,N_18354,N_18050);
nand U18560 (N_18560,N_18319,N_18193);
xor U18561 (N_18561,N_18240,N_18378);
or U18562 (N_18562,N_18334,N_18192);
nand U18563 (N_18563,N_18280,N_18205);
nand U18564 (N_18564,N_18249,N_18190);
and U18565 (N_18565,N_18146,N_18479);
xnor U18566 (N_18566,N_18075,N_18137);
nand U18567 (N_18567,N_18029,N_18418);
and U18568 (N_18568,N_18339,N_18057);
nor U18569 (N_18569,N_18447,N_18037);
nor U18570 (N_18570,N_18442,N_18004);
xor U18571 (N_18571,N_18109,N_18272);
or U18572 (N_18572,N_18326,N_18404);
nand U18573 (N_18573,N_18412,N_18445);
xor U18574 (N_18574,N_18283,N_18251);
or U18575 (N_18575,N_18472,N_18314);
nand U18576 (N_18576,N_18286,N_18225);
nand U18577 (N_18577,N_18318,N_18292);
xor U18578 (N_18578,N_18248,N_18375);
and U18579 (N_18579,N_18152,N_18048);
nand U18580 (N_18580,N_18342,N_18032);
nand U18581 (N_18581,N_18061,N_18276);
xor U18582 (N_18582,N_18080,N_18069);
xor U18583 (N_18583,N_18243,N_18265);
and U18584 (N_18584,N_18440,N_18382);
nand U18585 (N_18585,N_18414,N_18264);
or U18586 (N_18586,N_18232,N_18017);
nand U18587 (N_18587,N_18024,N_18485);
or U18588 (N_18588,N_18377,N_18135);
nor U18589 (N_18589,N_18299,N_18002);
and U18590 (N_18590,N_18391,N_18028);
and U18591 (N_18591,N_18187,N_18293);
nand U18592 (N_18592,N_18358,N_18060);
and U18593 (N_18593,N_18380,N_18115);
xor U18594 (N_18594,N_18481,N_18483);
nand U18595 (N_18595,N_18437,N_18177);
nor U18596 (N_18596,N_18180,N_18071);
or U18597 (N_18597,N_18281,N_18423);
xnor U18598 (N_18598,N_18194,N_18103);
nand U18599 (N_18599,N_18245,N_18023);
and U18600 (N_18600,N_18371,N_18114);
and U18601 (N_18601,N_18203,N_18031);
nand U18602 (N_18602,N_18419,N_18221);
or U18603 (N_18603,N_18348,N_18304);
nor U18604 (N_18604,N_18268,N_18040);
xnor U18605 (N_18605,N_18016,N_18034);
nand U18606 (N_18606,N_18408,N_18343);
xnor U18607 (N_18607,N_18059,N_18446);
and U18608 (N_18608,N_18138,N_18239);
or U18609 (N_18609,N_18450,N_18095);
xnor U18610 (N_18610,N_18374,N_18305);
or U18611 (N_18611,N_18211,N_18106);
nand U18612 (N_18612,N_18153,N_18218);
and U18613 (N_18613,N_18184,N_18227);
xnor U18614 (N_18614,N_18215,N_18496);
or U18615 (N_18615,N_18191,N_18329);
nand U18616 (N_18616,N_18422,N_18436);
or U18617 (N_18617,N_18309,N_18499);
xnor U18618 (N_18618,N_18136,N_18406);
xor U18619 (N_18619,N_18228,N_18369);
xnor U18620 (N_18620,N_18310,N_18282);
and U18621 (N_18621,N_18465,N_18410);
nor U18622 (N_18622,N_18258,N_18284);
xnor U18623 (N_18623,N_18006,N_18432);
and U18624 (N_18624,N_18476,N_18396);
nor U18625 (N_18625,N_18150,N_18489);
and U18626 (N_18626,N_18252,N_18068);
nor U18627 (N_18627,N_18434,N_18128);
and U18628 (N_18628,N_18212,N_18351);
nand U18629 (N_18629,N_18010,N_18111);
xnor U18630 (N_18630,N_18238,N_18160);
nor U18631 (N_18631,N_18131,N_18196);
nor U18632 (N_18632,N_18189,N_18066);
nor U18633 (N_18633,N_18303,N_18461);
and U18634 (N_18634,N_18025,N_18022);
or U18635 (N_18635,N_18038,N_18035);
and U18636 (N_18636,N_18054,N_18108);
or U18637 (N_18637,N_18441,N_18497);
nand U18638 (N_18638,N_18297,N_18486);
nand U18639 (N_18639,N_18083,N_18147);
nand U18640 (N_18640,N_18043,N_18122);
or U18641 (N_18641,N_18149,N_18011);
nor U18642 (N_18642,N_18405,N_18403);
and U18643 (N_18643,N_18498,N_18478);
or U18644 (N_18644,N_18246,N_18373);
or U18645 (N_18645,N_18233,N_18381);
xnor U18646 (N_18646,N_18475,N_18244);
and U18647 (N_18647,N_18019,N_18026);
xor U18648 (N_18648,N_18076,N_18466);
or U18649 (N_18649,N_18454,N_18091);
nor U18650 (N_18650,N_18356,N_18387);
nor U18651 (N_18651,N_18277,N_18336);
nand U18652 (N_18652,N_18015,N_18044);
nor U18653 (N_18653,N_18287,N_18301);
and U18654 (N_18654,N_18355,N_18039);
nand U18655 (N_18655,N_18313,N_18360);
nand U18656 (N_18656,N_18294,N_18364);
nand U18657 (N_18657,N_18163,N_18141);
nor U18658 (N_18658,N_18081,N_18469);
and U18659 (N_18659,N_18457,N_18130);
nor U18660 (N_18660,N_18317,N_18462);
or U18661 (N_18661,N_18217,N_18186);
nor U18662 (N_18662,N_18089,N_18344);
nand U18663 (N_18663,N_18162,N_18413);
and U18664 (N_18664,N_18133,N_18005);
and U18665 (N_18665,N_18359,N_18269);
and U18666 (N_18666,N_18036,N_18495);
or U18667 (N_18667,N_18142,N_18295);
nor U18668 (N_18668,N_18207,N_18328);
nor U18669 (N_18669,N_18030,N_18411);
or U18670 (N_18670,N_18402,N_18021);
nor U18671 (N_18671,N_18086,N_18353);
nor U18672 (N_18672,N_18231,N_18077);
or U18673 (N_18673,N_18312,N_18459);
nor U18674 (N_18674,N_18216,N_18121);
nor U18675 (N_18675,N_18430,N_18341);
nand U18676 (N_18676,N_18444,N_18053);
nand U18677 (N_18677,N_18098,N_18392);
nor U18678 (N_18678,N_18390,N_18159);
nand U18679 (N_18679,N_18397,N_18174);
nand U18680 (N_18680,N_18234,N_18197);
nand U18681 (N_18681,N_18209,N_18259);
xnor U18682 (N_18682,N_18051,N_18323);
nand U18683 (N_18683,N_18073,N_18335);
and U18684 (N_18684,N_18494,N_18428);
nand U18685 (N_18685,N_18235,N_18361);
nor U18686 (N_18686,N_18143,N_18172);
xor U18687 (N_18687,N_18416,N_18482);
nor U18688 (N_18688,N_18480,N_18333);
nor U18689 (N_18689,N_18220,N_18202);
and U18690 (N_18690,N_18471,N_18242);
or U18691 (N_18691,N_18070,N_18112);
and U18692 (N_18692,N_18033,N_18183);
nand U18693 (N_18693,N_18376,N_18110);
and U18694 (N_18694,N_18082,N_18157);
xor U18695 (N_18695,N_18093,N_18367);
and U18696 (N_18696,N_18262,N_18266);
xor U18697 (N_18697,N_18042,N_18102);
or U18698 (N_18698,N_18020,N_18097);
and U18699 (N_18699,N_18129,N_18074);
or U18700 (N_18700,N_18167,N_18182);
and U18701 (N_18701,N_18195,N_18267);
nand U18702 (N_18702,N_18401,N_18477);
nor U18703 (N_18703,N_18316,N_18296);
and U18704 (N_18704,N_18151,N_18370);
nor U18705 (N_18705,N_18096,N_18079);
nor U18706 (N_18706,N_18058,N_18302);
and U18707 (N_18707,N_18206,N_18288);
xnor U18708 (N_18708,N_18181,N_18368);
nand U18709 (N_18709,N_18052,N_18123);
and U18710 (N_18710,N_18156,N_18213);
or U18711 (N_18711,N_18385,N_18455);
xnor U18712 (N_18712,N_18175,N_18198);
nand U18713 (N_18713,N_18426,N_18275);
nand U18714 (N_18714,N_18330,N_18307);
nor U18715 (N_18715,N_18415,N_18224);
and U18716 (N_18716,N_18055,N_18458);
nor U18717 (N_18717,N_18250,N_18420);
nand U18718 (N_18718,N_18260,N_18349);
nand U18719 (N_18719,N_18072,N_18140);
nor U18720 (N_18720,N_18400,N_18139);
or U18721 (N_18721,N_18185,N_18433);
nor U18722 (N_18722,N_18208,N_18065);
and U18723 (N_18723,N_18322,N_18350);
nand U18724 (N_18724,N_18407,N_18214);
nand U18725 (N_18725,N_18256,N_18125);
nand U18726 (N_18726,N_18424,N_18067);
and U18727 (N_18727,N_18165,N_18383);
or U18728 (N_18728,N_18393,N_18199);
nand U18729 (N_18729,N_18427,N_18271);
xnor U18730 (N_18730,N_18105,N_18464);
and U18731 (N_18731,N_18467,N_18229);
xnor U18732 (N_18732,N_18166,N_18289);
and U18733 (N_18733,N_18170,N_18041);
xnor U18734 (N_18734,N_18308,N_18001);
xnor U18735 (N_18735,N_18300,N_18087);
and U18736 (N_18736,N_18389,N_18178);
or U18737 (N_18737,N_18421,N_18325);
or U18738 (N_18738,N_18487,N_18027);
nor U18739 (N_18739,N_18332,N_18164);
and U18740 (N_18740,N_18116,N_18443);
and U18741 (N_18741,N_18379,N_18078);
nor U18742 (N_18742,N_18179,N_18155);
nand U18743 (N_18743,N_18119,N_18320);
xnor U18744 (N_18744,N_18161,N_18347);
or U18745 (N_18745,N_18273,N_18014);
xnor U18746 (N_18746,N_18278,N_18124);
or U18747 (N_18747,N_18394,N_18094);
and U18748 (N_18748,N_18492,N_18470);
nand U18749 (N_18749,N_18365,N_18261);
xnor U18750 (N_18750,N_18126,N_18334);
and U18751 (N_18751,N_18432,N_18008);
and U18752 (N_18752,N_18484,N_18303);
and U18753 (N_18753,N_18006,N_18241);
or U18754 (N_18754,N_18330,N_18192);
xor U18755 (N_18755,N_18349,N_18292);
nand U18756 (N_18756,N_18057,N_18365);
or U18757 (N_18757,N_18417,N_18051);
or U18758 (N_18758,N_18273,N_18168);
and U18759 (N_18759,N_18216,N_18400);
nand U18760 (N_18760,N_18338,N_18132);
xnor U18761 (N_18761,N_18485,N_18445);
and U18762 (N_18762,N_18221,N_18232);
xor U18763 (N_18763,N_18343,N_18319);
nand U18764 (N_18764,N_18380,N_18172);
and U18765 (N_18765,N_18076,N_18034);
and U18766 (N_18766,N_18141,N_18354);
xor U18767 (N_18767,N_18245,N_18370);
xnor U18768 (N_18768,N_18292,N_18368);
or U18769 (N_18769,N_18005,N_18249);
or U18770 (N_18770,N_18207,N_18281);
xor U18771 (N_18771,N_18412,N_18129);
or U18772 (N_18772,N_18083,N_18361);
or U18773 (N_18773,N_18015,N_18404);
or U18774 (N_18774,N_18047,N_18010);
nand U18775 (N_18775,N_18415,N_18099);
nor U18776 (N_18776,N_18358,N_18134);
or U18777 (N_18777,N_18215,N_18391);
or U18778 (N_18778,N_18006,N_18169);
and U18779 (N_18779,N_18346,N_18048);
and U18780 (N_18780,N_18262,N_18069);
nand U18781 (N_18781,N_18021,N_18295);
xor U18782 (N_18782,N_18156,N_18466);
or U18783 (N_18783,N_18390,N_18264);
nand U18784 (N_18784,N_18047,N_18195);
and U18785 (N_18785,N_18328,N_18153);
and U18786 (N_18786,N_18297,N_18458);
nand U18787 (N_18787,N_18136,N_18314);
or U18788 (N_18788,N_18078,N_18240);
nor U18789 (N_18789,N_18206,N_18414);
and U18790 (N_18790,N_18328,N_18397);
or U18791 (N_18791,N_18397,N_18147);
nor U18792 (N_18792,N_18087,N_18238);
or U18793 (N_18793,N_18415,N_18263);
or U18794 (N_18794,N_18008,N_18044);
or U18795 (N_18795,N_18418,N_18420);
and U18796 (N_18796,N_18283,N_18346);
nand U18797 (N_18797,N_18211,N_18367);
nor U18798 (N_18798,N_18337,N_18391);
xor U18799 (N_18799,N_18434,N_18046);
xor U18800 (N_18800,N_18023,N_18496);
nor U18801 (N_18801,N_18257,N_18046);
nand U18802 (N_18802,N_18076,N_18406);
nand U18803 (N_18803,N_18442,N_18008);
nor U18804 (N_18804,N_18218,N_18444);
and U18805 (N_18805,N_18262,N_18264);
xor U18806 (N_18806,N_18377,N_18348);
xnor U18807 (N_18807,N_18248,N_18407);
nor U18808 (N_18808,N_18220,N_18460);
nor U18809 (N_18809,N_18061,N_18302);
nand U18810 (N_18810,N_18490,N_18006);
and U18811 (N_18811,N_18277,N_18335);
xor U18812 (N_18812,N_18066,N_18124);
nor U18813 (N_18813,N_18231,N_18291);
or U18814 (N_18814,N_18224,N_18287);
or U18815 (N_18815,N_18448,N_18188);
xnor U18816 (N_18816,N_18357,N_18399);
xnor U18817 (N_18817,N_18424,N_18307);
and U18818 (N_18818,N_18134,N_18111);
nor U18819 (N_18819,N_18026,N_18025);
xor U18820 (N_18820,N_18447,N_18290);
and U18821 (N_18821,N_18428,N_18369);
and U18822 (N_18822,N_18120,N_18350);
xor U18823 (N_18823,N_18182,N_18419);
xnor U18824 (N_18824,N_18015,N_18158);
xor U18825 (N_18825,N_18192,N_18225);
xnor U18826 (N_18826,N_18228,N_18035);
nand U18827 (N_18827,N_18419,N_18446);
and U18828 (N_18828,N_18491,N_18122);
xor U18829 (N_18829,N_18123,N_18375);
and U18830 (N_18830,N_18022,N_18334);
xnor U18831 (N_18831,N_18412,N_18260);
xor U18832 (N_18832,N_18026,N_18219);
or U18833 (N_18833,N_18005,N_18335);
nand U18834 (N_18834,N_18246,N_18150);
nor U18835 (N_18835,N_18377,N_18292);
or U18836 (N_18836,N_18304,N_18040);
nand U18837 (N_18837,N_18235,N_18191);
or U18838 (N_18838,N_18026,N_18042);
xnor U18839 (N_18839,N_18390,N_18140);
and U18840 (N_18840,N_18265,N_18449);
and U18841 (N_18841,N_18466,N_18260);
or U18842 (N_18842,N_18078,N_18012);
xnor U18843 (N_18843,N_18379,N_18276);
or U18844 (N_18844,N_18344,N_18429);
nor U18845 (N_18845,N_18179,N_18183);
xor U18846 (N_18846,N_18038,N_18018);
nand U18847 (N_18847,N_18328,N_18084);
nor U18848 (N_18848,N_18355,N_18340);
and U18849 (N_18849,N_18353,N_18035);
nor U18850 (N_18850,N_18327,N_18288);
nand U18851 (N_18851,N_18218,N_18333);
nor U18852 (N_18852,N_18225,N_18433);
xor U18853 (N_18853,N_18040,N_18088);
nor U18854 (N_18854,N_18301,N_18283);
nand U18855 (N_18855,N_18481,N_18289);
nand U18856 (N_18856,N_18473,N_18281);
and U18857 (N_18857,N_18401,N_18151);
and U18858 (N_18858,N_18064,N_18275);
nor U18859 (N_18859,N_18349,N_18430);
nand U18860 (N_18860,N_18162,N_18110);
and U18861 (N_18861,N_18088,N_18154);
nand U18862 (N_18862,N_18456,N_18203);
nor U18863 (N_18863,N_18494,N_18137);
nand U18864 (N_18864,N_18316,N_18416);
and U18865 (N_18865,N_18193,N_18364);
and U18866 (N_18866,N_18292,N_18314);
and U18867 (N_18867,N_18290,N_18363);
nor U18868 (N_18868,N_18087,N_18472);
xor U18869 (N_18869,N_18241,N_18318);
or U18870 (N_18870,N_18284,N_18105);
xor U18871 (N_18871,N_18427,N_18192);
nand U18872 (N_18872,N_18368,N_18039);
xnor U18873 (N_18873,N_18039,N_18119);
xnor U18874 (N_18874,N_18015,N_18318);
nand U18875 (N_18875,N_18278,N_18238);
nor U18876 (N_18876,N_18409,N_18312);
and U18877 (N_18877,N_18422,N_18419);
and U18878 (N_18878,N_18237,N_18458);
and U18879 (N_18879,N_18328,N_18466);
nand U18880 (N_18880,N_18096,N_18486);
or U18881 (N_18881,N_18140,N_18399);
nor U18882 (N_18882,N_18480,N_18370);
or U18883 (N_18883,N_18131,N_18234);
nand U18884 (N_18884,N_18001,N_18014);
nand U18885 (N_18885,N_18424,N_18176);
nor U18886 (N_18886,N_18192,N_18381);
nor U18887 (N_18887,N_18242,N_18115);
xnor U18888 (N_18888,N_18317,N_18387);
and U18889 (N_18889,N_18207,N_18253);
nand U18890 (N_18890,N_18371,N_18387);
xnor U18891 (N_18891,N_18090,N_18445);
xnor U18892 (N_18892,N_18240,N_18241);
or U18893 (N_18893,N_18238,N_18334);
xor U18894 (N_18894,N_18101,N_18036);
xnor U18895 (N_18895,N_18214,N_18165);
nor U18896 (N_18896,N_18028,N_18045);
or U18897 (N_18897,N_18290,N_18175);
nor U18898 (N_18898,N_18034,N_18228);
nor U18899 (N_18899,N_18389,N_18496);
or U18900 (N_18900,N_18306,N_18273);
and U18901 (N_18901,N_18101,N_18148);
nor U18902 (N_18902,N_18461,N_18016);
nor U18903 (N_18903,N_18489,N_18052);
and U18904 (N_18904,N_18238,N_18248);
nor U18905 (N_18905,N_18117,N_18044);
and U18906 (N_18906,N_18170,N_18188);
nand U18907 (N_18907,N_18120,N_18104);
xnor U18908 (N_18908,N_18082,N_18483);
and U18909 (N_18909,N_18343,N_18335);
or U18910 (N_18910,N_18380,N_18315);
nand U18911 (N_18911,N_18340,N_18127);
nor U18912 (N_18912,N_18121,N_18477);
or U18913 (N_18913,N_18115,N_18467);
xnor U18914 (N_18914,N_18361,N_18274);
nor U18915 (N_18915,N_18309,N_18298);
or U18916 (N_18916,N_18136,N_18420);
or U18917 (N_18917,N_18462,N_18095);
and U18918 (N_18918,N_18173,N_18004);
and U18919 (N_18919,N_18484,N_18323);
or U18920 (N_18920,N_18073,N_18258);
nand U18921 (N_18921,N_18483,N_18494);
xnor U18922 (N_18922,N_18469,N_18339);
nand U18923 (N_18923,N_18022,N_18001);
nand U18924 (N_18924,N_18067,N_18476);
nand U18925 (N_18925,N_18309,N_18485);
and U18926 (N_18926,N_18199,N_18209);
or U18927 (N_18927,N_18370,N_18471);
nor U18928 (N_18928,N_18076,N_18285);
or U18929 (N_18929,N_18485,N_18126);
or U18930 (N_18930,N_18229,N_18338);
or U18931 (N_18931,N_18401,N_18270);
and U18932 (N_18932,N_18334,N_18146);
nor U18933 (N_18933,N_18047,N_18361);
and U18934 (N_18934,N_18052,N_18132);
nor U18935 (N_18935,N_18124,N_18426);
xor U18936 (N_18936,N_18118,N_18321);
nor U18937 (N_18937,N_18028,N_18312);
nand U18938 (N_18938,N_18211,N_18471);
and U18939 (N_18939,N_18476,N_18109);
and U18940 (N_18940,N_18198,N_18033);
nor U18941 (N_18941,N_18481,N_18339);
and U18942 (N_18942,N_18413,N_18326);
or U18943 (N_18943,N_18202,N_18135);
or U18944 (N_18944,N_18427,N_18300);
xnor U18945 (N_18945,N_18191,N_18201);
nand U18946 (N_18946,N_18137,N_18482);
and U18947 (N_18947,N_18109,N_18271);
nand U18948 (N_18948,N_18163,N_18134);
xnor U18949 (N_18949,N_18154,N_18307);
nor U18950 (N_18950,N_18302,N_18493);
or U18951 (N_18951,N_18056,N_18159);
xor U18952 (N_18952,N_18190,N_18306);
nand U18953 (N_18953,N_18486,N_18078);
nor U18954 (N_18954,N_18059,N_18296);
or U18955 (N_18955,N_18412,N_18168);
or U18956 (N_18956,N_18049,N_18115);
or U18957 (N_18957,N_18135,N_18102);
xnor U18958 (N_18958,N_18206,N_18493);
nor U18959 (N_18959,N_18168,N_18344);
or U18960 (N_18960,N_18298,N_18231);
or U18961 (N_18961,N_18430,N_18342);
nand U18962 (N_18962,N_18292,N_18114);
xor U18963 (N_18963,N_18351,N_18470);
xnor U18964 (N_18964,N_18189,N_18188);
nor U18965 (N_18965,N_18325,N_18486);
and U18966 (N_18966,N_18426,N_18453);
or U18967 (N_18967,N_18217,N_18023);
xor U18968 (N_18968,N_18322,N_18082);
xnor U18969 (N_18969,N_18176,N_18345);
xor U18970 (N_18970,N_18439,N_18046);
nor U18971 (N_18971,N_18330,N_18393);
xnor U18972 (N_18972,N_18217,N_18231);
and U18973 (N_18973,N_18449,N_18011);
nor U18974 (N_18974,N_18373,N_18257);
nand U18975 (N_18975,N_18496,N_18108);
and U18976 (N_18976,N_18140,N_18371);
nor U18977 (N_18977,N_18321,N_18074);
nor U18978 (N_18978,N_18145,N_18227);
or U18979 (N_18979,N_18120,N_18442);
and U18980 (N_18980,N_18177,N_18089);
xnor U18981 (N_18981,N_18367,N_18276);
or U18982 (N_18982,N_18259,N_18112);
or U18983 (N_18983,N_18153,N_18202);
nor U18984 (N_18984,N_18139,N_18492);
nand U18985 (N_18985,N_18164,N_18224);
xnor U18986 (N_18986,N_18294,N_18102);
nor U18987 (N_18987,N_18410,N_18336);
nor U18988 (N_18988,N_18268,N_18270);
and U18989 (N_18989,N_18382,N_18071);
and U18990 (N_18990,N_18131,N_18187);
xnor U18991 (N_18991,N_18474,N_18246);
xor U18992 (N_18992,N_18082,N_18460);
and U18993 (N_18993,N_18380,N_18043);
or U18994 (N_18994,N_18463,N_18155);
nor U18995 (N_18995,N_18465,N_18012);
and U18996 (N_18996,N_18414,N_18456);
nor U18997 (N_18997,N_18017,N_18245);
and U18998 (N_18998,N_18036,N_18281);
or U18999 (N_18999,N_18338,N_18415);
or U19000 (N_19000,N_18655,N_18748);
nand U19001 (N_19001,N_18561,N_18906);
nand U19002 (N_19002,N_18733,N_18889);
or U19003 (N_19003,N_18738,N_18799);
or U19004 (N_19004,N_18705,N_18949);
and U19005 (N_19005,N_18873,N_18653);
or U19006 (N_19006,N_18529,N_18820);
nand U19007 (N_19007,N_18589,N_18780);
nor U19008 (N_19008,N_18965,N_18914);
xnor U19009 (N_19009,N_18755,N_18867);
xor U19010 (N_19010,N_18781,N_18538);
nor U19011 (N_19011,N_18552,N_18893);
xnor U19012 (N_19012,N_18632,N_18710);
and U19013 (N_19013,N_18721,N_18718);
or U19014 (N_19014,N_18610,N_18711);
and U19015 (N_19015,N_18809,N_18891);
nand U19016 (N_19016,N_18551,N_18570);
and U19017 (N_19017,N_18709,N_18514);
xnor U19018 (N_19018,N_18966,N_18872);
nand U19019 (N_19019,N_18801,N_18830);
xor U19020 (N_19020,N_18640,N_18811);
or U19021 (N_19021,N_18745,N_18904);
nand U19022 (N_19022,N_18600,N_18779);
and U19023 (N_19023,N_18909,N_18505);
or U19024 (N_19024,N_18871,N_18917);
xor U19025 (N_19025,N_18870,N_18998);
nand U19026 (N_19026,N_18928,N_18983);
and U19027 (N_19027,N_18866,N_18986);
or U19028 (N_19028,N_18817,N_18598);
and U19029 (N_19029,N_18689,N_18635);
nor U19030 (N_19030,N_18800,N_18833);
or U19031 (N_19031,N_18923,N_18730);
nand U19032 (N_19032,N_18701,N_18750);
and U19033 (N_19033,N_18937,N_18592);
and U19034 (N_19034,N_18775,N_18694);
nand U19035 (N_19035,N_18731,N_18760);
nand U19036 (N_19036,N_18617,N_18548);
and U19037 (N_19037,N_18740,N_18531);
nand U19038 (N_19038,N_18968,N_18677);
xor U19039 (N_19039,N_18956,N_18619);
nand U19040 (N_19040,N_18579,N_18686);
or U19041 (N_19041,N_18615,N_18708);
or U19042 (N_19042,N_18604,N_18868);
nand U19043 (N_19043,N_18757,N_18573);
and U19044 (N_19044,N_18970,N_18588);
xor U19045 (N_19045,N_18692,N_18631);
or U19046 (N_19046,N_18771,N_18887);
nor U19047 (N_19047,N_18574,N_18674);
xnor U19048 (N_19048,N_18825,N_18854);
and U19049 (N_19049,N_18667,N_18727);
xor U19050 (N_19050,N_18941,N_18668);
or U19051 (N_19051,N_18796,N_18582);
or U19052 (N_19052,N_18784,N_18783);
or U19053 (N_19053,N_18666,N_18533);
nand U19054 (N_19054,N_18879,N_18537);
or U19055 (N_19055,N_18860,N_18554);
and U19056 (N_19056,N_18915,N_18608);
or U19057 (N_19057,N_18584,N_18850);
and U19058 (N_19058,N_18782,N_18565);
and U19059 (N_19059,N_18650,N_18752);
xor U19060 (N_19060,N_18841,N_18581);
nor U19061 (N_19061,N_18777,N_18776);
xnor U19062 (N_19062,N_18735,N_18876);
nand U19063 (N_19063,N_18616,N_18568);
xor U19064 (N_19064,N_18687,N_18996);
nand U19065 (N_19065,N_18831,N_18766);
nand U19066 (N_19066,N_18654,N_18508);
and U19067 (N_19067,N_18770,N_18555);
xnor U19068 (N_19068,N_18746,N_18989);
or U19069 (N_19069,N_18549,N_18520);
nor U19070 (N_19070,N_18648,N_18821);
and U19071 (N_19071,N_18810,N_18652);
nor U19072 (N_19072,N_18834,N_18612);
xnor U19073 (N_19073,N_18994,N_18753);
or U19074 (N_19074,N_18892,N_18678);
nor U19075 (N_19075,N_18545,N_18975);
xor U19076 (N_19076,N_18501,N_18539);
and U19077 (N_19077,N_18544,N_18806);
xor U19078 (N_19078,N_18528,N_18944);
and U19079 (N_19079,N_18706,N_18702);
nand U19080 (N_19080,N_18717,N_18913);
nand U19081 (N_19081,N_18763,N_18695);
xor U19082 (N_19082,N_18563,N_18696);
and U19083 (N_19083,N_18601,N_18855);
nor U19084 (N_19084,N_18919,N_18997);
nor U19085 (N_19085,N_18844,N_18511);
xor U19086 (N_19086,N_18703,N_18865);
nand U19087 (N_19087,N_18808,N_18874);
or U19088 (N_19088,N_18851,N_18790);
nor U19089 (N_19089,N_18691,N_18826);
or U19090 (N_19090,N_18627,N_18762);
or U19091 (N_19091,N_18973,N_18823);
or U19092 (N_19092,N_18605,N_18785);
or U19093 (N_19093,N_18591,N_18723);
nor U19094 (N_19094,N_18629,N_18829);
nor U19095 (N_19095,N_18593,N_18990);
nor U19096 (N_19096,N_18580,N_18540);
nand U19097 (N_19097,N_18902,N_18535);
nor U19098 (N_19098,N_18951,N_18964);
and U19099 (N_19099,N_18958,N_18816);
xnor U19100 (N_19100,N_18840,N_18594);
nor U19101 (N_19101,N_18530,N_18947);
nor U19102 (N_19102,N_18791,N_18517);
or U19103 (N_19103,N_18962,N_18637);
and U19104 (N_19104,N_18862,N_18832);
nor U19105 (N_19105,N_18839,N_18805);
or U19106 (N_19106,N_18999,N_18736);
nor U19107 (N_19107,N_18522,N_18575);
or U19108 (N_19108,N_18633,N_18925);
and U19109 (N_19109,N_18795,N_18901);
xnor U19110 (N_19110,N_18741,N_18908);
nor U19111 (N_19111,N_18638,N_18792);
nand U19112 (N_19112,N_18649,N_18729);
or U19113 (N_19113,N_18659,N_18747);
nor U19114 (N_19114,N_18761,N_18897);
nor U19115 (N_19115,N_18793,N_18804);
or U19116 (N_19116,N_18722,N_18642);
and U19117 (N_19117,N_18559,N_18698);
and U19118 (N_19118,N_18859,N_18662);
and U19119 (N_19119,N_18972,N_18845);
or U19120 (N_19120,N_18715,N_18773);
nand U19121 (N_19121,N_18577,N_18646);
nor U19122 (N_19122,N_18807,N_18991);
nand U19123 (N_19123,N_18607,N_18869);
or U19124 (N_19124,N_18827,N_18506);
nor U19125 (N_19125,N_18510,N_18935);
nand U19126 (N_19126,N_18883,N_18950);
nand U19127 (N_19127,N_18553,N_18948);
nor U19128 (N_19128,N_18606,N_18819);
xor U19129 (N_19129,N_18907,N_18641);
nand U19130 (N_19130,N_18571,N_18945);
and U19131 (N_19131,N_18814,N_18885);
and U19132 (N_19132,N_18982,N_18620);
or U19133 (N_19133,N_18521,N_18758);
or U19134 (N_19134,N_18957,N_18683);
nand U19135 (N_19135,N_18961,N_18894);
or U19136 (N_19136,N_18828,N_18707);
xnor U19137 (N_19137,N_18987,N_18920);
nand U19138 (N_19138,N_18926,N_18534);
or U19139 (N_19139,N_18621,N_18679);
and U19140 (N_19140,N_18967,N_18503);
nor U19141 (N_19141,N_18504,N_18794);
and U19142 (N_19142,N_18590,N_18680);
and U19143 (N_19143,N_18884,N_18734);
or U19144 (N_19144,N_18963,N_18959);
nor U19145 (N_19145,N_18712,N_18911);
or U19146 (N_19146,N_18933,N_18651);
and U19147 (N_19147,N_18670,N_18769);
nor U19148 (N_19148,N_18942,N_18671);
nor U19149 (N_19149,N_18714,N_18664);
nand U19150 (N_19150,N_18527,N_18939);
nor U19151 (N_19151,N_18512,N_18921);
nor U19152 (N_19152,N_18556,N_18737);
and U19153 (N_19153,N_18977,N_18523);
xnor U19154 (N_19154,N_18797,N_18788);
nand U19155 (N_19155,N_18971,N_18697);
nor U19156 (N_19156,N_18672,N_18960);
and U19157 (N_19157,N_18586,N_18946);
xor U19158 (N_19158,N_18665,N_18532);
xnor U19159 (N_19159,N_18720,N_18864);
xnor U19160 (N_19160,N_18849,N_18918);
nor U19161 (N_19161,N_18846,N_18836);
nor U19162 (N_19162,N_18557,N_18622);
xor U19163 (N_19163,N_18988,N_18656);
nand U19164 (N_19164,N_18881,N_18603);
and U19165 (N_19165,N_18688,N_18910);
nor U19166 (N_19166,N_18912,N_18526);
nand U19167 (N_19167,N_18838,N_18550);
and U19168 (N_19168,N_18993,N_18609);
and U19169 (N_19169,N_18562,N_18599);
nor U19170 (N_19170,N_18681,N_18974);
xnor U19171 (N_19171,N_18954,N_18931);
or U19172 (N_19172,N_18930,N_18749);
nand U19173 (N_19173,N_18660,N_18848);
and U19174 (N_19174,N_18516,N_18583);
nand U19175 (N_19175,N_18847,N_18812);
nor U19176 (N_19176,N_18518,N_18756);
nor U19177 (N_19177,N_18863,N_18818);
xor U19178 (N_19178,N_18952,N_18613);
and U19179 (N_19179,N_18700,N_18618);
and U19180 (N_19180,N_18878,N_18858);
nor U19181 (N_19181,N_18595,N_18875);
nor U19182 (N_19182,N_18566,N_18842);
or U19183 (N_19183,N_18882,N_18542);
or U19184 (N_19184,N_18713,N_18587);
and U19185 (N_19185,N_18837,N_18597);
nor U19186 (N_19186,N_18896,N_18567);
and U19187 (N_19187,N_18623,N_18934);
nor U19188 (N_19188,N_18742,N_18978);
xnor U19189 (N_19189,N_18765,N_18645);
and U19190 (N_19190,N_18772,N_18900);
nand U19191 (N_19191,N_18682,N_18732);
xor U19192 (N_19192,N_18541,N_18690);
xnor U19193 (N_19193,N_18759,N_18853);
nand U19194 (N_19194,N_18895,N_18685);
and U19195 (N_19195,N_18569,N_18509);
xnor U19196 (N_19196,N_18955,N_18886);
nor U19197 (N_19197,N_18639,N_18979);
nor U19198 (N_19198,N_18813,N_18774);
and U19199 (N_19199,N_18676,N_18976);
nor U19200 (N_19200,N_18803,N_18744);
or U19201 (N_19201,N_18513,N_18852);
and U19202 (N_19202,N_18861,N_18719);
and U19203 (N_19203,N_18940,N_18663);
xor U19204 (N_19204,N_18558,N_18980);
nand U19205 (N_19205,N_18743,N_18754);
nand U19206 (N_19206,N_18936,N_18786);
or U19207 (N_19207,N_18500,N_18572);
or U19208 (N_19208,N_18643,N_18724);
nand U19209 (N_19209,N_18798,N_18995);
xor U19210 (N_19210,N_18824,N_18630);
nor U19211 (N_19211,N_18924,N_18547);
xor U19212 (N_19212,N_18835,N_18880);
nor U19213 (N_19213,N_18673,N_18787);
or U19214 (N_19214,N_18953,N_18802);
nor U19215 (N_19215,N_18693,N_18903);
nor U19216 (N_19216,N_18644,N_18519);
and U19217 (N_19217,N_18625,N_18898);
and U19218 (N_19218,N_18647,N_18596);
nor U19219 (N_19219,N_18916,N_18525);
nor U19220 (N_19220,N_18578,N_18992);
nor U19221 (N_19221,N_18856,N_18585);
nor U19222 (N_19222,N_18927,N_18726);
nor U19223 (N_19223,N_18564,N_18768);
xnor U19224 (N_19224,N_18704,N_18657);
nor U19225 (N_19225,N_18624,N_18661);
nor U19226 (N_19226,N_18943,N_18634);
xnor U19227 (N_19227,N_18932,N_18614);
xnor U19228 (N_19228,N_18675,N_18684);
nor U19229 (N_19229,N_18611,N_18628);
and U19230 (N_19230,N_18789,N_18502);
xnor U19231 (N_19231,N_18922,N_18546);
or U19232 (N_19232,N_18981,N_18938);
nor U19233 (N_19233,N_18626,N_18843);
nor U19234 (N_19234,N_18536,N_18857);
and U19235 (N_19235,N_18669,N_18543);
nand U19236 (N_19236,N_18751,N_18888);
or U19237 (N_19237,N_18636,N_18877);
nand U19238 (N_19238,N_18764,N_18890);
xor U19239 (N_19239,N_18699,N_18515);
nor U19240 (N_19240,N_18507,N_18929);
nor U19241 (N_19241,N_18899,N_18602);
or U19242 (N_19242,N_18739,N_18767);
nand U19243 (N_19243,N_18778,N_18658);
or U19244 (N_19244,N_18728,N_18969);
nor U19245 (N_19245,N_18725,N_18985);
or U19246 (N_19246,N_18905,N_18576);
or U19247 (N_19247,N_18822,N_18524);
or U19248 (N_19248,N_18815,N_18560);
and U19249 (N_19249,N_18716,N_18984);
nor U19250 (N_19250,N_18594,N_18792);
nor U19251 (N_19251,N_18939,N_18520);
nand U19252 (N_19252,N_18696,N_18940);
nand U19253 (N_19253,N_18851,N_18856);
nand U19254 (N_19254,N_18588,N_18965);
xnor U19255 (N_19255,N_18924,N_18782);
or U19256 (N_19256,N_18891,N_18781);
xnor U19257 (N_19257,N_18861,N_18786);
and U19258 (N_19258,N_18918,N_18744);
or U19259 (N_19259,N_18726,N_18893);
nand U19260 (N_19260,N_18965,N_18506);
nor U19261 (N_19261,N_18946,N_18572);
or U19262 (N_19262,N_18745,N_18668);
xor U19263 (N_19263,N_18988,N_18762);
xor U19264 (N_19264,N_18648,N_18928);
nor U19265 (N_19265,N_18933,N_18596);
xor U19266 (N_19266,N_18672,N_18762);
or U19267 (N_19267,N_18941,N_18834);
nand U19268 (N_19268,N_18773,N_18792);
or U19269 (N_19269,N_18690,N_18550);
nand U19270 (N_19270,N_18794,N_18914);
nor U19271 (N_19271,N_18556,N_18582);
nor U19272 (N_19272,N_18507,N_18604);
nand U19273 (N_19273,N_18746,N_18888);
nor U19274 (N_19274,N_18592,N_18820);
nand U19275 (N_19275,N_18945,N_18796);
xnor U19276 (N_19276,N_18507,N_18800);
nand U19277 (N_19277,N_18502,N_18509);
and U19278 (N_19278,N_18881,N_18651);
nor U19279 (N_19279,N_18808,N_18976);
nor U19280 (N_19280,N_18567,N_18504);
and U19281 (N_19281,N_18660,N_18546);
nor U19282 (N_19282,N_18645,N_18623);
nor U19283 (N_19283,N_18998,N_18817);
or U19284 (N_19284,N_18582,N_18944);
nor U19285 (N_19285,N_18933,N_18522);
xor U19286 (N_19286,N_18930,N_18546);
xnor U19287 (N_19287,N_18789,N_18868);
and U19288 (N_19288,N_18874,N_18973);
nor U19289 (N_19289,N_18658,N_18795);
xor U19290 (N_19290,N_18518,N_18597);
nand U19291 (N_19291,N_18518,N_18637);
or U19292 (N_19292,N_18862,N_18641);
and U19293 (N_19293,N_18865,N_18902);
nor U19294 (N_19294,N_18754,N_18987);
nor U19295 (N_19295,N_18677,N_18613);
or U19296 (N_19296,N_18694,N_18553);
and U19297 (N_19297,N_18612,N_18561);
nand U19298 (N_19298,N_18989,N_18953);
nor U19299 (N_19299,N_18514,N_18710);
nand U19300 (N_19300,N_18611,N_18799);
xnor U19301 (N_19301,N_18958,N_18662);
xnor U19302 (N_19302,N_18994,N_18926);
and U19303 (N_19303,N_18861,N_18809);
and U19304 (N_19304,N_18589,N_18662);
or U19305 (N_19305,N_18716,N_18699);
xor U19306 (N_19306,N_18542,N_18876);
xnor U19307 (N_19307,N_18990,N_18510);
or U19308 (N_19308,N_18677,N_18666);
nand U19309 (N_19309,N_18892,N_18866);
xor U19310 (N_19310,N_18916,N_18781);
xnor U19311 (N_19311,N_18889,N_18509);
or U19312 (N_19312,N_18562,N_18911);
or U19313 (N_19313,N_18820,N_18564);
nand U19314 (N_19314,N_18834,N_18617);
and U19315 (N_19315,N_18731,N_18630);
nor U19316 (N_19316,N_18541,N_18755);
xnor U19317 (N_19317,N_18974,N_18592);
nor U19318 (N_19318,N_18979,N_18559);
and U19319 (N_19319,N_18784,N_18804);
xnor U19320 (N_19320,N_18887,N_18906);
or U19321 (N_19321,N_18860,N_18765);
and U19322 (N_19322,N_18760,N_18825);
nor U19323 (N_19323,N_18859,N_18824);
nand U19324 (N_19324,N_18662,N_18700);
or U19325 (N_19325,N_18509,N_18513);
or U19326 (N_19326,N_18602,N_18615);
nand U19327 (N_19327,N_18678,N_18593);
nor U19328 (N_19328,N_18606,N_18590);
nor U19329 (N_19329,N_18809,N_18662);
nor U19330 (N_19330,N_18531,N_18516);
or U19331 (N_19331,N_18705,N_18527);
xor U19332 (N_19332,N_18833,N_18510);
or U19333 (N_19333,N_18694,N_18814);
xnor U19334 (N_19334,N_18874,N_18957);
xor U19335 (N_19335,N_18562,N_18604);
nand U19336 (N_19336,N_18830,N_18821);
and U19337 (N_19337,N_18536,N_18794);
nor U19338 (N_19338,N_18998,N_18556);
xnor U19339 (N_19339,N_18518,N_18893);
xnor U19340 (N_19340,N_18770,N_18766);
and U19341 (N_19341,N_18894,N_18953);
nor U19342 (N_19342,N_18588,N_18683);
nand U19343 (N_19343,N_18840,N_18676);
nand U19344 (N_19344,N_18786,N_18927);
or U19345 (N_19345,N_18982,N_18944);
or U19346 (N_19346,N_18792,N_18874);
nand U19347 (N_19347,N_18975,N_18773);
or U19348 (N_19348,N_18740,N_18698);
or U19349 (N_19349,N_18583,N_18509);
xor U19350 (N_19350,N_18689,N_18942);
nor U19351 (N_19351,N_18625,N_18767);
nor U19352 (N_19352,N_18833,N_18748);
or U19353 (N_19353,N_18854,N_18661);
nor U19354 (N_19354,N_18644,N_18807);
nor U19355 (N_19355,N_18559,N_18800);
nand U19356 (N_19356,N_18787,N_18983);
xor U19357 (N_19357,N_18766,N_18716);
xnor U19358 (N_19358,N_18557,N_18637);
or U19359 (N_19359,N_18974,N_18883);
xnor U19360 (N_19360,N_18799,N_18604);
nand U19361 (N_19361,N_18563,N_18564);
nor U19362 (N_19362,N_18504,N_18908);
xnor U19363 (N_19363,N_18544,N_18723);
or U19364 (N_19364,N_18674,N_18756);
or U19365 (N_19365,N_18535,N_18997);
nand U19366 (N_19366,N_18891,N_18963);
nor U19367 (N_19367,N_18908,N_18687);
or U19368 (N_19368,N_18738,N_18509);
or U19369 (N_19369,N_18647,N_18844);
nor U19370 (N_19370,N_18678,N_18964);
or U19371 (N_19371,N_18831,N_18940);
nor U19372 (N_19372,N_18516,N_18860);
nand U19373 (N_19373,N_18557,N_18806);
nand U19374 (N_19374,N_18542,N_18627);
nor U19375 (N_19375,N_18637,N_18798);
nor U19376 (N_19376,N_18764,N_18900);
xnor U19377 (N_19377,N_18675,N_18996);
nor U19378 (N_19378,N_18696,N_18569);
and U19379 (N_19379,N_18560,N_18607);
and U19380 (N_19380,N_18587,N_18641);
nand U19381 (N_19381,N_18968,N_18727);
nand U19382 (N_19382,N_18951,N_18599);
nand U19383 (N_19383,N_18614,N_18664);
xor U19384 (N_19384,N_18686,N_18723);
or U19385 (N_19385,N_18655,N_18892);
xor U19386 (N_19386,N_18604,N_18595);
nand U19387 (N_19387,N_18608,N_18673);
xor U19388 (N_19388,N_18715,N_18586);
nand U19389 (N_19389,N_18752,N_18876);
nor U19390 (N_19390,N_18655,N_18526);
and U19391 (N_19391,N_18562,N_18868);
nand U19392 (N_19392,N_18729,N_18770);
nor U19393 (N_19393,N_18760,N_18514);
xnor U19394 (N_19394,N_18797,N_18538);
or U19395 (N_19395,N_18758,N_18835);
nor U19396 (N_19396,N_18682,N_18526);
and U19397 (N_19397,N_18920,N_18732);
xnor U19398 (N_19398,N_18663,N_18738);
nand U19399 (N_19399,N_18643,N_18738);
and U19400 (N_19400,N_18564,N_18755);
nor U19401 (N_19401,N_18873,N_18981);
or U19402 (N_19402,N_18793,N_18991);
or U19403 (N_19403,N_18821,N_18564);
or U19404 (N_19404,N_18768,N_18616);
nand U19405 (N_19405,N_18757,N_18512);
and U19406 (N_19406,N_18870,N_18955);
and U19407 (N_19407,N_18575,N_18508);
and U19408 (N_19408,N_18870,N_18796);
and U19409 (N_19409,N_18886,N_18694);
nand U19410 (N_19410,N_18804,N_18860);
and U19411 (N_19411,N_18872,N_18856);
and U19412 (N_19412,N_18591,N_18933);
and U19413 (N_19413,N_18855,N_18925);
nor U19414 (N_19414,N_18518,N_18790);
and U19415 (N_19415,N_18733,N_18811);
nand U19416 (N_19416,N_18559,N_18630);
or U19417 (N_19417,N_18646,N_18859);
nand U19418 (N_19418,N_18754,N_18852);
xor U19419 (N_19419,N_18659,N_18547);
xnor U19420 (N_19420,N_18822,N_18970);
nor U19421 (N_19421,N_18598,N_18628);
and U19422 (N_19422,N_18771,N_18974);
or U19423 (N_19423,N_18624,N_18723);
or U19424 (N_19424,N_18876,N_18904);
nor U19425 (N_19425,N_18717,N_18542);
and U19426 (N_19426,N_18680,N_18576);
or U19427 (N_19427,N_18985,N_18643);
and U19428 (N_19428,N_18959,N_18828);
xnor U19429 (N_19429,N_18791,N_18681);
nand U19430 (N_19430,N_18811,N_18829);
xor U19431 (N_19431,N_18768,N_18925);
nand U19432 (N_19432,N_18513,N_18687);
nand U19433 (N_19433,N_18916,N_18888);
nor U19434 (N_19434,N_18949,N_18955);
or U19435 (N_19435,N_18554,N_18605);
or U19436 (N_19436,N_18856,N_18680);
and U19437 (N_19437,N_18886,N_18582);
and U19438 (N_19438,N_18611,N_18813);
xor U19439 (N_19439,N_18973,N_18904);
xnor U19440 (N_19440,N_18860,N_18763);
and U19441 (N_19441,N_18986,N_18751);
xor U19442 (N_19442,N_18787,N_18910);
and U19443 (N_19443,N_18843,N_18612);
and U19444 (N_19444,N_18629,N_18591);
or U19445 (N_19445,N_18662,N_18607);
nor U19446 (N_19446,N_18503,N_18984);
nand U19447 (N_19447,N_18559,N_18561);
xnor U19448 (N_19448,N_18904,N_18695);
xor U19449 (N_19449,N_18515,N_18596);
nand U19450 (N_19450,N_18688,N_18532);
or U19451 (N_19451,N_18777,N_18974);
xnor U19452 (N_19452,N_18731,N_18533);
nand U19453 (N_19453,N_18881,N_18884);
or U19454 (N_19454,N_18645,N_18752);
nand U19455 (N_19455,N_18687,N_18518);
and U19456 (N_19456,N_18599,N_18518);
or U19457 (N_19457,N_18521,N_18815);
xnor U19458 (N_19458,N_18990,N_18546);
or U19459 (N_19459,N_18961,N_18949);
nand U19460 (N_19460,N_18586,N_18834);
nor U19461 (N_19461,N_18913,N_18616);
nand U19462 (N_19462,N_18825,N_18603);
nor U19463 (N_19463,N_18786,N_18926);
and U19464 (N_19464,N_18796,N_18773);
or U19465 (N_19465,N_18867,N_18609);
nor U19466 (N_19466,N_18814,N_18630);
nand U19467 (N_19467,N_18683,N_18745);
nor U19468 (N_19468,N_18559,N_18973);
nand U19469 (N_19469,N_18621,N_18564);
nor U19470 (N_19470,N_18766,N_18610);
nor U19471 (N_19471,N_18767,N_18965);
or U19472 (N_19472,N_18999,N_18703);
xor U19473 (N_19473,N_18807,N_18999);
nor U19474 (N_19474,N_18598,N_18951);
and U19475 (N_19475,N_18948,N_18537);
nor U19476 (N_19476,N_18891,N_18805);
or U19477 (N_19477,N_18608,N_18935);
nor U19478 (N_19478,N_18534,N_18817);
xnor U19479 (N_19479,N_18887,N_18510);
nor U19480 (N_19480,N_18975,N_18672);
or U19481 (N_19481,N_18849,N_18645);
or U19482 (N_19482,N_18676,N_18624);
xor U19483 (N_19483,N_18996,N_18709);
nor U19484 (N_19484,N_18805,N_18736);
or U19485 (N_19485,N_18952,N_18939);
and U19486 (N_19486,N_18907,N_18679);
xor U19487 (N_19487,N_18845,N_18867);
or U19488 (N_19488,N_18794,N_18845);
xor U19489 (N_19489,N_18998,N_18706);
xor U19490 (N_19490,N_18640,N_18962);
or U19491 (N_19491,N_18915,N_18661);
and U19492 (N_19492,N_18739,N_18806);
nor U19493 (N_19493,N_18988,N_18506);
and U19494 (N_19494,N_18788,N_18713);
nor U19495 (N_19495,N_18847,N_18537);
xnor U19496 (N_19496,N_18767,N_18967);
or U19497 (N_19497,N_18684,N_18638);
or U19498 (N_19498,N_18603,N_18901);
xor U19499 (N_19499,N_18991,N_18920);
xor U19500 (N_19500,N_19485,N_19158);
or U19501 (N_19501,N_19046,N_19028);
xor U19502 (N_19502,N_19489,N_19159);
and U19503 (N_19503,N_19470,N_19473);
nand U19504 (N_19504,N_19318,N_19432);
xnor U19505 (N_19505,N_19193,N_19382);
xor U19506 (N_19506,N_19410,N_19341);
nor U19507 (N_19507,N_19371,N_19013);
xor U19508 (N_19508,N_19217,N_19173);
xnor U19509 (N_19509,N_19228,N_19294);
nand U19510 (N_19510,N_19076,N_19398);
nor U19511 (N_19511,N_19269,N_19167);
nand U19512 (N_19512,N_19429,N_19117);
nor U19513 (N_19513,N_19062,N_19165);
or U19514 (N_19514,N_19091,N_19266);
nor U19515 (N_19515,N_19408,N_19422);
and U19516 (N_19516,N_19312,N_19149);
and U19517 (N_19517,N_19019,N_19260);
or U19518 (N_19518,N_19134,N_19478);
and U19519 (N_19519,N_19094,N_19139);
xor U19520 (N_19520,N_19163,N_19125);
xor U19521 (N_19521,N_19348,N_19477);
or U19522 (N_19522,N_19301,N_19264);
nor U19523 (N_19523,N_19457,N_19452);
or U19524 (N_19524,N_19487,N_19176);
nor U19525 (N_19525,N_19435,N_19051);
and U19526 (N_19526,N_19071,N_19211);
or U19527 (N_19527,N_19395,N_19140);
xor U19528 (N_19528,N_19138,N_19175);
xnor U19529 (N_19529,N_19048,N_19106);
nand U19530 (N_19530,N_19381,N_19237);
nor U19531 (N_19531,N_19244,N_19010);
and U19532 (N_19532,N_19388,N_19396);
nor U19533 (N_19533,N_19359,N_19327);
or U19534 (N_19534,N_19430,N_19456);
and U19535 (N_19535,N_19070,N_19251);
nor U19536 (N_19536,N_19286,N_19290);
or U19537 (N_19537,N_19417,N_19340);
and U19538 (N_19538,N_19321,N_19412);
nor U19539 (N_19539,N_19225,N_19317);
and U19540 (N_19540,N_19267,N_19349);
or U19541 (N_19541,N_19461,N_19346);
nand U19542 (N_19542,N_19399,N_19235);
nand U19543 (N_19543,N_19250,N_19099);
nand U19544 (N_19544,N_19271,N_19001);
nor U19545 (N_19545,N_19233,N_19424);
and U19546 (N_19546,N_19052,N_19316);
xor U19547 (N_19547,N_19310,N_19330);
and U19548 (N_19548,N_19389,N_19127);
nor U19549 (N_19549,N_19130,N_19224);
nor U19550 (N_19550,N_19384,N_19463);
nand U19551 (N_19551,N_19448,N_19017);
nor U19552 (N_19552,N_19328,N_19113);
xnor U19553 (N_19553,N_19356,N_19352);
nand U19554 (N_19554,N_19445,N_19009);
nand U19555 (N_19555,N_19073,N_19192);
nor U19556 (N_19556,N_19105,N_19037);
nand U19557 (N_19557,N_19377,N_19108);
or U19558 (N_19558,N_19040,N_19087);
or U19559 (N_19559,N_19164,N_19168);
or U19560 (N_19560,N_19469,N_19004);
nor U19561 (N_19561,N_19136,N_19096);
nand U19562 (N_19562,N_19287,N_19351);
and U19563 (N_19563,N_19295,N_19218);
and U19564 (N_19564,N_19495,N_19302);
or U19565 (N_19565,N_19282,N_19147);
and U19566 (N_19566,N_19097,N_19213);
nor U19567 (N_19567,N_19481,N_19026);
nand U19568 (N_19568,N_19088,N_19488);
nand U19569 (N_19569,N_19261,N_19362);
or U19570 (N_19570,N_19187,N_19298);
nand U19571 (N_19571,N_19272,N_19216);
xor U19572 (N_19572,N_19236,N_19086);
xor U19573 (N_19573,N_19016,N_19323);
xor U19574 (N_19574,N_19363,N_19032);
or U19575 (N_19575,N_19433,N_19344);
xor U19576 (N_19576,N_19102,N_19472);
or U19577 (N_19577,N_19407,N_19181);
nor U19578 (N_19578,N_19154,N_19254);
nor U19579 (N_19579,N_19190,N_19393);
xor U19580 (N_19580,N_19484,N_19077);
xor U19581 (N_19581,N_19419,N_19006);
nand U19582 (N_19582,N_19036,N_19258);
xnor U19583 (N_19583,N_19129,N_19179);
or U19584 (N_19584,N_19441,N_19305);
nand U19585 (N_19585,N_19111,N_19297);
nor U19586 (N_19586,N_19423,N_19379);
nor U19587 (N_19587,N_19189,N_19355);
and U19588 (N_19588,N_19437,N_19372);
nor U19589 (N_19589,N_19119,N_19438);
nand U19590 (N_19590,N_19132,N_19498);
xor U19591 (N_19591,N_19378,N_19023);
or U19592 (N_19592,N_19171,N_19322);
xnor U19593 (N_19593,N_19338,N_19057);
or U19594 (N_19594,N_19146,N_19199);
xnor U19595 (N_19595,N_19143,N_19198);
and U19596 (N_19596,N_19243,N_19131);
and U19597 (N_19597,N_19162,N_19436);
nand U19598 (N_19598,N_19034,N_19405);
nand U19599 (N_19599,N_19380,N_19003);
nand U19600 (N_19600,N_19059,N_19263);
nand U19601 (N_19601,N_19103,N_19428);
nand U19602 (N_19602,N_19063,N_19242);
xnor U19603 (N_19603,N_19008,N_19358);
or U19604 (N_19604,N_19247,N_19311);
or U19605 (N_19605,N_19081,N_19033);
and U19606 (N_19606,N_19151,N_19259);
or U19607 (N_19607,N_19169,N_19174);
or U19608 (N_19608,N_19390,N_19232);
nor U19609 (N_19609,N_19234,N_19018);
nor U19610 (N_19610,N_19084,N_19426);
and U19611 (N_19611,N_19369,N_19208);
or U19612 (N_19612,N_19241,N_19279);
or U19613 (N_19613,N_19256,N_19172);
nor U19614 (N_19614,N_19126,N_19475);
nor U19615 (N_19615,N_19112,N_19280);
or U19616 (N_19616,N_19166,N_19462);
nand U19617 (N_19617,N_19354,N_19201);
xor U19618 (N_19618,N_19226,N_19152);
nand U19619 (N_19619,N_19066,N_19420);
nor U19620 (N_19620,N_19060,N_19289);
nor U19621 (N_19621,N_19157,N_19220);
xnor U19622 (N_19622,N_19347,N_19342);
nand U19623 (N_19623,N_19000,N_19418);
or U19624 (N_19624,N_19067,N_19496);
or U19625 (N_19625,N_19474,N_19148);
and U19626 (N_19626,N_19205,N_19494);
and U19627 (N_19627,N_19153,N_19367);
or U19628 (N_19628,N_19252,N_19011);
xor U19629 (N_19629,N_19265,N_19442);
nand U19630 (N_19630,N_19391,N_19101);
nand U19631 (N_19631,N_19024,N_19121);
nor U19632 (N_19632,N_19497,N_19303);
and U19633 (N_19633,N_19089,N_19299);
nor U19634 (N_19634,N_19184,N_19434);
nand U19635 (N_19635,N_19325,N_19332);
xor U19636 (N_19636,N_19118,N_19015);
or U19637 (N_19637,N_19392,N_19161);
nor U19638 (N_19638,N_19383,N_19284);
nor U19639 (N_19639,N_19386,N_19090);
and U19640 (N_19640,N_19406,N_19203);
or U19641 (N_19641,N_19002,N_19313);
or U19642 (N_19642,N_19042,N_19361);
and U19643 (N_19643,N_19466,N_19160);
xnor U19644 (N_19644,N_19409,N_19292);
nand U19645 (N_19645,N_19079,N_19020);
or U19646 (N_19646,N_19116,N_19476);
nor U19647 (N_19647,N_19440,N_19337);
nand U19648 (N_19648,N_19444,N_19012);
and U19649 (N_19649,N_19219,N_19025);
and U19650 (N_19650,N_19450,N_19364);
and U19651 (N_19651,N_19068,N_19182);
nor U19652 (N_19652,N_19183,N_19123);
nand U19653 (N_19653,N_19209,N_19464);
xnor U19654 (N_19654,N_19030,N_19291);
and U19655 (N_19655,N_19155,N_19145);
or U19656 (N_19656,N_19044,N_19360);
xor U19657 (N_19657,N_19465,N_19376);
or U19658 (N_19658,N_19230,N_19370);
or U19659 (N_19659,N_19069,N_19180);
nor U19660 (N_19660,N_19082,N_19142);
nor U19661 (N_19661,N_19221,N_19207);
xnor U19662 (N_19662,N_19061,N_19331);
or U19663 (N_19663,N_19270,N_19401);
and U19664 (N_19664,N_19306,N_19246);
nor U19665 (N_19665,N_19093,N_19482);
nand U19666 (N_19666,N_19064,N_19309);
xnor U19667 (N_19667,N_19277,N_19447);
xor U19668 (N_19668,N_19065,N_19202);
nor U19669 (N_19669,N_19114,N_19204);
and U19670 (N_19670,N_19137,N_19439);
nand U19671 (N_19671,N_19320,N_19459);
nand U19672 (N_19672,N_19120,N_19479);
xor U19673 (N_19673,N_19185,N_19486);
or U19674 (N_19674,N_19215,N_19248);
and U19675 (N_19675,N_19324,N_19038);
nor U19676 (N_19676,N_19304,N_19490);
and U19677 (N_19677,N_19308,N_19385);
nand U19678 (N_19678,N_19210,N_19483);
nand U19679 (N_19679,N_19333,N_19335);
xnor U19680 (N_19680,N_19115,N_19275);
xnor U19681 (N_19681,N_19245,N_19005);
xnor U19682 (N_19682,N_19449,N_19411);
xor U19683 (N_19683,N_19387,N_19098);
and U19684 (N_19684,N_19083,N_19056);
nand U19685 (N_19685,N_19281,N_19413);
and U19686 (N_19686,N_19455,N_19365);
xor U19687 (N_19687,N_19283,N_19339);
or U19688 (N_19688,N_19239,N_19334);
or U19689 (N_19689,N_19049,N_19357);
nor U19690 (N_19690,N_19415,N_19078);
and U19691 (N_19691,N_19039,N_19336);
nand U19692 (N_19692,N_19054,N_19374);
nor U19693 (N_19693,N_19041,N_19343);
nor U19694 (N_19694,N_19350,N_19454);
or U19695 (N_19695,N_19231,N_19249);
and U19696 (N_19696,N_19085,N_19326);
nor U19697 (N_19697,N_19397,N_19402);
and U19698 (N_19698,N_19141,N_19100);
or U19699 (N_19699,N_19196,N_19194);
nand U19700 (N_19700,N_19460,N_19022);
nand U19701 (N_19701,N_19253,N_19451);
or U19702 (N_19702,N_19471,N_19414);
or U19703 (N_19703,N_19373,N_19047);
and U19704 (N_19704,N_19446,N_19135);
nand U19705 (N_19705,N_19007,N_19421);
xnor U19706 (N_19706,N_19206,N_19195);
or U19707 (N_19707,N_19427,N_19031);
nor U19708 (N_19708,N_19014,N_19050);
nor U19709 (N_19709,N_19345,N_19431);
nand U19710 (N_19710,N_19214,N_19133);
and U19711 (N_19711,N_19107,N_19240);
and U19712 (N_19712,N_19296,N_19197);
and U19713 (N_19713,N_19403,N_19109);
nor U19714 (N_19714,N_19262,N_19178);
nor U19715 (N_19715,N_19110,N_19467);
xor U19716 (N_19716,N_19400,N_19074);
and U19717 (N_19717,N_19186,N_19453);
nand U19718 (N_19718,N_19425,N_19315);
or U19719 (N_19719,N_19375,N_19212);
xnor U19720 (N_19720,N_19200,N_19300);
and U19721 (N_19721,N_19124,N_19314);
nor U19722 (N_19722,N_19368,N_19353);
xnor U19723 (N_19723,N_19035,N_19122);
nor U19724 (N_19724,N_19072,N_19499);
xor U19725 (N_19725,N_19053,N_19170);
or U19726 (N_19726,N_19255,N_19319);
nor U19727 (N_19727,N_19043,N_19492);
nand U19728 (N_19728,N_19329,N_19480);
or U19729 (N_19729,N_19095,N_19055);
and U19730 (N_19730,N_19257,N_19104);
or U19731 (N_19731,N_19227,N_19223);
and U19732 (N_19732,N_19443,N_19128);
or U19733 (N_19733,N_19491,N_19222);
or U19734 (N_19734,N_19144,N_19273);
and U19735 (N_19735,N_19027,N_19493);
or U19736 (N_19736,N_19416,N_19092);
xnor U19737 (N_19737,N_19029,N_19229);
nand U19738 (N_19738,N_19150,N_19191);
nor U19739 (N_19739,N_19080,N_19276);
or U19740 (N_19740,N_19177,N_19278);
nand U19741 (N_19741,N_19045,N_19058);
nor U19742 (N_19742,N_19021,N_19188);
xnor U19743 (N_19743,N_19156,N_19268);
nand U19744 (N_19744,N_19468,N_19075);
or U19745 (N_19745,N_19288,N_19274);
nand U19746 (N_19746,N_19238,N_19293);
nor U19747 (N_19747,N_19404,N_19285);
nand U19748 (N_19748,N_19458,N_19307);
and U19749 (N_19749,N_19366,N_19394);
and U19750 (N_19750,N_19250,N_19356);
or U19751 (N_19751,N_19450,N_19245);
nand U19752 (N_19752,N_19230,N_19431);
or U19753 (N_19753,N_19224,N_19037);
or U19754 (N_19754,N_19067,N_19490);
or U19755 (N_19755,N_19175,N_19070);
or U19756 (N_19756,N_19448,N_19455);
or U19757 (N_19757,N_19433,N_19479);
xor U19758 (N_19758,N_19409,N_19150);
nor U19759 (N_19759,N_19315,N_19399);
nor U19760 (N_19760,N_19196,N_19313);
xnor U19761 (N_19761,N_19346,N_19269);
xor U19762 (N_19762,N_19030,N_19188);
or U19763 (N_19763,N_19466,N_19166);
nand U19764 (N_19764,N_19233,N_19040);
and U19765 (N_19765,N_19077,N_19135);
and U19766 (N_19766,N_19070,N_19322);
xnor U19767 (N_19767,N_19260,N_19281);
or U19768 (N_19768,N_19448,N_19344);
xnor U19769 (N_19769,N_19419,N_19066);
xnor U19770 (N_19770,N_19389,N_19272);
or U19771 (N_19771,N_19253,N_19236);
xnor U19772 (N_19772,N_19430,N_19480);
xor U19773 (N_19773,N_19006,N_19498);
and U19774 (N_19774,N_19446,N_19406);
nand U19775 (N_19775,N_19425,N_19126);
and U19776 (N_19776,N_19452,N_19461);
or U19777 (N_19777,N_19294,N_19044);
nor U19778 (N_19778,N_19136,N_19007);
and U19779 (N_19779,N_19399,N_19226);
xor U19780 (N_19780,N_19422,N_19203);
nand U19781 (N_19781,N_19085,N_19442);
nand U19782 (N_19782,N_19406,N_19368);
or U19783 (N_19783,N_19076,N_19311);
xnor U19784 (N_19784,N_19423,N_19041);
nand U19785 (N_19785,N_19497,N_19487);
and U19786 (N_19786,N_19012,N_19445);
nand U19787 (N_19787,N_19233,N_19446);
nand U19788 (N_19788,N_19395,N_19086);
and U19789 (N_19789,N_19268,N_19492);
xor U19790 (N_19790,N_19134,N_19027);
xor U19791 (N_19791,N_19183,N_19250);
nor U19792 (N_19792,N_19172,N_19478);
and U19793 (N_19793,N_19269,N_19126);
or U19794 (N_19794,N_19193,N_19024);
nor U19795 (N_19795,N_19406,N_19340);
xor U19796 (N_19796,N_19267,N_19379);
xnor U19797 (N_19797,N_19239,N_19484);
nand U19798 (N_19798,N_19447,N_19484);
nand U19799 (N_19799,N_19216,N_19016);
nor U19800 (N_19800,N_19107,N_19025);
xnor U19801 (N_19801,N_19402,N_19021);
and U19802 (N_19802,N_19450,N_19376);
xnor U19803 (N_19803,N_19424,N_19409);
or U19804 (N_19804,N_19483,N_19348);
nor U19805 (N_19805,N_19401,N_19097);
or U19806 (N_19806,N_19487,N_19111);
and U19807 (N_19807,N_19421,N_19453);
and U19808 (N_19808,N_19416,N_19479);
nand U19809 (N_19809,N_19289,N_19246);
or U19810 (N_19810,N_19213,N_19289);
nor U19811 (N_19811,N_19123,N_19364);
and U19812 (N_19812,N_19401,N_19457);
xnor U19813 (N_19813,N_19214,N_19384);
and U19814 (N_19814,N_19289,N_19459);
nor U19815 (N_19815,N_19032,N_19106);
and U19816 (N_19816,N_19203,N_19415);
xor U19817 (N_19817,N_19479,N_19115);
xnor U19818 (N_19818,N_19171,N_19415);
nand U19819 (N_19819,N_19134,N_19290);
nand U19820 (N_19820,N_19000,N_19156);
and U19821 (N_19821,N_19101,N_19095);
nand U19822 (N_19822,N_19129,N_19481);
xnor U19823 (N_19823,N_19082,N_19190);
nand U19824 (N_19824,N_19495,N_19246);
xnor U19825 (N_19825,N_19048,N_19350);
nor U19826 (N_19826,N_19217,N_19223);
nand U19827 (N_19827,N_19431,N_19341);
nand U19828 (N_19828,N_19268,N_19389);
nor U19829 (N_19829,N_19420,N_19335);
xnor U19830 (N_19830,N_19257,N_19359);
xnor U19831 (N_19831,N_19385,N_19195);
nand U19832 (N_19832,N_19429,N_19299);
and U19833 (N_19833,N_19137,N_19025);
or U19834 (N_19834,N_19119,N_19083);
or U19835 (N_19835,N_19207,N_19354);
and U19836 (N_19836,N_19105,N_19397);
xnor U19837 (N_19837,N_19143,N_19286);
or U19838 (N_19838,N_19433,N_19162);
and U19839 (N_19839,N_19254,N_19384);
and U19840 (N_19840,N_19280,N_19307);
or U19841 (N_19841,N_19039,N_19379);
nor U19842 (N_19842,N_19433,N_19280);
xor U19843 (N_19843,N_19458,N_19424);
xnor U19844 (N_19844,N_19461,N_19476);
xor U19845 (N_19845,N_19464,N_19407);
nand U19846 (N_19846,N_19159,N_19003);
nor U19847 (N_19847,N_19440,N_19471);
or U19848 (N_19848,N_19110,N_19185);
xor U19849 (N_19849,N_19017,N_19173);
xor U19850 (N_19850,N_19235,N_19211);
or U19851 (N_19851,N_19478,N_19186);
xnor U19852 (N_19852,N_19049,N_19170);
nand U19853 (N_19853,N_19481,N_19349);
xor U19854 (N_19854,N_19406,N_19020);
xor U19855 (N_19855,N_19451,N_19290);
and U19856 (N_19856,N_19457,N_19149);
and U19857 (N_19857,N_19032,N_19149);
nor U19858 (N_19858,N_19386,N_19431);
nor U19859 (N_19859,N_19308,N_19089);
nand U19860 (N_19860,N_19269,N_19320);
and U19861 (N_19861,N_19443,N_19359);
and U19862 (N_19862,N_19323,N_19291);
nand U19863 (N_19863,N_19109,N_19112);
and U19864 (N_19864,N_19327,N_19256);
nand U19865 (N_19865,N_19034,N_19443);
xor U19866 (N_19866,N_19388,N_19248);
nand U19867 (N_19867,N_19112,N_19151);
nor U19868 (N_19868,N_19468,N_19231);
nor U19869 (N_19869,N_19282,N_19214);
xor U19870 (N_19870,N_19161,N_19417);
and U19871 (N_19871,N_19367,N_19166);
nor U19872 (N_19872,N_19415,N_19128);
nor U19873 (N_19873,N_19298,N_19202);
nor U19874 (N_19874,N_19028,N_19135);
nor U19875 (N_19875,N_19179,N_19288);
nor U19876 (N_19876,N_19349,N_19484);
and U19877 (N_19877,N_19348,N_19037);
xnor U19878 (N_19878,N_19375,N_19255);
xnor U19879 (N_19879,N_19337,N_19457);
xnor U19880 (N_19880,N_19055,N_19365);
nor U19881 (N_19881,N_19097,N_19098);
nand U19882 (N_19882,N_19136,N_19004);
xnor U19883 (N_19883,N_19341,N_19214);
xor U19884 (N_19884,N_19422,N_19048);
nor U19885 (N_19885,N_19182,N_19463);
xor U19886 (N_19886,N_19098,N_19163);
xnor U19887 (N_19887,N_19153,N_19328);
or U19888 (N_19888,N_19219,N_19169);
or U19889 (N_19889,N_19008,N_19062);
nand U19890 (N_19890,N_19214,N_19467);
nand U19891 (N_19891,N_19418,N_19174);
or U19892 (N_19892,N_19075,N_19359);
or U19893 (N_19893,N_19270,N_19241);
nand U19894 (N_19894,N_19017,N_19377);
or U19895 (N_19895,N_19388,N_19301);
nor U19896 (N_19896,N_19227,N_19136);
nor U19897 (N_19897,N_19436,N_19170);
nor U19898 (N_19898,N_19259,N_19390);
and U19899 (N_19899,N_19191,N_19445);
and U19900 (N_19900,N_19485,N_19236);
nor U19901 (N_19901,N_19444,N_19306);
nor U19902 (N_19902,N_19046,N_19467);
nand U19903 (N_19903,N_19210,N_19041);
and U19904 (N_19904,N_19486,N_19203);
nor U19905 (N_19905,N_19324,N_19437);
nand U19906 (N_19906,N_19411,N_19393);
or U19907 (N_19907,N_19399,N_19254);
nor U19908 (N_19908,N_19068,N_19084);
xor U19909 (N_19909,N_19000,N_19391);
xor U19910 (N_19910,N_19023,N_19325);
or U19911 (N_19911,N_19141,N_19182);
nand U19912 (N_19912,N_19373,N_19403);
or U19913 (N_19913,N_19285,N_19044);
and U19914 (N_19914,N_19342,N_19236);
nor U19915 (N_19915,N_19028,N_19057);
xor U19916 (N_19916,N_19123,N_19421);
xnor U19917 (N_19917,N_19207,N_19355);
xnor U19918 (N_19918,N_19126,N_19421);
or U19919 (N_19919,N_19206,N_19277);
xnor U19920 (N_19920,N_19208,N_19066);
or U19921 (N_19921,N_19365,N_19021);
xnor U19922 (N_19922,N_19255,N_19391);
or U19923 (N_19923,N_19485,N_19288);
nor U19924 (N_19924,N_19037,N_19029);
nand U19925 (N_19925,N_19067,N_19031);
and U19926 (N_19926,N_19180,N_19295);
nor U19927 (N_19927,N_19222,N_19246);
and U19928 (N_19928,N_19098,N_19266);
nand U19929 (N_19929,N_19341,N_19203);
or U19930 (N_19930,N_19102,N_19465);
xnor U19931 (N_19931,N_19243,N_19188);
xnor U19932 (N_19932,N_19201,N_19260);
nand U19933 (N_19933,N_19299,N_19289);
nor U19934 (N_19934,N_19376,N_19155);
and U19935 (N_19935,N_19149,N_19214);
nand U19936 (N_19936,N_19123,N_19184);
xor U19937 (N_19937,N_19244,N_19452);
or U19938 (N_19938,N_19322,N_19032);
or U19939 (N_19939,N_19411,N_19350);
nor U19940 (N_19940,N_19382,N_19128);
nand U19941 (N_19941,N_19495,N_19152);
xor U19942 (N_19942,N_19175,N_19386);
nand U19943 (N_19943,N_19316,N_19419);
nand U19944 (N_19944,N_19008,N_19223);
nor U19945 (N_19945,N_19499,N_19270);
and U19946 (N_19946,N_19009,N_19190);
and U19947 (N_19947,N_19395,N_19438);
xnor U19948 (N_19948,N_19179,N_19035);
and U19949 (N_19949,N_19334,N_19084);
nor U19950 (N_19950,N_19193,N_19278);
nand U19951 (N_19951,N_19340,N_19221);
nor U19952 (N_19952,N_19208,N_19430);
nand U19953 (N_19953,N_19172,N_19236);
or U19954 (N_19954,N_19301,N_19176);
nor U19955 (N_19955,N_19430,N_19288);
nor U19956 (N_19956,N_19247,N_19417);
xnor U19957 (N_19957,N_19383,N_19167);
nor U19958 (N_19958,N_19258,N_19158);
nor U19959 (N_19959,N_19458,N_19342);
nor U19960 (N_19960,N_19359,N_19438);
or U19961 (N_19961,N_19429,N_19392);
or U19962 (N_19962,N_19409,N_19241);
nand U19963 (N_19963,N_19294,N_19156);
and U19964 (N_19964,N_19127,N_19053);
xnor U19965 (N_19965,N_19213,N_19071);
nor U19966 (N_19966,N_19225,N_19439);
and U19967 (N_19967,N_19210,N_19361);
xor U19968 (N_19968,N_19435,N_19343);
nand U19969 (N_19969,N_19284,N_19462);
nand U19970 (N_19970,N_19000,N_19492);
nand U19971 (N_19971,N_19203,N_19026);
and U19972 (N_19972,N_19047,N_19008);
or U19973 (N_19973,N_19419,N_19377);
xor U19974 (N_19974,N_19265,N_19483);
and U19975 (N_19975,N_19326,N_19409);
xnor U19976 (N_19976,N_19036,N_19084);
xor U19977 (N_19977,N_19243,N_19013);
nor U19978 (N_19978,N_19484,N_19007);
and U19979 (N_19979,N_19094,N_19117);
nand U19980 (N_19980,N_19357,N_19306);
nor U19981 (N_19981,N_19142,N_19208);
nor U19982 (N_19982,N_19195,N_19430);
or U19983 (N_19983,N_19212,N_19246);
nand U19984 (N_19984,N_19456,N_19009);
nand U19985 (N_19985,N_19225,N_19212);
nand U19986 (N_19986,N_19350,N_19125);
nand U19987 (N_19987,N_19093,N_19242);
nand U19988 (N_19988,N_19483,N_19174);
or U19989 (N_19989,N_19353,N_19049);
xnor U19990 (N_19990,N_19079,N_19333);
nand U19991 (N_19991,N_19379,N_19326);
xnor U19992 (N_19992,N_19112,N_19376);
xnor U19993 (N_19993,N_19314,N_19243);
or U19994 (N_19994,N_19277,N_19453);
and U19995 (N_19995,N_19211,N_19216);
and U19996 (N_19996,N_19335,N_19070);
and U19997 (N_19997,N_19162,N_19153);
nor U19998 (N_19998,N_19409,N_19412);
xnor U19999 (N_19999,N_19152,N_19305);
or UO_0 (O_0,N_19888,N_19910);
xnor UO_1 (O_1,N_19653,N_19514);
nand UO_2 (O_2,N_19786,N_19914);
xnor UO_3 (O_3,N_19646,N_19681);
or UO_4 (O_4,N_19995,N_19993);
and UO_5 (O_5,N_19637,N_19569);
nor UO_6 (O_6,N_19658,N_19610);
or UO_7 (O_7,N_19751,N_19544);
nor UO_8 (O_8,N_19567,N_19505);
xor UO_9 (O_9,N_19853,N_19813);
nor UO_10 (O_10,N_19971,N_19986);
nand UO_11 (O_11,N_19509,N_19873);
and UO_12 (O_12,N_19898,N_19600);
xnor UO_13 (O_13,N_19792,N_19860);
nor UO_14 (O_14,N_19584,N_19948);
and UO_15 (O_15,N_19533,N_19761);
nand UO_16 (O_16,N_19749,N_19589);
xnor UO_17 (O_17,N_19985,N_19883);
nand UO_18 (O_18,N_19691,N_19889);
nand UO_19 (O_19,N_19906,N_19818);
xor UO_20 (O_20,N_19819,N_19542);
nor UO_21 (O_21,N_19711,N_19679);
or UO_22 (O_22,N_19964,N_19942);
and UO_23 (O_23,N_19540,N_19790);
and UO_24 (O_24,N_19545,N_19603);
and UO_25 (O_25,N_19688,N_19904);
nand UO_26 (O_26,N_19619,N_19537);
or UO_27 (O_27,N_19586,N_19946);
nor UO_28 (O_28,N_19758,N_19922);
nor UO_29 (O_29,N_19908,N_19754);
nor UO_30 (O_30,N_19686,N_19780);
xnor UO_31 (O_31,N_19661,N_19793);
or UO_32 (O_32,N_19972,N_19809);
and UO_33 (O_33,N_19718,N_19650);
xnor UO_34 (O_34,N_19725,N_19893);
xnor UO_35 (O_35,N_19755,N_19775);
nand UO_36 (O_36,N_19601,N_19848);
and UO_37 (O_37,N_19762,N_19909);
xor UO_38 (O_38,N_19821,N_19998);
and UO_39 (O_39,N_19708,N_19732);
or UO_40 (O_40,N_19713,N_19735);
nand UO_41 (O_41,N_19785,N_19625);
nand UO_42 (O_42,N_19894,N_19561);
or UO_43 (O_43,N_19705,N_19825);
and UO_44 (O_44,N_19714,N_19842);
xnor UO_45 (O_45,N_19820,N_19823);
nand UO_46 (O_46,N_19558,N_19668);
or UO_47 (O_47,N_19741,N_19866);
or UO_48 (O_48,N_19945,N_19716);
nor UO_49 (O_49,N_19845,N_19768);
nor UO_50 (O_50,N_19683,N_19698);
or UO_51 (O_51,N_19521,N_19938);
and UO_52 (O_52,N_19664,N_19773);
and UO_53 (O_53,N_19847,N_19506);
nor UO_54 (O_54,N_19512,N_19885);
nand UO_55 (O_55,N_19608,N_19666);
nor UO_56 (O_56,N_19856,N_19704);
and UO_57 (O_57,N_19648,N_19837);
nor UO_58 (O_58,N_19543,N_19634);
nand UO_59 (O_59,N_19899,N_19674);
or UO_60 (O_60,N_19526,N_19555);
nor UO_61 (O_61,N_19576,N_19535);
nor UO_62 (O_62,N_19726,N_19877);
xor UO_63 (O_63,N_19811,N_19911);
or UO_64 (O_64,N_19531,N_19587);
or UO_65 (O_65,N_19654,N_19760);
xor UO_66 (O_66,N_19534,N_19801);
nor UO_67 (O_67,N_19816,N_19772);
and UO_68 (O_68,N_19722,N_19682);
and UO_69 (O_69,N_19748,N_19616);
xnor UO_70 (O_70,N_19869,N_19992);
and UO_71 (O_71,N_19947,N_19644);
xnor UO_72 (O_72,N_19886,N_19835);
xor UO_73 (O_73,N_19670,N_19795);
or UO_74 (O_74,N_19783,N_19578);
and UO_75 (O_75,N_19671,N_19913);
nand UO_76 (O_76,N_19730,N_19902);
nor UO_77 (O_77,N_19511,N_19936);
or UO_78 (O_78,N_19797,N_19896);
and UO_79 (O_79,N_19800,N_19782);
nand UO_80 (O_80,N_19943,N_19662);
nand UO_81 (O_81,N_19974,N_19724);
nand UO_82 (O_82,N_19846,N_19685);
nand UO_83 (O_83,N_19776,N_19630);
and UO_84 (O_84,N_19779,N_19996);
nand UO_85 (O_85,N_19639,N_19852);
and UO_86 (O_86,N_19887,N_19721);
nand UO_87 (O_87,N_19590,N_19565);
nor UO_88 (O_88,N_19568,N_19524);
nand UO_89 (O_89,N_19629,N_19541);
nor UO_90 (O_90,N_19609,N_19857);
nand UO_91 (O_91,N_19753,N_19982);
or UO_92 (O_92,N_19833,N_19752);
nor UO_93 (O_93,N_19960,N_19638);
nand UO_94 (O_94,N_19743,N_19504);
nor UO_95 (O_95,N_19966,N_19728);
or UO_96 (O_96,N_19593,N_19941);
or UO_97 (O_97,N_19777,N_19851);
or UO_98 (O_98,N_19962,N_19763);
and UO_99 (O_99,N_19613,N_19742);
nor UO_100 (O_100,N_19834,N_19766);
xnor UO_101 (O_101,N_19502,N_19510);
nor UO_102 (O_102,N_19710,N_19740);
and UO_103 (O_103,N_19917,N_19518);
nand UO_104 (O_104,N_19759,N_19604);
xor UO_105 (O_105,N_19921,N_19810);
or UO_106 (O_106,N_19627,N_19689);
or UO_107 (O_107,N_19756,N_19802);
and UO_108 (O_108,N_19861,N_19583);
or UO_109 (O_109,N_19932,N_19920);
or UO_110 (O_110,N_19701,N_19709);
and UO_111 (O_111,N_19696,N_19767);
and UO_112 (O_112,N_19699,N_19592);
or UO_113 (O_113,N_19642,N_19977);
nand UO_114 (O_114,N_19678,N_19965);
nor UO_115 (O_115,N_19874,N_19665);
nand UO_116 (O_116,N_19529,N_19539);
nand UO_117 (O_117,N_19607,N_19633);
xnor UO_118 (O_118,N_19798,N_19680);
and UO_119 (O_119,N_19647,N_19612);
nor UO_120 (O_120,N_19657,N_19547);
xor UO_121 (O_121,N_19826,N_19649);
nor UO_122 (O_122,N_19525,N_19538);
nand UO_123 (O_123,N_19978,N_19515);
or UO_124 (O_124,N_19684,N_19746);
and UO_125 (O_125,N_19702,N_19892);
nand UO_126 (O_126,N_19931,N_19553);
nor UO_127 (O_127,N_19994,N_19879);
and UO_128 (O_128,N_19831,N_19791);
nor UO_129 (O_129,N_19757,N_19929);
nor UO_130 (O_130,N_19789,N_19765);
xor UO_131 (O_131,N_19636,N_19912);
or UO_132 (O_132,N_19617,N_19803);
nand UO_133 (O_133,N_19675,N_19882);
or UO_134 (O_134,N_19585,N_19829);
nand UO_135 (O_135,N_19573,N_19855);
nand UO_136 (O_136,N_19717,N_19700);
and UO_137 (O_137,N_19527,N_19915);
or UO_138 (O_138,N_19643,N_19991);
xnor UO_139 (O_139,N_19673,N_19564);
or UO_140 (O_140,N_19507,N_19796);
nor UO_141 (O_141,N_19927,N_19687);
or UO_142 (O_142,N_19623,N_19552);
nor UO_143 (O_143,N_19631,N_19554);
xor UO_144 (O_144,N_19595,N_19695);
xnor UO_145 (O_145,N_19738,N_19919);
nor UO_146 (O_146,N_19975,N_19729);
nor UO_147 (O_147,N_19736,N_19956);
nor UO_148 (O_148,N_19944,N_19656);
nor UO_149 (O_149,N_19891,N_19651);
xnor UO_150 (O_150,N_19769,N_19669);
and UO_151 (O_151,N_19871,N_19655);
or UO_152 (O_152,N_19881,N_19676);
nand UO_153 (O_153,N_19580,N_19987);
xor UO_154 (O_154,N_19693,N_19870);
and UO_155 (O_155,N_19745,N_19880);
nor UO_156 (O_156,N_19771,N_19770);
nor UO_157 (O_157,N_19865,N_19550);
and UO_158 (O_158,N_19968,N_19961);
or UO_159 (O_159,N_19577,N_19875);
xor UO_160 (O_160,N_19516,N_19723);
nor UO_161 (O_161,N_19989,N_19918);
xnor UO_162 (O_162,N_19814,N_19519);
or UO_163 (O_163,N_19950,N_19596);
or UO_164 (O_164,N_19976,N_19984);
nand UO_165 (O_165,N_19839,N_19990);
nand UO_166 (O_166,N_19559,N_19707);
nand UO_167 (O_167,N_19614,N_19878);
or UO_168 (O_168,N_19794,N_19597);
or UO_169 (O_169,N_19884,N_19599);
nor UO_170 (O_170,N_19784,N_19532);
nand UO_171 (O_171,N_19764,N_19692);
and UO_172 (O_172,N_19508,N_19652);
nor UO_173 (O_173,N_19712,N_19844);
or UO_174 (O_174,N_19624,N_19677);
xor UO_175 (O_175,N_19854,N_19983);
nor UO_176 (O_176,N_19641,N_19933);
nand UO_177 (O_177,N_19574,N_19967);
or UO_178 (O_178,N_19868,N_19799);
nor UO_179 (O_179,N_19788,N_19621);
nor UO_180 (O_180,N_19958,N_19622);
or UO_181 (O_181,N_19581,N_19660);
and UO_182 (O_182,N_19734,N_19626);
xor UO_183 (O_183,N_19517,N_19720);
xor UO_184 (O_184,N_19727,N_19530);
nor UO_185 (O_185,N_19706,N_19566);
nand UO_186 (O_186,N_19859,N_19667);
xor UO_187 (O_187,N_19957,N_19719);
nand UO_188 (O_188,N_19579,N_19953);
or UO_189 (O_189,N_19963,N_19571);
nand UO_190 (O_190,N_19864,N_19895);
or UO_191 (O_191,N_19973,N_19697);
or UO_192 (O_192,N_19628,N_19618);
and UO_193 (O_193,N_19808,N_19602);
xor UO_194 (O_194,N_19959,N_19903);
nand UO_195 (O_195,N_19737,N_19556);
nor UO_196 (O_196,N_19605,N_19690);
and UO_197 (O_197,N_19549,N_19969);
nor UO_198 (O_198,N_19832,N_19715);
xnor UO_199 (O_199,N_19598,N_19522);
nor UO_200 (O_200,N_19807,N_19867);
and UO_201 (O_201,N_19632,N_19876);
nor UO_202 (O_202,N_19747,N_19582);
or UO_203 (O_203,N_19924,N_19694);
xor UO_204 (O_204,N_19804,N_19897);
or UO_205 (O_205,N_19659,N_19774);
and UO_206 (O_206,N_19827,N_19954);
nor UO_207 (O_207,N_19815,N_19949);
or UO_208 (O_208,N_19940,N_19905);
xor UO_209 (O_209,N_19787,N_19501);
or UO_210 (O_210,N_19563,N_19645);
nor UO_211 (O_211,N_19840,N_19930);
and UO_212 (O_212,N_19890,N_19575);
nand UO_213 (O_213,N_19588,N_19981);
and UO_214 (O_214,N_19520,N_19546);
and UO_215 (O_215,N_19548,N_19557);
nand UO_216 (O_216,N_19838,N_19620);
and UO_217 (O_217,N_19606,N_19594);
xor UO_218 (O_218,N_19615,N_19937);
nor UO_219 (O_219,N_19858,N_19900);
nor UO_220 (O_220,N_19980,N_19611);
and UO_221 (O_221,N_19733,N_19928);
xnor UO_222 (O_222,N_19843,N_19806);
or UO_223 (O_223,N_19536,N_19999);
nor UO_224 (O_224,N_19841,N_19939);
xnor UO_225 (O_225,N_19988,N_19781);
and UO_226 (O_226,N_19750,N_19830);
and UO_227 (O_227,N_19817,N_19997);
xor UO_228 (O_228,N_19952,N_19672);
and UO_229 (O_229,N_19731,N_19916);
nand UO_230 (O_230,N_19850,N_19805);
nand UO_231 (O_231,N_19572,N_19744);
nand UO_232 (O_232,N_19663,N_19500);
nand UO_233 (O_233,N_19812,N_19523);
and UO_234 (O_234,N_19822,N_19955);
nand UO_235 (O_235,N_19934,N_19562);
or UO_236 (O_236,N_19862,N_19901);
nand UO_237 (O_237,N_19503,N_19925);
nand UO_238 (O_238,N_19778,N_19640);
or UO_239 (O_239,N_19560,N_19863);
nor UO_240 (O_240,N_19824,N_19635);
nand UO_241 (O_241,N_19551,N_19703);
nor UO_242 (O_242,N_19828,N_19836);
or UO_243 (O_243,N_19970,N_19528);
nor UO_244 (O_244,N_19570,N_19951);
and UO_245 (O_245,N_19591,N_19923);
xnor UO_246 (O_246,N_19849,N_19926);
nand UO_247 (O_247,N_19907,N_19513);
or UO_248 (O_248,N_19872,N_19979);
or UO_249 (O_249,N_19739,N_19935);
or UO_250 (O_250,N_19699,N_19892);
xnor UO_251 (O_251,N_19984,N_19519);
nand UO_252 (O_252,N_19504,N_19785);
nor UO_253 (O_253,N_19789,N_19983);
nand UO_254 (O_254,N_19713,N_19532);
nand UO_255 (O_255,N_19602,N_19803);
nor UO_256 (O_256,N_19981,N_19835);
nor UO_257 (O_257,N_19565,N_19578);
nand UO_258 (O_258,N_19714,N_19616);
or UO_259 (O_259,N_19919,N_19847);
nor UO_260 (O_260,N_19901,N_19768);
nand UO_261 (O_261,N_19603,N_19696);
nor UO_262 (O_262,N_19801,N_19578);
and UO_263 (O_263,N_19597,N_19702);
and UO_264 (O_264,N_19613,N_19918);
and UO_265 (O_265,N_19728,N_19732);
and UO_266 (O_266,N_19616,N_19816);
nor UO_267 (O_267,N_19931,N_19867);
and UO_268 (O_268,N_19732,N_19872);
or UO_269 (O_269,N_19738,N_19762);
nor UO_270 (O_270,N_19654,N_19912);
nor UO_271 (O_271,N_19984,N_19604);
and UO_272 (O_272,N_19823,N_19771);
nor UO_273 (O_273,N_19666,N_19798);
or UO_274 (O_274,N_19934,N_19586);
or UO_275 (O_275,N_19763,N_19580);
nand UO_276 (O_276,N_19864,N_19889);
and UO_277 (O_277,N_19938,N_19715);
and UO_278 (O_278,N_19555,N_19996);
xor UO_279 (O_279,N_19664,N_19651);
nor UO_280 (O_280,N_19995,N_19534);
nand UO_281 (O_281,N_19894,N_19938);
nor UO_282 (O_282,N_19895,N_19634);
xnor UO_283 (O_283,N_19917,N_19944);
nand UO_284 (O_284,N_19730,N_19914);
xnor UO_285 (O_285,N_19772,N_19623);
xnor UO_286 (O_286,N_19934,N_19568);
nor UO_287 (O_287,N_19653,N_19587);
nor UO_288 (O_288,N_19642,N_19915);
nor UO_289 (O_289,N_19728,N_19741);
nor UO_290 (O_290,N_19703,N_19826);
or UO_291 (O_291,N_19793,N_19978);
or UO_292 (O_292,N_19577,N_19581);
and UO_293 (O_293,N_19828,N_19919);
or UO_294 (O_294,N_19500,N_19513);
and UO_295 (O_295,N_19989,N_19733);
nor UO_296 (O_296,N_19996,N_19752);
and UO_297 (O_297,N_19569,N_19918);
nor UO_298 (O_298,N_19739,N_19921);
xor UO_299 (O_299,N_19714,N_19610);
or UO_300 (O_300,N_19911,N_19986);
nor UO_301 (O_301,N_19771,N_19656);
nor UO_302 (O_302,N_19507,N_19807);
nand UO_303 (O_303,N_19631,N_19629);
xor UO_304 (O_304,N_19618,N_19848);
or UO_305 (O_305,N_19721,N_19508);
nand UO_306 (O_306,N_19842,N_19580);
nor UO_307 (O_307,N_19732,N_19919);
xor UO_308 (O_308,N_19646,N_19828);
nor UO_309 (O_309,N_19996,N_19749);
xor UO_310 (O_310,N_19639,N_19767);
or UO_311 (O_311,N_19537,N_19666);
or UO_312 (O_312,N_19824,N_19534);
nand UO_313 (O_313,N_19737,N_19862);
nor UO_314 (O_314,N_19849,N_19844);
nand UO_315 (O_315,N_19695,N_19661);
and UO_316 (O_316,N_19618,N_19715);
and UO_317 (O_317,N_19839,N_19989);
nand UO_318 (O_318,N_19699,N_19868);
and UO_319 (O_319,N_19574,N_19995);
nand UO_320 (O_320,N_19812,N_19746);
and UO_321 (O_321,N_19988,N_19539);
or UO_322 (O_322,N_19975,N_19759);
nor UO_323 (O_323,N_19735,N_19771);
xnor UO_324 (O_324,N_19847,N_19584);
nand UO_325 (O_325,N_19527,N_19572);
nor UO_326 (O_326,N_19741,N_19559);
and UO_327 (O_327,N_19896,N_19662);
xnor UO_328 (O_328,N_19592,N_19893);
xor UO_329 (O_329,N_19689,N_19618);
or UO_330 (O_330,N_19567,N_19694);
nand UO_331 (O_331,N_19834,N_19929);
nor UO_332 (O_332,N_19558,N_19791);
nand UO_333 (O_333,N_19585,N_19888);
xor UO_334 (O_334,N_19570,N_19898);
nand UO_335 (O_335,N_19959,N_19511);
nand UO_336 (O_336,N_19863,N_19855);
or UO_337 (O_337,N_19610,N_19979);
nand UO_338 (O_338,N_19994,N_19749);
xnor UO_339 (O_339,N_19579,N_19857);
xor UO_340 (O_340,N_19660,N_19760);
and UO_341 (O_341,N_19938,N_19783);
or UO_342 (O_342,N_19993,N_19562);
or UO_343 (O_343,N_19581,N_19700);
nand UO_344 (O_344,N_19946,N_19895);
nor UO_345 (O_345,N_19818,N_19872);
and UO_346 (O_346,N_19636,N_19804);
or UO_347 (O_347,N_19681,N_19674);
nand UO_348 (O_348,N_19947,N_19518);
nor UO_349 (O_349,N_19891,N_19861);
nor UO_350 (O_350,N_19677,N_19809);
nand UO_351 (O_351,N_19931,N_19835);
nand UO_352 (O_352,N_19533,N_19817);
and UO_353 (O_353,N_19835,N_19728);
nand UO_354 (O_354,N_19787,N_19970);
nand UO_355 (O_355,N_19981,N_19870);
nor UO_356 (O_356,N_19888,N_19826);
or UO_357 (O_357,N_19564,N_19721);
or UO_358 (O_358,N_19986,N_19898);
xor UO_359 (O_359,N_19668,N_19847);
nor UO_360 (O_360,N_19960,N_19964);
xnor UO_361 (O_361,N_19826,N_19831);
nand UO_362 (O_362,N_19698,N_19500);
nand UO_363 (O_363,N_19547,N_19847);
nand UO_364 (O_364,N_19704,N_19904);
nand UO_365 (O_365,N_19701,N_19967);
xnor UO_366 (O_366,N_19753,N_19913);
nand UO_367 (O_367,N_19647,N_19828);
xor UO_368 (O_368,N_19582,N_19788);
nor UO_369 (O_369,N_19991,N_19619);
nor UO_370 (O_370,N_19515,N_19992);
nor UO_371 (O_371,N_19617,N_19691);
and UO_372 (O_372,N_19852,N_19872);
and UO_373 (O_373,N_19677,N_19996);
xor UO_374 (O_374,N_19874,N_19506);
xor UO_375 (O_375,N_19964,N_19720);
or UO_376 (O_376,N_19779,N_19773);
or UO_377 (O_377,N_19738,N_19630);
and UO_378 (O_378,N_19687,N_19609);
nand UO_379 (O_379,N_19688,N_19598);
or UO_380 (O_380,N_19753,N_19816);
and UO_381 (O_381,N_19623,N_19658);
nor UO_382 (O_382,N_19814,N_19929);
nand UO_383 (O_383,N_19764,N_19945);
nand UO_384 (O_384,N_19888,N_19874);
xnor UO_385 (O_385,N_19663,N_19638);
or UO_386 (O_386,N_19514,N_19524);
and UO_387 (O_387,N_19597,N_19575);
or UO_388 (O_388,N_19809,N_19585);
or UO_389 (O_389,N_19809,N_19871);
nand UO_390 (O_390,N_19806,N_19723);
xor UO_391 (O_391,N_19662,N_19646);
and UO_392 (O_392,N_19525,N_19666);
and UO_393 (O_393,N_19904,N_19931);
nand UO_394 (O_394,N_19956,N_19565);
nor UO_395 (O_395,N_19799,N_19748);
nand UO_396 (O_396,N_19558,N_19821);
nand UO_397 (O_397,N_19960,N_19517);
or UO_398 (O_398,N_19729,N_19569);
or UO_399 (O_399,N_19717,N_19524);
xnor UO_400 (O_400,N_19536,N_19627);
and UO_401 (O_401,N_19528,N_19986);
xnor UO_402 (O_402,N_19849,N_19684);
nand UO_403 (O_403,N_19770,N_19536);
and UO_404 (O_404,N_19704,N_19752);
or UO_405 (O_405,N_19850,N_19754);
nor UO_406 (O_406,N_19533,N_19509);
and UO_407 (O_407,N_19813,N_19946);
and UO_408 (O_408,N_19862,N_19836);
or UO_409 (O_409,N_19505,N_19972);
nor UO_410 (O_410,N_19514,N_19547);
nor UO_411 (O_411,N_19821,N_19795);
nand UO_412 (O_412,N_19556,N_19519);
nor UO_413 (O_413,N_19594,N_19651);
and UO_414 (O_414,N_19970,N_19544);
nand UO_415 (O_415,N_19621,N_19823);
nor UO_416 (O_416,N_19502,N_19614);
nand UO_417 (O_417,N_19913,N_19711);
or UO_418 (O_418,N_19712,N_19766);
xnor UO_419 (O_419,N_19505,N_19846);
nand UO_420 (O_420,N_19643,N_19737);
nand UO_421 (O_421,N_19913,N_19977);
nand UO_422 (O_422,N_19943,N_19636);
nand UO_423 (O_423,N_19614,N_19974);
nand UO_424 (O_424,N_19581,N_19930);
nand UO_425 (O_425,N_19721,N_19669);
xnor UO_426 (O_426,N_19962,N_19837);
nor UO_427 (O_427,N_19904,N_19861);
nor UO_428 (O_428,N_19994,N_19847);
nor UO_429 (O_429,N_19507,N_19582);
or UO_430 (O_430,N_19944,N_19546);
or UO_431 (O_431,N_19848,N_19811);
or UO_432 (O_432,N_19719,N_19527);
or UO_433 (O_433,N_19924,N_19827);
nand UO_434 (O_434,N_19576,N_19847);
or UO_435 (O_435,N_19516,N_19933);
or UO_436 (O_436,N_19909,N_19597);
xnor UO_437 (O_437,N_19830,N_19994);
and UO_438 (O_438,N_19890,N_19866);
xnor UO_439 (O_439,N_19584,N_19690);
nor UO_440 (O_440,N_19614,N_19632);
or UO_441 (O_441,N_19547,N_19518);
xnor UO_442 (O_442,N_19626,N_19658);
or UO_443 (O_443,N_19690,N_19692);
or UO_444 (O_444,N_19546,N_19943);
or UO_445 (O_445,N_19641,N_19575);
nor UO_446 (O_446,N_19783,N_19704);
nand UO_447 (O_447,N_19885,N_19503);
nor UO_448 (O_448,N_19869,N_19929);
nor UO_449 (O_449,N_19515,N_19963);
nand UO_450 (O_450,N_19718,N_19819);
or UO_451 (O_451,N_19865,N_19845);
xor UO_452 (O_452,N_19521,N_19610);
and UO_453 (O_453,N_19725,N_19852);
nor UO_454 (O_454,N_19840,N_19740);
and UO_455 (O_455,N_19741,N_19544);
nand UO_456 (O_456,N_19698,N_19941);
xor UO_457 (O_457,N_19892,N_19559);
nand UO_458 (O_458,N_19770,N_19501);
and UO_459 (O_459,N_19860,N_19731);
nand UO_460 (O_460,N_19587,N_19621);
and UO_461 (O_461,N_19539,N_19646);
xor UO_462 (O_462,N_19716,N_19810);
xor UO_463 (O_463,N_19567,N_19904);
xnor UO_464 (O_464,N_19509,N_19518);
nand UO_465 (O_465,N_19731,N_19838);
xor UO_466 (O_466,N_19757,N_19816);
or UO_467 (O_467,N_19870,N_19797);
or UO_468 (O_468,N_19939,N_19846);
and UO_469 (O_469,N_19717,N_19968);
nand UO_470 (O_470,N_19966,N_19982);
nor UO_471 (O_471,N_19995,N_19673);
nand UO_472 (O_472,N_19878,N_19612);
or UO_473 (O_473,N_19621,N_19982);
and UO_474 (O_474,N_19960,N_19938);
and UO_475 (O_475,N_19961,N_19773);
or UO_476 (O_476,N_19940,N_19771);
nand UO_477 (O_477,N_19965,N_19812);
nor UO_478 (O_478,N_19852,N_19922);
nor UO_479 (O_479,N_19754,N_19962);
or UO_480 (O_480,N_19780,N_19679);
nand UO_481 (O_481,N_19683,N_19976);
xnor UO_482 (O_482,N_19631,N_19744);
or UO_483 (O_483,N_19834,N_19843);
and UO_484 (O_484,N_19614,N_19597);
and UO_485 (O_485,N_19556,N_19744);
or UO_486 (O_486,N_19515,N_19730);
or UO_487 (O_487,N_19631,N_19675);
xor UO_488 (O_488,N_19688,N_19534);
and UO_489 (O_489,N_19902,N_19782);
and UO_490 (O_490,N_19995,N_19867);
nand UO_491 (O_491,N_19932,N_19532);
or UO_492 (O_492,N_19604,N_19851);
and UO_493 (O_493,N_19870,N_19796);
and UO_494 (O_494,N_19601,N_19747);
nand UO_495 (O_495,N_19654,N_19765);
and UO_496 (O_496,N_19966,N_19721);
or UO_497 (O_497,N_19714,N_19871);
xor UO_498 (O_498,N_19963,N_19501);
nor UO_499 (O_499,N_19654,N_19801);
nor UO_500 (O_500,N_19653,N_19761);
and UO_501 (O_501,N_19777,N_19798);
or UO_502 (O_502,N_19957,N_19744);
nor UO_503 (O_503,N_19835,N_19748);
and UO_504 (O_504,N_19684,N_19628);
xor UO_505 (O_505,N_19642,N_19786);
nor UO_506 (O_506,N_19544,N_19895);
nor UO_507 (O_507,N_19790,N_19805);
or UO_508 (O_508,N_19737,N_19718);
nand UO_509 (O_509,N_19738,N_19888);
nand UO_510 (O_510,N_19627,N_19663);
nor UO_511 (O_511,N_19620,N_19507);
and UO_512 (O_512,N_19812,N_19531);
nor UO_513 (O_513,N_19692,N_19602);
and UO_514 (O_514,N_19847,N_19910);
and UO_515 (O_515,N_19786,N_19834);
nand UO_516 (O_516,N_19840,N_19945);
or UO_517 (O_517,N_19932,N_19949);
nand UO_518 (O_518,N_19718,N_19872);
or UO_519 (O_519,N_19600,N_19853);
and UO_520 (O_520,N_19879,N_19775);
xor UO_521 (O_521,N_19983,N_19865);
nor UO_522 (O_522,N_19687,N_19989);
nor UO_523 (O_523,N_19934,N_19781);
nand UO_524 (O_524,N_19536,N_19987);
or UO_525 (O_525,N_19639,N_19587);
xor UO_526 (O_526,N_19763,N_19545);
xor UO_527 (O_527,N_19632,N_19579);
or UO_528 (O_528,N_19514,N_19747);
nand UO_529 (O_529,N_19985,N_19721);
xnor UO_530 (O_530,N_19778,N_19674);
or UO_531 (O_531,N_19631,N_19848);
nand UO_532 (O_532,N_19611,N_19810);
or UO_533 (O_533,N_19665,N_19941);
or UO_534 (O_534,N_19660,N_19623);
or UO_535 (O_535,N_19729,N_19682);
or UO_536 (O_536,N_19769,N_19700);
and UO_537 (O_537,N_19922,N_19663);
nand UO_538 (O_538,N_19853,N_19582);
nor UO_539 (O_539,N_19606,N_19577);
or UO_540 (O_540,N_19637,N_19777);
nand UO_541 (O_541,N_19845,N_19733);
and UO_542 (O_542,N_19648,N_19948);
nor UO_543 (O_543,N_19813,N_19955);
and UO_544 (O_544,N_19532,N_19610);
or UO_545 (O_545,N_19641,N_19517);
or UO_546 (O_546,N_19811,N_19517);
or UO_547 (O_547,N_19836,N_19980);
and UO_548 (O_548,N_19819,N_19795);
or UO_549 (O_549,N_19754,N_19712);
and UO_550 (O_550,N_19556,N_19843);
nand UO_551 (O_551,N_19955,N_19972);
xnor UO_552 (O_552,N_19567,N_19736);
and UO_553 (O_553,N_19939,N_19929);
and UO_554 (O_554,N_19730,N_19597);
and UO_555 (O_555,N_19657,N_19679);
xor UO_556 (O_556,N_19694,N_19932);
and UO_557 (O_557,N_19930,N_19529);
nor UO_558 (O_558,N_19962,N_19607);
nor UO_559 (O_559,N_19924,N_19503);
or UO_560 (O_560,N_19905,N_19911);
and UO_561 (O_561,N_19672,N_19721);
and UO_562 (O_562,N_19746,N_19859);
and UO_563 (O_563,N_19836,N_19544);
nand UO_564 (O_564,N_19683,N_19860);
xnor UO_565 (O_565,N_19658,N_19533);
nor UO_566 (O_566,N_19957,N_19971);
xor UO_567 (O_567,N_19519,N_19983);
nor UO_568 (O_568,N_19512,N_19595);
or UO_569 (O_569,N_19921,N_19608);
xor UO_570 (O_570,N_19977,N_19899);
and UO_571 (O_571,N_19954,N_19516);
or UO_572 (O_572,N_19607,N_19676);
xnor UO_573 (O_573,N_19555,N_19698);
and UO_574 (O_574,N_19665,N_19523);
nor UO_575 (O_575,N_19783,N_19654);
nand UO_576 (O_576,N_19582,N_19908);
or UO_577 (O_577,N_19551,N_19599);
or UO_578 (O_578,N_19676,N_19728);
xor UO_579 (O_579,N_19661,N_19856);
xnor UO_580 (O_580,N_19656,N_19935);
or UO_581 (O_581,N_19844,N_19565);
and UO_582 (O_582,N_19646,N_19930);
nor UO_583 (O_583,N_19571,N_19510);
and UO_584 (O_584,N_19560,N_19816);
and UO_585 (O_585,N_19526,N_19549);
nand UO_586 (O_586,N_19598,N_19601);
nand UO_587 (O_587,N_19608,N_19698);
and UO_588 (O_588,N_19675,N_19903);
or UO_589 (O_589,N_19807,N_19614);
and UO_590 (O_590,N_19540,N_19707);
nor UO_591 (O_591,N_19587,N_19675);
and UO_592 (O_592,N_19606,N_19517);
and UO_593 (O_593,N_19890,N_19776);
nor UO_594 (O_594,N_19897,N_19836);
nor UO_595 (O_595,N_19667,N_19623);
nand UO_596 (O_596,N_19945,N_19528);
nor UO_597 (O_597,N_19876,N_19991);
xor UO_598 (O_598,N_19551,N_19670);
nor UO_599 (O_599,N_19698,N_19645);
and UO_600 (O_600,N_19856,N_19781);
nand UO_601 (O_601,N_19571,N_19620);
nand UO_602 (O_602,N_19861,N_19873);
and UO_603 (O_603,N_19549,N_19599);
nor UO_604 (O_604,N_19866,N_19697);
nor UO_605 (O_605,N_19972,N_19867);
and UO_606 (O_606,N_19626,N_19868);
and UO_607 (O_607,N_19551,N_19622);
nand UO_608 (O_608,N_19731,N_19554);
or UO_609 (O_609,N_19889,N_19626);
nor UO_610 (O_610,N_19967,N_19999);
nor UO_611 (O_611,N_19563,N_19702);
nor UO_612 (O_612,N_19880,N_19710);
or UO_613 (O_613,N_19628,N_19626);
xnor UO_614 (O_614,N_19993,N_19645);
and UO_615 (O_615,N_19782,N_19514);
and UO_616 (O_616,N_19640,N_19571);
or UO_617 (O_617,N_19718,N_19890);
xnor UO_618 (O_618,N_19583,N_19997);
nand UO_619 (O_619,N_19972,N_19673);
and UO_620 (O_620,N_19990,N_19622);
xnor UO_621 (O_621,N_19515,N_19763);
nor UO_622 (O_622,N_19934,N_19577);
nor UO_623 (O_623,N_19631,N_19804);
and UO_624 (O_624,N_19893,N_19678);
and UO_625 (O_625,N_19563,N_19958);
xor UO_626 (O_626,N_19524,N_19608);
xnor UO_627 (O_627,N_19597,N_19916);
and UO_628 (O_628,N_19886,N_19889);
xnor UO_629 (O_629,N_19549,N_19527);
nand UO_630 (O_630,N_19634,N_19715);
nor UO_631 (O_631,N_19935,N_19887);
and UO_632 (O_632,N_19661,N_19735);
and UO_633 (O_633,N_19516,N_19670);
or UO_634 (O_634,N_19588,N_19544);
xor UO_635 (O_635,N_19736,N_19891);
or UO_636 (O_636,N_19734,N_19691);
xnor UO_637 (O_637,N_19588,N_19598);
nor UO_638 (O_638,N_19799,N_19895);
nand UO_639 (O_639,N_19710,N_19651);
nand UO_640 (O_640,N_19670,N_19837);
and UO_641 (O_641,N_19585,N_19844);
or UO_642 (O_642,N_19605,N_19648);
xnor UO_643 (O_643,N_19938,N_19974);
nor UO_644 (O_644,N_19553,N_19657);
nand UO_645 (O_645,N_19756,N_19646);
nand UO_646 (O_646,N_19915,N_19673);
nand UO_647 (O_647,N_19719,N_19720);
xor UO_648 (O_648,N_19822,N_19960);
xor UO_649 (O_649,N_19689,N_19558);
and UO_650 (O_650,N_19932,N_19829);
nand UO_651 (O_651,N_19558,N_19671);
nand UO_652 (O_652,N_19641,N_19585);
xnor UO_653 (O_653,N_19988,N_19903);
nor UO_654 (O_654,N_19571,N_19554);
nor UO_655 (O_655,N_19851,N_19815);
xnor UO_656 (O_656,N_19927,N_19705);
xor UO_657 (O_657,N_19916,N_19937);
nor UO_658 (O_658,N_19536,N_19528);
and UO_659 (O_659,N_19974,N_19705);
nand UO_660 (O_660,N_19899,N_19646);
nand UO_661 (O_661,N_19908,N_19961);
nor UO_662 (O_662,N_19890,N_19536);
and UO_663 (O_663,N_19788,N_19655);
nand UO_664 (O_664,N_19896,N_19877);
or UO_665 (O_665,N_19772,N_19975);
nor UO_666 (O_666,N_19776,N_19864);
xnor UO_667 (O_667,N_19927,N_19545);
nand UO_668 (O_668,N_19562,N_19695);
nor UO_669 (O_669,N_19904,N_19949);
and UO_670 (O_670,N_19945,N_19993);
or UO_671 (O_671,N_19700,N_19956);
or UO_672 (O_672,N_19639,N_19678);
or UO_673 (O_673,N_19804,N_19986);
or UO_674 (O_674,N_19668,N_19768);
xor UO_675 (O_675,N_19618,N_19993);
nand UO_676 (O_676,N_19757,N_19526);
xnor UO_677 (O_677,N_19595,N_19928);
nor UO_678 (O_678,N_19722,N_19823);
and UO_679 (O_679,N_19850,N_19815);
nand UO_680 (O_680,N_19893,N_19700);
nor UO_681 (O_681,N_19933,N_19726);
nand UO_682 (O_682,N_19501,N_19510);
nor UO_683 (O_683,N_19901,N_19833);
xor UO_684 (O_684,N_19507,N_19551);
xnor UO_685 (O_685,N_19526,N_19697);
nand UO_686 (O_686,N_19562,N_19870);
nand UO_687 (O_687,N_19840,N_19601);
nand UO_688 (O_688,N_19706,N_19803);
and UO_689 (O_689,N_19865,N_19830);
nand UO_690 (O_690,N_19952,N_19555);
nor UO_691 (O_691,N_19888,N_19702);
or UO_692 (O_692,N_19720,N_19721);
xor UO_693 (O_693,N_19639,N_19765);
nor UO_694 (O_694,N_19658,N_19570);
or UO_695 (O_695,N_19609,N_19898);
and UO_696 (O_696,N_19605,N_19630);
xnor UO_697 (O_697,N_19608,N_19688);
nand UO_698 (O_698,N_19566,N_19923);
nor UO_699 (O_699,N_19766,N_19814);
and UO_700 (O_700,N_19623,N_19944);
nand UO_701 (O_701,N_19925,N_19783);
and UO_702 (O_702,N_19902,N_19577);
and UO_703 (O_703,N_19912,N_19738);
nor UO_704 (O_704,N_19779,N_19711);
xor UO_705 (O_705,N_19531,N_19839);
and UO_706 (O_706,N_19541,N_19820);
nand UO_707 (O_707,N_19810,N_19733);
nor UO_708 (O_708,N_19656,N_19713);
or UO_709 (O_709,N_19616,N_19618);
nand UO_710 (O_710,N_19530,N_19575);
xor UO_711 (O_711,N_19702,N_19893);
nand UO_712 (O_712,N_19934,N_19806);
or UO_713 (O_713,N_19786,N_19640);
and UO_714 (O_714,N_19993,N_19737);
xnor UO_715 (O_715,N_19704,N_19779);
or UO_716 (O_716,N_19919,N_19771);
xnor UO_717 (O_717,N_19868,N_19720);
and UO_718 (O_718,N_19711,N_19998);
xor UO_719 (O_719,N_19534,N_19617);
and UO_720 (O_720,N_19869,N_19534);
xnor UO_721 (O_721,N_19614,N_19500);
nand UO_722 (O_722,N_19789,N_19908);
xor UO_723 (O_723,N_19671,N_19959);
or UO_724 (O_724,N_19624,N_19559);
nor UO_725 (O_725,N_19744,N_19521);
and UO_726 (O_726,N_19593,N_19611);
nand UO_727 (O_727,N_19905,N_19725);
or UO_728 (O_728,N_19599,N_19518);
nand UO_729 (O_729,N_19869,N_19577);
nor UO_730 (O_730,N_19825,N_19683);
or UO_731 (O_731,N_19656,N_19600);
or UO_732 (O_732,N_19898,N_19510);
and UO_733 (O_733,N_19975,N_19764);
nor UO_734 (O_734,N_19866,N_19682);
nand UO_735 (O_735,N_19610,N_19924);
xor UO_736 (O_736,N_19721,N_19950);
nor UO_737 (O_737,N_19869,N_19595);
nor UO_738 (O_738,N_19841,N_19839);
xnor UO_739 (O_739,N_19660,N_19847);
or UO_740 (O_740,N_19850,N_19607);
nand UO_741 (O_741,N_19512,N_19815);
nand UO_742 (O_742,N_19796,N_19768);
xnor UO_743 (O_743,N_19739,N_19832);
or UO_744 (O_744,N_19501,N_19994);
nor UO_745 (O_745,N_19860,N_19530);
or UO_746 (O_746,N_19947,N_19513);
xor UO_747 (O_747,N_19618,N_19549);
or UO_748 (O_748,N_19557,N_19804);
nor UO_749 (O_749,N_19642,N_19820);
nand UO_750 (O_750,N_19763,N_19511);
nor UO_751 (O_751,N_19937,N_19605);
or UO_752 (O_752,N_19819,N_19618);
nand UO_753 (O_753,N_19584,N_19552);
nand UO_754 (O_754,N_19946,N_19518);
nand UO_755 (O_755,N_19702,N_19914);
nand UO_756 (O_756,N_19539,N_19854);
xnor UO_757 (O_757,N_19613,N_19507);
nand UO_758 (O_758,N_19971,N_19791);
nand UO_759 (O_759,N_19510,N_19551);
nand UO_760 (O_760,N_19865,N_19610);
nand UO_761 (O_761,N_19695,N_19776);
xor UO_762 (O_762,N_19844,N_19508);
nand UO_763 (O_763,N_19670,N_19972);
nor UO_764 (O_764,N_19918,N_19619);
nor UO_765 (O_765,N_19871,N_19776);
xor UO_766 (O_766,N_19836,N_19918);
nand UO_767 (O_767,N_19826,N_19660);
xor UO_768 (O_768,N_19616,N_19867);
and UO_769 (O_769,N_19594,N_19592);
nand UO_770 (O_770,N_19859,N_19931);
nand UO_771 (O_771,N_19964,N_19536);
and UO_772 (O_772,N_19936,N_19514);
or UO_773 (O_773,N_19560,N_19940);
nand UO_774 (O_774,N_19648,N_19853);
nand UO_775 (O_775,N_19550,N_19696);
nand UO_776 (O_776,N_19753,N_19708);
nand UO_777 (O_777,N_19974,N_19600);
nor UO_778 (O_778,N_19745,N_19947);
nand UO_779 (O_779,N_19534,N_19645);
or UO_780 (O_780,N_19808,N_19769);
xnor UO_781 (O_781,N_19638,N_19954);
nor UO_782 (O_782,N_19861,N_19960);
and UO_783 (O_783,N_19787,N_19500);
or UO_784 (O_784,N_19634,N_19628);
nand UO_785 (O_785,N_19786,N_19648);
and UO_786 (O_786,N_19579,N_19511);
or UO_787 (O_787,N_19559,N_19639);
and UO_788 (O_788,N_19628,N_19880);
or UO_789 (O_789,N_19937,N_19816);
nor UO_790 (O_790,N_19786,N_19584);
xnor UO_791 (O_791,N_19562,N_19675);
and UO_792 (O_792,N_19798,N_19936);
nand UO_793 (O_793,N_19779,N_19874);
xnor UO_794 (O_794,N_19841,N_19685);
nand UO_795 (O_795,N_19881,N_19925);
nor UO_796 (O_796,N_19889,N_19675);
and UO_797 (O_797,N_19512,N_19673);
or UO_798 (O_798,N_19646,N_19906);
nand UO_799 (O_799,N_19689,N_19810);
xor UO_800 (O_800,N_19988,N_19880);
nor UO_801 (O_801,N_19797,N_19659);
xor UO_802 (O_802,N_19672,N_19873);
nand UO_803 (O_803,N_19538,N_19598);
or UO_804 (O_804,N_19735,N_19985);
nor UO_805 (O_805,N_19990,N_19835);
nor UO_806 (O_806,N_19514,N_19954);
nand UO_807 (O_807,N_19888,N_19690);
or UO_808 (O_808,N_19683,N_19690);
nor UO_809 (O_809,N_19555,N_19623);
nor UO_810 (O_810,N_19701,N_19614);
xor UO_811 (O_811,N_19777,N_19860);
nor UO_812 (O_812,N_19879,N_19917);
nand UO_813 (O_813,N_19575,N_19538);
or UO_814 (O_814,N_19782,N_19725);
nor UO_815 (O_815,N_19882,N_19823);
and UO_816 (O_816,N_19760,N_19821);
xor UO_817 (O_817,N_19716,N_19864);
or UO_818 (O_818,N_19797,N_19920);
nor UO_819 (O_819,N_19867,N_19922);
nand UO_820 (O_820,N_19869,N_19847);
xnor UO_821 (O_821,N_19513,N_19943);
xor UO_822 (O_822,N_19619,N_19982);
or UO_823 (O_823,N_19792,N_19606);
or UO_824 (O_824,N_19753,N_19875);
xnor UO_825 (O_825,N_19767,N_19713);
or UO_826 (O_826,N_19800,N_19932);
or UO_827 (O_827,N_19886,N_19828);
nor UO_828 (O_828,N_19595,N_19915);
or UO_829 (O_829,N_19922,N_19989);
nand UO_830 (O_830,N_19865,N_19627);
and UO_831 (O_831,N_19653,N_19915);
nor UO_832 (O_832,N_19732,N_19700);
nand UO_833 (O_833,N_19799,N_19554);
and UO_834 (O_834,N_19713,N_19920);
nand UO_835 (O_835,N_19679,N_19555);
or UO_836 (O_836,N_19914,N_19983);
and UO_837 (O_837,N_19981,N_19974);
nor UO_838 (O_838,N_19847,N_19593);
or UO_839 (O_839,N_19574,N_19798);
nor UO_840 (O_840,N_19595,N_19790);
or UO_841 (O_841,N_19835,N_19549);
xor UO_842 (O_842,N_19973,N_19731);
xor UO_843 (O_843,N_19708,N_19793);
xor UO_844 (O_844,N_19637,N_19956);
and UO_845 (O_845,N_19828,N_19521);
nand UO_846 (O_846,N_19802,N_19674);
xnor UO_847 (O_847,N_19529,N_19941);
or UO_848 (O_848,N_19635,N_19512);
xnor UO_849 (O_849,N_19565,N_19725);
or UO_850 (O_850,N_19815,N_19714);
and UO_851 (O_851,N_19740,N_19593);
nand UO_852 (O_852,N_19888,N_19529);
nor UO_853 (O_853,N_19665,N_19909);
xnor UO_854 (O_854,N_19638,N_19791);
and UO_855 (O_855,N_19940,N_19801);
xnor UO_856 (O_856,N_19768,N_19912);
nand UO_857 (O_857,N_19763,N_19689);
nor UO_858 (O_858,N_19608,N_19781);
and UO_859 (O_859,N_19739,N_19594);
or UO_860 (O_860,N_19736,N_19515);
xnor UO_861 (O_861,N_19787,N_19867);
nand UO_862 (O_862,N_19940,N_19782);
or UO_863 (O_863,N_19998,N_19717);
or UO_864 (O_864,N_19777,N_19985);
and UO_865 (O_865,N_19731,N_19503);
nor UO_866 (O_866,N_19929,N_19692);
nor UO_867 (O_867,N_19573,N_19670);
nor UO_868 (O_868,N_19726,N_19701);
and UO_869 (O_869,N_19725,N_19545);
nand UO_870 (O_870,N_19912,N_19904);
and UO_871 (O_871,N_19851,N_19914);
nor UO_872 (O_872,N_19881,N_19621);
and UO_873 (O_873,N_19744,N_19597);
xor UO_874 (O_874,N_19883,N_19793);
nand UO_875 (O_875,N_19831,N_19919);
or UO_876 (O_876,N_19729,N_19642);
nor UO_877 (O_877,N_19856,N_19634);
or UO_878 (O_878,N_19533,N_19966);
or UO_879 (O_879,N_19808,N_19864);
nor UO_880 (O_880,N_19920,N_19661);
or UO_881 (O_881,N_19590,N_19730);
nand UO_882 (O_882,N_19761,N_19821);
xor UO_883 (O_883,N_19709,N_19961);
nor UO_884 (O_884,N_19782,N_19913);
or UO_885 (O_885,N_19988,N_19968);
or UO_886 (O_886,N_19771,N_19818);
nor UO_887 (O_887,N_19541,N_19512);
or UO_888 (O_888,N_19505,N_19895);
xor UO_889 (O_889,N_19614,N_19634);
nand UO_890 (O_890,N_19567,N_19792);
or UO_891 (O_891,N_19608,N_19592);
and UO_892 (O_892,N_19628,N_19822);
xor UO_893 (O_893,N_19660,N_19824);
nor UO_894 (O_894,N_19579,N_19990);
nor UO_895 (O_895,N_19912,N_19696);
nand UO_896 (O_896,N_19646,N_19861);
or UO_897 (O_897,N_19534,N_19993);
or UO_898 (O_898,N_19630,N_19758);
nor UO_899 (O_899,N_19532,N_19577);
or UO_900 (O_900,N_19614,N_19520);
xor UO_901 (O_901,N_19983,N_19583);
nand UO_902 (O_902,N_19923,N_19530);
xnor UO_903 (O_903,N_19885,N_19711);
or UO_904 (O_904,N_19706,N_19699);
nor UO_905 (O_905,N_19881,N_19552);
or UO_906 (O_906,N_19719,N_19874);
xor UO_907 (O_907,N_19694,N_19838);
nor UO_908 (O_908,N_19563,N_19865);
nand UO_909 (O_909,N_19781,N_19657);
nor UO_910 (O_910,N_19740,N_19882);
nor UO_911 (O_911,N_19933,N_19785);
and UO_912 (O_912,N_19630,N_19962);
xor UO_913 (O_913,N_19604,N_19699);
and UO_914 (O_914,N_19544,N_19669);
xnor UO_915 (O_915,N_19952,N_19714);
xnor UO_916 (O_916,N_19709,N_19934);
or UO_917 (O_917,N_19992,N_19844);
or UO_918 (O_918,N_19622,N_19560);
nor UO_919 (O_919,N_19673,N_19822);
nand UO_920 (O_920,N_19817,N_19846);
xnor UO_921 (O_921,N_19745,N_19861);
nand UO_922 (O_922,N_19961,N_19651);
and UO_923 (O_923,N_19721,N_19605);
nor UO_924 (O_924,N_19797,N_19550);
nor UO_925 (O_925,N_19515,N_19533);
and UO_926 (O_926,N_19901,N_19510);
and UO_927 (O_927,N_19934,N_19865);
or UO_928 (O_928,N_19654,N_19519);
xor UO_929 (O_929,N_19634,N_19923);
xor UO_930 (O_930,N_19582,N_19800);
nand UO_931 (O_931,N_19591,N_19928);
or UO_932 (O_932,N_19618,N_19638);
xor UO_933 (O_933,N_19914,N_19803);
or UO_934 (O_934,N_19591,N_19842);
and UO_935 (O_935,N_19502,N_19896);
or UO_936 (O_936,N_19978,N_19838);
or UO_937 (O_937,N_19837,N_19703);
nor UO_938 (O_938,N_19505,N_19600);
nor UO_939 (O_939,N_19973,N_19523);
nor UO_940 (O_940,N_19855,N_19718);
nor UO_941 (O_941,N_19776,N_19812);
or UO_942 (O_942,N_19970,N_19531);
nand UO_943 (O_943,N_19672,N_19982);
or UO_944 (O_944,N_19510,N_19872);
or UO_945 (O_945,N_19693,N_19561);
xnor UO_946 (O_946,N_19887,N_19664);
and UO_947 (O_947,N_19924,N_19616);
nand UO_948 (O_948,N_19826,N_19678);
and UO_949 (O_949,N_19818,N_19662);
nor UO_950 (O_950,N_19929,N_19563);
nor UO_951 (O_951,N_19862,N_19529);
nand UO_952 (O_952,N_19760,N_19904);
nand UO_953 (O_953,N_19643,N_19832);
or UO_954 (O_954,N_19840,N_19926);
xor UO_955 (O_955,N_19920,N_19523);
nor UO_956 (O_956,N_19735,N_19819);
nor UO_957 (O_957,N_19926,N_19608);
and UO_958 (O_958,N_19579,N_19680);
nor UO_959 (O_959,N_19698,N_19968);
nor UO_960 (O_960,N_19685,N_19767);
nand UO_961 (O_961,N_19923,N_19859);
nor UO_962 (O_962,N_19753,N_19634);
nand UO_963 (O_963,N_19912,N_19619);
or UO_964 (O_964,N_19994,N_19645);
nand UO_965 (O_965,N_19718,N_19514);
xor UO_966 (O_966,N_19676,N_19953);
nand UO_967 (O_967,N_19518,N_19638);
and UO_968 (O_968,N_19898,N_19665);
or UO_969 (O_969,N_19812,N_19706);
xnor UO_970 (O_970,N_19887,N_19875);
and UO_971 (O_971,N_19667,N_19675);
and UO_972 (O_972,N_19889,N_19727);
xor UO_973 (O_973,N_19612,N_19799);
xor UO_974 (O_974,N_19555,N_19752);
nand UO_975 (O_975,N_19896,N_19744);
or UO_976 (O_976,N_19786,N_19777);
nor UO_977 (O_977,N_19993,N_19905);
nand UO_978 (O_978,N_19878,N_19556);
or UO_979 (O_979,N_19967,N_19741);
or UO_980 (O_980,N_19655,N_19947);
nor UO_981 (O_981,N_19520,N_19908);
or UO_982 (O_982,N_19606,N_19873);
nand UO_983 (O_983,N_19740,N_19735);
nor UO_984 (O_984,N_19732,N_19512);
xor UO_985 (O_985,N_19630,N_19777);
or UO_986 (O_986,N_19691,N_19812);
nor UO_987 (O_987,N_19620,N_19895);
and UO_988 (O_988,N_19902,N_19693);
nand UO_989 (O_989,N_19769,N_19874);
nand UO_990 (O_990,N_19628,N_19532);
xor UO_991 (O_991,N_19803,N_19737);
or UO_992 (O_992,N_19823,N_19500);
or UO_993 (O_993,N_19932,N_19647);
or UO_994 (O_994,N_19628,N_19937);
xnor UO_995 (O_995,N_19742,N_19583);
xor UO_996 (O_996,N_19857,N_19945);
or UO_997 (O_997,N_19582,N_19531);
nor UO_998 (O_998,N_19806,N_19506);
or UO_999 (O_999,N_19661,N_19868);
nor UO_1000 (O_1000,N_19569,N_19987);
nand UO_1001 (O_1001,N_19821,N_19612);
nor UO_1002 (O_1002,N_19796,N_19604);
and UO_1003 (O_1003,N_19634,N_19886);
nor UO_1004 (O_1004,N_19967,N_19683);
and UO_1005 (O_1005,N_19864,N_19988);
or UO_1006 (O_1006,N_19503,N_19623);
nand UO_1007 (O_1007,N_19956,N_19595);
or UO_1008 (O_1008,N_19877,N_19562);
xnor UO_1009 (O_1009,N_19570,N_19930);
or UO_1010 (O_1010,N_19942,N_19962);
nand UO_1011 (O_1011,N_19567,N_19844);
or UO_1012 (O_1012,N_19741,N_19864);
nor UO_1013 (O_1013,N_19917,N_19548);
xor UO_1014 (O_1014,N_19902,N_19692);
and UO_1015 (O_1015,N_19974,N_19717);
or UO_1016 (O_1016,N_19876,N_19687);
and UO_1017 (O_1017,N_19843,N_19948);
and UO_1018 (O_1018,N_19684,N_19972);
and UO_1019 (O_1019,N_19587,N_19889);
xor UO_1020 (O_1020,N_19711,N_19607);
or UO_1021 (O_1021,N_19620,N_19927);
nor UO_1022 (O_1022,N_19517,N_19824);
nand UO_1023 (O_1023,N_19736,N_19987);
and UO_1024 (O_1024,N_19740,N_19649);
nor UO_1025 (O_1025,N_19685,N_19740);
and UO_1026 (O_1026,N_19774,N_19952);
nand UO_1027 (O_1027,N_19682,N_19519);
nand UO_1028 (O_1028,N_19810,N_19838);
and UO_1029 (O_1029,N_19991,N_19631);
xnor UO_1030 (O_1030,N_19978,N_19895);
and UO_1031 (O_1031,N_19897,N_19945);
or UO_1032 (O_1032,N_19770,N_19533);
nor UO_1033 (O_1033,N_19790,N_19591);
nor UO_1034 (O_1034,N_19921,N_19896);
or UO_1035 (O_1035,N_19904,N_19650);
nor UO_1036 (O_1036,N_19528,N_19527);
or UO_1037 (O_1037,N_19711,N_19619);
nor UO_1038 (O_1038,N_19797,N_19855);
or UO_1039 (O_1039,N_19992,N_19692);
or UO_1040 (O_1040,N_19500,N_19777);
xnor UO_1041 (O_1041,N_19604,N_19641);
xor UO_1042 (O_1042,N_19672,N_19647);
nand UO_1043 (O_1043,N_19602,N_19758);
or UO_1044 (O_1044,N_19646,N_19745);
xor UO_1045 (O_1045,N_19676,N_19965);
and UO_1046 (O_1046,N_19967,N_19692);
and UO_1047 (O_1047,N_19658,N_19686);
xor UO_1048 (O_1048,N_19510,N_19577);
xnor UO_1049 (O_1049,N_19888,N_19630);
nor UO_1050 (O_1050,N_19627,N_19934);
or UO_1051 (O_1051,N_19730,N_19622);
nor UO_1052 (O_1052,N_19957,N_19923);
nand UO_1053 (O_1053,N_19680,N_19733);
xor UO_1054 (O_1054,N_19930,N_19514);
and UO_1055 (O_1055,N_19545,N_19527);
and UO_1056 (O_1056,N_19676,N_19658);
nand UO_1057 (O_1057,N_19718,N_19984);
and UO_1058 (O_1058,N_19697,N_19751);
xnor UO_1059 (O_1059,N_19506,N_19890);
nand UO_1060 (O_1060,N_19888,N_19654);
or UO_1061 (O_1061,N_19644,N_19664);
nor UO_1062 (O_1062,N_19642,N_19860);
nand UO_1063 (O_1063,N_19635,N_19704);
nand UO_1064 (O_1064,N_19800,N_19694);
nor UO_1065 (O_1065,N_19741,N_19848);
xnor UO_1066 (O_1066,N_19813,N_19907);
or UO_1067 (O_1067,N_19767,N_19893);
and UO_1068 (O_1068,N_19936,N_19816);
or UO_1069 (O_1069,N_19577,N_19785);
nor UO_1070 (O_1070,N_19705,N_19907);
xor UO_1071 (O_1071,N_19949,N_19606);
xor UO_1072 (O_1072,N_19983,N_19912);
or UO_1073 (O_1073,N_19610,N_19508);
nor UO_1074 (O_1074,N_19644,N_19540);
nand UO_1075 (O_1075,N_19929,N_19642);
xor UO_1076 (O_1076,N_19774,N_19836);
and UO_1077 (O_1077,N_19723,N_19820);
and UO_1078 (O_1078,N_19945,N_19540);
xor UO_1079 (O_1079,N_19588,N_19821);
or UO_1080 (O_1080,N_19842,N_19672);
and UO_1081 (O_1081,N_19855,N_19525);
or UO_1082 (O_1082,N_19634,N_19850);
and UO_1083 (O_1083,N_19617,N_19781);
and UO_1084 (O_1084,N_19587,N_19502);
nor UO_1085 (O_1085,N_19708,N_19779);
nor UO_1086 (O_1086,N_19916,N_19650);
or UO_1087 (O_1087,N_19971,N_19714);
or UO_1088 (O_1088,N_19777,N_19709);
xnor UO_1089 (O_1089,N_19659,N_19879);
and UO_1090 (O_1090,N_19784,N_19647);
and UO_1091 (O_1091,N_19733,N_19866);
or UO_1092 (O_1092,N_19761,N_19760);
nor UO_1093 (O_1093,N_19626,N_19847);
and UO_1094 (O_1094,N_19913,N_19760);
and UO_1095 (O_1095,N_19558,N_19990);
or UO_1096 (O_1096,N_19671,N_19932);
xnor UO_1097 (O_1097,N_19969,N_19886);
xor UO_1098 (O_1098,N_19987,N_19582);
or UO_1099 (O_1099,N_19878,N_19548);
or UO_1100 (O_1100,N_19987,N_19776);
and UO_1101 (O_1101,N_19710,N_19895);
or UO_1102 (O_1102,N_19619,N_19564);
nand UO_1103 (O_1103,N_19564,N_19841);
or UO_1104 (O_1104,N_19521,N_19671);
or UO_1105 (O_1105,N_19904,N_19623);
xor UO_1106 (O_1106,N_19625,N_19534);
xnor UO_1107 (O_1107,N_19516,N_19937);
nand UO_1108 (O_1108,N_19651,N_19556);
or UO_1109 (O_1109,N_19749,N_19783);
xnor UO_1110 (O_1110,N_19842,N_19905);
nor UO_1111 (O_1111,N_19942,N_19622);
or UO_1112 (O_1112,N_19651,N_19902);
and UO_1113 (O_1113,N_19930,N_19857);
or UO_1114 (O_1114,N_19798,N_19985);
xor UO_1115 (O_1115,N_19591,N_19852);
and UO_1116 (O_1116,N_19820,N_19647);
nand UO_1117 (O_1117,N_19614,N_19892);
and UO_1118 (O_1118,N_19816,N_19614);
or UO_1119 (O_1119,N_19823,N_19736);
nand UO_1120 (O_1120,N_19620,N_19724);
or UO_1121 (O_1121,N_19709,N_19878);
and UO_1122 (O_1122,N_19882,N_19559);
nor UO_1123 (O_1123,N_19778,N_19801);
xnor UO_1124 (O_1124,N_19506,N_19850);
or UO_1125 (O_1125,N_19845,N_19722);
xnor UO_1126 (O_1126,N_19660,N_19976);
or UO_1127 (O_1127,N_19611,N_19648);
and UO_1128 (O_1128,N_19715,N_19721);
nor UO_1129 (O_1129,N_19540,N_19560);
or UO_1130 (O_1130,N_19779,N_19784);
nor UO_1131 (O_1131,N_19656,N_19777);
xnor UO_1132 (O_1132,N_19605,N_19934);
nand UO_1133 (O_1133,N_19953,N_19696);
xnor UO_1134 (O_1134,N_19641,N_19727);
nor UO_1135 (O_1135,N_19837,N_19528);
nor UO_1136 (O_1136,N_19523,N_19606);
and UO_1137 (O_1137,N_19535,N_19643);
nand UO_1138 (O_1138,N_19702,N_19841);
and UO_1139 (O_1139,N_19676,N_19747);
nand UO_1140 (O_1140,N_19783,N_19545);
xor UO_1141 (O_1141,N_19621,N_19975);
nand UO_1142 (O_1142,N_19649,N_19687);
and UO_1143 (O_1143,N_19804,N_19942);
nor UO_1144 (O_1144,N_19917,N_19500);
and UO_1145 (O_1145,N_19686,N_19676);
or UO_1146 (O_1146,N_19916,N_19725);
nor UO_1147 (O_1147,N_19786,N_19759);
and UO_1148 (O_1148,N_19780,N_19689);
and UO_1149 (O_1149,N_19804,N_19690);
nand UO_1150 (O_1150,N_19597,N_19974);
nand UO_1151 (O_1151,N_19507,N_19751);
or UO_1152 (O_1152,N_19506,N_19678);
nand UO_1153 (O_1153,N_19906,N_19891);
or UO_1154 (O_1154,N_19576,N_19897);
and UO_1155 (O_1155,N_19708,N_19758);
or UO_1156 (O_1156,N_19561,N_19699);
xnor UO_1157 (O_1157,N_19791,N_19685);
xnor UO_1158 (O_1158,N_19674,N_19689);
nor UO_1159 (O_1159,N_19529,N_19754);
or UO_1160 (O_1160,N_19812,N_19974);
or UO_1161 (O_1161,N_19744,N_19645);
xnor UO_1162 (O_1162,N_19696,N_19909);
xnor UO_1163 (O_1163,N_19781,N_19672);
nor UO_1164 (O_1164,N_19903,N_19545);
nor UO_1165 (O_1165,N_19599,N_19842);
nor UO_1166 (O_1166,N_19851,N_19671);
xor UO_1167 (O_1167,N_19955,N_19716);
xnor UO_1168 (O_1168,N_19676,N_19570);
xnor UO_1169 (O_1169,N_19551,N_19927);
nor UO_1170 (O_1170,N_19890,N_19994);
xnor UO_1171 (O_1171,N_19953,N_19834);
xnor UO_1172 (O_1172,N_19997,N_19753);
and UO_1173 (O_1173,N_19619,N_19806);
nand UO_1174 (O_1174,N_19883,N_19884);
xnor UO_1175 (O_1175,N_19709,N_19622);
nand UO_1176 (O_1176,N_19798,N_19566);
nand UO_1177 (O_1177,N_19504,N_19849);
nor UO_1178 (O_1178,N_19602,N_19825);
and UO_1179 (O_1179,N_19707,N_19870);
xnor UO_1180 (O_1180,N_19877,N_19786);
and UO_1181 (O_1181,N_19729,N_19508);
and UO_1182 (O_1182,N_19755,N_19766);
nand UO_1183 (O_1183,N_19846,N_19979);
nor UO_1184 (O_1184,N_19745,N_19652);
or UO_1185 (O_1185,N_19769,N_19511);
nor UO_1186 (O_1186,N_19734,N_19743);
or UO_1187 (O_1187,N_19872,N_19553);
nor UO_1188 (O_1188,N_19840,N_19563);
or UO_1189 (O_1189,N_19774,N_19922);
xnor UO_1190 (O_1190,N_19928,N_19801);
and UO_1191 (O_1191,N_19584,N_19583);
xnor UO_1192 (O_1192,N_19537,N_19572);
or UO_1193 (O_1193,N_19844,N_19518);
and UO_1194 (O_1194,N_19848,N_19908);
or UO_1195 (O_1195,N_19888,N_19775);
and UO_1196 (O_1196,N_19960,N_19981);
nand UO_1197 (O_1197,N_19619,N_19728);
and UO_1198 (O_1198,N_19740,N_19804);
or UO_1199 (O_1199,N_19504,N_19988);
and UO_1200 (O_1200,N_19904,N_19682);
or UO_1201 (O_1201,N_19659,N_19857);
and UO_1202 (O_1202,N_19925,N_19727);
nor UO_1203 (O_1203,N_19816,N_19872);
nand UO_1204 (O_1204,N_19857,N_19600);
nor UO_1205 (O_1205,N_19955,N_19978);
nand UO_1206 (O_1206,N_19835,N_19692);
and UO_1207 (O_1207,N_19525,N_19505);
and UO_1208 (O_1208,N_19865,N_19732);
nand UO_1209 (O_1209,N_19862,N_19621);
and UO_1210 (O_1210,N_19704,N_19677);
and UO_1211 (O_1211,N_19564,N_19748);
nand UO_1212 (O_1212,N_19563,N_19795);
nor UO_1213 (O_1213,N_19555,N_19979);
and UO_1214 (O_1214,N_19801,N_19567);
or UO_1215 (O_1215,N_19807,N_19961);
xnor UO_1216 (O_1216,N_19619,N_19582);
nand UO_1217 (O_1217,N_19529,N_19606);
or UO_1218 (O_1218,N_19601,N_19884);
nor UO_1219 (O_1219,N_19818,N_19924);
xor UO_1220 (O_1220,N_19750,N_19927);
xor UO_1221 (O_1221,N_19556,N_19907);
xor UO_1222 (O_1222,N_19521,N_19684);
or UO_1223 (O_1223,N_19784,N_19937);
nand UO_1224 (O_1224,N_19634,N_19907);
xor UO_1225 (O_1225,N_19835,N_19785);
nand UO_1226 (O_1226,N_19567,N_19799);
xor UO_1227 (O_1227,N_19877,N_19700);
xor UO_1228 (O_1228,N_19825,N_19890);
and UO_1229 (O_1229,N_19741,N_19743);
and UO_1230 (O_1230,N_19714,N_19754);
nand UO_1231 (O_1231,N_19628,N_19912);
and UO_1232 (O_1232,N_19891,N_19944);
and UO_1233 (O_1233,N_19570,N_19966);
xnor UO_1234 (O_1234,N_19776,N_19989);
nand UO_1235 (O_1235,N_19783,N_19830);
or UO_1236 (O_1236,N_19552,N_19886);
nor UO_1237 (O_1237,N_19756,N_19801);
and UO_1238 (O_1238,N_19848,N_19716);
nor UO_1239 (O_1239,N_19867,N_19608);
nor UO_1240 (O_1240,N_19552,N_19683);
or UO_1241 (O_1241,N_19959,N_19771);
nand UO_1242 (O_1242,N_19657,N_19870);
nor UO_1243 (O_1243,N_19748,N_19552);
nor UO_1244 (O_1244,N_19601,N_19850);
nor UO_1245 (O_1245,N_19539,N_19820);
nor UO_1246 (O_1246,N_19909,N_19671);
nand UO_1247 (O_1247,N_19620,N_19558);
or UO_1248 (O_1248,N_19959,N_19665);
xor UO_1249 (O_1249,N_19982,N_19913);
nand UO_1250 (O_1250,N_19931,N_19667);
nand UO_1251 (O_1251,N_19654,N_19767);
nand UO_1252 (O_1252,N_19834,N_19948);
xnor UO_1253 (O_1253,N_19885,N_19513);
xnor UO_1254 (O_1254,N_19666,N_19855);
xnor UO_1255 (O_1255,N_19595,N_19572);
nor UO_1256 (O_1256,N_19524,N_19762);
and UO_1257 (O_1257,N_19816,N_19825);
and UO_1258 (O_1258,N_19577,N_19583);
xnor UO_1259 (O_1259,N_19600,N_19924);
xnor UO_1260 (O_1260,N_19515,N_19942);
nand UO_1261 (O_1261,N_19713,N_19782);
xnor UO_1262 (O_1262,N_19554,N_19521);
nor UO_1263 (O_1263,N_19976,N_19925);
or UO_1264 (O_1264,N_19827,N_19786);
nor UO_1265 (O_1265,N_19560,N_19563);
xor UO_1266 (O_1266,N_19574,N_19520);
or UO_1267 (O_1267,N_19572,N_19891);
nor UO_1268 (O_1268,N_19565,N_19823);
or UO_1269 (O_1269,N_19878,N_19996);
xnor UO_1270 (O_1270,N_19905,N_19537);
xor UO_1271 (O_1271,N_19612,N_19898);
nor UO_1272 (O_1272,N_19750,N_19822);
or UO_1273 (O_1273,N_19957,N_19784);
xor UO_1274 (O_1274,N_19941,N_19922);
and UO_1275 (O_1275,N_19568,N_19842);
or UO_1276 (O_1276,N_19631,N_19834);
nand UO_1277 (O_1277,N_19954,N_19662);
xnor UO_1278 (O_1278,N_19844,N_19500);
xor UO_1279 (O_1279,N_19980,N_19625);
or UO_1280 (O_1280,N_19543,N_19522);
xnor UO_1281 (O_1281,N_19987,N_19717);
or UO_1282 (O_1282,N_19683,N_19998);
or UO_1283 (O_1283,N_19540,N_19677);
or UO_1284 (O_1284,N_19867,N_19872);
or UO_1285 (O_1285,N_19659,N_19619);
or UO_1286 (O_1286,N_19823,N_19770);
or UO_1287 (O_1287,N_19534,N_19676);
or UO_1288 (O_1288,N_19774,N_19851);
xnor UO_1289 (O_1289,N_19769,N_19901);
or UO_1290 (O_1290,N_19782,N_19720);
xnor UO_1291 (O_1291,N_19955,N_19993);
nor UO_1292 (O_1292,N_19915,N_19770);
xor UO_1293 (O_1293,N_19570,N_19706);
and UO_1294 (O_1294,N_19726,N_19742);
nor UO_1295 (O_1295,N_19912,N_19508);
nand UO_1296 (O_1296,N_19792,N_19996);
xor UO_1297 (O_1297,N_19805,N_19507);
xor UO_1298 (O_1298,N_19664,N_19627);
or UO_1299 (O_1299,N_19741,N_19746);
nand UO_1300 (O_1300,N_19646,N_19911);
and UO_1301 (O_1301,N_19927,N_19834);
and UO_1302 (O_1302,N_19511,N_19567);
or UO_1303 (O_1303,N_19834,N_19563);
nand UO_1304 (O_1304,N_19822,N_19593);
and UO_1305 (O_1305,N_19826,N_19580);
and UO_1306 (O_1306,N_19555,N_19690);
or UO_1307 (O_1307,N_19558,N_19597);
xnor UO_1308 (O_1308,N_19601,N_19520);
nand UO_1309 (O_1309,N_19635,N_19979);
xnor UO_1310 (O_1310,N_19652,N_19682);
nor UO_1311 (O_1311,N_19919,N_19577);
or UO_1312 (O_1312,N_19985,N_19724);
xnor UO_1313 (O_1313,N_19892,N_19529);
or UO_1314 (O_1314,N_19626,N_19586);
nor UO_1315 (O_1315,N_19522,N_19652);
xnor UO_1316 (O_1316,N_19589,N_19667);
xnor UO_1317 (O_1317,N_19812,N_19889);
or UO_1318 (O_1318,N_19712,N_19726);
xor UO_1319 (O_1319,N_19978,N_19557);
and UO_1320 (O_1320,N_19992,N_19532);
nor UO_1321 (O_1321,N_19760,N_19939);
or UO_1322 (O_1322,N_19851,N_19688);
nor UO_1323 (O_1323,N_19724,N_19971);
nand UO_1324 (O_1324,N_19739,N_19523);
nand UO_1325 (O_1325,N_19851,N_19664);
or UO_1326 (O_1326,N_19883,N_19592);
xnor UO_1327 (O_1327,N_19769,N_19836);
nor UO_1328 (O_1328,N_19865,N_19576);
or UO_1329 (O_1329,N_19684,N_19949);
xor UO_1330 (O_1330,N_19844,N_19534);
nand UO_1331 (O_1331,N_19520,N_19624);
nor UO_1332 (O_1332,N_19729,N_19677);
and UO_1333 (O_1333,N_19996,N_19744);
xnor UO_1334 (O_1334,N_19912,N_19585);
and UO_1335 (O_1335,N_19736,N_19518);
and UO_1336 (O_1336,N_19772,N_19608);
xnor UO_1337 (O_1337,N_19995,N_19799);
nand UO_1338 (O_1338,N_19644,N_19847);
nor UO_1339 (O_1339,N_19651,N_19759);
or UO_1340 (O_1340,N_19869,N_19715);
xnor UO_1341 (O_1341,N_19758,N_19751);
and UO_1342 (O_1342,N_19912,N_19786);
nor UO_1343 (O_1343,N_19585,N_19686);
nand UO_1344 (O_1344,N_19908,N_19540);
and UO_1345 (O_1345,N_19512,N_19886);
and UO_1346 (O_1346,N_19634,N_19560);
nand UO_1347 (O_1347,N_19749,N_19529);
and UO_1348 (O_1348,N_19812,N_19820);
or UO_1349 (O_1349,N_19500,N_19578);
or UO_1350 (O_1350,N_19854,N_19849);
nor UO_1351 (O_1351,N_19592,N_19748);
nand UO_1352 (O_1352,N_19704,N_19751);
nor UO_1353 (O_1353,N_19895,N_19664);
xor UO_1354 (O_1354,N_19755,N_19721);
xnor UO_1355 (O_1355,N_19918,N_19748);
and UO_1356 (O_1356,N_19705,N_19941);
xor UO_1357 (O_1357,N_19753,N_19805);
nor UO_1358 (O_1358,N_19986,N_19785);
or UO_1359 (O_1359,N_19530,N_19865);
xnor UO_1360 (O_1360,N_19876,N_19954);
and UO_1361 (O_1361,N_19812,N_19809);
nand UO_1362 (O_1362,N_19744,N_19940);
nand UO_1363 (O_1363,N_19890,N_19645);
nor UO_1364 (O_1364,N_19886,N_19617);
and UO_1365 (O_1365,N_19730,N_19775);
or UO_1366 (O_1366,N_19647,N_19829);
and UO_1367 (O_1367,N_19758,N_19853);
nand UO_1368 (O_1368,N_19977,N_19666);
nand UO_1369 (O_1369,N_19503,N_19703);
xor UO_1370 (O_1370,N_19518,N_19754);
and UO_1371 (O_1371,N_19603,N_19861);
and UO_1372 (O_1372,N_19695,N_19663);
nor UO_1373 (O_1373,N_19900,N_19846);
nor UO_1374 (O_1374,N_19568,N_19600);
nand UO_1375 (O_1375,N_19721,N_19579);
nand UO_1376 (O_1376,N_19721,N_19920);
and UO_1377 (O_1377,N_19709,N_19927);
nor UO_1378 (O_1378,N_19938,N_19806);
nand UO_1379 (O_1379,N_19709,N_19877);
or UO_1380 (O_1380,N_19627,N_19775);
nor UO_1381 (O_1381,N_19830,N_19611);
nand UO_1382 (O_1382,N_19843,N_19818);
or UO_1383 (O_1383,N_19749,N_19907);
and UO_1384 (O_1384,N_19833,N_19983);
nor UO_1385 (O_1385,N_19931,N_19713);
or UO_1386 (O_1386,N_19711,N_19819);
nand UO_1387 (O_1387,N_19861,N_19805);
nand UO_1388 (O_1388,N_19544,N_19978);
nand UO_1389 (O_1389,N_19667,N_19698);
and UO_1390 (O_1390,N_19716,N_19661);
nor UO_1391 (O_1391,N_19804,N_19849);
xnor UO_1392 (O_1392,N_19743,N_19846);
nor UO_1393 (O_1393,N_19975,N_19991);
nor UO_1394 (O_1394,N_19729,N_19586);
xor UO_1395 (O_1395,N_19782,N_19761);
and UO_1396 (O_1396,N_19807,N_19731);
xor UO_1397 (O_1397,N_19800,N_19785);
xnor UO_1398 (O_1398,N_19687,N_19845);
or UO_1399 (O_1399,N_19754,N_19647);
and UO_1400 (O_1400,N_19869,N_19799);
and UO_1401 (O_1401,N_19613,N_19990);
and UO_1402 (O_1402,N_19527,N_19574);
and UO_1403 (O_1403,N_19881,N_19845);
and UO_1404 (O_1404,N_19750,N_19952);
or UO_1405 (O_1405,N_19715,N_19971);
nor UO_1406 (O_1406,N_19623,N_19706);
xor UO_1407 (O_1407,N_19644,N_19665);
nand UO_1408 (O_1408,N_19829,N_19824);
or UO_1409 (O_1409,N_19510,N_19669);
and UO_1410 (O_1410,N_19580,N_19805);
nor UO_1411 (O_1411,N_19557,N_19923);
xnor UO_1412 (O_1412,N_19953,N_19684);
or UO_1413 (O_1413,N_19917,N_19679);
nand UO_1414 (O_1414,N_19909,N_19809);
nor UO_1415 (O_1415,N_19907,N_19646);
and UO_1416 (O_1416,N_19876,N_19657);
or UO_1417 (O_1417,N_19875,N_19526);
xnor UO_1418 (O_1418,N_19603,N_19979);
nor UO_1419 (O_1419,N_19709,N_19626);
nand UO_1420 (O_1420,N_19504,N_19773);
or UO_1421 (O_1421,N_19709,N_19867);
nor UO_1422 (O_1422,N_19844,N_19881);
nor UO_1423 (O_1423,N_19883,N_19826);
or UO_1424 (O_1424,N_19716,N_19725);
xnor UO_1425 (O_1425,N_19942,N_19587);
and UO_1426 (O_1426,N_19559,N_19623);
or UO_1427 (O_1427,N_19996,N_19575);
nand UO_1428 (O_1428,N_19869,N_19567);
and UO_1429 (O_1429,N_19836,N_19759);
nor UO_1430 (O_1430,N_19858,N_19924);
nor UO_1431 (O_1431,N_19571,N_19745);
or UO_1432 (O_1432,N_19710,N_19610);
and UO_1433 (O_1433,N_19740,N_19973);
nand UO_1434 (O_1434,N_19647,N_19695);
nor UO_1435 (O_1435,N_19533,N_19668);
nand UO_1436 (O_1436,N_19998,N_19710);
nand UO_1437 (O_1437,N_19794,N_19749);
and UO_1438 (O_1438,N_19955,N_19674);
and UO_1439 (O_1439,N_19944,N_19943);
nand UO_1440 (O_1440,N_19762,N_19705);
nor UO_1441 (O_1441,N_19761,N_19945);
nand UO_1442 (O_1442,N_19554,N_19561);
xor UO_1443 (O_1443,N_19897,N_19649);
xnor UO_1444 (O_1444,N_19627,N_19895);
nor UO_1445 (O_1445,N_19828,N_19902);
nor UO_1446 (O_1446,N_19558,N_19606);
and UO_1447 (O_1447,N_19883,N_19924);
or UO_1448 (O_1448,N_19718,N_19907);
xnor UO_1449 (O_1449,N_19538,N_19524);
nand UO_1450 (O_1450,N_19815,N_19782);
nand UO_1451 (O_1451,N_19980,N_19698);
or UO_1452 (O_1452,N_19808,N_19729);
xor UO_1453 (O_1453,N_19792,N_19856);
nor UO_1454 (O_1454,N_19678,N_19709);
xnor UO_1455 (O_1455,N_19770,N_19921);
nor UO_1456 (O_1456,N_19964,N_19932);
nand UO_1457 (O_1457,N_19828,N_19600);
and UO_1458 (O_1458,N_19635,N_19972);
xor UO_1459 (O_1459,N_19554,N_19541);
nand UO_1460 (O_1460,N_19994,N_19921);
xnor UO_1461 (O_1461,N_19514,N_19751);
xor UO_1462 (O_1462,N_19879,N_19568);
xor UO_1463 (O_1463,N_19646,N_19771);
nand UO_1464 (O_1464,N_19946,N_19552);
and UO_1465 (O_1465,N_19793,N_19600);
xnor UO_1466 (O_1466,N_19542,N_19592);
nor UO_1467 (O_1467,N_19989,N_19941);
xnor UO_1468 (O_1468,N_19642,N_19604);
xor UO_1469 (O_1469,N_19958,N_19911);
xor UO_1470 (O_1470,N_19979,N_19830);
or UO_1471 (O_1471,N_19749,N_19639);
and UO_1472 (O_1472,N_19824,N_19928);
xnor UO_1473 (O_1473,N_19528,N_19999);
or UO_1474 (O_1474,N_19637,N_19748);
nor UO_1475 (O_1475,N_19845,N_19985);
nor UO_1476 (O_1476,N_19553,N_19703);
xor UO_1477 (O_1477,N_19921,N_19527);
xor UO_1478 (O_1478,N_19853,N_19903);
or UO_1479 (O_1479,N_19615,N_19778);
xor UO_1480 (O_1480,N_19669,N_19689);
xnor UO_1481 (O_1481,N_19975,N_19663);
or UO_1482 (O_1482,N_19652,N_19765);
nand UO_1483 (O_1483,N_19711,N_19576);
xor UO_1484 (O_1484,N_19831,N_19903);
nand UO_1485 (O_1485,N_19974,N_19761);
nand UO_1486 (O_1486,N_19649,N_19788);
xnor UO_1487 (O_1487,N_19527,N_19925);
nor UO_1488 (O_1488,N_19938,N_19850);
and UO_1489 (O_1489,N_19909,N_19578);
or UO_1490 (O_1490,N_19724,N_19713);
nand UO_1491 (O_1491,N_19641,N_19600);
xor UO_1492 (O_1492,N_19777,N_19756);
or UO_1493 (O_1493,N_19529,N_19694);
xor UO_1494 (O_1494,N_19914,N_19787);
or UO_1495 (O_1495,N_19861,N_19768);
xnor UO_1496 (O_1496,N_19589,N_19712);
and UO_1497 (O_1497,N_19842,N_19746);
or UO_1498 (O_1498,N_19723,N_19821);
or UO_1499 (O_1499,N_19684,N_19519);
and UO_1500 (O_1500,N_19614,N_19552);
or UO_1501 (O_1501,N_19564,N_19585);
or UO_1502 (O_1502,N_19816,N_19735);
and UO_1503 (O_1503,N_19884,N_19794);
or UO_1504 (O_1504,N_19753,N_19586);
and UO_1505 (O_1505,N_19530,N_19588);
or UO_1506 (O_1506,N_19731,N_19610);
or UO_1507 (O_1507,N_19654,N_19814);
or UO_1508 (O_1508,N_19507,N_19850);
nand UO_1509 (O_1509,N_19640,N_19746);
or UO_1510 (O_1510,N_19877,N_19721);
nor UO_1511 (O_1511,N_19704,N_19995);
and UO_1512 (O_1512,N_19959,N_19767);
nor UO_1513 (O_1513,N_19568,N_19702);
or UO_1514 (O_1514,N_19873,N_19562);
or UO_1515 (O_1515,N_19954,N_19574);
or UO_1516 (O_1516,N_19720,N_19620);
nand UO_1517 (O_1517,N_19711,N_19633);
nor UO_1518 (O_1518,N_19532,N_19625);
and UO_1519 (O_1519,N_19769,N_19743);
or UO_1520 (O_1520,N_19515,N_19555);
nand UO_1521 (O_1521,N_19571,N_19708);
nor UO_1522 (O_1522,N_19655,N_19622);
and UO_1523 (O_1523,N_19807,N_19604);
and UO_1524 (O_1524,N_19987,N_19506);
or UO_1525 (O_1525,N_19555,N_19745);
xnor UO_1526 (O_1526,N_19885,N_19994);
xor UO_1527 (O_1527,N_19541,N_19688);
xor UO_1528 (O_1528,N_19839,N_19823);
nor UO_1529 (O_1529,N_19926,N_19699);
xnor UO_1530 (O_1530,N_19522,N_19706);
and UO_1531 (O_1531,N_19618,N_19538);
or UO_1532 (O_1532,N_19842,N_19698);
nor UO_1533 (O_1533,N_19633,N_19509);
nor UO_1534 (O_1534,N_19760,N_19753);
xnor UO_1535 (O_1535,N_19501,N_19791);
nand UO_1536 (O_1536,N_19971,N_19570);
xnor UO_1537 (O_1537,N_19723,N_19735);
nor UO_1538 (O_1538,N_19966,N_19501);
xor UO_1539 (O_1539,N_19641,N_19584);
nor UO_1540 (O_1540,N_19798,N_19855);
xor UO_1541 (O_1541,N_19862,N_19667);
xor UO_1542 (O_1542,N_19745,N_19991);
nor UO_1543 (O_1543,N_19815,N_19786);
nor UO_1544 (O_1544,N_19639,N_19592);
nor UO_1545 (O_1545,N_19807,N_19940);
nand UO_1546 (O_1546,N_19554,N_19546);
nand UO_1547 (O_1547,N_19813,N_19944);
nand UO_1548 (O_1548,N_19903,N_19806);
and UO_1549 (O_1549,N_19779,N_19567);
nor UO_1550 (O_1550,N_19511,N_19954);
or UO_1551 (O_1551,N_19932,N_19530);
xnor UO_1552 (O_1552,N_19977,N_19829);
xor UO_1553 (O_1553,N_19799,N_19824);
nor UO_1554 (O_1554,N_19628,N_19746);
nand UO_1555 (O_1555,N_19678,N_19799);
nor UO_1556 (O_1556,N_19720,N_19830);
and UO_1557 (O_1557,N_19822,N_19560);
xor UO_1558 (O_1558,N_19502,N_19690);
nand UO_1559 (O_1559,N_19672,N_19597);
xor UO_1560 (O_1560,N_19882,N_19701);
xnor UO_1561 (O_1561,N_19623,N_19837);
xnor UO_1562 (O_1562,N_19689,N_19549);
or UO_1563 (O_1563,N_19903,N_19699);
and UO_1564 (O_1564,N_19665,N_19916);
and UO_1565 (O_1565,N_19911,N_19787);
xnor UO_1566 (O_1566,N_19759,N_19655);
and UO_1567 (O_1567,N_19548,N_19817);
or UO_1568 (O_1568,N_19950,N_19625);
and UO_1569 (O_1569,N_19587,N_19775);
xnor UO_1570 (O_1570,N_19576,N_19814);
nor UO_1571 (O_1571,N_19670,N_19529);
nand UO_1572 (O_1572,N_19522,N_19601);
xnor UO_1573 (O_1573,N_19879,N_19774);
xor UO_1574 (O_1574,N_19705,N_19555);
nor UO_1575 (O_1575,N_19758,N_19735);
nor UO_1576 (O_1576,N_19794,N_19786);
xnor UO_1577 (O_1577,N_19699,N_19690);
xor UO_1578 (O_1578,N_19773,N_19547);
nand UO_1579 (O_1579,N_19562,N_19933);
nor UO_1580 (O_1580,N_19595,N_19514);
and UO_1581 (O_1581,N_19939,N_19890);
xor UO_1582 (O_1582,N_19685,N_19631);
nand UO_1583 (O_1583,N_19984,N_19567);
xor UO_1584 (O_1584,N_19515,N_19620);
and UO_1585 (O_1585,N_19894,N_19962);
and UO_1586 (O_1586,N_19800,N_19908);
or UO_1587 (O_1587,N_19998,N_19818);
nand UO_1588 (O_1588,N_19894,N_19869);
xor UO_1589 (O_1589,N_19596,N_19900);
or UO_1590 (O_1590,N_19880,N_19835);
and UO_1591 (O_1591,N_19724,N_19806);
and UO_1592 (O_1592,N_19579,N_19763);
and UO_1593 (O_1593,N_19551,N_19987);
nand UO_1594 (O_1594,N_19579,N_19547);
nor UO_1595 (O_1595,N_19627,N_19684);
and UO_1596 (O_1596,N_19653,N_19788);
nand UO_1597 (O_1597,N_19866,N_19842);
and UO_1598 (O_1598,N_19964,N_19812);
nand UO_1599 (O_1599,N_19854,N_19548);
nand UO_1600 (O_1600,N_19846,N_19972);
nand UO_1601 (O_1601,N_19915,N_19555);
and UO_1602 (O_1602,N_19757,N_19861);
nor UO_1603 (O_1603,N_19689,N_19716);
xnor UO_1604 (O_1604,N_19965,N_19971);
xor UO_1605 (O_1605,N_19600,N_19968);
nand UO_1606 (O_1606,N_19738,N_19774);
nand UO_1607 (O_1607,N_19898,N_19554);
xor UO_1608 (O_1608,N_19936,N_19755);
and UO_1609 (O_1609,N_19963,N_19578);
or UO_1610 (O_1610,N_19707,N_19526);
xor UO_1611 (O_1611,N_19704,N_19820);
nand UO_1612 (O_1612,N_19986,N_19629);
or UO_1613 (O_1613,N_19952,N_19563);
or UO_1614 (O_1614,N_19921,N_19662);
nand UO_1615 (O_1615,N_19818,N_19752);
xnor UO_1616 (O_1616,N_19519,N_19632);
and UO_1617 (O_1617,N_19544,N_19501);
and UO_1618 (O_1618,N_19691,N_19950);
xor UO_1619 (O_1619,N_19729,N_19685);
nor UO_1620 (O_1620,N_19848,N_19841);
xor UO_1621 (O_1621,N_19984,N_19621);
xnor UO_1622 (O_1622,N_19920,N_19885);
xnor UO_1623 (O_1623,N_19686,N_19902);
nor UO_1624 (O_1624,N_19629,N_19800);
xnor UO_1625 (O_1625,N_19940,N_19701);
or UO_1626 (O_1626,N_19517,N_19687);
or UO_1627 (O_1627,N_19677,N_19863);
or UO_1628 (O_1628,N_19551,N_19967);
nor UO_1629 (O_1629,N_19611,N_19771);
nand UO_1630 (O_1630,N_19859,N_19890);
and UO_1631 (O_1631,N_19998,N_19803);
nor UO_1632 (O_1632,N_19615,N_19752);
or UO_1633 (O_1633,N_19747,N_19893);
nor UO_1634 (O_1634,N_19839,N_19826);
xnor UO_1635 (O_1635,N_19630,N_19546);
nand UO_1636 (O_1636,N_19733,N_19912);
and UO_1637 (O_1637,N_19781,N_19530);
nor UO_1638 (O_1638,N_19598,N_19554);
and UO_1639 (O_1639,N_19569,N_19917);
or UO_1640 (O_1640,N_19739,N_19991);
or UO_1641 (O_1641,N_19730,N_19767);
or UO_1642 (O_1642,N_19988,N_19727);
nand UO_1643 (O_1643,N_19702,N_19762);
xnor UO_1644 (O_1644,N_19986,N_19851);
nand UO_1645 (O_1645,N_19657,N_19791);
nor UO_1646 (O_1646,N_19990,N_19655);
and UO_1647 (O_1647,N_19953,N_19584);
nor UO_1648 (O_1648,N_19629,N_19820);
nand UO_1649 (O_1649,N_19817,N_19913);
nand UO_1650 (O_1650,N_19839,N_19858);
nor UO_1651 (O_1651,N_19583,N_19809);
and UO_1652 (O_1652,N_19707,N_19611);
xnor UO_1653 (O_1653,N_19991,N_19974);
nand UO_1654 (O_1654,N_19519,N_19897);
or UO_1655 (O_1655,N_19695,N_19934);
or UO_1656 (O_1656,N_19593,N_19972);
nand UO_1657 (O_1657,N_19788,N_19889);
nand UO_1658 (O_1658,N_19655,N_19781);
nor UO_1659 (O_1659,N_19926,N_19538);
and UO_1660 (O_1660,N_19850,N_19721);
or UO_1661 (O_1661,N_19999,N_19962);
nor UO_1662 (O_1662,N_19675,N_19574);
nor UO_1663 (O_1663,N_19915,N_19501);
or UO_1664 (O_1664,N_19698,N_19521);
or UO_1665 (O_1665,N_19663,N_19998);
nand UO_1666 (O_1666,N_19556,N_19707);
or UO_1667 (O_1667,N_19947,N_19554);
nor UO_1668 (O_1668,N_19706,N_19800);
nand UO_1669 (O_1669,N_19680,N_19714);
nand UO_1670 (O_1670,N_19993,N_19642);
nand UO_1671 (O_1671,N_19627,N_19944);
xor UO_1672 (O_1672,N_19832,N_19817);
or UO_1673 (O_1673,N_19841,N_19747);
or UO_1674 (O_1674,N_19933,N_19865);
or UO_1675 (O_1675,N_19529,N_19712);
nor UO_1676 (O_1676,N_19997,N_19764);
or UO_1677 (O_1677,N_19671,N_19869);
nor UO_1678 (O_1678,N_19511,N_19867);
or UO_1679 (O_1679,N_19819,N_19864);
or UO_1680 (O_1680,N_19661,N_19861);
xnor UO_1681 (O_1681,N_19618,N_19530);
nand UO_1682 (O_1682,N_19965,N_19567);
nand UO_1683 (O_1683,N_19969,N_19687);
and UO_1684 (O_1684,N_19624,N_19598);
xor UO_1685 (O_1685,N_19652,N_19729);
nor UO_1686 (O_1686,N_19718,N_19944);
nor UO_1687 (O_1687,N_19797,N_19813);
and UO_1688 (O_1688,N_19678,N_19861);
nor UO_1689 (O_1689,N_19712,N_19558);
nand UO_1690 (O_1690,N_19605,N_19563);
nand UO_1691 (O_1691,N_19641,N_19974);
or UO_1692 (O_1692,N_19685,N_19799);
nor UO_1693 (O_1693,N_19804,N_19783);
and UO_1694 (O_1694,N_19781,N_19995);
or UO_1695 (O_1695,N_19842,N_19785);
and UO_1696 (O_1696,N_19963,N_19921);
or UO_1697 (O_1697,N_19643,N_19523);
nor UO_1698 (O_1698,N_19841,N_19899);
nand UO_1699 (O_1699,N_19583,N_19547);
nand UO_1700 (O_1700,N_19941,N_19522);
nand UO_1701 (O_1701,N_19580,N_19572);
nand UO_1702 (O_1702,N_19962,N_19980);
or UO_1703 (O_1703,N_19533,N_19856);
nor UO_1704 (O_1704,N_19536,N_19556);
nor UO_1705 (O_1705,N_19692,N_19968);
or UO_1706 (O_1706,N_19713,N_19617);
or UO_1707 (O_1707,N_19516,N_19606);
and UO_1708 (O_1708,N_19517,N_19692);
and UO_1709 (O_1709,N_19851,N_19575);
nand UO_1710 (O_1710,N_19621,N_19663);
xor UO_1711 (O_1711,N_19918,N_19599);
xor UO_1712 (O_1712,N_19632,N_19776);
or UO_1713 (O_1713,N_19503,N_19565);
nor UO_1714 (O_1714,N_19944,N_19875);
xnor UO_1715 (O_1715,N_19777,N_19945);
nand UO_1716 (O_1716,N_19808,N_19904);
or UO_1717 (O_1717,N_19845,N_19534);
and UO_1718 (O_1718,N_19590,N_19514);
nand UO_1719 (O_1719,N_19534,N_19500);
or UO_1720 (O_1720,N_19697,N_19543);
or UO_1721 (O_1721,N_19540,N_19891);
and UO_1722 (O_1722,N_19606,N_19920);
nor UO_1723 (O_1723,N_19962,N_19602);
and UO_1724 (O_1724,N_19547,N_19887);
xnor UO_1725 (O_1725,N_19946,N_19861);
nor UO_1726 (O_1726,N_19712,N_19626);
nand UO_1727 (O_1727,N_19923,N_19595);
nand UO_1728 (O_1728,N_19802,N_19857);
nand UO_1729 (O_1729,N_19939,N_19689);
and UO_1730 (O_1730,N_19706,N_19893);
nand UO_1731 (O_1731,N_19753,N_19746);
or UO_1732 (O_1732,N_19656,N_19871);
or UO_1733 (O_1733,N_19981,N_19842);
or UO_1734 (O_1734,N_19527,N_19663);
xnor UO_1735 (O_1735,N_19833,N_19779);
or UO_1736 (O_1736,N_19693,N_19510);
and UO_1737 (O_1737,N_19809,N_19790);
and UO_1738 (O_1738,N_19942,N_19675);
or UO_1739 (O_1739,N_19880,N_19555);
nor UO_1740 (O_1740,N_19990,N_19695);
and UO_1741 (O_1741,N_19773,N_19537);
nand UO_1742 (O_1742,N_19823,N_19707);
nor UO_1743 (O_1743,N_19696,N_19925);
nor UO_1744 (O_1744,N_19766,N_19943);
or UO_1745 (O_1745,N_19650,N_19731);
xnor UO_1746 (O_1746,N_19953,N_19934);
nor UO_1747 (O_1747,N_19513,N_19978);
nand UO_1748 (O_1748,N_19937,N_19696);
or UO_1749 (O_1749,N_19505,N_19919);
nor UO_1750 (O_1750,N_19876,N_19932);
nor UO_1751 (O_1751,N_19822,N_19825);
nand UO_1752 (O_1752,N_19727,N_19633);
nor UO_1753 (O_1753,N_19779,N_19776);
nor UO_1754 (O_1754,N_19559,N_19618);
nand UO_1755 (O_1755,N_19549,N_19713);
xor UO_1756 (O_1756,N_19684,N_19991);
xor UO_1757 (O_1757,N_19733,N_19615);
nand UO_1758 (O_1758,N_19960,N_19620);
nor UO_1759 (O_1759,N_19676,N_19553);
and UO_1760 (O_1760,N_19707,N_19619);
or UO_1761 (O_1761,N_19692,N_19715);
nand UO_1762 (O_1762,N_19583,N_19713);
xnor UO_1763 (O_1763,N_19727,N_19936);
nor UO_1764 (O_1764,N_19528,N_19794);
xnor UO_1765 (O_1765,N_19937,N_19815);
nor UO_1766 (O_1766,N_19590,N_19898);
or UO_1767 (O_1767,N_19615,N_19589);
xnor UO_1768 (O_1768,N_19574,N_19502);
xor UO_1769 (O_1769,N_19898,N_19760);
and UO_1770 (O_1770,N_19960,N_19536);
and UO_1771 (O_1771,N_19510,N_19689);
nor UO_1772 (O_1772,N_19633,N_19732);
nor UO_1773 (O_1773,N_19780,N_19598);
nand UO_1774 (O_1774,N_19825,N_19949);
and UO_1775 (O_1775,N_19516,N_19712);
xnor UO_1776 (O_1776,N_19955,N_19659);
and UO_1777 (O_1777,N_19562,N_19842);
or UO_1778 (O_1778,N_19839,N_19680);
or UO_1779 (O_1779,N_19884,N_19516);
and UO_1780 (O_1780,N_19811,N_19983);
nand UO_1781 (O_1781,N_19539,N_19835);
nand UO_1782 (O_1782,N_19765,N_19585);
and UO_1783 (O_1783,N_19967,N_19816);
nor UO_1784 (O_1784,N_19797,N_19716);
nand UO_1785 (O_1785,N_19671,N_19875);
xor UO_1786 (O_1786,N_19893,N_19515);
xor UO_1787 (O_1787,N_19654,N_19694);
xor UO_1788 (O_1788,N_19530,N_19774);
nor UO_1789 (O_1789,N_19719,N_19821);
or UO_1790 (O_1790,N_19579,N_19590);
nand UO_1791 (O_1791,N_19628,N_19669);
nor UO_1792 (O_1792,N_19658,N_19548);
or UO_1793 (O_1793,N_19830,N_19625);
nor UO_1794 (O_1794,N_19552,N_19674);
or UO_1795 (O_1795,N_19533,N_19661);
nand UO_1796 (O_1796,N_19545,N_19509);
or UO_1797 (O_1797,N_19852,N_19961);
nand UO_1798 (O_1798,N_19699,N_19553);
nor UO_1799 (O_1799,N_19649,N_19777);
xor UO_1800 (O_1800,N_19594,N_19794);
xnor UO_1801 (O_1801,N_19860,N_19560);
xnor UO_1802 (O_1802,N_19547,N_19662);
xor UO_1803 (O_1803,N_19722,N_19605);
or UO_1804 (O_1804,N_19637,N_19757);
xor UO_1805 (O_1805,N_19852,N_19696);
and UO_1806 (O_1806,N_19591,N_19794);
xor UO_1807 (O_1807,N_19894,N_19644);
nand UO_1808 (O_1808,N_19797,N_19698);
nand UO_1809 (O_1809,N_19726,N_19782);
and UO_1810 (O_1810,N_19817,N_19709);
and UO_1811 (O_1811,N_19631,N_19515);
nor UO_1812 (O_1812,N_19971,N_19963);
nor UO_1813 (O_1813,N_19508,N_19956);
or UO_1814 (O_1814,N_19847,N_19632);
xnor UO_1815 (O_1815,N_19893,N_19558);
or UO_1816 (O_1816,N_19734,N_19904);
or UO_1817 (O_1817,N_19698,N_19927);
nand UO_1818 (O_1818,N_19673,N_19962);
and UO_1819 (O_1819,N_19776,N_19599);
nor UO_1820 (O_1820,N_19583,N_19591);
nand UO_1821 (O_1821,N_19664,N_19761);
and UO_1822 (O_1822,N_19783,N_19750);
nand UO_1823 (O_1823,N_19587,N_19694);
nor UO_1824 (O_1824,N_19809,N_19752);
or UO_1825 (O_1825,N_19937,N_19541);
and UO_1826 (O_1826,N_19842,N_19897);
nand UO_1827 (O_1827,N_19856,N_19714);
xor UO_1828 (O_1828,N_19646,N_19723);
or UO_1829 (O_1829,N_19549,N_19538);
xor UO_1830 (O_1830,N_19736,N_19558);
and UO_1831 (O_1831,N_19512,N_19562);
nand UO_1832 (O_1832,N_19776,N_19590);
xor UO_1833 (O_1833,N_19526,N_19753);
nor UO_1834 (O_1834,N_19554,N_19985);
nand UO_1835 (O_1835,N_19680,N_19706);
nor UO_1836 (O_1836,N_19565,N_19558);
xnor UO_1837 (O_1837,N_19847,N_19535);
nand UO_1838 (O_1838,N_19951,N_19968);
or UO_1839 (O_1839,N_19980,N_19568);
nor UO_1840 (O_1840,N_19747,N_19564);
nand UO_1841 (O_1841,N_19859,N_19633);
or UO_1842 (O_1842,N_19797,N_19833);
and UO_1843 (O_1843,N_19810,N_19950);
or UO_1844 (O_1844,N_19656,N_19797);
nor UO_1845 (O_1845,N_19969,N_19786);
and UO_1846 (O_1846,N_19946,N_19906);
and UO_1847 (O_1847,N_19552,N_19793);
or UO_1848 (O_1848,N_19750,N_19805);
or UO_1849 (O_1849,N_19501,N_19718);
nand UO_1850 (O_1850,N_19647,N_19546);
nor UO_1851 (O_1851,N_19532,N_19588);
or UO_1852 (O_1852,N_19599,N_19981);
nand UO_1853 (O_1853,N_19919,N_19891);
nand UO_1854 (O_1854,N_19905,N_19645);
or UO_1855 (O_1855,N_19605,N_19795);
nor UO_1856 (O_1856,N_19903,N_19727);
or UO_1857 (O_1857,N_19800,N_19500);
or UO_1858 (O_1858,N_19971,N_19512);
or UO_1859 (O_1859,N_19810,N_19637);
and UO_1860 (O_1860,N_19864,N_19779);
and UO_1861 (O_1861,N_19732,N_19804);
or UO_1862 (O_1862,N_19661,N_19602);
xnor UO_1863 (O_1863,N_19967,N_19832);
and UO_1864 (O_1864,N_19637,N_19594);
nand UO_1865 (O_1865,N_19592,N_19664);
xnor UO_1866 (O_1866,N_19986,N_19814);
or UO_1867 (O_1867,N_19919,N_19602);
and UO_1868 (O_1868,N_19609,N_19979);
and UO_1869 (O_1869,N_19799,N_19653);
nand UO_1870 (O_1870,N_19851,N_19866);
or UO_1871 (O_1871,N_19852,N_19510);
and UO_1872 (O_1872,N_19582,N_19672);
nor UO_1873 (O_1873,N_19908,N_19512);
or UO_1874 (O_1874,N_19875,N_19579);
and UO_1875 (O_1875,N_19578,N_19607);
or UO_1876 (O_1876,N_19632,N_19762);
nor UO_1877 (O_1877,N_19564,N_19679);
xnor UO_1878 (O_1878,N_19697,N_19906);
xor UO_1879 (O_1879,N_19841,N_19663);
or UO_1880 (O_1880,N_19932,N_19767);
nand UO_1881 (O_1881,N_19854,N_19503);
nand UO_1882 (O_1882,N_19973,N_19915);
nand UO_1883 (O_1883,N_19675,N_19893);
nand UO_1884 (O_1884,N_19848,N_19777);
or UO_1885 (O_1885,N_19588,N_19933);
nor UO_1886 (O_1886,N_19886,N_19736);
xor UO_1887 (O_1887,N_19715,N_19770);
nand UO_1888 (O_1888,N_19840,N_19866);
and UO_1889 (O_1889,N_19664,N_19970);
or UO_1890 (O_1890,N_19524,N_19872);
or UO_1891 (O_1891,N_19618,N_19546);
nor UO_1892 (O_1892,N_19777,N_19738);
nor UO_1893 (O_1893,N_19954,N_19627);
nor UO_1894 (O_1894,N_19857,N_19910);
xnor UO_1895 (O_1895,N_19764,N_19874);
nor UO_1896 (O_1896,N_19638,N_19667);
nand UO_1897 (O_1897,N_19964,N_19824);
xor UO_1898 (O_1898,N_19623,N_19681);
nor UO_1899 (O_1899,N_19620,N_19772);
nor UO_1900 (O_1900,N_19885,N_19808);
and UO_1901 (O_1901,N_19817,N_19779);
and UO_1902 (O_1902,N_19678,N_19735);
xor UO_1903 (O_1903,N_19709,N_19676);
xor UO_1904 (O_1904,N_19519,N_19997);
or UO_1905 (O_1905,N_19573,N_19850);
xnor UO_1906 (O_1906,N_19619,N_19676);
xnor UO_1907 (O_1907,N_19998,N_19874);
nor UO_1908 (O_1908,N_19633,N_19969);
xnor UO_1909 (O_1909,N_19631,N_19625);
xnor UO_1910 (O_1910,N_19861,N_19952);
and UO_1911 (O_1911,N_19950,N_19555);
nand UO_1912 (O_1912,N_19613,N_19527);
nand UO_1913 (O_1913,N_19523,N_19708);
nand UO_1914 (O_1914,N_19736,N_19516);
and UO_1915 (O_1915,N_19573,N_19870);
nand UO_1916 (O_1916,N_19975,N_19837);
xnor UO_1917 (O_1917,N_19962,N_19992);
or UO_1918 (O_1918,N_19851,N_19731);
and UO_1919 (O_1919,N_19592,N_19744);
and UO_1920 (O_1920,N_19529,N_19969);
nand UO_1921 (O_1921,N_19781,N_19845);
nand UO_1922 (O_1922,N_19956,N_19582);
and UO_1923 (O_1923,N_19944,N_19503);
or UO_1924 (O_1924,N_19529,N_19613);
nor UO_1925 (O_1925,N_19781,N_19772);
xor UO_1926 (O_1926,N_19562,N_19570);
nand UO_1927 (O_1927,N_19636,N_19886);
nor UO_1928 (O_1928,N_19841,N_19631);
xor UO_1929 (O_1929,N_19809,N_19581);
nand UO_1930 (O_1930,N_19856,N_19576);
xnor UO_1931 (O_1931,N_19775,N_19679);
or UO_1932 (O_1932,N_19679,N_19552);
xnor UO_1933 (O_1933,N_19759,N_19774);
or UO_1934 (O_1934,N_19985,N_19938);
xor UO_1935 (O_1935,N_19674,N_19500);
and UO_1936 (O_1936,N_19505,N_19774);
or UO_1937 (O_1937,N_19929,N_19681);
xor UO_1938 (O_1938,N_19787,N_19696);
xnor UO_1939 (O_1939,N_19993,N_19842);
nand UO_1940 (O_1940,N_19973,N_19673);
nor UO_1941 (O_1941,N_19627,N_19500);
or UO_1942 (O_1942,N_19624,N_19672);
or UO_1943 (O_1943,N_19665,N_19885);
or UO_1944 (O_1944,N_19552,N_19595);
nor UO_1945 (O_1945,N_19781,N_19872);
xnor UO_1946 (O_1946,N_19600,N_19523);
and UO_1947 (O_1947,N_19964,N_19830);
nand UO_1948 (O_1948,N_19918,N_19728);
and UO_1949 (O_1949,N_19775,N_19869);
xnor UO_1950 (O_1950,N_19534,N_19608);
and UO_1951 (O_1951,N_19537,N_19521);
nor UO_1952 (O_1952,N_19728,N_19655);
or UO_1953 (O_1953,N_19844,N_19672);
xnor UO_1954 (O_1954,N_19543,N_19822);
nand UO_1955 (O_1955,N_19849,N_19701);
xor UO_1956 (O_1956,N_19986,N_19908);
and UO_1957 (O_1957,N_19583,N_19795);
nand UO_1958 (O_1958,N_19565,N_19905);
nand UO_1959 (O_1959,N_19999,N_19766);
nand UO_1960 (O_1960,N_19969,N_19877);
and UO_1961 (O_1961,N_19566,N_19571);
xnor UO_1962 (O_1962,N_19796,N_19692);
nand UO_1963 (O_1963,N_19513,N_19722);
xor UO_1964 (O_1964,N_19793,N_19517);
and UO_1965 (O_1965,N_19580,N_19648);
nor UO_1966 (O_1966,N_19839,N_19831);
xnor UO_1967 (O_1967,N_19898,N_19646);
nand UO_1968 (O_1968,N_19507,N_19577);
and UO_1969 (O_1969,N_19813,N_19986);
nor UO_1970 (O_1970,N_19873,N_19693);
xor UO_1971 (O_1971,N_19562,N_19730);
xnor UO_1972 (O_1972,N_19975,N_19955);
nor UO_1973 (O_1973,N_19824,N_19675);
nand UO_1974 (O_1974,N_19676,N_19852);
nor UO_1975 (O_1975,N_19532,N_19809);
xnor UO_1976 (O_1976,N_19531,N_19661);
nor UO_1977 (O_1977,N_19857,N_19515);
nor UO_1978 (O_1978,N_19790,N_19864);
xor UO_1979 (O_1979,N_19911,N_19515);
nand UO_1980 (O_1980,N_19759,N_19867);
or UO_1981 (O_1981,N_19638,N_19783);
and UO_1982 (O_1982,N_19785,N_19706);
nor UO_1983 (O_1983,N_19530,N_19769);
nand UO_1984 (O_1984,N_19958,N_19711);
xnor UO_1985 (O_1985,N_19800,N_19747);
and UO_1986 (O_1986,N_19941,N_19595);
and UO_1987 (O_1987,N_19699,N_19836);
nand UO_1988 (O_1988,N_19511,N_19944);
xor UO_1989 (O_1989,N_19977,N_19707);
xor UO_1990 (O_1990,N_19693,N_19772);
xnor UO_1991 (O_1991,N_19676,N_19954);
and UO_1992 (O_1992,N_19887,N_19852);
or UO_1993 (O_1993,N_19819,N_19587);
xor UO_1994 (O_1994,N_19746,N_19707);
nand UO_1995 (O_1995,N_19990,N_19951);
nor UO_1996 (O_1996,N_19836,N_19665);
xor UO_1997 (O_1997,N_19881,N_19623);
nor UO_1998 (O_1998,N_19726,N_19554);
nor UO_1999 (O_1999,N_19680,N_19906);
xnor UO_2000 (O_2000,N_19824,N_19546);
nand UO_2001 (O_2001,N_19643,N_19597);
and UO_2002 (O_2002,N_19579,N_19805);
or UO_2003 (O_2003,N_19641,N_19626);
xnor UO_2004 (O_2004,N_19820,N_19854);
and UO_2005 (O_2005,N_19535,N_19590);
xnor UO_2006 (O_2006,N_19972,N_19750);
or UO_2007 (O_2007,N_19520,N_19652);
or UO_2008 (O_2008,N_19550,N_19969);
nand UO_2009 (O_2009,N_19846,N_19572);
xor UO_2010 (O_2010,N_19570,N_19692);
or UO_2011 (O_2011,N_19519,N_19736);
or UO_2012 (O_2012,N_19958,N_19977);
nor UO_2013 (O_2013,N_19918,N_19944);
nand UO_2014 (O_2014,N_19705,N_19831);
or UO_2015 (O_2015,N_19869,N_19586);
nand UO_2016 (O_2016,N_19754,N_19577);
nand UO_2017 (O_2017,N_19785,N_19554);
and UO_2018 (O_2018,N_19838,N_19669);
nor UO_2019 (O_2019,N_19703,N_19926);
xnor UO_2020 (O_2020,N_19738,N_19764);
and UO_2021 (O_2021,N_19617,N_19574);
nor UO_2022 (O_2022,N_19711,N_19522);
and UO_2023 (O_2023,N_19627,N_19847);
nor UO_2024 (O_2024,N_19771,N_19935);
nand UO_2025 (O_2025,N_19516,N_19659);
nand UO_2026 (O_2026,N_19628,N_19770);
nor UO_2027 (O_2027,N_19764,N_19590);
nor UO_2028 (O_2028,N_19874,N_19504);
nand UO_2029 (O_2029,N_19997,N_19804);
and UO_2030 (O_2030,N_19825,N_19623);
nand UO_2031 (O_2031,N_19741,N_19618);
nor UO_2032 (O_2032,N_19527,N_19958);
nand UO_2033 (O_2033,N_19729,N_19659);
xnor UO_2034 (O_2034,N_19847,N_19954);
xor UO_2035 (O_2035,N_19780,N_19810);
nand UO_2036 (O_2036,N_19814,N_19802);
and UO_2037 (O_2037,N_19800,N_19522);
nor UO_2038 (O_2038,N_19977,N_19896);
nor UO_2039 (O_2039,N_19949,N_19930);
nand UO_2040 (O_2040,N_19581,N_19589);
and UO_2041 (O_2041,N_19899,N_19658);
xor UO_2042 (O_2042,N_19558,N_19756);
and UO_2043 (O_2043,N_19993,N_19775);
nand UO_2044 (O_2044,N_19534,N_19527);
or UO_2045 (O_2045,N_19541,N_19623);
nand UO_2046 (O_2046,N_19606,N_19718);
or UO_2047 (O_2047,N_19625,N_19752);
and UO_2048 (O_2048,N_19917,N_19922);
and UO_2049 (O_2049,N_19587,N_19773);
nor UO_2050 (O_2050,N_19575,N_19618);
nor UO_2051 (O_2051,N_19536,N_19889);
or UO_2052 (O_2052,N_19734,N_19620);
or UO_2053 (O_2053,N_19506,N_19507);
nor UO_2054 (O_2054,N_19920,N_19639);
nand UO_2055 (O_2055,N_19528,N_19570);
or UO_2056 (O_2056,N_19557,N_19606);
nor UO_2057 (O_2057,N_19726,N_19659);
nand UO_2058 (O_2058,N_19953,N_19883);
nor UO_2059 (O_2059,N_19967,N_19957);
or UO_2060 (O_2060,N_19888,N_19976);
xnor UO_2061 (O_2061,N_19977,N_19727);
and UO_2062 (O_2062,N_19787,N_19945);
xor UO_2063 (O_2063,N_19556,N_19742);
nand UO_2064 (O_2064,N_19843,N_19820);
nand UO_2065 (O_2065,N_19777,N_19593);
nor UO_2066 (O_2066,N_19879,N_19938);
or UO_2067 (O_2067,N_19962,N_19950);
or UO_2068 (O_2068,N_19702,N_19528);
xnor UO_2069 (O_2069,N_19943,N_19514);
nand UO_2070 (O_2070,N_19835,N_19898);
xnor UO_2071 (O_2071,N_19764,N_19899);
nor UO_2072 (O_2072,N_19694,N_19911);
nor UO_2073 (O_2073,N_19546,N_19501);
nand UO_2074 (O_2074,N_19894,N_19920);
nor UO_2075 (O_2075,N_19522,N_19688);
nand UO_2076 (O_2076,N_19807,N_19817);
nor UO_2077 (O_2077,N_19712,N_19706);
and UO_2078 (O_2078,N_19705,N_19521);
nor UO_2079 (O_2079,N_19903,N_19936);
and UO_2080 (O_2080,N_19870,N_19650);
and UO_2081 (O_2081,N_19514,N_19618);
or UO_2082 (O_2082,N_19858,N_19639);
xor UO_2083 (O_2083,N_19954,N_19693);
and UO_2084 (O_2084,N_19982,N_19961);
xnor UO_2085 (O_2085,N_19910,N_19964);
and UO_2086 (O_2086,N_19612,N_19989);
or UO_2087 (O_2087,N_19643,N_19922);
xor UO_2088 (O_2088,N_19881,N_19960);
nor UO_2089 (O_2089,N_19640,N_19852);
xnor UO_2090 (O_2090,N_19533,N_19561);
or UO_2091 (O_2091,N_19708,N_19946);
nand UO_2092 (O_2092,N_19561,N_19826);
and UO_2093 (O_2093,N_19656,N_19503);
nand UO_2094 (O_2094,N_19562,N_19515);
and UO_2095 (O_2095,N_19774,N_19569);
xor UO_2096 (O_2096,N_19598,N_19762);
xnor UO_2097 (O_2097,N_19788,N_19827);
nand UO_2098 (O_2098,N_19582,N_19655);
or UO_2099 (O_2099,N_19966,N_19863);
or UO_2100 (O_2100,N_19694,N_19641);
and UO_2101 (O_2101,N_19646,N_19613);
nand UO_2102 (O_2102,N_19812,N_19588);
nor UO_2103 (O_2103,N_19831,N_19644);
and UO_2104 (O_2104,N_19888,N_19968);
nor UO_2105 (O_2105,N_19827,N_19567);
or UO_2106 (O_2106,N_19843,N_19505);
or UO_2107 (O_2107,N_19921,N_19632);
and UO_2108 (O_2108,N_19849,N_19954);
nor UO_2109 (O_2109,N_19898,N_19714);
and UO_2110 (O_2110,N_19737,N_19886);
xor UO_2111 (O_2111,N_19910,N_19622);
and UO_2112 (O_2112,N_19599,N_19959);
xor UO_2113 (O_2113,N_19608,N_19890);
nor UO_2114 (O_2114,N_19803,N_19794);
nor UO_2115 (O_2115,N_19995,N_19847);
xnor UO_2116 (O_2116,N_19563,N_19847);
or UO_2117 (O_2117,N_19911,N_19785);
nor UO_2118 (O_2118,N_19517,N_19601);
nand UO_2119 (O_2119,N_19790,N_19876);
xor UO_2120 (O_2120,N_19883,N_19632);
and UO_2121 (O_2121,N_19608,N_19593);
or UO_2122 (O_2122,N_19890,N_19586);
or UO_2123 (O_2123,N_19621,N_19561);
or UO_2124 (O_2124,N_19735,N_19676);
or UO_2125 (O_2125,N_19817,N_19650);
xor UO_2126 (O_2126,N_19705,N_19864);
nor UO_2127 (O_2127,N_19872,N_19758);
or UO_2128 (O_2128,N_19534,N_19807);
or UO_2129 (O_2129,N_19600,N_19607);
nand UO_2130 (O_2130,N_19643,N_19927);
or UO_2131 (O_2131,N_19636,N_19704);
xnor UO_2132 (O_2132,N_19725,N_19989);
nand UO_2133 (O_2133,N_19638,N_19740);
and UO_2134 (O_2134,N_19798,N_19871);
nor UO_2135 (O_2135,N_19828,N_19944);
and UO_2136 (O_2136,N_19830,N_19725);
nand UO_2137 (O_2137,N_19976,N_19918);
or UO_2138 (O_2138,N_19590,N_19729);
nor UO_2139 (O_2139,N_19777,N_19563);
and UO_2140 (O_2140,N_19647,N_19915);
and UO_2141 (O_2141,N_19742,N_19821);
xor UO_2142 (O_2142,N_19883,N_19952);
and UO_2143 (O_2143,N_19800,N_19570);
nand UO_2144 (O_2144,N_19535,N_19828);
or UO_2145 (O_2145,N_19534,N_19573);
nor UO_2146 (O_2146,N_19822,N_19839);
nand UO_2147 (O_2147,N_19558,N_19952);
or UO_2148 (O_2148,N_19930,N_19697);
xor UO_2149 (O_2149,N_19927,N_19794);
nand UO_2150 (O_2150,N_19867,N_19693);
and UO_2151 (O_2151,N_19592,N_19859);
or UO_2152 (O_2152,N_19532,N_19729);
or UO_2153 (O_2153,N_19653,N_19685);
nand UO_2154 (O_2154,N_19891,N_19654);
or UO_2155 (O_2155,N_19694,N_19927);
or UO_2156 (O_2156,N_19934,N_19997);
nand UO_2157 (O_2157,N_19732,N_19871);
or UO_2158 (O_2158,N_19505,N_19860);
xnor UO_2159 (O_2159,N_19642,N_19848);
and UO_2160 (O_2160,N_19863,N_19817);
and UO_2161 (O_2161,N_19984,N_19506);
xor UO_2162 (O_2162,N_19548,N_19969);
or UO_2163 (O_2163,N_19832,N_19553);
and UO_2164 (O_2164,N_19662,N_19722);
and UO_2165 (O_2165,N_19566,N_19710);
and UO_2166 (O_2166,N_19880,N_19909);
and UO_2167 (O_2167,N_19881,N_19692);
or UO_2168 (O_2168,N_19744,N_19871);
nor UO_2169 (O_2169,N_19575,N_19987);
and UO_2170 (O_2170,N_19546,N_19597);
nand UO_2171 (O_2171,N_19745,N_19876);
nor UO_2172 (O_2172,N_19640,N_19772);
and UO_2173 (O_2173,N_19687,N_19891);
and UO_2174 (O_2174,N_19646,N_19619);
and UO_2175 (O_2175,N_19732,N_19972);
or UO_2176 (O_2176,N_19574,N_19615);
xnor UO_2177 (O_2177,N_19860,N_19596);
nor UO_2178 (O_2178,N_19577,N_19960);
or UO_2179 (O_2179,N_19507,N_19857);
nor UO_2180 (O_2180,N_19998,N_19854);
xnor UO_2181 (O_2181,N_19763,N_19724);
xnor UO_2182 (O_2182,N_19750,N_19582);
and UO_2183 (O_2183,N_19514,N_19893);
xnor UO_2184 (O_2184,N_19592,N_19733);
xor UO_2185 (O_2185,N_19719,N_19815);
nand UO_2186 (O_2186,N_19647,N_19645);
xnor UO_2187 (O_2187,N_19966,N_19937);
and UO_2188 (O_2188,N_19845,N_19852);
nor UO_2189 (O_2189,N_19549,N_19719);
xnor UO_2190 (O_2190,N_19664,N_19943);
nor UO_2191 (O_2191,N_19976,N_19554);
xor UO_2192 (O_2192,N_19619,N_19851);
xnor UO_2193 (O_2193,N_19976,N_19682);
nand UO_2194 (O_2194,N_19983,N_19692);
xor UO_2195 (O_2195,N_19573,N_19763);
and UO_2196 (O_2196,N_19680,N_19691);
xnor UO_2197 (O_2197,N_19681,N_19721);
nand UO_2198 (O_2198,N_19584,N_19809);
nor UO_2199 (O_2199,N_19982,N_19645);
xor UO_2200 (O_2200,N_19716,N_19614);
and UO_2201 (O_2201,N_19644,N_19873);
xnor UO_2202 (O_2202,N_19816,N_19898);
and UO_2203 (O_2203,N_19896,N_19567);
or UO_2204 (O_2204,N_19657,N_19566);
and UO_2205 (O_2205,N_19640,N_19540);
nand UO_2206 (O_2206,N_19609,N_19795);
xor UO_2207 (O_2207,N_19613,N_19582);
and UO_2208 (O_2208,N_19872,N_19522);
nor UO_2209 (O_2209,N_19789,N_19690);
xor UO_2210 (O_2210,N_19779,N_19731);
xnor UO_2211 (O_2211,N_19938,N_19551);
nor UO_2212 (O_2212,N_19794,N_19763);
xnor UO_2213 (O_2213,N_19503,N_19899);
nand UO_2214 (O_2214,N_19669,N_19867);
nand UO_2215 (O_2215,N_19604,N_19973);
or UO_2216 (O_2216,N_19879,N_19531);
and UO_2217 (O_2217,N_19863,N_19725);
or UO_2218 (O_2218,N_19705,N_19554);
nor UO_2219 (O_2219,N_19705,N_19631);
xor UO_2220 (O_2220,N_19844,N_19897);
nor UO_2221 (O_2221,N_19856,N_19518);
and UO_2222 (O_2222,N_19811,N_19686);
or UO_2223 (O_2223,N_19522,N_19984);
nor UO_2224 (O_2224,N_19891,N_19772);
or UO_2225 (O_2225,N_19917,N_19840);
xnor UO_2226 (O_2226,N_19910,N_19606);
nand UO_2227 (O_2227,N_19654,N_19942);
nand UO_2228 (O_2228,N_19800,N_19767);
xnor UO_2229 (O_2229,N_19615,N_19662);
and UO_2230 (O_2230,N_19709,N_19896);
nor UO_2231 (O_2231,N_19971,N_19712);
xnor UO_2232 (O_2232,N_19513,N_19516);
nand UO_2233 (O_2233,N_19981,N_19715);
or UO_2234 (O_2234,N_19865,N_19711);
xor UO_2235 (O_2235,N_19574,N_19923);
or UO_2236 (O_2236,N_19836,N_19896);
xnor UO_2237 (O_2237,N_19607,N_19522);
xnor UO_2238 (O_2238,N_19956,N_19714);
and UO_2239 (O_2239,N_19585,N_19559);
or UO_2240 (O_2240,N_19852,N_19853);
nor UO_2241 (O_2241,N_19903,N_19880);
xor UO_2242 (O_2242,N_19552,N_19790);
nor UO_2243 (O_2243,N_19504,N_19811);
nor UO_2244 (O_2244,N_19794,N_19926);
nand UO_2245 (O_2245,N_19520,N_19619);
and UO_2246 (O_2246,N_19881,N_19629);
xor UO_2247 (O_2247,N_19520,N_19783);
xor UO_2248 (O_2248,N_19740,N_19521);
or UO_2249 (O_2249,N_19685,N_19613);
nor UO_2250 (O_2250,N_19540,N_19743);
xnor UO_2251 (O_2251,N_19818,N_19614);
and UO_2252 (O_2252,N_19842,N_19899);
xor UO_2253 (O_2253,N_19607,N_19698);
nor UO_2254 (O_2254,N_19661,N_19973);
xor UO_2255 (O_2255,N_19948,N_19846);
or UO_2256 (O_2256,N_19768,N_19740);
nand UO_2257 (O_2257,N_19683,N_19859);
and UO_2258 (O_2258,N_19634,N_19624);
or UO_2259 (O_2259,N_19594,N_19608);
nor UO_2260 (O_2260,N_19981,N_19661);
and UO_2261 (O_2261,N_19616,N_19920);
nor UO_2262 (O_2262,N_19615,N_19630);
xor UO_2263 (O_2263,N_19720,N_19594);
xnor UO_2264 (O_2264,N_19669,N_19659);
and UO_2265 (O_2265,N_19515,N_19542);
nand UO_2266 (O_2266,N_19725,N_19969);
or UO_2267 (O_2267,N_19802,N_19911);
nand UO_2268 (O_2268,N_19503,N_19582);
or UO_2269 (O_2269,N_19878,N_19611);
nand UO_2270 (O_2270,N_19814,N_19588);
and UO_2271 (O_2271,N_19599,N_19524);
nor UO_2272 (O_2272,N_19905,N_19740);
nand UO_2273 (O_2273,N_19736,N_19871);
nand UO_2274 (O_2274,N_19865,N_19537);
nor UO_2275 (O_2275,N_19713,N_19591);
xnor UO_2276 (O_2276,N_19855,N_19734);
or UO_2277 (O_2277,N_19903,N_19553);
nand UO_2278 (O_2278,N_19625,N_19736);
nand UO_2279 (O_2279,N_19565,N_19652);
nand UO_2280 (O_2280,N_19854,N_19929);
xor UO_2281 (O_2281,N_19685,N_19728);
xnor UO_2282 (O_2282,N_19892,N_19579);
nor UO_2283 (O_2283,N_19548,N_19526);
xnor UO_2284 (O_2284,N_19545,N_19853);
and UO_2285 (O_2285,N_19801,N_19855);
or UO_2286 (O_2286,N_19989,N_19601);
nand UO_2287 (O_2287,N_19819,N_19784);
and UO_2288 (O_2288,N_19955,N_19537);
or UO_2289 (O_2289,N_19646,N_19920);
and UO_2290 (O_2290,N_19839,N_19723);
and UO_2291 (O_2291,N_19920,N_19759);
xnor UO_2292 (O_2292,N_19803,N_19870);
nand UO_2293 (O_2293,N_19884,N_19944);
xnor UO_2294 (O_2294,N_19777,N_19809);
xor UO_2295 (O_2295,N_19784,N_19835);
or UO_2296 (O_2296,N_19543,N_19551);
and UO_2297 (O_2297,N_19909,N_19770);
nor UO_2298 (O_2298,N_19668,N_19692);
xnor UO_2299 (O_2299,N_19865,N_19808);
nor UO_2300 (O_2300,N_19858,N_19760);
nand UO_2301 (O_2301,N_19542,N_19716);
nand UO_2302 (O_2302,N_19981,N_19604);
xor UO_2303 (O_2303,N_19688,N_19973);
nand UO_2304 (O_2304,N_19727,N_19743);
and UO_2305 (O_2305,N_19993,N_19779);
nor UO_2306 (O_2306,N_19992,N_19825);
xnor UO_2307 (O_2307,N_19675,N_19685);
xnor UO_2308 (O_2308,N_19967,N_19820);
and UO_2309 (O_2309,N_19822,N_19990);
nor UO_2310 (O_2310,N_19544,N_19863);
nor UO_2311 (O_2311,N_19792,N_19711);
or UO_2312 (O_2312,N_19836,N_19875);
and UO_2313 (O_2313,N_19843,N_19930);
nor UO_2314 (O_2314,N_19621,N_19906);
nor UO_2315 (O_2315,N_19662,N_19726);
nor UO_2316 (O_2316,N_19947,N_19542);
and UO_2317 (O_2317,N_19702,N_19942);
and UO_2318 (O_2318,N_19580,N_19749);
xnor UO_2319 (O_2319,N_19629,N_19759);
nor UO_2320 (O_2320,N_19812,N_19760);
or UO_2321 (O_2321,N_19891,N_19786);
nor UO_2322 (O_2322,N_19853,N_19888);
nor UO_2323 (O_2323,N_19869,N_19748);
and UO_2324 (O_2324,N_19637,N_19805);
xor UO_2325 (O_2325,N_19952,N_19918);
xor UO_2326 (O_2326,N_19898,N_19670);
and UO_2327 (O_2327,N_19585,N_19773);
nor UO_2328 (O_2328,N_19683,N_19774);
nand UO_2329 (O_2329,N_19899,N_19932);
xor UO_2330 (O_2330,N_19642,N_19524);
or UO_2331 (O_2331,N_19689,N_19571);
nor UO_2332 (O_2332,N_19921,N_19792);
and UO_2333 (O_2333,N_19975,N_19728);
and UO_2334 (O_2334,N_19747,N_19765);
xnor UO_2335 (O_2335,N_19520,N_19568);
xnor UO_2336 (O_2336,N_19802,N_19554);
nand UO_2337 (O_2337,N_19504,N_19640);
xnor UO_2338 (O_2338,N_19662,N_19705);
or UO_2339 (O_2339,N_19575,N_19850);
nand UO_2340 (O_2340,N_19790,N_19877);
and UO_2341 (O_2341,N_19735,N_19850);
or UO_2342 (O_2342,N_19608,N_19861);
nand UO_2343 (O_2343,N_19766,N_19737);
nor UO_2344 (O_2344,N_19847,N_19548);
and UO_2345 (O_2345,N_19681,N_19817);
nand UO_2346 (O_2346,N_19765,N_19844);
or UO_2347 (O_2347,N_19887,N_19986);
xnor UO_2348 (O_2348,N_19960,N_19950);
and UO_2349 (O_2349,N_19642,N_19587);
xnor UO_2350 (O_2350,N_19749,N_19776);
xnor UO_2351 (O_2351,N_19955,N_19629);
or UO_2352 (O_2352,N_19542,N_19831);
and UO_2353 (O_2353,N_19804,N_19782);
or UO_2354 (O_2354,N_19985,N_19949);
or UO_2355 (O_2355,N_19560,N_19660);
or UO_2356 (O_2356,N_19777,N_19757);
or UO_2357 (O_2357,N_19676,N_19890);
nand UO_2358 (O_2358,N_19832,N_19695);
nor UO_2359 (O_2359,N_19697,N_19990);
nor UO_2360 (O_2360,N_19585,N_19883);
nor UO_2361 (O_2361,N_19959,N_19660);
and UO_2362 (O_2362,N_19748,N_19859);
nand UO_2363 (O_2363,N_19921,N_19774);
xor UO_2364 (O_2364,N_19700,N_19736);
or UO_2365 (O_2365,N_19571,N_19829);
nor UO_2366 (O_2366,N_19915,N_19721);
and UO_2367 (O_2367,N_19674,N_19949);
or UO_2368 (O_2368,N_19587,N_19941);
nand UO_2369 (O_2369,N_19558,N_19644);
xor UO_2370 (O_2370,N_19992,N_19720);
xnor UO_2371 (O_2371,N_19785,N_19749);
xor UO_2372 (O_2372,N_19936,N_19843);
xnor UO_2373 (O_2373,N_19858,N_19943);
nor UO_2374 (O_2374,N_19507,N_19774);
nor UO_2375 (O_2375,N_19574,N_19608);
nand UO_2376 (O_2376,N_19683,N_19811);
xnor UO_2377 (O_2377,N_19756,N_19622);
xor UO_2378 (O_2378,N_19662,N_19827);
xor UO_2379 (O_2379,N_19998,N_19909);
nor UO_2380 (O_2380,N_19875,N_19622);
nand UO_2381 (O_2381,N_19910,N_19572);
or UO_2382 (O_2382,N_19759,N_19712);
nand UO_2383 (O_2383,N_19647,N_19749);
nor UO_2384 (O_2384,N_19988,N_19906);
nand UO_2385 (O_2385,N_19507,N_19647);
nand UO_2386 (O_2386,N_19999,N_19619);
or UO_2387 (O_2387,N_19662,N_19851);
or UO_2388 (O_2388,N_19976,N_19803);
and UO_2389 (O_2389,N_19596,N_19843);
nand UO_2390 (O_2390,N_19551,N_19789);
and UO_2391 (O_2391,N_19639,N_19731);
nand UO_2392 (O_2392,N_19851,N_19764);
or UO_2393 (O_2393,N_19859,N_19870);
or UO_2394 (O_2394,N_19596,N_19872);
and UO_2395 (O_2395,N_19839,N_19898);
nor UO_2396 (O_2396,N_19972,N_19960);
nand UO_2397 (O_2397,N_19513,N_19863);
xor UO_2398 (O_2398,N_19952,N_19795);
nand UO_2399 (O_2399,N_19533,N_19795);
or UO_2400 (O_2400,N_19906,N_19548);
nor UO_2401 (O_2401,N_19827,N_19587);
nor UO_2402 (O_2402,N_19797,N_19928);
or UO_2403 (O_2403,N_19533,N_19627);
xnor UO_2404 (O_2404,N_19525,N_19925);
nand UO_2405 (O_2405,N_19680,N_19785);
and UO_2406 (O_2406,N_19919,N_19616);
nand UO_2407 (O_2407,N_19607,N_19512);
nor UO_2408 (O_2408,N_19723,N_19771);
nor UO_2409 (O_2409,N_19926,N_19905);
nand UO_2410 (O_2410,N_19664,N_19989);
xnor UO_2411 (O_2411,N_19528,N_19611);
or UO_2412 (O_2412,N_19980,N_19697);
nand UO_2413 (O_2413,N_19505,N_19706);
and UO_2414 (O_2414,N_19696,N_19919);
and UO_2415 (O_2415,N_19946,N_19826);
and UO_2416 (O_2416,N_19552,N_19698);
nand UO_2417 (O_2417,N_19835,N_19540);
or UO_2418 (O_2418,N_19904,N_19575);
nand UO_2419 (O_2419,N_19545,N_19712);
xnor UO_2420 (O_2420,N_19926,N_19615);
or UO_2421 (O_2421,N_19780,N_19808);
nor UO_2422 (O_2422,N_19709,N_19635);
nand UO_2423 (O_2423,N_19510,N_19864);
nand UO_2424 (O_2424,N_19772,N_19947);
and UO_2425 (O_2425,N_19694,N_19673);
xnor UO_2426 (O_2426,N_19963,N_19905);
nand UO_2427 (O_2427,N_19688,N_19540);
xor UO_2428 (O_2428,N_19749,N_19823);
and UO_2429 (O_2429,N_19650,N_19573);
xor UO_2430 (O_2430,N_19968,N_19945);
nand UO_2431 (O_2431,N_19891,N_19859);
nand UO_2432 (O_2432,N_19920,N_19543);
or UO_2433 (O_2433,N_19778,N_19741);
nor UO_2434 (O_2434,N_19721,N_19514);
or UO_2435 (O_2435,N_19626,N_19563);
or UO_2436 (O_2436,N_19904,N_19672);
nor UO_2437 (O_2437,N_19855,N_19724);
or UO_2438 (O_2438,N_19525,N_19799);
and UO_2439 (O_2439,N_19730,N_19517);
nand UO_2440 (O_2440,N_19927,N_19865);
or UO_2441 (O_2441,N_19817,N_19841);
nor UO_2442 (O_2442,N_19541,N_19905);
xnor UO_2443 (O_2443,N_19730,N_19542);
or UO_2444 (O_2444,N_19762,N_19557);
or UO_2445 (O_2445,N_19724,N_19694);
or UO_2446 (O_2446,N_19842,N_19898);
nand UO_2447 (O_2447,N_19654,N_19917);
and UO_2448 (O_2448,N_19741,N_19678);
or UO_2449 (O_2449,N_19558,N_19967);
xnor UO_2450 (O_2450,N_19800,N_19794);
nor UO_2451 (O_2451,N_19744,N_19776);
or UO_2452 (O_2452,N_19707,N_19904);
or UO_2453 (O_2453,N_19526,N_19661);
and UO_2454 (O_2454,N_19614,N_19996);
and UO_2455 (O_2455,N_19909,N_19547);
and UO_2456 (O_2456,N_19548,N_19834);
or UO_2457 (O_2457,N_19999,N_19557);
xnor UO_2458 (O_2458,N_19933,N_19630);
xor UO_2459 (O_2459,N_19957,N_19814);
xor UO_2460 (O_2460,N_19705,N_19973);
or UO_2461 (O_2461,N_19615,N_19546);
nand UO_2462 (O_2462,N_19587,N_19646);
or UO_2463 (O_2463,N_19535,N_19919);
or UO_2464 (O_2464,N_19667,N_19630);
nor UO_2465 (O_2465,N_19938,N_19795);
or UO_2466 (O_2466,N_19808,N_19876);
and UO_2467 (O_2467,N_19869,N_19850);
nand UO_2468 (O_2468,N_19978,N_19903);
or UO_2469 (O_2469,N_19933,N_19997);
xnor UO_2470 (O_2470,N_19899,N_19866);
xnor UO_2471 (O_2471,N_19892,N_19786);
xnor UO_2472 (O_2472,N_19609,N_19500);
or UO_2473 (O_2473,N_19502,N_19528);
and UO_2474 (O_2474,N_19659,N_19807);
nor UO_2475 (O_2475,N_19683,N_19760);
nor UO_2476 (O_2476,N_19510,N_19918);
and UO_2477 (O_2477,N_19881,N_19652);
xnor UO_2478 (O_2478,N_19903,N_19825);
and UO_2479 (O_2479,N_19569,N_19863);
xor UO_2480 (O_2480,N_19738,N_19708);
nor UO_2481 (O_2481,N_19526,N_19845);
xnor UO_2482 (O_2482,N_19826,N_19852);
or UO_2483 (O_2483,N_19915,N_19734);
nor UO_2484 (O_2484,N_19724,N_19692);
nor UO_2485 (O_2485,N_19746,N_19679);
xor UO_2486 (O_2486,N_19760,N_19631);
or UO_2487 (O_2487,N_19513,N_19964);
xor UO_2488 (O_2488,N_19528,N_19873);
and UO_2489 (O_2489,N_19756,N_19830);
xnor UO_2490 (O_2490,N_19853,N_19807);
xnor UO_2491 (O_2491,N_19747,N_19678);
nor UO_2492 (O_2492,N_19590,N_19627);
nand UO_2493 (O_2493,N_19872,N_19750);
nand UO_2494 (O_2494,N_19745,N_19701);
and UO_2495 (O_2495,N_19683,N_19876);
nand UO_2496 (O_2496,N_19603,N_19996);
xnor UO_2497 (O_2497,N_19652,N_19937);
nand UO_2498 (O_2498,N_19654,N_19819);
nand UO_2499 (O_2499,N_19835,N_19831);
endmodule