module basic_3000_30000_3500_10_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_235,In_2893);
nand U1 (N_1,In_2391,In_1998);
and U2 (N_2,In_2687,In_580);
xor U3 (N_3,In_733,In_800);
or U4 (N_4,In_1790,In_2002);
or U5 (N_5,In_1230,In_1403);
and U6 (N_6,In_2357,In_1139);
and U7 (N_7,In_2888,In_1959);
and U8 (N_8,In_1570,In_1762);
or U9 (N_9,In_946,In_344);
or U10 (N_10,In_2285,In_1127);
and U11 (N_11,In_2151,In_2952);
or U12 (N_12,In_914,In_2602);
and U13 (N_13,In_2239,In_2695);
nand U14 (N_14,In_1591,In_1303);
nor U15 (N_15,In_2551,In_1114);
and U16 (N_16,In_384,In_2286);
or U17 (N_17,In_2934,In_1386);
nor U18 (N_18,In_1796,In_1081);
or U19 (N_19,In_2069,In_2953);
or U20 (N_20,In_2675,In_744);
nand U21 (N_21,In_2577,In_1256);
and U22 (N_22,In_1971,In_939);
nor U23 (N_23,In_988,In_2057);
nor U24 (N_24,In_538,In_2631);
xnor U25 (N_25,In_2298,In_2146);
nand U26 (N_26,In_2714,In_1445);
xnor U27 (N_27,In_2763,In_1311);
nor U28 (N_28,In_984,In_1004);
nand U29 (N_29,In_2486,In_6);
xor U30 (N_30,In_2067,In_2643);
and U31 (N_31,In_2564,In_1773);
xnor U32 (N_32,In_1382,In_2931);
nor U33 (N_33,In_1600,In_58);
nor U34 (N_34,In_2407,In_2751);
xor U35 (N_35,In_2333,In_1638);
or U36 (N_36,In_506,In_743);
nor U37 (N_37,In_1288,In_2670);
nand U38 (N_38,In_481,In_767);
nand U39 (N_39,In_2827,In_1877);
or U40 (N_40,In_1460,In_2375);
nand U41 (N_41,In_2647,In_2388);
and U42 (N_42,In_1070,In_2563);
xnor U43 (N_43,In_1327,In_2196);
nand U44 (N_44,In_992,In_776);
xnor U45 (N_45,In_690,In_2149);
or U46 (N_46,In_1434,In_2024);
and U47 (N_47,In_1952,In_1118);
and U48 (N_48,In_1574,In_2083);
nor U49 (N_49,In_1791,In_868);
and U50 (N_50,In_485,In_1618);
nand U51 (N_51,In_2716,In_2937);
or U52 (N_52,In_1598,In_1116);
nor U53 (N_53,In_704,In_671);
nand U54 (N_54,In_1851,In_106);
xor U55 (N_55,In_1199,In_2955);
xnor U56 (N_56,In_1060,In_127);
xnor U57 (N_57,In_2105,In_53);
xnor U58 (N_58,In_1861,In_1117);
nor U59 (N_59,In_2053,In_1677);
nand U60 (N_60,In_1431,In_2193);
xnor U61 (N_61,In_1398,In_2976);
or U62 (N_62,In_2147,In_1261);
and U63 (N_63,In_2126,In_2240);
and U64 (N_64,In_303,In_634);
or U65 (N_65,In_2543,In_2529);
nand U66 (N_66,In_1358,In_365);
or U67 (N_67,In_172,In_1158);
or U68 (N_68,In_2632,In_2129);
or U69 (N_69,In_2197,In_498);
and U70 (N_70,In_996,In_175);
nand U71 (N_71,In_1897,In_1009);
and U72 (N_72,In_1641,In_537);
and U73 (N_73,In_1713,In_1527);
and U74 (N_74,In_2251,In_624);
nor U75 (N_75,In_1626,In_448);
xnor U76 (N_76,In_1494,In_959);
nand U77 (N_77,In_2779,In_52);
nor U78 (N_78,In_1917,In_19);
or U79 (N_79,In_1976,In_1704);
or U80 (N_80,In_1874,In_1633);
or U81 (N_81,In_846,In_1143);
or U82 (N_82,In_1953,In_1934);
nor U83 (N_83,In_394,In_620);
or U84 (N_84,In_519,In_1340);
xnor U85 (N_85,In_2609,In_1505);
xor U86 (N_86,In_1504,In_1103);
nor U87 (N_87,In_2904,In_281);
nor U88 (N_88,In_663,In_2981);
nand U89 (N_89,In_969,In_760);
and U90 (N_90,In_554,In_1383);
xnor U91 (N_91,In_480,In_551);
and U92 (N_92,In_246,In_1301);
nand U93 (N_93,In_2454,In_525);
xor U94 (N_94,In_1844,In_2153);
nor U95 (N_95,In_1669,In_1548);
nand U96 (N_96,In_2512,In_1599);
nand U97 (N_97,In_2195,In_465);
nor U98 (N_98,In_918,In_2493);
xor U99 (N_99,In_1688,In_129);
or U100 (N_100,In_2079,In_544);
or U101 (N_101,In_120,In_2371);
and U102 (N_102,In_192,In_2299);
nor U103 (N_103,In_2782,In_85);
nand U104 (N_104,In_759,In_1239);
nand U105 (N_105,In_2102,In_37);
or U106 (N_106,In_904,In_247);
and U107 (N_107,In_1942,In_2718);
and U108 (N_108,In_226,In_1449);
or U109 (N_109,In_186,In_1853);
xnor U110 (N_110,In_517,In_131);
xor U111 (N_111,In_2004,In_2132);
nand U112 (N_112,In_1259,In_1663);
nand U113 (N_113,In_524,In_1520);
nor U114 (N_114,In_2206,In_2785);
or U115 (N_115,In_1833,In_2618);
and U116 (N_116,In_2739,In_1958);
nor U117 (N_117,In_2170,In_1067);
xnor U118 (N_118,In_1993,In_732);
nor U119 (N_119,In_2074,In_2294);
or U120 (N_120,In_1296,In_999);
nor U121 (N_121,In_1898,In_2096);
nor U122 (N_122,In_1904,In_1332);
and U123 (N_123,In_1001,In_1342);
nand U124 (N_124,In_1219,In_2844);
nor U125 (N_125,In_169,In_689);
xor U126 (N_126,In_335,In_605);
nand U127 (N_127,In_2379,In_2430);
xor U128 (N_128,In_2778,In_1372);
or U129 (N_129,In_1517,In_1651);
or U130 (N_130,In_266,In_686);
nor U131 (N_131,In_1882,In_1229);
xnor U132 (N_132,In_1975,In_536);
nand U133 (N_133,In_165,In_2011);
or U134 (N_134,In_963,In_2830);
or U135 (N_135,In_2172,In_1203);
xnor U136 (N_136,In_794,In_2982);
nand U137 (N_137,In_2499,In_2709);
nor U138 (N_138,In_2527,In_2349);
or U139 (N_139,In_1888,In_30);
and U140 (N_140,In_463,In_2596);
and U141 (N_141,In_275,In_2732);
nand U142 (N_142,In_2615,In_2317);
nand U143 (N_143,In_63,In_492);
and U144 (N_144,In_1852,In_2015);
nand U145 (N_145,In_2496,In_895);
xnor U146 (N_146,In_2044,In_1606);
or U147 (N_147,In_1472,In_495);
and U148 (N_148,In_2509,In_1697);
nand U149 (N_149,In_3,In_2826);
xnor U150 (N_150,In_39,In_1648);
and U151 (N_151,In_215,In_2211);
nand U152 (N_152,In_156,In_1341);
or U153 (N_153,In_2300,In_190);
nor U154 (N_154,In_2930,In_1385);
and U155 (N_155,In_2429,In_2235);
or U156 (N_156,In_1490,In_66);
nand U157 (N_157,In_137,In_2710);
xnor U158 (N_158,In_1801,In_433);
nand U159 (N_159,In_203,In_1605);
or U160 (N_160,In_1566,In_1929);
or U161 (N_161,In_2896,In_1660);
xor U162 (N_162,In_1152,In_1981);
and U163 (N_163,In_1192,In_881);
xor U164 (N_164,In_2447,In_1918);
xor U165 (N_165,In_726,In_684);
nor U166 (N_166,In_1878,In_1147);
and U167 (N_167,In_483,In_859);
and U168 (N_168,In_1161,In_1830);
and U169 (N_169,In_1099,In_1503);
xor U170 (N_170,In_2162,In_278);
nor U171 (N_171,In_2238,In_1933);
and U172 (N_172,In_807,In_1226);
and U173 (N_173,In_1337,In_429);
xnor U174 (N_174,In_1113,In_1587);
or U175 (N_175,In_673,In_371);
nand U176 (N_176,In_792,In_2503);
and U177 (N_177,In_417,In_936);
nand U178 (N_178,In_2065,In_2008);
nand U179 (N_179,In_602,In_2699);
and U180 (N_180,In_651,In_2702);
nand U181 (N_181,In_2051,In_2722);
xor U182 (N_182,In_7,In_1772);
and U183 (N_183,In_1731,In_1072);
and U184 (N_184,In_2620,In_1642);
and U185 (N_185,In_332,In_450);
nor U186 (N_186,In_2772,In_427);
nor U187 (N_187,In_1565,In_1623);
xnor U188 (N_188,In_228,In_1588);
or U189 (N_189,In_1691,In_2340);
or U190 (N_190,In_1656,In_1695);
and U191 (N_191,In_1966,In_2671);
or U192 (N_192,In_2075,In_2628);
or U193 (N_193,In_665,In_2208);
nor U194 (N_194,In_33,In_2851);
nand U195 (N_195,In_2380,In_2054);
nand U196 (N_196,In_1846,In_2607);
nor U197 (N_197,In_1157,In_1531);
xor U198 (N_198,In_0,In_2591);
xor U199 (N_199,In_1278,In_1196);
nand U200 (N_200,In_2191,In_901);
or U201 (N_201,In_2050,In_2749);
and U202 (N_202,In_2408,In_196);
nor U203 (N_203,In_2917,In_2787);
nor U204 (N_204,In_230,In_2823);
and U205 (N_205,In_1346,In_1041);
nor U206 (N_206,In_2879,In_729);
nor U207 (N_207,In_1115,In_1857);
and U208 (N_208,In_1907,In_900);
nand U209 (N_209,In_2555,In_1859);
and U210 (N_210,In_2692,In_2325);
and U211 (N_211,In_1987,In_1397);
or U212 (N_212,In_73,In_2005);
nor U213 (N_213,In_870,In_415);
nor U214 (N_214,In_557,In_103);
nor U215 (N_215,In_872,In_2320);
or U216 (N_216,In_1596,In_2528);
nand U217 (N_217,In_2436,In_589);
or U218 (N_218,In_1657,In_1951);
xor U219 (N_219,In_2664,In_1568);
xnor U220 (N_220,In_47,In_2201);
or U221 (N_221,In_929,In_838);
nor U222 (N_222,In_979,In_132);
xor U223 (N_223,In_2076,In_2427);
and U224 (N_224,In_82,In_361);
or U225 (N_225,In_750,In_1776);
nor U226 (N_226,In_1572,In_262);
and U227 (N_227,In_385,In_29);
xnor U228 (N_228,In_2257,In_627);
or U229 (N_229,In_1112,In_459);
or U230 (N_230,In_2588,In_507);
or U231 (N_231,In_2434,In_951);
or U232 (N_232,In_2852,In_2979);
or U233 (N_233,In_738,In_314);
nand U234 (N_234,In_2092,In_662);
xnor U235 (N_235,In_2387,In_1575);
xnor U236 (N_236,In_104,In_2167);
nand U237 (N_237,In_1381,In_1124);
xor U238 (N_238,In_2464,In_768);
nand U239 (N_239,In_348,In_380);
nor U240 (N_240,In_326,In_1048);
xnor U241 (N_241,In_2334,In_1206);
xor U242 (N_242,In_143,In_1577);
nor U243 (N_243,In_708,In_1040);
nand U244 (N_244,In_1827,In_421);
and U245 (N_245,In_600,In_1593);
and U246 (N_246,In_1578,In_158);
and U247 (N_247,In_2544,In_1930);
and U248 (N_248,In_721,In_568);
and U249 (N_249,In_2495,In_42);
nor U250 (N_250,In_490,In_840);
nand U251 (N_251,In_1707,In_2697);
nor U252 (N_252,In_1845,In_205);
nor U253 (N_253,In_1684,In_1905);
and U254 (N_254,In_438,In_748);
xnor U255 (N_255,In_76,In_290);
nor U256 (N_256,In_1011,In_173);
or U257 (N_257,In_2541,In_2913);
xor U258 (N_258,In_2255,In_1245);
nor U259 (N_259,In_2237,In_1685);
xor U260 (N_260,In_2242,In_973);
xor U261 (N_261,In_1010,In_2439);
or U262 (N_262,In_112,In_916);
nand U263 (N_263,In_1093,In_2534);
nand U264 (N_264,In_2256,In_256);
or U265 (N_265,In_1780,In_2474);
xnor U266 (N_266,In_224,In_1996);
or U267 (N_267,In_2525,In_234);
nor U268 (N_268,In_2846,In_697);
xor U269 (N_269,In_2225,In_1284);
nand U270 (N_270,In_2222,In_1207);
nor U271 (N_271,In_2511,In_619);
nor U272 (N_272,In_13,In_1002);
or U273 (N_273,In_20,In_2884);
or U274 (N_274,In_1896,In_886);
or U275 (N_275,In_2983,In_2614);
and U276 (N_276,In_2727,In_705);
nand U277 (N_277,In_1887,In_2258);
or U278 (N_278,In_1369,In_2766);
and U279 (N_279,In_1287,In_334);
and U280 (N_280,In_1122,In_1409);
nand U281 (N_281,In_436,In_54);
nor U282 (N_282,In_2022,In_935);
and U283 (N_283,In_2243,In_860);
or U284 (N_284,In_1184,In_2556);
or U285 (N_285,In_2624,In_2154);
nor U286 (N_286,In_390,In_328);
or U287 (N_287,In_640,In_1558);
nor U288 (N_288,In_1603,In_2420);
and U289 (N_289,In_1813,In_1283);
nand U290 (N_290,In_615,In_21);
nand U291 (N_291,In_894,In_55);
xor U292 (N_292,In_2397,In_2677);
nand U293 (N_293,In_1345,In_788);
or U294 (N_294,In_308,In_2794);
or U295 (N_295,In_2106,In_453);
or U296 (N_296,In_2662,In_1266);
xor U297 (N_297,In_1890,In_1766);
and U298 (N_298,In_1077,In_2326);
nand U299 (N_299,In_258,In_231);
and U300 (N_300,In_337,In_2691);
and U301 (N_301,In_1003,In_680);
xor U302 (N_302,In_1995,In_1761);
xnor U303 (N_303,In_1640,In_1771);
nand U304 (N_304,In_995,In_830);
nand U305 (N_305,In_2085,In_786);
and U306 (N_306,In_2116,In_2686);
nor U307 (N_307,In_770,In_1499);
and U308 (N_308,In_608,In_1065);
nor U309 (N_309,In_177,In_631);
nor U310 (N_310,In_577,In_2650);
nor U311 (N_311,In_1734,In_457);
xnor U312 (N_312,In_2306,In_2314);
or U313 (N_313,In_1871,In_116);
and U314 (N_314,In_1592,In_1650);
and U315 (N_315,In_1185,In_787);
nor U316 (N_316,In_1254,In_1447);
or U317 (N_317,In_454,In_2655);
or U318 (N_318,In_820,In_790);
or U319 (N_319,In_410,In_1526);
nand U320 (N_320,In_1849,In_954);
nor U321 (N_321,In_2854,In_2924);
xor U322 (N_322,In_2275,In_1549);
xor U323 (N_323,In_1175,In_2338);
and U324 (N_324,In_1176,In_2033);
nor U325 (N_325,In_724,In_871);
and U326 (N_326,In_312,In_2038);
and U327 (N_327,In_2941,In_1492);
nor U328 (N_328,In_1729,In_353);
and U329 (N_329,In_115,In_2214);
and U330 (N_330,In_796,In_245);
xor U331 (N_331,In_1968,In_1823);
nor U332 (N_332,In_336,In_1220);
nand U333 (N_333,In_2292,In_155);
nor U334 (N_334,In_696,In_771);
xnor U335 (N_335,In_284,In_878);
xor U336 (N_336,In_5,In_2674);
xor U337 (N_337,In_2589,In_2767);
nor U338 (N_338,In_2090,In_700);
nor U339 (N_339,In_2109,In_254);
xnor U340 (N_340,In_289,In_307);
xnor U341 (N_341,In_635,In_2254);
or U342 (N_342,In_906,In_2249);
and U343 (N_343,In_494,In_2121);
nand U344 (N_344,In_1553,In_1310);
nor U345 (N_345,In_1424,In_2426);
xor U346 (N_346,In_730,In_1546);
or U347 (N_347,In_1444,In_1954);
xnor U348 (N_348,In_2019,In_1211);
xnor U349 (N_349,In_1148,In_2756);
nor U350 (N_350,In_502,In_2020);
and U351 (N_351,In_1415,In_2324);
nor U352 (N_352,In_191,In_377);
nor U353 (N_353,In_727,In_1715);
nor U354 (N_354,In_2743,In_473);
and U355 (N_355,In_563,In_1421);
nand U356 (N_356,In_1906,In_86);
nand U357 (N_357,In_1679,In_2419);
xnor U358 (N_358,In_464,In_882);
xor U359 (N_359,In_1810,In_2335);
nor U360 (N_360,In_576,In_1709);
nor U361 (N_361,In_1661,In_2453);
and U362 (N_362,In_822,In_2890);
or U363 (N_363,In_2568,In_2142);
xor U364 (N_364,In_1380,In_2706);
and U365 (N_365,In_88,In_1529);
or U366 (N_366,In_1292,In_1328);
nor U367 (N_367,In_2369,In_720);
xnor U368 (N_368,In_2745,In_2030);
nor U369 (N_369,In_2048,In_2703);
or U370 (N_370,In_2322,In_2497);
and U371 (N_371,In_614,In_1560);
and U372 (N_372,In_1649,In_2283);
nand U373 (N_373,In_1454,In_2409);
nor U374 (N_374,In_2361,In_1528);
xor U375 (N_375,In_220,In_2392);
nand U376 (N_376,In_2797,In_531);
or U377 (N_377,In_1957,In_599);
nand U378 (N_378,In_1330,In_1412);
or U379 (N_379,In_783,In_2715);
xor U380 (N_380,In_123,In_2875);
xor U381 (N_381,In_818,In_1443);
nor U382 (N_382,In_2733,In_823);
and U383 (N_383,In_1921,In_2232);
nor U384 (N_384,In_2344,In_2470);
nand U385 (N_385,In_1052,In_2549);
nor U386 (N_386,In_1702,In_1567);
and U387 (N_387,In_277,In_943);
or U388 (N_388,In_2127,In_342);
or U389 (N_389,In_2672,In_813);
or U390 (N_390,In_1094,In_2049);
nand U391 (N_391,In_675,In_435);
nand U392 (N_392,In_2789,In_2803);
xnor U393 (N_393,In_2784,In_2578);
or U394 (N_394,In_72,In_304);
nor U395 (N_395,In_1922,In_2707);
xnor U396 (N_396,In_296,In_2712);
or U397 (N_397,In_897,In_956);
nor U398 (N_398,In_1119,In_2894);
or U399 (N_399,In_714,In_539);
nand U400 (N_400,In_2180,In_2939);
nand U401 (N_401,In_285,In_1071);
or U402 (N_402,In_1274,In_2912);
nor U403 (N_403,In_409,In_2911);
nand U404 (N_404,In_1387,In_975);
nand U405 (N_405,In_2989,In_2708);
or U406 (N_406,In_1891,In_843);
nand U407 (N_407,In_2422,In_2942);
xnor U408 (N_408,In_808,In_2754);
xnor U409 (N_409,In_1672,In_2533);
and U410 (N_410,In_2035,In_2213);
nand U411 (N_411,In_401,In_1613);
xnor U412 (N_412,In_1585,In_135);
and U413 (N_413,In_2310,In_1051);
nand U414 (N_414,In_1299,In_1498);
nand U415 (N_415,In_1193,In_722);
xor U416 (N_416,In_276,In_2669);
or U417 (N_417,In_2831,In_408);
or U418 (N_418,In_2961,In_562);
and U419 (N_419,In_2762,In_2757);
nand U420 (N_420,In_2156,In_2342);
and U421 (N_421,In_1326,In_2402);
and U422 (N_422,In_1822,In_1180);
nor U423 (N_423,In_2818,In_2176);
and U424 (N_424,In_2508,In_757);
or U425 (N_425,In_2424,In_1120);
nor U426 (N_426,In_319,In_981);
xnor U427 (N_427,In_2560,In_1181);
or U428 (N_428,In_445,In_1769);
and U429 (N_429,In_831,In_1105);
xor U430 (N_430,In_2567,In_1726);
nand U431 (N_431,In_844,In_357);
xnor U432 (N_432,In_18,In_188);
xnor U433 (N_433,In_617,In_2309);
or U434 (N_434,In_2077,In_2903);
and U435 (N_435,In_1485,In_2561);
xor U436 (N_436,In_397,In_148);
or U437 (N_437,In_793,In_2483);
and U438 (N_438,In_236,In_2052);
xor U439 (N_439,In_1418,In_1422);
or U440 (N_440,In_2363,In_1440);
and U441 (N_441,In_1255,In_1770);
xor U442 (N_442,In_2218,In_214);
xnor U443 (N_443,In_1614,In_402);
xor U444 (N_444,In_1243,In_1389);
xnor U445 (N_445,In_1322,In_1821);
nor U446 (N_446,In_10,In_2312);
or U447 (N_447,In_934,In_2362);
xor U448 (N_448,In_2274,In_628);
and U449 (N_449,In_1928,In_1043);
and U450 (N_450,In_2036,In_164);
and U451 (N_451,In_1435,In_1100);
xnor U452 (N_452,In_2804,In_1564);
nor U453 (N_453,In_681,In_1066);
nand U454 (N_454,In_1260,In_171);
nand U455 (N_455,In_2413,In_1069);
nand U456 (N_456,In_1324,In_1583);
nor U457 (N_457,In_734,In_1532);
nor U458 (N_458,In_183,In_755);
or U459 (N_459,In_648,In_2446);
nand U460 (N_460,In_1267,In_1817);
nor U461 (N_461,In_2513,In_287);
xor U462 (N_462,In_2644,In_2223);
xnor U463 (N_463,In_574,In_623);
or U464 (N_464,In_2629,In_1579);
nand U465 (N_465,In_2623,In_1514);
and U466 (N_466,In_1920,In_32);
xnor U467 (N_467,In_508,In_1355);
and U468 (N_468,In_883,In_1559);
and U469 (N_469,In_2788,In_2164);
nor U470 (N_470,In_1253,In_2343);
or U471 (N_471,In_1451,In_2110);
nand U472 (N_472,In_924,In_1076);
and U473 (N_473,In_2452,In_350);
or U474 (N_474,In_251,In_542);
nand U475 (N_475,In_1982,In_2773);
xnor U476 (N_476,In_2072,In_2456);
nand U477 (N_477,In_2117,In_133);
nand U478 (N_478,In_678,In_2954);
or U479 (N_479,In_108,In_2595);
nor U480 (N_480,In_2936,In_1007);
xor U481 (N_481,In_2502,In_2080);
or U482 (N_482,In_828,In_1482);
nor U483 (N_483,In_283,In_2565);
and U484 (N_484,In_2705,In_1123);
xnor U485 (N_485,In_1194,In_1913);
nand U486 (N_486,In_2457,In_1838);
nand U487 (N_487,In_374,In_913);
nor U488 (N_488,In_1885,In_2128);
xnor U489 (N_489,In_105,In_2330);
nor U490 (N_490,In_656,In_2969);
xnor U491 (N_491,In_1902,In_2460);
nor U492 (N_492,In_1997,In_2231);
and U493 (N_493,In_719,In_2832);
or U494 (N_494,In_948,In_889);
or U495 (N_495,In_2667,In_2580);
nand U496 (N_496,In_2160,In_1738);
nand U497 (N_497,In_1252,In_2721);
nor U498 (N_498,In_2995,In_461);
or U499 (N_499,In_499,In_2381);
xnor U500 (N_500,In_1227,In_1733);
or U501 (N_501,In_1536,In_2104);
nand U502 (N_502,In_763,In_1163);
nand U503 (N_503,In_178,In_17);
and U504 (N_504,In_27,In_970);
xor U505 (N_505,In_1675,In_1384);
nand U506 (N_506,In_2654,In_2347);
nand U507 (N_507,In_2498,In_372);
xor U508 (N_508,In_2524,In_921);
or U509 (N_509,In_638,In_399);
nor U510 (N_510,In_211,In_2611);
or U511 (N_511,In_146,In_643);
nand U512 (N_512,In_1487,In_185);
or U513 (N_513,In_2122,In_56);
nor U514 (N_514,In_565,In_2482);
or U515 (N_515,In_735,In_2806);
and U516 (N_516,In_1458,In_1475);
nor U517 (N_517,In_799,In_1319);
or U518 (N_518,In_2210,In_509);
and U519 (N_519,In_2592,In_2130);
nand U520 (N_520,In_2437,In_1883);
and U521 (N_521,In_273,In_1231);
nor U522 (N_522,In_1017,In_543);
nand U523 (N_523,In_2881,In_141);
or U524 (N_524,In_1016,In_1716);
xnor U525 (N_525,In_1742,In_2501);
or U526 (N_526,In_1291,In_1177);
or U527 (N_527,In_219,In_102);
or U528 (N_528,In_1257,In_2405);
or U529 (N_529,In_2451,In_34);
nand U530 (N_530,In_1831,In_1625);
nand U531 (N_531,In_2886,In_1144);
or U532 (N_532,In_902,In_751);
xnor U533 (N_533,In_2382,In_611);
nand U534 (N_534,In_1753,In_2966);
xor U535 (N_535,In_937,In_1818);
xnor U536 (N_536,In_1711,In_325);
xnor U537 (N_537,In_1700,In_676);
nand U538 (N_538,In_1031,In_2481);
or U539 (N_539,In_2421,In_1323);
xor U540 (N_540,In_1765,In_1969);
and U541 (N_541,In_613,In_2895);
xor U542 (N_542,In_2571,In_249);
nor U543 (N_543,In_947,In_90);
and U544 (N_544,In_1825,In_610);
nor U545 (N_545,In_1994,In_815);
and U546 (N_546,In_1343,In_1875);
or U547 (N_547,In_2505,In_1521);
nand U548 (N_548,In_839,In_2858);
nor U549 (N_549,In_2139,In_51);
and U550 (N_550,In_2269,In_2720);
nor U551 (N_551,In_2582,In_1515);
and U552 (N_552,In_98,In_2212);
nor U553 (N_553,In_2780,In_1732);
nand U554 (N_554,In_841,In_1581);
xor U555 (N_555,In_1881,In_316);
or U556 (N_556,In_2847,In_1130);
nand U557 (N_557,In_569,In_2270);
nor U558 (N_558,In_2037,In_805);
nand U559 (N_559,In_2849,In_65);
nor U560 (N_560,In_64,In_779);
nand U561 (N_561,In_1561,In_2475);
nand U562 (N_562,In_1378,In_534);
xor U563 (N_563,In_87,In_2207);
nor U564 (N_564,In_93,In_821);
nor U565 (N_565,In_1850,In_218);
xor U566 (N_566,In_1061,In_572);
xnor U567 (N_567,In_2236,In_60);
and U568 (N_568,In_1644,In_1151);
nand U569 (N_569,In_1645,In_1293);
nand U570 (N_570,In_2821,In_2178);
xnor U571 (N_571,In_1962,In_479);
and U572 (N_572,In_405,In_932);
nor U573 (N_573,In_2459,In_2431);
and U574 (N_574,In_89,In_1104);
xor U575 (N_575,In_2145,In_2865);
nor U576 (N_576,In_1800,In_1502);
and U577 (N_577,In_1014,In_1535);
or U578 (N_578,In_1647,In_2805);
nand U579 (N_579,In_1044,In_1719);
and U580 (N_580,In_515,In_297);
nor U581 (N_581,In_1804,In_466);
and U582 (N_582,In_661,In_873);
nand U583 (N_583,In_1699,In_2028);
and U584 (N_584,In_1735,In_2769);
nor U585 (N_585,In_2617,In_1235);
nor U586 (N_586,In_1428,In_2965);
nor U587 (N_587,In_1209,In_2867);
nor U588 (N_588,In_1584,In_1432);
and U589 (N_589,In_2169,In_1828);
and U590 (N_590,In_1414,In_1604);
nor U591 (N_591,In_1989,In_955);
and U592 (N_592,In_1658,In_125);
xnor U593 (N_593,In_2328,In_2668);
nor U594 (N_594,In_997,In_961);
xor U595 (N_595,In_920,In_2438);
nor U596 (N_596,In_305,In_657);
xnor U597 (N_597,In_892,In_1478);
and U598 (N_598,In_2234,In_2467);
xnor U599 (N_599,In_612,In_2143);
nand U600 (N_600,In_92,In_96);
nor U601 (N_601,In_1571,In_298);
or U602 (N_602,In_802,In_1550);
xnor U603 (N_603,In_816,In_324);
or U604 (N_604,In_2007,In_286);
or U605 (N_605,In_862,In_1946);
and U606 (N_606,In_1038,In_2148);
or U607 (N_607,In_927,In_1698);
nand U608 (N_608,In_2689,In_81);
and U609 (N_609,In_1889,In_2850);
nand U610 (N_610,In_2711,In_520);
nor U611 (N_611,In_2747,In_1868);
xor U612 (N_612,In_35,In_2205);
or U613 (N_613,In_2777,In_2071);
and U614 (N_614,In_1617,In_1903);
or U615 (N_615,In_827,In_1210);
or U616 (N_616,In_2994,In_2368);
nand U617 (N_617,In_2659,In_2259);
nor U618 (N_618,In_585,In_345);
and U619 (N_619,In_381,In_2155);
nor U620 (N_620,In_2358,In_2835);
or U621 (N_621,In_2260,In_2217);
or U622 (N_622,In_1943,In_134);
xnor U623 (N_623,In_739,In_1168);
xnor U624 (N_624,In_1448,In_2443);
or U625 (N_625,In_1637,In_982);
and U626 (N_626,In_2279,In_2938);
and U627 (N_627,In_2593,In_45);
nand U628 (N_628,In_1019,In_4);
xnor U629 (N_629,In_654,In_1134);
nand U630 (N_630,In_1189,In_255);
or U631 (N_631,In_1608,In_1664);
nor U632 (N_632,In_124,In_1602);
xnor U633 (N_633,In_986,In_482);
and U634 (N_634,In_2833,In_2653);
and U635 (N_635,In_2590,In_819);
nor U636 (N_636,In_2313,In_1523);
or U637 (N_637,In_1941,In_1855);
nor U638 (N_638,In_1459,In_877);
nand U639 (N_639,In_232,In_2819);
and U640 (N_640,In_1784,In_2303);
and U641 (N_641,In_1840,In_2390);
nand U642 (N_642,In_582,In_2730);
or U643 (N_643,In_709,In_940);
nand U644 (N_644,In_242,In_2698);
xnor U645 (N_645,In_2316,In_1681);
nand U646 (N_646,In_1068,In_1522);
xor U647 (N_647,In_2101,In_824);
nor U648 (N_648,In_2550,In_1980);
or U649 (N_649,In_978,In_2723);
and U650 (N_650,In_2758,In_2056);
xor U651 (N_651,In_1030,In_666);
xor U652 (N_652,In_1834,In_695);
and U653 (N_653,In_777,In_238);
nor U654 (N_654,In_2393,In_1465);
nor U655 (N_655,In_2046,In_2463);
xor U656 (N_656,In_1972,In_1353);
nor U657 (N_657,In_2377,In_1965);
xnor U658 (N_658,In_1086,In_1717);
xor U659 (N_659,In_2370,In_2001);
nand U660 (N_660,In_1634,In_1142);
nor U661 (N_661,In_2182,In_682);
and U662 (N_662,In_1137,In_2909);
nor U663 (N_663,In_2,In_1106);
nor U664 (N_664,In_2837,In_378);
or U665 (N_665,In_2520,In_1400);
nor U666 (N_666,In_1622,In_206);
and U667 (N_667,In_1036,In_176);
xnor U668 (N_668,In_1511,In_2531);
xor U669 (N_669,In_2776,In_1111);
nor U670 (N_670,In_1005,In_1080);
xor U671 (N_671,In_1268,In_1507);
or U672 (N_672,In_2267,In_355);
and U673 (N_673,In_2095,In_2014);
xnor U674 (N_674,In_2790,In_552);
and U675 (N_675,In_1563,In_718);
or U676 (N_676,In_2250,In_1805);
nor U677 (N_677,In_1493,In_976);
xnor U678 (N_678,In_1325,In_1555);
and U679 (N_679,In_2119,In_1429);
xnor U680 (N_680,In_1950,In_279);
and U681 (N_681,In_2103,In_692);
and U682 (N_682,In_359,In_2017);
nor U683 (N_683,In_896,In_885);
xnor U684 (N_684,In_2253,In_2323);
and U685 (N_685,In_1961,In_2066);
nor U686 (N_686,In_1474,In_1978);
nand U687 (N_687,In_1215,In_1926);
and U688 (N_688,In_2332,In_2651);
and U689 (N_689,In_1131,In_265);
or U690 (N_690,In_658,In_363);
and U691 (N_691,In_452,In_1673);
xor U692 (N_692,In_2152,In_271);
nand U693 (N_693,In_1393,In_2341);
or U694 (N_694,In_2972,In_2440);
nor U695 (N_695,In_626,In_930);
xnor U696 (N_696,In_2535,In_468);
xor U697 (N_697,In_61,In_2599);
or U698 (N_698,In_1710,In_826);
nand U699 (N_699,In_2948,In_1167);
and U700 (N_700,In_2753,In_411);
or U701 (N_701,In_1983,In_1307);
xor U702 (N_702,In_2638,In_2355);
nor U703 (N_703,In_586,In_1159);
or U704 (N_704,In_75,In_2023);
xor U705 (N_705,In_694,In_1870);
or U706 (N_706,In_2064,In_1225);
nor U707 (N_707,In_2282,In_908);
or U708 (N_708,In_139,In_1275);
and U709 (N_709,In_197,In_2799);
nor U710 (N_710,In_2575,In_413);
nand U711 (N_711,In_1329,In_2016);
nor U712 (N_712,In_2553,In_550);
xor U713 (N_713,In_1867,In_579);
and U714 (N_714,In_1973,In_1178);
nor U715 (N_715,In_655,In_2868);
nor U716 (N_716,In_987,In_36);
and U717 (N_717,In_2228,In_23);
xnor U718 (N_718,In_46,In_2834);
xor U719 (N_719,In_1573,In_477);
nand U720 (N_720,In_1228,In_2569);
and U721 (N_721,In_1541,In_1078);
or U722 (N_722,In_299,In_1156);
xnor U723 (N_723,In_2423,In_2308);
or U724 (N_724,In_1869,In_1356);
or U725 (N_725,In_100,In_1250);
and U726 (N_726,In_1034,In_2971);
and U727 (N_727,In_1615,In_269);
and U728 (N_728,In_180,In_163);
and U729 (N_729,In_2791,In_1000);
nand U730 (N_730,In_2645,In_2731);
nor U731 (N_731,In_1305,In_2059);
nor U732 (N_732,In_2857,In_2786);
xnor U733 (N_733,In_474,In_1282);
xor U734 (N_734,In_618,In_2417);
nand U735 (N_735,In_1362,In_68);
xor U736 (N_736,In_1368,In_1399);
and U737 (N_737,In_2441,In_725);
and U738 (N_738,In_1491,In_77);
xor U739 (N_739,In_1408,In_1457);
and U740 (N_740,In_1812,In_2013);
and U741 (N_741,In_1510,In_1542);
and U742 (N_742,In_797,In_548);
and U743 (N_743,In_1763,In_2098);
and U744 (N_744,In_2500,In_2478);
xor U745 (N_745,In_1102,In_1630);
and U746 (N_746,In_740,In_321);
or U747 (N_747,In_833,In_766);
nor U748 (N_748,In_2673,In_2539);
xnor U749 (N_749,In_2658,In_583);
and U750 (N_750,In_434,In_1162);
nor U751 (N_751,In_2018,In_594);
nor U752 (N_752,In_879,In_2750);
nor U753 (N_753,In_44,In_2842);
nand U754 (N_754,In_1331,In_998);
nand U755 (N_755,In_2871,In_1866);
or U756 (N_756,In_1121,In_2226);
nor U757 (N_757,In_1880,In_2108);
or U758 (N_758,In_1635,In_1165);
nor U759 (N_759,In_221,In_1361);
nor U760 (N_760,In_2998,In_2947);
nor U761 (N_761,In_1028,In_2039);
and U762 (N_762,In_669,In_1513);
xor U763 (N_763,In_2277,In_346);
and U764 (N_764,In_1621,In_1468);
xor U765 (N_765,In_1188,In_227);
nand U766 (N_766,In_2978,In_923);
nor U767 (N_767,In_198,In_1171);
xor U768 (N_768,In_439,In_1814);
nand U769 (N_769,In_446,In_2468);
and U770 (N_770,In_566,In_746);
nor U771 (N_771,In_2633,In_1488);
xor U772 (N_772,In_323,In_1352);
or U773 (N_773,In_1751,In_2783);
xor U774 (N_774,In_851,In_2946);
and U775 (N_775,In_2725,In_2935);
nor U776 (N_776,In_1300,In_2630);
or U777 (N_777,In_1097,In_2032);
xor U778 (N_778,In_801,In_1653);
xor U779 (N_779,In_2975,In_1204);
and U780 (N_780,In_194,In_1063);
nand U781 (N_781,In_1682,In_2605);
nor U782 (N_782,In_2376,In_1879);
nand U783 (N_783,In_253,In_1438);
and U784 (N_784,In_2365,In_2450);
nand U785 (N_785,In_2869,In_2021);
xnor U786 (N_786,In_1674,In_1837);
xor U787 (N_787,In_2993,In_1955);
nor U788 (N_788,In_1556,In_1924);
nand U789 (N_789,In_814,In_2494);
xor U790 (N_790,In_2774,In_1586);
nand U791 (N_791,In_431,In_1678);
xnor U792 (N_792,In_687,In_2068);
xor U793 (N_793,In_488,In_1258);
or U794 (N_794,In_1013,In_2252);
and U795 (N_795,In_1208,In_1027);
or U796 (N_796,In_14,In_1554);
nor U797 (N_797,In_15,In_1285);
nor U798 (N_798,In_2428,In_2186);
nand U799 (N_799,In_2862,In_2523);
nor U800 (N_800,In_2266,In_527);
and U801 (N_801,In_778,In_309);
or U802 (N_802,In_2685,In_968);
nand U803 (N_803,In_1683,In_810);
or U804 (N_804,In_240,In_688);
or U805 (N_805,In_2557,In_1433);
and U806 (N_806,In_2719,In_2684);
nor U807 (N_807,In_2399,In_2383);
or U808 (N_808,In_1666,In_2606);
or U809 (N_809,In_1794,In_2960);
xor U810 (N_810,In_564,In_2885);
nor U811 (N_811,In_208,In_1609);
or U812 (N_812,In_313,In_1538);
and U813 (N_813,In_1160,In_2907);
or U814 (N_814,In_1037,In_1450);
xnor U815 (N_815,In_2041,In_749);
and U816 (N_816,In_629,In_1947);
or U817 (N_817,In_2537,In_2820);
nor U818 (N_818,In_1741,In_2418);
and U819 (N_819,In_1872,In_1788);
xnor U820 (N_820,In_2181,In_1084);
nor U821 (N_821,In_782,In_2681);
nand U822 (N_822,In_2877,In_412);
nand U823 (N_823,In_128,In_373);
nand U824 (N_824,In_2957,In_2696);
nor U825 (N_825,In_2741,In_57);
and U826 (N_826,In_723,In_1018);
xnor U827 (N_827,In_1940,In_990);
nand U828 (N_828,In_2202,In_553);
xor U829 (N_829,In_1348,In_672);
or U830 (N_830,In_370,In_216);
nand U831 (N_831,In_1516,In_532);
nor U832 (N_832,In_2768,In_1864);
nor U833 (N_833,In_48,In_912);
nor U834 (N_834,In_2746,In_2150);
or U835 (N_835,In_379,In_2648);
and U836 (N_836,In_160,In_2940);
or U837 (N_837,In_2838,In_1477);
and U838 (N_838,In_1595,In_2801);
and U839 (N_839,In_288,In_2276);
and U840 (N_840,In_2811,In_2619);
and U841 (N_841,In_261,In_2123);
and U842 (N_842,In_587,In_2740);
and U843 (N_843,In_1149,In_1944);
and U844 (N_844,In_2959,In_122);
nand U845 (N_845,In_117,In_237);
nor U846 (N_846,In_917,In_1544);
and U847 (N_847,In_1723,In_1439);
nor U848 (N_848,In_1109,In_145);
or U849 (N_849,In_83,In_193);
nor U850 (N_850,In_2688,In_2189);
nor U851 (N_851,In_2866,In_1012);
nor U852 (N_852,In_2522,In_2530);
xnor U853 (N_853,In_2538,In_1486);
or U854 (N_854,In_478,In_578);
and U855 (N_855,In_693,In_2245);
xnor U856 (N_856,In_1777,In_2336);
nor U857 (N_857,In_761,In_356);
and U858 (N_858,In_1335,In_1132);
nor U859 (N_859,In_1452,In_510);
xor U860 (N_860,In_931,In_136);
xor U861 (N_861,In_364,In_2744);
xor U862 (N_862,In_1365,In_184);
or U863 (N_863,In_2752,In_1756);
nand U864 (N_864,In_1101,In_1096);
nand U865 (N_865,In_1775,In_1778);
nand U866 (N_866,In_1271,In_2159);
and U867 (N_867,In_1893,In_1154);
nand U868 (N_868,In_1338,In_1786);
nand U869 (N_869,In_1476,In_1407);
and U870 (N_870,In_2086,In_2175);
nand U871 (N_871,In_2872,In_2639);
or U872 (N_872,In_2188,In_1923);
nor U873 (N_873,In_1725,In_1829);
and U874 (N_874,In_2491,In_1655);
nand U875 (N_875,In_1949,In_1714);
and U876 (N_876,In_1281,In_2855);
xor U877 (N_877,In_547,In_69);
and U878 (N_878,In_2581,In_945);
or U879 (N_879,In_1899,In_1313);
nand U880 (N_880,In_2061,In_1269);
and U881 (N_881,In_2465,In_1524);
nand U882 (N_882,In_2813,In_1847);
nand U883 (N_883,In_2385,In_949);
nand U884 (N_884,In_2625,In_1767);
nand U885 (N_885,In_652,In_2348);
and U886 (N_886,In_1092,In_606);
xnor U887 (N_887,In_907,In_94);
xor U888 (N_888,In_2802,In_1360);
nor U889 (N_889,In_179,In_716);
and U890 (N_890,In_764,In_2043);
nand U891 (N_891,In_2131,In_2107);
and U892 (N_892,In_1779,In_2968);
or U893 (N_893,In_2403,In_1806);
xnor U894 (N_894,In_1318,In_1543);
nor U895 (N_895,In_1597,In_1024);
nor U896 (N_896,In_2353,In_1347);
nor U897 (N_897,In_16,In_1755);
nand U898 (N_898,In_848,In_1787);
or U899 (N_899,In_2635,In_274);
or U900 (N_900,In_368,In_660);
nor U901 (N_901,In_1436,In_2009);
nand U902 (N_902,In_1055,In_2171);
or U903 (N_903,In_2949,In_260);
or U904 (N_904,In_1213,In_1411);
and U905 (N_905,In_2812,In_1224);
nand U906 (N_906,In_774,In_500);
or U907 (N_907,In_1547,In_1936);
and U908 (N_908,In_2248,In_1856);
or U909 (N_909,In_1125,In_25);
nor U910 (N_910,In_2680,In_2729);
and U911 (N_911,In_317,In_223);
xnor U912 (N_912,In_187,In_1396);
and U913 (N_913,In_1760,In_604);
xnor U914 (N_914,In_239,In_181);
nand U915 (N_915,In_424,In_944);
nor U916 (N_916,In_2389,In_1442);
nor U917 (N_917,In_2646,In_1616);
or U918 (N_918,In_556,In_388);
and U919 (N_919,In_590,In_1562);
or U920 (N_920,In_2374,In_1636);
or U921 (N_921,In_455,In_376);
nor U922 (N_922,In_329,In_2289);
xnor U923 (N_923,In_2091,In_2810);
or U924 (N_924,In_1500,In_153);
or U925 (N_925,In_2489,In_1816);
nand U926 (N_926,In_1839,In_2916);
xor U927 (N_927,In_1249,In_856);
nand U928 (N_928,In_1540,In_1053);
nor U929 (N_929,In_2327,In_467);
nand U930 (N_930,In_1525,In_2860);
nand U931 (N_931,In_1594,In_2247);
xor U932 (N_932,In_2781,In_341);
or U933 (N_933,In_1991,In_440);
nand U934 (N_934,In_291,In_980);
nor U935 (N_935,In_11,In_637);
nor U936 (N_936,In_2227,In_1232);
xnor U937 (N_937,In_2900,In_1308);
and U938 (N_938,In_2807,In_2244);
or U939 (N_939,In_2287,In_1789);
nand U940 (N_940,In_470,In_1079);
or U941 (N_941,In_1512,In_2297);
nor U942 (N_942,In_715,In_1357);
or U943 (N_943,In_1795,In_2199);
and U944 (N_944,In_22,In_1819);
nand U945 (N_945,In_2933,In_1911);
and U946 (N_946,In_442,In_1694);
or U947 (N_947,In_1712,In_974);
or U948 (N_948,In_1692,In_942);
and U949 (N_949,In_1333,In_149);
or U950 (N_950,In_1835,In_1091);
and U951 (N_951,In_2124,In_1937);
or U952 (N_952,In_903,In_717);
and U953 (N_953,In_866,In_369);
and U954 (N_954,In_301,In_1265);
xnor U955 (N_955,In_2305,In_2587);
xnor U956 (N_956,In_857,In_1153);
or U957 (N_957,In_1150,In_2547);
nand U958 (N_958,In_2278,In_1262);
nor U959 (N_959,In_809,In_1133);
or U960 (N_960,In_1720,In_1627);
nand U961 (N_961,In_418,In_683);
and U962 (N_962,In_967,In_1020);
nand U963 (N_963,In_1484,In_2874);
and U964 (N_964,In_1708,In_1582);
xor U965 (N_965,In_2471,In_789);
xor U966 (N_966,In_1128,In_2765);
nand U967 (N_967,In_1841,In_1273);
or U968 (N_968,In_1580,In_869);
or U969 (N_969,In_853,In_1317);
nor U970 (N_970,In_670,In_2597);
nand U971 (N_971,In_1910,In_784);
nor U972 (N_972,In_2764,In_1785);
and U973 (N_973,In_2485,In_267);
nor U974 (N_974,In_710,In_2649);
nor U975 (N_975,In_1690,In_1216);
and U976 (N_976,In_642,In_78);
or U977 (N_977,In_1015,In_2462);
or U978 (N_978,In_737,In_957);
nor U979 (N_979,In_1774,In_1826);
nand U980 (N_980,In_1843,In_2634);
and U981 (N_981,In_2863,In_1701);
or U982 (N_982,In_157,In_1098);
or U983 (N_983,In_2891,In_2514);
xnor U984 (N_984,In_2552,In_1915);
nor U985 (N_985,In_2800,In_622);
or U986 (N_986,In_1748,In_2822);
nand U987 (N_987,In_2187,In_2906);
xnor U988 (N_988,In_1286,In_1799);
or U989 (N_989,In_2586,In_268);
xor U990 (N_990,In_49,In_1802);
nor U991 (N_991,In_765,In_213);
nand U992 (N_992,In_2656,In_834);
or U993 (N_993,In_1033,In_2853);
xor U994 (N_994,In_2925,In_1280);
or U995 (N_995,In_182,In_2682);
nor U996 (N_996,In_2570,In_1047);
and U997 (N_997,In_1807,In_691);
or U998 (N_998,In_1576,In_1489);
or U999 (N_999,In_832,In_1042);
nor U1000 (N_1000,In_310,In_1590);
xnor U1001 (N_1001,In_2610,In_659);
and U1002 (N_1002,In_2444,In_2905);
or U1003 (N_1003,In_2873,In_2141);
and U1004 (N_1004,In_909,In_2366);
nor U1005 (N_1005,In_150,In_1057);
and U1006 (N_1006,In_2882,In_919);
or U1007 (N_1007,In_775,In_2337);
and U1008 (N_1008,In_1025,In_2657);
xnor U1009 (N_1009,In_867,In_1956);
nor U1010 (N_1010,In_1276,In_395);
and U1011 (N_1011,In_2999,In_2484);
and U1012 (N_1012,In_292,In_189);
xor U1013 (N_1013,In_2986,In_2280);
xnor U1014 (N_1014,In_1620,In_741);
and U1015 (N_1015,In_607,In_521);
xor U1016 (N_1016,In_1687,In_1242);
xnor U1017 (N_1017,In_2713,In_109);
and U1018 (N_1018,In_795,In_233);
nand U1019 (N_1019,In_2401,In_698);
and U1020 (N_1020,In_2166,In_1272);
nand U1021 (N_1021,In_2089,In_1964);
and U1022 (N_1022,In_414,In_1464);
and U1023 (N_1023,In_151,In_2506);
nand U1024 (N_1024,In_1985,In_2613);
or U1025 (N_1025,In_2433,In_280);
xor U1026 (N_1026,In_2137,In_1863);
nand U1027 (N_1027,In_1534,In_2724);
nor U1028 (N_1028,In_170,In_217);
nor U1029 (N_1029,In_1388,In_259);
nand U1030 (N_1030,In_1083,In_144);
or U1031 (N_1031,In_1290,In_1212);
nor U1032 (N_1032,In_1074,In_1730);
or U1033 (N_1033,In_2573,In_1750);
nor U1034 (N_1034,In_1811,In_2395);
nor U1035 (N_1035,In_1251,In_28);
or U1036 (N_1036,In_2839,In_2622);
and U1037 (N_1037,In_1992,In_1064);
xor U1038 (N_1038,In_989,In_898);
nand U1039 (N_1039,In_2598,In_1557);
or U1040 (N_1040,In_858,In_2134);
nand U1041 (N_1041,In_2760,In_1744);
and U1042 (N_1042,In_2815,In_581);
xor U1043 (N_1043,In_2058,In_747);
or U1044 (N_1044,In_2923,In_875);
and U1045 (N_1045,In_701,In_1759);
nand U1046 (N_1046,In_2519,In_1140);
xor U1047 (N_1047,In_79,In_1876);
and U1048 (N_1048,In_1461,In_850);
nand U1049 (N_1049,In_2579,In_2093);
xnor U1050 (N_1050,In_209,In_2737);
and U1051 (N_1051,In_1960,In_1483);
nor U1052 (N_1052,In_2082,In_318);
nand U1053 (N_1053,In_2183,In_650);
xnor U1054 (N_1054,In_471,In_1607);
nand U1055 (N_1055,In_2958,In_540);
and U1056 (N_1056,In_1508,In_2356);
nand U1057 (N_1057,In_2136,In_1136);
nand U1058 (N_1058,In_2734,In_1832);
nor U1059 (N_1059,In_2824,In_2521);
xor U1060 (N_1060,In_1289,In_1624);
nor U1061 (N_1061,In_1551,In_2414);
or U1062 (N_1062,In_2572,In_97);
nand U1063 (N_1063,In_1931,In_505);
xor U1064 (N_1064,In_202,In_863);
nand U1065 (N_1065,In_1334,In_630);
nand U1066 (N_1066,In_295,In_2548);
nor U1067 (N_1067,In_1999,In_849);
nand U1068 (N_1068,In_1404,In_756);
or U1069 (N_1069,In_1238,In_1705);
nor U1070 (N_1070,In_2404,In_2165);
and U1071 (N_1071,In_829,In_2554);
or U1072 (N_1072,In_911,In_2616);
xnor U1073 (N_1073,In_603,In_1316);
nand U1074 (N_1074,In_962,In_855);
xor U1075 (N_1075,In_2704,In_983);
or U1076 (N_1076,In_1509,In_167);
nand U1077 (N_1077,In_496,In_2748);
or U1078 (N_1078,In_668,In_2073);
xor U1079 (N_1079,In_113,In_168);
nand U1080 (N_1080,In_1198,In_2661);
or U1081 (N_1081,In_1848,In_593);
xnor U1082 (N_1082,In_1886,In_2472);
xnor U1083 (N_1083,In_837,In_67);
nor U1084 (N_1084,In_2157,In_2603);
nor U1085 (N_1085,In_2793,In_1234);
and U1086 (N_1086,In_2194,In_2411);
or U1087 (N_1087,In_1430,In_703);
and U1088 (N_1088,In_1533,In_1315);
nand U1089 (N_1089,In_1706,In_2480);
nand U1090 (N_1090,In_426,In_200);
or U1091 (N_1091,In_2261,In_512);
nand U1092 (N_1092,In_1039,In_559);
nand U1093 (N_1093,In_99,In_2663);
or U1094 (N_1094,In_2627,In_1463);
nand U1095 (N_1095,In_2542,In_1842);
nand U1096 (N_1096,In_2997,In_584);
and U1097 (N_1097,In_2026,In_306);
nor U1098 (N_1098,In_1456,In_1183);
xnor U1099 (N_1099,In_854,In_516);
nor U1100 (N_1100,In_1611,In_2386);
or U1101 (N_1101,In_811,In_327);
nor U1102 (N_1102,In_1646,In_159);
xor U1103 (N_1103,In_2876,In_2345);
or U1104 (N_1104,In_728,In_423);
nor U1105 (N_1105,In_404,In_1746);
nor U1106 (N_1106,In_1737,In_1241);
nand U1107 (N_1107,In_649,In_1696);
or U1108 (N_1108,In_26,In_2173);
or U1109 (N_1109,In_742,In_2728);
nor U1110 (N_1110,In_1628,In_2951);
nor U1111 (N_1111,In_1277,In_1901);
or U1112 (N_1112,In_2458,In_398);
and U1113 (N_1113,In_762,In_847);
nand U1114 (N_1114,In_2135,In_2224);
and U1115 (N_1115,In_965,In_570);
nand U1116 (N_1116,In_382,In_360);
nand U1117 (N_1117,In_1900,In_2840);
or U1118 (N_1118,In_501,In_2229);
xor U1119 (N_1119,In_416,In_1394);
nand U1120 (N_1120,In_161,In_2062);
xor U1121 (N_1121,In_2284,In_425);
or U1122 (N_1122,In_2536,In_2448);
nor U1123 (N_1123,In_2410,In_2608);
xnor U1124 (N_1124,In_2271,In_1420);
nor U1125 (N_1125,In_1473,In_549);
xor U1126 (N_1126,In_804,In_1908);
or U1127 (N_1127,In_1240,In_2488);
nor U1128 (N_1128,In_2504,In_1395);
and U1129 (N_1129,In_1884,In_2311);
and U1130 (N_1130,In_2559,In_993);
nor U1131 (N_1131,In_1197,In_2771);
xnor U1132 (N_1132,In_1894,In_864);
nand U1133 (N_1133,In_110,In_817);
nand U1134 (N_1134,In_1495,In_2897);
xor U1135 (N_1135,In_1689,In_1059);
and U1136 (N_1136,In_80,In_2288);
and U1137 (N_1137,In_1749,In_43);
xnor U1138 (N_1138,In_1873,In_1945);
or U1139 (N_1139,In_2246,In_451);
or U1140 (N_1140,In_1752,In_130);
nor U1141 (N_1141,In_971,In_140);
nor U1142 (N_1142,In_1087,In_351);
and U1143 (N_1143,In_2601,In_915);
and U1144 (N_1144,In_1129,In_1470);
nand U1145 (N_1145,In_2990,In_558);
and U1146 (N_1146,In_1743,In_1373);
nand U1147 (N_1147,In_2466,In_711);
or U1148 (N_1148,In_2870,In_2604);
nand U1149 (N_1149,In_523,In_2841);
and U1150 (N_1150,In_2042,In_2922);
nor U1151 (N_1151,In_2113,In_2825);
nor U1152 (N_1152,In_1506,In_2795);
and U1153 (N_1153,In_419,In_546);
and U1154 (N_1154,In_1191,In_2461);
xor U1155 (N_1155,In_358,In_835);
nand U1156 (N_1156,In_953,In_2359);
xnor U1157 (N_1157,In_2665,In_560);
or U1158 (N_1158,In_1126,In_1050);
or U1159 (N_1159,In_2003,In_1233);
nand U1160 (N_1160,In_2510,In_2678);
nor U1161 (N_1161,In_596,In_1721);
nand U1162 (N_1162,In_444,In_1174);
nand U1163 (N_1163,In_893,In_702);
and U1164 (N_1164,In_2373,In_2690);
nor U1165 (N_1165,In_2070,In_2215);
or U1166 (N_1166,In_1218,In_71);
nor U1167 (N_1167,In_2219,In_59);
nand U1168 (N_1168,In_9,In_1364);
and U1169 (N_1169,In_674,In_2996);
or U1170 (N_1170,In_1029,In_2144);
and U1171 (N_1171,In_2412,In_212);
nor U1172 (N_1172,In_486,In_2962);
and U1173 (N_1173,In_195,In_2700);
xnor U1174 (N_1174,In_2984,In_1026);
nor U1175 (N_1175,In_2220,In_2339);
or U1176 (N_1176,In_1990,In_1481);
nand U1177 (N_1177,In_2473,In_320);
and U1178 (N_1178,In_2360,In_1023);
nand U1179 (N_1179,In_2378,In_282);
nand U1180 (N_1180,In_74,In_2293);
nand U1181 (N_1181,In_1589,In_2562);
nand U1182 (N_1182,In_1237,In_1423);
and U1183 (N_1183,In_111,In_1632);
xor U1184 (N_1184,In_667,In_713);
and U1185 (N_1185,In_1643,In_571);
or U1186 (N_1186,In_2755,In_845);
nor U1187 (N_1187,In_2761,In_2272);
and U1188 (N_1188,In_1865,In_2950);
and U1189 (N_1189,In_1798,In_891);
and U1190 (N_1190,In_204,In_322);
nor U1191 (N_1191,In_1367,In_541);
nand U1192 (N_1192,In_2400,In_533);
and U1193 (N_1193,In_890,In_1803);
nand U1194 (N_1194,In_2321,In_2515);
nand U1195 (N_1195,In_8,In_2792);
nand U1196 (N_1196,In_781,In_1919);
nor U1197 (N_1197,In_2901,In_1601);
or U1198 (N_1198,In_2814,In_545);
nor U1199 (N_1199,In_2406,In_2432);
or U1200 (N_1200,In_2174,In_1754);
or U1201 (N_1201,In_347,In_952);
nor U1202 (N_1202,In_2140,In_2992);
and U1203 (N_1203,In_2435,In_1914);
nand U1204 (N_1204,In_1693,In_2031);
xor U1205 (N_1205,In_1426,In_1792);
and U1206 (N_1206,In_1304,In_2676);
nor U1207 (N_1207,In_2956,In_1740);
and U1208 (N_1208,In_1667,In_994);
nand U1209 (N_1209,In_2817,In_616);
or U1210 (N_1210,In_1392,In_1195);
nor U1211 (N_1211,In_1977,In_1349);
nand U1212 (N_1212,In_2927,In_1035);
nand U1213 (N_1213,In_2168,In_2262);
nor U1214 (N_1214,In_2012,In_252);
nor U1215 (N_1215,In_1416,In_754);
xnor U1216 (N_1216,In_1170,In_2679);
nor U1217 (N_1217,In_2179,In_1757);
or U1218 (N_1218,In_2114,In_806);
xnor U1219 (N_1219,In_2775,In_2558);
xor U1220 (N_1220,In_2735,In_354);
nand U1221 (N_1221,In_2120,In_2230);
or U1222 (N_1222,In_960,In_315);
xnor U1223 (N_1223,In_1302,In_2177);
and U1224 (N_1224,In_1612,In_1264);
xnor U1225 (N_1225,In_646,In_1462);
nor U1226 (N_1226,In_1294,In_528);
or U1227 (N_1227,In_1820,In_2883);
or U1228 (N_1228,In_437,In_977);
and U1229 (N_1229,In_2479,In_1164);
nor U1230 (N_1230,In_1862,In_2796);
xor U1231 (N_1231,In_2087,In_1075);
or U1232 (N_1232,In_985,In_422);
or U1233 (N_1233,In_1925,In_1552);
nand U1234 (N_1234,In_2967,In_264);
nor U1235 (N_1235,In_2425,In_1391);
nor U1236 (N_1236,In_2845,In_1747);
or U1237 (N_1237,In_1479,In_1745);
xnor U1238 (N_1238,In_529,In_575);
or U1239 (N_1239,In_812,In_1480);
or U1240 (N_1240,In_1662,In_1201);
nor U1241 (N_1241,In_333,In_1);
nand U1242 (N_1242,In_1190,In_383);
xnor U1243 (N_1243,In_403,In_2221);
xnor U1244 (N_1244,In_1248,In_2034);
nand U1245 (N_1245,In_852,In_644);
nor U1246 (N_1246,In_330,In_201);
or U1247 (N_1247,In_475,In_119);
nor U1248 (N_1248,In_609,In_1200);
nand U1249 (N_1249,In_526,In_1073);
or U1250 (N_1250,In_706,In_2636);
or U1251 (N_1251,In_2477,In_456);
nor U1252 (N_1252,In_653,In_339);
nor U1253 (N_1253,In_1545,In_625);
and U1254 (N_1254,In_601,In_2926);
nand U1255 (N_1255,In_1860,In_2025);
and U1256 (N_1256,In_1022,In_2920);
nand U1257 (N_1257,In_1186,In_966);
nor U1258 (N_1258,In_2887,In_2029);
or U1259 (N_1259,In_2241,In_400);
or U1260 (N_1260,In_1339,In_294);
or U1261 (N_1261,In_1979,In_2233);
nand U1262 (N_1262,In_489,In_1783);
or U1263 (N_1263,In_664,In_2290);
or U1264 (N_1264,In_1728,In_991);
and U1265 (N_1265,In_1537,In_2892);
nor U1266 (N_1266,In_785,In_1496);
xnor U1267 (N_1267,In_1781,In_2899);
nand U1268 (N_1268,In_2263,In_2928);
or U1269 (N_1269,In_1935,In_2111);
xor U1270 (N_1270,In_2487,In_1021);
or U1271 (N_1271,In_933,In_2045);
nor U1272 (N_1272,In_302,In_2836);
xnor U1273 (N_1273,In_362,In_2919);
nor U1274 (N_1274,In_865,In_162);
and U1275 (N_1275,In_107,In_2442);
xor U1276 (N_1276,In_1854,In_2914);
nor U1277 (N_1277,In_2864,In_1088);
nor U1278 (N_1278,In_1182,In_2843);
nor U1279 (N_1279,In_352,In_1909);
and U1280 (N_1280,In_1963,In_588);
and U1281 (N_1281,In_2115,In_430);
nand U1282 (N_1282,In_1406,In_469);
xor U1283 (N_1283,In_1410,In_922);
or U1284 (N_1284,In_1085,In_1824);
and U1285 (N_1285,In_270,In_2469);
nor U1286 (N_1286,In_2848,In_41);
nor U1287 (N_1287,In_366,In_349);
or U1288 (N_1288,In_2198,In_1419);
nand U1289 (N_1289,In_2517,In_1758);
or U1290 (N_1290,In_1320,In_1169);
xor U1291 (N_1291,In_1058,In_407);
or U1292 (N_1292,In_406,In_1441);
xnor U1293 (N_1293,In_925,In_803);
or U1294 (N_1294,In_1453,In_2055);
nand U1295 (N_1295,In_31,In_836);
and U1296 (N_1296,In_2200,In_1497);
and U1297 (N_1297,In_887,In_699);
xor U1298 (N_1298,In_147,In_1056);
xor U1299 (N_1299,In_1321,In_1089);
and U1300 (N_1300,In_1722,In_1363);
or U1301 (N_1301,In_2915,In_2097);
nand U1302 (N_1302,In_677,In_2331);
nor U1303 (N_1303,In_2736,In_2770);
and U1304 (N_1304,In_1046,In_487);
and U1305 (N_1305,In_2963,In_1110);
or U1306 (N_1306,In_1008,In_2693);
and U1307 (N_1307,In_1932,In_2660);
or U1308 (N_1308,In_1671,In_2945);
xnor U1309 (N_1309,In_1654,In_632);
nor U1310 (N_1310,In_928,In_2518);
nand U1311 (N_1311,In_1703,In_2545);
xor U1312 (N_1312,In_152,In_2354);
nand U1313 (N_1313,In_514,In_1501);
or U1314 (N_1314,In_2980,In_598);
and U1315 (N_1315,In_343,In_842);
and U1316 (N_1316,In_2304,In_2880);
or U1317 (N_1317,In_166,In_1095);
nand U1318 (N_1318,In_1466,In_2209);
xnor U1319 (N_1319,In_1793,In_1619);
nand U1320 (N_1320,In_50,In_1427);
or U1321 (N_1321,In_2742,In_1988);
xor U1322 (N_1322,In_1652,In_752);
nand U1323 (N_1323,In_1970,In_462);
nand U1324 (N_1324,In_1727,In_2302);
or U1325 (N_1325,In_1244,In_2273);
or U1326 (N_1326,In_1246,In_1927);
xor U1327 (N_1327,In_1739,In_2859);
nor U1328 (N_1328,In_449,In_338);
nor U1329 (N_1329,In_1797,In_1455);
nor U1330 (N_1330,In_340,In_1006);
nor U1331 (N_1331,In_1768,In_1377);
nand U1332 (N_1332,In_1135,In_2507);
and U1333 (N_1333,In_2902,In_522);
or U1334 (N_1334,In_331,In_645);
or U1335 (N_1335,In_2991,In_1967);
nand U1336 (N_1336,In_1808,In_2307);
xor U1337 (N_1337,In_1306,In_2546);
xnor U1338 (N_1338,In_1858,In_392);
and U1339 (N_1339,In_2585,In_958);
xor U1340 (N_1340,In_2084,In_2717);
nand U1341 (N_1341,In_2372,In_2081);
nand U1342 (N_1342,In_876,In_2264);
xor U1343 (N_1343,In_647,In_2612);
or U1344 (N_1344,In_24,In_1082);
nor U1345 (N_1345,In_1895,In_2060);
nor U1346 (N_1346,In_2594,In_1782);
and U1347 (N_1347,In_1836,In_458);
nor U1348 (N_1348,In_263,In_229);
and U1349 (N_1349,In_2977,In_1629);
nand U1350 (N_1350,In_2929,In_84);
nand U1351 (N_1351,In_1108,In_1344);
or U1352 (N_1352,In_2384,In_70);
or U1353 (N_1353,In_2642,In_2898);
or U1354 (N_1354,In_772,In_1446);
xor U1355 (N_1355,In_2918,In_1379);
and U1356 (N_1356,In_1912,In_2944);
nor U1357 (N_1357,In_460,In_2576);
or U1358 (N_1358,In_1062,In_222);
nand U1359 (N_1359,In_2268,In_2319);
nor U1360 (N_1360,In_493,In_210);
nand U1361 (N_1361,In_1155,In_2125);
nand U1362 (N_1362,In_2455,In_798);
or U1363 (N_1363,In_2396,In_199);
xor U1364 (N_1364,In_2726,In_2932);
or U1365 (N_1365,In_1351,In_2985);
or U1366 (N_1366,In_2816,In_592);
nor U1367 (N_1367,In_138,In_1370);
xor U1368 (N_1368,In_1665,In_1425);
or U1369 (N_1369,In_2158,In_38);
or U1370 (N_1370,In_1309,In_95);
nor U1371 (N_1371,In_391,In_387);
nand U1372 (N_1372,In_861,In_504);
or U1373 (N_1373,In_1916,In_2291);
and U1374 (N_1374,In_2112,In_1413);
and U1375 (N_1375,In_1359,In_2352);
nor U1376 (N_1376,In_2641,In_2185);
or U1377 (N_1377,In_884,In_2047);
xnor U1378 (N_1378,In_1214,In_386);
or U1379 (N_1379,In_791,In_2701);
xor U1380 (N_1380,In_2566,In_2759);
xor U1381 (N_1381,In_1138,In_2878);
nand U1382 (N_1382,In_1297,In_1680);
or U1383 (N_1383,In_769,In_1312);
or U1384 (N_1384,In_2318,In_1314);
xor U1385 (N_1385,In_2351,In_1467);
xor U1386 (N_1386,In_555,In_1518);
xnor U1387 (N_1387,In_1610,In_428);
and U1388 (N_1388,In_1146,In_1336);
nand U1389 (N_1389,In_1172,In_535);
and U1390 (N_1390,In_1938,In_2010);
xnor U1391 (N_1391,In_899,In_2445);
or U1392 (N_1392,In_126,In_1539);
nor U1393 (N_1393,In_2398,In_941);
or U1394 (N_1394,In_1145,In_2943);
xnor U1395 (N_1395,In_926,In_511);
nor U1396 (N_1396,In_1045,In_1724);
xor U1397 (N_1397,In_2476,In_591);
nor U1398 (N_1398,In_91,In_905);
nand U1399 (N_1399,In_375,In_2415);
and U1400 (N_1400,In_1401,In_1187);
and U1401 (N_1401,In_1718,In_272);
xor U1402 (N_1402,In_2889,In_938);
or U1403 (N_1403,In_1298,In_2184);
or U1404 (N_1404,In_1371,In_2640);
nor U1405 (N_1405,In_2973,In_476);
nor U1406 (N_1406,In_432,In_2006);
xnor U1407 (N_1407,In_2910,In_2265);
nand U1408 (N_1408,In_1437,In_1417);
and U1409 (N_1409,In_736,In_758);
and U1410 (N_1410,In_2281,In_393);
and U1411 (N_1411,In_2532,In_503);
nand U1412 (N_1412,In_2100,In_300);
xor U1413 (N_1413,In_1974,In_567);
nand U1414 (N_1414,In_1374,In_2987);
xnor U1415 (N_1415,In_731,In_2583);
xnor U1416 (N_1416,In_1984,In_2088);
or U1417 (N_1417,In_2161,In_2626);
or U1418 (N_1418,In_2190,In_243);
nand U1419 (N_1419,In_2118,In_1223);
or U1420 (N_1420,In_518,In_1263);
xnor U1421 (N_1421,In_1054,In_396);
and U1422 (N_1422,In_174,In_121);
xor U1423 (N_1423,In_2163,In_2828);
xnor U1424 (N_1424,In_1659,In_1736);
xnor U1425 (N_1425,In_441,In_2000);
xnor U1426 (N_1426,In_2394,In_1686);
nor U1427 (N_1427,In_257,In_1221);
and U1428 (N_1428,In_1354,In_2204);
or U1429 (N_1429,In_497,In_2516);
or U1430 (N_1430,In_2192,In_888);
and U1431 (N_1431,In_367,In_2063);
or U1432 (N_1432,In_2295,In_2301);
nor U1433 (N_1433,In_2600,In_825);
xnor U1434 (N_1434,In_1530,In_1390);
nand U1435 (N_1435,In_1090,In_2964);
or U1436 (N_1436,In_447,In_2798);
nor U1437 (N_1437,In_1376,In_1519);
xor U1438 (N_1438,In_2574,In_2296);
or U1439 (N_1439,In_154,In_2367);
xor U1440 (N_1440,In_2694,In_2449);
and U1441 (N_1441,In_1948,In_621);
nand U1442 (N_1442,In_2203,In_2683);
nor U1443 (N_1443,In_1471,In_244);
xor U1444 (N_1444,In_2490,In_1247);
and U1445 (N_1445,In_773,In_513);
nor U1446 (N_1446,In_2988,In_2974);
and U1447 (N_1447,In_2027,In_389);
nor U1448 (N_1448,In_2652,In_241);
xnor U1449 (N_1449,In_1569,In_142);
nand U1450 (N_1450,In_2138,In_2970);
nor U1451 (N_1451,In_2315,In_910);
nand U1452 (N_1452,In_2094,In_2829);
nand U1453 (N_1453,In_1631,In_753);
or U1454 (N_1454,In_2040,In_561);
and U1455 (N_1455,In_1222,In_712);
xnor U1456 (N_1456,In_880,In_573);
nand U1457 (N_1457,In_62,In_40);
or U1458 (N_1458,In_874,In_250);
or U1459 (N_1459,In_1217,In_1049);
or U1460 (N_1460,In_1279,In_1402);
xor U1461 (N_1461,In_1141,In_2584);
and U1462 (N_1462,In_1236,In_707);
or U1463 (N_1463,In_420,In_597);
or U1464 (N_1464,In_2856,In_641);
and U1465 (N_1465,In_1668,In_2808);
nor U1466 (N_1466,In_293,In_101);
xor U1467 (N_1467,In_1639,In_2133);
nand U1468 (N_1468,In_685,In_780);
or U1469 (N_1469,In_950,In_2216);
or U1470 (N_1470,In_2861,In_2540);
nor U1471 (N_1471,In_484,In_1892);
xor U1472 (N_1472,In_1366,In_1670);
nor U1473 (N_1473,In_2621,In_2346);
nand U1474 (N_1474,In_964,In_1405);
and U1475 (N_1475,In_1676,In_443);
xor U1476 (N_1476,In_2526,In_207);
nand U1477 (N_1477,In_2099,In_595);
nand U1478 (N_1478,In_2921,In_118);
nor U1479 (N_1479,In_225,In_2364);
nor U1480 (N_1480,In_1764,In_1179);
nor U1481 (N_1481,In_530,In_679);
xor U1482 (N_1482,In_1173,In_248);
nor U1483 (N_1483,In_1986,In_745);
and U1484 (N_1484,In_1032,In_2809);
xor U1485 (N_1485,In_2637,In_2078);
or U1486 (N_1486,In_1295,In_1469);
xor U1487 (N_1487,In_2416,In_2666);
nor U1488 (N_1488,In_2738,In_1809);
nand U1489 (N_1489,In_1166,In_491);
or U1490 (N_1490,In_2350,In_1375);
xnor U1491 (N_1491,In_2329,In_2908);
xnor U1492 (N_1492,In_633,In_1815);
xnor U1493 (N_1493,In_1350,In_1205);
or U1494 (N_1494,In_1270,In_2492);
nor U1495 (N_1495,In_311,In_972);
or U1496 (N_1496,In_636,In_114);
nand U1497 (N_1497,In_1107,In_639);
or U1498 (N_1498,In_1202,In_472);
or U1499 (N_1499,In_12,In_1939);
xor U1500 (N_1500,In_1757,In_1170);
or U1501 (N_1501,In_331,In_367);
or U1502 (N_1502,In_385,In_2383);
and U1503 (N_1503,In_1933,In_1423);
or U1504 (N_1504,In_2001,In_277);
xor U1505 (N_1505,In_653,In_1094);
xnor U1506 (N_1506,In_747,In_1719);
nand U1507 (N_1507,In_143,In_553);
or U1508 (N_1508,In_1379,In_198);
xor U1509 (N_1509,In_1774,In_2433);
xor U1510 (N_1510,In_747,In_99);
nand U1511 (N_1511,In_2018,In_2176);
nand U1512 (N_1512,In_790,In_130);
or U1513 (N_1513,In_1934,In_978);
nand U1514 (N_1514,In_1805,In_936);
nand U1515 (N_1515,In_958,In_2520);
nand U1516 (N_1516,In_198,In_2760);
nand U1517 (N_1517,In_1859,In_559);
nor U1518 (N_1518,In_1181,In_826);
nand U1519 (N_1519,In_878,In_430);
or U1520 (N_1520,In_2256,In_1720);
nand U1521 (N_1521,In_2646,In_1194);
and U1522 (N_1522,In_1957,In_2735);
nor U1523 (N_1523,In_176,In_2267);
and U1524 (N_1524,In_542,In_2501);
nand U1525 (N_1525,In_2221,In_2630);
xor U1526 (N_1526,In_570,In_47);
nor U1527 (N_1527,In_343,In_1248);
or U1528 (N_1528,In_1162,In_1786);
and U1529 (N_1529,In_236,In_1705);
and U1530 (N_1530,In_1035,In_538);
or U1531 (N_1531,In_1071,In_2302);
or U1532 (N_1532,In_228,In_9);
or U1533 (N_1533,In_1344,In_2977);
xor U1534 (N_1534,In_2461,In_2638);
nand U1535 (N_1535,In_881,In_1488);
and U1536 (N_1536,In_1202,In_942);
and U1537 (N_1537,In_1620,In_2841);
xor U1538 (N_1538,In_2407,In_2302);
nor U1539 (N_1539,In_2387,In_1936);
nor U1540 (N_1540,In_1941,In_1270);
xor U1541 (N_1541,In_2879,In_7);
or U1542 (N_1542,In_1025,In_2132);
nor U1543 (N_1543,In_2782,In_2465);
nor U1544 (N_1544,In_2210,In_2759);
nand U1545 (N_1545,In_1778,In_2643);
and U1546 (N_1546,In_996,In_869);
and U1547 (N_1547,In_982,In_1724);
xor U1548 (N_1548,In_1351,In_2405);
xor U1549 (N_1549,In_338,In_633);
or U1550 (N_1550,In_1501,In_2982);
xnor U1551 (N_1551,In_1587,In_497);
or U1552 (N_1552,In_596,In_1203);
or U1553 (N_1553,In_1639,In_2804);
xnor U1554 (N_1554,In_2510,In_256);
and U1555 (N_1555,In_513,In_2470);
and U1556 (N_1556,In_2092,In_780);
nor U1557 (N_1557,In_2301,In_1834);
xor U1558 (N_1558,In_154,In_2697);
nand U1559 (N_1559,In_1350,In_2722);
nand U1560 (N_1560,In_1734,In_2269);
nor U1561 (N_1561,In_2828,In_81);
xnor U1562 (N_1562,In_2941,In_190);
nor U1563 (N_1563,In_838,In_170);
xnor U1564 (N_1564,In_976,In_2291);
xnor U1565 (N_1565,In_2673,In_2770);
nand U1566 (N_1566,In_1308,In_1810);
nor U1567 (N_1567,In_2065,In_1436);
xor U1568 (N_1568,In_2790,In_1409);
nor U1569 (N_1569,In_1213,In_1963);
and U1570 (N_1570,In_1708,In_2149);
nand U1571 (N_1571,In_2986,In_2912);
and U1572 (N_1572,In_1729,In_1330);
or U1573 (N_1573,In_1659,In_1853);
xor U1574 (N_1574,In_2584,In_2228);
nor U1575 (N_1575,In_1396,In_1527);
or U1576 (N_1576,In_263,In_2309);
or U1577 (N_1577,In_310,In_1354);
or U1578 (N_1578,In_147,In_1055);
and U1579 (N_1579,In_1126,In_2697);
or U1580 (N_1580,In_2956,In_640);
nor U1581 (N_1581,In_1984,In_803);
or U1582 (N_1582,In_565,In_1193);
xnor U1583 (N_1583,In_1975,In_1785);
nand U1584 (N_1584,In_2759,In_1188);
nor U1585 (N_1585,In_358,In_2909);
nor U1586 (N_1586,In_1242,In_1798);
and U1587 (N_1587,In_1399,In_2037);
and U1588 (N_1588,In_26,In_1328);
or U1589 (N_1589,In_2395,In_2901);
nor U1590 (N_1590,In_37,In_795);
nand U1591 (N_1591,In_761,In_318);
nor U1592 (N_1592,In_754,In_299);
or U1593 (N_1593,In_2271,In_1455);
and U1594 (N_1594,In_2374,In_1599);
or U1595 (N_1595,In_2562,In_2535);
nor U1596 (N_1596,In_1315,In_629);
nor U1597 (N_1597,In_736,In_82);
nand U1598 (N_1598,In_1462,In_1854);
xnor U1599 (N_1599,In_760,In_599);
or U1600 (N_1600,In_752,In_1788);
and U1601 (N_1601,In_646,In_1872);
nand U1602 (N_1602,In_1348,In_2858);
nor U1603 (N_1603,In_1391,In_43);
nor U1604 (N_1604,In_1327,In_529);
nand U1605 (N_1605,In_935,In_244);
nor U1606 (N_1606,In_1982,In_851);
xnor U1607 (N_1607,In_2633,In_1708);
or U1608 (N_1608,In_632,In_1675);
nand U1609 (N_1609,In_2943,In_1348);
and U1610 (N_1610,In_2752,In_3);
nor U1611 (N_1611,In_2626,In_1534);
or U1612 (N_1612,In_1863,In_737);
or U1613 (N_1613,In_1132,In_2963);
or U1614 (N_1614,In_1269,In_1720);
nand U1615 (N_1615,In_2898,In_1491);
or U1616 (N_1616,In_2251,In_1132);
and U1617 (N_1617,In_115,In_54);
nand U1618 (N_1618,In_2216,In_899);
or U1619 (N_1619,In_2031,In_2539);
nor U1620 (N_1620,In_1214,In_1556);
and U1621 (N_1621,In_2565,In_1193);
or U1622 (N_1622,In_2653,In_2991);
or U1623 (N_1623,In_564,In_272);
nor U1624 (N_1624,In_258,In_1010);
nand U1625 (N_1625,In_231,In_708);
or U1626 (N_1626,In_1337,In_2335);
nor U1627 (N_1627,In_1850,In_2734);
xor U1628 (N_1628,In_1238,In_188);
or U1629 (N_1629,In_1336,In_1272);
nor U1630 (N_1630,In_1205,In_1553);
and U1631 (N_1631,In_1605,In_1058);
nand U1632 (N_1632,In_487,In_67);
nand U1633 (N_1633,In_2100,In_2291);
nor U1634 (N_1634,In_1197,In_2687);
nand U1635 (N_1635,In_2251,In_2637);
or U1636 (N_1636,In_1538,In_854);
xor U1637 (N_1637,In_2895,In_2274);
or U1638 (N_1638,In_177,In_2715);
nor U1639 (N_1639,In_2555,In_1400);
xnor U1640 (N_1640,In_1377,In_2185);
nand U1641 (N_1641,In_565,In_1409);
nor U1642 (N_1642,In_44,In_965);
or U1643 (N_1643,In_68,In_2826);
and U1644 (N_1644,In_2620,In_158);
xor U1645 (N_1645,In_585,In_2453);
nand U1646 (N_1646,In_2842,In_2042);
nand U1647 (N_1647,In_585,In_697);
nor U1648 (N_1648,In_2328,In_491);
nor U1649 (N_1649,In_1154,In_2755);
or U1650 (N_1650,In_218,In_65);
nor U1651 (N_1651,In_1697,In_708);
nand U1652 (N_1652,In_2248,In_550);
xor U1653 (N_1653,In_716,In_1363);
or U1654 (N_1654,In_1194,In_496);
xnor U1655 (N_1655,In_1150,In_2546);
nand U1656 (N_1656,In_952,In_988);
nor U1657 (N_1657,In_174,In_1621);
xor U1658 (N_1658,In_747,In_736);
or U1659 (N_1659,In_1345,In_2068);
nand U1660 (N_1660,In_795,In_2298);
and U1661 (N_1661,In_2482,In_2819);
nand U1662 (N_1662,In_1099,In_1837);
or U1663 (N_1663,In_840,In_308);
xor U1664 (N_1664,In_1899,In_924);
and U1665 (N_1665,In_1430,In_2111);
nor U1666 (N_1666,In_1400,In_2791);
nand U1667 (N_1667,In_1390,In_875);
xnor U1668 (N_1668,In_2001,In_2487);
or U1669 (N_1669,In_1863,In_911);
or U1670 (N_1670,In_163,In_280);
and U1671 (N_1671,In_911,In_1888);
and U1672 (N_1672,In_1167,In_815);
or U1673 (N_1673,In_216,In_929);
xor U1674 (N_1674,In_213,In_965);
nor U1675 (N_1675,In_2741,In_1957);
nand U1676 (N_1676,In_435,In_162);
nand U1677 (N_1677,In_2919,In_617);
and U1678 (N_1678,In_675,In_1716);
xnor U1679 (N_1679,In_852,In_2205);
nand U1680 (N_1680,In_2054,In_2309);
nor U1681 (N_1681,In_1602,In_1081);
and U1682 (N_1682,In_2596,In_1673);
and U1683 (N_1683,In_1024,In_1283);
nand U1684 (N_1684,In_535,In_1328);
or U1685 (N_1685,In_2012,In_2134);
nand U1686 (N_1686,In_1352,In_1271);
xnor U1687 (N_1687,In_2330,In_794);
and U1688 (N_1688,In_2762,In_1191);
nand U1689 (N_1689,In_793,In_2027);
xnor U1690 (N_1690,In_1518,In_2002);
nor U1691 (N_1691,In_1225,In_26);
and U1692 (N_1692,In_2533,In_847);
and U1693 (N_1693,In_2624,In_2873);
nor U1694 (N_1694,In_462,In_1724);
or U1695 (N_1695,In_1029,In_947);
or U1696 (N_1696,In_2467,In_2570);
and U1697 (N_1697,In_752,In_1064);
nand U1698 (N_1698,In_1006,In_2375);
xnor U1699 (N_1699,In_1628,In_630);
and U1700 (N_1700,In_1534,In_2344);
nor U1701 (N_1701,In_2016,In_2463);
or U1702 (N_1702,In_2119,In_2156);
xnor U1703 (N_1703,In_1306,In_1300);
nand U1704 (N_1704,In_1680,In_395);
xor U1705 (N_1705,In_1393,In_332);
and U1706 (N_1706,In_2851,In_2970);
nand U1707 (N_1707,In_2319,In_2640);
nand U1708 (N_1708,In_1414,In_2681);
nand U1709 (N_1709,In_44,In_2457);
xnor U1710 (N_1710,In_18,In_1973);
nand U1711 (N_1711,In_2572,In_2425);
nand U1712 (N_1712,In_27,In_1176);
and U1713 (N_1713,In_1652,In_70);
xor U1714 (N_1714,In_1474,In_785);
and U1715 (N_1715,In_129,In_1621);
nor U1716 (N_1716,In_2728,In_2771);
or U1717 (N_1717,In_254,In_2111);
and U1718 (N_1718,In_2792,In_2429);
xor U1719 (N_1719,In_2737,In_1240);
and U1720 (N_1720,In_48,In_2203);
and U1721 (N_1721,In_2602,In_2135);
xor U1722 (N_1722,In_2819,In_1380);
nor U1723 (N_1723,In_907,In_2927);
xnor U1724 (N_1724,In_1720,In_265);
or U1725 (N_1725,In_594,In_562);
xor U1726 (N_1726,In_206,In_1331);
xor U1727 (N_1727,In_150,In_2311);
nand U1728 (N_1728,In_1835,In_1148);
nand U1729 (N_1729,In_1581,In_1281);
nand U1730 (N_1730,In_1932,In_2510);
xor U1731 (N_1731,In_2342,In_32);
and U1732 (N_1732,In_2578,In_979);
nor U1733 (N_1733,In_2058,In_1947);
or U1734 (N_1734,In_1926,In_1230);
nand U1735 (N_1735,In_2143,In_91);
nor U1736 (N_1736,In_2089,In_1095);
nand U1737 (N_1737,In_443,In_1914);
or U1738 (N_1738,In_870,In_1168);
nand U1739 (N_1739,In_665,In_935);
nor U1740 (N_1740,In_1631,In_1228);
and U1741 (N_1741,In_11,In_2846);
xnor U1742 (N_1742,In_1431,In_936);
and U1743 (N_1743,In_206,In_2427);
nand U1744 (N_1744,In_1420,In_946);
nor U1745 (N_1745,In_1475,In_2076);
nor U1746 (N_1746,In_2119,In_697);
and U1747 (N_1747,In_2485,In_2529);
or U1748 (N_1748,In_2309,In_1768);
and U1749 (N_1749,In_309,In_2687);
and U1750 (N_1750,In_1085,In_2004);
xnor U1751 (N_1751,In_2361,In_2236);
nand U1752 (N_1752,In_1504,In_163);
nor U1753 (N_1753,In_954,In_1472);
xnor U1754 (N_1754,In_1449,In_1361);
and U1755 (N_1755,In_119,In_782);
and U1756 (N_1756,In_1184,In_2790);
nand U1757 (N_1757,In_621,In_1376);
nor U1758 (N_1758,In_2731,In_1108);
nand U1759 (N_1759,In_1822,In_2253);
nand U1760 (N_1760,In_1037,In_1089);
xor U1761 (N_1761,In_2263,In_2064);
or U1762 (N_1762,In_1226,In_470);
nor U1763 (N_1763,In_2194,In_888);
or U1764 (N_1764,In_2717,In_304);
or U1765 (N_1765,In_110,In_2038);
or U1766 (N_1766,In_1938,In_2795);
xor U1767 (N_1767,In_1673,In_1200);
and U1768 (N_1768,In_2456,In_215);
or U1769 (N_1769,In_1168,In_2808);
nor U1770 (N_1770,In_359,In_1722);
nor U1771 (N_1771,In_1438,In_602);
and U1772 (N_1772,In_729,In_1230);
or U1773 (N_1773,In_1844,In_2918);
xnor U1774 (N_1774,In_2894,In_963);
nor U1775 (N_1775,In_610,In_2577);
and U1776 (N_1776,In_1918,In_286);
and U1777 (N_1777,In_1857,In_961);
nor U1778 (N_1778,In_1678,In_416);
nand U1779 (N_1779,In_62,In_1949);
and U1780 (N_1780,In_1494,In_81);
or U1781 (N_1781,In_589,In_1515);
or U1782 (N_1782,In_836,In_1371);
or U1783 (N_1783,In_2884,In_1151);
xnor U1784 (N_1784,In_1605,In_2305);
nand U1785 (N_1785,In_2894,In_97);
xnor U1786 (N_1786,In_2115,In_2456);
and U1787 (N_1787,In_1903,In_391);
or U1788 (N_1788,In_1537,In_33);
nand U1789 (N_1789,In_964,In_2184);
nor U1790 (N_1790,In_141,In_2677);
and U1791 (N_1791,In_479,In_170);
and U1792 (N_1792,In_2813,In_332);
nor U1793 (N_1793,In_2494,In_2968);
and U1794 (N_1794,In_1133,In_2929);
xnor U1795 (N_1795,In_1716,In_1565);
xor U1796 (N_1796,In_1968,In_561);
and U1797 (N_1797,In_1928,In_1946);
xnor U1798 (N_1798,In_1853,In_2297);
or U1799 (N_1799,In_1037,In_669);
nand U1800 (N_1800,In_2724,In_1700);
nand U1801 (N_1801,In_2682,In_517);
nor U1802 (N_1802,In_634,In_2682);
or U1803 (N_1803,In_2131,In_2385);
or U1804 (N_1804,In_1832,In_1000);
or U1805 (N_1805,In_2617,In_2108);
and U1806 (N_1806,In_342,In_2375);
or U1807 (N_1807,In_427,In_882);
and U1808 (N_1808,In_130,In_1464);
xnor U1809 (N_1809,In_1588,In_937);
nor U1810 (N_1810,In_2041,In_2453);
nand U1811 (N_1811,In_2162,In_1553);
and U1812 (N_1812,In_744,In_2850);
or U1813 (N_1813,In_295,In_2835);
and U1814 (N_1814,In_2592,In_2258);
and U1815 (N_1815,In_1807,In_2827);
nand U1816 (N_1816,In_2931,In_1456);
nor U1817 (N_1817,In_1430,In_2618);
nor U1818 (N_1818,In_251,In_2467);
nand U1819 (N_1819,In_2431,In_1112);
nor U1820 (N_1820,In_1262,In_636);
nor U1821 (N_1821,In_336,In_2018);
or U1822 (N_1822,In_1227,In_101);
nor U1823 (N_1823,In_2231,In_2956);
or U1824 (N_1824,In_2140,In_1322);
or U1825 (N_1825,In_1334,In_1710);
xor U1826 (N_1826,In_2883,In_1466);
xnor U1827 (N_1827,In_1063,In_963);
nor U1828 (N_1828,In_2802,In_504);
nand U1829 (N_1829,In_2311,In_2775);
nor U1830 (N_1830,In_1808,In_475);
nor U1831 (N_1831,In_857,In_21);
xor U1832 (N_1832,In_1129,In_943);
and U1833 (N_1833,In_994,In_2853);
nor U1834 (N_1834,In_1873,In_598);
or U1835 (N_1835,In_2265,In_2881);
nand U1836 (N_1836,In_2565,In_2851);
or U1837 (N_1837,In_1038,In_1070);
or U1838 (N_1838,In_1185,In_2457);
and U1839 (N_1839,In_1847,In_2306);
or U1840 (N_1840,In_1327,In_2160);
xnor U1841 (N_1841,In_312,In_311);
nor U1842 (N_1842,In_989,In_1072);
and U1843 (N_1843,In_1125,In_587);
and U1844 (N_1844,In_1374,In_30);
xor U1845 (N_1845,In_1294,In_2540);
xnor U1846 (N_1846,In_1694,In_2547);
or U1847 (N_1847,In_889,In_239);
nand U1848 (N_1848,In_2307,In_2453);
or U1849 (N_1849,In_1968,In_1117);
and U1850 (N_1850,In_671,In_2196);
or U1851 (N_1851,In_2844,In_335);
nand U1852 (N_1852,In_1168,In_1067);
xnor U1853 (N_1853,In_426,In_567);
and U1854 (N_1854,In_636,In_565);
or U1855 (N_1855,In_2248,In_2279);
nor U1856 (N_1856,In_857,In_11);
nand U1857 (N_1857,In_1464,In_1236);
xnor U1858 (N_1858,In_2387,In_968);
nand U1859 (N_1859,In_1213,In_747);
and U1860 (N_1860,In_1715,In_2057);
and U1861 (N_1861,In_1912,In_316);
or U1862 (N_1862,In_1853,In_1856);
and U1863 (N_1863,In_2139,In_2393);
nand U1864 (N_1864,In_1039,In_1427);
or U1865 (N_1865,In_1193,In_1488);
xnor U1866 (N_1866,In_1752,In_700);
or U1867 (N_1867,In_2993,In_1717);
and U1868 (N_1868,In_2884,In_2660);
nor U1869 (N_1869,In_459,In_754);
nor U1870 (N_1870,In_383,In_1546);
nor U1871 (N_1871,In_2893,In_609);
or U1872 (N_1872,In_2209,In_1148);
and U1873 (N_1873,In_1306,In_829);
and U1874 (N_1874,In_1570,In_2678);
nor U1875 (N_1875,In_2532,In_486);
and U1876 (N_1876,In_2727,In_807);
nor U1877 (N_1877,In_1750,In_1084);
nor U1878 (N_1878,In_1016,In_1401);
and U1879 (N_1879,In_2685,In_1181);
nor U1880 (N_1880,In_762,In_176);
xor U1881 (N_1881,In_1581,In_1090);
and U1882 (N_1882,In_1754,In_2319);
nand U1883 (N_1883,In_564,In_1187);
nand U1884 (N_1884,In_1092,In_1070);
or U1885 (N_1885,In_412,In_481);
and U1886 (N_1886,In_1601,In_1447);
nor U1887 (N_1887,In_1691,In_868);
and U1888 (N_1888,In_416,In_1672);
nand U1889 (N_1889,In_712,In_285);
nand U1890 (N_1890,In_48,In_1082);
nor U1891 (N_1891,In_1728,In_676);
xor U1892 (N_1892,In_692,In_1586);
xnor U1893 (N_1893,In_1370,In_813);
or U1894 (N_1894,In_2828,In_2784);
and U1895 (N_1895,In_2004,In_150);
xnor U1896 (N_1896,In_2025,In_2833);
and U1897 (N_1897,In_1226,In_1578);
nor U1898 (N_1898,In_2607,In_124);
nor U1899 (N_1899,In_487,In_814);
xnor U1900 (N_1900,In_2279,In_2631);
nand U1901 (N_1901,In_1999,In_1529);
nor U1902 (N_1902,In_1296,In_2662);
or U1903 (N_1903,In_2653,In_2477);
nor U1904 (N_1904,In_1564,In_2872);
nor U1905 (N_1905,In_1177,In_2308);
or U1906 (N_1906,In_2806,In_390);
xnor U1907 (N_1907,In_1311,In_759);
and U1908 (N_1908,In_124,In_1345);
or U1909 (N_1909,In_1527,In_1543);
nand U1910 (N_1910,In_276,In_1652);
nand U1911 (N_1911,In_702,In_1852);
nor U1912 (N_1912,In_1326,In_2506);
or U1913 (N_1913,In_34,In_395);
nand U1914 (N_1914,In_1197,In_831);
or U1915 (N_1915,In_2156,In_505);
nor U1916 (N_1916,In_1962,In_2143);
and U1917 (N_1917,In_2546,In_1136);
xnor U1918 (N_1918,In_2916,In_109);
or U1919 (N_1919,In_224,In_242);
xor U1920 (N_1920,In_2408,In_1705);
xor U1921 (N_1921,In_2822,In_667);
xnor U1922 (N_1922,In_1941,In_2708);
nor U1923 (N_1923,In_765,In_908);
nor U1924 (N_1924,In_812,In_2446);
and U1925 (N_1925,In_2306,In_804);
nor U1926 (N_1926,In_1941,In_1728);
or U1927 (N_1927,In_1150,In_1274);
nand U1928 (N_1928,In_1352,In_2926);
nand U1929 (N_1929,In_2494,In_872);
or U1930 (N_1930,In_780,In_1229);
or U1931 (N_1931,In_2654,In_2096);
and U1932 (N_1932,In_1402,In_1419);
nand U1933 (N_1933,In_604,In_1521);
xor U1934 (N_1934,In_832,In_2513);
and U1935 (N_1935,In_1927,In_1252);
and U1936 (N_1936,In_2500,In_59);
nor U1937 (N_1937,In_1457,In_2272);
or U1938 (N_1938,In_347,In_1441);
nand U1939 (N_1939,In_2250,In_1377);
nor U1940 (N_1940,In_2023,In_2292);
nand U1941 (N_1941,In_1926,In_2865);
or U1942 (N_1942,In_2994,In_1527);
nand U1943 (N_1943,In_2678,In_269);
or U1944 (N_1944,In_2240,In_2998);
nand U1945 (N_1945,In_1273,In_2434);
xor U1946 (N_1946,In_2527,In_1129);
or U1947 (N_1947,In_2390,In_2333);
xnor U1948 (N_1948,In_2424,In_1759);
xor U1949 (N_1949,In_1773,In_272);
and U1950 (N_1950,In_52,In_1748);
xor U1951 (N_1951,In_1855,In_1243);
nand U1952 (N_1952,In_1163,In_2182);
nand U1953 (N_1953,In_1957,In_1049);
and U1954 (N_1954,In_838,In_2297);
nand U1955 (N_1955,In_991,In_2339);
nor U1956 (N_1956,In_1125,In_1898);
and U1957 (N_1957,In_204,In_484);
nand U1958 (N_1958,In_2227,In_1810);
or U1959 (N_1959,In_663,In_2320);
nor U1960 (N_1960,In_1858,In_2096);
xor U1961 (N_1961,In_875,In_1400);
or U1962 (N_1962,In_314,In_508);
nor U1963 (N_1963,In_2993,In_1976);
or U1964 (N_1964,In_694,In_1827);
nor U1965 (N_1965,In_2305,In_1545);
nor U1966 (N_1966,In_1016,In_2886);
nor U1967 (N_1967,In_2853,In_2260);
or U1968 (N_1968,In_2509,In_1018);
xnor U1969 (N_1969,In_2932,In_2156);
nor U1970 (N_1970,In_1240,In_363);
nand U1971 (N_1971,In_2407,In_2949);
and U1972 (N_1972,In_2021,In_1923);
and U1973 (N_1973,In_2589,In_2879);
xor U1974 (N_1974,In_2494,In_1992);
and U1975 (N_1975,In_358,In_882);
nand U1976 (N_1976,In_1094,In_2547);
nand U1977 (N_1977,In_594,In_2143);
nor U1978 (N_1978,In_807,In_2407);
nor U1979 (N_1979,In_350,In_165);
xor U1980 (N_1980,In_111,In_232);
xor U1981 (N_1981,In_174,In_1391);
nor U1982 (N_1982,In_1692,In_1015);
nor U1983 (N_1983,In_2983,In_1101);
nor U1984 (N_1984,In_457,In_2155);
and U1985 (N_1985,In_2085,In_2606);
nand U1986 (N_1986,In_1412,In_861);
xor U1987 (N_1987,In_1619,In_2005);
xnor U1988 (N_1988,In_2733,In_1529);
nor U1989 (N_1989,In_980,In_1604);
and U1990 (N_1990,In_227,In_1730);
or U1991 (N_1991,In_192,In_1893);
xnor U1992 (N_1992,In_2561,In_340);
xnor U1993 (N_1993,In_2512,In_1318);
and U1994 (N_1994,In_1397,In_1052);
xnor U1995 (N_1995,In_1135,In_1326);
nor U1996 (N_1996,In_1870,In_1320);
nand U1997 (N_1997,In_1038,In_1253);
nor U1998 (N_1998,In_2165,In_574);
nor U1999 (N_1999,In_469,In_2221);
or U2000 (N_2000,In_388,In_286);
nor U2001 (N_2001,In_2619,In_391);
xnor U2002 (N_2002,In_1044,In_792);
nand U2003 (N_2003,In_2358,In_444);
and U2004 (N_2004,In_2341,In_2903);
and U2005 (N_2005,In_1623,In_1029);
and U2006 (N_2006,In_1961,In_1582);
nand U2007 (N_2007,In_2948,In_584);
nand U2008 (N_2008,In_1423,In_2878);
nand U2009 (N_2009,In_2714,In_1406);
nor U2010 (N_2010,In_376,In_1247);
xnor U2011 (N_2011,In_1139,In_277);
and U2012 (N_2012,In_1057,In_1427);
nor U2013 (N_2013,In_1524,In_2783);
nor U2014 (N_2014,In_2930,In_1375);
xor U2015 (N_2015,In_938,In_1485);
nor U2016 (N_2016,In_476,In_2386);
and U2017 (N_2017,In_2625,In_1332);
nor U2018 (N_2018,In_243,In_2640);
xor U2019 (N_2019,In_1733,In_780);
or U2020 (N_2020,In_1506,In_1955);
nor U2021 (N_2021,In_1560,In_356);
or U2022 (N_2022,In_2999,In_836);
nor U2023 (N_2023,In_2354,In_1781);
xnor U2024 (N_2024,In_274,In_2567);
or U2025 (N_2025,In_63,In_608);
and U2026 (N_2026,In_1021,In_1115);
or U2027 (N_2027,In_1869,In_2463);
and U2028 (N_2028,In_2650,In_1092);
or U2029 (N_2029,In_2766,In_912);
xnor U2030 (N_2030,In_1685,In_1003);
or U2031 (N_2031,In_436,In_2490);
and U2032 (N_2032,In_1139,In_887);
and U2033 (N_2033,In_503,In_2404);
xor U2034 (N_2034,In_1728,In_1483);
or U2035 (N_2035,In_2006,In_2294);
or U2036 (N_2036,In_844,In_2309);
and U2037 (N_2037,In_1116,In_1016);
nor U2038 (N_2038,In_2200,In_2014);
nand U2039 (N_2039,In_2814,In_983);
xor U2040 (N_2040,In_1629,In_472);
nand U2041 (N_2041,In_1306,In_2531);
nor U2042 (N_2042,In_1363,In_1571);
or U2043 (N_2043,In_2486,In_2831);
or U2044 (N_2044,In_497,In_2697);
or U2045 (N_2045,In_1133,In_883);
or U2046 (N_2046,In_1848,In_2352);
nor U2047 (N_2047,In_210,In_2162);
and U2048 (N_2048,In_1307,In_1080);
or U2049 (N_2049,In_2613,In_1677);
xnor U2050 (N_2050,In_1401,In_761);
nor U2051 (N_2051,In_172,In_2655);
nor U2052 (N_2052,In_2863,In_1036);
or U2053 (N_2053,In_2051,In_359);
or U2054 (N_2054,In_1121,In_788);
or U2055 (N_2055,In_821,In_1010);
nand U2056 (N_2056,In_43,In_1373);
or U2057 (N_2057,In_385,In_748);
xnor U2058 (N_2058,In_270,In_1680);
xor U2059 (N_2059,In_2014,In_1570);
xor U2060 (N_2060,In_1608,In_541);
and U2061 (N_2061,In_944,In_2103);
nand U2062 (N_2062,In_2321,In_437);
and U2063 (N_2063,In_2711,In_1919);
nor U2064 (N_2064,In_483,In_2039);
and U2065 (N_2065,In_43,In_2886);
and U2066 (N_2066,In_483,In_826);
or U2067 (N_2067,In_1605,In_1304);
nand U2068 (N_2068,In_2682,In_2445);
xor U2069 (N_2069,In_1437,In_1969);
nand U2070 (N_2070,In_408,In_2925);
xnor U2071 (N_2071,In_964,In_103);
nor U2072 (N_2072,In_601,In_158);
and U2073 (N_2073,In_1578,In_2316);
nor U2074 (N_2074,In_1292,In_2213);
nand U2075 (N_2075,In_2434,In_632);
or U2076 (N_2076,In_759,In_2939);
nand U2077 (N_2077,In_193,In_900);
nor U2078 (N_2078,In_2931,In_1106);
and U2079 (N_2079,In_799,In_1930);
nor U2080 (N_2080,In_97,In_2392);
and U2081 (N_2081,In_306,In_1235);
nor U2082 (N_2082,In_1730,In_655);
or U2083 (N_2083,In_271,In_2135);
and U2084 (N_2084,In_2387,In_1793);
xnor U2085 (N_2085,In_1323,In_1217);
xor U2086 (N_2086,In_1354,In_2669);
nand U2087 (N_2087,In_349,In_2873);
nand U2088 (N_2088,In_2298,In_565);
or U2089 (N_2089,In_2569,In_2502);
nand U2090 (N_2090,In_1649,In_2924);
nand U2091 (N_2091,In_1380,In_484);
and U2092 (N_2092,In_2298,In_777);
nand U2093 (N_2093,In_2432,In_279);
nor U2094 (N_2094,In_706,In_2793);
nand U2095 (N_2095,In_1474,In_2157);
and U2096 (N_2096,In_2897,In_2738);
and U2097 (N_2097,In_361,In_2026);
xnor U2098 (N_2098,In_2438,In_1834);
nor U2099 (N_2099,In_1670,In_1250);
xnor U2100 (N_2100,In_1912,In_133);
or U2101 (N_2101,In_1646,In_1258);
or U2102 (N_2102,In_2246,In_582);
nand U2103 (N_2103,In_1827,In_721);
nor U2104 (N_2104,In_683,In_2059);
nor U2105 (N_2105,In_2854,In_2565);
and U2106 (N_2106,In_429,In_1454);
xor U2107 (N_2107,In_2175,In_2330);
nor U2108 (N_2108,In_1545,In_2683);
and U2109 (N_2109,In_1688,In_1953);
or U2110 (N_2110,In_1513,In_1290);
xnor U2111 (N_2111,In_2673,In_1186);
and U2112 (N_2112,In_2236,In_2326);
and U2113 (N_2113,In_37,In_1297);
xor U2114 (N_2114,In_1144,In_1445);
nor U2115 (N_2115,In_1046,In_2869);
and U2116 (N_2116,In_392,In_759);
xnor U2117 (N_2117,In_2586,In_79);
or U2118 (N_2118,In_1731,In_977);
xnor U2119 (N_2119,In_786,In_1396);
nor U2120 (N_2120,In_1292,In_2053);
nand U2121 (N_2121,In_2743,In_1958);
and U2122 (N_2122,In_111,In_188);
xor U2123 (N_2123,In_1311,In_373);
and U2124 (N_2124,In_225,In_2383);
or U2125 (N_2125,In_2553,In_654);
or U2126 (N_2126,In_1387,In_1193);
nand U2127 (N_2127,In_2279,In_1138);
nand U2128 (N_2128,In_1658,In_1979);
and U2129 (N_2129,In_149,In_975);
and U2130 (N_2130,In_2739,In_878);
or U2131 (N_2131,In_0,In_97);
nand U2132 (N_2132,In_7,In_2781);
and U2133 (N_2133,In_759,In_2911);
nor U2134 (N_2134,In_2193,In_2432);
nor U2135 (N_2135,In_1891,In_2969);
nand U2136 (N_2136,In_500,In_846);
and U2137 (N_2137,In_1664,In_2436);
nand U2138 (N_2138,In_499,In_2250);
nor U2139 (N_2139,In_32,In_1510);
nor U2140 (N_2140,In_2843,In_462);
nor U2141 (N_2141,In_1583,In_2099);
and U2142 (N_2142,In_391,In_2621);
nand U2143 (N_2143,In_1727,In_2848);
and U2144 (N_2144,In_1407,In_1671);
nor U2145 (N_2145,In_2171,In_1007);
or U2146 (N_2146,In_976,In_1230);
xor U2147 (N_2147,In_832,In_2433);
and U2148 (N_2148,In_443,In_2329);
nand U2149 (N_2149,In_2386,In_1344);
nand U2150 (N_2150,In_825,In_2229);
or U2151 (N_2151,In_2208,In_691);
nand U2152 (N_2152,In_1312,In_1975);
nor U2153 (N_2153,In_614,In_1124);
xnor U2154 (N_2154,In_1851,In_593);
nor U2155 (N_2155,In_1330,In_459);
nand U2156 (N_2156,In_695,In_1748);
and U2157 (N_2157,In_312,In_133);
or U2158 (N_2158,In_1808,In_2889);
nor U2159 (N_2159,In_216,In_1656);
nand U2160 (N_2160,In_900,In_1144);
and U2161 (N_2161,In_2115,In_1016);
nand U2162 (N_2162,In_348,In_2221);
and U2163 (N_2163,In_903,In_1977);
and U2164 (N_2164,In_2780,In_2561);
nand U2165 (N_2165,In_2986,In_420);
xnor U2166 (N_2166,In_2173,In_1323);
xor U2167 (N_2167,In_1018,In_54);
or U2168 (N_2168,In_1365,In_2917);
xnor U2169 (N_2169,In_1081,In_1178);
and U2170 (N_2170,In_765,In_1320);
xnor U2171 (N_2171,In_494,In_1317);
nand U2172 (N_2172,In_1753,In_382);
nand U2173 (N_2173,In_1240,In_1045);
or U2174 (N_2174,In_887,In_2682);
nand U2175 (N_2175,In_183,In_2305);
xnor U2176 (N_2176,In_172,In_1692);
and U2177 (N_2177,In_577,In_171);
nor U2178 (N_2178,In_2724,In_1721);
and U2179 (N_2179,In_2017,In_1899);
or U2180 (N_2180,In_1879,In_1767);
and U2181 (N_2181,In_702,In_1734);
xnor U2182 (N_2182,In_1524,In_2662);
or U2183 (N_2183,In_750,In_2493);
and U2184 (N_2184,In_1229,In_319);
or U2185 (N_2185,In_739,In_152);
nor U2186 (N_2186,In_575,In_2251);
nand U2187 (N_2187,In_1693,In_33);
nand U2188 (N_2188,In_405,In_1884);
or U2189 (N_2189,In_2965,In_1385);
nand U2190 (N_2190,In_714,In_2736);
nor U2191 (N_2191,In_1695,In_1488);
and U2192 (N_2192,In_700,In_317);
or U2193 (N_2193,In_2321,In_1943);
nor U2194 (N_2194,In_2939,In_260);
and U2195 (N_2195,In_413,In_377);
xor U2196 (N_2196,In_1389,In_2604);
nand U2197 (N_2197,In_1891,In_539);
or U2198 (N_2198,In_930,In_1717);
or U2199 (N_2199,In_1455,In_2546);
nand U2200 (N_2200,In_2418,In_2434);
xor U2201 (N_2201,In_854,In_1450);
and U2202 (N_2202,In_1127,In_336);
xor U2203 (N_2203,In_942,In_1760);
nor U2204 (N_2204,In_2545,In_2188);
xor U2205 (N_2205,In_753,In_2915);
or U2206 (N_2206,In_1742,In_12);
xor U2207 (N_2207,In_1362,In_1666);
xor U2208 (N_2208,In_569,In_1981);
nor U2209 (N_2209,In_313,In_2201);
xnor U2210 (N_2210,In_1170,In_2971);
xor U2211 (N_2211,In_1791,In_1466);
and U2212 (N_2212,In_1542,In_2489);
or U2213 (N_2213,In_2053,In_2530);
and U2214 (N_2214,In_2183,In_1388);
xnor U2215 (N_2215,In_279,In_2122);
or U2216 (N_2216,In_593,In_2377);
and U2217 (N_2217,In_2386,In_2297);
xnor U2218 (N_2218,In_2669,In_570);
xor U2219 (N_2219,In_2210,In_385);
xor U2220 (N_2220,In_2011,In_1147);
nand U2221 (N_2221,In_2038,In_2135);
nand U2222 (N_2222,In_2497,In_1298);
and U2223 (N_2223,In_2271,In_2021);
nor U2224 (N_2224,In_611,In_906);
and U2225 (N_2225,In_2935,In_1060);
xnor U2226 (N_2226,In_1804,In_853);
nor U2227 (N_2227,In_1444,In_1577);
nand U2228 (N_2228,In_620,In_222);
xnor U2229 (N_2229,In_2129,In_2723);
nor U2230 (N_2230,In_1293,In_1926);
and U2231 (N_2231,In_1461,In_1316);
xor U2232 (N_2232,In_746,In_2162);
nor U2233 (N_2233,In_2194,In_2289);
xnor U2234 (N_2234,In_644,In_1031);
xor U2235 (N_2235,In_1822,In_2370);
or U2236 (N_2236,In_619,In_1428);
nor U2237 (N_2237,In_1479,In_1314);
or U2238 (N_2238,In_1515,In_2003);
nor U2239 (N_2239,In_1177,In_2887);
or U2240 (N_2240,In_2433,In_1766);
nor U2241 (N_2241,In_788,In_2827);
nor U2242 (N_2242,In_2802,In_1473);
nand U2243 (N_2243,In_2254,In_2532);
nand U2244 (N_2244,In_2570,In_2681);
xnor U2245 (N_2245,In_1989,In_2002);
nand U2246 (N_2246,In_2747,In_291);
xor U2247 (N_2247,In_157,In_1049);
nand U2248 (N_2248,In_1558,In_2318);
or U2249 (N_2249,In_905,In_2320);
or U2250 (N_2250,In_1876,In_89);
nand U2251 (N_2251,In_2122,In_1555);
or U2252 (N_2252,In_2084,In_2581);
nand U2253 (N_2253,In_1851,In_2956);
nand U2254 (N_2254,In_2644,In_749);
xnor U2255 (N_2255,In_2604,In_1837);
xor U2256 (N_2256,In_1891,In_839);
nand U2257 (N_2257,In_36,In_1540);
nor U2258 (N_2258,In_1413,In_1009);
or U2259 (N_2259,In_1057,In_425);
nand U2260 (N_2260,In_900,In_2152);
xnor U2261 (N_2261,In_46,In_626);
and U2262 (N_2262,In_2102,In_689);
or U2263 (N_2263,In_388,In_2910);
nand U2264 (N_2264,In_234,In_817);
xor U2265 (N_2265,In_1756,In_342);
or U2266 (N_2266,In_2524,In_776);
xor U2267 (N_2267,In_2895,In_2953);
nand U2268 (N_2268,In_2939,In_2704);
xnor U2269 (N_2269,In_2248,In_78);
xnor U2270 (N_2270,In_1478,In_2493);
nor U2271 (N_2271,In_570,In_1075);
or U2272 (N_2272,In_1978,In_2202);
xnor U2273 (N_2273,In_901,In_91);
nand U2274 (N_2274,In_1890,In_778);
and U2275 (N_2275,In_1804,In_777);
nand U2276 (N_2276,In_1237,In_854);
xor U2277 (N_2277,In_136,In_2456);
nand U2278 (N_2278,In_581,In_2066);
or U2279 (N_2279,In_145,In_951);
and U2280 (N_2280,In_2227,In_2829);
nor U2281 (N_2281,In_292,In_1915);
nor U2282 (N_2282,In_2729,In_1707);
or U2283 (N_2283,In_2245,In_1617);
and U2284 (N_2284,In_2316,In_1400);
xnor U2285 (N_2285,In_1317,In_2519);
or U2286 (N_2286,In_2661,In_1309);
xnor U2287 (N_2287,In_1858,In_1983);
xor U2288 (N_2288,In_2440,In_973);
nand U2289 (N_2289,In_342,In_903);
and U2290 (N_2290,In_874,In_1548);
xor U2291 (N_2291,In_170,In_2422);
xnor U2292 (N_2292,In_1096,In_365);
and U2293 (N_2293,In_1770,In_1386);
xnor U2294 (N_2294,In_1148,In_1397);
and U2295 (N_2295,In_1344,In_2922);
xnor U2296 (N_2296,In_593,In_2370);
nand U2297 (N_2297,In_268,In_1594);
xor U2298 (N_2298,In_2374,In_2492);
and U2299 (N_2299,In_243,In_1937);
nand U2300 (N_2300,In_629,In_1395);
or U2301 (N_2301,In_794,In_2592);
and U2302 (N_2302,In_2637,In_885);
and U2303 (N_2303,In_1902,In_1639);
and U2304 (N_2304,In_2270,In_2156);
nor U2305 (N_2305,In_987,In_2992);
or U2306 (N_2306,In_2563,In_898);
nor U2307 (N_2307,In_1722,In_2684);
and U2308 (N_2308,In_387,In_661);
xnor U2309 (N_2309,In_2663,In_2943);
or U2310 (N_2310,In_1241,In_164);
nor U2311 (N_2311,In_582,In_2698);
nor U2312 (N_2312,In_996,In_514);
nor U2313 (N_2313,In_2382,In_1730);
or U2314 (N_2314,In_2278,In_893);
xnor U2315 (N_2315,In_2515,In_39);
nor U2316 (N_2316,In_909,In_2909);
or U2317 (N_2317,In_2352,In_41);
nand U2318 (N_2318,In_1899,In_369);
or U2319 (N_2319,In_2695,In_1966);
nor U2320 (N_2320,In_1692,In_1673);
nand U2321 (N_2321,In_1870,In_873);
nand U2322 (N_2322,In_1404,In_1293);
and U2323 (N_2323,In_2792,In_56);
xnor U2324 (N_2324,In_2048,In_1166);
nand U2325 (N_2325,In_1284,In_1185);
xor U2326 (N_2326,In_2975,In_1945);
nand U2327 (N_2327,In_1459,In_1029);
or U2328 (N_2328,In_566,In_2164);
and U2329 (N_2329,In_1903,In_754);
or U2330 (N_2330,In_1986,In_63);
nand U2331 (N_2331,In_952,In_2744);
xor U2332 (N_2332,In_2536,In_2169);
nor U2333 (N_2333,In_455,In_1700);
or U2334 (N_2334,In_1747,In_157);
xnor U2335 (N_2335,In_1387,In_1562);
xor U2336 (N_2336,In_1092,In_1687);
and U2337 (N_2337,In_2585,In_1057);
nor U2338 (N_2338,In_1733,In_1379);
xor U2339 (N_2339,In_2409,In_370);
nand U2340 (N_2340,In_2644,In_1928);
nor U2341 (N_2341,In_1088,In_286);
xor U2342 (N_2342,In_2172,In_1081);
nand U2343 (N_2343,In_509,In_2687);
xor U2344 (N_2344,In_1958,In_722);
nand U2345 (N_2345,In_2749,In_2281);
xor U2346 (N_2346,In_1952,In_2565);
or U2347 (N_2347,In_1744,In_1342);
and U2348 (N_2348,In_232,In_1271);
and U2349 (N_2349,In_2896,In_148);
xnor U2350 (N_2350,In_879,In_1276);
nand U2351 (N_2351,In_520,In_1640);
and U2352 (N_2352,In_2571,In_1470);
nand U2353 (N_2353,In_1053,In_2493);
or U2354 (N_2354,In_2882,In_220);
xor U2355 (N_2355,In_424,In_2155);
nand U2356 (N_2356,In_1730,In_1020);
and U2357 (N_2357,In_2960,In_2426);
nand U2358 (N_2358,In_2479,In_2328);
nand U2359 (N_2359,In_2069,In_1199);
and U2360 (N_2360,In_2430,In_2081);
or U2361 (N_2361,In_2991,In_243);
or U2362 (N_2362,In_741,In_2493);
xnor U2363 (N_2363,In_1020,In_1401);
nor U2364 (N_2364,In_2506,In_1640);
nand U2365 (N_2365,In_639,In_2290);
xnor U2366 (N_2366,In_560,In_1124);
or U2367 (N_2367,In_1142,In_1279);
and U2368 (N_2368,In_815,In_2554);
and U2369 (N_2369,In_1946,In_1804);
or U2370 (N_2370,In_2633,In_46);
or U2371 (N_2371,In_2000,In_627);
nor U2372 (N_2372,In_635,In_2599);
and U2373 (N_2373,In_956,In_2025);
nand U2374 (N_2374,In_3,In_675);
and U2375 (N_2375,In_458,In_1073);
and U2376 (N_2376,In_1459,In_1020);
or U2377 (N_2377,In_2008,In_2191);
xor U2378 (N_2378,In_1836,In_1673);
nor U2379 (N_2379,In_2112,In_2534);
xnor U2380 (N_2380,In_1542,In_337);
and U2381 (N_2381,In_2596,In_1349);
and U2382 (N_2382,In_2208,In_1686);
or U2383 (N_2383,In_1510,In_1473);
and U2384 (N_2384,In_113,In_2545);
nor U2385 (N_2385,In_2180,In_2811);
nor U2386 (N_2386,In_2,In_773);
xor U2387 (N_2387,In_2527,In_2529);
nand U2388 (N_2388,In_1387,In_2613);
xnor U2389 (N_2389,In_2701,In_266);
or U2390 (N_2390,In_1471,In_1966);
or U2391 (N_2391,In_1934,In_1504);
nand U2392 (N_2392,In_744,In_1130);
nand U2393 (N_2393,In_1346,In_1633);
and U2394 (N_2394,In_680,In_2944);
or U2395 (N_2395,In_411,In_1449);
nor U2396 (N_2396,In_1908,In_2798);
nand U2397 (N_2397,In_1005,In_1748);
and U2398 (N_2398,In_2311,In_2821);
and U2399 (N_2399,In_1277,In_2976);
xnor U2400 (N_2400,In_1086,In_339);
and U2401 (N_2401,In_628,In_1724);
or U2402 (N_2402,In_1741,In_2437);
nand U2403 (N_2403,In_2323,In_2013);
and U2404 (N_2404,In_753,In_1120);
or U2405 (N_2405,In_1358,In_2159);
xor U2406 (N_2406,In_2564,In_2462);
or U2407 (N_2407,In_2915,In_2606);
xor U2408 (N_2408,In_1818,In_600);
and U2409 (N_2409,In_2213,In_2045);
nor U2410 (N_2410,In_924,In_2312);
nor U2411 (N_2411,In_750,In_2280);
or U2412 (N_2412,In_2446,In_1339);
nor U2413 (N_2413,In_2377,In_2422);
xnor U2414 (N_2414,In_2753,In_2672);
xor U2415 (N_2415,In_1151,In_2091);
xnor U2416 (N_2416,In_1953,In_1910);
or U2417 (N_2417,In_310,In_1249);
nor U2418 (N_2418,In_1411,In_2745);
and U2419 (N_2419,In_1483,In_2797);
and U2420 (N_2420,In_2669,In_119);
nor U2421 (N_2421,In_739,In_2093);
nor U2422 (N_2422,In_1297,In_1825);
and U2423 (N_2423,In_1641,In_2174);
or U2424 (N_2424,In_552,In_303);
nor U2425 (N_2425,In_1653,In_2606);
and U2426 (N_2426,In_2175,In_2323);
nor U2427 (N_2427,In_2047,In_2834);
nand U2428 (N_2428,In_2934,In_1517);
nand U2429 (N_2429,In_2874,In_1281);
nor U2430 (N_2430,In_2145,In_2814);
nor U2431 (N_2431,In_641,In_749);
nand U2432 (N_2432,In_60,In_1187);
xor U2433 (N_2433,In_2939,In_240);
xnor U2434 (N_2434,In_1303,In_2270);
xor U2435 (N_2435,In_1033,In_493);
and U2436 (N_2436,In_1325,In_2940);
nand U2437 (N_2437,In_149,In_468);
nor U2438 (N_2438,In_2568,In_2243);
nor U2439 (N_2439,In_2254,In_2294);
or U2440 (N_2440,In_489,In_1557);
and U2441 (N_2441,In_2979,In_1526);
and U2442 (N_2442,In_2702,In_2960);
and U2443 (N_2443,In_1270,In_1161);
and U2444 (N_2444,In_258,In_1107);
nand U2445 (N_2445,In_467,In_2288);
nand U2446 (N_2446,In_385,In_980);
nor U2447 (N_2447,In_1067,In_2665);
xor U2448 (N_2448,In_2912,In_1094);
nand U2449 (N_2449,In_1952,In_1902);
or U2450 (N_2450,In_2812,In_585);
or U2451 (N_2451,In_175,In_1580);
nand U2452 (N_2452,In_342,In_395);
or U2453 (N_2453,In_67,In_1586);
nand U2454 (N_2454,In_186,In_2234);
xnor U2455 (N_2455,In_1911,In_2561);
xnor U2456 (N_2456,In_2412,In_1932);
xor U2457 (N_2457,In_1322,In_2714);
xnor U2458 (N_2458,In_967,In_387);
xnor U2459 (N_2459,In_454,In_2797);
and U2460 (N_2460,In_2886,In_351);
and U2461 (N_2461,In_1462,In_2040);
nand U2462 (N_2462,In_752,In_2212);
or U2463 (N_2463,In_267,In_2181);
nand U2464 (N_2464,In_2413,In_2537);
nor U2465 (N_2465,In_1991,In_1749);
xor U2466 (N_2466,In_919,In_474);
or U2467 (N_2467,In_2109,In_1174);
nand U2468 (N_2468,In_633,In_1242);
xnor U2469 (N_2469,In_2802,In_2458);
nand U2470 (N_2470,In_2247,In_2171);
xor U2471 (N_2471,In_615,In_2169);
xor U2472 (N_2472,In_356,In_2435);
or U2473 (N_2473,In_2360,In_1122);
and U2474 (N_2474,In_1308,In_2562);
or U2475 (N_2475,In_1249,In_2559);
and U2476 (N_2476,In_584,In_1965);
xnor U2477 (N_2477,In_1336,In_409);
xnor U2478 (N_2478,In_148,In_1337);
nor U2479 (N_2479,In_832,In_2161);
nor U2480 (N_2480,In_1435,In_983);
nand U2481 (N_2481,In_481,In_694);
or U2482 (N_2482,In_906,In_629);
nand U2483 (N_2483,In_1702,In_372);
nand U2484 (N_2484,In_468,In_1269);
and U2485 (N_2485,In_1301,In_352);
nor U2486 (N_2486,In_558,In_459);
xor U2487 (N_2487,In_531,In_275);
xnor U2488 (N_2488,In_864,In_278);
and U2489 (N_2489,In_424,In_897);
nor U2490 (N_2490,In_2546,In_2615);
nand U2491 (N_2491,In_2705,In_1572);
or U2492 (N_2492,In_1675,In_1240);
xnor U2493 (N_2493,In_1498,In_810);
and U2494 (N_2494,In_2909,In_2887);
nor U2495 (N_2495,In_2105,In_2202);
or U2496 (N_2496,In_685,In_1158);
or U2497 (N_2497,In_1046,In_145);
xor U2498 (N_2498,In_2320,In_1953);
xor U2499 (N_2499,In_733,In_262);
or U2500 (N_2500,In_76,In_1201);
nand U2501 (N_2501,In_2607,In_439);
xnor U2502 (N_2502,In_1813,In_2605);
xnor U2503 (N_2503,In_2261,In_2772);
nand U2504 (N_2504,In_2540,In_2561);
xnor U2505 (N_2505,In_1153,In_1904);
xor U2506 (N_2506,In_2731,In_1106);
nand U2507 (N_2507,In_2683,In_1966);
nand U2508 (N_2508,In_512,In_1502);
nand U2509 (N_2509,In_2512,In_2623);
nand U2510 (N_2510,In_2021,In_1943);
or U2511 (N_2511,In_1903,In_1142);
nor U2512 (N_2512,In_84,In_463);
xnor U2513 (N_2513,In_2645,In_321);
or U2514 (N_2514,In_2264,In_1612);
nor U2515 (N_2515,In_2627,In_815);
nor U2516 (N_2516,In_2571,In_2413);
and U2517 (N_2517,In_2675,In_239);
nand U2518 (N_2518,In_1846,In_2529);
xnor U2519 (N_2519,In_2572,In_241);
nand U2520 (N_2520,In_2572,In_199);
nand U2521 (N_2521,In_1547,In_215);
nor U2522 (N_2522,In_1603,In_1235);
or U2523 (N_2523,In_2080,In_1912);
xnor U2524 (N_2524,In_680,In_235);
nor U2525 (N_2525,In_2244,In_961);
or U2526 (N_2526,In_1030,In_2958);
or U2527 (N_2527,In_2464,In_477);
or U2528 (N_2528,In_1449,In_1701);
xnor U2529 (N_2529,In_2836,In_856);
xor U2530 (N_2530,In_2220,In_34);
nor U2531 (N_2531,In_782,In_712);
and U2532 (N_2532,In_1507,In_2795);
nand U2533 (N_2533,In_1833,In_2878);
nand U2534 (N_2534,In_1659,In_1057);
xnor U2535 (N_2535,In_1523,In_2958);
or U2536 (N_2536,In_2468,In_2120);
or U2537 (N_2537,In_841,In_1702);
or U2538 (N_2538,In_1167,In_935);
xor U2539 (N_2539,In_2145,In_2966);
or U2540 (N_2540,In_1631,In_1235);
nor U2541 (N_2541,In_214,In_2131);
or U2542 (N_2542,In_533,In_923);
nor U2543 (N_2543,In_2889,In_779);
nand U2544 (N_2544,In_557,In_583);
nor U2545 (N_2545,In_981,In_1024);
nand U2546 (N_2546,In_2078,In_113);
xnor U2547 (N_2547,In_2726,In_1855);
or U2548 (N_2548,In_643,In_2607);
nand U2549 (N_2549,In_2288,In_2245);
nor U2550 (N_2550,In_1805,In_1626);
xnor U2551 (N_2551,In_2953,In_224);
nor U2552 (N_2552,In_643,In_493);
or U2553 (N_2553,In_2475,In_2969);
and U2554 (N_2554,In_2146,In_1976);
nand U2555 (N_2555,In_478,In_2733);
nor U2556 (N_2556,In_2374,In_2464);
nor U2557 (N_2557,In_2364,In_374);
nand U2558 (N_2558,In_2236,In_1277);
nand U2559 (N_2559,In_2026,In_1162);
or U2560 (N_2560,In_2769,In_2191);
and U2561 (N_2561,In_1569,In_2128);
and U2562 (N_2562,In_2338,In_2842);
or U2563 (N_2563,In_1376,In_1703);
and U2564 (N_2564,In_826,In_1996);
nor U2565 (N_2565,In_2355,In_2232);
nor U2566 (N_2566,In_594,In_2684);
xor U2567 (N_2567,In_489,In_2785);
and U2568 (N_2568,In_1539,In_1251);
nand U2569 (N_2569,In_2644,In_2185);
and U2570 (N_2570,In_2615,In_1144);
or U2571 (N_2571,In_231,In_1451);
nand U2572 (N_2572,In_2190,In_656);
or U2573 (N_2573,In_2069,In_28);
and U2574 (N_2574,In_1561,In_2580);
xor U2575 (N_2575,In_502,In_2287);
nand U2576 (N_2576,In_1004,In_2472);
or U2577 (N_2577,In_2780,In_416);
and U2578 (N_2578,In_1262,In_175);
nand U2579 (N_2579,In_37,In_2893);
xor U2580 (N_2580,In_1856,In_2153);
nor U2581 (N_2581,In_2788,In_2902);
xnor U2582 (N_2582,In_1049,In_731);
nor U2583 (N_2583,In_2709,In_361);
nor U2584 (N_2584,In_2217,In_1918);
xor U2585 (N_2585,In_2215,In_626);
nand U2586 (N_2586,In_1099,In_909);
or U2587 (N_2587,In_776,In_848);
or U2588 (N_2588,In_2282,In_1636);
and U2589 (N_2589,In_2276,In_644);
nand U2590 (N_2590,In_2163,In_1983);
xor U2591 (N_2591,In_920,In_1868);
nand U2592 (N_2592,In_2646,In_1590);
nand U2593 (N_2593,In_2320,In_90);
nor U2594 (N_2594,In_1108,In_306);
and U2595 (N_2595,In_2414,In_678);
nand U2596 (N_2596,In_2653,In_734);
nand U2597 (N_2597,In_2154,In_462);
xnor U2598 (N_2598,In_2692,In_2512);
xnor U2599 (N_2599,In_2145,In_1949);
xnor U2600 (N_2600,In_924,In_1339);
or U2601 (N_2601,In_759,In_2594);
nor U2602 (N_2602,In_1342,In_2057);
nor U2603 (N_2603,In_1303,In_795);
xnor U2604 (N_2604,In_2866,In_459);
nor U2605 (N_2605,In_2844,In_2463);
or U2606 (N_2606,In_949,In_312);
nand U2607 (N_2607,In_2108,In_2502);
xor U2608 (N_2608,In_488,In_1378);
or U2609 (N_2609,In_2816,In_2191);
or U2610 (N_2610,In_217,In_2391);
nand U2611 (N_2611,In_2518,In_1296);
nand U2612 (N_2612,In_2513,In_1450);
nor U2613 (N_2613,In_318,In_2088);
xnor U2614 (N_2614,In_876,In_1007);
xor U2615 (N_2615,In_2438,In_1195);
and U2616 (N_2616,In_2315,In_196);
xnor U2617 (N_2617,In_1618,In_668);
and U2618 (N_2618,In_2949,In_2074);
nand U2619 (N_2619,In_1867,In_1564);
or U2620 (N_2620,In_1926,In_2361);
nor U2621 (N_2621,In_2987,In_1568);
nand U2622 (N_2622,In_1358,In_1597);
nand U2623 (N_2623,In_2224,In_639);
nor U2624 (N_2624,In_1350,In_1256);
nor U2625 (N_2625,In_2419,In_1483);
and U2626 (N_2626,In_716,In_1692);
and U2627 (N_2627,In_238,In_667);
or U2628 (N_2628,In_93,In_1934);
xnor U2629 (N_2629,In_1835,In_2591);
or U2630 (N_2630,In_1793,In_1261);
or U2631 (N_2631,In_68,In_1004);
nor U2632 (N_2632,In_126,In_2453);
nand U2633 (N_2633,In_2830,In_2429);
or U2634 (N_2634,In_352,In_1660);
nor U2635 (N_2635,In_70,In_838);
nor U2636 (N_2636,In_2452,In_597);
and U2637 (N_2637,In_2177,In_52);
xnor U2638 (N_2638,In_202,In_928);
and U2639 (N_2639,In_1116,In_743);
and U2640 (N_2640,In_324,In_1152);
nand U2641 (N_2641,In_1673,In_134);
nand U2642 (N_2642,In_271,In_826);
nand U2643 (N_2643,In_2418,In_2619);
xnor U2644 (N_2644,In_1479,In_641);
xnor U2645 (N_2645,In_1996,In_4);
nor U2646 (N_2646,In_2826,In_71);
xnor U2647 (N_2647,In_2725,In_1383);
or U2648 (N_2648,In_337,In_2301);
xor U2649 (N_2649,In_512,In_2644);
or U2650 (N_2650,In_1758,In_1854);
or U2651 (N_2651,In_1173,In_368);
xnor U2652 (N_2652,In_1444,In_856);
xor U2653 (N_2653,In_902,In_388);
and U2654 (N_2654,In_902,In_250);
nor U2655 (N_2655,In_1475,In_2483);
and U2656 (N_2656,In_1141,In_1468);
or U2657 (N_2657,In_2837,In_597);
or U2658 (N_2658,In_1148,In_828);
nand U2659 (N_2659,In_2142,In_636);
nor U2660 (N_2660,In_300,In_169);
nor U2661 (N_2661,In_870,In_2437);
and U2662 (N_2662,In_299,In_2539);
nor U2663 (N_2663,In_425,In_85);
and U2664 (N_2664,In_2870,In_102);
or U2665 (N_2665,In_2667,In_2199);
xnor U2666 (N_2666,In_848,In_2500);
or U2667 (N_2667,In_2740,In_2544);
and U2668 (N_2668,In_1349,In_2330);
xor U2669 (N_2669,In_1077,In_43);
nand U2670 (N_2670,In_2799,In_1643);
nand U2671 (N_2671,In_2447,In_2795);
nor U2672 (N_2672,In_1864,In_2766);
nor U2673 (N_2673,In_2708,In_2994);
nor U2674 (N_2674,In_1168,In_67);
xor U2675 (N_2675,In_1141,In_2535);
xor U2676 (N_2676,In_1830,In_2612);
or U2677 (N_2677,In_361,In_569);
and U2678 (N_2678,In_2309,In_2167);
nand U2679 (N_2679,In_1899,In_1617);
or U2680 (N_2680,In_1580,In_423);
xnor U2681 (N_2681,In_940,In_2438);
or U2682 (N_2682,In_2882,In_2993);
and U2683 (N_2683,In_203,In_2529);
nor U2684 (N_2684,In_1495,In_990);
xnor U2685 (N_2685,In_2488,In_1812);
or U2686 (N_2686,In_988,In_2291);
and U2687 (N_2687,In_1730,In_568);
nor U2688 (N_2688,In_2938,In_2400);
xor U2689 (N_2689,In_1278,In_2489);
or U2690 (N_2690,In_2659,In_625);
xnor U2691 (N_2691,In_2545,In_317);
nor U2692 (N_2692,In_81,In_2623);
or U2693 (N_2693,In_2166,In_1681);
or U2694 (N_2694,In_1697,In_422);
or U2695 (N_2695,In_606,In_396);
and U2696 (N_2696,In_212,In_2192);
nor U2697 (N_2697,In_2202,In_1846);
and U2698 (N_2698,In_1676,In_782);
or U2699 (N_2699,In_1389,In_1550);
and U2700 (N_2700,In_2441,In_57);
and U2701 (N_2701,In_99,In_790);
nor U2702 (N_2702,In_328,In_942);
or U2703 (N_2703,In_2519,In_2025);
or U2704 (N_2704,In_2196,In_2926);
xor U2705 (N_2705,In_1848,In_1405);
and U2706 (N_2706,In_1524,In_2018);
or U2707 (N_2707,In_1981,In_791);
nand U2708 (N_2708,In_2295,In_826);
nand U2709 (N_2709,In_1015,In_2208);
and U2710 (N_2710,In_1735,In_725);
and U2711 (N_2711,In_173,In_1562);
nor U2712 (N_2712,In_2986,In_1362);
nand U2713 (N_2713,In_535,In_1949);
nor U2714 (N_2714,In_1993,In_2214);
and U2715 (N_2715,In_2709,In_2383);
and U2716 (N_2716,In_810,In_2260);
nand U2717 (N_2717,In_1276,In_1469);
nand U2718 (N_2718,In_2759,In_945);
xnor U2719 (N_2719,In_2020,In_1856);
nand U2720 (N_2720,In_2802,In_1288);
and U2721 (N_2721,In_686,In_1496);
xnor U2722 (N_2722,In_1070,In_2082);
nand U2723 (N_2723,In_1239,In_2017);
or U2724 (N_2724,In_1467,In_1711);
nor U2725 (N_2725,In_1011,In_1842);
xor U2726 (N_2726,In_1564,In_276);
or U2727 (N_2727,In_2236,In_2823);
or U2728 (N_2728,In_767,In_1270);
and U2729 (N_2729,In_874,In_614);
xor U2730 (N_2730,In_2825,In_2231);
nor U2731 (N_2731,In_822,In_1617);
nand U2732 (N_2732,In_917,In_532);
nor U2733 (N_2733,In_1651,In_2735);
and U2734 (N_2734,In_1510,In_1639);
nand U2735 (N_2735,In_313,In_508);
and U2736 (N_2736,In_32,In_1926);
nand U2737 (N_2737,In_1863,In_2042);
xnor U2738 (N_2738,In_1905,In_1028);
xor U2739 (N_2739,In_911,In_1277);
nand U2740 (N_2740,In_333,In_2983);
and U2741 (N_2741,In_2703,In_2095);
and U2742 (N_2742,In_751,In_1191);
xor U2743 (N_2743,In_2299,In_339);
and U2744 (N_2744,In_852,In_144);
nand U2745 (N_2745,In_2758,In_1590);
nand U2746 (N_2746,In_1633,In_440);
nand U2747 (N_2747,In_953,In_2140);
xnor U2748 (N_2748,In_2226,In_1922);
nor U2749 (N_2749,In_638,In_968);
or U2750 (N_2750,In_575,In_1723);
and U2751 (N_2751,In_1856,In_1113);
xnor U2752 (N_2752,In_1030,In_2026);
xnor U2753 (N_2753,In_2406,In_1399);
and U2754 (N_2754,In_1753,In_2875);
or U2755 (N_2755,In_425,In_1407);
xnor U2756 (N_2756,In_2004,In_2946);
xor U2757 (N_2757,In_1252,In_1834);
or U2758 (N_2758,In_623,In_1330);
and U2759 (N_2759,In_799,In_1158);
nand U2760 (N_2760,In_2607,In_2559);
nand U2761 (N_2761,In_1465,In_103);
nand U2762 (N_2762,In_504,In_1384);
nor U2763 (N_2763,In_1983,In_2496);
xor U2764 (N_2764,In_573,In_898);
and U2765 (N_2765,In_1280,In_2631);
or U2766 (N_2766,In_2854,In_2974);
nand U2767 (N_2767,In_188,In_2247);
or U2768 (N_2768,In_978,In_1804);
and U2769 (N_2769,In_1333,In_250);
and U2770 (N_2770,In_1474,In_2886);
and U2771 (N_2771,In_519,In_1527);
and U2772 (N_2772,In_381,In_812);
xor U2773 (N_2773,In_537,In_1063);
or U2774 (N_2774,In_1578,In_2027);
and U2775 (N_2775,In_1443,In_166);
xor U2776 (N_2776,In_133,In_2338);
or U2777 (N_2777,In_365,In_2647);
nor U2778 (N_2778,In_2889,In_2570);
and U2779 (N_2779,In_2644,In_848);
xnor U2780 (N_2780,In_278,In_279);
nor U2781 (N_2781,In_898,In_151);
or U2782 (N_2782,In_1666,In_2686);
and U2783 (N_2783,In_256,In_444);
and U2784 (N_2784,In_2278,In_2165);
xnor U2785 (N_2785,In_2937,In_1346);
nand U2786 (N_2786,In_896,In_54);
xor U2787 (N_2787,In_117,In_460);
nand U2788 (N_2788,In_578,In_2486);
and U2789 (N_2789,In_1811,In_2556);
xnor U2790 (N_2790,In_2789,In_699);
nor U2791 (N_2791,In_2298,In_1849);
nand U2792 (N_2792,In_700,In_2623);
nand U2793 (N_2793,In_354,In_1075);
or U2794 (N_2794,In_402,In_1198);
nor U2795 (N_2795,In_2490,In_2771);
nand U2796 (N_2796,In_2704,In_1142);
and U2797 (N_2797,In_2725,In_236);
and U2798 (N_2798,In_2952,In_1638);
nand U2799 (N_2799,In_443,In_2311);
and U2800 (N_2800,In_163,In_2467);
and U2801 (N_2801,In_2888,In_2301);
and U2802 (N_2802,In_1043,In_1818);
nor U2803 (N_2803,In_168,In_1785);
or U2804 (N_2804,In_520,In_2816);
nor U2805 (N_2805,In_1247,In_472);
nor U2806 (N_2806,In_1605,In_820);
xor U2807 (N_2807,In_2751,In_628);
nor U2808 (N_2808,In_975,In_1783);
nand U2809 (N_2809,In_939,In_2321);
nor U2810 (N_2810,In_510,In_2520);
nand U2811 (N_2811,In_1514,In_1336);
xor U2812 (N_2812,In_2395,In_2830);
xor U2813 (N_2813,In_1767,In_512);
nand U2814 (N_2814,In_2770,In_181);
nand U2815 (N_2815,In_2945,In_2380);
or U2816 (N_2816,In_2382,In_549);
xnor U2817 (N_2817,In_1535,In_1735);
nand U2818 (N_2818,In_1012,In_2561);
nand U2819 (N_2819,In_37,In_2892);
xor U2820 (N_2820,In_368,In_2301);
xor U2821 (N_2821,In_484,In_2087);
or U2822 (N_2822,In_1957,In_1211);
nor U2823 (N_2823,In_1440,In_1025);
nand U2824 (N_2824,In_2402,In_1925);
xnor U2825 (N_2825,In_1339,In_506);
and U2826 (N_2826,In_2563,In_2203);
nand U2827 (N_2827,In_2052,In_487);
nand U2828 (N_2828,In_1112,In_456);
or U2829 (N_2829,In_2377,In_2969);
or U2830 (N_2830,In_702,In_1184);
and U2831 (N_2831,In_2503,In_593);
nand U2832 (N_2832,In_2222,In_2681);
or U2833 (N_2833,In_2181,In_376);
nand U2834 (N_2834,In_2983,In_763);
or U2835 (N_2835,In_783,In_1253);
and U2836 (N_2836,In_101,In_2748);
xnor U2837 (N_2837,In_1064,In_2222);
xor U2838 (N_2838,In_836,In_1430);
and U2839 (N_2839,In_2330,In_788);
and U2840 (N_2840,In_2023,In_1420);
nor U2841 (N_2841,In_2648,In_905);
and U2842 (N_2842,In_1854,In_2410);
nor U2843 (N_2843,In_2215,In_89);
xor U2844 (N_2844,In_2849,In_2176);
or U2845 (N_2845,In_2081,In_2802);
and U2846 (N_2846,In_2966,In_1651);
or U2847 (N_2847,In_450,In_2160);
and U2848 (N_2848,In_2170,In_2164);
or U2849 (N_2849,In_1169,In_1418);
xnor U2850 (N_2850,In_2989,In_2794);
or U2851 (N_2851,In_625,In_1104);
nand U2852 (N_2852,In_501,In_752);
or U2853 (N_2853,In_1592,In_1826);
and U2854 (N_2854,In_1688,In_2931);
nand U2855 (N_2855,In_1705,In_869);
or U2856 (N_2856,In_2223,In_1147);
xnor U2857 (N_2857,In_919,In_2962);
and U2858 (N_2858,In_730,In_2356);
and U2859 (N_2859,In_1590,In_2793);
xnor U2860 (N_2860,In_2167,In_1498);
and U2861 (N_2861,In_1444,In_2509);
xnor U2862 (N_2862,In_25,In_2326);
xor U2863 (N_2863,In_816,In_1285);
nor U2864 (N_2864,In_434,In_2645);
nor U2865 (N_2865,In_2381,In_1111);
xnor U2866 (N_2866,In_2612,In_1656);
or U2867 (N_2867,In_2928,In_926);
xor U2868 (N_2868,In_775,In_1859);
and U2869 (N_2869,In_1690,In_913);
nand U2870 (N_2870,In_228,In_2136);
and U2871 (N_2871,In_2821,In_2087);
or U2872 (N_2872,In_2662,In_95);
xnor U2873 (N_2873,In_889,In_774);
and U2874 (N_2874,In_310,In_561);
nor U2875 (N_2875,In_106,In_1601);
nor U2876 (N_2876,In_366,In_1238);
nor U2877 (N_2877,In_228,In_592);
nor U2878 (N_2878,In_1125,In_2133);
or U2879 (N_2879,In_1642,In_1240);
or U2880 (N_2880,In_241,In_1304);
and U2881 (N_2881,In_1423,In_796);
nand U2882 (N_2882,In_2881,In_1264);
nor U2883 (N_2883,In_424,In_1467);
nand U2884 (N_2884,In_1864,In_2998);
nand U2885 (N_2885,In_2392,In_2017);
or U2886 (N_2886,In_1906,In_2898);
or U2887 (N_2887,In_2717,In_226);
xor U2888 (N_2888,In_1619,In_1789);
and U2889 (N_2889,In_2842,In_361);
or U2890 (N_2890,In_530,In_2041);
xnor U2891 (N_2891,In_176,In_397);
xor U2892 (N_2892,In_612,In_2184);
nand U2893 (N_2893,In_2874,In_358);
or U2894 (N_2894,In_1949,In_1469);
nor U2895 (N_2895,In_539,In_1339);
xnor U2896 (N_2896,In_1228,In_1853);
or U2897 (N_2897,In_1272,In_39);
xor U2898 (N_2898,In_386,In_2340);
xnor U2899 (N_2899,In_2752,In_1137);
xnor U2900 (N_2900,In_748,In_260);
nand U2901 (N_2901,In_270,In_1824);
nand U2902 (N_2902,In_1097,In_571);
or U2903 (N_2903,In_1994,In_1570);
xnor U2904 (N_2904,In_739,In_2979);
or U2905 (N_2905,In_767,In_414);
nand U2906 (N_2906,In_2905,In_225);
nor U2907 (N_2907,In_1793,In_868);
nand U2908 (N_2908,In_2289,In_2290);
xor U2909 (N_2909,In_2017,In_2196);
or U2910 (N_2910,In_2178,In_1427);
and U2911 (N_2911,In_2518,In_167);
nor U2912 (N_2912,In_1180,In_2687);
or U2913 (N_2913,In_1420,In_2882);
xnor U2914 (N_2914,In_1097,In_1360);
nand U2915 (N_2915,In_1802,In_1439);
or U2916 (N_2916,In_755,In_1665);
xnor U2917 (N_2917,In_681,In_1190);
nand U2918 (N_2918,In_2729,In_2184);
or U2919 (N_2919,In_281,In_1036);
nand U2920 (N_2920,In_2045,In_1971);
xnor U2921 (N_2921,In_854,In_871);
nand U2922 (N_2922,In_239,In_899);
and U2923 (N_2923,In_2232,In_1315);
xnor U2924 (N_2924,In_1753,In_1723);
nand U2925 (N_2925,In_1057,In_665);
nor U2926 (N_2926,In_495,In_2742);
xor U2927 (N_2927,In_2969,In_2804);
nor U2928 (N_2928,In_2695,In_596);
or U2929 (N_2929,In_1525,In_1661);
or U2930 (N_2930,In_1528,In_304);
and U2931 (N_2931,In_1164,In_117);
nand U2932 (N_2932,In_2885,In_1278);
nand U2933 (N_2933,In_2014,In_1565);
nand U2934 (N_2934,In_1066,In_2153);
nand U2935 (N_2935,In_40,In_1498);
xnor U2936 (N_2936,In_1917,In_2068);
or U2937 (N_2937,In_375,In_66);
nor U2938 (N_2938,In_2199,In_563);
and U2939 (N_2939,In_1152,In_200);
xor U2940 (N_2940,In_913,In_410);
xor U2941 (N_2941,In_2580,In_325);
nand U2942 (N_2942,In_1170,In_2830);
xor U2943 (N_2943,In_1422,In_130);
nor U2944 (N_2944,In_1915,In_1501);
or U2945 (N_2945,In_1044,In_841);
nor U2946 (N_2946,In_2962,In_24);
and U2947 (N_2947,In_1118,In_1329);
and U2948 (N_2948,In_2358,In_2659);
xor U2949 (N_2949,In_1233,In_2173);
and U2950 (N_2950,In_876,In_2062);
or U2951 (N_2951,In_2220,In_1639);
nand U2952 (N_2952,In_866,In_675);
and U2953 (N_2953,In_2366,In_709);
and U2954 (N_2954,In_686,In_1090);
and U2955 (N_2955,In_2941,In_647);
xor U2956 (N_2956,In_45,In_1795);
and U2957 (N_2957,In_918,In_1707);
nor U2958 (N_2958,In_1488,In_92);
xor U2959 (N_2959,In_1785,In_1254);
xnor U2960 (N_2960,In_1881,In_1730);
nand U2961 (N_2961,In_1155,In_1981);
or U2962 (N_2962,In_1329,In_2341);
xor U2963 (N_2963,In_1697,In_1902);
and U2964 (N_2964,In_1107,In_2973);
and U2965 (N_2965,In_2478,In_879);
nor U2966 (N_2966,In_12,In_2979);
and U2967 (N_2967,In_1879,In_1496);
xor U2968 (N_2968,In_1257,In_2953);
or U2969 (N_2969,In_1858,In_1166);
or U2970 (N_2970,In_44,In_1952);
xor U2971 (N_2971,In_1698,In_2003);
nand U2972 (N_2972,In_251,In_626);
or U2973 (N_2973,In_593,In_1231);
nor U2974 (N_2974,In_2939,In_317);
nor U2975 (N_2975,In_32,In_1971);
or U2976 (N_2976,In_1588,In_1676);
or U2977 (N_2977,In_1449,In_2639);
and U2978 (N_2978,In_285,In_902);
xnor U2979 (N_2979,In_479,In_2679);
or U2980 (N_2980,In_576,In_2351);
or U2981 (N_2981,In_697,In_2042);
or U2982 (N_2982,In_543,In_499);
nand U2983 (N_2983,In_1868,In_1872);
or U2984 (N_2984,In_2079,In_1393);
nand U2985 (N_2985,In_2972,In_1332);
or U2986 (N_2986,In_1539,In_763);
nand U2987 (N_2987,In_593,In_939);
nand U2988 (N_2988,In_948,In_2646);
and U2989 (N_2989,In_445,In_2777);
or U2990 (N_2990,In_1852,In_660);
and U2991 (N_2991,In_2328,In_2785);
nand U2992 (N_2992,In_1157,In_2821);
xor U2993 (N_2993,In_93,In_1767);
or U2994 (N_2994,In_932,In_2620);
and U2995 (N_2995,In_720,In_1165);
xor U2996 (N_2996,In_763,In_2477);
xnor U2997 (N_2997,In_1455,In_1701);
nand U2998 (N_2998,In_430,In_311);
nor U2999 (N_2999,In_2277,In_2777);
xnor U3000 (N_3000,N_1540,N_2753);
xnor U3001 (N_3001,N_2280,N_696);
xnor U3002 (N_3002,N_634,N_2078);
nor U3003 (N_3003,N_2223,N_2289);
xnor U3004 (N_3004,N_1180,N_405);
nor U3005 (N_3005,N_2844,N_1516);
and U3006 (N_3006,N_1442,N_2936);
or U3007 (N_3007,N_2946,N_156);
nor U3008 (N_3008,N_1880,N_1052);
xnor U3009 (N_3009,N_2443,N_2402);
or U3010 (N_3010,N_856,N_700);
nand U3011 (N_3011,N_751,N_2530);
and U3012 (N_3012,N_671,N_1847);
xor U3013 (N_3013,N_692,N_1168);
nor U3014 (N_3014,N_30,N_2645);
or U3015 (N_3015,N_348,N_698);
nand U3016 (N_3016,N_2252,N_250);
xor U3017 (N_3017,N_1494,N_2145);
or U3018 (N_3018,N_609,N_1688);
nor U3019 (N_3019,N_943,N_1261);
nor U3020 (N_3020,N_799,N_212);
nor U3021 (N_3021,N_782,N_2096);
and U3022 (N_3022,N_529,N_2260);
nor U3023 (N_3023,N_1267,N_1395);
nor U3024 (N_3024,N_1003,N_1697);
xor U3025 (N_3025,N_2425,N_594);
nand U3026 (N_3026,N_1485,N_1088);
xnor U3027 (N_3027,N_849,N_2056);
and U3028 (N_3028,N_226,N_2921);
nand U3029 (N_3029,N_1557,N_711);
nor U3030 (N_3030,N_2549,N_2864);
xor U3031 (N_3031,N_1200,N_1407);
and U3032 (N_3032,N_738,N_1080);
nor U3033 (N_3033,N_2878,N_658);
or U3034 (N_3034,N_2734,N_2849);
and U3035 (N_3035,N_666,N_1888);
or U3036 (N_3036,N_1171,N_320);
nand U3037 (N_3037,N_651,N_1372);
or U3038 (N_3038,N_1857,N_1574);
nor U3039 (N_3039,N_688,N_999);
and U3040 (N_3040,N_1464,N_2118);
xor U3041 (N_3041,N_1301,N_520);
nor U3042 (N_3042,N_2546,N_2344);
xnor U3043 (N_3043,N_2746,N_884);
nor U3044 (N_3044,N_191,N_456);
or U3045 (N_3045,N_1678,N_2342);
and U3046 (N_3046,N_495,N_558);
xnor U3047 (N_3047,N_19,N_926);
nor U3048 (N_3048,N_1863,N_1957);
nand U3049 (N_3049,N_141,N_79);
nand U3050 (N_3050,N_2710,N_2042);
nor U3051 (N_3051,N_1791,N_915);
and U3052 (N_3052,N_1138,N_2147);
xor U3053 (N_3053,N_2677,N_1446);
or U3054 (N_3054,N_2744,N_483);
nand U3055 (N_3055,N_112,N_961);
xnor U3056 (N_3056,N_531,N_2940);
nand U3057 (N_3057,N_1081,N_1854);
nor U3058 (N_3058,N_2156,N_2200);
nand U3059 (N_3059,N_177,N_2061);
and U3060 (N_3060,N_794,N_1490);
and U3061 (N_3061,N_2644,N_1876);
or U3062 (N_3062,N_218,N_693);
nor U3063 (N_3063,N_2025,N_619);
nor U3064 (N_3064,N_1103,N_1815);
nor U3065 (N_3065,N_1367,N_1821);
xnor U3066 (N_3066,N_822,N_1343);
or U3067 (N_3067,N_874,N_2509);
nor U3068 (N_3068,N_2621,N_2304);
or U3069 (N_3069,N_290,N_1762);
nor U3070 (N_3070,N_2384,N_304);
nand U3071 (N_3071,N_2949,N_633);
and U3072 (N_3072,N_2133,N_2616);
nor U3073 (N_3073,N_1070,N_970);
or U3074 (N_3074,N_1443,N_121);
xnor U3075 (N_3075,N_2323,N_1590);
nand U3076 (N_3076,N_2081,N_2293);
or U3077 (N_3077,N_942,N_154);
nand U3078 (N_3078,N_2242,N_2122);
or U3079 (N_3079,N_418,N_2937);
nand U3080 (N_3080,N_1513,N_2092);
nor U3081 (N_3081,N_1592,N_2718);
xor U3082 (N_3082,N_2682,N_2222);
nor U3083 (N_3083,N_78,N_287);
nor U3084 (N_3084,N_65,N_2015);
nor U3085 (N_3085,N_1227,N_229);
or U3086 (N_3086,N_727,N_1292);
nor U3087 (N_3087,N_1403,N_1561);
nand U3088 (N_3088,N_244,N_1056);
or U3089 (N_3089,N_1046,N_2451);
nor U3090 (N_3090,N_1584,N_302);
and U3091 (N_3091,N_1351,N_385);
or U3092 (N_3092,N_2121,N_1541);
or U3093 (N_3093,N_2310,N_2766);
nor U3094 (N_3094,N_2972,N_1708);
nand U3095 (N_3095,N_1458,N_99);
nor U3096 (N_3096,N_2050,N_446);
nand U3097 (N_3097,N_1444,N_1441);
nand U3098 (N_3098,N_1251,N_1600);
nand U3099 (N_3099,N_2899,N_1648);
nand U3100 (N_3100,N_2841,N_2966);
nand U3101 (N_3101,N_323,N_2129);
and U3102 (N_3102,N_1693,N_754);
and U3103 (N_3103,N_2307,N_2220);
or U3104 (N_3104,N_1189,N_2195);
nor U3105 (N_3105,N_1657,N_424);
nand U3106 (N_3106,N_840,N_2435);
xor U3107 (N_3107,N_2205,N_2194);
nand U3108 (N_3108,N_847,N_1994);
and U3109 (N_3109,N_863,N_114);
or U3110 (N_3110,N_1448,N_917);
or U3111 (N_3111,N_1624,N_2089);
xnor U3112 (N_3112,N_2218,N_243);
and U3113 (N_3113,N_51,N_438);
and U3114 (N_3114,N_4,N_491);
and U3115 (N_3115,N_1828,N_480);
and U3116 (N_3116,N_997,N_901);
nand U3117 (N_3117,N_538,N_2005);
nand U3118 (N_3118,N_1698,N_629);
and U3119 (N_3119,N_1755,N_182);
nor U3120 (N_3120,N_1431,N_861);
and U3121 (N_3121,N_2641,N_518);
nand U3122 (N_3122,N_1342,N_360);
xnor U3123 (N_3123,N_2582,N_1986);
or U3124 (N_3124,N_2700,N_2320);
xnor U3125 (N_3125,N_2594,N_1113);
or U3126 (N_3126,N_2519,N_956);
or U3127 (N_3127,N_1595,N_1997);
nand U3128 (N_3128,N_878,N_1996);
and U3129 (N_3129,N_2680,N_1398);
or U3130 (N_3130,N_2774,N_1029);
nand U3131 (N_3131,N_268,N_1521);
xnor U3132 (N_3132,N_398,N_1535);
nand U3133 (N_3133,N_1026,N_2484);
or U3134 (N_3134,N_625,N_703);
xor U3135 (N_3135,N_1417,N_1701);
nor U3136 (N_3136,N_1524,N_2593);
xnor U3137 (N_3137,N_1706,N_477);
nor U3138 (N_3138,N_2747,N_967);
or U3139 (N_3139,N_1900,N_2836);
or U3140 (N_3140,N_953,N_1047);
nand U3141 (N_3141,N_2834,N_195);
nor U3142 (N_3142,N_2748,N_932);
and U3143 (N_3143,N_1817,N_1651);
nand U3144 (N_3144,N_329,N_1157);
xor U3145 (N_3145,N_2498,N_353);
and U3146 (N_3146,N_1622,N_138);
nor U3147 (N_3147,N_2206,N_2625);
nor U3148 (N_3148,N_68,N_2591);
xnor U3149 (N_3149,N_399,N_2894);
or U3150 (N_3150,N_2948,N_1747);
nor U3151 (N_3151,N_725,N_2552);
nand U3152 (N_3152,N_2770,N_2910);
xnor U3153 (N_3153,N_2571,N_1455);
xor U3154 (N_3154,N_2230,N_2165);
xnor U3155 (N_3155,N_2555,N_1898);
xnor U3156 (N_3156,N_2161,N_2455);
xor U3157 (N_3157,N_2332,N_1468);
nand U3158 (N_3158,N_1575,N_110);
or U3159 (N_3159,N_2995,N_325);
nand U3160 (N_3160,N_2866,N_1314);
xnor U3161 (N_3161,N_2634,N_172);
and U3162 (N_3162,N_1077,N_2450);
nor U3163 (N_3163,N_1843,N_1633);
nand U3164 (N_3164,N_784,N_139);
and U3165 (N_3165,N_463,N_1288);
nor U3166 (N_3166,N_548,N_2904);
or U3167 (N_3167,N_41,N_2462);
xor U3168 (N_3168,N_663,N_2011);
or U3169 (N_3169,N_1718,N_769);
nand U3170 (N_3170,N_2742,N_2655);
nor U3171 (N_3171,N_2585,N_277);
nand U3172 (N_3172,N_1366,N_1766);
nand U3173 (N_3173,N_789,N_2422);
and U3174 (N_3174,N_1660,N_2236);
xnor U3175 (N_3175,N_1319,N_1296);
nand U3176 (N_3176,N_2523,N_1385);
nor U3177 (N_3177,N_437,N_1761);
xor U3178 (N_3178,N_1445,N_2597);
or U3179 (N_3179,N_337,N_2541);
nand U3180 (N_3180,N_1040,N_507);
or U3181 (N_3181,N_931,N_2590);
nor U3182 (N_3182,N_2690,N_2883);
or U3183 (N_3183,N_1402,N_1093);
nand U3184 (N_3184,N_339,N_1944);
nand U3185 (N_3185,N_321,N_2939);
and U3186 (N_3186,N_860,N_2798);
xnor U3187 (N_3187,N_36,N_1379);
nand U3188 (N_3188,N_2146,N_188);
and U3189 (N_3189,N_149,N_2279);
nand U3190 (N_3190,N_1938,N_285);
or U3191 (N_3191,N_1105,N_2855);
xnor U3192 (N_3192,N_793,N_1325);
and U3193 (N_3193,N_1998,N_1295);
nor U3194 (N_3194,N_1545,N_88);
nor U3195 (N_3195,N_2657,N_2814);
nand U3196 (N_3196,N_659,N_1069);
nor U3197 (N_3197,N_905,N_2415);
nor U3198 (N_3198,N_2013,N_2363);
and U3199 (N_3199,N_642,N_1065);
xnor U3200 (N_3200,N_26,N_1289);
nand U3201 (N_3201,N_755,N_1714);
or U3202 (N_3202,N_610,N_275);
xor U3203 (N_3203,N_2063,N_20);
nor U3204 (N_3204,N_2232,N_1038);
nand U3205 (N_3205,N_2022,N_836);
nand U3206 (N_3206,N_2067,N_1582);
and U3207 (N_3207,N_1330,N_2369);
nor U3208 (N_3208,N_983,N_2857);
nand U3209 (N_3209,N_1753,N_1045);
xnor U3210 (N_3210,N_1087,N_924);
nor U3211 (N_3211,N_717,N_591);
and U3212 (N_3212,N_2362,N_1016);
nand U3213 (N_3213,N_2475,N_1380);
xor U3214 (N_3214,N_1376,N_39);
and U3215 (N_3215,N_307,N_1836);
xor U3216 (N_3216,N_1341,N_1119);
or U3217 (N_3217,N_2665,N_862);
xor U3218 (N_3218,N_572,N_873);
or U3219 (N_3219,N_1223,N_2326);
or U3220 (N_3220,N_2557,N_387);
xor U3221 (N_3221,N_1160,N_1118);
and U3222 (N_3222,N_165,N_912);
or U3223 (N_3223,N_2752,N_1306);
xor U3224 (N_3224,N_2155,N_221);
xnor U3225 (N_3225,N_222,N_1043);
nor U3226 (N_3226,N_220,N_371);
xor U3227 (N_3227,N_1750,N_1902);
nand U3228 (N_3228,N_240,N_1084);
and U3229 (N_3229,N_301,N_2273);
xor U3230 (N_3230,N_2970,N_971);
nor U3231 (N_3231,N_1795,N_649);
or U3232 (N_3232,N_723,N_305);
xor U3233 (N_3233,N_1129,N_2292);
or U3234 (N_3234,N_1484,N_1155);
nor U3235 (N_3235,N_994,N_1941);
nor U3236 (N_3236,N_1014,N_2378);
nor U3237 (N_3237,N_1619,N_2704);
nand U3238 (N_3238,N_2691,N_1775);
or U3239 (N_3239,N_1260,N_8);
and U3240 (N_3240,N_1607,N_2882);
nand U3241 (N_3241,N_1601,N_2246);
and U3242 (N_3242,N_1765,N_2652);
nor U3243 (N_3243,N_2167,N_179);
nor U3244 (N_3244,N_2745,N_1165);
nor U3245 (N_3245,N_2901,N_1790);
nor U3246 (N_3246,N_365,N_313);
and U3247 (N_3247,N_1562,N_473);
nor U3248 (N_3248,N_429,N_330);
nor U3249 (N_3249,N_1573,N_2642);
nor U3250 (N_3250,N_1375,N_780);
or U3251 (N_3251,N_2932,N_1534);
and U3252 (N_3252,N_2938,N_656);
or U3253 (N_3253,N_498,N_1426);
or U3254 (N_3254,N_2202,N_13);
or U3255 (N_3255,N_426,N_823);
xor U3256 (N_3256,N_270,N_271);
and U3257 (N_3257,N_1886,N_45);
nor U3258 (N_3258,N_181,N_2446);
and U3259 (N_3259,N_1659,N_2093);
and U3260 (N_3260,N_600,N_1694);
nand U3261 (N_3261,N_2391,N_2083);
nor U3262 (N_3262,N_601,N_344);
nand U3263 (N_3263,N_2695,N_2674);
and U3264 (N_3264,N_621,N_2076);
xor U3265 (N_3265,N_362,N_544);
xnor U3266 (N_3266,N_1020,N_208);
xnor U3267 (N_3267,N_1671,N_959);
nor U3268 (N_3268,N_273,N_1699);
xnor U3269 (N_3269,N_1895,N_1037);
and U3270 (N_3270,N_567,N_2379);
xor U3271 (N_3271,N_2701,N_1005);
and U3272 (N_3272,N_2685,N_1391);
or U3273 (N_3273,N_1856,N_939);
nand U3274 (N_3274,N_2812,N_1629);
xnor U3275 (N_3275,N_389,N_1917);
or U3276 (N_3276,N_2683,N_1191);
xnor U3277 (N_3277,N_1906,N_1277);
or U3278 (N_3278,N_11,N_2912);
nor U3279 (N_3279,N_962,N_2891);
nor U3280 (N_3280,N_1204,N_1705);
xnor U3281 (N_3281,N_257,N_1304);
xor U3282 (N_3282,N_1309,N_2653);
xor U3283 (N_3283,N_23,N_2212);
or U3284 (N_3284,N_2851,N_1335);
and U3285 (N_3285,N_644,N_2012);
or U3286 (N_3286,N_2009,N_1550);
nand U3287 (N_3287,N_537,N_2113);
and U3288 (N_3288,N_74,N_982);
nor U3289 (N_3289,N_1058,N_2268);
and U3290 (N_3290,N_710,N_687);
or U3291 (N_3291,N_2233,N_70);
nand U3292 (N_3292,N_234,N_826);
xor U3293 (N_3293,N_71,N_2054);
xnor U3294 (N_3294,N_2244,N_660);
nor U3295 (N_3295,N_318,N_2299);
and U3296 (N_3296,N_664,N_811);
and U3297 (N_3297,N_2565,N_233);
and U3298 (N_3298,N_167,N_2470);
xor U3299 (N_3299,N_1672,N_963);
nand U3300 (N_3300,N_311,N_2262);
and U3301 (N_3301,N_2296,N_1499);
xnor U3302 (N_3302,N_771,N_2333);
and U3303 (N_3303,N_260,N_2478);
nand U3304 (N_3304,N_1389,N_2278);
nand U3305 (N_3305,N_1780,N_1411);
or U3306 (N_3306,N_2285,N_2860);
or U3307 (N_3307,N_2238,N_2809);
and U3308 (N_3308,N_2783,N_2131);
and U3309 (N_3309,N_2769,N_2908);
xnor U3310 (N_3310,N_1787,N_2623);
or U3311 (N_3311,N_124,N_1415);
and U3312 (N_3312,N_2397,N_1337);
and U3313 (N_3313,N_207,N_2713);
and U3314 (N_3314,N_185,N_2294);
nand U3315 (N_3315,N_2420,N_1572);
nand U3316 (N_3316,N_204,N_2457);
nor U3317 (N_3317,N_2771,N_1220);
or U3318 (N_3318,N_1205,N_2465);
and U3319 (N_3319,N_2108,N_487);
nor U3320 (N_3320,N_2620,N_2466);
xnor U3321 (N_3321,N_1800,N_408);
xnor U3322 (N_3322,N_1209,N_80);
or U3323 (N_3323,N_109,N_2884);
xnor U3324 (N_3324,N_1523,N_2082);
nand U3325 (N_3325,N_1814,N_2804);
xnor U3326 (N_3326,N_331,N_800);
and U3327 (N_3327,N_2002,N_2302);
xor U3328 (N_3328,N_2309,N_2241);
xnor U3329 (N_3329,N_388,N_2168);
and U3330 (N_3330,N_841,N_2432);
xnor U3331 (N_3331,N_582,N_2417);
nand U3332 (N_3332,N_1300,N_338);
nor U3333 (N_3333,N_486,N_702);
nor U3334 (N_3334,N_872,N_460);
nand U3335 (N_3335,N_1109,N_2749);
nand U3336 (N_3336,N_2149,N_383);
nor U3337 (N_3337,N_1438,N_173);
nor U3338 (N_3338,N_433,N_731);
nand U3339 (N_3339,N_2604,N_1684);
nand U3340 (N_3340,N_1594,N_1786);
nor U3341 (N_3341,N_1918,N_364);
nand U3342 (N_3342,N_81,N_1569);
and U3343 (N_3343,N_2351,N_361);
xnor U3344 (N_3344,N_1675,N_380);
and U3345 (N_3345,N_411,N_401);
or U3346 (N_3346,N_2654,N_2984);
nand U3347 (N_3347,N_2837,N_1329);
and U3348 (N_3348,N_1782,N_2576);
nor U3349 (N_3349,N_1525,N_458);
nor U3350 (N_3350,N_1263,N_527);
nor U3351 (N_3351,N_464,N_1641);
nand U3352 (N_3352,N_1988,N_1636);
or U3353 (N_3353,N_1646,N_1454);
nand U3354 (N_3354,N_2255,N_1152);
or U3355 (N_3355,N_2761,N_2471);
xnor U3356 (N_3356,N_2449,N_607);
nor U3357 (N_3357,N_2479,N_2322);
and U3358 (N_3358,N_2324,N_1608);
nor U3359 (N_3359,N_1252,N_2992);
nand U3360 (N_3360,N_540,N_231);
nor U3361 (N_3361,N_2787,N_804);
or U3362 (N_3362,N_2057,N_1015);
xor U3363 (N_3363,N_1502,N_535);
xor U3364 (N_3364,N_2338,N_2711);
xnor U3365 (N_3365,N_1363,N_984);
or U3366 (N_3366,N_2829,N_1127);
xnor U3367 (N_3367,N_470,N_2876);
xor U3368 (N_3368,N_2068,N_1169);
nor U3369 (N_3369,N_707,N_2215);
or U3370 (N_3370,N_239,N_118);
xor U3371 (N_3371,N_201,N_369);
nor U3372 (N_3372,N_1825,N_2073);
xor U3373 (N_3373,N_1617,N_1982);
nand U3374 (N_3374,N_2234,N_1203);
or U3375 (N_3375,N_1228,N_1433);
and U3376 (N_3376,N_1298,N_249);
nor U3377 (N_3377,N_1001,N_2825);
or U3378 (N_3378,N_1222,N_837);
xnor U3379 (N_3379,N_1456,N_1831);
and U3380 (N_3380,N_2403,N_1471);
and U3381 (N_3381,N_1904,N_779);
and U3382 (N_3382,N_1849,N_1007);
nor U3383 (N_3383,N_1287,N_131);
xor U3384 (N_3384,N_2738,N_2724);
and U3385 (N_3385,N_35,N_2335);
xnor U3386 (N_3386,N_363,N_263);
and U3387 (N_3387,N_2612,N_2835);
nor U3388 (N_3388,N_2157,N_569);
xor U3389 (N_3389,N_1530,N_1870);
nor U3390 (N_3390,N_2491,N_1509);
nor U3391 (N_3391,N_1842,N_2586);
nor U3392 (N_3392,N_1560,N_2980);
and U3393 (N_3393,N_1235,N_2132);
nand U3394 (N_3394,N_562,N_2003);
nand U3395 (N_3395,N_2705,N_1593);
and U3396 (N_3396,N_2914,N_1409);
nand U3397 (N_3397,N_868,N_1793);
xnor U3398 (N_3398,N_695,N_922);
nor U3399 (N_3399,N_76,N_1949);
and U3400 (N_3400,N_1334,N_1776);
xor U3401 (N_3401,N_1618,N_772);
nor U3402 (N_3402,N_2865,N_791);
and U3403 (N_3403,N_989,N_2563);
xnor U3404 (N_3404,N_620,N_876);
or U3405 (N_3405,N_1019,N_2381);
xnor U3406 (N_3406,N_504,N_596);
and U3407 (N_3407,N_1835,N_1023);
xnor U3408 (N_3408,N_1242,N_266);
nand U3409 (N_3409,N_1208,N_2201);
or U3410 (N_3410,N_2554,N_2024);
and U3411 (N_3411,N_1769,N_1808);
xor U3412 (N_3412,N_2085,N_386);
or U3413 (N_3413,N_1278,N_816);
xnor U3414 (N_3414,N_2021,N_91);
and U3415 (N_3415,N_194,N_2906);
or U3416 (N_3416,N_357,N_2447);
xnor U3417 (N_3417,N_1813,N_1217);
nand U3418 (N_3418,N_1489,N_2830);
or U3419 (N_3419,N_393,N_603);
or U3420 (N_3420,N_449,N_52);
or U3421 (N_3421,N_1905,N_1115);
xor U3422 (N_3422,N_828,N_2151);
nand U3423 (N_3423,N_2848,N_2524);
or U3424 (N_3424,N_102,N_1172);
nand U3425 (N_3425,N_1491,N_825);
nor U3426 (N_3426,N_2315,N_1164);
and U3427 (N_3427,N_2531,N_2072);
nor U3428 (N_3428,N_2956,N_973);
or U3429 (N_3429,N_1819,N_299);
xnor U3430 (N_3430,N_1274,N_2030);
or U3431 (N_3431,N_2567,N_1);
nand U3432 (N_3432,N_1744,N_467);
or U3433 (N_3433,N_734,N_713);
xnor U3434 (N_3434,N_579,N_2365);
nand U3435 (N_3435,N_2895,N_199);
xnor U3436 (N_3436,N_2510,N_2873);
nor U3437 (N_3437,N_683,N_98);
nand U3438 (N_3438,N_103,N_2803);
or U3439 (N_3439,N_728,N_47);
nand U3440 (N_3440,N_2224,N_2460);
nand U3441 (N_3441,N_1211,N_2091);
nor U3442 (N_3442,N_1789,N_210);
or U3443 (N_3443,N_1554,N_2330);
nor U3444 (N_3444,N_1614,N_1925);
nor U3445 (N_3445,N_701,N_2776);
xnor U3446 (N_3446,N_2395,N_2796);
nand U3447 (N_3447,N_1658,N_281);
nor U3448 (N_3448,N_2094,N_245);
and U3449 (N_3449,N_2823,N_729);
or U3450 (N_3450,N_2660,N_359);
xor U3451 (N_3451,N_2144,N_1885);
or U3452 (N_3452,N_1627,N_632);
or U3453 (N_3453,N_1632,N_2917);
xor U3454 (N_3454,N_1059,N_190);
nor U3455 (N_3455,N_536,N_1585);
and U3456 (N_3456,N_3,N_180);
xnor U3457 (N_3457,N_1686,N_2400);
or U3458 (N_3458,N_1867,N_2649);
nor U3459 (N_3459,N_500,N_974);
nand U3460 (N_3460,N_2055,N_2473);
xnor U3461 (N_3461,N_2811,N_2556);
nor U3462 (N_3462,N_740,N_272);
and U3463 (N_3463,N_1841,N_2628);
xnor U3464 (N_3464,N_1929,N_946);
or U3465 (N_3465,N_1432,N_309);
and U3466 (N_3466,N_2547,N_1044);
and U3467 (N_3467,N_1060,N_888);
nand U3468 (N_3468,N_1427,N_1071);
xor U3469 (N_3469,N_2458,N_2308);
and U3470 (N_3470,N_546,N_1816);
nor U3471 (N_3471,N_1810,N_2633);
xnor U3472 (N_3472,N_1186,N_748);
nor U3473 (N_3473,N_17,N_1935);
and U3474 (N_3474,N_2944,N_77);
nand U3475 (N_3475,N_434,N_2999);
or U3476 (N_3476,N_143,N_1284);
and U3477 (N_3477,N_413,N_1230);
nor U3478 (N_3478,N_2854,N_2592);
nand U3479 (N_3479,N_247,N_1979);
xnor U3480 (N_3480,N_2440,N_1096);
or U3481 (N_3481,N_889,N_1853);
xor U3482 (N_3482,N_2784,N_1262);
and U3483 (N_3483,N_2902,N_1269);
or U3484 (N_3484,N_1591,N_101);
and U3485 (N_3485,N_2756,N_1921);
nand U3486 (N_3486,N_2243,N_1995);
nor U3487 (N_3487,N_2943,N_2905);
nand U3488 (N_3488,N_1482,N_1662);
nand U3489 (N_3489,N_1803,N_1645);
nand U3490 (N_3490,N_2824,N_1745);
or U3491 (N_3491,N_639,N_2225);
nor U3492 (N_3492,N_1511,N_1146);
and U3493 (N_3493,N_1599,N_265);
xnor U3494 (N_3494,N_1374,N_1357);
nand U3495 (N_3495,N_871,N_1072);
nand U3496 (N_3496,N_817,N_2916);
nand U3497 (N_3497,N_134,N_454);
xnor U3498 (N_3498,N_1067,N_564);
xnor U3499 (N_3499,N_376,N_2903);
and U3500 (N_3500,N_1259,N_1156);
xnor U3501 (N_3501,N_1650,N_801);
or U3502 (N_3502,N_928,N_1805);
or U3503 (N_3503,N_2964,N_1449);
xnor U3504 (N_3504,N_170,N_1830);
nand U3505 (N_3505,N_1392,N_2116);
or U3506 (N_3506,N_1307,N_528);
and U3507 (N_3507,N_2605,N_2689);
nand U3508 (N_3508,N_1669,N_2659);
xor U3509 (N_3509,N_451,N_499);
nand U3510 (N_3510,N_2210,N_1095);
xor U3511 (N_3511,N_2269,N_2303);
and U3512 (N_3512,N_1634,N_2253);
nor U3513 (N_3513,N_1009,N_2639);
nand U3514 (N_3514,N_2788,N_1587);
xnor U3515 (N_3515,N_897,N_1476);
and U3516 (N_3516,N_147,N_892);
and U3517 (N_3517,N_778,N_2707);
nor U3518 (N_3518,N_798,N_2990);
xor U3519 (N_3519,N_1954,N_264);
and U3520 (N_3520,N_2931,N_2859);
and U3521 (N_3521,N_1838,N_2062);
and U3522 (N_3522,N_2007,N_1723);
nand U3523 (N_3523,N_2584,N_2717);
xor U3524 (N_3524,N_2885,N_501);
xor U3525 (N_3525,N_18,N_2482);
or U3526 (N_3526,N_1159,N_818);
or U3527 (N_3527,N_1664,N_2404);
nand U3528 (N_3528,N_2383,N_1899);
and U3529 (N_3529,N_16,N_1350);
nor U3530 (N_3530,N_957,N_745);
nand U3531 (N_3531,N_914,N_2773);
nor U3532 (N_3532,N_1360,N_1420);
nor U3533 (N_3533,N_1518,N_830);
nor U3534 (N_3534,N_2152,N_2401);
or U3535 (N_3535,N_764,N_274);
nand U3536 (N_3536,N_435,N_0);
nor U3537 (N_3537,N_2512,N_602);
nand U3538 (N_3538,N_2598,N_1283);
and U3539 (N_3539,N_677,N_584);
or U3540 (N_3540,N_2545,N_851);
or U3541 (N_3541,N_1216,N_902);
nand U3542 (N_3542,N_1537,N_2553);
and U3543 (N_3543,N_614,N_2272);
xnor U3544 (N_3544,N_2953,N_189);
xnor U3545 (N_3545,N_1151,N_2719);
nand U3546 (N_3546,N_227,N_877);
nor U3547 (N_3547,N_414,N_2095);
nor U3548 (N_3548,N_373,N_724);
nor U3549 (N_3549,N_2575,N_2712);
xor U3550 (N_3550,N_1031,N_162);
or U3551 (N_3551,N_298,N_1355);
or U3552 (N_3552,N_2474,N_2688);
and U3553 (N_3553,N_2892,N_1543);
xor U3554 (N_3554,N_1352,N_948);
and U3555 (N_3555,N_1596,N_2153);
nand U3556 (N_3556,N_469,N_2636);
nand U3557 (N_3557,N_106,N_56);
xnor U3558 (N_3558,N_1233,N_2044);
or U3559 (N_3559,N_2040,N_1757);
xor U3560 (N_3560,N_2254,N_598);
nor U3561 (N_3561,N_2137,N_1520);
and U3562 (N_3562,N_2373,N_2010);
and U3563 (N_3563,N_524,N_2918);
nor U3564 (N_3564,N_2331,N_1879);
nand U3565 (N_3565,N_2786,N_2375);
xnor U3566 (N_3566,N_1408,N_1422);
or U3567 (N_3567,N_214,N_2270);
xnor U3568 (N_3568,N_1924,N_1275);
or U3569 (N_3569,N_2314,N_2416);
nor U3570 (N_3570,N_2227,N_916);
and U3571 (N_3571,N_815,N_1128);
xor U3572 (N_3572,N_2023,N_2480);
nor U3573 (N_3573,N_1013,N_1201);
and U3574 (N_3574,N_1239,N_2101);
or U3575 (N_3575,N_1294,N_1498);
or U3576 (N_3576,N_1397,N_48);
xnor U3577 (N_3577,N_1036,N_2897);
and U3578 (N_3578,N_2481,N_1492);
xnor U3579 (N_3579,N_2679,N_2382);
nor U3580 (N_3580,N_1967,N_186);
nand U3581 (N_3581,N_1394,N_845);
nand U3582 (N_3582,N_2536,N_920);
or U3583 (N_3583,N_705,N_1091);
xor U3584 (N_3584,N_282,N_2228);
or U3585 (N_3585,N_829,N_1042);
and U3586 (N_3586,N_489,N_1971);
xor U3587 (N_3587,N_2877,N_150);
xor U3588 (N_3588,N_2818,N_718);
xnor U3589 (N_3589,N_2764,N_2295);
nor U3590 (N_3590,N_2613,N_144);
xor U3591 (N_3591,N_1193,N_1365);
nand U3592 (N_3592,N_1139,N_184);
nor U3593 (N_3593,N_853,N_958);
and U3594 (N_3594,N_2130,N_699);
and U3595 (N_3595,N_256,N_2539);
or U3596 (N_3596,N_661,N_402);
nand U3597 (N_3597,N_1101,N_1361);
or U3598 (N_3598,N_1655,N_1715);
or U3599 (N_3599,N_1666,N_2433);
or U3600 (N_3600,N_1860,N_1947);
and U3601 (N_3601,N_576,N_2164);
xor U3602 (N_3602,N_812,N_648);
or U3603 (N_3603,N_2638,N_904);
xor U3604 (N_3604,N_1048,N_883);
xnor U3605 (N_3605,N_1923,N_2485);
xor U3606 (N_3606,N_541,N_2573);
or U3607 (N_3607,N_315,N_107);
nor U3608 (N_3608,N_2951,N_2434);
xnor U3609 (N_3609,N_2368,N_1952);
or U3610 (N_3610,N_2502,N_1002);
nor U3611 (N_3611,N_2123,N_616);
or U3612 (N_3612,N_1099,N_2352);
nor U3613 (N_3613,N_1192,N_1735);
xnor U3614 (N_3614,N_2399,N_203);
nor U3615 (N_3615,N_108,N_2842);
nand U3616 (N_3616,N_1570,N_2204);
nand U3617 (N_3617,N_1567,N_2551);
nand U3618 (N_3618,N_2431,N_2821);
xor U3619 (N_3619,N_1248,N_2240);
or U3620 (N_3620,N_2740,N_2669);
or U3621 (N_3621,N_137,N_2698);
nand U3622 (N_3622,N_1308,N_1054);
nand U3623 (N_3623,N_899,N_462);
and U3624 (N_3624,N_1090,N_2175);
and U3625 (N_3625,N_117,N_1625);
or U3626 (N_3626,N_237,N_2799);
nor U3627 (N_3627,N_136,N_749);
nor U3628 (N_3628,N_606,N_2110);
nand U3629 (N_3629,N_21,N_2736);
nand U3630 (N_3630,N_288,N_57);
and U3631 (N_3631,N_1290,N_228);
or U3632 (N_3632,N_2961,N_2780);
nor U3633 (N_3633,N_479,N_267);
or U3634 (N_3634,N_1637,N_2406);
xnor U3635 (N_3635,N_2316,N_838);
xnor U3636 (N_3636,N_773,N_2467);
and U3637 (N_3637,N_720,N_1506);
xor U3638 (N_3638,N_291,N_1317);
and U3639 (N_3639,N_511,N_1527);
and U3640 (N_3640,N_1396,N_1089);
or U3641 (N_3641,N_1920,N_2495);
nand U3642 (N_3642,N_84,N_1927);
nor U3643 (N_3643,N_623,N_503);
or U3644 (N_3644,N_2978,N_2472);
and U3645 (N_3645,N_2800,N_1772);
xor U3646 (N_3646,N_2806,N_1400);
and U3647 (N_3647,N_690,N_1362);
nand U3648 (N_3648,N_1558,N_89);
nand U3649 (N_3649,N_1187,N_910);
nor U3650 (N_3650,N_2128,N_708);
nor U3651 (N_3651,N_410,N_1206);
and U3652 (N_3652,N_1677,N_2900);
xnor U3653 (N_3653,N_2596,N_2488);
and U3654 (N_3654,N_2358,N_1597);
xor U3655 (N_3655,N_157,N_542);
nand U3656 (N_3656,N_1977,N_1388);
and U3657 (N_3657,N_43,N_1640);
or U3658 (N_3658,N_1852,N_1401);
xor U3659 (N_3659,N_15,N_938);
nor U3660 (N_3660,N_1344,N_471);
nand U3661 (N_3661,N_834,N_2436);
nand U3662 (N_3662,N_1167,N_2927);
nor U3663 (N_3663,N_977,N_797);
or U3664 (N_3664,N_295,N_2182);
or U3665 (N_3665,N_1406,N_918);
and U3666 (N_3666,N_1066,N_1194);
nand U3667 (N_3667,N_2199,N_2611);
nand U3668 (N_3668,N_882,N_640);
nand U3669 (N_3669,N_2993,N_2987);
nor U3670 (N_3670,N_732,N_1881);
and U3671 (N_3671,N_2709,N_1215);
or U3672 (N_3672,N_2935,N_2615);
nor U3673 (N_3673,N_317,N_608);
and U3674 (N_3674,N_762,N_349);
xnor U3675 (N_3675,N_382,N_1690);
nand U3676 (N_3676,N_404,N_523);
and U3677 (N_3677,N_1626,N_796);
xor U3678 (N_3678,N_1487,N_1707);
xnor U3679 (N_3679,N_1279,N_911);
nand U3680 (N_3680,N_1429,N_1313);
xnor U3681 (N_3681,N_2911,N_2257);
nand U3682 (N_3682,N_1751,N_2192);
and U3683 (N_3683,N_2359,N_1726);
and U3684 (N_3684,N_492,N_176);
nor U3685 (N_3685,N_2163,N_421);
and U3686 (N_3686,N_2059,N_2245);
nor U3687 (N_3687,N_2656,N_2869);
or U3688 (N_3688,N_2439,N_2832);
or U3689 (N_3689,N_2881,N_2208);
and U3690 (N_3690,N_891,N_1345);
and U3691 (N_3691,N_526,N_308);
nor U3692 (N_3692,N_2696,N_1983);
and U3693 (N_3693,N_1926,N_776);
or U3694 (N_3694,N_2329,N_2052);
nand U3695 (N_3695,N_341,N_2751);
nor U3696 (N_3696,N_2513,N_1844);
nor U3697 (N_3697,N_969,N_1804);
xor U3698 (N_3698,N_2924,N_354);
nor U3699 (N_3699,N_2725,N_1875);
and U3700 (N_3700,N_1889,N_280);
nor U3701 (N_3701,N_1654,N_2544);
nor U3702 (N_3702,N_954,N_1387);
nor U3703 (N_3703,N_1551,N_907);
or U3704 (N_3704,N_1890,N_1945);
and U3705 (N_3705,N_209,N_1124);
and U3706 (N_3706,N_1249,N_1579);
nand U3707 (N_3707,N_1333,N_1531);
nand U3708 (N_3708,N_1234,N_1237);
xor U3709 (N_3709,N_2261,N_1848);
xnor U3710 (N_3710,N_2650,N_2708);
nand U3711 (N_3711,N_1725,N_650);
xnor U3712 (N_3712,N_2077,N_1685);
nand U3713 (N_3713,N_1488,N_1990);
and U3714 (N_3714,N_2341,N_1145);
nor U3715 (N_3715,N_253,N_757);
nor U3716 (N_3716,N_2568,N_2098);
or U3717 (N_3717,N_2423,N_1131);
nor U3718 (N_3718,N_232,N_921);
nor U3719 (N_3719,N_1612,N_2136);
nor U3720 (N_3720,N_1086,N_33);
and U3721 (N_3721,N_2640,N_1989);
nand U3722 (N_3722,N_1851,N_1111);
xnor U3723 (N_3723,N_2726,N_366);
xor U3724 (N_3724,N_783,N_1613);
or U3725 (N_3725,N_1555,N_1656);
xor U3726 (N_3726,N_1504,N_2618);
xor U3727 (N_3727,N_1332,N_1508);
and U3728 (N_3728,N_372,N_857);
nor U3729 (N_3729,N_1273,N_187);
nor U3730 (N_3730,N_40,N_1428);
nor U3731 (N_3731,N_1229,N_1801);
and U3732 (N_3732,N_164,N_1829);
nor U3733 (N_3733,N_2686,N_1547);
and U3734 (N_3734,N_604,N_1225);
and U3735 (N_3735,N_2452,N_950);
and U3736 (N_3736,N_662,N_976);
nor U3737 (N_3737,N_428,N_1536);
nor U3738 (N_3738,N_390,N_1670);
xor U3739 (N_3739,N_1720,N_2981);
nor U3740 (N_3740,N_1754,N_1074);
xnor U3741 (N_3741,N_1377,N_668);
xnor U3742 (N_3742,N_2380,N_327);
nand U3743 (N_3743,N_2364,N_2276);
nand U3744 (N_3744,N_1779,N_2374);
nor U3745 (N_3745,N_92,N_680);
or U3746 (N_3746,N_2781,N_2410);
xnor U3747 (N_3747,N_2492,N_790);
xnor U3748 (N_3748,N_1068,N_864);
or U3749 (N_3749,N_58,N_1430);
and U3750 (N_3750,N_2064,N_2933);
xor U3751 (N_3751,N_611,N_2750);
xnor U3752 (N_3752,N_1256,N_2274);
or U3753 (N_3753,N_2564,N_515);
nand U3754 (N_3754,N_2020,N_1948);
xnor U3755 (N_3755,N_1497,N_1616);
xnor U3756 (N_3756,N_116,N_2186);
nor U3757 (N_3757,N_2782,N_2394);
and U3758 (N_3758,N_1955,N_259);
nor U3759 (N_3759,N_2355,N_674);
and U3760 (N_3760,N_1964,N_115);
nand U3761 (N_3761,N_806,N_1033);
nor U3762 (N_3762,N_1719,N_2856);
xor U3763 (N_3763,N_368,N_419);
nor U3764 (N_3764,N_1501,N_2448);
nand U3765 (N_3765,N_2772,N_588);
xnor U3766 (N_3766,N_1773,N_1603);
and U3767 (N_3767,N_1353,N_1174);
nor U3768 (N_3768,N_557,N_2561);
nor U3769 (N_3769,N_775,N_1532);
nor U3770 (N_3770,N_2337,N_2666);
xor U3771 (N_3771,N_2071,N_1121);
nor U3772 (N_3772,N_978,N_450);
xor U3773 (N_3773,N_2730,N_1472);
nand U3774 (N_3774,N_2515,N_27);
xor U3775 (N_3775,N_1276,N_1486);
nand U3776 (N_3776,N_2871,N_1028);
nor U3777 (N_3777,N_1758,N_1148);
or U3778 (N_3778,N_1199,N_530);
or U3779 (N_3779,N_2847,N_1100);
xor U3780 (N_3780,N_2499,N_630);
or U3781 (N_3781,N_2203,N_1667);
nand U3782 (N_3782,N_1615,N_2277);
nor U3783 (N_3783,N_2504,N_2217);
and U3784 (N_3784,N_2514,N_2727);
or U3785 (N_3785,N_824,N_1827);
xor U3786 (N_3786,N_2287,N_269);
or U3787 (N_3787,N_563,N_2828);
or U3788 (N_3788,N_2,N_2714);
or U3789 (N_3789,N_552,N_1894);
xnor U3790 (N_3790,N_2115,N_2925);
xor U3791 (N_3791,N_2619,N_2079);
nand U3792 (N_3792,N_758,N_1010);
or U3793 (N_3793,N_1855,N_886);
nor U3794 (N_3794,N_739,N_587);
or U3795 (N_3795,N_2027,N_988);
nor U3796 (N_3796,N_2583,N_2760);
and U3797 (N_3797,N_1611,N_945);
nand U3798 (N_3798,N_1245,N_1478);
nor U3799 (N_3799,N_1942,N_1865);
nor U3800 (N_3800,N_2630,N_2412);
xnor U3801 (N_3801,N_1323,N_2046);
nand U3802 (N_3802,N_1928,N_676);
and U3803 (N_3803,N_2353,N_1144);
nand U3804 (N_3804,N_2159,N_2671);
nor U3805 (N_3805,N_1919,N_2229);
nand U3806 (N_3806,N_37,N_1937);
nor U3807 (N_3807,N_2265,N_908);
nor U3808 (N_3808,N_2794,N_2648);
nand U3809 (N_3809,N_378,N_1721);
or U3810 (N_3810,N_455,N_2879);
nand U3811 (N_3811,N_2543,N_626);
xnor U3812 (N_3812,N_1126,N_597);
xnor U3813 (N_3813,N_506,N_2453);
nand U3814 (N_3814,N_2737,N_235);
nand U3815 (N_3815,N_2532,N_543);
and U3816 (N_3816,N_1459,N_1057);
nor U3817 (N_3817,N_936,N_1250);
nand U3818 (N_3818,N_2388,N_1177);
xor U3819 (N_3819,N_843,N_1709);
or U3820 (N_3820,N_252,N_2075);
nor U3821 (N_3821,N_94,N_2231);
and U3822 (N_3822,N_10,N_1682);
nand U3823 (N_3823,N_2386,N_533);
or U3824 (N_3824,N_2249,N_1514);
and U3825 (N_3825,N_1727,N_2697);
and U3826 (N_3826,N_996,N_986);
nand U3827 (N_3827,N_551,N_2569);
nand U3828 (N_3828,N_681,N_1286);
nor U3829 (N_3829,N_1642,N_447);
nor U3830 (N_3830,N_665,N_2741);
or U3831 (N_3831,N_595,N_2792);
nor U3832 (N_3832,N_1526,N_465);
nor U3833 (N_3833,N_1781,N_5);
or U3834 (N_3834,N_935,N_627);
nand U3835 (N_3835,N_453,N_2213);
nand U3836 (N_3836,N_2572,N_2031);
nor U3837 (N_3837,N_1978,N_1922);
xor U3838 (N_3838,N_32,N_2500);
nor U3839 (N_3839,N_53,N_29);
or U3840 (N_3840,N_1291,N_1770);
and U3841 (N_3841,N_586,N_142);
nand U3842 (N_3842,N_719,N_2336);
nand U3843 (N_3843,N_1807,N_839);
xor U3844 (N_3844,N_2171,N_1628);
nor U3845 (N_3845,N_2489,N_1243);
and U3846 (N_3846,N_2958,N_197);
nand U3847 (N_3847,N_1163,N_123);
and U3848 (N_3848,N_1696,N_2954);
xor U3849 (N_3849,N_1732,N_571);
xor U3850 (N_3850,N_1457,N_1872);
or U3851 (N_3851,N_2998,N_512);
or U3852 (N_3852,N_774,N_2518);
or U3853 (N_3853,N_2036,N_1493);
and U3854 (N_3854,N_1214,N_539);
and U3855 (N_3855,N_1195,N_2039);
xor U3856 (N_3856,N_1946,N_2635);
nor U3857 (N_3857,N_1739,N_1008);
nand U3858 (N_3858,N_679,N_1258);
nor U3859 (N_3859,N_2609,N_178);
nor U3860 (N_3860,N_2424,N_1064);
nor U3861 (N_3861,N_379,N_2340);
and U3862 (N_3862,N_63,N_1120);
and U3863 (N_3863,N_2426,N_689);
nor U3864 (N_3864,N_686,N_1130);
nand U3865 (N_3865,N_1652,N_2209);
and U3866 (N_3866,N_215,N_2810);
nand U3867 (N_3867,N_2047,N_97);
or U3868 (N_3868,N_397,N_356);
nor U3869 (N_3869,N_1909,N_1915);
nand U3870 (N_3870,N_2494,N_1577);
and U3871 (N_3871,N_2820,N_1908);
xnor U3872 (N_3872,N_1110,N_1210);
or U3873 (N_3873,N_1140,N_2247);
nand U3874 (N_3874,N_2148,N_1950);
or U3875 (N_3875,N_1418,N_2282);
nor U3876 (N_3876,N_622,N_1011);
xor U3877 (N_3877,N_2360,N_1866);
and U3878 (N_3878,N_1238,N_1303);
xnor U3879 (N_3879,N_2318,N_2173);
or U3880 (N_3880,N_2694,N_2120);
or U3881 (N_3881,N_1861,N_1984);
xor U3882 (N_3882,N_2486,N_2134);
nand U3883 (N_3883,N_374,N_1034);
nor U3884 (N_3884,N_2833,N_90);
nor U3885 (N_3885,N_2839,N_2405);
nor U3886 (N_3886,N_2893,N_1030);
nand U3887 (N_3887,N_2928,N_1437);
nand U3888 (N_3888,N_409,N_2602);
xor U3889 (N_3889,N_2527,N_1102);
nand U3890 (N_3890,N_343,N_1752);
or U3891 (N_3891,N_2258,N_2994);
xnor U3892 (N_3892,N_1897,N_712);
and U3893 (N_3893,N_2237,N_2111);
nand U3894 (N_3894,N_1606,N_306);
nand U3895 (N_3895,N_2977,N_1749);
or U3896 (N_3896,N_64,N_2430);
nand U3897 (N_3897,N_2154,N_2507);
and U3898 (N_3898,N_2516,N_242);
xor U3899 (N_3899,N_2348,N_1837);
and U3900 (N_3900,N_490,N_1812);
xnor U3901 (N_3901,N_335,N_1310);
or U3902 (N_3902,N_1871,N_2376);
and U3903 (N_3903,N_2387,N_2763);
or U3904 (N_3904,N_709,N_2367);
nor U3905 (N_3905,N_2312,N_2221);
xnor U3906 (N_3906,N_1373,N_1474);
or U3907 (N_3907,N_647,N_1257);
nor U3908 (N_3908,N_2398,N_1820);
xnor U3909 (N_3909,N_1522,N_577);
and U3910 (N_3910,N_1673,N_1510);
nand U3911 (N_3911,N_1271,N_1901);
nand U3912 (N_3912,N_1198,N_2385);
nor U3913 (N_3913,N_1185,N_2185);
or U3914 (N_3914,N_1049,N_1777);
and U3915 (N_3915,N_635,N_2235);
or U3916 (N_3916,N_1649,N_1461);
xor U3917 (N_3917,N_1181,N_508);
or U3918 (N_3918,N_133,N_613);
and U3919 (N_3919,N_2627,N_1731);
nor U3920 (N_3920,N_14,N_2305);
nand U3921 (N_3921,N_205,N_1134);
and U3922 (N_3922,N_2143,N_2845);
and U3923 (N_3923,N_1000,N_554);
or U3924 (N_3924,N_163,N_358);
nand U3925 (N_3925,N_2915,N_1563);
nor U3926 (N_3926,N_654,N_2162);
nor U3927 (N_3927,N_2038,N_2126);
xor U3928 (N_3928,N_2444,N_1383);
nor U3929 (N_3929,N_1463,N_1980);
xor U3930 (N_3930,N_347,N_2196);
and U3931 (N_3931,N_2357,N_2284);
xnor U3932 (N_3932,N_1877,N_1170);
or U3933 (N_3933,N_514,N_550);
nor U3934 (N_3934,N_2442,N_2290);
nand U3935 (N_3935,N_422,N_1452);
nand U3936 (N_3936,N_1713,N_1236);
nand U3937 (N_3937,N_2138,N_1006);
xnor U3938 (N_3938,N_1987,N_1533);
nand U3939 (N_3939,N_787,N_2032);
or U3940 (N_3940,N_2775,N_615);
and U3941 (N_3941,N_1393,N_1733);
xnor U3942 (N_3942,N_2919,N_599);
and U3943 (N_3943,N_2962,N_1700);
nor U3944 (N_3944,N_1869,N_852);
nand U3945 (N_3945,N_2929,N_95);
xor U3946 (N_3946,N_406,N_2926);
nand U3947 (N_3947,N_741,N_1039);
nand U3948 (N_3948,N_1312,N_2437);
nand U3949 (N_3949,N_865,N_1178);
nor U3950 (N_3950,N_2767,N_750);
or U3951 (N_3951,N_352,N_805);
nand U3952 (N_3952,N_2045,N_292);
or U3953 (N_3953,N_2319,N_547);
nand U3954 (N_3954,N_2505,N_1737);
xnor U3955 (N_3955,N_175,N_1097);
nand U3956 (N_3956,N_2084,N_2647);
nand U3957 (N_3957,N_2867,N_746);
or U3958 (N_3958,N_146,N_1085);
nand U3959 (N_3959,N_12,N_923);
xor U3960 (N_3960,N_276,N_236);
nor U3961 (N_3961,N_168,N_2060);
and U3962 (N_3962,N_855,N_2589);
and U3963 (N_3963,N_2214,N_2890);
or U3964 (N_3964,N_722,N_49);
nand U3965 (N_3965,N_1639,N_2886);
or U3966 (N_3966,N_1728,N_870);
xor U3967 (N_3967,N_1137,N_1571);
and U3968 (N_3968,N_1495,N_2807);
nor U3969 (N_3969,N_375,N_1265);
xnor U3970 (N_3970,N_2000,N_2960);
and U3971 (N_3971,N_1999,N_821);
xnor U3972 (N_3972,N_766,N_1348);
nor U3973 (N_3973,N_2058,N_1823);
nor U3974 (N_3974,N_2170,N_22);
xor U3975 (N_3975,N_1104,N_431);
xnor U3976 (N_3976,N_9,N_2560);
and U3977 (N_3977,N_1302,N_425);
nor U3978 (N_3978,N_258,N_1840);
or U3979 (N_3979,N_1326,N_1436);
and U3980 (N_3980,N_1602,N_655);
and U3981 (N_3981,N_2762,N_1564);
nor U3982 (N_3982,N_2207,N_1021);
or U3983 (N_3983,N_2826,N_767);
or U3984 (N_3984,N_820,N_1190);
or U3985 (N_3985,N_964,N_2907);
and U3986 (N_3986,N_2862,N_2150);
or U3987 (N_3987,N_1785,N_104);
xnor U3988 (N_3988,N_761,N_1240);
xor U3989 (N_3989,N_1378,N_246);
and U3990 (N_3990,N_75,N_427);
or U3991 (N_3991,N_132,N_2184);
or U3992 (N_3992,N_618,N_858);
nor U3993 (N_3993,N_129,N_1760);
xnor U3994 (N_3994,N_2692,N_2099);
and U3995 (N_3995,N_2041,N_2019);
xnor U3996 (N_3996,N_2574,N_493);
nor U3997 (N_3997,N_1973,N_394);
xnor U3998 (N_3998,N_819,N_2969);
nand U3999 (N_3999,N_684,N_2838);
nor U4000 (N_4000,N_1384,N_1811);
and U4001 (N_4001,N_1370,N_585);
xnor U4002 (N_4002,N_2548,N_2074);
or U4003 (N_4003,N_2872,N_1565);
nor U4004 (N_4004,N_1142,N_1741);
or U4005 (N_4005,N_198,N_2651);
xor U4006 (N_4006,N_583,N_284);
xnor U4007 (N_4007,N_1473,N_2913);
nand U4008 (N_4008,N_1960,N_2327);
nand U4009 (N_4009,N_126,N_1605);
and U4010 (N_4010,N_2790,N_183);
xor U4011 (N_4011,N_1588,N_1878);
and U4012 (N_4012,N_2661,N_135);
nor U4013 (N_4013,N_1017,N_432);
nand U4014 (N_4014,N_1903,N_1179);
nor U4015 (N_4015,N_2941,N_2699);
nand U4016 (N_4016,N_1959,N_66);
or U4017 (N_4017,N_1371,N_255);
and U4018 (N_4018,N_2874,N_1891);
nand U4019 (N_4019,N_2300,N_1784);
nor U4020 (N_4020,N_1425,N_2570);
and U4021 (N_4021,N_1232,N_1566);
nor U4022 (N_4022,N_2822,N_1280);
and U4023 (N_4023,N_605,N_1993);
or U4024 (N_4024,N_589,N_2107);
and U4025 (N_4025,N_2577,N_2735);
xor U4026 (N_4026,N_128,N_2321);
nand U4027 (N_4027,N_105,N_652);
and U4028 (N_4028,N_1858,N_1410);
nand U4029 (N_4029,N_113,N_2759);
xnor U4030 (N_4030,N_1122,N_2070);
nor U4031 (N_4031,N_1414,N_2017);
xnor U4032 (N_4032,N_1358,N_2346);
nand U4033 (N_4033,N_1035,N_1538);
nand U4034 (N_4034,N_565,N_423);
nor U4035 (N_4035,N_403,N_2256);
nand U4036 (N_4036,N_2950,N_2643);
nor U4037 (N_4037,N_549,N_1768);
nor U4038 (N_4038,N_2517,N_342);
nor U4039 (N_4039,N_1743,N_568);
xnor U4040 (N_4040,N_2001,N_1892);
nand U4041 (N_4041,N_866,N_513);
nor U4042 (N_4042,N_1297,N_312);
nand U4043 (N_4043,N_2942,N_879);
nand U4044 (N_4044,N_960,N_1460);
or U4045 (N_4045,N_1724,N_2673);
xnor U4046 (N_4046,N_2722,N_981);
nand U4047 (N_4047,N_111,N_2004);
or U4048 (N_4048,N_2779,N_392);
xnor U4049 (N_4049,N_391,N_1695);
and U4050 (N_4050,N_2599,N_2266);
xnor U4051 (N_4051,N_2427,N_1063);
nand U4052 (N_4052,N_2562,N_1704);
xor U4053 (N_4053,N_1767,N_2180);
and U4054 (N_4054,N_2733,N_2483);
nand U4055 (N_4055,N_1500,N_1519);
nor U4056 (N_4056,N_2716,N_83);
nand U4057 (N_4057,N_2124,N_1759);
and U4058 (N_4058,N_1832,N_1012);
or U4059 (N_4059,N_2550,N_646);
or U4060 (N_4060,N_979,N_1143);
xnor U4061 (N_4061,N_2361,N_2033);
or U4062 (N_4062,N_2662,N_412);
or U4063 (N_4063,N_122,N_2037);
or U4064 (N_4064,N_846,N_1076);
xor U4065 (N_4065,N_350,N_396);
or U4066 (N_4066,N_1386,N_2693);
nor U4067 (N_4067,N_532,N_169);
nor U4068 (N_4068,N_1910,N_2097);
and U4069 (N_4069,N_2139,N_159);
nand U4070 (N_4070,N_1053,N_1188);
or U4071 (N_4071,N_1676,N_2497);
or U4072 (N_4072,N_1528,N_560);
nand U4073 (N_4073,N_213,N_2103);
or U4074 (N_4074,N_1025,N_521);
or U4075 (N_4075,N_416,N_2198);
nor U4076 (N_4076,N_965,N_2271);
or U4077 (N_4077,N_1161,N_814);
or U4078 (N_4078,N_1638,N_452);
nand U4079 (N_4079,N_2889,N_2861);
or U4080 (N_4080,N_1623,N_2372);
and U4081 (N_4081,N_991,N_200);
nand U4082 (N_4082,N_1799,N_1246);
or U4083 (N_4083,N_7,N_1419);
or U4084 (N_4084,N_1966,N_2026);
nand U4085 (N_4085,N_1668,N_810);
nand U4086 (N_4086,N_319,N_87);
nor U4087 (N_4087,N_1716,N_2754);
nand U4088 (N_4088,N_384,N_1299);
or U4089 (N_4089,N_2982,N_795);
xor U4090 (N_4090,N_2035,N_192);
nand U4091 (N_4091,N_261,N_842);
nor U4092 (N_4092,N_1991,N_440);
xnor U4093 (N_4093,N_2193,N_2298);
nand U4094 (N_4094,N_1794,N_1680);
nand U4095 (N_4095,N_1756,N_1542);
nor U4096 (N_4096,N_2347,N_509);
or U4097 (N_4097,N_1985,N_296);
xor U4098 (N_4098,N_2538,N_1970);
nor U4099 (N_4099,N_2930,N_1197);
nor U4100 (N_4100,N_1936,N_944);
xor U4101 (N_4101,N_641,N_1846);
nand U4102 (N_4102,N_900,N_786);
xor U4103 (N_4103,N_919,N_1578);
nor U4104 (N_4104,N_1679,N_1293);
nand U4105 (N_4105,N_1055,N_1364);
nand U4106 (N_4106,N_502,N_1092);
and U4107 (N_4107,N_1413,N_1969);
xnor U4108 (N_4108,N_1883,N_1125);
or U4109 (N_4109,N_1850,N_1586);
or U4110 (N_4110,N_1253,N_2102);
nor U4111 (N_4111,N_934,N_1475);
and U4112 (N_4112,N_1315,N_62);
or U4113 (N_4113,N_2493,N_2501);
nor U4114 (N_4114,N_2112,N_947);
nand U4115 (N_4115,N_1266,N_248);
nor U4116 (N_4116,N_2963,N_1907);
nand U4117 (N_4117,N_415,N_1024);
nor U4118 (N_4118,N_2542,N_1465);
nor U4119 (N_4119,N_1450,N_1213);
nor U4120 (N_4120,N_581,N_1285);
and U4121 (N_4121,N_1798,N_193);
xor U4122 (N_4122,N_1176,N_1975);
xor U4123 (N_4123,N_2414,N_2968);
or U4124 (N_4124,N_1255,N_1736);
and U4125 (N_4125,N_1311,N_1559);
or U4126 (N_4126,N_322,N_1368);
nor U4127 (N_4127,N_763,N_1149);
and U4128 (N_4128,N_2393,N_2409);
xnor U4129 (N_4129,N_2454,N_2967);
or U4130 (N_4130,N_148,N_1075);
nor U4131 (N_4131,N_2566,N_2863);
xnor U4132 (N_4132,N_1094,N_2429);
nor U4133 (N_4133,N_1467,N_1150);
xor U4134 (N_4134,N_476,N_1620);
xor U4135 (N_4135,N_145,N_1635);
nand U4136 (N_4136,N_1349,N_417);
nand U4137 (N_4137,N_1175,N_1691);
xor U4138 (N_4138,N_2755,N_2588);
nand U4139 (N_4139,N_1653,N_2286);
or U4140 (N_4140,N_1824,N_1647);
nand U4141 (N_4141,N_788,N_2188);
xnor U4142 (N_4142,N_2629,N_44);
or U4143 (N_4143,N_802,N_2739);
nand U4144 (N_4144,N_2817,N_933);
nand U4145 (N_4145,N_1405,N_2034);
nor U4146 (N_4146,N_1338,N_2805);
nand U4147 (N_4147,N_716,N_2106);
and U4148 (N_4148,N_2226,N_1884);
nor U4149 (N_4149,N_1503,N_96);
xor U4150 (N_4150,N_637,N_1328);
xnor U4151 (N_4151,N_370,N_1796);
xor U4152 (N_4152,N_160,N_2317);
nor U4153 (N_4153,N_672,N_1107);
and U4154 (N_4154,N_1183,N_241);
and U4155 (N_4155,N_2601,N_559);
nor U4156 (N_4156,N_1589,N_1079);
xor U4157 (N_4157,N_2006,N_638);
or U4158 (N_4158,N_2016,N_279);
nor U4159 (N_4159,N_1712,N_593);
nor U4160 (N_4160,N_742,N_2610);
nor U4161 (N_4161,N_2819,N_1318);
and U4162 (N_4162,N_2947,N_516);
or U4163 (N_4163,N_968,N_980);
nand U4164 (N_4164,N_286,N_925);
nor U4165 (N_4165,N_2664,N_1027);
and U4166 (N_4166,N_1548,N_2211);
xor U4167 (N_4167,N_781,N_225);
or U4168 (N_4168,N_2985,N_1806);
or U4169 (N_4169,N_1771,N_2728);
nor U4170 (N_4170,N_1462,N_894);
xnor U4171 (N_4171,N_2777,N_351);
xor U4172 (N_4172,N_1158,N_2334);
or U4173 (N_4173,N_161,N_2311);
or U4174 (N_4174,N_340,N_1305);
and U4175 (N_4175,N_575,N_1992);
and U4176 (N_4176,N_1845,N_752);
and U4177 (N_4177,N_333,N_2922);
xnor U4178 (N_4178,N_1083,N_278);
nor U4179 (N_4179,N_505,N_430);
or U4180 (N_4180,N_657,N_2578);
nor U4181 (N_4181,N_2177,N_2793);
nor U4182 (N_4182,N_2607,N_1219);
nand U4183 (N_4183,N_1711,N_675);
and U4184 (N_4184,N_807,N_1687);
nor U4185 (N_4185,N_2975,N_2181);
nor U4186 (N_4186,N_1583,N_570);
nand U4187 (N_4187,N_2868,N_1477);
or U4188 (N_4188,N_482,N_617);
and U4189 (N_4189,N_1515,N_1061);
nor U4190 (N_4190,N_445,N_1316);
xor U4191 (N_4191,N_2008,N_835);
nor U4192 (N_4192,N_2976,N_367);
xnor U4193 (N_4193,N_1581,N_1517);
xnor U4194 (N_4194,N_119,N_895);
or U4195 (N_4195,N_2166,N_706);
nand U4196 (N_4196,N_2476,N_1404);
or U4197 (N_4197,N_2525,N_1416);
and U4198 (N_4198,N_653,N_678);
xnor U4199 (N_4199,N_2988,N_785);
xor U4200 (N_4200,N_223,N_466);
and U4201 (N_4201,N_2959,N_1221);
or U4202 (N_4202,N_293,N_2757);
nand U4203 (N_4203,N_238,N_1507);
and U4204 (N_4204,N_316,N_667);
or U4205 (N_4205,N_2069,N_326);
nor U4206 (N_4206,N_1610,N_314);
or U4207 (N_4207,N_2600,N_61);
or U4208 (N_4208,N_1231,N_59);
or U4209 (N_4209,N_2104,N_612);
and U4210 (N_4210,N_130,N_1934);
and U4211 (N_4211,N_628,N_1336);
nor U4212 (N_4212,N_2687,N_2114);
nor U4213 (N_4213,N_2675,N_952);
nand U4214 (N_4214,N_2370,N_2765);
and U4215 (N_4215,N_2172,N_2468);
nor U4216 (N_4216,N_151,N_1763);
nor U4217 (N_4217,N_2670,N_844);
nor U4218 (N_4218,N_1778,N_2197);
nor U4219 (N_4219,N_1479,N_753);
nor U4220 (N_4220,N_2053,N_1939);
xor U4221 (N_4221,N_2827,N_2952);
xor U4222 (N_4222,N_1833,N_481);
nor U4223 (N_4223,N_1481,N_1322);
nand U4224 (N_4224,N_1809,N_25);
or U4225 (N_4225,N_1839,N_2328);
nand U4226 (N_4226,N_848,N_442);
and U4227 (N_4227,N_1576,N_1665);
nand U4228 (N_4228,N_1356,N_120);
xnor U4229 (N_4229,N_2350,N_1382);
or U4230 (N_4230,N_2520,N_510);
nand U4231 (N_4231,N_2880,N_2029);
and U4232 (N_4232,N_328,N_1282);
nand U4233 (N_4233,N_2721,N_2301);
xnor U4234 (N_4234,N_2974,N_2503);
xor U4235 (N_4235,N_251,N_1440);
xor U4236 (N_4236,N_881,N_2603);
and U4237 (N_4237,N_2345,N_448);
xor U4238 (N_4238,N_1621,N_2127);
and U4239 (N_4239,N_1112,N_82);
or U4240 (N_4240,N_496,N_893);
nor U4241 (N_4241,N_2105,N_1496);
nor U4242 (N_4242,N_1321,N_332);
or U4243 (N_4243,N_972,N_2141);
xnor U4244 (N_4244,N_985,N_885);
and U4245 (N_4245,N_1132,N_475);
nor U4246 (N_4246,N_2624,N_1424);
or U4247 (N_4247,N_859,N_93);
nand U4248 (N_4248,N_896,N_2668);
nand U4249 (N_4249,N_2646,N_927);
and U4250 (N_4250,N_2343,N_1051);
nor U4251 (N_4251,N_929,N_2581);
and U4252 (N_4252,N_1218,N_2875);
and U4253 (N_4253,N_478,N_2813);
or U4254 (N_4254,N_1734,N_1822);
and U4255 (N_4255,N_1913,N_2259);
nor U4256 (N_4256,N_1331,N_1041);
xor U4257 (N_4257,N_2178,N_2088);
nand U4258 (N_4258,N_694,N_2658);
nand U4259 (N_4259,N_2896,N_2049);
nand U4260 (N_4260,N_1268,N_2846);
nor U4261 (N_4261,N_355,N_2945);
xnor U4262 (N_4262,N_2535,N_1544);
xor U4263 (N_4263,N_202,N_2508);
nor U4264 (N_4264,N_2461,N_1434);
and U4265 (N_4265,N_747,N_439);
xor U4266 (N_4266,N_2066,N_1965);
nand U4267 (N_4267,N_735,N_2681);
nor U4268 (N_4268,N_85,N_2703);
and U4269 (N_4269,N_1631,N_645);
or U4270 (N_4270,N_1196,N_2816);
xor U4271 (N_4271,N_1399,N_887);
or U4272 (N_4272,N_1117,N_1272);
nand U4273 (N_4273,N_2858,N_765);
or U4274 (N_4274,N_2100,N_2117);
and U4275 (N_4275,N_809,N_294);
xor U4276 (N_4276,N_2853,N_484);
or U4277 (N_4277,N_1764,N_2411);
nor U4278 (N_4278,N_803,N_2090);
nor U4279 (N_4279,N_721,N_1212);
nor U4280 (N_4280,N_174,N_561);
xor U4281 (N_4281,N_643,N_1480);
and U4282 (N_4282,N_1951,N_72);
nand U4283 (N_4283,N_556,N_1390);
xnor U4284 (N_4284,N_2989,N_60);
or U4285 (N_4285,N_1439,N_715);
or U4286 (N_4286,N_975,N_1896);
and U4287 (N_4287,N_2048,N_1022);
or U4288 (N_4288,N_590,N_573);
or U4289 (N_4289,N_494,N_2463);
nor U4290 (N_4290,N_1916,N_2789);
and U4291 (N_4291,N_1340,N_1661);
nor U4292 (N_4292,N_1681,N_2971);
xor U4293 (N_4293,N_2720,N_67);
and U4294 (N_4294,N_808,N_2371);
nand U4295 (N_4295,N_2396,N_2768);
nor U4296 (N_4296,N_2743,N_995);
or U4297 (N_4297,N_2996,N_1887);
xor U4298 (N_4298,N_2390,N_682);
or U4299 (N_4299,N_1703,N_2676);
and U4300 (N_4300,N_1873,N_2297);
or U4301 (N_4301,N_2534,N_517);
nand U4302 (N_4302,N_903,N_1932);
and U4303 (N_4303,N_2142,N_2732);
or U4304 (N_4304,N_2275,N_2464);
or U4305 (N_4305,N_457,N_1893);
nand U4306 (N_4306,N_1327,N_254);
nor U4307 (N_4307,N_230,N_2986);
nor U4308 (N_4308,N_2528,N_1381);
xnor U4309 (N_4309,N_1802,N_792);
and U4310 (N_4310,N_2477,N_833);
or U4311 (N_4311,N_1568,N_1435);
nor U4312 (N_4312,N_2366,N_50);
xnor U4313 (N_4313,N_1882,N_2617);
or U4314 (N_4314,N_2176,N_217);
xor U4315 (N_4315,N_444,N_1933);
xnor U4316 (N_4316,N_2291,N_2413);
and U4317 (N_4317,N_497,N_1423);
or U4318 (N_4318,N_955,N_951);
nand U4319 (N_4319,N_1346,N_2802);
nor U4320 (N_4320,N_407,N_2526);
or U4321 (N_4321,N_1116,N_2216);
nand U4322 (N_4322,N_211,N_850);
nor U4323 (N_4323,N_345,N_2587);
or U4324 (N_4324,N_1580,N_1742);
or U4325 (N_4325,N_2419,N_2537);
or U4326 (N_4326,N_2264,N_566);
nand U4327 (N_4327,N_2955,N_1683);
xnor U4328 (N_4328,N_1147,N_140);
or U4329 (N_4329,N_443,N_2791);
or U4330 (N_4330,N_1598,N_737);
and U4331 (N_4331,N_2356,N_1604);
or U4332 (N_4332,N_670,N_2219);
xor U4333 (N_4333,N_1032,N_155);
or U4334 (N_4334,N_2339,N_2808);
and U4335 (N_4335,N_2795,N_1644);
nor U4336 (N_4336,N_324,N_2706);
nor U4337 (N_4337,N_1412,N_2441);
nand U4338 (N_4338,N_1153,N_744);
nor U4339 (N_4339,N_770,N_1451);
or U4340 (N_4340,N_2606,N_2281);
and U4341 (N_4341,N_1466,N_73);
xnor U4342 (N_4342,N_669,N_1868);
or U4343 (N_4343,N_196,N_1943);
and U4344 (N_4344,N_909,N_24);
nor U4345 (N_4345,N_990,N_697);
and U4346 (N_4346,N_1062,N_2715);
nand U4347 (N_4347,N_2251,N_2983);
nand U4348 (N_4348,N_2189,N_1826);
and U4349 (N_4349,N_1797,N_1792);
xor U4350 (N_4350,N_1783,N_1974);
nor U4351 (N_4351,N_522,N_1774);
nand U4352 (N_4352,N_2663,N_1663);
nand U4353 (N_4353,N_336,N_459);
nand U4354 (N_4354,N_869,N_400);
nand U4355 (N_4355,N_2158,N_1247);
nor U4356 (N_4356,N_2014,N_987);
nor U4357 (N_4357,N_1166,N_992);
and U4358 (N_4358,N_1320,N_381);
or U4359 (N_4359,N_283,N_153);
nand U4360 (N_4360,N_880,N_949);
and U4361 (N_4361,N_1270,N_55);
nor U4362 (N_4362,N_166,N_395);
or U4363 (N_4363,N_1702,N_1674);
nor U4364 (N_4364,N_726,N_1447);
nor U4365 (N_4365,N_756,N_685);
and U4366 (N_4366,N_2456,N_867);
or U4367 (N_4367,N_1226,N_2187);
nor U4368 (N_4368,N_2843,N_1512);
xnor U4369 (N_4369,N_1553,N_28);
nor U4370 (N_4370,N_631,N_216);
and U4371 (N_4371,N_574,N_2392);
or U4372 (N_4372,N_2407,N_420);
xor U4373 (N_4373,N_1722,N_2631);
or U4374 (N_4374,N_488,N_1202);
xnor U4375 (N_4375,N_303,N_2080);
and U4376 (N_4376,N_854,N_2428);
or U4377 (N_4377,N_930,N_1643);
or U4378 (N_4378,N_2135,N_2043);
nand U4379 (N_4379,N_2684,N_1469);
nand U4380 (N_4380,N_2160,N_624);
or U4381 (N_4381,N_1862,N_2263);
or U4382 (N_4382,N_580,N_2920);
nand U4383 (N_4383,N_2051,N_768);
xnor U4384 (N_4384,N_704,N_940);
nand U4385 (N_4385,N_2731,N_1968);
xor U4386 (N_4386,N_736,N_2313);
or U4387 (N_4387,N_461,N_2522);
and U4388 (N_4388,N_1369,N_1241);
nand U4389 (N_4389,N_46,N_1505);
or U4390 (N_4390,N_2459,N_6);
xor U4391 (N_4391,N_578,N_2840);
and U4392 (N_4392,N_2028,N_346);
xor U4393 (N_4393,N_1106,N_2239);
xor U4394 (N_4394,N_2529,N_534);
xnor U4395 (N_4395,N_813,N_2065);
nor U4396 (N_4396,N_2672,N_2614);
nor U4397 (N_4397,N_2973,N_1281);
nand U4398 (N_4398,N_310,N_2626);
xnor U4399 (N_4399,N_2506,N_2667);
nor U4400 (N_4400,N_1859,N_86);
or U4401 (N_4401,N_2637,N_334);
xor U4402 (N_4402,N_2934,N_1254);
or U4403 (N_4403,N_1347,N_1154);
xor U4404 (N_4404,N_1073,N_2190);
nand U4405 (N_4405,N_1740,N_1324);
and U4406 (N_4406,N_2815,N_125);
or U4407 (N_4407,N_1729,N_1162);
xnor U4408 (N_4408,N_1141,N_555);
nor U4409 (N_4409,N_2169,N_898);
xnor U4410 (N_4410,N_289,N_2965);
or U4411 (N_4411,N_69,N_300);
nor U4412 (N_4412,N_171,N_2579);
nor U4413 (N_4413,N_1453,N_1050);
and U4414 (N_4414,N_1976,N_2389);
or U4415 (N_4415,N_875,N_673);
nor U4416 (N_4416,N_2418,N_730);
xor U4417 (N_4417,N_1609,N_34);
xor U4418 (N_4418,N_1834,N_2183);
and U4419 (N_4419,N_38,N_1748);
xnor U4420 (N_4420,N_158,N_1359);
nand U4421 (N_4421,N_743,N_1552);
nand U4422 (N_4422,N_2540,N_2490);
xor U4423 (N_4423,N_2850,N_1078);
xnor U4424 (N_4424,N_760,N_1710);
nand U4425 (N_4425,N_2469,N_993);
nand U4426 (N_4426,N_2250,N_553);
and U4427 (N_4427,N_2174,N_2119);
nand U4428 (N_4428,N_1864,N_219);
xnor U4429 (N_4429,N_1958,N_127);
nand U4430 (N_4430,N_2445,N_474);
or U4431 (N_4431,N_2678,N_441);
nand U4432 (N_4432,N_1123,N_1746);
xor U4433 (N_4433,N_1717,N_262);
nor U4434 (N_4434,N_2496,N_2533);
or U4435 (N_4435,N_1549,N_2979);
xor U4436 (N_4436,N_2608,N_966);
and U4437 (N_4437,N_636,N_906);
nand U4438 (N_4438,N_2831,N_2785);
and U4439 (N_4439,N_224,N_1098);
nand U4440 (N_4440,N_206,N_1818);
nand U4441 (N_4441,N_2086,N_2723);
or U4442 (N_4442,N_1940,N_2248);
xor U4443 (N_4443,N_777,N_2595);
or U4444 (N_4444,N_1630,N_2377);
nor U4445 (N_4445,N_2559,N_1182);
and U4446 (N_4446,N_2852,N_1114);
xor U4447 (N_4447,N_1556,N_54);
xnor U4448 (N_4448,N_525,N_1224);
and U4449 (N_4449,N_2997,N_1914);
nand U4450 (N_4450,N_2521,N_1004);
and U4451 (N_4451,N_831,N_2558);
nand U4452 (N_4452,N_1546,N_941);
nand U4453 (N_4453,N_1483,N_2909);
nand U4454 (N_4454,N_1788,N_890);
or U4455 (N_4455,N_100,N_2702);
and U4456 (N_4456,N_2887,N_1911);
xnor U4457 (N_4457,N_592,N_1018);
nand U4458 (N_4458,N_2087,N_468);
nand U4459 (N_4459,N_1539,N_2580);
nand U4460 (N_4460,N_759,N_2288);
xor U4461 (N_4461,N_2191,N_485);
nor U4462 (N_4462,N_1874,N_1173);
nand U4463 (N_4463,N_2267,N_2306);
or U4464 (N_4464,N_913,N_2888);
xor U4465 (N_4465,N_714,N_297);
xor U4466 (N_4466,N_472,N_2421);
or U4467 (N_4467,N_2957,N_1470);
nor U4468 (N_4468,N_377,N_2487);
xor U4469 (N_4469,N_1730,N_42);
and U4470 (N_4470,N_2325,N_519);
or U4471 (N_4471,N_1135,N_2801);
nand U4472 (N_4472,N_1963,N_1930);
xnor U4473 (N_4473,N_2632,N_1912);
or U4474 (N_4474,N_1264,N_2140);
nand U4475 (N_4475,N_1244,N_998);
nor U4476 (N_4476,N_152,N_1962);
xor U4477 (N_4477,N_1108,N_2898);
and U4478 (N_4478,N_827,N_2511);
xnor U4479 (N_4479,N_2125,N_1689);
nor U4480 (N_4480,N_2729,N_2438);
nand U4481 (N_4481,N_2408,N_691);
xor U4482 (N_4482,N_832,N_1972);
or U4483 (N_4483,N_1207,N_1692);
or U4484 (N_4484,N_1956,N_2758);
nand U4485 (N_4485,N_1421,N_1133);
or U4486 (N_4486,N_2179,N_2109);
nor U4487 (N_4487,N_1953,N_1354);
xnor U4488 (N_4488,N_1738,N_2354);
and U4489 (N_4489,N_733,N_1136);
nor U4490 (N_4490,N_2923,N_2622);
nand U4491 (N_4491,N_2778,N_2991);
nand U4492 (N_4492,N_1184,N_1961);
nand U4493 (N_4493,N_1981,N_937);
nand U4494 (N_4494,N_1931,N_1339);
xnor U4495 (N_4495,N_545,N_1082);
xor U4496 (N_4496,N_2283,N_2870);
and U4497 (N_4497,N_2349,N_1529);
nand U4498 (N_4498,N_2018,N_436);
xor U4499 (N_4499,N_31,N_2797);
and U4500 (N_4500,N_1342,N_1214);
and U4501 (N_4501,N_678,N_1454);
nand U4502 (N_4502,N_2166,N_1761);
and U4503 (N_4503,N_2016,N_2442);
nor U4504 (N_4504,N_520,N_2266);
nand U4505 (N_4505,N_2402,N_1280);
nand U4506 (N_4506,N_1681,N_489);
or U4507 (N_4507,N_384,N_2464);
and U4508 (N_4508,N_849,N_87);
or U4509 (N_4509,N_2194,N_1830);
xor U4510 (N_4510,N_212,N_2527);
nor U4511 (N_4511,N_240,N_2649);
nor U4512 (N_4512,N_2977,N_2949);
nand U4513 (N_4513,N_119,N_2794);
or U4514 (N_4514,N_2141,N_1250);
or U4515 (N_4515,N_1817,N_2199);
or U4516 (N_4516,N_2703,N_2461);
or U4517 (N_4517,N_1119,N_2293);
and U4518 (N_4518,N_193,N_1204);
nand U4519 (N_4519,N_780,N_310);
nand U4520 (N_4520,N_1949,N_133);
or U4521 (N_4521,N_755,N_1320);
or U4522 (N_4522,N_1361,N_2302);
or U4523 (N_4523,N_2208,N_2652);
or U4524 (N_4524,N_1615,N_663);
xnor U4525 (N_4525,N_207,N_2356);
nand U4526 (N_4526,N_2688,N_1364);
nor U4527 (N_4527,N_162,N_2051);
xor U4528 (N_4528,N_2767,N_512);
nor U4529 (N_4529,N_758,N_115);
and U4530 (N_4530,N_1161,N_434);
nor U4531 (N_4531,N_2962,N_2463);
and U4532 (N_4532,N_1919,N_203);
nand U4533 (N_4533,N_1706,N_274);
nand U4534 (N_4534,N_1000,N_591);
and U4535 (N_4535,N_2097,N_770);
nand U4536 (N_4536,N_817,N_1826);
xnor U4537 (N_4537,N_132,N_2308);
nand U4538 (N_4538,N_413,N_61);
or U4539 (N_4539,N_232,N_2320);
nand U4540 (N_4540,N_342,N_2624);
and U4541 (N_4541,N_147,N_789);
nor U4542 (N_4542,N_134,N_2340);
nor U4543 (N_4543,N_1484,N_836);
nor U4544 (N_4544,N_1244,N_2509);
nor U4545 (N_4545,N_1802,N_106);
xor U4546 (N_4546,N_321,N_495);
and U4547 (N_4547,N_1489,N_1876);
nor U4548 (N_4548,N_2187,N_2708);
nor U4549 (N_4549,N_874,N_2648);
nand U4550 (N_4550,N_1937,N_384);
nor U4551 (N_4551,N_2058,N_1312);
nand U4552 (N_4552,N_2054,N_2057);
and U4553 (N_4553,N_1058,N_1422);
or U4554 (N_4554,N_1989,N_2946);
xor U4555 (N_4555,N_1555,N_1543);
xnor U4556 (N_4556,N_277,N_2042);
nand U4557 (N_4557,N_1950,N_812);
xor U4558 (N_4558,N_2398,N_1135);
or U4559 (N_4559,N_2984,N_2459);
nand U4560 (N_4560,N_300,N_2939);
and U4561 (N_4561,N_1488,N_2455);
or U4562 (N_4562,N_1864,N_1163);
nor U4563 (N_4563,N_910,N_1707);
nor U4564 (N_4564,N_2928,N_108);
nor U4565 (N_4565,N_800,N_1855);
nand U4566 (N_4566,N_2046,N_1865);
or U4567 (N_4567,N_864,N_1622);
or U4568 (N_4568,N_2100,N_2718);
xnor U4569 (N_4569,N_1030,N_355);
xnor U4570 (N_4570,N_2815,N_1619);
and U4571 (N_4571,N_526,N_301);
xnor U4572 (N_4572,N_534,N_136);
and U4573 (N_4573,N_2868,N_2927);
xnor U4574 (N_4574,N_2585,N_1091);
or U4575 (N_4575,N_703,N_2330);
nor U4576 (N_4576,N_57,N_468);
nand U4577 (N_4577,N_2503,N_1973);
and U4578 (N_4578,N_2263,N_1426);
xnor U4579 (N_4579,N_1154,N_2513);
or U4580 (N_4580,N_1886,N_2920);
or U4581 (N_4581,N_811,N_1842);
nor U4582 (N_4582,N_1464,N_906);
and U4583 (N_4583,N_61,N_1139);
nand U4584 (N_4584,N_767,N_2580);
nand U4585 (N_4585,N_120,N_2828);
and U4586 (N_4586,N_2077,N_1446);
and U4587 (N_4587,N_564,N_2504);
nand U4588 (N_4588,N_2570,N_2765);
and U4589 (N_4589,N_1668,N_1803);
or U4590 (N_4590,N_9,N_2378);
and U4591 (N_4591,N_1851,N_2718);
nand U4592 (N_4592,N_544,N_64);
nor U4593 (N_4593,N_1414,N_1131);
nor U4594 (N_4594,N_2625,N_2865);
nand U4595 (N_4595,N_2288,N_2110);
and U4596 (N_4596,N_1681,N_1270);
nor U4597 (N_4597,N_36,N_308);
or U4598 (N_4598,N_1436,N_2244);
and U4599 (N_4599,N_1468,N_1315);
or U4600 (N_4600,N_2454,N_865);
and U4601 (N_4601,N_683,N_1396);
xor U4602 (N_4602,N_1283,N_847);
and U4603 (N_4603,N_1231,N_2404);
xor U4604 (N_4604,N_2640,N_372);
nor U4605 (N_4605,N_2160,N_93);
or U4606 (N_4606,N_633,N_674);
nor U4607 (N_4607,N_524,N_2273);
nor U4608 (N_4608,N_2833,N_1928);
or U4609 (N_4609,N_53,N_1017);
nand U4610 (N_4610,N_174,N_1446);
xnor U4611 (N_4611,N_2898,N_2666);
xnor U4612 (N_4612,N_1294,N_2727);
nor U4613 (N_4613,N_2776,N_299);
nor U4614 (N_4614,N_1370,N_328);
and U4615 (N_4615,N_2872,N_572);
and U4616 (N_4616,N_804,N_674);
or U4617 (N_4617,N_2255,N_1557);
nand U4618 (N_4618,N_2400,N_783);
or U4619 (N_4619,N_1027,N_1113);
nand U4620 (N_4620,N_1738,N_2466);
nor U4621 (N_4621,N_2116,N_2502);
and U4622 (N_4622,N_1950,N_1170);
or U4623 (N_4623,N_2537,N_1427);
xor U4624 (N_4624,N_540,N_2232);
and U4625 (N_4625,N_1241,N_198);
or U4626 (N_4626,N_2129,N_2081);
or U4627 (N_4627,N_1664,N_2984);
nand U4628 (N_4628,N_285,N_2810);
and U4629 (N_4629,N_2794,N_914);
nor U4630 (N_4630,N_1555,N_173);
xor U4631 (N_4631,N_2757,N_1772);
xnor U4632 (N_4632,N_390,N_1885);
nand U4633 (N_4633,N_677,N_1430);
nand U4634 (N_4634,N_1159,N_2812);
and U4635 (N_4635,N_1118,N_668);
and U4636 (N_4636,N_1924,N_2213);
or U4637 (N_4637,N_1157,N_1473);
nand U4638 (N_4638,N_2725,N_375);
and U4639 (N_4639,N_2907,N_1606);
and U4640 (N_4640,N_418,N_1570);
and U4641 (N_4641,N_1245,N_622);
xor U4642 (N_4642,N_1305,N_2921);
nor U4643 (N_4643,N_145,N_485);
and U4644 (N_4644,N_1206,N_1823);
and U4645 (N_4645,N_2289,N_685);
nor U4646 (N_4646,N_1009,N_2765);
and U4647 (N_4647,N_1509,N_409);
nor U4648 (N_4648,N_1864,N_1965);
or U4649 (N_4649,N_2222,N_1935);
nand U4650 (N_4650,N_527,N_2105);
xor U4651 (N_4651,N_2745,N_275);
and U4652 (N_4652,N_1578,N_1715);
xor U4653 (N_4653,N_1640,N_748);
nor U4654 (N_4654,N_351,N_87);
or U4655 (N_4655,N_2071,N_993);
nand U4656 (N_4656,N_942,N_2600);
nand U4657 (N_4657,N_1831,N_1295);
and U4658 (N_4658,N_731,N_2302);
xor U4659 (N_4659,N_1976,N_2030);
xor U4660 (N_4660,N_2148,N_2741);
or U4661 (N_4661,N_873,N_280);
nor U4662 (N_4662,N_545,N_2719);
and U4663 (N_4663,N_2752,N_1474);
nand U4664 (N_4664,N_1349,N_429);
nor U4665 (N_4665,N_216,N_1791);
xor U4666 (N_4666,N_1599,N_1755);
nor U4667 (N_4667,N_2657,N_2414);
nor U4668 (N_4668,N_309,N_360);
xor U4669 (N_4669,N_2868,N_625);
xor U4670 (N_4670,N_1145,N_747);
nor U4671 (N_4671,N_2339,N_71);
or U4672 (N_4672,N_59,N_2038);
nand U4673 (N_4673,N_1660,N_943);
and U4674 (N_4674,N_1710,N_2762);
and U4675 (N_4675,N_1079,N_961);
nand U4676 (N_4676,N_1921,N_2424);
and U4677 (N_4677,N_1449,N_2026);
nand U4678 (N_4678,N_2772,N_293);
nand U4679 (N_4679,N_325,N_2377);
nand U4680 (N_4680,N_804,N_1744);
nand U4681 (N_4681,N_2027,N_1270);
nor U4682 (N_4682,N_2330,N_2480);
nand U4683 (N_4683,N_1493,N_2295);
and U4684 (N_4684,N_1324,N_593);
and U4685 (N_4685,N_2914,N_2567);
or U4686 (N_4686,N_2449,N_1184);
and U4687 (N_4687,N_2580,N_479);
and U4688 (N_4688,N_2452,N_88);
nand U4689 (N_4689,N_2749,N_2786);
or U4690 (N_4690,N_400,N_1469);
xnor U4691 (N_4691,N_1279,N_181);
or U4692 (N_4692,N_1849,N_1830);
nand U4693 (N_4693,N_588,N_2912);
and U4694 (N_4694,N_1598,N_2203);
xnor U4695 (N_4695,N_1894,N_23);
nand U4696 (N_4696,N_2690,N_1395);
nor U4697 (N_4697,N_2366,N_2606);
nand U4698 (N_4698,N_2973,N_1982);
and U4699 (N_4699,N_669,N_2805);
and U4700 (N_4700,N_2379,N_1999);
nor U4701 (N_4701,N_1204,N_1816);
nand U4702 (N_4702,N_1597,N_355);
nand U4703 (N_4703,N_1929,N_317);
xor U4704 (N_4704,N_2428,N_967);
xnor U4705 (N_4705,N_1982,N_1696);
and U4706 (N_4706,N_34,N_208);
or U4707 (N_4707,N_2984,N_644);
or U4708 (N_4708,N_669,N_719);
nor U4709 (N_4709,N_2522,N_906);
nor U4710 (N_4710,N_1106,N_1916);
and U4711 (N_4711,N_940,N_2214);
xor U4712 (N_4712,N_2025,N_302);
nand U4713 (N_4713,N_209,N_2877);
nand U4714 (N_4714,N_1797,N_1988);
nor U4715 (N_4715,N_1783,N_6);
and U4716 (N_4716,N_402,N_1086);
or U4717 (N_4717,N_1044,N_1946);
nand U4718 (N_4718,N_2297,N_2173);
nand U4719 (N_4719,N_2680,N_2398);
or U4720 (N_4720,N_2846,N_2265);
nand U4721 (N_4721,N_2585,N_875);
nand U4722 (N_4722,N_2618,N_221);
or U4723 (N_4723,N_1949,N_1132);
and U4724 (N_4724,N_296,N_2198);
and U4725 (N_4725,N_591,N_1984);
nand U4726 (N_4726,N_1992,N_544);
nand U4727 (N_4727,N_2608,N_2032);
nor U4728 (N_4728,N_270,N_535);
or U4729 (N_4729,N_1161,N_2371);
nor U4730 (N_4730,N_2791,N_1767);
nor U4731 (N_4731,N_66,N_2155);
and U4732 (N_4732,N_2642,N_431);
nor U4733 (N_4733,N_1269,N_1958);
and U4734 (N_4734,N_561,N_57);
nand U4735 (N_4735,N_1534,N_257);
nand U4736 (N_4736,N_2448,N_2171);
nor U4737 (N_4737,N_857,N_1719);
or U4738 (N_4738,N_467,N_2089);
or U4739 (N_4739,N_2925,N_292);
and U4740 (N_4740,N_2389,N_5);
and U4741 (N_4741,N_2969,N_1292);
or U4742 (N_4742,N_2777,N_1833);
xnor U4743 (N_4743,N_333,N_662);
or U4744 (N_4744,N_500,N_2863);
or U4745 (N_4745,N_2029,N_131);
and U4746 (N_4746,N_758,N_1561);
or U4747 (N_4747,N_93,N_47);
xor U4748 (N_4748,N_419,N_381);
or U4749 (N_4749,N_1495,N_2213);
nand U4750 (N_4750,N_1345,N_1175);
xor U4751 (N_4751,N_1518,N_401);
nor U4752 (N_4752,N_254,N_1169);
xor U4753 (N_4753,N_86,N_2468);
xnor U4754 (N_4754,N_2077,N_1179);
nor U4755 (N_4755,N_960,N_1772);
and U4756 (N_4756,N_1373,N_1408);
or U4757 (N_4757,N_1172,N_2384);
and U4758 (N_4758,N_903,N_832);
xnor U4759 (N_4759,N_1208,N_922);
nand U4760 (N_4760,N_1840,N_47);
nor U4761 (N_4761,N_1760,N_2764);
nor U4762 (N_4762,N_2485,N_902);
xnor U4763 (N_4763,N_406,N_2490);
nand U4764 (N_4764,N_810,N_1767);
nor U4765 (N_4765,N_2992,N_1891);
or U4766 (N_4766,N_2726,N_2201);
nor U4767 (N_4767,N_768,N_1995);
or U4768 (N_4768,N_802,N_2631);
and U4769 (N_4769,N_1276,N_289);
and U4770 (N_4770,N_33,N_424);
and U4771 (N_4771,N_1472,N_107);
nand U4772 (N_4772,N_2523,N_2057);
nand U4773 (N_4773,N_619,N_679);
nor U4774 (N_4774,N_1637,N_2786);
nand U4775 (N_4775,N_963,N_1843);
or U4776 (N_4776,N_1471,N_1134);
or U4777 (N_4777,N_668,N_2347);
and U4778 (N_4778,N_1667,N_1980);
nor U4779 (N_4779,N_1614,N_1209);
nor U4780 (N_4780,N_2451,N_614);
nand U4781 (N_4781,N_173,N_977);
nand U4782 (N_4782,N_1814,N_158);
nand U4783 (N_4783,N_75,N_1063);
xnor U4784 (N_4784,N_279,N_1423);
xor U4785 (N_4785,N_2838,N_2089);
xnor U4786 (N_4786,N_1978,N_2177);
and U4787 (N_4787,N_2845,N_717);
nor U4788 (N_4788,N_568,N_2381);
xor U4789 (N_4789,N_2532,N_1787);
xnor U4790 (N_4790,N_496,N_2089);
and U4791 (N_4791,N_1089,N_1763);
xnor U4792 (N_4792,N_2902,N_540);
xor U4793 (N_4793,N_1683,N_220);
xnor U4794 (N_4794,N_1069,N_990);
nand U4795 (N_4795,N_1301,N_2262);
xor U4796 (N_4796,N_2889,N_2687);
and U4797 (N_4797,N_1266,N_2424);
or U4798 (N_4798,N_907,N_2113);
xor U4799 (N_4799,N_1094,N_506);
xor U4800 (N_4800,N_476,N_1553);
and U4801 (N_4801,N_2223,N_900);
xnor U4802 (N_4802,N_2309,N_162);
nor U4803 (N_4803,N_2882,N_344);
or U4804 (N_4804,N_16,N_1868);
xnor U4805 (N_4805,N_686,N_747);
nor U4806 (N_4806,N_1922,N_1915);
or U4807 (N_4807,N_2577,N_2094);
xnor U4808 (N_4808,N_2316,N_2245);
xnor U4809 (N_4809,N_2806,N_1206);
and U4810 (N_4810,N_937,N_1438);
or U4811 (N_4811,N_1727,N_853);
nand U4812 (N_4812,N_2044,N_400);
nand U4813 (N_4813,N_839,N_2041);
nand U4814 (N_4814,N_1048,N_196);
or U4815 (N_4815,N_615,N_150);
nand U4816 (N_4816,N_651,N_47);
nand U4817 (N_4817,N_1393,N_42);
and U4818 (N_4818,N_842,N_1156);
or U4819 (N_4819,N_1467,N_1619);
nor U4820 (N_4820,N_1194,N_2419);
nor U4821 (N_4821,N_969,N_2622);
or U4822 (N_4822,N_1784,N_1269);
and U4823 (N_4823,N_2181,N_2454);
and U4824 (N_4824,N_2726,N_51);
or U4825 (N_4825,N_128,N_1850);
or U4826 (N_4826,N_1300,N_253);
and U4827 (N_4827,N_2271,N_1281);
nor U4828 (N_4828,N_916,N_1929);
nand U4829 (N_4829,N_2913,N_1519);
xor U4830 (N_4830,N_2340,N_456);
or U4831 (N_4831,N_1559,N_1927);
nand U4832 (N_4832,N_1936,N_2388);
nand U4833 (N_4833,N_1895,N_724);
nor U4834 (N_4834,N_1972,N_1334);
nor U4835 (N_4835,N_1474,N_940);
nor U4836 (N_4836,N_2413,N_859);
nand U4837 (N_4837,N_2573,N_1756);
and U4838 (N_4838,N_586,N_2256);
xnor U4839 (N_4839,N_578,N_1975);
nand U4840 (N_4840,N_650,N_1234);
nor U4841 (N_4841,N_2409,N_2460);
nor U4842 (N_4842,N_920,N_1221);
or U4843 (N_4843,N_886,N_1365);
nand U4844 (N_4844,N_2158,N_2788);
nand U4845 (N_4845,N_694,N_9);
xor U4846 (N_4846,N_1294,N_30);
nor U4847 (N_4847,N_574,N_2702);
nor U4848 (N_4848,N_1558,N_1001);
nor U4849 (N_4849,N_75,N_1815);
nand U4850 (N_4850,N_2729,N_1821);
or U4851 (N_4851,N_1508,N_1789);
xnor U4852 (N_4852,N_2769,N_2751);
nor U4853 (N_4853,N_473,N_2867);
and U4854 (N_4854,N_1592,N_2492);
xor U4855 (N_4855,N_561,N_1430);
and U4856 (N_4856,N_220,N_2126);
and U4857 (N_4857,N_398,N_2111);
xor U4858 (N_4858,N_501,N_2006);
nor U4859 (N_4859,N_523,N_1533);
nor U4860 (N_4860,N_1360,N_1336);
nand U4861 (N_4861,N_2668,N_1686);
nand U4862 (N_4862,N_1209,N_1738);
or U4863 (N_4863,N_1537,N_1879);
nand U4864 (N_4864,N_2251,N_1971);
nor U4865 (N_4865,N_2574,N_2381);
or U4866 (N_4866,N_2724,N_1189);
and U4867 (N_4867,N_1360,N_812);
and U4868 (N_4868,N_1064,N_2195);
nor U4869 (N_4869,N_1198,N_1390);
and U4870 (N_4870,N_1560,N_1387);
xnor U4871 (N_4871,N_2696,N_677);
and U4872 (N_4872,N_84,N_2163);
nand U4873 (N_4873,N_668,N_803);
xnor U4874 (N_4874,N_1428,N_2367);
nor U4875 (N_4875,N_272,N_1973);
and U4876 (N_4876,N_1979,N_2697);
nand U4877 (N_4877,N_1737,N_1908);
or U4878 (N_4878,N_2123,N_1562);
and U4879 (N_4879,N_371,N_1926);
xor U4880 (N_4880,N_1935,N_160);
nor U4881 (N_4881,N_680,N_2324);
or U4882 (N_4882,N_461,N_1757);
nand U4883 (N_4883,N_368,N_2089);
and U4884 (N_4884,N_2856,N_2763);
nor U4885 (N_4885,N_2814,N_148);
nor U4886 (N_4886,N_2596,N_121);
or U4887 (N_4887,N_857,N_560);
nor U4888 (N_4888,N_1337,N_2792);
and U4889 (N_4889,N_2302,N_1532);
nand U4890 (N_4890,N_1466,N_2500);
or U4891 (N_4891,N_2085,N_2867);
nand U4892 (N_4892,N_2587,N_1516);
nand U4893 (N_4893,N_1490,N_808);
nand U4894 (N_4894,N_1374,N_2336);
nand U4895 (N_4895,N_2924,N_1413);
nand U4896 (N_4896,N_908,N_239);
nand U4897 (N_4897,N_218,N_650);
nand U4898 (N_4898,N_362,N_904);
and U4899 (N_4899,N_2838,N_1433);
or U4900 (N_4900,N_1867,N_1215);
and U4901 (N_4901,N_302,N_2494);
xor U4902 (N_4902,N_2642,N_1234);
and U4903 (N_4903,N_24,N_142);
and U4904 (N_4904,N_1491,N_1722);
nand U4905 (N_4905,N_1636,N_2276);
nor U4906 (N_4906,N_2185,N_713);
or U4907 (N_4907,N_1036,N_2352);
nor U4908 (N_4908,N_2204,N_433);
or U4909 (N_4909,N_2431,N_153);
nand U4910 (N_4910,N_1949,N_2474);
or U4911 (N_4911,N_1074,N_545);
and U4912 (N_4912,N_237,N_880);
xor U4913 (N_4913,N_1445,N_1808);
nor U4914 (N_4914,N_401,N_206);
xor U4915 (N_4915,N_1012,N_2672);
xor U4916 (N_4916,N_2174,N_554);
nor U4917 (N_4917,N_2554,N_729);
xor U4918 (N_4918,N_1555,N_2299);
nor U4919 (N_4919,N_970,N_533);
and U4920 (N_4920,N_1753,N_2810);
nand U4921 (N_4921,N_964,N_2647);
or U4922 (N_4922,N_1852,N_306);
nand U4923 (N_4923,N_1032,N_363);
and U4924 (N_4924,N_1998,N_1197);
xor U4925 (N_4925,N_2350,N_303);
nand U4926 (N_4926,N_164,N_1955);
and U4927 (N_4927,N_1560,N_2373);
nand U4928 (N_4928,N_2887,N_127);
and U4929 (N_4929,N_1483,N_1983);
xor U4930 (N_4930,N_2179,N_1625);
nor U4931 (N_4931,N_2256,N_2873);
or U4932 (N_4932,N_209,N_2858);
and U4933 (N_4933,N_771,N_594);
nor U4934 (N_4934,N_883,N_146);
nor U4935 (N_4935,N_2383,N_1541);
xor U4936 (N_4936,N_2240,N_393);
nand U4937 (N_4937,N_94,N_957);
nand U4938 (N_4938,N_60,N_2551);
nand U4939 (N_4939,N_1191,N_2937);
or U4940 (N_4940,N_711,N_2645);
xnor U4941 (N_4941,N_560,N_68);
nand U4942 (N_4942,N_764,N_1917);
or U4943 (N_4943,N_558,N_657);
nand U4944 (N_4944,N_2596,N_2418);
and U4945 (N_4945,N_388,N_1105);
and U4946 (N_4946,N_2306,N_1283);
or U4947 (N_4947,N_700,N_2131);
nand U4948 (N_4948,N_2464,N_122);
nand U4949 (N_4949,N_177,N_886);
and U4950 (N_4950,N_315,N_2144);
nor U4951 (N_4951,N_647,N_778);
or U4952 (N_4952,N_2591,N_1970);
and U4953 (N_4953,N_29,N_1840);
nand U4954 (N_4954,N_1342,N_357);
nor U4955 (N_4955,N_602,N_1220);
nor U4956 (N_4956,N_1010,N_1481);
nand U4957 (N_4957,N_457,N_2420);
nand U4958 (N_4958,N_898,N_478);
nand U4959 (N_4959,N_585,N_1781);
nor U4960 (N_4960,N_2012,N_216);
and U4961 (N_4961,N_1666,N_849);
nor U4962 (N_4962,N_502,N_2591);
or U4963 (N_4963,N_2463,N_310);
nand U4964 (N_4964,N_2875,N_814);
xor U4965 (N_4965,N_1886,N_2671);
nor U4966 (N_4966,N_1944,N_574);
and U4967 (N_4967,N_2823,N_1350);
nor U4968 (N_4968,N_1033,N_1889);
or U4969 (N_4969,N_257,N_660);
xnor U4970 (N_4970,N_2275,N_2023);
nor U4971 (N_4971,N_2994,N_2878);
nand U4972 (N_4972,N_351,N_792);
nor U4973 (N_4973,N_773,N_1174);
nor U4974 (N_4974,N_1614,N_909);
or U4975 (N_4975,N_510,N_1418);
xor U4976 (N_4976,N_1614,N_975);
nor U4977 (N_4977,N_1919,N_2427);
nor U4978 (N_4978,N_1964,N_2041);
or U4979 (N_4979,N_515,N_516);
xor U4980 (N_4980,N_2997,N_2133);
and U4981 (N_4981,N_1008,N_182);
or U4982 (N_4982,N_2609,N_1993);
or U4983 (N_4983,N_1092,N_2575);
and U4984 (N_4984,N_2440,N_267);
nand U4985 (N_4985,N_393,N_315);
and U4986 (N_4986,N_1528,N_130);
nand U4987 (N_4987,N_1757,N_677);
and U4988 (N_4988,N_1934,N_1690);
or U4989 (N_4989,N_2441,N_2723);
nand U4990 (N_4990,N_1286,N_1573);
or U4991 (N_4991,N_1940,N_448);
xnor U4992 (N_4992,N_182,N_1489);
nor U4993 (N_4993,N_488,N_1471);
nand U4994 (N_4994,N_1232,N_1107);
xor U4995 (N_4995,N_2454,N_1585);
and U4996 (N_4996,N_2239,N_732);
nor U4997 (N_4997,N_2762,N_1479);
xnor U4998 (N_4998,N_2650,N_742);
and U4999 (N_4999,N_2720,N_2809);
or U5000 (N_5000,N_2368,N_1545);
xnor U5001 (N_5001,N_975,N_81);
xor U5002 (N_5002,N_2805,N_1340);
nor U5003 (N_5003,N_1855,N_763);
or U5004 (N_5004,N_1562,N_2832);
nand U5005 (N_5005,N_1484,N_1091);
xor U5006 (N_5006,N_1688,N_1269);
nand U5007 (N_5007,N_870,N_2321);
or U5008 (N_5008,N_2190,N_2793);
nand U5009 (N_5009,N_2817,N_55);
nor U5010 (N_5010,N_1010,N_1442);
xnor U5011 (N_5011,N_1998,N_1672);
and U5012 (N_5012,N_1586,N_2505);
nand U5013 (N_5013,N_2824,N_1639);
nor U5014 (N_5014,N_1330,N_391);
and U5015 (N_5015,N_1319,N_1348);
xnor U5016 (N_5016,N_2633,N_191);
nor U5017 (N_5017,N_1700,N_1721);
nand U5018 (N_5018,N_2000,N_1689);
or U5019 (N_5019,N_682,N_775);
nor U5020 (N_5020,N_1263,N_2502);
and U5021 (N_5021,N_2649,N_2089);
nand U5022 (N_5022,N_290,N_1631);
or U5023 (N_5023,N_1789,N_833);
or U5024 (N_5024,N_179,N_2889);
and U5025 (N_5025,N_681,N_2458);
nor U5026 (N_5026,N_2392,N_802);
xor U5027 (N_5027,N_661,N_1681);
or U5028 (N_5028,N_2385,N_2255);
nor U5029 (N_5029,N_104,N_1150);
xnor U5030 (N_5030,N_2705,N_1434);
nor U5031 (N_5031,N_2178,N_134);
nor U5032 (N_5032,N_372,N_919);
or U5033 (N_5033,N_958,N_2152);
or U5034 (N_5034,N_2671,N_128);
and U5035 (N_5035,N_1571,N_1996);
xor U5036 (N_5036,N_135,N_2128);
nand U5037 (N_5037,N_266,N_600);
and U5038 (N_5038,N_641,N_1500);
nand U5039 (N_5039,N_2702,N_2515);
xnor U5040 (N_5040,N_2183,N_1009);
and U5041 (N_5041,N_1016,N_2743);
nor U5042 (N_5042,N_487,N_533);
and U5043 (N_5043,N_1689,N_1511);
nor U5044 (N_5044,N_908,N_2094);
nor U5045 (N_5045,N_1149,N_1635);
nand U5046 (N_5046,N_2030,N_1460);
nor U5047 (N_5047,N_263,N_2559);
and U5048 (N_5048,N_2447,N_1670);
and U5049 (N_5049,N_1618,N_1478);
nand U5050 (N_5050,N_1312,N_186);
xnor U5051 (N_5051,N_2664,N_1126);
and U5052 (N_5052,N_22,N_1370);
nand U5053 (N_5053,N_1757,N_1413);
nand U5054 (N_5054,N_157,N_1652);
and U5055 (N_5055,N_305,N_2246);
or U5056 (N_5056,N_84,N_2839);
and U5057 (N_5057,N_686,N_2329);
and U5058 (N_5058,N_2635,N_33);
xor U5059 (N_5059,N_1042,N_1528);
xnor U5060 (N_5060,N_2917,N_2706);
and U5061 (N_5061,N_715,N_1874);
and U5062 (N_5062,N_296,N_2371);
nand U5063 (N_5063,N_1367,N_666);
and U5064 (N_5064,N_2188,N_2394);
or U5065 (N_5065,N_1158,N_525);
and U5066 (N_5066,N_2032,N_697);
xnor U5067 (N_5067,N_2688,N_2596);
xnor U5068 (N_5068,N_1226,N_1387);
nand U5069 (N_5069,N_1825,N_1025);
nor U5070 (N_5070,N_2729,N_2856);
xnor U5071 (N_5071,N_2485,N_309);
xor U5072 (N_5072,N_1352,N_2153);
nor U5073 (N_5073,N_327,N_2942);
xor U5074 (N_5074,N_2017,N_1194);
or U5075 (N_5075,N_2798,N_1848);
nand U5076 (N_5076,N_2005,N_1500);
or U5077 (N_5077,N_2371,N_1528);
and U5078 (N_5078,N_927,N_322);
or U5079 (N_5079,N_1523,N_2290);
and U5080 (N_5080,N_838,N_2647);
and U5081 (N_5081,N_2619,N_1836);
or U5082 (N_5082,N_2639,N_1010);
or U5083 (N_5083,N_1592,N_1050);
nor U5084 (N_5084,N_986,N_472);
nand U5085 (N_5085,N_2829,N_393);
nand U5086 (N_5086,N_681,N_1788);
xor U5087 (N_5087,N_2811,N_1410);
or U5088 (N_5088,N_276,N_582);
or U5089 (N_5089,N_802,N_1747);
xnor U5090 (N_5090,N_2036,N_1862);
xnor U5091 (N_5091,N_873,N_1087);
xor U5092 (N_5092,N_78,N_1900);
or U5093 (N_5093,N_1220,N_2033);
nor U5094 (N_5094,N_394,N_1454);
nor U5095 (N_5095,N_946,N_655);
nand U5096 (N_5096,N_1318,N_2869);
nand U5097 (N_5097,N_1821,N_2924);
xor U5098 (N_5098,N_353,N_2337);
and U5099 (N_5099,N_2878,N_662);
or U5100 (N_5100,N_2208,N_329);
nor U5101 (N_5101,N_2009,N_1168);
and U5102 (N_5102,N_630,N_2206);
nand U5103 (N_5103,N_2226,N_1239);
or U5104 (N_5104,N_237,N_1139);
nor U5105 (N_5105,N_326,N_414);
and U5106 (N_5106,N_559,N_9);
and U5107 (N_5107,N_1355,N_638);
nor U5108 (N_5108,N_2221,N_1547);
nand U5109 (N_5109,N_658,N_127);
nand U5110 (N_5110,N_1621,N_1664);
or U5111 (N_5111,N_111,N_772);
and U5112 (N_5112,N_1727,N_2757);
nor U5113 (N_5113,N_321,N_553);
nand U5114 (N_5114,N_962,N_1474);
nor U5115 (N_5115,N_771,N_2782);
nor U5116 (N_5116,N_28,N_74);
or U5117 (N_5117,N_1641,N_1122);
nor U5118 (N_5118,N_1315,N_611);
xnor U5119 (N_5119,N_2085,N_2899);
and U5120 (N_5120,N_330,N_663);
and U5121 (N_5121,N_2199,N_1472);
xor U5122 (N_5122,N_2560,N_386);
nor U5123 (N_5123,N_2592,N_1188);
and U5124 (N_5124,N_1089,N_2686);
nand U5125 (N_5125,N_1092,N_2169);
nand U5126 (N_5126,N_2189,N_2185);
xor U5127 (N_5127,N_379,N_2833);
xnor U5128 (N_5128,N_433,N_329);
and U5129 (N_5129,N_1300,N_2310);
or U5130 (N_5130,N_763,N_628);
xor U5131 (N_5131,N_683,N_732);
xnor U5132 (N_5132,N_1476,N_1236);
or U5133 (N_5133,N_2088,N_77);
and U5134 (N_5134,N_1280,N_2990);
nand U5135 (N_5135,N_1112,N_233);
and U5136 (N_5136,N_824,N_1743);
nand U5137 (N_5137,N_677,N_595);
xor U5138 (N_5138,N_2304,N_87);
or U5139 (N_5139,N_1067,N_1003);
xor U5140 (N_5140,N_1173,N_785);
nor U5141 (N_5141,N_2631,N_990);
or U5142 (N_5142,N_932,N_1998);
nor U5143 (N_5143,N_1167,N_985);
or U5144 (N_5144,N_775,N_1235);
nor U5145 (N_5145,N_123,N_2206);
nor U5146 (N_5146,N_123,N_2816);
or U5147 (N_5147,N_1697,N_1517);
or U5148 (N_5148,N_570,N_499);
or U5149 (N_5149,N_2493,N_251);
xor U5150 (N_5150,N_2769,N_1620);
and U5151 (N_5151,N_2035,N_1152);
nor U5152 (N_5152,N_539,N_80);
nor U5153 (N_5153,N_179,N_244);
nor U5154 (N_5154,N_1678,N_1814);
or U5155 (N_5155,N_1339,N_2569);
or U5156 (N_5156,N_329,N_1664);
or U5157 (N_5157,N_2640,N_2624);
xor U5158 (N_5158,N_887,N_143);
nand U5159 (N_5159,N_1947,N_1590);
or U5160 (N_5160,N_2085,N_1869);
nor U5161 (N_5161,N_440,N_2154);
nand U5162 (N_5162,N_259,N_431);
nor U5163 (N_5163,N_1570,N_673);
nand U5164 (N_5164,N_550,N_1948);
or U5165 (N_5165,N_443,N_2604);
xor U5166 (N_5166,N_372,N_209);
xor U5167 (N_5167,N_179,N_2688);
and U5168 (N_5168,N_384,N_1311);
and U5169 (N_5169,N_1537,N_2782);
xor U5170 (N_5170,N_1738,N_1617);
nor U5171 (N_5171,N_2967,N_1013);
nor U5172 (N_5172,N_186,N_2816);
nor U5173 (N_5173,N_1821,N_1405);
nand U5174 (N_5174,N_2804,N_455);
and U5175 (N_5175,N_2260,N_1311);
xor U5176 (N_5176,N_1417,N_239);
xnor U5177 (N_5177,N_2389,N_2485);
nor U5178 (N_5178,N_1421,N_704);
xnor U5179 (N_5179,N_2381,N_2161);
nor U5180 (N_5180,N_1061,N_1044);
and U5181 (N_5181,N_2095,N_2754);
or U5182 (N_5182,N_2426,N_2259);
xnor U5183 (N_5183,N_2382,N_2328);
and U5184 (N_5184,N_773,N_2347);
and U5185 (N_5185,N_1428,N_2438);
or U5186 (N_5186,N_1768,N_1737);
nand U5187 (N_5187,N_176,N_922);
nand U5188 (N_5188,N_1175,N_1354);
nor U5189 (N_5189,N_2468,N_822);
or U5190 (N_5190,N_1814,N_1303);
nand U5191 (N_5191,N_2053,N_2804);
or U5192 (N_5192,N_1205,N_2277);
nor U5193 (N_5193,N_662,N_1963);
and U5194 (N_5194,N_2241,N_1652);
xor U5195 (N_5195,N_2709,N_1002);
or U5196 (N_5196,N_143,N_860);
or U5197 (N_5197,N_711,N_1926);
and U5198 (N_5198,N_876,N_748);
and U5199 (N_5199,N_2913,N_81);
nand U5200 (N_5200,N_2846,N_2666);
and U5201 (N_5201,N_413,N_1713);
and U5202 (N_5202,N_2298,N_40);
xnor U5203 (N_5203,N_886,N_1816);
and U5204 (N_5204,N_1209,N_1649);
or U5205 (N_5205,N_1540,N_280);
xor U5206 (N_5206,N_1814,N_1214);
nor U5207 (N_5207,N_1841,N_1898);
or U5208 (N_5208,N_2041,N_150);
and U5209 (N_5209,N_1463,N_2617);
xor U5210 (N_5210,N_2158,N_1161);
and U5211 (N_5211,N_616,N_1155);
and U5212 (N_5212,N_245,N_111);
xor U5213 (N_5213,N_1544,N_1665);
nor U5214 (N_5214,N_381,N_1739);
nor U5215 (N_5215,N_2740,N_1950);
xor U5216 (N_5216,N_2008,N_2978);
xor U5217 (N_5217,N_9,N_533);
and U5218 (N_5218,N_1194,N_234);
nor U5219 (N_5219,N_974,N_2721);
nor U5220 (N_5220,N_1425,N_1146);
or U5221 (N_5221,N_698,N_112);
or U5222 (N_5222,N_685,N_536);
and U5223 (N_5223,N_365,N_851);
or U5224 (N_5224,N_1803,N_442);
or U5225 (N_5225,N_2549,N_303);
and U5226 (N_5226,N_1459,N_1670);
and U5227 (N_5227,N_1253,N_818);
or U5228 (N_5228,N_751,N_919);
nand U5229 (N_5229,N_365,N_1908);
nand U5230 (N_5230,N_1111,N_2242);
nand U5231 (N_5231,N_2687,N_754);
nor U5232 (N_5232,N_626,N_257);
and U5233 (N_5233,N_2521,N_2039);
nor U5234 (N_5234,N_2861,N_1752);
nor U5235 (N_5235,N_65,N_1782);
or U5236 (N_5236,N_750,N_582);
xor U5237 (N_5237,N_989,N_1792);
and U5238 (N_5238,N_1252,N_2595);
nand U5239 (N_5239,N_1577,N_2029);
nor U5240 (N_5240,N_2770,N_2661);
and U5241 (N_5241,N_2179,N_303);
and U5242 (N_5242,N_2185,N_1000);
nor U5243 (N_5243,N_2203,N_478);
and U5244 (N_5244,N_1536,N_803);
or U5245 (N_5245,N_1393,N_1908);
nor U5246 (N_5246,N_969,N_306);
and U5247 (N_5247,N_2194,N_19);
nor U5248 (N_5248,N_1460,N_1442);
xnor U5249 (N_5249,N_2162,N_1940);
nor U5250 (N_5250,N_1123,N_1235);
nor U5251 (N_5251,N_1612,N_567);
xor U5252 (N_5252,N_2525,N_1803);
and U5253 (N_5253,N_1963,N_1018);
nor U5254 (N_5254,N_144,N_2371);
xnor U5255 (N_5255,N_2364,N_952);
nand U5256 (N_5256,N_2411,N_1254);
nand U5257 (N_5257,N_2199,N_957);
nor U5258 (N_5258,N_2493,N_1398);
nor U5259 (N_5259,N_52,N_2757);
xor U5260 (N_5260,N_2374,N_194);
xnor U5261 (N_5261,N_2922,N_691);
or U5262 (N_5262,N_1981,N_1435);
or U5263 (N_5263,N_658,N_2672);
nand U5264 (N_5264,N_2313,N_2873);
or U5265 (N_5265,N_2566,N_277);
or U5266 (N_5266,N_997,N_1899);
and U5267 (N_5267,N_2445,N_2093);
xnor U5268 (N_5268,N_2578,N_2694);
xor U5269 (N_5269,N_1889,N_1894);
nand U5270 (N_5270,N_1657,N_2566);
and U5271 (N_5271,N_233,N_933);
and U5272 (N_5272,N_1195,N_808);
or U5273 (N_5273,N_2258,N_48);
or U5274 (N_5274,N_1387,N_1172);
nor U5275 (N_5275,N_1412,N_1712);
xor U5276 (N_5276,N_2018,N_2337);
and U5277 (N_5277,N_2248,N_2565);
nor U5278 (N_5278,N_335,N_1952);
xor U5279 (N_5279,N_1222,N_394);
or U5280 (N_5280,N_2846,N_695);
nand U5281 (N_5281,N_2505,N_1449);
and U5282 (N_5282,N_2375,N_2992);
nor U5283 (N_5283,N_2963,N_1533);
nand U5284 (N_5284,N_1714,N_1054);
xor U5285 (N_5285,N_140,N_1481);
xor U5286 (N_5286,N_129,N_1698);
nor U5287 (N_5287,N_2724,N_990);
or U5288 (N_5288,N_1877,N_2821);
nor U5289 (N_5289,N_177,N_2792);
xnor U5290 (N_5290,N_2010,N_989);
xnor U5291 (N_5291,N_2369,N_589);
nand U5292 (N_5292,N_1104,N_994);
and U5293 (N_5293,N_255,N_1046);
xor U5294 (N_5294,N_1119,N_2715);
nand U5295 (N_5295,N_1877,N_2532);
and U5296 (N_5296,N_1963,N_2603);
or U5297 (N_5297,N_572,N_486);
and U5298 (N_5298,N_1303,N_244);
xor U5299 (N_5299,N_2213,N_591);
nor U5300 (N_5300,N_1115,N_1432);
nor U5301 (N_5301,N_360,N_2019);
and U5302 (N_5302,N_2092,N_855);
nand U5303 (N_5303,N_626,N_1085);
or U5304 (N_5304,N_805,N_1805);
and U5305 (N_5305,N_1060,N_2479);
xnor U5306 (N_5306,N_1546,N_2671);
nand U5307 (N_5307,N_2191,N_2955);
xor U5308 (N_5308,N_294,N_2255);
nand U5309 (N_5309,N_707,N_2537);
nand U5310 (N_5310,N_1764,N_490);
nand U5311 (N_5311,N_1015,N_1144);
nand U5312 (N_5312,N_2427,N_177);
and U5313 (N_5313,N_391,N_2148);
or U5314 (N_5314,N_2287,N_989);
or U5315 (N_5315,N_1620,N_288);
nand U5316 (N_5316,N_313,N_1983);
nand U5317 (N_5317,N_1129,N_1305);
nor U5318 (N_5318,N_1874,N_1846);
or U5319 (N_5319,N_2843,N_536);
or U5320 (N_5320,N_852,N_717);
nand U5321 (N_5321,N_1649,N_354);
and U5322 (N_5322,N_2457,N_948);
or U5323 (N_5323,N_2643,N_1045);
and U5324 (N_5324,N_2413,N_46);
and U5325 (N_5325,N_2305,N_1967);
or U5326 (N_5326,N_1628,N_995);
xnor U5327 (N_5327,N_1984,N_999);
xor U5328 (N_5328,N_1300,N_2884);
and U5329 (N_5329,N_1422,N_1999);
nor U5330 (N_5330,N_2537,N_2354);
nor U5331 (N_5331,N_1711,N_2028);
or U5332 (N_5332,N_1525,N_992);
xor U5333 (N_5333,N_1623,N_2020);
nand U5334 (N_5334,N_1223,N_2631);
nor U5335 (N_5335,N_2336,N_1214);
xnor U5336 (N_5336,N_2692,N_17);
xor U5337 (N_5337,N_822,N_1225);
xnor U5338 (N_5338,N_1271,N_29);
xnor U5339 (N_5339,N_2852,N_2992);
xor U5340 (N_5340,N_1549,N_824);
nor U5341 (N_5341,N_1172,N_2957);
nor U5342 (N_5342,N_1365,N_2424);
or U5343 (N_5343,N_2104,N_1956);
or U5344 (N_5344,N_2515,N_334);
xor U5345 (N_5345,N_1738,N_1228);
and U5346 (N_5346,N_1800,N_2378);
nand U5347 (N_5347,N_152,N_2480);
and U5348 (N_5348,N_2869,N_812);
nand U5349 (N_5349,N_2882,N_2985);
nor U5350 (N_5350,N_161,N_722);
and U5351 (N_5351,N_585,N_601);
and U5352 (N_5352,N_2539,N_2915);
nand U5353 (N_5353,N_1176,N_2081);
nor U5354 (N_5354,N_716,N_1042);
xor U5355 (N_5355,N_61,N_935);
and U5356 (N_5356,N_1616,N_399);
xnor U5357 (N_5357,N_1762,N_2823);
and U5358 (N_5358,N_313,N_777);
xor U5359 (N_5359,N_2688,N_273);
nand U5360 (N_5360,N_139,N_563);
nand U5361 (N_5361,N_329,N_795);
or U5362 (N_5362,N_1060,N_1013);
and U5363 (N_5363,N_390,N_1442);
and U5364 (N_5364,N_1658,N_2319);
or U5365 (N_5365,N_2424,N_330);
nor U5366 (N_5366,N_2074,N_1238);
or U5367 (N_5367,N_513,N_996);
or U5368 (N_5368,N_1841,N_2068);
nor U5369 (N_5369,N_1521,N_364);
nand U5370 (N_5370,N_1613,N_2234);
nor U5371 (N_5371,N_265,N_2450);
xnor U5372 (N_5372,N_245,N_1756);
nor U5373 (N_5373,N_370,N_1716);
xor U5374 (N_5374,N_954,N_2418);
xor U5375 (N_5375,N_572,N_2767);
and U5376 (N_5376,N_865,N_1297);
and U5377 (N_5377,N_297,N_1335);
xnor U5378 (N_5378,N_1786,N_883);
or U5379 (N_5379,N_499,N_1769);
nand U5380 (N_5380,N_2913,N_2556);
or U5381 (N_5381,N_1696,N_2311);
and U5382 (N_5382,N_1961,N_1220);
or U5383 (N_5383,N_2523,N_1172);
and U5384 (N_5384,N_1572,N_1047);
nand U5385 (N_5385,N_429,N_1003);
and U5386 (N_5386,N_351,N_2917);
xor U5387 (N_5387,N_213,N_1753);
or U5388 (N_5388,N_2290,N_2520);
or U5389 (N_5389,N_1444,N_2081);
nand U5390 (N_5390,N_1543,N_2743);
nor U5391 (N_5391,N_977,N_421);
nand U5392 (N_5392,N_719,N_743);
nand U5393 (N_5393,N_276,N_759);
nand U5394 (N_5394,N_1304,N_333);
nor U5395 (N_5395,N_1408,N_2104);
xor U5396 (N_5396,N_2450,N_2170);
or U5397 (N_5397,N_2527,N_1492);
nor U5398 (N_5398,N_612,N_124);
or U5399 (N_5399,N_2999,N_1834);
and U5400 (N_5400,N_1305,N_2523);
nand U5401 (N_5401,N_2030,N_2828);
and U5402 (N_5402,N_2086,N_1546);
or U5403 (N_5403,N_878,N_2035);
nand U5404 (N_5404,N_1452,N_1887);
nand U5405 (N_5405,N_2261,N_2688);
nor U5406 (N_5406,N_1226,N_1183);
nand U5407 (N_5407,N_291,N_2281);
xnor U5408 (N_5408,N_429,N_514);
nand U5409 (N_5409,N_2768,N_1627);
and U5410 (N_5410,N_2779,N_1498);
xnor U5411 (N_5411,N_2189,N_1729);
and U5412 (N_5412,N_1395,N_1970);
and U5413 (N_5413,N_487,N_819);
nand U5414 (N_5414,N_505,N_1173);
nor U5415 (N_5415,N_306,N_1338);
nand U5416 (N_5416,N_392,N_2029);
nor U5417 (N_5417,N_1652,N_1120);
nor U5418 (N_5418,N_1685,N_1403);
and U5419 (N_5419,N_1630,N_2452);
or U5420 (N_5420,N_2873,N_1083);
and U5421 (N_5421,N_1468,N_41);
nand U5422 (N_5422,N_1823,N_272);
nand U5423 (N_5423,N_760,N_363);
nand U5424 (N_5424,N_1959,N_1761);
or U5425 (N_5425,N_355,N_78);
and U5426 (N_5426,N_513,N_1403);
nor U5427 (N_5427,N_375,N_2202);
nor U5428 (N_5428,N_2394,N_937);
nand U5429 (N_5429,N_281,N_1442);
nand U5430 (N_5430,N_375,N_2300);
nor U5431 (N_5431,N_1149,N_1756);
or U5432 (N_5432,N_2454,N_1447);
xor U5433 (N_5433,N_1077,N_2970);
xor U5434 (N_5434,N_2407,N_1181);
nor U5435 (N_5435,N_2733,N_647);
and U5436 (N_5436,N_1661,N_1189);
and U5437 (N_5437,N_826,N_2017);
and U5438 (N_5438,N_1854,N_2210);
nor U5439 (N_5439,N_2255,N_2153);
nor U5440 (N_5440,N_564,N_2819);
and U5441 (N_5441,N_1601,N_179);
nand U5442 (N_5442,N_186,N_441);
and U5443 (N_5443,N_389,N_1554);
xnor U5444 (N_5444,N_1828,N_2068);
xnor U5445 (N_5445,N_932,N_2547);
nand U5446 (N_5446,N_1745,N_1304);
xnor U5447 (N_5447,N_30,N_126);
or U5448 (N_5448,N_53,N_1834);
nor U5449 (N_5449,N_2802,N_2331);
or U5450 (N_5450,N_370,N_1760);
nor U5451 (N_5451,N_2507,N_1703);
or U5452 (N_5452,N_915,N_287);
nand U5453 (N_5453,N_2154,N_1271);
nand U5454 (N_5454,N_1219,N_2678);
xnor U5455 (N_5455,N_1518,N_2800);
or U5456 (N_5456,N_2419,N_418);
nor U5457 (N_5457,N_1793,N_1278);
nor U5458 (N_5458,N_1772,N_1479);
xnor U5459 (N_5459,N_2532,N_1805);
xor U5460 (N_5460,N_1552,N_1380);
and U5461 (N_5461,N_853,N_2246);
xnor U5462 (N_5462,N_1961,N_395);
nand U5463 (N_5463,N_1589,N_2475);
xnor U5464 (N_5464,N_378,N_1444);
or U5465 (N_5465,N_1859,N_2163);
or U5466 (N_5466,N_2934,N_512);
nand U5467 (N_5467,N_2233,N_77);
nor U5468 (N_5468,N_297,N_2374);
or U5469 (N_5469,N_2828,N_2136);
nor U5470 (N_5470,N_2638,N_1871);
or U5471 (N_5471,N_2455,N_2874);
xor U5472 (N_5472,N_1838,N_2275);
nand U5473 (N_5473,N_461,N_1184);
or U5474 (N_5474,N_326,N_2249);
nor U5475 (N_5475,N_835,N_63);
nor U5476 (N_5476,N_9,N_944);
xor U5477 (N_5477,N_2362,N_1736);
or U5478 (N_5478,N_1603,N_2563);
nand U5479 (N_5479,N_1697,N_1244);
xor U5480 (N_5480,N_2998,N_287);
xnor U5481 (N_5481,N_198,N_1040);
nand U5482 (N_5482,N_2769,N_2942);
nand U5483 (N_5483,N_2024,N_2692);
xnor U5484 (N_5484,N_662,N_2001);
nand U5485 (N_5485,N_473,N_1119);
nand U5486 (N_5486,N_832,N_1812);
or U5487 (N_5487,N_1849,N_1153);
xor U5488 (N_5488,N_1391,N_1543);
nand U5489 (N_5489,N_2742,N_1206);
xor U5490 (N_5490,N_2180,N_1241);
and U5491 (N_5491,N_1996,N_1939);
xor U5492 (N_5492,N_2368,N_2866);
nor U5493 (N_5493,N_935,N_686);
nand U5494 (N_5494,N_748,N_1854);
and U5495 (N_5495,N_957,N_2047);
and U5496 (N_5496,N_1102,N_1710);
xor U5497 (N_5497,N_850,N_1806);
nand U5498 (N_5498,N_2755,N_1711);
or U5499 (N_5499,N_1116,N_2344);
nor U5500 (N_5500,N_1181,N_2950);
nand U5501 (N_5501,N_1584,N_2727);
xor U5502 (N_5502,N_2649,N_2027);
nand U5503 (N_5503,N_2598,N_2884);
and U5504 (N_5504,N_384,N_2372);
nand U5505 (N_5505,N_2115,N_1098);
nor U5506 (N_5506,N_2808,N_2374);
nor U5507 (N_5507,N_2538,N_1593);
nor U5508 (N_5508,N_2476,N_2562);
xnor U5509 (N_5509,N_37,N_1921);
nor U5510 (N_5510,N_2100,N_2511);
or U5511 (N_5511,N_2535,N_2061);
or U5512 (N_5512,N_2677,N_2288);
or U5513 (N_5513,N_744,N_755);
xor U5514 (N_5514,N_1046,N_250);
xnor U5515 (N_5515,N_1273,N_1953);
xor U5516 (N_5516,N_585,N_327);
xor U5517 (N_5517,N_436,N_1534);
nand U5518 (N_5518,N_172,N_2965);
or U5519 (N_5519,N_2243,N_1687);
xor U5520 (N_5520,N_764,N_36);
or U5521 (N_5521,N_1952,N_2596);
or U5522 (N_5522,N_1644,N_270);
nor U5523 (N_5523,N_337,N_2481);
or U5524 (N_5524,N_2563,N_1538);
or U5525 (N_5525,N_359,N_1827);
xnor U5526 (N_5526,N_1498,N_402);
xnor U5527 (N_5527,N_1274,N_1190);
xnor U5528 (N_5528,N_1343,N_1007);
nand U5529 (N_5529,N_1289,N_2262);
xor U5530 (N_5530,N_2934,N_1190);
or U5531 (N_5531,N_2169,N_2135);
nand U5532 (N_5532,N_1159,N_1042);
xor U5533 (N_5533,N_2419,N_2174);
xnor U5534 (N_5534,N_2213,N_875);
and U5535 (N_5535,N_2828,N_255);
and U5536 (N_5536,N_146,N_1481);
and U5537 (N_5537,N_1625,N_1597);
nand U5538 (N_5538,N_2404,N_457);
xor U5539 (N_5539,N_1537,N_2995);
nor U5540 (N_5540,N_381,N_705);
xor U5541 (N_5541,N_1331,N_2323);
nand U5542 (N_5542,N_1442,N_2899);
nand U5543 (N_5543,N_35,N_850);
and U5544 (N_5544,N_260,N_562);
nand U5545 (N_5545,N_1871,N_2797);
and U5546 (N_5546,N_2796,N_962);
nand U5547 (N_5547,N_1593,N_97);
and U5548 (N_5548,N_1543,N_514);
nand U5549 (N_5549,N_206,N_2572);
xor U5550 (N_5550,N_743,N_2854);
nand U5551 (N_5551,N_2737,N_1016);
nand U5552 (N_5552,N_2217,N_2861);
nand U5553 (N_5553,N_827,N_2731);
xnor U5554 (N_5554,N_2013,N_277);
and U5555 (N_5555,N_2639,N_2159);
xnor U5556 (N_5556,N_1198,N_1604);
or U5557 (N_5557,N_233,N_1063);
xnor U5558 (N_5558,N_2033,N_1398);
and U5559 (N_5559,N_2918,N_1370);
xnor U5560 (N_5560,N_143,N_62);
and U5561 (N_5561,N_2291,N_2983);
nor U5562 (N_5562,N_657,N_523);
nor U5563 (N_5563,N_743,N_2498);
nor U5564 (N_5564,N_1165,N_1054);
or U5565 (N_5565,N_350,N_1315);
nand U5566 (N_5566,N_2667,N_1618);
and U5567 (N_5567,N_2254,N_1621);
nand U5568 (N_5568,N_84,N_1136);
nor U5569 (N_5569,N_945,N_107);
nand U5570 (N_5570,N_2689,N_1045);
nand U5571 (N_5571,N_781,N_2329);
nor U5572 (N_5572,N_1443,N_1455);
nor U5573 (N_5573,N_19,N_2852);
nand U5574 (N_5574,N_2927,N_957);
and U5575 (N_5575,N_383,N_1084);
xor U5576 (N_5576,N_2601,N_1863);
and U5577 (N_5577,N_2468,N_207);
xnor U5578 (N_5578,N_1657,N_309);
xor U5579 (N_5579,N_1015,N_561);
xor U5580 (N_5580,N_2833,N_2344);
and U5581 (N_5581,N_1004,N_1011);
nor U5582 (N_5582,N_888,N_1673);
nand U5583 (N_5583,N_181,N_2692);
nor U5584 (N_5584,N_1176,N_516);
or U5585 (N_5585,N_1834,N_2196);
xor U5586 (N_5586,N_127,N_644);
and U5587 (N_5587,N_2045,N_1725);
or U5588 (N_5588,N_2390,N_2498);
and U5589 (N_5589,N_292,N_1885);
nor U5590 (N_5590,N_1563,N_468);
nand U5591 (N_5591,N_1397,N_685);
nor U5592 (N_5592,N_884,N_1555);
nor U5593 (N_5593,N_487,N_2559);
and U5594 (N_5594,N_1278,N_1058);
nor U5595 (N_5595,N_1457,N_1454);
and U5596 (N_5596,N_270,N_1996);
nor U5597 (N_5597,N_821,N_184);
or U5598 (N_5598,N_210,N_2675);
nor U5599 (N_5599,N_692,N_1650);
xor U5600 (N_5600,N_1503,N_2420);
xor U5601 (N_5601,N_1881,N_171);
nand U5602 (N_5602,N_1261,N_1165);
nand U5603 (N_5603,N_954,N_2963);
nand U5604 (N_5604,N_2869,N_1028);
nor U5605 (N_5605,N_2511,N_2669);
nor U5606 (N_5606,N_478,N_1168);
nand U5607 (N_5607,N_2626,N_1967);
nand U5608 (N_5608,N_2363,N_2714);
nand U5609 (N_5609,N_1985,N_2056);
nand U5610 (N_5610,N_1248,N_1765);
nand U5611 (N_5611,N_2812,N_734);
nor U5612 (N_5612,N_1916,N_316);
and U5613 (N_5613,N_796,N_239);
nor U5614 (N_5614,N_66,N_1070);
and U5615 (N_5615,N_2502,N_1241);
nand U5616 (N_5616,N_338,N_2372);
nand U5617 (N_5617,N_1818,N_1476);
and U5618 (N_5618,N_361,N_896);
or U5619 (N_5619,N_1350,N_1923);
nor U5620 (N_5620,N_1615,N_2082);
nand U5621 (N_5621,N_1935,N_269);
and U5622 (N_5622,N_1542,N_549);
or U5623 (N_5623,N_304,N_1061);
nor U5624 (N_5624,N_2111,N_2035);
xor U5625 (N_5625,N_2342,N_836);
and U5626 (N_5626,N_888,N_2754);
or U5627 (N_5627,N_714,N_555);
xor U5628 (N_5628,N_1090,N_1905);
nor U5629 (N_5629,N_1084,N_2168);
and U5630 (N_5630,N_2663,N_2149);
and U5631 (N_5631,N_81,N_1108);
xor U5632 (N_5632,N_328,N_1231);
and U5633 (N_5633,N_1849,N_2968);
nand U5634 (N_5634,N_2304,N_2173);
or U5635 (N_5635,N_846,N_1731);
or U5636 (N_5636,N_870,N_1935);
xor U5637 (N_5637,N_1189,N_1874);
or U5638 (N_5638,N_1600,N_568);
nand U5639 (N_5639,N_2879,N_2269);
or U5640 (N_5640,N_2273,N_2278);
and U5641 (N_5641,N_2201,N_2363);
xor U5642 (N_5642,N_54,N_2957);
and U5643 (N_5643,N_2296,N_2505);
and U5644 (N_5644,N_719,N_2974);
xnor U5645 (N_5645,N_1557,N_1498);
nor U5646 (N_5646,N_2966,N_2471);
nand U5647 (N_5647,N_651,N_2210);
or U5648 (N_5648,N_596,N_1006);
or U5649 (N_5649,N_718,N_1069);
nand U5650 (N_5650,N_2496,N_1457);
xor U5651 (N_5651,N_2092,N_2640);
nand U5652 (N_5652,N_1009,N_2153);
or U5653 (N_5653,N_2377,N_1818);
and U5654 (N_5654,N_1036,N_711);
and U5655 (N_5655,N_2683,N_1983);
and U5656 (N_5656,N_2430,N_1092);
xnor U5657 (N_5657,N_101,N_1367);
or U5658 (N_5658,N_193,N_1533);
xor U5659 (N_5659,N_2266,N_899);
nor U5660 (N_5660,N_2311,N_624);
and U5661 (N_5661,N_676,N_2016);
xor U5662 (N_5662,N_2730,N_2074);
nor U5663 (N_5663,N_940,N_498);
xor U5664 (N_5664,N_1941,N_364);
and U5665 (N_5665,N_976,N_387);
and U5666 (N_5666,N_2548,N_2961);
or U5667 (N_5667,N_778,N_2582);
and U5668 (N_5668,N_1996,N_1544);
xor U5669 (N_5669,N_1892,N_1832);
xnor U5670 (N_5670,N_2332,N_427);
nand U5671 (N_5671,N_1244,N_9);
xor U5672 (N_5672,N_1154,N_2560);
xnor U5673 (N_5673,N_1098,N_2720);
or U5674 (N_5674,N_2444,N_922);
xnor U5675 (N_5675,N_1059,N_2949);
or U5676 (N_5676,N_1790,N_1324);
nor U5677 (N_5677,N_947,N_2209);
nand U5678 (N_5678,N_1180,N_1759);
nand U5679 (N_5679,N_1376,N_2293);
xor U5680 (N_5680,N_2390,N_1483);
and U5681 (N_5681,N_2360,N_1991);
nor U5682 (N_5682,N_1806,N_1005);
and U5683 (N_5683,N_1804,N_2398);
or U5684 (N_5684,N_351,N_511);
nand U5685 (N_5685,N_87,N_2982);
or U5686 (N_5686,N_1524,N_2017);
xnor U5687 (N_5687,N_1377,N_1740);
xnor U5688 (N_5688,N_821,N_2689);
or U5689 (N_5689,N_805,N_1052);
nor U5690 (N_5690,N_2203,N_1313);
nand U5691 (N_5691,N_1187,N_2039);
xor U5692 (N_5692,N_592,N_1541);
or U5693 (N_5693,N_2693,N_2246);
nand U5694 (N_5694,N_2470,N_2461);
and U5695 (N_5695,N_12,N_2434);
nand U5696 (N_5696,N_1758,N_1118);
nand U5697 (N_5697,N_885,N_853);
and U5698 (N_5698,N_2693,N_1488);
and U5699 (N_5699,N_2943,N_1539);
and U5700 (N_5700,N_633,N_1322);
xnor U5701 (N_5701,N_2151,N_1042);
and U5702 (N_5702,N_666,N_1437);
nand U5703 (N_5703,N_1578,N_1681);
nand U5704 (N_5704,N_443,N_1050);
nand U5705 (N_5705,N_2811,N_97);
xnor U5706 (N_5706,N_876,N_2279);
or U5707 (N_5707,N_488,N_2742);
and U5708 (N_5708,N_495,N_2546);
and U5709 (N_5709,N_1727,N_1915);
xnor U5710 (N_5710,N_116,N_1670);
and U5711 (N_5711,N_670,N_494);
or U5712 (N_5712,N_1584,N_2785);
or U5713 (N_5713,N_1414,N_2284);
nand U5714 (N_5714,N_1584,N_850);
and U5715 (N_5715,N_2607,N_1338);
nor U5716 (N_5716,N_2119,N_786);
nor U5717 (N_5717,N_1667,N_1163);
or U5718 (N_5718,N_115,N_2330);
nor U5719 (N_5719,N_1485,N_1599);
or U5720 (N_5720,N_2202,N_963);
or U5721 (N_5721,N_1752,N_1028);
or U5722 (N_5722,N_1163,N_1005);
xor U5723 (N_5723,N_930,N_2118);
xnor U5724 (N_5724,N_2350,N_2980);
xnor U5725 (N_5725,N_2144,N_2246);
or U5726 (N_5726,N_1911,N_938);
nand U5727 (N_5727,N_1258,N_994);
and U5728 (N_5728,N_492,N_2244);
or U5729 (N_5729,N_2709,N_1157);
nor U5730 (N_5730,N_713,N_2907);
or U5731 (N_5731,N_952,N_718);
nand U5732 (N_5732,N_579,N_639);
nor U5733 (N_5733,N_2263,N_216);
or U5734 (N_5734,N_1799,N_1232);
nand U5735 (N_5735,N_1648,N_2774);
or U5736 (N_5736,N_612,N_1711);
nand U5737 (N_5737,N_727,N_111);
nor U5738 (N_5738,N_1449,N_865);
nor U5739 (N_5739,N_607,N_899);
nor U5740 (N_5740,N_1630,N_2175);
xnor U5741 (N_5741,N_309,N_383);
nand U5742 (N_5742,N_1351,N_409);
and U5743 (N_5743,N_2658,N_1496);
and U5744 (N_5744,N_676,N_2811);
and U5745 (N_5745,N_1180,N_1478);
nor U5746 (N_5746,N_1710,N_2991);
and U5747 (N_5747,N_1893,N_1261);
xor U5748 (N_5748,N_1772,N_2457);
and U5749 (N_5749,N_871,N_2083);
and U5750 (N_5750,N_1512,N_113);
and U5751 (N_5751,N_2748,N_269);
xor U5752 (N_5752,N_888,N_2115);
or U5753 (N_5753,N_2465,N_448);
and U5754 (N_5754,N_106,N_2546);
nor U5755 (N_5755,N_1689,N_147);
or U5756 (N_5756,N_1805,N_2489);
xnor U5757 (N_5757,N_974,N_727);
and U5758 (N_5758,N_2018,N_2755);
and U5759 (N_5759,N_2335,N_2423);
and U5760 (N_5760,N_32,N_847);
and U5761 (N_5761,N_835,N_1352);
and U5762 (N_5762,N_1316,N_1908);
and U5763 (N_5763,N_1647,N_1189);
or U5764 (N_5764,N_2080,N_1898);
xnor U5765 (N_5765,N_2268,N_579);
nand U5766 (N_5766,N_1565,N_692);
nor U5767 (N_5767,N_520,N_138);
xor U5768 (N_5768,N_719,N_348);
and U5769 (N_5769,N_1533,N_1078);
and U5770 (N_5770,N_2646,N_2006);
or U5771 (N_5771,N_2440,N_801);
xnor U5772 (N_5772,N_1999,N_1253);
xnor U5773 (N_5773,N_1655,N_2690);
or U5774 (N_5774,N_1643,N_1280);
nand U5775 (N_5775,N_2945,N_2350);
or U5776 (N_5776,N_2876,N_2051);
nand U5777 (N_5777,N_1030,N_2766);
nand U5778 (N_5778,N_921,N_2830);
xor U5779 (N_5779,N_2138,N_576);
xor U5780 (N_5780,N_446,N_1903);
and U5781 (N_5781,N_2661,N_1849);
and U5782 (N_5782,N_2953,N_1640);
nand U5783 (N_5783,N_378,N_1917);
or U5784 (N_5784,N_1219,N_1551);
nand U5785 (N_5785,N_107,N_924);
and U5786 (N_5786,N_1341,N_131);
nand U5787 (N_5787,N_2055,N_958);
xnor U5788 (N_5788,N_1713,N_2504);
or U5789 (N_5789,N_2859,N_1062);
or U5790 (N_5790,N_2845,N_2022);
and U5791 (N_5791,N_556,N_306);
and U5792 (N_5792,N_694,N_780);
and U5793 (N_5793,N_287,N_279);
or U5794 (N_5794,N_2091,N_34);
nand U5795 (N_5795,N_2135,N_292);
nand U5796 (N_5796,N_1000,N_1758);
xor U5797 (N_5797,N_386,N_1612);
or U5798 (N_5798,N_1452,N_2911);
xor U5799 (N_5799,N_1661,N_1531);
nor U5800 (N_5800,N_2722,N_401);
nor U5801 (N_5801,N_2742,N_1941);
or U5802 (N_5802,N_1703,N_200);
or U5803 (N_5803,N_1955,N_2456);
nor U5804 (N_5804,N_1116,N_2203);
xnor U5805 (N_5805,N_40,N_299);
nor U5806 (N_5806,N_1443,N_1681);
and U5807 (N_5807,N_1990,N_781);
and U5808 (N_5808,N_1356,N_2287);
xnor U5809 (N_5809,N_2859,N_2964);
nor U5810 (N_5810,N_65,N_57);
nand U5811 (N_5811,N_2932,N_2995);
or U5812 (N_5812,N_2865,N_555);
and U5813 (N_5813,N_2543,N_1423);
or U5814 (N_5814,N_894,N_2557);
nand U5815 (N_5815,N_2911,N_723);
and U5816 (N_5816,N_2411,N_2457);
and U5817 (N_5817,N_1157,N_2154);
or U5818 (N_5818,N_1292,N_1046);
xor U5819 (N_5819,N_1561,N_2515);
or U5820 (N_5820,N_1519,N_966);
nor U5821 (N_5821,N_1488,N_1066);
nand U5822 (N_5822,N_1491,N_1095);
nor U5823 (N_5823,N_2005,N_983);
nor U5824 (N_5824,N_1672,N_77);
nand U5825 (N_5825,N_947,N_1226);
or U5826 (N_5826,N_99,N_2891);
nor U5827 (N_5827,N_575,N_887);
and U5828 (N_5828,N_2596,N_1310);
xnor U5829 (N_5829,N_2814,N_195);
and U5830 (N_5830,N_2494,N_2008);
and U5831 (N_5831,N_2720,N_1411);
nand U5832 (N_5832,N_580,N_845);
xnor U5833 (N_5833,N_576,N_406);
or U5834 (N_5834,N_432,N_2644);
or U5835 (N_5835,N_631,N_2878);
xnor U5836 (N_5836,N_507,N_1152);
nand U5837 (N_5837,N_2827,N_565);
nor U5838 (N_5838,N_2882,N_680);
nand U5839 (N_5839,N_1229,N_441);
or U5840 (N_5840,N_623,N_1400);
nor U5841 (N_5841,N_1548,N_1590);
nand U5842 (N_5842,N_527,N_37);
xor U5843 (N_5843,N_545,N_1465);
and U5844 (N_5844,N_494,N_312);
nand U5845 (N_5845,N_2843,N_2145);
nor U5846 (N_5846,N_882,N_2530);
xnor U5847 (N_5847,N_1522,N_2401);
or U5848 (N_5848,N_895,N_736);
nor U5849 (N_5849,N_2014,N_199);
xor U5850 (N_5850,N_1527,N_311);
nand U5851 (N_5851,N_1106,N_1583);
nor U5852 (N_5852,N_563,N_2202);
xnor U5853 (N_5853,N_2091,N_545);
or U5854 (N_5854,N_342,N_599);
nor U5855 (N_5855,N_696,N_421);
and U5856 (N_5856,N_1105,N_2615);
nand U5857 (N_5857,N_2461,N_933);
or U5858 (N_5858,N_2266,N_1855);
xor U5859 (N_5859,N_261,N_1471);
nand U5860 (N_5860,N_826,N_1974);
or U5861 (N_5861,N_1756,N_679);
or U5862 (N_5862,N_496,N_1815);
nand U5863 (N_5863,N_2542,N_1382);
and U5864 (N_5864,N_2836,N_317);
or U5865 (N_5865,N_1603,N_51);
xor U5866 (N_5866,N_2790,N_1034);
xor U5867 (N_5867,N_978,N_1484);
xor U5868 (N_5868,N_850,N_474);
nor U5869 (N_5869,N_640,N_1457);
nand U5870 (N_5870,N_640,N_30);
or U5871 (N_5871,N_2989,N_382);
nor U5872 (N_5872,N_1899,N_296);
and U5873 (N_5873,N_1261,N_561);
and U5874 (N_5874,N_475,N_1277);
and U5875 (N_5875,N_1726,N_889);
or U5876 (N_5876,N_2887,N_2761);
xor U5877 (N_5877,N_1060,N_983);
and U5878 (N_5878,N_324,N_1092);
or U5879 (N_5879,N_451,N_429);
nand U5880 (N_5880,N_2477,N_914);
nor U5881 (N_5881,N_924,N_695);
or U5882 (N_5882,N_1529,N_1128);
nand U5883 (N_5883,N_351,N_1120);
nand U5884 (N_5884,N_1373,N_1825);
nand U5885 (N_5885,N_1166,N_2851);
and U5886 (N_5886,N_2188,N_978);
nor U5887 (N_5887,N_2530,N_2119);
xnor U5888 (N_5888,N_2427,N_1869);
nor U5889 (N_5889,N_762,N_1403);
or U5890 (N_5890,N_2650,N_512);
or U5891 (N_5891,N_344,N_262);
or U5892 (N_5892,N_234,N_1690);
xnor U5893 (N_5893,N_2462,N_1018);
nand U5894 (N_5894,N_2238,N_2601);
and U5895 (N_5895,N_331,N_1097);
nor U5896 (N_5896,N_2120,N_1169);
and U5897 (N_5897,N_1470,N_1013);
or U5898 (N_5898,N_1228,N_1368);
or U5899 (N_5899,N_2681,N_2689);
xnor U5900 (N_5900,N_1530,N_1769);
xor U5901 (N_5901,N_923,N_1525);
xnor U5902 (N_5902,N_292,N_428);
xnor U5903 (N_5903,N_576,N_522);
and U5904 (N_5904,N_2842,N_1223);
nor U5905 (N_5905,N_2545,N_2493);
xor U5906 (N_5906,N_766,N_1047);
xnor U5907 (N_5907,N_1513,N_2072);
and U5908 (N_5908,N_405,N_532);
xnor U5909 (N_5909,N_1435,N_526);
nand U5910 (N_5910,N_2986,N_1525);
xnor U5911 (N_5911,N_364,N_1742);
xnor U5912 (N_5912,N_1133,N_2895);
nor U5913 (N_5913,N_2184,N_1306);
nor U5914 (N_5914,N_2884,N_703);
xnor U5915 (N_5915,N_2408,N_121);
or U5916 (N_5916,N_1509,N_790);
xor U5917 (N_5917,N_2503,N_1494);
nor U5918 (N_5918,N_2343,N_630);
or U5919 (N_5919,N_927,N_1981);
nor U5920 (N_5920,N_207,N_2154);
nand U5921 (N_5921,N_2662,N_620);
and U5922 (N_5922,N_1199,N_564);
xor U5923 (N_5923,N_1772,N_158);
or U5924 (N_5924,N_2663,N_72);
and U5925 (N_5925,N_212,N_2936);
and U5926 (N_5926,N_468,N_53);
and U5927 (N_5927,N_2332,N_140);
and U5928 (N_5928,N_413,N_2894);
xnor U5929 (N_5929,N_1221,N_2137);
nor U5930 (N_5930,N_1563,N_1883);
nor U5931 (N_5931,N_652,N_2338);
and U5932 (N_5932,N_2754,N_1698);
nand U5933 (N_5933,N_2005,N_2302);
or U5934 (N_5934,N_2119,N_1383);
xor U5935 (N_5935,N_1320,N_1016);
or U5936 (N_5936,N_2354,N_2393);
xnor U5937 (N_5937,N_723,N_2661);
nand U5938 (N_5938,N_2023,N_38);
nand U5939 (N_5939,N_242,N_2921);
xor U5940 (N_5940,N_2776,N_2213);
or U5941 (N_5941,N_906,N_1388);
nor U5942 (N_5942,N_2442,N_1708);
xor U5943 (N_5943,N_148,N_2038);
nor U5944 (N_5944,N_1673,N_1950);
or U5945 (N_5945,N_337,N_883);
xnor U5946 (N_5946,N_2359,N_469);
or U5947 (N_5947,N_1060,N_1625);
nand U5948 (N_5948,N_775,N_2533);
nor U5949 (N_5949,N_594,N_1719);
nor U5950 (N_5950,N_578,N_2460);
nor U5951 (N_5951,N_1171,N_2790);
nand U5952 (N_5952,N_1834,N_2469);
or U5953 (N_5953,N_863,N_2049);
xor U5954 (N_5954,N_567,N_1805);
xnor U5955 (N_5955,N_2495,N_2797);
and U5956 (N_5956,N_1512,N_1646);
or U5957 (N_5957,N_778,N_327);
nor U5958 (N_5958,N_2344,N_2419);
nor U5959 (N_5959,N_1286,N_629);
nand U5960 (N_5960,N_1709,N_1542);
nand U5961 (N_5961,N_308,N_2798);
and U5962 (N_5962,N_922,N_2587);
xor U5963 (N_5963,N_1414,N_331);
nand U5964 (N_5964,N_2603,N_2483);
nand U5965 (N_5965,N_356,N_2264);
nor U5966 (N_5966,N_19,N_2764);
nand U5967 (N_5967,N_2507,N_2969);
xnor U5968 (N_5968,N_868,N_205);
or U5969 (N_5969,N_104,N_1732);
or U5970 (N_5970,N_903,N_2436);
nor U5971 (N_5971,N_806,N_364);
nand U5972 (N_5972,N_1571,N_2671);
xnor U5973 (N_5973,N_148,N_1788);
and U5974 (N_5974,N_1298,N_2434);
xnor U5975 (N_5975,N_446,N_1080);
nand U5976 (N_5976,N_1460,N_171);
xnor U5977 (N_5977,N_2446,N_2037);
and U5978 (N_5978,N_1211,N_265);
nand U5979 (N_5979,N_2558,N_1589);
and U5980 (N_5980,N_1710,N_2031);
or U5981 (N_5981,N_779,N_2902);
nand U5982 (N_5982,N_1439,N_206);
nor U5983 (N_5983,N_1336,N_1838);
or U5984 (N_5984,N_29,N_1358);
nand U5985 (N_5985,N_382,N_1188);
nand U5986 (N_5986,N_2651,N_492);
and U5987 (N_5987,N_1503,N_1856);
nor U5988 (N_5988,N_1955,N_2712);
xnor U5989 (N_5989,N_2665,N_2216);
xnor U5990 (N_5990,N_1545,N_2411);
nand U5991 (N_5991,N_770,N_1763);
or U5992 (N_5992,N_657,N_2961);
and U5993 (N_5993,N_615,N_2736);
xnor U5994 (N_5994,N_2893,N_1572);
nor U5995 (N_5995,N_2251,N_2381);
and U5996 (N_5996,N_280,N_1032);
or U5997 (N_5997,N_1292,N_58);
nand U5998 (N_5998,N_2069,N_2004);
xor U5999 (N_5999,N_2801,N_1031);
or U6000 (N_6000,N_3110,N_4172);
xor U6001 (N_6001,N_5442,N_3339);
or U6002 (N_6002,N_4528,N_5639);
or U6003 (N_6003,N_3822,N_4268);
and U6004 (N_6004,N_5596,N_5505);
nand U6005 (N_6005,N_3687,N_3338);
or U6006 (N_6006,N_4343,N_3962);
nor U6007 (N_6007,N_3460,N_5806);
xnor U6008 (N_6008,N_5357,N_3375);
nand U6009 (N_6009,N_4787,N_3917);
and U6010 (N_6010,N_5562,N_5075);
or U6011 (N_6011,N_4582,N_3794);
nor U6012 (N_6012,N_5480,N_4157);
xnor U6013 (N_6013,N_5172,N_3480);
and U6014 (N_6014,N_4457,N_3587);
or U6015 (N_6015,N_3040,N_5324);
nand U6016 (N_6016,N_4399,N_5615);
and U6017 (N_6017,N_4694,N_5311);
xor U6018 (N_6018,N_4580,N_5692);
xor U6019 (N_6019,N_3751,N_3087);
and U6020 (N_6020,N_4448,N_4319);
nor U6021 (N_6021,N_5120,N_5927);
nand U6022 (N_6022,N_5429,N_3179);
xnor U6023 (N_6023,N_3564,N_3944);
nor U6024 (N_6024,N_4931,N_3019);
and U6025 (N_6025,N_3972,N_3256);
xor U6026 (N_6026,N_5732,N_3829);
and U6027 (N_6027,N_5059,N_4379);
or U6028 (N_6028,N_3578,N_3346);
nor U6029 (N_6029,N_3837,N_5452);
or U6030 (N_6030,N_5125,N_5537);
nand U6031 (N_6031,N_5568,N_4653);
or U6032 (N_6032,N_4291,N_3580);
nor U6033 (N_6033,N_5550,N_3952);
nand U6034 (N_6034,N_5360,N_4017);
nand U6035 (N_6035,N_4565,N_3327);
nand U6036 (N_6036,N_5974,N_5473);
xnor U6037 (N_6037,N_3843,N_5791);
nor U6038 (N_6038,N_5418,N_5833);
and U6039 (N_6039,N_4733,N_5684);
nand U6040 (N_6040,N_3471,N_3393);
or U6041 (N_6041,N_3558,N_3656);
and U6042 (N_6042,N_4445,N_5467);
nand U6043 (N_6043,N_3693,N_5619);
and U6044 (N_6044,N_5551,N_5618);
xor U6045 (N_6045,N_5033,N_5933);
xnor U6046 (N_6046,N_5738,N_5487);
or U6047 (N_6047,N_3995,N_3918);
xnor U6048 (N_6048,N_3444,N_5877);
or U6049 (N_6049,N_5097,N_5265);
nand U6050 (N_6050,N_3807,N_5001);
xnor U6051 (N_6051,N_4530,N_4654);
or U6052 (N_6052,N_5836,N_5347);
nor U6053 (N_6053,N_4896,N_5016);
nor U6054 (N_6054,N_3386,N_5681);
nand U6055 (N_6055,N_5611,N_3595);
or U6056 (N_6056,N_5542,N_4375);
and U6057 (N_6057,N_3431,N_3536);
xnor U6058 (N_6058,N_4856,N_5175);
nor U6059 (N_6059,N_5346,N_4977);
nand U6060 (N_6060,N_5285,N_3686);
nor U6061 (N_6061,N_3284,N_3163);
and U6062 (N_6062,N_4267,N_4855);
or U6063 (N_6063,N_5525,N_5051);
nor U6064 (N_6064,N_4921,N_5603);
nand U6065 (N_6065,N_3313,N_3806);
and U6066 (N_6066,N_5306,N_4747);
xnor U6067 (N_6067,N_5645,N_5246);
nor U6068 (N_6068,N_3907,N_4161);
nor U6069 (N_6069,N_3482,N_4998);
and U6070 (N_6070,N_4254,N_3382);
xnor U6071 (N_6071,N_3508,N_4119);
or U6072 (N_6072,N_5975,N_5762);
xor U6073 (N_6073,N_5793,N_5412);
nand U6074 (N_6074,N_5401,N_4550);
and U6075 (N_6075,N_3208,N_4970);
xnor U6076 (N_6076,N_4933,N_4926);
nor U6077 (N_6077,N_4667,N_3187);
and U6078 (N_6078,N_4934,N_5581);
nand U6079 (N_6079,N_3452,N_5163);
nand U6080 (N_6080,N_3928,N_4133);
or U6081 (N_6081,N_5516,N_5610);
or U6082 (N_6082,N_4063,N_5041);
or U6083 (N_6083,N_3671,N_3394);
and U6084 (N_6084,N_5432,N_3232);
nor U6085 (N_6085,N_3203,N_4302);
nor U6086 (N_6086,N_3416,N_5068);
nand U6087 (N_6087,N_5902,N_5935);
nand U6088 (N_6088,N_3285,N_4831);
and U6089 (N_6089,N_5155,N_3144);
or U6090 (N_6090,N_3763,N_5392);
nor U6091 (N_6091,N_3152,N_3045);
xor U6092 (N_6092,N_4489,N_4173);
or U6093 (N_6093,N_3505,N_3609);
nor U6094 (N_6094,N_3987,N_3241);
and U6095 (N_6095,N_4630,N_4811);
xor U6096 (N_6096,N_3639,N_3887);
xnor U6097 (N_6097,N_5904,N_5252);
xnor U6098 (N_6098,N_4808,N_3056);
or U6099 (N_6099,N_4591,N_4615);
and U6100 (N_6100,N_3079,N_5850);
xor U6101 (N_6101,N_5636,N_3638);
and U6102 (N_6102,N_4083,N_3511);
or U6103 (N_6103,N_3601,N_4416);
and U6104 (N_6104,N_5954,N_3621);
nor U6105 (N_6105,N_4819,N_3545);
xnor U6106 (N_6106,N_3497,N_4010);
nand U6107 (N_6107,N_4853,N_3903);
or U6108 (N_6108,N_4289,N_5063);
and U6109 (N_6109,N_5803,N_4231);
nor U6110 (N_6110,N_3184,N_4158);
nand U6111 (N_6111,N_3105,N_3640);
nand U6112 (N_6112,N_5647,N_3582);
xnor U6113 (N_6113,N_3757,N_3809);
and U6114 (N_6114,N_3075,N_4164);
xnor U6115 (N_6115,N_3205,N_3661);
nor U6116 (N_6116,N_4942,N_5196);
nand U6117 (N_6117,N_4039,N_4308);
or U6118 (N_6118,N_5188,N_3142);
nand U6119 (N_6119,N_5896,N_5664);
xor U6120 (N_6120,N_4065,N_5190);
or U6121 (N_6121,N_3585,N_3695);
or U6122 (N_6122,N_3438,N_3373);
xnor U6123 (N_6123,N_3466,N_5873);
nor U6124 (N_6124,N_3311,N_3344);
xnor U6125 (N_6125,N_4559,N_5454);
or U6126 (N_6126,N_5272,N_3439);
xnor U6127 (N_6127,N_3857,N_5569);
nor U6128 (N_6128,N_3235,N_5079);
or U6129 (N_6129,N_3780,N_4508);
xnor U6130 (N_6130,N_3930,N_5286);
nor U6131 (N_6131,N_4848,N_5846);
and U6132 (N_6132,N_3989,N_3739);
and U6133 (N_6133,N_4480,N_3157);
nand U6134 (N_6134,N_4219,N_3043);
and U6135 (N_6135,N_5228,N_4908);
and U6136 (N_6136,N_3306,N_4409);
and U6137 (N_6137,N_3145,N_4067);
and U6138 (N_6138,N_3692,N_5049);
xor U6139 (N_6139,N_5410,N_5519);
xnor U6140 (N_6140,N_5866,N_3015);
xor U6141 (N_6141,N_5187,N_3617);
xor U6142 (N_6142,N_3424,N_3769);
and U6143 (N_6143,N_3270,N_3553);
nand U6144 (N_6144,N_4093,N_5340);
or U6145 (N_6145,N_3978,N_3124);
or U6146 (N_6146,N_5184,N_4007);
nand U6147 (N_6147,N_3248,N_5822);
xor U6148 (N_6148,N_3217,N_3421);
nor U6149 (N_6149,N_5817,N_3795);
nor U6150 (N_6150,N_4165,N_3941);
xnor U6151 (N_6151,N_4110,N_5443);
nand U6152 (N_6152,N_5081,N_4042);
nand U6153 (N_6153,N_3588,N_4128);
and U6154 (N_6154,N_4222,N_5250);
nand U6155 (N_6155,N_5703,N_3499);
or U6156 (N_6156,N_4805,N_3598);
and U6157 (N_6157,N_5881,N_3334);
or U6158 (N_6158,N_4506,N_5992);
or U6159 (N_6159,N_3247,N_5457);
nor U6160 (N_6160,N_4206,N_3679);
and U6161 (N_6161,N_5740,N_3834);
and U6162 (N_6162,N_3865,N_4396);
nand U6163 (N_6163,N_4084,N_3914);
nand U6164 (N_6164,N_5310,N_3518);
nor U6165 (N_6165,N_3921,N_3657);
or U6166 (N_6166,N_3026,N_3803);
and U6167 (N_6167,N_4122,N_5751);
nand U6168 (N_6168,N_5594,N_5509);
or U6169 (N_6169,N_5654,N_4973);
and U6170 (N_6170,N_4752,N_5229);
or U6171 (N_6171,N_3817,N_5185);
and U6172 (N_6172,N_5011,N_3959);
and U6173 (N_6173,N_5691,N_5225);
and U6174 (N_6174,N_4835,N_5281);
or U6175 (N_6175,N_4576,N_4452);
and U6176 (N_6176,N_3402,N_3961);
xor U6177 (N_6177,N_3703,N_5783);
nor U6178 (N_6178,N_4186,N_4804);
xor U6179 (N_6179,N_5005,N_4418);
and U6180 (N_6180,N_3141,N_3852);
xnor U6181 (N_6181,N_3747,N_4769);
and U6182 (N_6182,N_4761,N_5157);
and U6183 (N_6183,N_4383,N_5243);
nor U6184 (N_6184,N_4387,N_4721);
nor U6185 (N_6185,N_3008,N_5220);
nor U6186 (N_6186,N_5917,N_4046);
nor U6187 (N_6187,N_4179,N_5165);
or U6188 (N_6188,N_4710,N_3287);
xor U6189 (N_6189,N_5508,N_4767);
and U6190 (N_6190,N_3027,N_4441);
xnor U6191 (N_6191,N_3410,N_4812);
or U6192 (N_6192,N_3396,N_4979);
and U6193 (N_6193,N_3859,N_5990);
nor U6194 (N_6194,N_4311,N_4753);
and U6195 (N_6195,N_3197,N_3006);
nand U6196 (N_6196,N_3167,N_4729);
xor U6197 (N_6197,N_5604,N_3413);
xnor U6198 (N_6198,N_3150,N_5488);
or U6199 (N_6199,N_5029,N_3282);
and U6200 (N_6200,N_5774,N_3533);
and U6201 (N_6201,N_4688,N_5642);
xor U6202 (N_6202,N_5366,N_5109);
nor U6203 (N_6203,N_4913,N_5032);
and U6204 (N_6204,N_4124,N_3674);
and U6205 (N_6205,N_4462,N_3622);
nor U6206 (N_6206,N_3500,N_4583);
or U6207 (N_6207,N_4539,N_4872);
nand U6208 (N_6208,N_3294,N_5458);
or U6209 (N_6209,N_5962,N_3159);
nand U6210 (N_6210,N_4505,N_5658);
xnor U6211 (N_6211,N_3273,N_4339);
or U6212 (N_6212,N_3754,N_5140);
nand U6213 (N_6213,N_3559,N_3155);
nand U6214 (N_6214,N_4703,N_3364);
xor U6215 (N_6215,N_3569,N_4648);
xor U6216 (N_6216,N_5966,N_5119);
and U6217 (N_6217,N_4689,N_4290);
xor U6218 (N_6218,N_3919,N_4572);
or U6219 (N_6219,N_3797,N_3352);
nor U6220 (N_6220,N_4193,N_3435);
xor U6221 (N_6221,N_3690,N_4765);
xor U6222 (N_6222,N_3229,N_5323);
or U6223 (N_6223,N_4672,N_4704);
and U6224 (N_6224,N_3391,N_3618);
nand U6225 (N_6225,N_5160,N_3140);
or U6226 (N_6226,N_4880,N_3745);
or U6227 (N_6227,N_5820,N_3331);
nand U6228 (N_6228,N_5960,N_4148);
nor U6229 (N_6229,N_4235,N_4874);
and U6230 (N_6230,N_3986,N_4044);
nand U6231 (N_6231,N_4213,N_3324);
nand U6232 (N_6232,N_3529,N_5829);
and U6233 (N_6233,N_4365,N_5115);
nor U6234 (N_6234,N_4912,N_4336);
xor U6235 (N_6235,N_5650,N_4300);
nor U6236 (N_6236,N_3672,N_4958);
nor U6237 (N_6237,N_3727,N_5143);
or U6238 (N_6238,N_3860,N_5828);
and U6239 (N_6239,N_4551,N_5223);
nand U6240 (N_6240,N_5199,N_3204);
and U6241 (N_6241,N_5937,N_4952);
xnor U6242 (N_6242,N_5224,N_3997);
nor U6243 (N_6243,N_3554,N_5095);
xor U6244 (N_6244,N_5755,N_3309);
and U6245 (N_6245,N_4001,N_5192);
and U6246 (N_6246,N_4679,N_3746);
xnor U6247 (N_6247,N_5583,N_5775);
or U6248 (N_6248,N_3268,N_4947);
xor U6249 (N_6249,N_5789,N_4734);
nand U6250 (N_6250,N_5781,N_4668);
xor U6251 (N_6251,N_3539,N_4946);
or U6252 (N_6252,N_4281,N_5078);
and U6253 (N_6253,N_4027,N_3355);
or U6254 (N_6254,N_5414,N_3635);
or U6255 (N_6255,N_3428,N_5393);
nand U6256 (N_6256,N_4446,N_4820);
nor U6257 (N_6257,N_5767,N_5816);
and U6258 (N_6258,N_5717,N_5970);
nor U6259 (N_6259,N_4382,N_5276);
or U6260 (N_6260,N_4829,N_4159);
nor U6261 (N_6261,N_4279,N_5133);
and U6262 (N_6262,N_3092,N_5168);
xor U6263 (N_6263,N_3329,N_3243);
or U6264 (N_6264,N_4728,N_5034);
and U6265 (N_6265,N_3960,N_4190);
nand U6266 (N_6266,N_3422,N_5996);
nor U6267 (N_6267,N_3905,N_5908);
or U6268 (N_6268,N_3429,N_4038);
or U6269 (N_6269,N_4184,N_4113);
nand U6270 (N_6270,N_4810,N_3594);
or U6271 (N_6271,N_3362,N_4756);
and U6272 (N_6272,N_3383,N_3648);
or U6273 (N_6273,N_3390,N_5289);
nor U6274 (N_6274,N_4652,N_3090);
xor U6275 (N_6275,N_3081,N_3652);
nand U6276 (N_6276,N_5395,N_3810);
xnor U6277 (N_6277,N_4760,N_5556);
or U6278 (N_6278,N_4871,N_3862);
xor U6279 (N_6279,N_5827,N_4025);
nor U6280 (N_6280,N_3254,N_5823);
and U6281 (N_6281,N_4132,N_4377);
nand U6282 (N_6282,N_4822,N_5154);
or U6283 (N_6283,N_5819,N_3778);
or U6284 (N_6284,N_3567,N_5938);
or U6285 (N_6285,N_3651,N_5858);
xnor U6286 (N_6286,N_3607,N_3550);
or U6287 (N_6287,N_4243,N_4090);
nand U6288 (N_6288,N_4833,N_3634);
or U6289 (N_6289,N_3670,N_5061);
nor U6290 (N_6290,N_4229,N_3713);
nor U6291 (N_6291,N_3450,N_5560);
or U6292 (N_6292,N_5065,N_3946);
nand U6293 (N_6293,N_5318,N_3073);
nor U6294 (N_6294,N_5054,N_3784);
or U6295 (N_6295,N_4324,N_4949);
nor U6296 (N_6296,N_5446,N_5646);
nand U6297 (N_6297,N_5624,N_3602);
nand U6298 (N_6298,N_5589,N_3117);
and U6299 (N_6299,N_3964,N_3202);
nor U6300 (N_6300,N_3504,N_4023);
xor U6301 (N_6301,N_3789,N_4274);
xnor U6302 (N_6302,N_3246,N_5719);
nor U6303 (N_6303,N_3283,N_4455);
and U6304 (N_6304,N_4209,N_4500);
xnor U6305 (N_6305,N_3908,N_5936);
nor U6306 (N_6306,N_3631,N_3696);
and U6307 (N_6307,N_5530,N_4350);
nor U6308 (N_6308,N_4002,N_3792);
and U6309 (N_6309,N_3178,N_3351);
nor U6310 (N_6310,N_3341,N_4182);
nor U6311 (N_6311,N_4656,N_3082);
xnor U6312 (N_6312,N_4537,N_5338);
xnor U6313 (N_6313,N_3615,N_3024);
or U6314 (N_6314,N_5352,N_4304);
nand U6315 (N_6315,N_5251,N_3174);
or U6316 (N_6316,N_4072,N_5471);
or U6317 (N_6317,N_5675,N_4830);
and U6318 (N_6318,N_5815,N_5290);
xor U6319 (N_6319,N_5574,N_5930);
nor U6320 (N_6320,N_4873,N_5267);
xnor U6321 (N_6321,N_3872,N_4482);
nand U6322 (N_6322,N_5763,N_4696);
xnor U6323 (N_6323,N_5907,N_5475);
or U6324 (N_6324,N_3733,N_5745);
and U6325 (N_6325,N_5279,N_5137);
nor U6326 (N_6326,N_3328,N_3719);
nor U6327 (N_6327,N_3314,N_4902);
and U6328 (N_6328,N_5756,N_4707);
and U6329 (N_6329,N_4204,N_4601);
or U6330 (N_6330,N_3994,N_3787);
nor U6331 (N_6331,N_5439,N_5230);
and U6332 (N_6332,N_5300,N_4437);
nand U6333 (N_6333,N_3199,N_3227);
nor U6334 (N_6334,N_4863,N_5420);
and U6335 (N_6335,N_4955,N_5538);
nor U6336 (N_6336,N_3377,N_5649);
xnor U6337 (N_6337,N_5247,N_4192);
or U6338 (N_6338,N_5351,N_4363);
nor U6339 (N_6339,N_4599,N_3212);
nor U6340 (N_6340,N_4661,N_4139);
nor U6341 (N_6341,N_4659,N_3293);
nor U6342 (N_6342,N_4348,N_4087);
and U6343 (N_6343,N_5812,N_5784);
or U6344 (N_6344,N_3401,N_5811);
nand U6345 (N_6345,N_4251,N_4813);
xor U6346 (N_6346,N_3704,N_5129);
or U6347 (N_6347,N_5824,N_5678);
nand U6348 (N_6348,N_4684,N_3723);
and U6349 (N_6349,N_3625,N_4643);
nand U6350 (N_6350,N_3737,N_5561);
or U6351 (N_6351,N_5106,N_5606);
nand U6352 (N_6352,N_3762,N_3158);
nand U6353 (N_6353,N_4378,N_5999);
nor U6354 (N_6354,N_3104,N_4356);
nand U6355 (N_6355,N_3552,N_4012);
xor U6356 (N_6356,N_4344,N_5534);
and U6357 (N_6357,N_3534,N_3400);
xnor U6358 (N_6358,N_3649,N_4837);
and U6359 (N_6359,N_5128,N_4494);
or U6360 (N_6360,N_4341,N_5727);
nor U6361 (N_6361,N_5768,N_3688);
nand U6362 (N_6362,N_3376,N_3201);
nand U6363 (N_6363,N_5808,N_5942);
or U6364 (N_6364,N_4675,N_4015);
nor U6365 (N_6365,N_5659,N_3035);
nor U6366 (N_6366,N_5166,N_4697);
and U6367 (N_6367,N_3211,N_3074);
nand U6368 (N_6368,N_5386,N_3219);
nor U6369 (N_6369,N_3221,N_4359);
nand U6370 (N_6370,N_5734,N_5474);
nand U6371 (N_6371,N_3838,N_3280);
nand U6372 (N_6372,N_4030,N_5102);
nor U6373 (N_6373,N_3419,N_3708);
and U6374 (N_6374,N_3985,N_5069);
nor U6375 (N_6375,N_5046,N_4784);
and U6376 (N_6376,N_3893,N_5441);
xnor U6377 (N_6377,N_4980,N_5814);
and U6378 (N_6378,N_4868,N_4748);
xnor U6379 (N_6379,N_4658,N_4419);
or U6380 (N_6380,N_4791,N_4212);
and U6381 (N_6381,N_3374,N_4996);
xor U6382 (N_6382,N_5067,N_5098);
xnor U6383 (N_6383,N_5946,N_5022);
and U6384 (N_6384,N_5771,N_4900);
and U6385 (N_6385,N_5979,N_3705);
nor U6386 (N_6386,N_5421,N_5609);
xor U6387 (N_6387,N_4466,N_4162);
nand U6388 (N_6388,N_4968,N_3927);
xnor U6389 (N_6389,N_3732,N_5982);
or U6390 (N_6390,N_5482,N_3593);
and U6391 (N_6391,N_3775,N_4285);
nand U6392 (N_6392,N_4080,N_4320);
nor U6393 (N_6393,N_4282,N_5437);
xor U6394 (N_6394,N_3108,N_5014);
nand U6395 (N_6395,N_3023,N_5950);
and U6396 (N_6396,N_4687,N_5219);
nor U6397 (N_6397,N_3522,N_4497);
nand U6398 (N_6398,N_4956,N_5991);
xor U6399 (N_6399,N_4841,N_4226);
and U6400 (N_6400,N_5752,N_4994);
and U6401 (N_6401,N_3408,N_3999);
or U6402 (N_6402,N_4496,N_3236);
nand U6403 (N_6403,N_4107,N_4532);
xor U6404 (N_6404,N_5852,N_5124);
and U6405 (N_6405,N_5345,N_5264);
and U6406 (N_6406,N_3387,N_3849);
xor U6407 (N_6407,N_5632,N_4013);
or U6408 (N_6408,N_4925,N_5723);
xor U6409 (N_6409,N_4138,N_5579);
or U6410 (N_6410,N_3209,N_3059);
xor U6411 (N_6411,N_5660,N_3641);
nand U6412 (N_6412,N_3646,N_3911);
xnor U6413 (N_6413,N_4031,N_5683);
nand U6414 (N_6414,N_3901,N_4623);
nand U6415 (N_6415,N_3425,N_5704);
and U6416 (N_6416,N_4376,N_4858);
nand U6417 (N_6417,N_4847,N_4217);
and U6418 (N_6418,N_3031,N_5030);
and U6419 (N_6419,N_5100,N_5799);
nor U6420 (N_6420,N_5073,N_3654);
xnor U6421 (N_6421,N_4775,N_4111);
nand U6422 (N_6422,N_5070,N_4669);
nand U6423 (N_6423,N_5554,N_3537);
xnor U6424 (N_6424,N_3766,N_3094);
and U6425 (N_6425,N_3194,N_5263);
nor U6426 (N_6426,N_4789,N_5709);
nand U6427 (N_6427,N_4590,N_5880);
nand U6428 (N_6428,N_5080,N_3397);
or U6429 (N_6429,N_4008,N_5641);
nand U6430 (N_6430,N_3895,N_5389);
xor U6431 (N_6431,N_3028,N_4857);
or U6432 (N_6432,N_5552,N_4678);
or U6433 (N_6433,N_4258,N_4272);
nand U6434 (N_6434,N_5766,N_5411);
xor U6435 (N_6435,N_4470,N_4066);
nor U6436 (N_6436,N_3575,N_3047);
or U6437 (N_6437,N_5909,N_5456);
xnor U6438 (N_6438,N_5677,N_4892);
or U6439 (N_6439,N_3488,N_4930);
and U6440 (N_6440,N_3619,N_5177);
nor U6441 (N_6441,N_5695,N_3321);
nand U6442 (N_6442,N_3561,N_4169);
xnor U6443 (N_6443,N_5234,N_4726);
nor U6444 (N_6444,N_5330,N_5708);
and U6445 (N_6445,N_4467,N_3451);
or U6446 (N_6446,N_3811,N_4766);
and U6447 (N_6447,N_5644,N_4384);
and U6448 (N_6448,N_5674,N_4944);
nor U6449 (N_6449,N_3170,N_5667);
nand U6450 (N_6450,N_3207,N_5301);
nand U6451 (N_6451,N_5179,N_3523);
xnor U6452 (N_6452,N_3267,N_4032);
nand U6453 (N_6453,N_4657,N_5914);
nand U6454 (N_6454,N_5287,N_4064);
or U6455 (N_6455,N_4711,N_3096);
xor U6456 (N_6456,N_5787,N_5919);
xor U6457 (N_6457,N_5720,N_4545);
nor U6458 (N_6458,N_4163,N_4420);
nor U6459 (N_6459,N_4298,N_4269);
nand U6460 (N_6460,N_4589,N_5668);
or U6461 (N_6461,N_5331,N_3065);
nand U6462 (N_6462,N_3604,N_4230);
nand U6463 (N_6463,N_4417,N_4567);
or U6464 (N_6464,N_5628,N_4102);
nor U6465 (N_6465,N_3667,N_4620);
or U6466 (N_6466,N_3813,N_5744);
and U6467 (N_6467,N_4909,N_5132);
and U6468 (N_6468,N_3098,N_4708);
and U6469 (N_6469,N_4168,N_5580);
or U6470 (N_6470,N_4743,N_4649);
nand U6471 (N_6471,N_4089,N_4883);
xor U6472 (N_6472,N_4296,N_5350);
or U6473 (N_6473,N_5159,N_5705);
nor U6474 (N_6474,N_4088,N_4690);
nand U6475 (N_6475,N_4614,N_3304);
and U6476 (N_6476,N_4585,N_4788);
xnor U6477 (N_6477,N_5375,N_4331);
xor U6478 (N_6478,N_3061,N_3126);
nor U6479 (N_6479,N_5321,N_5447);
or U6480 (N_6480,N_4076,N_5094);
xor U6481 (N_6481,N_5540,N_4610);
nor U6482 (N_6482,N_5653,N_5316);
or U6483 (N_6483,N_5216,N_4422);
nor U6484 (N_6484,N_3965,N_5385);
and U6485 (N_6485,N_5248,N_3606);
nand U6486 (N_6486,N_5558,N_5566);
nor U6487 (N_6487,N_5592,N_5277);
and U6488 (N_6488,N_3274,N_5804);
nand U6489 (N_6489,N_4862,N_4504);
xnor U6490 (N_6490,N_5087,N_3278);
and U6491 (N_6491,N_5138,N_5058);
or U6492 (N_6492,N_5890,N_4962);
and U6493 (N_6493,N_5209,N_4569);
nand U6494 (N_6494,N_4408,N_5736);
and U6495 (N_6495,N_3399,N_5004);
nand U6496 (N_6496,N_3916,N_3876);
xor U6497 (N_6497,N_3469,N_5655);
or U6498 (N_6498,N_5494,N_4197);
or U6499 (N_6499,N_5012,N_5213);
or U6500 (N_6500,N_3748,N_5912);
nor U6501 (N_6501,N_5969,N_4779);
nor U6502 (N_6502,N_5964,N_3509);
and U6503 (N_6503,N_5661,N_5498);
nand U6504 (N_6504,N_4861,N_4412);
and U6505 (N_6505,N_5370,N_4793);
nand U6506 (N_6506,N_3562,N_5490);
nand U6507 (N_6507,N_4778,N_4625);
nand U6508 (N_6508,N_3353,N_4402);
or U6509 (N_6509,N_5593,N_4199);
nor U6510 (N_6510,N_5202,N_4995);
or U6511 (N_6511,N_4520,N_5894);
nor U6512 (N_6512,N_3501,N_4203);
nand U6513 (N_6513,N_4893,N_5131);
nand U6514 (N_6514,N_4593,N_4922);
and U6515 (N_6515,N_4233,N_5888);
xor U6516 (N_6516,N_3642,N_4056);
nor U6517 (N_6517,N_3835,N_4535);
and U6518 (N_6518,N_3326,N_4105);
and U6519 (N_6519,N_5024,N_3468);
xor U6520 (N_6520,N_4509,N_5780);
nand U6521 (N_6521,N_5015,N_5754);
nand U6522 (N_6522,N_5210,N_4176);
xnor U6523 (N_6523,N_5472,N_4626);
or U6524 (N_6524,N_3525,N_5354);
xor U6525 (N_6525,N_4003,N_5423);
xor U6526 (N_6526,N_5895,N_3894);
and U6527 (N_6527,N_5634,N_5008);
nor U6528 (N_6528,N_4353,N_5368);
nor U6529 (N_6529,N_3049,N_5786);
xnor U6530 (N_6530,N_5023,N_4940);
or U6531 (N_6531,N_5725,N_5391);
or U6532 (N_6532,N_5548,N_5260);
and U6533 (N_6533,N_4096,N_4058);
nor U6534 (N_6534,N_3867,N_5963);
and U6535 (N_6535,N_5597,N_5813);
nand U6536 (N_6536,N_4034,N_3255);
xnor U6537 (N_6537,N_5961,N_5397);
and U6538 (N_6538,N_3442,N_4214);
xnor U6539 (N_6539,N_3407,N_4510);
xnor U6540 (N_6540,N_4877,N_4759);
xnor U6541 (N_6541,N_5564,N_3771);
or U6542 (N_6542,N_4638,N_3725);
xor U6543 (N_6543,N_4011,N_4352);
nor U6544 (N_6544,N_5953,N_4531);
nand U6545 (N_6545,N_3953,N_5303);
or U6546 (N_6546,N_5503,N_4048);
and U6547 (N_6547,N_4121,N_3086);
and U6548 (N_6548,N_3070,N_3405);
or U6549 (N_6549,N_4112,N_4646);
or U6550 (N_6550,N_5344,N_5257);
nor U6551 (N_6551,N_5320,N_4373);
or U6552 (N_6552,N_4629,N_3741);
nand U6553 (N_6553,N_3779,N_5702);
or U6554 (N_6554,N_3540,N_3447);
nor U6555 (N_6555,N_4981,N_3939);
and U6556 (N_6556,N_3519,N_4882);
or U6557 (N_6557,N_3669,N_3138);
or U6558 (N_6558,N_5268,N_4337);
nand U6559 (N_6559,N_3276,N_5750);
nor U6560 (N_6560,N_5461,N_3166);
nand U6561 (N_6561,N_4818,N_4957);
nand U6562 (N_6562,N_4205,N_5088);
nor U6563 (N_6563,N_3557,N_3234);
or U6564 (N_6564,N_4181,N_3744);
and U6565 (N_6565,N_4553,N_4501);
nor U6566 (N_6566,N_4828,N_3574);
nand U6567 (N_6567,N_5334,N_3330);
or U6568 (N_6568,N_5152,N_4987);
xnor U6569 (N_6569,N_4665,N_5524);
xor U6570 (N_6570,N_5835,N_5685);
and U6571 (N_6571,N_5801,N_4425);
xor U6572 (N_6572,N_5770,N_3764);
nand U6573 (N_6573,N_4366,N_3804);
nor U6574 (N_6574,N_5591,N_3812);
or U6575 (N_6575,N_5863,N_5772);
xor U6576 (N_6576,N_4109,N_3682);
or U6577 (N_6577,N_5864,N_4836);
and U6578 (N_6578,N_5139,N_4634);
and U6579 (N_6579,N_5275,N_4680);
xor U6580 (N_6580,N_5066,N_5342);
and U6581 (N_6581,N_4511,N_3967);
nor U6582 (N_6582,N_3343,N_4389);
or U6583 (N_6583,N_3128,N_3160);
nor U6584 (N_6584,N_3636,N_5361);
nor U6585 (N_6585,N_5531,N_4471);
nor U6586 (N_6586,N_4195,N_3620);
nand U6587 (N_6587,N_5502,N_3563);
and U6588 (N_6588,N_4318,N_4283);
nand U6589 (N_6589,N_4777,N_3710);
xor U6590 (N_6590,N_3542,N_5007);
nor U6591 (N_6591,N_5897,N_5818);
and U6592 (N_6592,N_4476,N_4305);
nand U6593 (N_6593,N_5565,N_4604);
xnor U6594 (N_6594,N_4491,N_4976);
and U6595 (N_6595,N_5925,N_5924);
nand U6596 (N_6596,N_4000,N_3003);
nor U6597 (N_6597,N_3434,N_5957);
nand U6598 (N_6598,N_5071,N_4938);
xor U6599 (N_6599,N_5795,N_5200);
and U6600 (N_6600,N_5453,N_3067);
nand U6601 (N_6601,N_3066,N_5686);
or U6602 (N_6602,N_4252,N_5497);
nand U6603 (N_6603,N_5955,N_3963);
nor U6604 (N_6604,N_3161,N_3038);
and U6605 (N_6605,N_3955,N_5359);
nand U6606 (N_6606,N_4499,N_4347);
nand U6607 (N_6607,N_4033,N_4587);
nor U6608 (N_6608,N_5096,N_3464);
nor U6609 (N_6609,N_4763,N_5117);
and U6610 (N_6610,N_4685,N_3206);
nand U6611 (N_6611,N_5557,N_4662);
xnor U6612 (N_6612,N_5884,N_5869);
nor U6613 (N_6613,N_3951,N_3685);
xnor U6614 (N_6614,N_4240,N_3699);
or U6615 (N_6615,N_3080,N_5878);
and U6616 (N_6616,N_4988,N_5500);
xor U6617 (N_6617,N_4218,N_3418);
nor U6618 (N_6618,N_3627,N_5578);
xor U6619 (N_6619,N_5616,N_3802);
and U6620 (N_6620,N_4238,N_5572);
or U6621 (N_6621,N_4727,N_3898);
or U6622 (N_6622,N_3189,N_5782);
or U6623 (N_6623,N_5204,N_3583);
and U6624 (N_6624,N_4519,N_4732);
or U6625 (N_6625,N_4415,N_4709);
nand U6626 (N_6626,N_5319,N_4421);
xor U6627 (N_6627,N_5178,N_3350);
nor U6628 (N_6628,N_4594,N_4737);
or U6629 (N_6629,N_4566,N_3915);
or U6630 (N_6630,N_5906,N_3643);
or U6631 (N_6631,N_4906,N_4832);
and U6632 (N_6632,N_4189,N_4449);
xor U6633 (N_6633,N_3077,N_4198);
or U6634 (N_6634,N_4091,N_5167);
or U6635 (N_6635,N_5036,N_5620);
and U6636 (N_6636,N_5180,N_4432);
and U6637 (N_6637,N_5796,N_5476);
xnor U6638 (N_6638,N_5026,N_4160);
and U6639 (N_6639,N_5341,N_3153);
and U6640 (N_6640,N_4540,N_4194);
xnor U6641 (N_6641,N_4866,N_5273);
and U6642 (N_6642,N_3758,N_4796);
or U6643 (N_6643,N_4349,N_3181);
nand U6644 (N_6644,N_3808,N_3659);
nand U6645 (N_6645,N_4859,N_3379);
nand U6646 (N_6646,N_4472,N_4237);
nand U6647 (N_6647,N_3291,N_4749);
xor U6648 (N_6648,N_3934,N_4698);
and U6649 (N_6649,N_3465,N_3029);
nor U6650 (N_6650,N_5424,N_4114);
nand U6651 (N_6651,N_3357,N_3281);
and U6652 (N_6652,N_5637,N_4809);
nand U6653 (N_6653,N_5194,N_3702);
and U6654 (N_6654,N_4256,N_4923);
nor U6655 (N_6655,N_4651,N_3531);
nand U6656 (N_6656,N_4406,N_4975);
or U6657 (N_6657,N_5269,N_4071);
or U6658 (N_6658,N_4242,N_3337);
nor U6659 (N_6659,N_4022,N_4936);
nor U6660 (N_6660,N_3738,N_4963);
nand U6661 (N_6661,N_5515,N_5055);
xnor U6662 (N_6662,N_4024,N_4562);
and U6663 (N_6663,N_5425,N_5746);
nor U6664 (N_6664,N_3544,N_3292);
or U6665 (N_6665,N_4959,N_3629);
and U6666 (N_6666,N_3890,N_5309);
nor U6667 (N_6667,N_4380,N_3022);
nand U6668 (N_6668,N_3814,N_3191);
or U6669 (N_6669,N_4745,N_4322);
or U6670 (N_6670,N_4277,N_5976);
and U6671 (N_6671,N_5212,N_4953);
nor U6672 (N_6672,N_5249,N_5536);
nor U6673 (N_6673,N_5528,N_3507);
nand U6674 (N_6674,N_3180,N_3121);
xor U6675 (N_6675,N_4321,N_4068);
nor U6676 (N_6676,N_4674,N_5355);
xor U6677 (N_6677,N_5983,N_4681);
nor U6678 (N_6678,N_5769,N_3240);
nand U6679 (N_6679,N_4911,N_4262);
or U6680 (N_6680,N_5690,N_4965);
or U6681 (N_6681,N_4473,N_5047);
nand U6682 (N_6682,N_3009,N_3437);
xor U6683 (N_6683,N_4826,N_3251);
nand U6684 (N_6684,N_3665,N_3215);
xor U6685 (N_6685,N_5892,N_5003);
xor U6686 (N_6686,N_5843,N_4478);
xnor U6687 (N_6687,N_3520,N_4079);
nand U6688 (N_6688,N_4081,N_4786);
nor U6689 (N_6689,N_4991,N_4392);
and U6690 (N_6690,N_5875,N_4723);
and U6691 (N_6691,N_5173,N_5266);
or U6692 (N_6692,N_5887,N_5009);
nand U6693 (N_6693,N_4573,N_3632);
nor U6694 (N_6694,N_5838,N_3112);
or U6695 (N_6695,N_4487,N_3445);
and U6696 (N_6696,N_4525,N_5761);
or U6697 (N_6697,N_4405,N_5805);
nor U6698 (N_6698,N_4803,N_4621);
xor U6699 (N_6699,N_4884,N_4202);
nor U6700 (N_6700,N_3164,N_3454);
nand U6701 (N_6701,N_5122,N_4750);
or U6702 (N_6702,N_3380,N_3913);
nor U6703 (N_6703,N_5031,N_4918);
xor U6704 (N_6704,N_3981,N_3000);
nor U6705 (N_6705,N_3259,N_5995);
nand U6706 (N_6706,N_3143,N_5092);
or U6707 (N_6707,N_4307,N_5282);
nand U6708 (N_6708,N_5270,N_4660);
and U6709 (N_6709,N_4800,N_5136);
and U6710 (N_6710,N_5911,N_3245);
xor U6711 (N_6711,N_3900,N_5899);
nand U6712 (N_6712,N_5062,N_4411);
nand U6713 (N_6713,N_3973,N_4622);
nand U6714 (N_6714,N_5084,N_5701);
or U6715 (N_6715,N_3877,N_3122);
xnor U6716 (N_6716,N_5294,N_3146);
or U6717 (N_6717,N_5688,N_5757);
and U6718 (N_6718,N_3071,N_5956);
nand U6719 (N_6719,N_3459,N_3171);
nand U6720 (N_6720,N_4313,N_4150);
xor U6721 (N_6721,N_3177,N_3185);
xnor U6722 (N_6722,N_4507,N_3947);
nand U6723 (N_6723,N_5083,N_4433);
nand U6724 (N_6724,N_3717,N_3225);
nand U6725 (N_6725,N_4887,N_3840);
and U6726 (N_6726,N_3319,N_3060);
nand U6727 (N_6727,N_4639,N_4574);
nand U6728 (N_6728,N_4641,N_5918);
xnor U6729 (N_6729,N_3224,N_5987);
nand U6730 (N_6730,N_3712,N_5586);
xor U6731 (N_6731,N_5127,N_4677);
and U6732 (N_6732,N_3198,N_5356);
xor U6733 (N_6733,N_5623,N_4309);
nor U6734 (N_6734,N_3524,N_5399);
nor U6735 (N_6735,N_4702,N_4029);
or U6736 (N_6736,N_4670,N_3005);
nor U6737 (N_6737,N_5737,N_4864);
nor U6738 (N_6738,N_5240,N_4450);
and U6739 (N_6739,N_3546,N_5479);
or U6740 (N_6740,N_5765,N_3312);
nor U6741 (N_6741,N_3770,N_5753);
xnor U6742 (N_6742,N_3776,N_4345);
or U6743 (N_6743,N_4327,N_5086);
or U6744 (N_6744,N_3348,N_5495);
nor U6745 (N_6745,N_5025,N_4171);
nand U6746 (N_6746,N_4954,N_4293);
and U6747 (N_6747,N_5394,N_5326);
nand U6748 (N_6748,N_3756,N_3154);
xnor U6749 (N_6749,N_4435,N_5147);
xnor U6750 (N_6750,N_3368,N_3214);
or U6751 (N_6751,N_5697,N_5121);
nand U6752 (N_6752,N_3586,N_4407);
or U6753 (N_6753,N_4236,N_3261);
nor U6754 (N_6754,N_3885,N_4891);
xnor U6755 (N_6755,N_4317,N_4261);
nor U6756 (N_6756,N_5107,N_3740);
or U6757 (N_6757,N_3301,N_4577);
or U6758 (N_6758,N_4842,N_5327);
nor U6759 (N_6759,N_5759,N_4554);
xnor U6760 (N_6760,N_4468,N_5253);
nand U6761 (N_6761,N_3816,N_5680);
nor U6762 (N_6762,N_5037,N_4596);
nand U6763 (N_6763,N_4586,N_3316);
xnor U6764 (N_6764,N_3735,N_5170);
and U6765 (N_6765,N_3663,N_4722);
nand U6766 (N_6766,N_4117,N_3743);
nor U6767 (N_6767,N_5130,N_4428);
or U6768 (N_6768,N_4635,N_3495);
nor U6769 (N_6769,N_3440,N_4253);
xnor U6770 (N_6770,N_3018,N_4974);
nor U6771 (N_6771,N_3998,N_4401);
xor U6772 (N_6772,N_3866,N_3992);
or U6773 (N_6773,N_4901,N_3100);
or U6774 (N_6774,N_5978,N_4137);
or U6775 (N_6775,N_4640,N_3868);
xnor U6776 (N_6776,N_5231,N_5629);
nor U6777 (N_6777,N_3231,N_5191);
or U6778 (N_6778,N_3372,N_3931);
or U6779 (N_6779,N_3384,N_3839);
xor U6780 (N_6780,N_5459,N_5052);
xnor U6781 (N_6781,N_3230,N_5682);
xnor U6782 (N_6782,N_3490,N_3091);
and U6783 (N_6783,N_4783,N_5000);
or U6784 (N_6784,N_5042,N_5535);
xor U6785 (N_6785,N_3369,N_5913);
nor U6786 (N_6786,N_3472,N_3423);
xor U6787 (N_6787,N_5056,N_4972);
nand U6788 (N_6788,N_5706,N_4082);
xnor U6789 (N_6789,N_5072,N_3021);
xor U6790 (N_6790,N_5810,N_4724);
and U6791 (N_6791,N_3793,N_4984);
xor U6792 (N_6792,N_5716,N_5463);
nor U6793 (N_6793,N_4568,N_4718);
and U6794 (N_6794,N_3449,N_4983);
nand U6795 (N_6795,N_4438,N_5718);
or U6796 (N_6796,N_3759,N_3644);
nand U6797 (N_6797,N_4292,N_3315);
xor U6798 (N_6798,N_4286,N_4328);
nand U6799 (N_6799,N_3173,N_3749);
or U6800 (N_6800,N_3614,N_4578);
or U6801 (N_6801,N_3768,N_3370);
and U6802 (N_6802,N_4790,N_3791);
xor U6803 (N_6803,N_3922,N_4780);
or U6804 (N_6804,N_4521,N_5337);
nand U6805 (N_6805,N_5236,N_3411);
nor U6806 (N_6806,N_5362,N_4990);
nor U6807 (N_6807,N_4014,N_5466);
and U6808 (N_6808,N_4579,N_3134);
nor U6809 (N_6809,N_3076,N_5112);
nand U6810 (N_6810,N_3136,N_3596);
xnor U6811 (N_6811,N_5872,N_3361);
xor U6812 (N_6812,N_4999,N_4776);
or U6813 (N_6813,N_5156,N_4581);
xor U6814 (N_6814,N_4802,N_5460);
xor U6815 (N_6815,N_3929,N_4095);
nand U6816 (N_6816,N_5948,N_4762);
nor U6817 (N_6817,N_3731,N_5903);
xor U6818 (N_6818,N_3902,N_5141);
or U6819 (N_6819,N_5943,N_3513);
or U6820 (N_6820,N_4917,N_4004);
nor U6821 (N_6821,N_4663,N_5045);
or U6822 (N_6822,N_4143,N_3186);
nor U6823 (N_6823,N_3305,N_4469);
or U6824 (N_6824,N_5207,N_3730);
nand U6825 (N_6825,N_4888,N_3755);
or U6826 (N_6826,N_3645,N_4644);
and U6827 (N_6827,N_5602,N_5889);
and U6828 (N_6828,N_3752,N_5730);
nand U6829 (N_6829,N_4155,N_4706);
nor U6830 (N_6830,N_5436,N_5587);
or U6831 (N_6831,N_3660,N_5567);
and U6832 (N_6832,N_5237,N_3237);
nand U6833 (N_6833,N_4486,N_3935);
and U6834 (N_6834,N_5091,N_3481);
and U6835 (N_6835,N_3566,N_3881);
and U6836 (N_6836,N_3286,N_3874);
xor U6837 (N_6837,N_4314,N_5940);
xnor U6838 (N_6838,N_5484,N_5278);
nand U6839 (N_6839,N_4939,N_4773);
xor U6840 (N_6840,N_4794,N_3068);
xor U6841 (N_6841,N_3183,N_4598);
nor U6842 (N_6842,N_5865,N_5440);
and U6843 (N_6843,N_4515,N_5501);
and U6844 (N_6844,N_5217,N_5742);
and U6845 (N_6845,N_3453,N_5377);
or U6846 (N_6846,N_5074,N_5485);
nand U6847 (N_6847,N_4951,N_3014);
and U6848 (N_6848,N_5193,N_4919);
nor U6849 (N_6849,N_5977,N_5040);
nand U6850 (N_6850,N_4054,N_5932);
nor U6851 (N_6851,N_3033,N_3841);
nor U6852 (N_6852,N_5293,N_5339);
nor U6853 (N_6853,N_3532,N_4127);
nand U6854 (N_6854,N_4897,N_3937);
xnor U6855 (N_6855,N_4484,N_5292);
and U6856 (N_6856,N_3680,N_4126);
or U6857 (N_6857,N_5809,N_5665);
nand U6858 (N_6858,N_5222,N_5855);
xor U6859 (N_6859,N_3815,N_5673);
and U6860 (N_6860,N_5384,N_4323);
nand U6861 (N_6861,N_3782,N_4021);
nand U6862 (N_6862,N_3673,N_5547);
xor U6863 (N_6863,N_4993,N_4603);
xor U6864 (N_6864,N_4522,N_5039);
and U6865 (N_6865,N_3116,N_4595);
nor U6866 (N_6866,N_4686,N_4611);
nand U6867 (N_6867,N_3605,N_5798);
nor U6868 (N_6868,N_3677,N_3020);
xnor U6869 (N_6869,N_3530,N_3427);
nor U6870 (N_6870,N_4315,N_4937);
xnor U6871 (N_6871,N_3783,N_4717);
xnor U6872 (N_6872,N_5959,N_4174);
or U6873 (N_6873,N_4271,N_4541);
and U6874 (N_6874,N_5853,N_4560);
and U6875 (N_6875,N_5048,N_4255);
and U6876 (N_6876,N_3878,N_4374);
xor U6877 (N_6877,N_4390,N_5396);
nor U6878 (N_6878,N_4440,N_4059);
nor U6879 (N_6879,N_5020,N_4633);
nand U6880 (N_6880,N_5158,N_5111);
nand U6881 (N_6881,N_4092,N_3502);
nor U6882 (N_6882,N_5886,N_3714);
nor U6883 (N_6883,N_5885,N_5522);
or U6884 (N_6884,N_4050,N_3528);
nor U6885 (N_6885,N_4216,N_5860);
xnor U6886 (N_6886,N_5035,N_3303);
xor U6887 (N_6887,N_3565,N_4456);
nand U6888 (N_6888,N_3589,N_4683);
or U6889 (N_6889,N_5218,N_5626);
and U6890 (N_6890,N_5612,N_5206);
nand U6891 (N_6891,N_5343,N_4393);
or U6892 (N_6892,N_5698,N_4120);
and U6893 (N_6893,N_4278,N_4246);
nor U6894 (N_6894,N_4465,N_3088);
xnor U6895 (N_6895,N_3172,N_3093);
and U6896 (N_6896,N_3233,N_4854);
or U6897 (N_6897,N_3716,N_3054);
nor U6898 (N_6898,N_3991,N_4355);
nor U6899 (N_6899,N_5367,N_4666);
nand U6900 (N_6900,N_5893,N_5057);
nor U6901 (N_6901,N_4085,N_4890);
and U6902 (N_6902,N_5462,N_4036);
or U6903 (N_6903,N_5614,N_5427);
nor U6904 (N_6904,N_3734,N_3943);
xnor U6905 (N_6905,N_5105,N_4086);
nand U6906 (N_6906,N_4414,N_3095);
and U6907 (N_6907,N_5445,N_4817);
and U6908 (N_6908,N_4388,N_5842);
nor U6909 (N_6909,N_3448,N_5714);
or U6910 (N_6910,N_4624,N_3591);
and U6911 (N_6911,N_5700,N_3983);
and U6912 (N_6912,N_5867,N_5743);
and U6913 (N_6913,N_5146,N_4849);
and U6914 (N_6914,N_3700,N_3949);
and U6915 (N_6915,N_3290,N_4175);
nor U6916 (N_6916,N_5076,N_5965);
or U6917 (N_6917,N_3932,N_5238);
nor U6918 (N_6918,N_3975,N_4259);
nor U6919 (N_6919,N_5707,N_5176);
xor U6920 (N_6920,N_3503,N_5837);
and U6921 (N_6921,N_4221,N_5870);
xnor U6922 (N_6922,N_4073,N_3101);
xor U6923 (N_6923,N_4060,N_3041);
xnor U6924 (N_6924,N_4823,N_5010);
xnor U6925 (N_6925,N_4824,N_3675);
and U6926 (N_6926,N_5434,N_5724);
or U6927 (N_6927,N_5640,N_3597);
or U6928 (N_6928,N_4430,N_4606);
and U6929 (N_6929,N_4280,N_3069);
nor U6930 (N_6930,N_3767,N_4705);
and U6931 (N_6931,N_5526,N_4334);
or U6932 (N_6932,N_5986,N_4671);
nor U6933 (N_6933,N_5496,N_3891);
nand U6934 (N_6934,N_4167,N_4894);
xor U6935 (N_6935,N_5539,N_4655);
nor U6936 (N_6936,N_3216,N_3266);
or U6937 (N_6937,N_4878,N_4713);
nor U6938 (N_6938,N_5013,N_5486);
and U6939 (N_6939,N_4928,N_3252);
nor U6940 (N_6940,N_4920,N_5599);
nand U6941 (N_6941,N_3958,N_3307);
nor U6942 (N_6942,N_3455,N_3359);
nor U6943 (N_6943,N_3072,N_4047);
and U6944 (N_6944,N_4404,N_3016);
and U6945 (N_6945,N_5545,N_3956);
or U6946 (N_6946,N_3263,N_4429);
nand U6947 (N_6947,N_5363,N_4798);
or U6948 (N_6948,N_4879,N_5722);
xnor U6949 (N_6949,N_3012,N_4673);
xnor U6950 (N_6950,N_4295,N_5090);
nor U6951 (N_6951,N_3249,N_3861);
nor U6952 (N_6952,N_3988,N_5945);
nor U6953 (N_6953,N_3137,N_3486);
and U6954 (N_6954,N_3551,N_3653);
nand U6955 (N_6955,N_5949,N_3613);
and U6956 (N_6956,N_3129,N_4257);
xor U6957 (N_6957,N_4154,N_3980);
or U6958 (N_6958,N_5244,N_3168);
nand U6959 (N_6959,N_4886,N_5422);
and U6960 (N_6960,N_5648,N_5985);
nor U6961 (N_6961,N_4588,N_3836);
nand U6962 (N_6962,N_3299,N_4241);
nor U6963 (N_6963,N_3264,N_3996);
nor U6964 (N_6964,N_3856,N_4739);
nor U6965 (N_6965,N_4564,N_5349);
xor U6966 (N_6966,N_3265,N_3801);
nor U6967 (N_6967,N_5922,N_4517);
or U6968 (N_6968,N_3828,N_4605);
or U6969 (N_6969,N_4223,N_3148);
or U6970 (N_6970,N_3623,N_4746);
nor U6971 (N_6971,N_3773,N_5598);
nor U6972 (N_6972,N_3924,N_5600);
or U6973 (N_6973,N_5186,N_5435);
xor U6974 (N_6974,N_4135,N_3560);
or U6975 (N_6975,N_3576,N_4493);
or U6976 (N_6976,N_5656,N_4795);
and U6977 (N_6977,N_3720,N_3135);
nand U6978 (N_6978,N_5262,N_3538);
xor U6979 (N_6979,N_5481,N_3200);
or U6980 (N_6980,N_4130,N_4463);
and U6981 (N_6981,N_3371,N_4607);
and U6982 (N_6982,N_4910,N_5404);
xnor U6983 (N_6983,N_4266,N_5512);
and U6984 (N_6984,N_5417,N_5171);
nor U6985 (N_6985,N_4701,N_3356);
nor U6986 (N_6986,N_4693,N_5825);
nor U6987 (N_6987,N_4730,N_3662);
nor U6988 (N_6988,N_5988,N_4239);
nand U6989 (N_6989,N_3409,N_5951);
or U6990 (N_6990,N_4263,N_4529);
xnor U6991 (N_6991,N_4052,N_4715);
or U6992 (N_6992,N_5532,N_4009);
xor U6993 (N_6993,N_5328,N_5426);
nand U6994 (N_6994,N_4273,N_5788);
nor U6995 (N_6995,N_3886,N_3340);
and U6996 (N_6996,N_3847,N_3262);
nand U6997 (N_6997,N_4632,N_4005);
nand U6998 (N_6998,N_3851,N_3084);
or U6999 (N_6999,N_3412,N_5915);
nand U7000 (N_7000,N_4094,N_4108);
and U7001 (N_7001,N_4971,N_3850);
nand U7002 (N_7002,N_5465,N_4969);
nand U7003 (N_7003,N_5651,N_5313);
or U7004 (N_7004,N_4224,N_3149);
nand U7005 (N_7005,N_3945,N_5118);
and U7006 (N_7006,N_3950,N_3871);
xor U7007 (N_7007,N_5390,N_4276);
nand U7008 (N_7008,N_5438,N_5582);
or U7009 (N_7009,N_4895,N_3349);
or U7010 (N_7010,N_5947,N_3496);
or U7011 (N_7011,N_3477,N_5862);
xnor U7012 (N_7012,N_5104,N_5777);
nor U7013 (N_7013,N_4310,N_5994);
nor U7014 (N_7014,N_5726,N_4916);
and U7015 (N_7015,N_4020,N_3366);
xor U7016 (N_7016,N_5711,N_5898);
xnor U7017 (N_7017,N_3827,N_3676);
xnor U7018 (N_7018,N_5239,N_5335);
nor U7019 (N_7019,N_3971,N_4492);
nand U7020 (N_7020,N_3139,N_5733);
xor U7021 (N_7021,N_3492,N_4297);
and U7022 (N_7022,N_5792,N_5546);
nand U7023 (N_7023,N_3603,N_4699);
xnor U7024 (N_7024,N_5364,N_3004);
and U7025 (N_7025,N_3805,N_5038);
xnor U7026 (N_7026,N_5430,N_3238);
and U7027 (N_7027,N_5135,N_5521);
or U7028 (N_7028,N_4742,N_4288);
nor U7029 (N_7029,N_3684,N_4538);
xor U7030 (N_7030,N_5901,N_5211);
and U7031 (N_7031,N_5571,N_4650);
and U7032 (N_7032,N_5405,N_3378);
xnor U7033 (N_7033,N_4536,N_3823);
nor U7034 (N_7034,N_3335,N_4782);
nor U7035 (N_7035,N_5099,N_4518);
or U7036 (N_7036,N_4208,N_4369);
xor U7037 (N_7037,N_3131,N_4700);
nor U7038 (N_7038,N_3333,N_4774);
nor U7039 (N_7039,N_5844,N_5891);
nor U7040 (N_7040,N_3176,N_5478);
nor U7041 (N_7041,N_4514,N_3365);
xnor U7042 (N_7042,N_5671,N_3250);
nand U7043 (N_7043,N_5093,N_5643);
or U7044 (N_7044,N_4400,N_4227);
xnor U7045 (N_7045,N_3036,N_4967);
or U7046 (N_7046,N_4846,N_4618);
and U7047 (N_7047,N_3345,N_3406);
or U7048 (N_7048,N_5369,N_3332);
or U7049 (N_7049,N_3433,N_3175);
and U7050 (N_7050,N_5201,N_5584);
and U7051 (N_7051,N_5570,N_4284);
or U7052 (N_7052,N_4294,N_5840);
and U7053 (N_7053,N_5299,N_4875);
or U7054 (N_7054,N_4474,N_5541);
xor U7055 (N_7055,N_5967,N_4043);
or U7056 (N_7056,N_3323,N_4544);
or U7057 (N_7057,N_3514,N_3707);
nor U7058 (N_7058,N_3938,N_3398);
xor U7059 (N_7059,N_5715,N_3089);
and U7060 (N_7060,N_4485,N_5735);
and U7061 (N_7061,N_4869,N_4006);
nand U7062 (N_7062,N_3788,N_5235);
xnor U7063 (N_7063,N_5169,N_3106);
nand U7064 (N_7064,N_4228,N_4035);
nor U7065 (N_7065,N_5431,N_3483);
nand U7066 (N_7066,N_3879,N_3119);
or U7067 (N_7067,N_5998,N_5255);
or U7068 (N_7068,N_4592,N_4772);
nand U7069 (N_7069,N_5741,N_5876);
nor U7070 (N_7070,N_3476,N_4442);
nand U7071 (N_7071,N_5464,N_5696);
nand U7072 (N_7072,N_3367,N_3258);
nor U7073 (N_7073,N_5415,N_3736);
xor U7074 (N_7074,N_5044,N_5529);
nor U7075 (N_7075,N_5103,N_4372);
xor U7076 (N_7076,N_5523,N_3063);
xnor U7077 (N_7077,N_4045,N_3633);
nor U7078 (N_7078,N_5489,N_5028);
xor U7079 (N_7079,N_5672,N_3123);
and U7080 (N_7080,N_5444,N_3798);
nand U7081 (N_7081,N_4852,N_4423);
nor U7082 (N_7082,N_4434,N_5398);
nor U7083 (N_7083,N_4098,N_3543);
xnor U7084 (N_7084,N_5874,N_3162);
or U7085 (N_7085,N_4185,N_4556);
nor U7086 (N_7086,N_4141,N_5573);
xor U7087 (N_7087,N_4755,N_4851);
and U7088 (N_7088,N_3853,N_4645);
nor U7089 (N_7089,N_4757,N_5699);
nor U7090 (N_7090,N_5595,N_5254);
or U7091 (N_7091,N_4207,N_4914);
or U7092 (N_7092,N_5241,N_5790);
nor U7093 (N_7093,N_5261,N_5518);
nor U7094 (N_7094,N_3113,N_4147);
and U7095 (N_7095,N_4905,N_4552);
or U7096 (N_7096,N_5764,N_5150);
nor U7097 (N_7097,N_4397,N_3571);
and U7098 (N_7098,N_5064,N_5181);
and U7099 (N_7099,N_4178,N_3515);
xor U7100 (N_7100,N_4490,N_3489);
or U7101 (N_7101,N_5929,N_5841);
and U7102 (N_7102,N_5295,N_5332);
nor U7103 (N_7103,N_5633,N_5208);
and U7104 (N_7104,N_3668,N_4140);
nor U7105 (N_7105,N_5183,N_3388);
and U7106 (N_7106,N_4338,N_4249);
and U7107 (N_7107,N_3395,N_3308);
nand U7108 (N_7108,N_5372,N_5151);
nand U7109 (N_7109,N_3034,N_5297);
nor U7110 (N_7110,N_4546,N_3970);
and U7111 (N_7111,N_5511,N_3777);
nor U7112 (N_7112,N_4631,N_5403);
nand U7113 (N_7113,N_3320,N_4329);
xnor U7114 (N_7114,N_3698,N_3218);
and U7115 (N_7115,N_5749,N_3590);
and U7116 (N_7116,N_3300,N_4037);
xor U7117 (N_7117,N_3584,N_3889);
xor U7118 (N_7118,N_3875,N_4966);
xor U7119 (N_7119,N_4210,N_3821);
or U7120 (N_7120,N_5713,N_4682);
nor U7121 (N_7121,N_5856,N_4053);
or U7122 (N_7122,N_3420,N_3446);
xnor U7123 (N_7123,N_3830,N_5679);
and U7124 (N_7124,N_5779,N_4825);
and U7125 (N_7125,N_4860,N_4616);
and U7126 (N_7126,N_3494,N_3630);
or U7127 (N_7127,N_3053,N_5006);
or U7128 (N_7128,N_4303,N_4584);
and U7129 (N_7129,N_5543,N_4326);
nand U7130 (N_7130,N_4152,N_4361);
and U7131 (N_7131,N_4570,N_3151);
xnor U7132 (N_7132,N_4028,N_3521);
and U7133 (N_7133,N_3342,N_4104);
nor U7134 (N_7134,N_4116,N_4927);
and U7135 (N_7135,N_5302,N_5149);
xnor U7136 (N_7136,N_4475,N_3050);
or U7137 (N_7137,N_5627,N_4744);
xor U7138 (N_7138,N_5358,N_4516);
xor U7139 (N_7139,N_5400,N_5851);
xor U7140 (N_7140,N_5778,N_4558);
or U7141 (N_7141,N_4211,N_3288);
nand U7142 (N_7142,N_3322,N_4403);
and U7143 (N_7143,N_4929,N_4346);
nand U7144 (N_7144,N_5017,N_3926);
nand U7145 (N_7145,N_5968,N_3436);
xor U7146 (N_7146,N_5108,N_3826);
nand U7147 (N_7147,N_5470,N_4997);
and U7148 (N_7148,N_3831,N_4354);
nor U7149 (N_7149,N_5879,N_4870);
nand U7150 (N_7150,N_5848,N_3888);
xnor U7151 (N_7151,N_5721,N_5483);
or U7152 (N_7152,N_3940,N_3432);
xnor U7153 (N_7153,N_3347,N_5861);
and U7154 (N_7154,N_5197,N_3880);
xnor U7155 (N_7155,N_3647,N_5785);
or U7156 (N_7156,N_5662,N_4170);
and U7157 (N_7157,N_3715,N_5544);
xor U7158 (N_7158,N_3664,N_4542);
or U7159 (N_7159,N_3147,N_4398);
nand U7160 (N_7160,N_4547,N_3354);
nand U7161 (N_7161,N_3403,N_4843);
xnor U7162 (N_7162,N_3064,N_5921);
and U7163 (N_7163,N_4225,N_3317);
or U7164 (N_7164,N_5760,N_4943);
xor U7165 (N_7165,N_5981,N_3954);
nand U7166 (N_7166,N_3385,N_3820);
and U7167 (N_7167,N_3512,N_3318);
nand U7168 (N_7168,N_3426,N_3269);
or U7169 (N_7169,N_4461,N_4460);
nor U7170 (N_7170,N_3228,N_5871);
and U7171 (N_7171,N_5256,N_5625);
nand U7172 (N_7172,N_4935,N_5174);
or U7173 (N_7173,N_3193,N_5800);
nor U7174 (N_7174,N_3742,N_5305);
xor U7175 (N_7175,N_5952,N_4041);
nand U7176 (N_7176,N_5298,N_4306);
xnor U7177 (N_7177,N_5428,N_4575);
or U7178 (N_7178,N_4549,N_3781);
and U7179 (N_7179,N_5980,N_3869);
xnor U7180 (N_7180,N_4498,N_5153);
xor U7181 (N_7181,N_5314,N_4018);
xnor U7182 (N_7182,N_5144,N_5407);
and U7183 (N_7183,N_5832,N_4335);
xnor U7184 (N_7184,N_3516,N_4731);
and U7185 (N_7185,N_4250,N_5142);
nor U7186 (N_7186,N_5493,N_3051);
xor U7187 (N_7187,N_4439,N_3007);
xor U7188 (N_7188,N_5382,N_3132);
and U7189 (N_7189,N_3718,N_3058);
xor U7190 (N_7190,N_4427,N_5520);
nand U7191 (N_7191,N_3527,N_4136);
nand U7192 (N_7192,N_3210,N_3253);
nand U7193 (N_7193,N_3846,N_5728);
xnor U7194 (N_7194,N_4200,N_3485);
nand U7195 (N_7195,N_5984,N_5513);
nor U7196 (N_7196,N_3899,N_3165);
xor U7197 (N_7197,N_5666,N_5336);
or U7198 (N_7198,N_3722,N_3242);
or U7199 (N_7199,N_3599,N_5296);
nand U7200 (N_7200,N_4876,N_4453);
xor U7201 (N_7201,N_5972,N_3701);
or U7202 (N_7202,N_4714,N_3125);
xnor U7203 (N_7203,N_3711,N_5492);
xor U7204 (N_7204,N_5608,N_4597);
nand U7205 (N_7205,N_3470,N_3726);
nor U7206 (N_7206,N_3133,N_5928);
or U7207 (N_7207,N_4436,N_3102);
nand U7208 (N_7208,N_3925,N_4156);
nand U7209 (N_7209,N_4513,N_5993);
nor U7210 (N_7210,N_3011,N_4153);
nand U7211 (N_7211,N_3222,N_3078);
or U7212 (N_7212,N_5288,N_5797);
and U7213 (N_7213,N_3325,N_5920);
or U7214 (N_7214,N_3882,N_4385);
and U7215 (N_7215,N_5776,N_4016);
xnor U7216 (N_7216,N_3295,N_5134);
and U7217 (N_7217,N_5926,N_3417);
and U7218 (N_7218,N_4040,N_4074);
nand U7219 (N_7219,N_5607,N_5116);
and U7220 (N_7220,N_4357,N_4118);
xor U7221 (N_7221,N_4691,N_5577);
nor U7222 (N_7222,N_5882,N_4247);
xor U7223 (N_7223,N_5381,N_5635);
nor U7224 (N_7224,N_3573,N_3848);
nand U7225 (N_7225,N_4815,N_3825);
nor U7226 (N_7226,N_5110,N_4627);
or U7227 (N_7227,N_3298,N_5590);
nand U7228 (N_7228,N_3681,N_4664);
nor U7229 (N_7229,N_4885,N_4245);
nor U7230 (N_7230,N_3666,N_4785);
nand U7231 (N_7231,N_5549,N_4123);
or U7232 (N_7232,N_3966,N_3042);
and U7233 (N_7233,N_5114,N_4070);
or U7234 (N_7234,N_3942,N_3577);
and U7235 (N_7235,N_5468,N_3957);
xnor U7236 (N_7236,N_3608,N_3296);
xor U7237 (N_7237,N_5652,N_3360);
nor U7238 (N_7238,N_5849,N_4637);
xnor U7239 (N_7239,N_5834,N_4692);
nand U7240 (N_7240,N_4196,N_5315);
or U7241 (N_7241,N_4444,N_3655);
or U7242 (N_7242,N_4287,N_3824);
nor U7243 (N_7243,N_3678,N_4850);
and U7244 (N_7244,N_4898,N_5162);
and U7245 (N_7245,N_3244,N_4533);
or U7246 (N_7246,N_4144,N_5308);
and U7247 (N_7247,N_4134,N_5221);
and U7248 (N_7248,N_3085,N_4781);
and U7249 (N_7249,N_4924,N_4904);
xor U7250 (N_7250,N_3114,N_3728);
nand U7251 (N_7251,N_5413,N_4719);
or U7252 (N_7252,N_3990,N_5227);
nor U7253 (N_7253,N_3786,N_3109);
nor U7254 (N_7254,N_5857,N_5694);
nand U7255 (N_7255,N_3404,N_5631);
xor U7256 (N_7256,N_3979,N_5729);
xnor U7257 (N_7257,N_3796,N_4608);
and U7258 (N_7258,N_3896,N_4451);
nor U7259 (N_7259,N_4770,N_5284);
nand U7260 (N_7260,N_3048,N_4333);
and U7261 (N_7261,N_3818,N_5514);
xnor U7262 (N_7262,N_4557,N_5934);
nor U7263 (N_7263,N_4960,N_4736);
xnor U7264 (N_7264,N_4738,N_4950);
xnor U7265 (N_7265,N_5794,N_3761);
xnor U7266 (N_7266,N_4115,N_4806);
and U7267 (N_7267,N_4051,N_3592);
and U7268 (N_7268,N_3556,N_3279);
or U7269 (N_7269,N_5506,N_3226);
and U7270 (N_7270,N_3785,N_5588);
nand U7271 (N_7271,N_5380,N_5997);
xnor U7272 (N_7272,N_4265,N_3772);
or U7273 (N_7273,N_4371,N_5419);
nor U7274 (N_7274,N_5910,N_3057);
xor U7275 (N_7275,N_3870,N_5259);
and U7276 (N_7276,N_4978,N_4180);
or U7277 (N_7277,N_4725,N_4386);
xnor U7278 (N_7278,N_3062,N_4915);
xnor U7279 (N_7279,N_5145,N_5019);
or U7280 (N_7280,N_4764,N_4301);
and U7281 (N_7281,N_3260,N_4395);
nor U7282 (N_7282,N_4534,N_3389);
nand U7283 (N_7283,N_3467,N_4889);
xor U7284 (N_7284,N_4191,N_5883);
xnor U7285 (N_7285,N_5605,N_4807);
or U7286 (N_7286,N_3883,N_3721);
or U7287 (N_7287,N_4151,N_4814);
nand U7288 (N_7288,N_4057,N_5409);
and U7289 (N_7289,N_4816,N_3456);
xor U7290 (N_7290,N_4758,N_5232);
or U7291 (N_7291,N_5387,N_5989);
or U7292 (N_7292,N_3570,N_3549);
and U7293 (N_7293,N_3010,N_5773);
nor U7294 (N_7294,N_4099,N_4636);
xnor U7295 (N_7295,N_4479,N_4187);
nor U7296 (N_7296,N_5507,N_3195);
or U7297 (N_7297,N_4932,N_5826);
nor U7298 (N_7298,N_5807,N_4483);
nand U7299 (N_7299,N_3506,N_3993);
and U7300 (N_7300,N_3555,N_5739);
nand U7301 (N_7301,N_4100,N_5198);
and U7302 (N_7302,N_4275,N_3474);
or U7303 (N_7303,N_3127,N_4367);
or U7304 (N_7304,N_5402,N_4075);
or U7305 (N_7305,N_4647,N_3819);
or U7306 (N_7306,N_5089,N_5845);
nand U7307 (N_7307,N_5517,N_3510);
nor U7308 (N_7308,N_4771,N_4845);
nand U7309 (N_7309,N_3897,N_3579);
nand U7310 (N_7310,N_4555,N_5027);
xor U7311 (N_7311,N_3909,N_5973);
nor U7312 (N_7312,N_5383,N_4989);
nand U7313 (N_7313,N_5406,N_4106);
nand U7314 (N_7314,N_5931,N_3855);
or U7315 (N_7315,N_5002,N_4827);
or U7316 (N_7316,N_3920,N_5214);
xor U7317 (N_7317,N_3535,N_4821);
and U7318 (N_7318,N_3706,N_4477);
or U7319 (N_7319,N_4424,N_5559);
xor U7320 (N_7320,N_3257,N_5416);
nor U7321 (N_7321,N_5448,N_5317);
and U7322 (N_7322,N_5050,N_3118);
nand U7323 (N_7323,N_5274,N_3441);
or U7324 (N_7324,N_4613,N_3628);
nor U7325 (N_7325,N_5905,N_5499);
nor U7326 (N_7326,N_4865,N_4410);
or U7327 (N_7327,N_3892,N_3336);
nand U7328 (N_7328,N_4061,N_3790);
and U7329 (N_7329,N_4248,N_3541);
nand U7330 (N_7330,N_3484,N_3572);
or U7331 (N_7331,N_4523,N_4903);
or U7332 (N_7332,N_4458,N_5958);
and U7333 (N_7333,N_5085,N_5371);
and U7334 (N_7334,N_4426,N_3581);
and U7335 (N_7335,N_3156,N_3473);
or U7336 (N_7336,N_3487,N_5450);
or U7337 (N_7337,N_5021,N_3858);
nor U7338 (N_7338,N_3381,N_3842);
nor U7339 (N_7339,N_4899,N_5164);
nand U7340 (N_7340,N_5280,N_3974);
xor U7341 (N_7341,N_5923,N_3196);
xor U7342 (N_7342,N_5731,N_4234);
xnor U7343 (N_7343,N_5944,N_3863);
and U7344 (N_7344,N_4961,N_3272);
or U7345 (N_7345,N_4201,N_3694);
xnor U7346 (N_7346,N_5215,N_4838);
and U7347 (N_7347,N_4342,N_3037);
nor U7348 (N_7348,N_4799,N_4146);
xor U7349 (N_7349,N_5242,N_5053);
xor U7350 (N_7350,N_5226,N_3729);
or U7351 (N_7351,N_5575,N_4325);
or U7352 (N_7352,N_3611,N_4768);
and U7353 (N_7353,N_5689,N_4792);
xor U7354 (N_7354,N_3624,N_4351);
nand U7355 (N_7355,N_3099,N_5101);
and U7356 (N_7356,N_3845,N_5182);
nand U7357 (N_7357,N_3984,N_4062);
or U7358 (N_7358,N_3750,N_4103);
and U7359 (N_7359,N_5854,N_4503);
and U7360 (N_7360,N_3457,N_3933);
nor U7361 (N_7361,N_5663,N_4177);
nor U7362 (N_7362,N_5601,N_4602);
and U7363 (N_7363,N_5868,N_3310);
nand U7364 (N_7364,N_5077,N_4754);
nand U7365 (N_7365,N_3936,N_5748);
and U7366 (N_7366,N_4907,N_3044);
xor U7367 (N_7367,N_4612,N_5195);
or U7368 (N_7368,N_5847,N_3697);
and U7369 (N_7369,N_4488,N_5859);
or U7370 (N_7370,N_5113,N_5043);
nand U7371 (N_7371,N_4548,N_5510);
nand U7372 (N_7372,N_5060,N_4840);
or U7373 (N_7373,N_3548,N_4125);
nand U7374 (N_7374,N_4527,N_4797);
xnor U7375 (N_7375,N_5189,N_5304);
or U7376 (N_7376,N_4069,N_5758);
and U7377 (N_7377,N_3103,N_5126);
or U7378 (N_7378,N_3547,N_3491);
or U7379 (N_7379,N_5376,N_3120);
nand U7380 (N_7380,N_5617,N_3612);
nand U7381 (N_7381,N_3760,N_3462);
xnor U7382 (N_7382,N_3239,N_5802);
nor U7383 (N_7383,N_3461,N_4628);
nor U7384 (N_7384,N_4526,N_4360);
nor U7385 (N_7385,N_3600,N_5348);
or U7386 (N_7386,N_3463,N_3220);
xnor U7387 (N_7387,N_3302,N_4524);
and U7388 (N_7388,N_3013,N_3192);
or U7389 (N_7389,N_4142,N_5329);
or U7390 (N_7390,N_5830,N_3277);
and U7391 (N_7391,N_5271,N_4299);
or U7392 (N_7392,N_4166,N_4619);
nor U7393 (N_7393,N_4561,N_5747);
nand U7394 (N_7394,N_5533,N_3844);
xnor U7395 (N_7395,N_4563,N_5971);
and U7396 (N_7396,N_4712,N_4447);
or U7397 (N_7397,N_4609,N_3650);
and U7398 (N_7398,N_4834,N_3689);
and U7399 (N_7399,N_4183,N_5621);
nor U7400 (N_7400,N_3906,N_5455);
xnor U7401 (N_7401,N_5018,N_3765);
nor U7402 (N_7402,N_5449,N_4055);
and U7403 (N_7403,N_3271,N_4495);
or U7404 (N_7404,N_3854,N_5148);
xnor U7405 (N_7405,N_5622,N_3982);
nand U7406 (N_7406,N_3910,N_3052);
or U7407 (N_7407,N_5161,N_5939);
and U7408 (N_7408,N_4358,N_3223);
and U7409 (N_7409,N_4881,N_4600);
nand U7410 (N_7410,N_5374,N_4720);
and U7411 (N_7411,N_5563,N_3458);
nor U7412 (N_7412,N_3275,N_5941);
and U7413 (N_7413,N_5576,N_3637);
xnor U7414 (N_7414,N_4695,N_5283);
nor U7415 (N_7415,N_3864,N_3392);
and U7416 (N_7416,N_4394,N_5831);
or U7417 (N_7417,N_3297,N_3923);
or U7418 (N_7418,N_5333,N_3032);
nor U7419 (N_7419,N_3969,N_3873);
nor U7420 (N_7420,N_3568,N_5670);
nand U7421 (N_7421,N_5123,N_4220);
nand U7422 (N_7422,N_5712,N_3799);
or U7423 (N_7423,N_4676,N_5613);
xor U7424 (N_7424,N_4391,N_3610);
or U7425 (N_7425,N_3443,N_3658);
xnor U7426 (N_7426,N_4751,N_3115);
nand U7427 (N_7427,N_4149,N_3493);
nand U7428 (N_7428,N_5555,N_4340);
or U7429 (N_7429,N_4215,N_5373);
or U7430 (N_7430,N_5451,N_5638);
nor U7431 (N_7431,N_4642,N_3130);
and U7432 (N_7432,N_3430,N_5203);
nand U7433 (N_7433,N_5365,N_4844);
xor U7434 (N_7434,N_4502,N_4941);
nor U7435 (N_7435,N_5916,N_5258);
nand U7436 (N_7436,N_3616,N_3190);
nand U7437 (N_7437,N_5307,N_3948);
or U7438 (N_7438,N_4312,N_4454);
nand U7439 (N_7439,N_5325,N_4049);
and U7440 (N_7440,N_3188,N_3107);
xor U7441 (N_7441,N_3111,N_5657);
xnor U7442 (N_7442,N_5553,N_5687);
or U7443 (N_7443,N_3097,N_3039);
and U7444 (N_7444,N_5312,N_5527);
xnor U7445 (N_7445,N_4443,N_4986);
nor U7446 (N_7446,N_5433,N_4316);
and U7447 (N_7447,N_4264,N_5821);
nor U7448 (N_7448,N_4019,N_5477);
nand U7449 (N_7449,N_4543,N_3002);
xnor U7450 (N_7450,N_4370,N_4413);
and U7451 (N_7451,N_3055,N_4839);
and U7452 (N_7452,N_3626,N_4992);
xnor U7453 (N_7453,N_4945,N_5693);
and U7454 (N_7454,N_5388,N_5379);
xor U7455 (N_7455,N_5710,N_4101);
nand U7456 (N_7456,N_5205,N_3289);
and U7457 (N_7457,N_3001,N_4985);
nand U7458 (N_7458,N_4330,N_3832);
nand U7459 (N_7459,N_4260,N_3017);
nand U7460 (N_7460,N_5469,N_4270);
and U7461 (N_7461,N_3976,N_3912);
nand U7462 (N_7462,N_4244,N_4571);
and U7463 (N_7463,N_3025,N_3475);
xor U7464 (N_7464,N_4964,N_4801);
nor U7465 (N_7465,N_4362,N_5353);
or U7466 (N_7466,N_4431,N_5900);
nor U7467 (N_7467,N_5630,N_3363);
or U7468 (N_7468,N_3968,N_3709);
and U7469 (N_7469,N_4381,N_3753);
and U7470 (N_7470,N_4145,N_4617);
nor U7471 (N_7471,N_3479,N_3724);
and U7472 (N_7472,N_5585,N_4129);
or U7473 (N_7473,N_4077,N_4364);
and U7474 (N_7474,N_3774,N_4741);
xor U7475 (N_7475,N_3083,N_5408);
nor U7476 (N_7476,N_4368,N_3030);
or U7477 (N_7477,N_3182,N_5245);
and U7478 (N_7478,N_5082,N_3169);
and U7479 (N_7479,N_4078,N_5233);
nor U7480 (N_7480,N_4131,N_3683);
or U7481 (N_7481,N_3884,N_3358);
xor U7482 (N_7482,N_4188,N_5839);
nor U7483 (N_7483,N_4512,N_4464);
nor U7484 (N_7484,N_5669,N_3478);
nand U7485 (N_7485,N_3517,N_3498);
or U7486 (N_7486,N_4982,N_3414);
xor U7487 (N_7487,N_3691,N_4097);
nand U7488 (N_7488,N_5491,N_3977);
or U7489 (N_7489,N_5504,N_4459);
or U7490 (N_7490,N_5322,N_3800);
xnor U7491 (N_7491,N_4232,N_4948);
or U7492 (N_7492,N_4716,N_4481);
nand U7493 (N_7493,N_5378,N_3526);
or U7494 (N_7494,N_3415,N_3904);
and U7495 (N_7495,N_3046,N_3833);
xor U7496 (N_7496,N_3213,N_4735);
nand U7497 (N_7497,N_4332,N_5676);
xnor U7498 (N_7498,N_4026,N_5291);
nor U7499 (N_7499,N_4740,N_4867);
or U7500 (N_7500,N_3027,N_5689);
nor U7501 (N_7501,N_3725,N_5414);
nand U7502 (N_7502,N_5695,N_5872);
and U7503 (N_7503,N_3671,N_4718);
nand U7504 (N_7504,N_5444,N_5151);
nor U7505 (N_7505,N_3827,N_3156);
or U7506 (N_7506,N_3456,N_5139);
or U7507 (N_7507,N_5127,N_5261);
nand U7508 (N_7508,N_3507,N_5629);
or U7509 (N_7509,N_4897,N_3769);
and U7510 (N_7510,N_4935,N_4209);
or U7511 (N_7511,N_4507,N_4573);
and U7512 (N_7512,N_4763,N_5105);
or U7513 (N_7513,N_4071,N_3868);
nand U7514 (N_7514,N_5787,N_4074);
xor U7515 (N_7515,N_3997,N_5664);
and U7516 (N_7516,N_3286,N_4446);
nand U7517 (N_7517,N_5510,N_4956);
nand U7518 (N_7518,N_3701,N_4322);
or U7519 (N_7519,N_3741,N_3489);
xor U7520 (N_7520,N_4829,N_4497);
or U7521 (N_7521,N_3690,N_5582);
nand U7522 (N_7522,N_5454,N_4115);
nor U7523 (N_7523,N_3905,N_4425);
and U7524 (N_7524,N_4204,N_5752);
and U7525 (N_7525,N_4811,N_5326);
xor U7526 (N_7526,N_3082,N_5366);
nor U7527 (N_7527,N_4605,N_4197);
or U7528 (N_7528,N_3392,N_4881);
and U7529 (N_7529,N_5862,N_5443);
xor U7530 (N_7530,N_4664,N_4118);
xnor U7531 (N_7531,N_3009,N_5209);
or U7532 (N_7532,N_5265,N_5491);
and U7533 (N_7533,N_5249,N_4576);
or U7534 (N_7534,N_3982,N_3282);
or U7535 (N_7535,N_5570,N_4168);
nor U7536 (N_7536,N_5767,N_5490);
and U7537 (N_7537,N_4592,N_5707);
and U7538 (N_7538,N_3913,N_4222);
xnor U7539 (N_7539,N_4731,N_3548);
nor U7540 (N_7540,N_3677,N_5268);
nand U7541 (N_7541,N_3779,N_5128);
or U7542 (N_7542,N_5142,N_4598);
nand U7543 (N_7543,N_3663,N_3660);
and U7544 (N_7544,N_5860,N_3359);
xor U7545 (N_7545,N_4081,N_3787);
nor U7546 (N_7546,N_5802,N_4561);
nand U7547 (N_7547,N_3453,N_4677);
and U7548 (N_7548,N_5207,N_5555);
nand U7549 (N_7549,N_5087,N_4498);
nand U7550 (N_7550,N_5945,N_3047);
or U7551 (N_7551,N_3980,N_3795);
nand U7552 (N_7552,N_4036,N_3305);
xor U7553 (N_7553,N_3287,N_4478);
nand U7554 (N_7554,N_4759,N_4298);
nand U7555 (N_7555,N_3177,N_5133);
and U7556 (N_7556,N_3360,N_4056);
nor U7557 (N_7557,N_5912,N_4248);
or U7558 (N_7558,N_4260,N_4325);
xor U7559 (N_7559,N_5033,N_5328);
nand U7560 (N_7560,N_4499,N_5659);
and U7561 (N_7561,N_3471,N_3944);
nand U7562 (N_7562,N_5872,N_3327);
xor U7563 (N_7563,N_5236,N_3358);
and U7564 (N_7564,N_5135,N_5903);
xor U7565 (N_7565,N_3432,N_4726);
nand U7566 (N_7566,N_5715,N_4633);
nand U7567 (N_7567,N_3599,N_3469);
nand U7568 (N_7568,N_4219,N_5277);
xor U7569 (N_7569,N_4220,N_5446);
and U7570 (N_7570,N_3295,N_5698);
and U7571 (N_7571,N_5982,N_5649);
or U7572 (N_7572,N_5152,N_4924);
xor U7573 (N_7573,N_5682,N_5922);
and U7574 (N_7574,N_3450,N_4097);
nand U7575 (N_7575,N_3868,N_3102);
or U7576 (N_7576,N_5844,N_4399);
nand U7577 (N_7577,N_4229,N_4964);
or U7578 (N_7578,N_5054,N_3398);
nand U7579 (N_7579,N_5732,N_4638);
and U7580 (N_7580,N_4128,N_5727);
or U7581 (N_7581,N_4901,N_3271);
or U7582 (N_7582,N_5811,N_3290);
nor U7583 (N_7583,N_3845,N_4616);
or U7584 (N_7584,N_4407,N_4102);
nand U7585 (N_7585,N_5926,N_5631);
and U7586 (N_7586,N_5312,N_3236);
nand U7587 (N_7587,N_5569,N_3230);
or U7588 (N_7588,N_4770,N_4210);
nand U7589 (N_7589,N_4322,N_3531);
xor U7590 (N_7590,N_5064,N_5451);
xnor U7591 (N_7591,N_3060,N_4153);
nor U7592 (N_7592,N_3020,N_3662);
or U7593 (N_7593,N_5958,N_5125);
and U7594 (N_7594,N_4754,N_5107);
or U7595 (N_7595,N_5230,N_3077);
nor U7596 (N_7596,N_5631,N_4334);
xnor U7597 (N_7597,N_3306,N_5518);
or U7598 (N_7598,N_5992,N_4125);
nand U7599 (N_7599,N_4543,N_4420);
or U7600 (N_7600,N_5497,N_3136);
or U7601 (N_7601,N_5134,N_4425);
and U7602 (N_7602,N_3525,N_3582);
nor U7603 (N_7603,N_4132,N_3445);
and U7604 (N_7604,N_5693,N_4631);
or U7605 (N_7605,N_5607,N_5128);
or U7606 (N_7606,N_5878,N_3524);
xor U7607 (N_7607,N_4502,N_4191);
and U7608 (N_7608,N_4279,N_3302);
and U7609 (N_7609,N_5045,N_5499);
nand U7610 (N_7610,N_3249,N_5923);
xnor U7611 (N_7611,N_4338,N_3861);
xor U7612 (N_7612,N_5067,N_5345);
or U7613 (N_7613,N_4066,N_3312);
xnor U7614 (N_7614,N_3559,N_5034);
xnor U7615 (N_7615,N_5856,N_5220);
nor U7616 (N_7616,N_3653,N_3113);
xnor U7617 (N_7617,N_4425,N_4284);
nand U7618 (N_7618,N_5383,N_4431);
or U7619 (N_7619,N_5717,N_5853);
xnor U7620 (N_7620,N_3805,N_4628);
or U7621 (N_7621,N_5170,N_3802);
or U7622 (N_7622,N_5391,N_3031);
nor U7623 (N_7623,N_3638,N_4787);
nor U7624 (N_7624,N_5471,N_3319);
and U7625 (N_7625,N_4238,N_3099);
and U7626 (N_7626,N_3033,N_3150);
nor U7627 (N_7627,N_3148,N_4002);
or U7628 (N_7628,N_5074,N_3909);
and U7629 (N_7629,N_5277,N_3301);
nor U7630 (N_7630,N_4458,N_4568);
nor U7631 (N_7631,N_3717,N_3884);
xor U7632 (N_7632,N_3744,N_4018);
nand U7633 (N_7633,N_4981,N_4987);
nand U7634 (N_7634,N_3468,N_5315);
nor U7635 (N_7635,N_5189,N_5571);
or U7636 (N_7636,N_3627,N_3351);
and U7637 (N_7637,N_3701,N_4496);
xnor U7638 (N_7638,N_5492,N_5156);
xor U7639 (N_7639,N_3912,N_5586);
or U7640 (N_7640,N_3691,N_3730);
nor U7641 (N_7641,N_3717,N_4769);
and U7642 (N_7642,N_4796,N_3591);
and U7643 (N_7643,N_5208,N_4398);
nand U7644 (N_7644,N_3831,N_4436);
xor U7645 (N_7645,N_3354,N_4106);
xor U7646 (N_7646,N_5201,N_3443);
and U7647 (N_7647,N_3248,N_5169);
xnor U7648 (N_7648,N_4041,N_5423);
and U7649 (N_7649,N_5373,N_3029);
nand U7650 (N_7650,N_5664,N_4364);
nor U7651 (N_7651,N_3626,N_4136);
or U7652 (N_7652,N_5375,N_4159);
or U7653 (N_7653,N_5646,N_3046);
and U7654 (N_7654,N_4436,N_3369);
or U7655 (N_7655,N_4210,N_4735);
nor U7656 (N_7656,N_5756,N_3918);
xnor U7657 (N_7657,N_4458,N_4662);
xor U7658 (N_7658,N_5781,N_5101);
nand U7659 (N_7659,N_3807,N_4464);
nor U7660 (N_7660,N_5384,N_5169);
nand U7661 (N_7661,N_4721,N_4306);
and U7662 (N_7662,N_3772,N_4077);
nor U7663 (N_7663,N_3915,N_4672);
nor U7664 (N_7664,N_3971,N_3995);
xor U7665 (N_7665,N_3617,N_3038);
or U7666 (N_7666,N_3860,N_3738);
nor U7667 (N_7667,N_4428,N_5380);
or U7668 (N_7668,N_4768,N_4105);
nand U7669 (N_7669,N_4349,N_3197);
xor U7670 (N_7670,N_3966,N_3752);
nand U7671 (N_7671,N_4216,N_4639);
xnor U7672 (N_7672,N_5851,N_4087);
and U7673 (N_7673,N_3787,N_4463);
xnor U7674 (N_7674,N_3298,N_3197);
or U7675 (N_7675,N_4453,N_3890);
or U7676 (N_7676,N_5270,N_3640);
xnor U7677 (N_7677,N_5505,N_4264);
or U7678 (N_7678,N_4581,N_3741);
xnor U7679 (N_7679,N_5313,N_4964);
xnor U7680 (N_7680,N_3096,N_4686);
or U7681 (N_7681,N_4241,N_4534);
nor U7682 (N_7682,N_5176,N_4939);
or U7683 (N_7683,N_3554,N_5290);
nand U7684 (N_7684,N_3730,N_5920);
and U7685 (N_7685,N_3403,N_5745);
or U7686 (N_7686,N_5548,N_4700);
xnor U7687 (N_7687,N_5993,N_3682);
nand U7688 (N_7688,N_5826,N_4534);
nor U7689 (N_7689,N_5805,N_4797);
nor U7690 (N_7690,N_5098,N_4138);
and U7691 (N_7691,N_5003,N_5279);
nor U7692 (N_7692,N_4504,N_5625);
nor U7693 (N_7693,N_3183,N_5181);
xor U7694 (N_7694,N_3317,N_5064);
and U7695 (N_7695,N_3303,N_3633);
nand U7696 (N_7696,N_5348,N_4173);
and U7697 (N_7697,N_4952,N_5878);
nor U7698 (N_7698,N_3251,N_4122);
or U7699 (N_7699,N_3513,N_5723);
nand U7700 (N_7700,N_5800,N_4929);
and U7701 (N_7701,N_3857,N_5065);
nand U7702 (N_7702,N_4412,N_3910);
xnor U7703 (N_7703,N_5825,N_5565);
xor U7704 (N_7704,N_5628,N_4755);
nor U7705 (N_7705,N_3523,N_4022);
and U7706 (N_7706,N_3586,N_5423);
nor U7707 (N_7707,N_4681,N_3315);
nand U7708 (N_7708,N_5483,N_3077);
and U7709 (N_7709,N_4673,N_5418);
nor U7710 (N_7710,N_5943,N_3991);
or U7711 (N_7711,N_3419,N_3917);
nor U7712 (N_7712,N_4282,N_3258);
and U7713 (N_7713,N_3716,N_4730);
nor U7714 (N_7714,N_3329,N_3499);
and U7715 (N_7715,N_3623,N_3870);
nor U7716 (N_7716,N_4330,N_3666);
xor U7717 (N_7717,N_5557,N_5443);
or U7718 (N_7718,N_5997,N_3656);
or U7719 (N_7719,N_5967,N_5392);
or U7720 (N_7720,N_4088,N_4348);
nor U7721 (N_7721,N_5286,N_3217);
xnor U7722 (N_7722,N_4695,N_3758);
or U7723 (N_7723,N_3314,N_5432);
and U7724 (N_7724,N_4250,N_3353);
nand U7725 (N_7725,N_4072,N_4760);
and U7726 (N_7726,N_3761,N_4969);
nor U7727 (N_7727,N_3663,N_5893);
and U7728 (N_7728,N_5252,N_3374);
and U7729 (N_7729,N_5935,N_3858);
nand U7730 (N_7730,N_3587,N_5505);
or U7731 (N_7731,N_3036,N_5706);
xor U7732 (N_7732,N_5347,N_4001);
and U7733 (N_7733,N_4691,N_3407);
nand U7734 (N_7734,N_4373,N_4695);
or U7735 (N_7735,N_4883,N_5064);
or U7736 (N_7736,N_5019,N_4835);
or U7737 (N_7737,N_4473,N_4513);
xnor U7738 (N_7738,N_4923,N_3231);
nand U7739 (N_7739,N_4696,N_5359);
nor U7740 (N_7740,N_5738,N_4897);
nand U7741 (N_7741,N_5194,N_5013);
xor U7742 (N_7742,N_5276,N_5393);
xor U7743 (N_7743,N_5876,N_4546);
or U7744 (N_7744,N_5408,N_3880);
nor U7745 (N_7745,N_5067,N_5960);
and U7746 (N_7746,N_3869,N_3309);
nand U7747 (N_7747,N_3446,N_4879);
and U7748 (N_7748,N_4857,N_3093);
nand U7749 (N_7749,N_3873,N_5506);
or U7750 (N_7750,N_4362,N_4156);
or U7751 (N_7751,N_5824,N_4774);
nor U7752 (N_7752,N_4332,N_3181);
or U7753 (N_7753,N_5446,N_3630);
nor U7754 (N_7754,N_4567,N_3200);
nor U7755 (N_7755,N_4351,N_4444);
nand U7756 (N_7756,N_3159,N_5456);
or U7757 (N_7757,N_3474,N_5676);
or U7758 (N_7758,N_4219,N_5652);
nor U7759 (N_7759,N_5675,N_3029);
nand U7760 (N_7760,N_5086,N_5984);
or U7761 (N_7761,N_3381,N_3155);
or U7762 (N_7762,N_3603,N_4408);
nand U7763 (N_7763,N_5253,N_5287);
or U7764 (N_7764,N_5523,N_4406);
nand U7765 (N_7765,N_3923,N_4149);
xor U7766 (N_7766,N_4924,N_5107);
or U7767 (N_7767,N_5424,N_4843);
or U7768 (N_7768,N_5023,N_3373);
and U7769 (N_7769,N_5962,N_5169);
and U7770 (N_7770,N_5435,N_3567);
or U7771 (N_7771,N_3549,N_4830);
nor U7772 (N_7772,N_5738,N_3170);
or U7773 (N_7773,N_5288,N_5951);
or U7774 (N_7774,N_5352,N_5765);
xnor U7775 (N_7775,N_3415,N_5852);
xnor U7776 (N_7776,N_3287,N_5183);
nand U7777 (N_7777,N_3569,N_3845);
xnor U7778 (N_7778,N_5708,N_4547);
xor U7779 (N_7779,N_4513,N_5095);
xnor U7780 (N_7780,N_4526,N_5456);
xnor U7781 (N_7781,N_3787,N_3013);
nor U7782 (N_7782,N_3187,N_5146);
nand U7783 (N_7783,N_3030,N_4597);
nand U7784 (N_7784,N_4417,N_4195);
nor U7785 (N_7785,N_5222,N_4527);
nand U7786 (N_7786,N_5129,N_3429);
and U7787 (N_7787,N_3819,N_4018);
nor U7788 (N_7788,N_3534,N_5916);
nand U7789 (N_7789,N_3207,N_5340);
nor U7790 (N_7790,N_3579,N_5277);
nand U7791 (N_7791,N_3878,N_3602);
nor U7792 (N_7792,N_5460,N_3159);
xor U7793 (N_7793,N_4239,N_3449);
xor U7794 (N_7794,N_4632,N_3269);
and U7795 (N_7795,N_3078,N_5314);
nor U7796 (N_7796,N_3768,N_4733);
and U7797 (N_7797,N_3584,N_3189);
nor U7798 (N_7798,N_5096,N_3822);
nand U7799 (N_7799,N_5942,N_5885);
nor U7800 (N_7800,N_3126,N_4293);
or U7801 (N_7801,N_5093,N_5976);
xor U7802 (N_7802,N_3842,N_4774);
or U7803 (N_7803,N_5465,N_3949);
and U7804 (N_7804,N_5953,N_5693);
nor U7805 (N_7805,N_5831,N_3398);
nand U7806 (N_7806,N_3911,N_3111);
nand U7807 (N_7807,N_3969,N_5925);
nor U7808 (N_7808,N_3674,N_4952);
nand U7809 (N_7809,N_3259,N_5930);
and U7810 (N_7810,N_5109,N_4885);
or U7811 (N_7811,N_4976,N_5235);
or U7812 (N_7812,N_4932,N_5130);
nor U7813 (N_7813,N_3962,N_3480);
or U7814 (N_7814,N_3098,N_4327);
or U7815 (N_7815,N_4158,N_4246);
or U7816 (N_7816,N_4979,N_3608);
nor U7817 (N_7817,N_5290,N_4793);
nand U7818 (N_7818,N_4568,N_5054);
nand U7819 (N_7819,N_4313,N_3031);
nor U7820 (N_7820,N_4185,N_5038);
or U7821 (N_7821,N_5729,N_5649);
nand U7822 (N_7822,N_5877,N_3469);
and U7823 (N_7823,N_3367,N_5039);
and U7824 (N_7824,N_3735,N_4758);
nand U7825 (N_7825,N_4267,N_5021);
or U7826 (N_7826,N_3973,N_4517);
or U7827 (N_7827,N_3251,N_5674);
and U7828 (N_7828,N_5539,N_5560);
nor U7829 (N_7829,N_5701,N_5779);
nand U7830 (N_7830,N_5105,N_3133);
xnor U7831 (N_7831,N_4060,N_3278);
and U7832 (N_7832,N_5105,N_3041);
nand U7833 (N_7833,N_4258,N_4734);
nor U7834 (N_7834,N_3589,N_5766);
or U7835 (N_7835,N_5152,N_3969);
xor U7836 (N_7836,N_5966,N_4240);
or U7837 (N_7837,N_5519,N_3903);
and U7838 (N_7838,N_3863,N_5430);
or U7839 (N_7839,N_3066,N_5625);
xnor U7840 (N_7840,N_4944,N_5550);
or U7841 (N_7841,N_3131,N_4154);
xor U7842 (N_7842,N_5691,N_5668);
nand U7843 (N_7843,N_3980,N_4526);
or U7844 (N_7844,N_4160,N_5773);
nand U7845 (N_7845,N_5123,N_4713);
xor U7846 (N_7846,N_4644,N_5619);
and U7847 (N_7847,N_3804,N_4971);
xor U7848 (N_7848,N_4299,N_5593);
nor U7849 (N_7849,N_3170,N_5994);
nor U7850 (N_7850,N_4276,N_4848);
nor U7851 (N_7851,N_5889,N_3896);
nor U7852 (N_7852,N_3025,N_3699);
nand U7853 (N_7853,N_5158,N_5935);
and U7854 (N_7854,N_5245,N_4158);
nor U7855 (N_7855,N_3982,N_4673);
or U7856 (N_7856,N_5453,N_3279);
nand U7857 (N_7857,N_5676,N_5279);
or U7858 (N_7858,N_3608,N_5901);
nand U7859 (N_7859,N_3857,N_3083);
or U7860 (N_7860,N_3160,N_3420);
or U7861 (N_7861,N_4126,N_3763);
nor U7862 (N_7862,N_5383,N_5040);
nor U7863 (N_7863,N_3413,N_4938);
xnor U7864 (N_7864,N_5417,N_3739);
nor U7865 (N_7865,N_5877,N_5111);
nand U7866 (N_7866,N_3548,N_5028);
and U7867 (N_7867,N_3021,N_4383);
and U7868 (N_7868,N_3286,N_3363);
xor U7869 (N_7869,N_5749,N_3234);
nand U7870 (N_7870,N_5882,N_3917);
or U7871 (N_7871,N_3415,N_5197);
nand U7872 (N_7872,N_4818,N_4013);
nor U7873 (N_7873,N_5162,N_4667);
xor U7874 (N_7874,N_3854,N_4830);
or U7875 (N_7875,N_3843,N_3236);
and U7876 (N_7876,N_4453,N_5258);
and U7877 (N_7877,N_4180,N_4315);
and U7878 (N_7878,N_4472,N_4119);
nand U7879 (N_7879,N_3435,N_3916);
or U7880 (N_7880,N_3480,N_4746);
or U7881 (N_7881,N_4196,N_4034);
nor U7882 (N_7882,N_5768,N_5301);
nand U7883 (N_7883,N_3846,N_4255);
and U7884 (N_7884,N_4539,N_3085);
and U7885 (N_7885,N_4775,N_5528);
or U7886 (N_7886,N_5948,N_4230);
or U7887 (N_7887,N_4060,N_5880);
and U7888 (N_7888,N_3778,N_5828);
xor U7889 (N_7889,N_5535,N_4787);
nand U7890 (N_7890,N_5195,N_4643);
xnor U7891 (N_7891,N_5806,N_4631);
nand U7892 (N_7892,N_4550,N_4940);
nand U7893 (N_7893,N_3551,N_3009);
nand U7894 (N_7894,N_4097,N_3443);
nand U7895 (N_7895,N_5000,N_5857);
or U7896 (N_7896,N_5091,N_5660);
nor U7897 (N_7897,N_3207,N_4148);
and U7898 (N_7898,N_4230,N_3257);
or U7899 (N_7899,N_3695,N_3985);
nor U7900 (N_7900,N_5370,N_4204);
and U7901 (N_7901,N_3945,N_4440);
or U7902 (N_7902,N_4569,N_3706);
nand U7903 (N_7903,N_5024,N_5448);
nand U7904 (N_7904,N_3048,N_4741);
nor U7905 (N_7905,N_3358,N_4688);
xnor U7906 (N_7906,N_5805,N_5627);
nand U7907 (N_7907,N_4609,N_4429);
and U7908 (N_7908,N_3707,N_3860);
and U7909 (N_7909,N_5443,N_3164);
nor U7910 (N_7910,N_3712,N_3823);
nor U7911 (N_7911,N_3876,N_3738);
xor U7912 (N_7912,N_5324,N_4242);
xor U7913 (N_7913,N_3875,N_4380);
or U7914 (N_7914,N_5701,N_5444);
and U7915 (N_7915,N_4532,N_5126);
nor U7916 (N_7916,N_4330,N_4957);
and U7917 (N_7917,N_3367,N_4978);
xor U7918 (N_7918,N_3774,N_4484);
and U7919 (N_7919,N_3047,N_5644);
nand U7920 (N_7920,N_5232,N_4209);
nor U7921 (N_7921,N_3820,N_5426);
or U7922 (N_7922,N_3661,N_4695);
or U7923 (N_7923,N_5801,N_4426);
or U7924 (N_7924,N_4091,N_5407);
nand U7925 (N_7925,N_4226,N_4252);
and U7926 (N_7926,N_4902,N_3176);
xor U7927 (N_7927,N_5735,N_5083);
and U7928 (N_7928,N_5827,N_3723);
nor U7929 (N_7929,N_4015,N_5878);
nand U7930 (N_7930,N_5878,N_3060);
nand U7931 (N_7931,N_3190,N_5956);
and U7932 (N_7932,N_3624,N_5319);
or U7933 (N_7933,N_3245,N_5210);
or U7934 (N_7934,N_3415,N_5787);
xnor U7935 (N_7935,N_3075,N_4153);
and U7936 (N_7936,N_5618,N_5422);
xnor U7937 (N_7937,N_3856,N_3166);
xnor U7938 (N_7938,N_3006,N_5505);
xnor U7939 (N_7939,N_3238,N_4200);
nand U7940 (N_7940,N_5739,N_4499);
or U7941 (N_7941,N_5327,N_3339);
and U7942 (N_7942,N_3144,N_5504);
nor U7943 (N_7943,N_4741,N_4587);
xor U7944 (N_7944,N_3498,N_5941);
and U7945 (N_7945,N_5304,N_3618);
and U7946 (N_7946,N_5436,N_3269);
xnor U7947 (N_7947,N_3806,N_5134);
and U7948 (N_7948,N_3416,N_4222);
nor U7949 (N_7949,N_3032,N_4165);
and U7950 (N_7950,N_4569,N_3256);
or U7951 (N_7951,N_5087,N_4891);
and U7952 (N_7952,N_4778,N_4017);
and U7953 (N_7953,N_3859,N_5966);
or U7954 (N_7954,N_5777,N_3012);
or U7955 (N_7955,N_5919,N_5062);
nor U7956 (N_7956,N_5150,N_3795);
xor U7957 (N_7957,N_5160,N_5857);
or U7958 (N_7958,N_4898,N_5850);
nand U7959 (N_7959,N_3518,N_4533);
xor U7960 (N_7960,N_4559,N_3748);
nor U7961 (N_7961,N_4950,N_3835);
or U7962 (N_7962,N_3862,N_4384);
nand U7963 (N_7963,N_5121,N_5858);
nand U7964 (N_7964,N_4153,N_5673);
or U7965 (N_7965,N_4722,N_5597);
and U7966 (N_7966,N_4831,N_3671);
or U7967 (N_7967,N_3373,N_4879);
nand U7968 (N_7968,N_3499,N_4586);
nand U7969 (N_7969,N_5968,N_4965);
nor U7970 (N_7970,N_4751,N_5419);
nor U7971 (N_7971,N_4575,N_3786);
or U7972 (N_7972,N_3213,N_5471);
xnor U7973 (N_7973,N_5072,N_5906);
and U7974 (N_7974,N_4709,N_5003);
or U7975 (N_7975,N_5821,N_4727);
and U7976 (N_7976,N_5456,N_5046);
nand U7977 (N_7977,N_5766,N_4221);
and U7978 (N_7978,N_3472,N_5194);
nand U7979 (N_7979,N_3773,N_3205);
or U7980 (N_7980,N_5676,N_4762);
nor U7981 (N_7981,N_3102,N_4568);
nor U7982 (N_7982,N_5620,N_5710);
or U7983 (N_7983,N_4764,N_3272);
xor U7984 (N_7984,N_4948,N_3993);
and U7985 (N_7985,N_5115,N_3934);
nand U7986 (N_7986,N_3588,N_5332);
or U7987 (N_7987,N_3961,N_5958);
and U7988 (N_7988,N_4015,N_5671);
nand U7989 (N_7989,N_5957,N_3177);
or U7990 (N_7990,N_4705,N_5166);
nor U7991 (N_7991,N_3437,N_3177);
nand U7992 (N_7992,N_3369,N_5531);
and U7993 (N_7993,N_4375,N_3548);
and U7994 (N_7994,N_3320,N_3861);
nand U7995 (N_7995,N_3940,N_5458);
or U7996 (N_7996,N_4186,N_5031);
nand U7997 (N_7997,N_3531,N_4995);
nor U7998 (N_7998,N_5232,N_3023);
and U7999 (N_7999,N_5629,N_4801);
and U8000 (N_8000,N_3409,N_4629);
nand U8001 (N_8001,N_3592,N_4545);
or U8002 (N_8002,N_4886,N_3861);
nor U8003 (N_8003,N_5027,N_5462);
and U8004 (N_8004,N_5491,N_5739);
nor U8005 (N_8005,N_5860,N_4854);
xnor U8006 (N_8006,N_3577,N_5693);
xnor U8007 (N_8007,N_3516,N_4869);
xnor U8008 (N_8008,N_5962,N_3827);
nand U8009 (N_8009,N_5318,N_5696);
and U8010 (N_8010,N_4495,N_5666);
xor U8011 (N_8011,N_5515,N_5360);
nand U8012 (N_8012,N_4126,N_5905);
xnor U8013 (N_8013,N_5229,N_5124);
nand U8014 (N_8014,N_3730,N_5926);
or U8015 (N_8015,N_4665,N_4601);
xnor U8016 (N_8016,N_4204,N_3651);
and U8017 (N_8017,N_5643,N_3964);
nor U8018 (N_8018,N_3438,N_4725);
and U8019 (N_8019,N_5049,N_4285);
xor U8020 (N_8020,N_5756,N_3776);
nand U8021 (N_8021,N_4180,N_4517);
and U8022 (N_8022,N_5844,N_5761);
or U8023 (N_8023,N_5408,N_5401);
nand U8024 (N_8024,N_3072,N_4675);
or U8025 (N_8025,N_3201,N_5472);
nand U8026 (N_8026,N_4984,N_5045);
and U8027 (N_8027,N_4116,N_4016);
xnor U8028 (N_8028,N_3413,N_5772);
nor U8029 (N_8029,N_3190,N_4392);
nand U8030 (N_8030,N_5454,N_4968);
nor U8031 (N_8031,N_5755,N_5840);
nand U8032 (N_8032,N_3090,N_3154);
and U8033 (N_8033,N_4365,N_4977);
or U8034 (N_8034,N_5611,N_3786);
xor U8035 (N_8035,N_3450,N_4546);
or U8036 (N_8036,N_5344,N_5431);
or U8037 (N_8037,N_5711,N_5261);
or U8038 (N_8038,N_4791,N_5452);
xnor U8039 (N_8039,N_5716,N_3360);
and U8040 (N_8040,N_5982,N_4481);
or U8041 (N_8041,N_4791,N_4761);
xnor U8042 (N_8042,N_4867,N_3645);
xnor U8043 (N_8043,N_3877,N_3256);
xnor U8044 (N_8044,N_3567,N_4033);
xnor U8045 (N_8045,N_4061,N_4995);
nor U8046 (N_8046,N_5835,N_3937);
xnor U8047 (N_8047,N_4316,N_4536);
xnor U8048 (N_8048,N_4595,N_3888);
nand U8049 (N_8049,N_5197,N_5368);
xor U8050 (N_8050,N_3512,N_5544);
nor U8051 (N_8051,N_5332,N_5113);
nor U8052 (N_8052,N_5706,N_3128);
nand U8053 (N_8053,N_5349,N_3293);
nand U8054 (N_8054,N_4952,N_3697);
nor U8055 (N_8055,N_5028,N_4670);
and U8056 (N_8056,N_3852,N_5821);
nor U8057 (N_8057,N_5282,N_3277);
nand U8058 (N_8058,N_5484,N_3233);
or U8059 (N_8059,N_5208,N_5270);
nor U8060 (N_8060,N_5093,N_3108);
xnor U8061 (N_8061,N_4807,N_3902);
nand U8062 (N_8062,N_5108,N_4588);
and U8063 (N_8063,N_5183,N_3888);
or U8064 (N_8064,N_5263,N_4625);
nand U8065 (N_8065,N_4751,N_3962);
xnor U8066 (N_8066,N_3922,N_5229);
nand U8067 (N_8067,N_4864,N_3928);
and U8068 (N_8068,N_3362,N_3972);
nor U8069 (N_8069,N_4272,N_5992);
nor U8070 (N_8070,N_3449,N_4952);
nor U8071 (N_8071,N_5841,N_4361);
nand U8072 (N_8072,N_3305,N_4693);
or U8073 (N_8073,N_5694,N_4417);
and U8074 (N_8074,N_5788,N_3887);
and U8075 (N_8075,N_4820,N_3842);
nand U8076 (N_8076,N_5339,N_4896);
or U8077 (N_8077,N_5801,N_5045);
nor U8078 (N_8078,N_5412,N_4953);
or U8079 (N_8079,N_4678,N_4972);
xnor U8080 (N_8080,N_4608,N_4547);
xor U8081 (N_8081,N_5246,N_4973);
and U8082 (N_8082,N_4781,N_3774);
or U8083 (N_8083,N_3423,N_3800);
or U8084 (N_8084,N_3475,N_3611);
xor U8085 (N_8085,N_3654,N_4334);
nor U8086 (N_8086,N_5117,N_5208);
nor U8087 (N_8087,N_4089,N_4266);
xor U8088 (N_8088,N_3558,N_5364);
nand U8089 (N_8089,N_4452,N_3088);
nand U8090 (N_8090,N_4791,N_4315);
nand U8091 (N_8091,N_3469,N_5401);
or U8092 (N_8092,N_3332,N_5547);
and U8093 (N_8093,N_5461,N_5862);
xnor U8094 (N_8094,N_4422,N_5975);
nor U8095 (N_8095,N_5036,N_4194);
nor U8096 (N_8096,N_3088,N_5093);
or U8097 (N_8097,N_5118,N_3606);
and U8098 (N_8098,N_3914,N_5735);
xor U8099 (N_8099,N_5557,N_5552);
and U8100 (N_8100,N_3199,N_4157);
nor U8101 (N_8101,N_4511,N_3616);
or U8102 (N_8102,N_3780,N_4251);
nand U8103 (N_8103,N_4356,N_4687);
nor U8104 (N_8104,N_4126,N_5084);
or U8105 (N_8105,N_4272,N_4634);
nor U8106 (N_8106,N_4511,N_3420);
and U8107 (N_8107,N_4946,N_3208);
nand U8108 (N_8108,N_4288,N_5366);
nand U8109 (N_8109,N_5058,N_4042);
and U8110 (N_8110,N_4655,N_5630);
xnor U8111 (N_8111,N_3540,N_4339);
and U8112 (N_8112,N_3853,N_3647);
nor U8113 (N_8113,N_3419,N_4987);
or U8114 (N_8114,N_3668,N_4360);
nand U8115 (N_8115,N_3013,N_3863);
and U8116 (N_8116,N_5459,N_3272);
xor U8117 (N_8117,N_5505,N_4626);
and U8118 (N_8118,N_5767,N_3769);
and U8119 (N_8119,N_3644,N_3791);
nand U8120 (N_8120,N_4105,N_3060);
or U8121 (N_8121,N_4436,N_5251);
and U8122 (N_8122,N_3078,N_4666);
nand U8123 (N_8123,N_3369,N_5823);
or U8124 (N_8124,N_4513,N_5069);
or U8125 (N_8125,N_3524,N_4269);
and U8126 (N_8126,N_3640,N_4147);
or U8127 (N_8127,N_5481,N_4997);
nor U8128 (N_8128,N_4380,N_4316);
nor U8129 (N_8129,N_4329,N_5316);
xnor U8130 (N_8130,N_5660,N_3731);
nand U8131 (N_8131,N_3459,N_4998);
nor U8132 (N_8132,N_3844,N_3649);
or U8133 (N_8133,N_4748,N_4090);
or U8134 (N_8134,N_4967,N_3110);
xor U8135 (N_8135,N_5956,N_3770);
or U8136 (N_8136,N_5443,N_3205);
xnor U8137 (N_8137,N_3647,N_3843);
nor U8138 (N_8138,N_3990,N_5228);
nor U8139 (N_8139,N_5486,N_5865);
xor U8140 (N_8140,N_3813,N_3549);
or U8141 (N_8141,N_5378,N_5107);
or U8142 (N_8142,N_4910,N_3365);
nor U8143 (N_8143,N_5244,N_4990);
nand U8144 (N_8144,N_4419,N_3846);
xnor U8145 (N_8145,N_4856,N_5260);
or U8146 (N_8146,N_3826,N_5302);
or U8147 (N_8147,N_4748,N_5358);
or U8148 (N_8148,N_3289,N_5196);
xor U8149 (N_8149,N_5565,N_3869);
nor U8150 (N_8150,N_3743,N_4212);
nand U8151 (N_8151,N_5810,N_5563);
or U8152 (N_8152,N_3208,N_5246);
xor U8153 (N_8153,N_4927,N_4724);
nand U8154 (N_8154,N_4560,N_3582);
nand U8155 (N_8155,N_3263,N_4055);
and U8156 (N_8156,N_5656,N_3839);
nor U8157 (N_8157,N_5726,N_5218);
xor U8158 (N_8158,N_3757,N_3085);
or U8159 (N_8159,N_3798,N_3432);
and U8160 (N_8160,N_3669,N_5633);
nor U8161 (N_8161,N_4652,N_5870);
xor U8162 (N_8162,N_4625,N_3609);
and U8163 (N_8163,N_4979,N_4475);
nand U8164 (N_8164,N_4299,N_4284);
and U8165 (N_8165,N_5637,N_4514);
or U8166 (N_8166,N_3758,N_5397);
nor U8167 (N_8167,N_5221,N_4565);
xnor U8168 (N_8168,N_5370,N_5229);
and U8169 (N_8169,N_4407,N_5012);
xor U8170 (N_8170,N_5201,N_5829);
and U8171 (N_8171,N_3958,N_5903);
xor U8172 (N_8172,N_5593,N_4979);
or U8173 (N_8173,N_3091,N_3433);
nand U8174 (N_8174,N_4349,N_5416);
nor U8175 (N_8175,N_5530,N_3680);
nor U8176 (N_8176,N_4172,N_5966);
nand U8177 (N_8177,N_5139,N_3498);
nand U8178 (N_8178,N_4348,N_3068);
nand U8179 (N_8179,N_4889,N_3216);
nor U8180 (N_8180,N_5462,N_3437);
xor U8181 (N_8181,N_3817,N_3823);
nor U8182 (N_8182,N_3668,N_5322);
or U8183 (N_8183,N_5741,N_5522);
nand U8184 (N_8184,N_3491,N_4625);
nor U8185 (N_8185,N_4948,N_4009);
nand U8186 (N_8186,N_5924,N_4555);
nand U8187 (N_8187,N_3901,N_5687);
or U8188 (N_8188,N_5249,N_4769);
and U8189 (N_8189,N_5916,N_4275);
or U8190 (N_8190,N_4858,N_5730);
or U8191 (N_8191,N_5865,N_3348);
xnor U8192 (N_8192,N_3617,N_4553);
xnor U8193 (N_8193,N_4306,N_3264);
nor U8194 (N_8194,N_4214,N_4576);
nand U8195 (N_8195,N_3786,N_3353);
nor U8196 (N_8196,N_5771,N_3149);
nand U8197 (N_8197,N_5570,N_5225);
or U8198 (N_8198,N_4216,N_5486);
xnor U8199 (N_8199,N_3681,N_5389);
and U8200 (N_8200,N_4555,N_5291);
or U8201 (N_8201,N_4669,N_3425);
xnor U8202 (N_8202,N_5348,N_5133);
and U8203 (N_8203,N_3914,N_4341);
or U8204 (N_8204,N_4341,N_3624);
nand U8205 (N_8205,N_3851,N_5867);
and U8206 (N_8206,N_3478,N_3901);
nor U8207 (N_8207,N_3623,N_4306);
or U8208 (N_8208,N_5024,N_5306);
xor U8209 (N_8209,N_4396,N_5700);
nor U8210 (N_8210,N_4137,N_3714);
xnor U8211 (N_8211,N_4322,N_5376);
and U8212 (N_8212,N_5178,N_3620);
nand U8213 (N_8213,N_5412,N_5650);
or U8214 (N_8214,N_5842,N_5118);
xnor U8215 (N_8215,N_5235,N_5073);
and U8216 (N_8216,N_5691,N_4420);
and U8217 (N_8217,N_5604,N_5010);
nor U8218 (N_8218,N_5873,N_4032);
nor U8219 (N_8219,N_3537,N_4971);
nor U8220 (N_8220,N_4298,N_3636);
nand U8221 (N_8221,N_3920,N_4341);
nand U8222 (N_8222,N_3298,N_5799);
and U8223 (N_8223,N_5612,N_3397);
and U8224 (N_8224,N_5685,N_3971);
xor U8225 (N_8225,N_3489,N_3155);
nand U8226 (N_8226,N_3700,N_4409);
or U8227 (N_8227,N_4309,N_5369);
and U8228 (N_8228,N_5796,N_3391);
or U8229 (N_8229,N_4982,N_4475);
nand U8230 (N_8230,N_4744,N_4155);
and U8231 (N_8231,N_3567,N_4785);
nor U8232 (N_8232,N_4527,N_5910);
xnor U8233 (N_8233,N_4543,N_3078);
nor U8234 (N_8234,N_4360,N_4943);
nand U8235 (N_8235,N_3543,N_5470);
and U8236 (N_8236,N_5930,N_4726);
xnor U8237 (N_8237,N_5089,N_3875);
xor U8238 (N_8238,N_5351,N_3568);
xor U8239 (N_8239,N_4162,N_4365);
or U8240 (N_8240,N_4195,N_5493);
or U8241 (N_8241,N_3016,N_5854);
and U8242 (N_8242,N_4054,N_3315);
nand U8243 (N_8243,N_4812,N_4771);
and U8244 (N_8244,N_5742,N_5523);
or U8245 (N_8245,N_4830,N_4078);
nand U8246 (N_8246,N_4691,N_5599);
nor U8247 (N_8247,N_4837,N_4372);
nor U8248 (N_8248,N_4295,N_4938);
nor U8249 (N_8249,N_5983,N_3799);
or U8250 (N_8250,N_3168,N_4383);
xor U8251 (N_8251,N_3779,N_5748);
and U8252 (N_8252,N_5101,N_5210);
nand U8253 (N_8253,N_4288,N_4941);
xor U8254 (N_8254,N_3345,N_5176);
nor U8255 (N_8255,N_3703,N_5460);
or U8256 (N_8256,N_3908,N_3957);
xnor U8257 (N_8257,N_4587,N_4319);
nor U8258 (N_8258,N_4933,N_4177);
and U8259 (N_8259,N_5451,N_5555);
and U8260 (N_8260,N_4922,N_3201);
or U8261 (N_8261,N_5718,N_4120);
nor U8262 (N_8262,N_5753,N_5685);
nor U8263 (N_8263,N_4797,N_5019);
and U8264 (N_8264,N_5622,N_4408);
or U8265 (N_8265,N_5857,N_5608);
and U8266 (N_8266,N_4076,N_3294);
and U8267 (N_8267,N_3492,N_3745);
nor U8268 (N_8268,N_3476,N_4833);
xnor U8269 (N_8269,N_5588,N_4884);
xor U8270 (N_8270,N_4832,N_4581);
nor U8271 (N_8271,N_5071,N_4748);
nand U8272 (N_8272,N_4653,N_3107);
nor U8273 (N_8273,N_5198,N_4727);
xnor U8274 (N_8274,N_4312,N_5533);
and U8275 (N_8275,N_3819,N_5107);
nor U8276 (N_8276,N_4796,N_3009);
or U8277 (N_8277,N_3729,N_5161);
and U8278 (N_8278,N_4988,N_3659);
xor U8279 (N_8279,N_3257,N_4885);
or U8280 (N_8280,N_3520,N_3719);
nand U8281 (N_8281,N_3403,N_4385);
nand U8282 (N_8282,N_4451,N_5822);
nand U8283 (N_8283,N_4270,N_3232);
xnor U8284 (N_8284,N_4618,N_3004);
nor U8285 (N_8285,N_5001,N_5432);
and U8286 (N_8286,N_3534,N_4876);
nand U8287 (N_8287,N_4421,N_4039);
or U8288 (N_8288,N_5422,N_3607);
nor U8289 (N_8289,N_3414,N_4034);
xor U8290 (N_8290,N_4472,N_5252);
and U8291 (N_8291,N_5591,N_4672);
or U8292 (N_8292,N_5819,N_4997);
xnor U8293 (N_8293,N_3762,N_4273);
nor U8294 (N_8294,N_5817,N_5182);
or U8295 (N_8295,N_4791,N_5047);
xor U8296 (N_8296,N_5950,N_5624);
or U8297 (N_8297,N_4085,N_5763);
xnor U8298 (N_8298,N_5252,N_5278);
and U8299 (N_8299,N_3241,N_3100);
xnor U8300 (N_8300,N_4421,N_5694);
or U8301 (N_8301,N_5343,N_3878);
xor U8302 (N_8302,N_3399,N_4963);
xor U8303 (N_8303,N_3363,N_5474);
nor U8304 (N_8304,N_3234,N_5271);
nand U8305 (N_8305,N_3998,N_5287);
nand U8306 (N_8306,N_3812,N_4793);
nand U8307 (N_8307,N_5409,N_4900);
nand U8308 (N_8308,N_5871,N_5367);
and U8309 (N_8309,N_3296,N_4904);
nand U8310 (N_8310,N_3867,N_5624);
nor U8311 (N_8311,N_3511,N_5841);
nor U8312 (N_8312,N_3241,N_3733);
nor U8313 (N_8313,N_3251,N_3425);
xnor U8314 (N_8314,N_4374,N_4409);
xnor U8315 (N_8315,N_3991,N_3366);
or U8316 (N_8316,N_3798,N_3879);
or U8317 (N_8317,N_5541,N_4638);
and U8318 (N_8318,N_3152,N_5211);
or U8319 (N_8319,N_4627,N_4469);
xor U8320 (N_8320,N_3249,N_3738);
and U8321 (N_8321,N_4004,N_5825);
or U8322 (N_8322,N_3385,N_5702);
xor U8323 (N_8323,N_3994,N_5390);
and U8324 (N_8324,N_4277,N_4509);
nor U8325 (N_8325,N_3756,N_5921);
nor U8326 (N_8326,N_5915,N_3392);
nor U8327 (N_8327,N_3742,N_5901);
or U8328 (N_8328,N_3691,N_5483);
xor U8329 (N_8329,N_5299,N_5143);
nand U8330 (N_8330,N_4965,N_5145);
xor U8331 (N_8331,N_5359,N_5498);
nand U8332 (N_8332,N_5192,N_4668);
nand U8333 (N_8333,N_4526,N_4037);
nor U8334 (N_8334,N_4810,N_5895);
nor U8335 (N_8335,N_3790,N_4047);
xnor U8336 (N_8336,N_4880,N_5417);
and U8337 (N_8337,N_3045,N_3515);
nor U8338 (N_8338,N_4184,N_3767);
or U8339 (N_8339,N_3005,N_4384);
nand U8340 (N_8340,N_5449,N_3206);
xnor U8341 (N_8341,N_3969,N_4042);
nand U8342 (N_8342,N_5848,N_4030);
xor U8343 (N_8343,N_4297,N_4565);
and U8344 (N_8344,N_4169,N_5322);
and U8345 (N_8345,N_3665,N_4212);
xor U8346 (N_8346,N_3892,N_3519);
nand U8347 (N_8347,N_5857,N_5646);
nand U8348 (N_8348,N_5463,N_5745);
or U8349 (N_8349,N_5108,N_5221);
and U8350 (N_8350,N_3601,N_3857);
nor U8351 (N_8351,N_3620,N_5044);
and U8352 (N_8352,N_4116,N_3980);
and U8353 (N_8353,N_4390,N_4973);
xor U8354 (N_8354,N_5742,N_3429);
nor U8355 (N_8355,N_3687,N_5367);
nand U8356 (N_8356,N_4959,N_4124);
xnor U8357 (N_8357,N_3222,N_5548);
or U8358 (N_8358,N_3472,N_3616);
or U8359 (N_8359,N_5874,N_3293);
xor U8360 (N_8360,N_4206,N_5525);
nand U8361 (N_8361,N_3822,N_3827);
or U8362 (N_8362,N_5851,N_5552);
nor U8363 (N_8363,N_4546,N_4044);
nand U8364 (N_8364,N_5905,N_4586);
and U8365 (N_8365,N_3665,N_4513);
xor U8366 (N_8366,N_5520,N_4199);
nand U8367 (N_8367,N_4459,N_4423);
xor U8368 (N_8368,N_4361,N_3841);
and U8369 (N_8369,N_4491,N_4053);
nand U8370 (N_8370,N_4608,N_3308);
nor U8371 (N_8371,N_4609,N_4341);
or U8372 (N_8372,N_5683,N_3244);
nand U8373 (N_8373,N_5705,N_3277);
and U8374 (N_8374,N_4491,N_5937);
nand U8375 (N_8375,N_4342,N_5881);
nand U8376 (N_8376,N_3321,N_4892);
or U8377 (N_8377,N_4828,N_5790);
or U8378 (N_8378,N_3286,N_4547);
xor U8379 (N_8379,N_5313,N_5583);
nor U8380 (N_8380,N_3826,N_5895);
nor U8381 (N_8381,N_4704,N_5994);
xor U8382 (N_8382,N_3091,N_4614);
or U8383 (N_8383,N_5427,N_5381);
or U8384 (N_8384,N_4682,N_3619);
and U8385 (N_8385,N_5590,N_4922);
and U8386 (N_8386,N_5929,N_4684);
xnor U8387 (N_8387,N_4129,N_5964);
xor U8388 (N_8388,N_4159,N_4365);
and U8389 (N_8389,N_3583,N_3050);
or U8390 (N_8390,N_3446,N_4113);
xnor U8391 (N_8391,N_3273,N_4121);
xor U8392 (N_8392,N_5330,N_3573);
nand U8393 (N_8393,N_5965,N_3501);
xnor U8394 (N_8394,N_4420,N_4119);
nand U8395 (N_8395,N_3900,N_4334);
xor U8396 (N_8396,N_5710,N_4688);
xor U8397 (N_8397,N_3409,N_3587);
xor U8398 (N_8398,N_4304,N_4822);
and U8399 (N_8399,N_4175,N_5905);
nand U8400 (N_8400,N_4878,N_4692);
and U8401 (N_8401,N_5435,N_5181);
or U8402 (N_8402,N_5601,N_4765);
nand U8403 (N_8403,N_4425,N_3735);
nand U8404 (N_8404,N_3519,N_3821);
nand U8405 (N_8405,N_4918,N_4957);
nor U8406 (N_8406,N_3426,N_5862);
xor U8407 (N_8407,N_5386,N_3634);
or U8408 (N_8408,N_5737,N_4781);
or U8409 (N_8409,N_3762,N_5171);
or U8410 (N_8410,N_4293,N_5018);
and U8411 (N_8411,N_3907,N_5143);
nor U8412 (N_8412,N_5404,N_3699);
xnor U8413 (N_8413,N_4284,N_4071);
or U8414 (N_8414,N_3006,N_4519);
nand U8415 (N_8415,N_3212,N_3319);
nand U8416 (N_8416,N_5295,N_4681);
nand U8417 (N_8417,N_4848,N_5738);
nor U8418 (N_8418,N_3660,N_5551);
nand U8419 (N_8419,N_4920,N_4162);
xor U8420 (N_8420,N_3901,N_5466);
xor U8421 (N_8421,N_4412,N_4956);
nand U8422 (N_8422,N_4060,N_4580);
nand U8423 (N_8423,N_5612,N_5395);
xnor U8424 (N_8424,N_3176,N_4934);
nor U8425 (N_8425,N_4094,N_5041);
and U8426 (N_8426,N_5546,N_4838);
xor U8427 (N_8427,N_5511,N_5299);
xnor U8428 (N_8428,N_3219,N_5100);
nand U8429 (N_8429,N_5388,N_4637);
or U8430 (N_8430,N_3316,N_3354);
xnor U8431 (N_8431,N_5001,N_4883);
or U8432 (N_8432,N_3583,N_4399);
xnor U8433 (N_8433,N_5501,N_5480);
or U8434 (N_8434,N_4129,N_4371);
nand U8435 (N_8435,N_4007,N_3618);
xor U8436 (N_8436,N_5299,N_4988);
nor U8437 (N_8437,N_4534,N_5255);
and U8438 (N_8438,N_5809,N_4760);
xnor U8439 (N_8439,N_4724,N_3857);
nor U8440 (N_8440,N_5576,N_5692);
nand U8441 (N_8441,N_5151,N_5180);
xnor U8442 (N_8442,N_4279,N_4259);
and U8443 (N_8443,N_3422,N_5679);
nor U8444 (N_8444,N_3042,N_3274);
xor U8445 (N_8445,N_4492,N_4331);
or U8446 (N_8446,N_5140,N_5174);
nand U8447 (N_8447,N_4466,N_3460);
nand U8448 (N_8448,N_3118,N_4737);
and U8449 (N_8449,N_4702,N_3064);
and U8450 (N_8450,N_3590,N_3160);
nor U8451 (N_8451,N_5086,N_5645);
xor U8452 (N_8452,N_5500,N_4683);
nand U8453 (N_8453,N_4793,N_3383);
nor U8454 (N_8454,N_5065,N_4049);
and U8455 (N_8455,N_5691,N_5130);
nor U8456 (N_8456,N_5961,N_3326);
and U8457 (N_8457,N_5983,N_4879);
and U8458 (N_8458,N_4971,N_4912);
or U8459 (N_8459,N_4172,N_3353);
nand U8460 (N_8460,N_5131,N_4201);
and U8461 (N_8461,N_4031,N_5447);
nand U8462 (N_8462,N_3935,N_4766);
xnor U8463 (N_8463,N_5402,N_3383);
nand U8464 (N_8464,N_4492,N_5986);
nand U8465 (N_8465,N_3570,N_4119);
nor U8466 (N_8466,N_5768,N_3579);
and U8467 (N_8467,N_4997,N_5716);
xor U8468 (N_8468,N_3162,N_5483);
nand U8469 (N_8469,N_5950,N_5248);
nor U8470 (N_8470,N_3611,N_3848);
and U8471 (N_8471,N_3639,N_3959);
and U8472 (N_8472,N_3159,N_5413);
xor U8473 (N_8473,N_4092,N_3226);
xnor U8474 (N_8474,N_5343,N_3322);
nor U8475 (N_8475,N_3194,N_3192);
or U8476 (N_8476,N_4770,N_5156);
xnor U8477 (N_8477,N_4985,N_4738);
xnor U8478 (N_8478,N_5981,N_5674);
and U8479 (N_8479,N_3593,N_4305);
or U8480 (N_8480,N_5528,N_3380);
or U8481 (N_8481,N_3393,N_4787);
or U8482 (N_8482,N_3387,N_4568);
and U8483 (N_8483,N_3971,N_5330);
or U8484 (N_8484,N_5350,N_3808);
nand U8485 (N_8485,N_4075,N_5520);
nor U8486 (N_8486,N_4168,N_3409);
nand U8487 (N_8487,N_5256,N_4808);
and U8488 (N_8488,N_5117,N_5754);
or U8489 (N_8489,N_5116,N_5401);
nor U8490 (N_8490,N_5122,N_3725);
nand U8491 (N_8491,N_4735,N_5867);
and U8492 (N_8492,N_4428,N_4313);
xor U8493 (N_8493,N_3639,N_3297);
nor U8494 (N_8494,N_4572,N_5443);
nand U8495 (N_8495,N_3386,N_5073);
and U8496 (N_8496,N_3708,N_4360);
nand U8497 (N_8497,N_4536,N_3481);
xnor U8498 (N_8498,N_4812,N_4665);
and U8499 (N_8499,N_5075,N_3466);
xor U8500 (N_8500,N_4207,N_4395);
and U8501 (N_8501,N_5972,N_5854);
nand U8502 (N_8502,N_4678,N_3609);
nand U8503 (N_8503,N_4167,N_3966);
and U8504 (N_8504,N_4311,N_3162);
and U8505 (N_8505,N_5301,N_5816);
and U8506 (N_8506,N_4977,N_4862);
nand U8507 (N_8507,N_4988,N_5291);
nand U8508 (N_8508,N_5613,N_4521);
and U8509 (N_8509,N_4351,N_5617);
or U8510 (N_8510,N_5024,N_5428);
xor U8511 (N_8511,N_3346,N_5898);
xnor U8512 (N_8512,N_3371,N_5333);
nor U8513 (N_8513,N_5257,N_4313);
or U8514 (N_8514,N_5169,N_4684);
xor U8515 (N_8515,N_3057,N_4127);
nand U8516 (N_8516,N_5857,N_5008);
and U8517 (N_8517,N_4021,N_5753);
xnor U8518 (N_8518,N_3548,N_4657);
nor U8519 (N_8519,N_5308,N_5184);
nand U8520 (N_8520,N_3753,N_3389);
and U8521 (N_8521,N_5841,N_4355);
nor U8522 (N_8522,N_3342,N_3072);
nor U8523 (N_8523,N_4397,N_4642);
and U8524 (N_8524,N_4239,N_4512);
nor U8525 (N_8525,N_3500,N_3511);
xnor U8526 (N_8526,N_5029,N_5176);
nor U8527 (N_8527,N_3035,N_5142);
or U8528 (N_8528,N_3196,N_3976);
xor U8529 (N_8529,N_3176,N_3986);
or U8530 (N_8530,N_3986,N_3935);
xnor U8531 (N_8531,N_5580,N_5346);
or U8532 (N_8532,N_4051,N_3456);
xor U8533 (N_8533,N_5991,N_4716);
xor U8534 (N_8534,N_3693,N_5134);
or U8535 (N_8535,N_5480,N_5534);
xor U8536 (N_8536,N_3186,N_3166);
xor U8537 (N_8537,N_3880,N_3209);
nor U8538 (N_8538,N_3315,N_5681);
nor U8539 (N_8539,N_3974,N_5463);
nand U8540 (N_8540,N_3270,N_4055);
xor U8541 (N_8541,N_3555,N_4487);
xor U8542 (N_8542,N_3771,N_4921);
nor U8543 (N_8543,N_5654,N_4770);
nand U8544 (N_8544,N_3539,N_3946);
and U8545 (N_8545,N_3053,N_3799);
xnor U8546 (N_8546,N_4917,N_5900);
nand U8547 (N_8547,N_5182,N_3213);
and U8548 (N_8548,N_5897,N_4175);
nand U8549 (N_8549,N_4227,N_4182);
or U8550 (N_8550,N_5990,N_5175);
or U8551 (N_8551,N_3484,N_4992);
nor U8552 (N_8552,N_3823,N_4759);
and U8553 (N_8553,N_5464,N_4327);
nand U8554 (N_8554,N_4077,N_3673);
and U8555 (N_8555,N_5473,N_5045);
nor U8556 (N_8556,N_3836,N_3854);
xor U8557 (N_8557,N_3795,N_5774);
nor U8558 (N_8558,N_4923,N_5257);
nand U8559 (N_8559,N_4426,N_3149);
nand U8560 (N_8560,N_5335,N_3117);
nand U8561 (N_8561,N_4194,N_3334);
or U8562 (N_8562,N_3213,N_3262);
and U8563 (N_8563,N_5786,N_5848);
xnor U8564 (N_8564,N_4483,N_5982);
or U8565 (N_8565,N_4188,N_3846);
xor U8566 (N_8566,N_3488,N_3224);
xor U8567 (N_8567,N_5773,N_3147);
xnor U8568 (N_8568,N_4061,N_5944);
and U8569 (N_8569,N_4105,N_5276);
nor U8570 (N_8570,N_4812,N_5229);
and U8571 (N_8571,N_5670,N_3022);
or U8572 (N_8572,N_4302,N_5813);
nand U8573 (N_8573,N_5391,N_5703);
and U8574 (N_8574,N_5788,N_3618);
nand U8575 (N_8575,N_4351,N_5360);
and U8576 (N_8576,N_4426,N_3228);
xnor U8577 (N_8577,N_3253,N_4324);
xnor U8578 (N_8578,N_4043,N_5179);
nand U8579 (N_8579,N_5668,N_5194);
nor U8580 (N_8580,N_3340,N_3293);
xor U8581 (N_8581,N_4503,N_4634);
nand U8582 (N_8582,N_5585,N_4988);
xnor U8583 (N_8583,N_5962,N_3557);
nor U8584 (N_8584,N_4437,N_3579);
nand U8585 (N_8585,N_3187,N_3366);
or U8586 (N_8586,N_3136,N_4342);
or U8587 (N_8587,N_5616,N_4781);
nor U8588 (N_8588,N_4976,N_4826);
and U8589 (N_8589,N_4028,N_4852);
xnor U8590 (N_8590,N_5539,N_3040);
nand U8591 (N_8591,N_3035,N_5108);
or U8592 (N_8592,N_4308,N_4056);
nand U8593 (N_8593,N_5207,N_3590);
nand U8594 (N_8594,N_4911,N_5111);
or U8595 (N_8595,N_3876,N_5387);
or U8596 (N_8596,N_5024,N_5956);
and U8597 (N_8597,N_3090,N_5381);
nor U8598 (N_8598,N_4919,N_3717);
or U8599 (N_8599,N_3306,N_4517);
and U8600 (N_8600,N_3027,N_5318);
nor U8601 (N_8601,N_4674,N_4416);
or U8602 (N_8602,N_4113,N_5399);
and U8603 (N_8603,N_3616,N_3283);
xor U8604 (N_8604,N_4528,N_3103);
or U8605 (N_8605,N_4577,N_3373);
or U8606 (N_8606,N_4033,N_3561);
xnor U8607 (N_8607,N_3005,N_4300);
and U8608 (N_8608,N_5168,N_5329);
or U8609 (N_8609,N_3180,N_4675);
or U8610 (N_8610,N_3904,N_4138);
and U8611 (N_8611,N_4313,N_5818);
xnor U8612 (N_8612,N_5013,N_4839);
nand U8613 (N_8613,N_3230,N_3195);
or U8614 (N_8614,N_4848,N_4655);
xor U8615 (N_8615,N_3506,N_3720);
xor U8616 (N_8616,N_5668,N_5613);
and U8617 (N_8617,N_4073,N_3648);
nand U8618 (N_8618,N_5259,N_3730);
and U8619 (N_8619,N_4644,N_3546);
or U8620 (N_8620,N_5091,N_3733);
nor U8621 (N_8621,N_5966,N_3536);
xor U8622 (N_8622,N_3600,N_5829);
nand U8623 (N_8623,N_4042,N_4244);
or U8624 (N_8624,N_4220,N_5857);
nor U8625 (N_8625,N_5173,N_5486);
nand U8626 (N_8626,N_4840,N_4976);
nor U8627 (N_8627,N_5468,N_3328);
xor U8628 (N_8628,N_5768,N_3810);
and U8629 (N_8629,N_3654,N_5399);
nor U8630 (N_8630,N_4700,N_5567);
xnor U8631 (N_8631,N_5974,N_5773);
nor U8632 (N_8632,N_5046,N_3107);
nor U8633 (N_8633,N_4285,N_4394);
nand U8634 (N_8634,N_4615,N_5609);
and U8635 (N_8635,N_3498,N_4736);
nand U8636 (N_8636,N_4903,N_4453);
xnor U8637 (N_8637,N_4110,N_4940);
xor U8638 (N_8638,N_4887,N_4871);
xor U8639 (N_8639,N_4831,N_5894);
or U8640 (N_8640,N_4840,N_3829);
nor U8641 (N_8641,N_5515,N_4753);
nor U8642 (N_8642,N_5474,N_4861);
or U8643 (N_8643,N_4245,N_4150);
nand U8644 (N_8644,N_5318,N_3539);
or U8645 (N_8645,N_3513,N_4558);
and U8646 (N_8646,N_3922,N_4275);
or U8647 (N_8647,N_5060,N_4256);
or U8648 (N_8648,N_4900,N_3612);
and U8649 (N_8649,N_4752,N_5325);
xnor U8650 (N_8650,N_3204,N_5323);
nor U8651 (N_8651,N_4566,N_3738);
xnor U8652 (N_8652,N_5999,N_3140);
xor U8653 (N_8653,N_4186,N_5908);
or U8654 (N_8654,N_5783,N_4359);
nor U8655 (N_8655,N_5533,N_3705);
or U8656 (N_8656,N_4518,N_3162);
xnor U8657 (N_8657,N_3198,N_3751);
nand U8658 (N_8658,N_3988,N_5092);
nand U8659 (N_8659,N_5881,N_3282);
xor U8660 (N_8660,N_5655,N_5238);
and U8661 (N_8661,N_5603,N_4018);
nor U8662 (N_8662,N_5241,N_4594);
nand U8663 (N_8663,N_3946,N_5049);
or U8664 (N_8664,N_3138,N_4092);
nor U8665 (N_8665,N_5588,N_4469);
and U8666 (N_8666,N_4591,N_4538);
or U8667 (N_8667,N_4159,N_3218);
and U8668 (N_8668,N_3125,N_5375);
or U8669 (N_8669,N_5849,N_4937);
and U8670 (N_8670,N_3148,N_3218);
or U8671 (N_8671,N_4907,N_3933);
or U8672 (N_8672,N_3150,N_4926);
and U8673 (N_8673,N_5732,N_5319);
xor U8674 (N_8674,N_4775,N_4211);
and U8675 (N_8675,N_4693,N_3372);
xor U8676 (N_8676,N_3595,N_4224);
and U8677 (N_8677,N_3412,N_4691);
xor U8678 (N_8678,N_3187,N_5068);
or U8679 (N_8679,N_5321,N_5022);
xor U8680 (N_8680,N_4161,N_4582);
nand U8681 (N_8681,N_5819,N_4304);
and U8682 (N_8682,N_5005,N_4235);
or U8683 (N_8683,N_3150,N_3992);
nand U8684 (N_8684,N_3921,N_4749);
nor U8685 (N_8685,N_4933,N_5667);
xnor U8686 (N_8686,N_3640,N_3019);
nand U8687 (N_8687,N_4318,N_5666);
or U8688 (N_8688,N_4226,N_4050);
nand U8689 (N_8689,N_4922,N_4316);
nor U8690 (N_8690,N_3925,N_4612);
xor U8691 (N_8691,N_4997,N_5010);
nor U8692 (N_8692,N_4619,N_5514);
nor U8693 (N_8693,N_4958,N_3531);
and U8694 (N_8694,N_3679,N_5199);
and U8695 (N_8695,N_5781,N_3893);
nor U8696 (N_8696,N_5542,N_4528);
xor U8697 (N_8697,N_4936,N_5502);
xnor U8698 (N_8698,N_3795,N_4979);
nor U8699 (N_8699,N_4705,N_3606);
nand U8700 (N_8700,N_4710,N_4287);
and U8701 (N_8701,N_4134,N_4350);
and U8702 (N_8702,N_3937,N_3719);
or U8703 (N_8703,N_3722,N_3889);
or U8704 (N_8704,N_3488,N_4558);
and U8705 (N_8705,N_4327,N_5599);
and U8706 (N_8706,N_5328,N_4265);
or U8707 (N_8707,N_4324,N_5998);
nand U8708 (N_8708,N_4616,N_4284);
nand U8709 (N_8709,N_5721,N_3333);
nand U8710 (N_8710,N_5517,N_3368);
or U8711 (N_8711,N_4532,N_4327);
xor U8712 (N_8712,N_5691,N_4779);
xor U8713 (N_8713,N_4711,N_5256);
and U8714 (N_8714,N_3267,N_5675);
xor U8715 (N_8715,N_4593,N_3688);
and U8716 (N_8716,N_4828,N_3742);
nand U8717 (N_8717,N_3738,N_5858);
xor U8718 (N_8718,N_3602,N_3576);
and U8719 (N_8719,N_4142,N_4546);
or U8720 (N_8720,N_5625,N_3946);
xnor U8721 (N_8721,N_5104,N_4414);
and U8722 (N_8722,N_3516,N_5047);
nand U8723 (N_8723,N_5583,N_3478);
and U8724 (N_8724,N_5303,N_4883);
xnor U8725 (N_8725,N_5140,N_5250);
xnor U8726 (N_8726,N_5236,N_5295);
nand U8727 (N_8727,N_4129,N_3921);
or U8728 (N_8728,N_5915,N_4280);
or U8729 (N_8729,N_3533,N_3422);
xor U8730 (N_8730,N_4226,N_5828);
nand U8731 (N_8731,N_4200,N_5070);
nand U8732 (N_8732,N_4143,N_5247);
nor U8733 (N_8733,N_3785,N_5547);
nand U8734 (N_8734,N_5830,N_4328);
nor U8735 (N_8735,N_3927,N_3442);
nor U8736 (N_8736,N_4998,N_3936);
nor U8737 (N_8737,N_3193,N_3389);
and U8738 (N_8738,N_5185,N_4872);
nor U8739 (N_8739,N_4677,N_5144);
or U8740 (N_8740,N_3991,N_5372);
nand U8741 (N_8741,N_5654,N_3011);
or U8742 (N_8742,N_5196,N_5579);
or U8743 (N_8743,N_3581,N_4896);
or U8744 (N_8744,N_3629,N_5591);
xnor U8745 (N_8745,N_3786,N_5989);
and U8746 (N_8746,N_5381,N_5442);
or U8747 (N_8747,N_3025,N_3505);
and U8748 (N_8748,N_5321,N_5395);
and U8749 (N_8749,N_5404,N_3223);
nor U8750 (N_8750,N_4247,N_3644);
xor U8751 (N_8751,N_3216,N_5174);
and U8752 (N_8752,N_5430,N_4802);
and U8753 (N_8753,N_3914,N_3369);
nand U8754 (N_8754,N_5348,N_3908);
or U8755 (N_8755,N_3245,N_5251);
or U8756 (N_8756,N_4367,N_3568);
xor U8757 (N_8757,N_3631,N_3192);
or U8758 (N_8758,N_5054,N_4941);
or U8759 (N_8759,N_5406,N_3179);
nand U8760 (N_8760,N_4864,N_5680);
xor U8761 (N_8761,N_4794,N_4890);
nor U8762 (N_8762,N_5171,N_3177);
xnor U8763 (N_8763,N_5238,N_3326);
or U8764 (N_8764,N_5220,N_4070);
nand U8765 (N_8765,N_5096,N_4670);
xor U8766 (N_8766,N_4414,N_4233);
or U8767 (N_8767,N_3044,N_5860);
and U8768 (N_8768,N_3421,N_5266);
nand U8769 (N_8769,N_4509,N_3821);
or U8770 (N_8770,N_4160,N_4075);
and U8771 (N_8771,N_3359,N_4378);
nand U8772 (N_8772,N_5652,N_5801);
or U8773 (N_8773,N_3481,N_4809);
or U8774 (N_8774,N_3829,N_5692);
nor U8775 (N_8775,N_5675,N_3351);
nand U8776 (N_8776,N_5246,N_3194);
xor U8777 (N_8777,N_3898,N_5089);
xnor U8778 (N_8778,N_3956,N_4149);
xnor U8779 (N_8779,N_3410,N_5168);
nand U8780 (N_8780,N_4599,N_5187);
nor U8781 (N_8781,N_5477,N_5211);
and U8782 (N_8782,N_5995,N_3238);
or U8783 (N_8783,N_4523,N_4977);
and U8784 (N_8784,N_3621,N_4965);
xnor U8785 (N_8785,N_3345,N_5046);
or U8786 (N_8786,N_5467,N_5261);
and U8787 (N_8787,N_4754,N_5877);
nor U8788 (N_8788,N_5613,N_4265);
xnor U8789 (N_8789,N_4973,N_4208);
nand U8790 (N_8790,N_3888,N_3044);
nor U8791 (N_8791,N_3769,N_5007);
and U8792 (N_8792,N_3205,N_4789);
xnor U8793 (N_8793,N_4518,N_3409);
or U8794 (N_8794,N_5942,N_3158);
nand U8795 (N_8795,N_4369,N_4183);
and U8796 (N_8796,N_5699,N_3816);
xnor U8797 (N_8797,N_5515,N_4393);
xnor U8798 (N_8798,N_5618,N_5194);
nor U8799 (N_8799,N_4479,N_5569);
and U8800 (N_8800,N_5142,N_5618);
and U8801 (N_8801,N_4462,N_3399);
or U8802 (N_8802,N_3908,N_5440);
nor U8803 (N_8803,N_5250,N_4676);
xnor U8804 (N_8804,N_4298,N_4634);
or U8805 (N_8805,N_5786,N_5317);
and U8806 (N_8806,N_3156,N_4114);
and U8807 (N_8807,N_3869,N_3167);
and U8808 (N_8808,N_5722,N_5632);
xor U8809 (N_8809,N_4115,N_4261);
nand U8810 (N_8810,N_3099,N_4010);
nor U8811 (N_8811,N_3722,N_4072);
nand U8812 (N_8812,N_5564,N_5909);
nor U8813 (N_8813,N_5623,N_4642);
nand U8814 (N_8814,N_5018,N_5268);
and U8815 (N_8815,N_3868,N_5992);
nor U8816 (N_8816,N_4524,N_3068);
and U8817 (N_8817,N_3731,N_5183);
or U8818 (N_8818,N_3979,N_4893);
and U8819 (N_8819,N_5057,N_4814);
nand U8820 (N_8820,N_4981,N_4097);
and U8821 (N_8821,N_4377,N_3624);
and U8822 (N_8822,N_5855,N_3606);
nor U8823 (N_8823,N_3124,N_4734);
or U8824 (N_8824,N_3472,N_4503);
and U8825 (N_8825,N_5833,N_3161);
nand U8826 (N_8826,N_3003,N_3869);
xnor U8827 (N_8827,N_4263,N_3910);
nor U8828 (N_8828,N_4827,N_4501);
nand U8829 (N_8829,N_4069,N_5052);
xor U8830 (N_8830,N_5050,N_3286);
xor U8831 (N_8831,N_3520,N_5906);
and U8832 (N_8832,N_3469,N_5029);
xnor U8833 (N_8833,N_3128,N_5833);
nand U8834 (N_8834,N_4203,N_5759);
nand U8835 (N_8835,N_3534,N_3775);
nand U8836 (N_8836,N_3985,N_5854);
nand U8837 (N_8837,N_3566,N_4189);
xor U8838 (N_8838,N_4347,N_4378);
or U8839 (N_8839,N_5345,N_4686);
nor U8840 (N_8840,N_3576,N_3206);
and U8841 (N_8841,N_3202,N_4209);
and U8842 (N_8842,N_5270,N_5445);
and U8843 (N_8843,N_4982,N_3408);
nand U8844 (N_8844,N_3995,N_4175);
nor U8845 (N_8845,N_3470,N_5599);
nand U8846 (N_8846,N_3754,N_3002);
xnor U8847 (N_8847,N_4289,N_3603);
xnor U8848 (N_8848,N_4073,N_5132);
or U8849 (N_8849,N_5219,N_5749);
or U8850 (N_8850,N_3398,N_3726);
xnor U8851 (N_8851,N_5905,N_3295);
xnor U8852 (N_8852,N_3793,N_4516);
and U8853 (N_8853,N_4389,N_3916);
nand U8854 (N_8854,N_4825,N_4674);
xor U8855 (N_8855,N_5289,N_4796);
nand U8856 (N_8856,N_3655,N_3745);
nor U8857 (N_8857,N_3579,N_3178);
nor U8858 (N_8858,N_4669,N_3852);
or U8859 (N_8859,N_4052,N_4770);
nand U8860 (N_8860,N_3098,N_4968);
nor U8861 (N_8861,N_5509,N_5979);
or U8862 (N_8862,N_4156,N_3692);
nor U8863 (N_8863,N_3210,N_4259);
nand U8864 (N_8864,N_3570,N_4935);
nor U8865 (N_8865,N_5366,N_4060);
or U8866 (N_8866,N_5587,N_3921);
nor U8867 (N_8867,N_3900,N_4448);
nand U8868 (N_8868,N_3736,N_5063);
nand U8869 (N_8869,N_5710,N_4385);
or U8870 (N_8870,N_5876,N_4729);
xor U8871 (N_8871,N_3730,N_4327);
and U8872 (N_8872,N_5335,N_3532);
or U8873 (N_8873,N_5173,N_4777);
nand U8874 (N_8874,N_3896,N_5108);
nor U8875 (N_8875,N_5210,N_4020);
nor U8876 (N_8876,N_4147,N_4653);
and U8877 (N_8877,N_3405,N_5678);
nand U8878 (N_8878,N_4621,N_4014);
or U8879 (N_8879,N_4745,N_5336);
and U8880 (N_8880,N_5569,N_3189);
nand U8881 (N_8881,N_5104,N_3016);
xor U8882 (N_8882,N_4912,N_4526);
nand U8883 (N_8883,N_4164,N_5010);
nand U8884 (N_8884,N_3100,N_3382);
xor U8885 (N_8885,N_4723,N_4115);
nor U8886 (N_8886,N_4988,N_4810);
and U8887 (N_8887,N_5662,N_5165);
or U8888 (N_8888,N_3508,N_5005);
xnor U8889 (N_8889,N_3102,N_5769);
xor U8890 (N_8890,N_5073,N_3605);
nand U8891 (N_8891,N_5080,N_3840);
and U8892 (N_8892,N_3985,N_4599);
or U8893 (N_8893,N_5865,N_5022);
and U8894 (N_8894,N_4117,N_4229);
nor U8895 (N_8895,N_4203,N_3418);
nor U8896 (N_8896,N_5700,N_3178);
nor U8897 (N_8897,N_3067,N_4391);
and U8898 (N_8898,N_5708,N_4488);
or U8899 (N_8899,N_4837,N_3390);
xnor U8900 (N_8900,N_3804,N_5752);
or U8901 (N_8901,N_4921,N_5873);
or U8902 (N_8902,N_4118,N_3548);
nor U8903 (N_8903,N_4557,N_3795);
nor U8904 (N_8904,N_4917,N_4073);
and U8905 (N_8905,N_3007,N_5463);
nor U8906 (N_8906,N_3616,N_5441);
or U8907 (N_8907,N_3789,N_4031);
xnor U8908 (N_8908,N_4939,N_5236);
nor U8909 (N_8909,N_4036,N_5525);
or U8910 (N_8910,N_4299,N_5487);
nand U8911 (N_8911,N_3141,N_4922);
or U8912 (N_8912,N_4119,N_4628);
or U8913 (N_8913,N_5833,N_5043);
nor U8914 (N_8914,N_4027,N_3186);
nand U8915 (N_8915,N_4520,N_3404);
or U8916 (N_8916,N_5311,N_4553);
xnor U8917 (N_8917,N_4377,N_3423);
xor U8918 (N_8918,N_4473,N_5763);
xnor U8919 (N_8919,N_3588,N_4325);
nor U8920 (N_8920,N_4968,N_3181);
xor U8921 (N_8921,N_5677,N_3719);
xor U8922 (N_8922,N_5096,N_3782);
and U8923 (N_8923,N_4780,N_3262);
nand U8924 (N_8924,N_5329,N_4657);
or U8925 (N_8925,N_4244,N_3371);
xor U8926 (N_8926,N_5742,N_4549);
nand U8927 (N_8927,N_3876,N_4653);
xnor U8928 (N_8928,N_5476,N_4165);
nand U8929 (N_8929,N_5907,N_3418);
or U8930 (N_8930,N_5679,N_4387);
nand U8931 (N_8931,N_3278,N_3480);
xnor U8932 (N_8932,N_4840,N_4212);
or U8933 (N_8933,N_4112,N_3809);
or U8934 (N_8934,N_3364,N_3674);
and U8935 (N_8935,N_4236,N_3815);
nor U8936 (N_8936,N_5243,N_5824);
xnor U8937 (N_8937,N_3612,N_4963);
nand U8938 (N_8938,N_3282,N_4412);
nand U8939 (N_8939,N_3499,N_4990);
xor U8940 (N_8940,N_3277,N_5140);
xnor U8941 (N_8941,N_3176,N_4666);
or U8942 (N_8942,N_4697,N_4796);
nor U8943 (N_8943,N_5476,N_3030);
and U8944 (N_8944,N_4615,N_4074);
xnor U8945 (N_8945,N_4558,N_3826);
nor U8946 (N_8946,N_4325,N_4889);
nand U8947 (N_8947,N_5164,N_4587);
xor U8948 (N_8948,N_5111,N_5662);
xor U8949 (N_8949,N_3605,N_3472);
nor U8950 (N_8950,N_4247,N_3017);
xor U8951 (N_8951,N_3027,N_4644);
xor U8952 (N_8952,N_3613,N_3183);
and U8953 (N_8953,N_3145,N_3998);
nand U8954 (N_8954,N_5949,N_4189);
xnor U8955 (N_8955,N_3813,N_4414);
or U8956 (N_8956,N_3548,N_5127);
and U8957 (N_8957,N_5321,N_4220);
nand U8958 (N_8958,N_5999,N_5247);
nand U8959 (N_8959,N_4435,N_4838);
or U8960 (N_8960,N_5937,N_5538);
or U8961 (N_8961,N_5073,N_5519);
or U8962 (N_8962,N_5219,N_5600);
or U8963 (N_8963,N_3346,N_5622);
or U8964 (N_8964,N_5749,N_3406);
nor U8965 (N_8965,N_5704,N_3226);
nor U8966 (N_8966,N_5780,N_4168);
xnor U8967 (N_8967,N_4252,N_4976);
nor U8968 (N_8968,N_3060,N_4538);
and U8969 (N_8969,N_4251,N_4137);
and U8970 (N_8970,N_4240,N_4006);
and U8971 (N_8971,N_4477,N_3038);
or U8972 (N_8972,N_4081,N_4437);
and U8973 (N_8973,N_5478,N_4448);
or U8974 (N_8974,N_4184,N_3219);
nand U8975 (N_8975,N_4897,N_3540);
or U8976 (N_8976,N_3776,N_5145);
or U8977 (N_8977,N_4540,N_5682);
and U8978 (N_8978,N_5720,N_4352);
and U8979 (N_8979,N_5520,N_4983);
nand U8980 (N_8980,N_5955,N_3074);
nor U8981 (N_8981,N_5123,N_4143);
and U8982 (N_8982,N_5374,N_5646);
nand U8983 (N_8983,N_3319,N_4357);
nor U8984 (N_8984,N_4055,N_5290);
and U8985 (N_8985,N_3667,N_3060);
or U8986 (N_8986,N_4041,N_3959);
nand U8987 (N_8987,N_5522,N_5026);
nor U8988 (N_8988,N_4281,N_3202);
nand U8989 (N_8989,N_4484,N_3664);
nand U8990 (N_8990,N_3414,N_5044);
and U8991 (N_8991,N_5385,N_3929);
nand U8992 (N_8992,N_3626,N_4720);
or U8993 (N_8993,N_3002,N_3960);
and U8994 (N_8994,N_3948,N_3760);
xnor U8995 (N_8995,N_4276,N_5414);
xor U8996 (N_8996,N_3398,N_5626);
or U8997 (N_8997,N_4343,N_3561);
and U8998 (N_8998,N_3558,N_3001);
or U8999 (N_8999,N_3709,N_3233);
nor U9000 (N_9000,N_7478,N_7303);
xor U9001 (N_9001,N_6823,N_7875);
nand U9002 (N_9002,N_7445,N_8050);
nand U9003 (N_9003,N_8773,N_7547);
or U9004 (N_9004,N_7997,N_6187);
nor U9005 (N_9005,N_8019,N_8783);
nand U9006 (N_9006,N_6092,N_8674);
and U9007 (N_9007,N_8653,N_6000);
nor U9008 (N_9008,N_8903,N_7385);
and U9009 (N_9009,N_7496,N_8741);
or U9010 (N_9010,N_8716,N_7971);
nor U9011 (N_9011,N_7325,N_7469);
nor U9012 (N_9012,N_6393,N_8769);
or U9013 (N_9013,N_6637,N_6297);
nor U9014 (N_9014,N_7017,N_7881);
nor U9015 (N_9015,N_7624,N_8968);
xor U9016 (N_9016,N_8371,N_7969);
or U9017 (N_9017,N_6373,N_6719);
and U9018 (N_9018,N_6062,N_8486);
or U9019 (N_9019,N_6327,N_6502);
xnor U9020 (N_9020,N_6715,N_7336);
nand U9021 (N_9021,N_6009,N_8384);
and U9022 (N_9022,N_6809,N_7748);
or U9023 (N_9023,N_6237,N_8094);
or U9024 (N_9024,N_6457,N_6850);
xnor U9025 (N_9025,N_8839,N_6467);
and U9026 (N_9026,N_7894,N_8591);
nand U9027 (N_9027,N_7514,N_6746);
or U9028 (N_9028,N_6911,N_7441);
nor U9029 (N_9029,N_6053,N_8363);
nand U9030 (N_9030,N_7225,N_7529);
and U9031 (N_9031,N_7028,N_8237);
xnor U9032 (N_9032,N_7286,N_8836);
and U9033 (N_9033,N_6376,N_6822);
and U9034 (N_9034,N_7470,N_8243);
or U9035 (N_9035,N_8885,N_6937);
nor U9036 (N_9036,N_6930,N_8712);
or U9037 (N_9037,N_6088,N_6303);
nand U9038 (N_9038,N_8487,N_7666);
or U9039 (N_9039,N_8660,N_7690);
nor U9040 (N_9040,N_6029,N_8454);
nand U9041 (N_9041,N_6629,N_6131);
nor U9042 (N_9042,N_6154,N_6568);
nand U9043 (N_9043,N_8075,N_6331);
or U9044 (N_9044,N_7981,N_7835);
nor U9045 (N_9045,N_6641,N_7825);
and U9046 (N_9046,N_8684,N_8287);
xor U9047 (N_9047,N_7412,N_6229);
nor U9048 (N_9048,N_8328,N_8303);
nand U9049 (N_9049,N_6898,N_7654);
or U9050 (N_9050,N_7551,N_7783);
nor U9051 (N_9051,N_6665,N_6804);
nor U9052 (N_9052,N_6343,N_7903);
nand U9053 (N_9053,N_7192,N_8664);
or U9054 (N_9054,N_7570,N_7444);
xor U9055 (N_9055,N_6946,N_7956);
nand U9056 (N_9056,N_7952,N_6975);
nor U9057 (N_9057,N_6864,N_7662);
or U9058 (N_9058,N_7697,N_6744);
nand U9059 (N_9059,N_6006,N_8045);
nor U9060 (N_9060,N_7269,N_6593);
xor U9061 (N_9061,N_8990,N_7837);
nor U9062 (N_9062,N_8670,N_7241);
and U9063 (N_9063,N_7742,N_6477);
nor U9064 (N_9064,N_8085,N_8004);
xor U9065 (N_9065,N_7562,N_7647);
and U9066 (N_9066,N_7129,N_8008);
nor U9067 (N_9067,N_6957,N_8060);
xor U9068 (N_9068,N_7604,N_6535);
xnor U9069 (N_9069,N_8518,N_6033);
or U9070 (N_9070,N_8582,N_6623);
xnor U9071 (N_9071,N_6317,N_8629);
or U9072 (N_9072,N_8809,N_8916);
and U9073 (N_9073,N_7576,N_6562);
nor U9074 (N_9074,N_7806,N_7611);
and U9075 (N_9075,N_8465,N_8392);
and U9076 (N_9076,N_8522,N_8801);
or U9077 (N_9077,N_8269,N_7630);
or U9078 (N_9078,N_8079,N_7261);
nor U9079 (N_9079,N_6344,N_7097);
xor U9080 (N_9080,N_6288,N_7904);
or U9081 (N_9081,N_6319,N_7585);
or U9082 (N_9082,N_6969,N_8166);
or U9083 (N_9083,N_8647,N_8271);
nor U9084 (N_9084,N_7644,N_8370);
and U9085 (N_9085,N_8665,N_7553);
or U9086 (N_9086,N_6639,N_6789);
or U9087 (N_9087,N_7155,N_7479);
and U9088 (N_9088,N_6359,N_6291);
or U9089 (N_9089,N_8135,N_7781);
xnor U9090 (N_9090,N_8059,N_7632);
or U9091 (N_9091,N_7517,N_7379);
xnor U9092 (N_9092,N_7146,N_8567);
xnor U9093 (N_9093,N_8093,N_8889);
nor U9094 (N_9094,N_7143,N_6602);
nor U9095 (N_9095,N_6175,N_7824);
nor U9096 (N_9096,N_7826,N_6314);
nor U9097 (N_9097,N_7572,N_8497);
nand U9098 (N_9098,N_7628,N_7617);
and U9099 (N_9099,N_6616,N_6674);
nor U9100 (N_9100,N_7150,N_6948);
and U9101 (N_9101,N_7432,N_7649);
nand U9102 (N_9102,N_8230,N_6614);
and U9103 (N_9103,N_8192,N_8387);
or U9104 (N_9104,N_7382,N_8991);
and U9105 (N_9105,N_6382,N_8214);
nor U9106 (N_9106,N_6523,N_7926);
or U9107 (N_9107,N_8410,N_7450);
nand U9108 (N_9108,N_6923,N_7987);
xnor U9109 (N_9109,N_6992,N_6790);
nand U9110 (N_9110,N_8734,N_7142);
nor U9111 (N_9111,N_7565,N_6251);
xnor U9112 (N_9112,N_7646,N_8097);
nor U9113 (N_9113,N_6067,N_7564);
or U9114 (N_9114,N_6759,N_6463);
nand U9115 (N_9115,N_7465,N_8729);
nand U9116 (N_9116,N_8270,N_7148);
nand U9117 (N_9117,N_6375,N_6916);
and U9118 (N_9118,N_8613,N_6632);
xor U9119 (N_9119,N_8025,N_6571);
xnor U9120 (N_9120,N_7104,N_6444);
xor U9121 (N_9121,N_6466,N_7503);
xnor U9122 (N_9122,N_8541,N_8309);
nor U9123 (N_9123,N_6398,N_6401);
nand U9124 (N_9124,N_7897,N_6378);
and U9125 (N_9125,N_7242,N_8178);
nand U9126 (N_9126,N_7116,N_7531);
nand U9127 (N_9127,N_6583,N_6200);
and U9128 (N_9128,N_8056,N_6416);
xor U9129 (N_9129,N_6193,N_6439);
or U9130 (N_9130,N_8218,N_7065);
nor U9131 (N_9131,N_6732,N_8543);
nand U9132 (N_9132,N_6144,N_6945);
and U9133 (N_9133,N_7640,N_8492);
nand U9134 (N_9134,N_7795,N_7100);
or U9135 (N_9135,N_7607,N_6046);
or U9136 (N_9136,N_6260,N_6280);
nand U9137 (N_9137,N_6871,N_8251);
nand U9138 (N_9138,N_8703,N_6436);
xnor U9139 (N_9139,N_7995,N_6914);
and U9140 (N_9140,N_8907,N_7831);
nor U9141 (N_9141,N_7822,N_6471);
nor U9142 (N_9142,N_8606,N_6565);
nor U9143 (N_9143,N_7345,N_6064);
xor U9144 (N_9144,N_8708,N_8277);
nand U9145 (N_9145,N_6908,N_6970);
or U9146 (N_9146,N_6377,N_7235);
and U9147 (N_9147,N_6509,N_7859);
xor U9148 (N_9148,N_8944,N_6702);
xor U9149 (N_9149,N_8354,N_7679);
nor U9150 (N_9150,N_8141,N_6627);
and U9151 (N_9151,N_7718,N_7988);
and U9152 (N_9152,N_6569,N_8255);
nor U9153 (N_9153,N_7056,N_8584);
or U9154 (N_9154,N_7486,N_7307);
xor U9155 (N_9155,N_7184,N_7110);
xnor U9156 (N_9156,N_6592,N_8161);
nor U9157 (N_9157,N_7488,N_6972);
nand U9158 (N_9158,N_8088,N_6302);
or U9159 (N_9159,N_6407,N_8369);
nor U9160 (N_9160,N_8510,N_6054);
nand U9161 (N_9161,N_8391,N_8203);
or U9162 (N_9162,N_6717,N_6532);
xor U9163 (N_9163,N_7049,N_7291);
and U9164 (N_9164,N_8940,N_8559);
nand U9165 (N_9165,N_8331,N_7058);
or U9166 (N_9166,N_7180,N_6638);
and U9167 (N_9167,N_6005,N_7886);
xnor U9168 (N_9168,N_7297,N_7168);
and U9169 (N_9169,N_6501,N_7800);
xnor U9170 (N_9170,N_6815,N_7392);
or U9171 (N_9171,N_6932,N_8129);
nor U9172 (N_9172,N_7153,N_8471);
or U9173 (N_9173,N_8039,N_8174);
or U9174 (N_9174,N_7052,N_7317);
nor U9175 (N_9175,N_8780,N_7902);
and U9176 (N_9176,N_6897,N_6472);
or U9177 (N_9177,N_7850,N_7590);
or U9178 (N_9178,N_8546,N_7292);
nor U9179 (N_9179,N_7435,N_6423);
and U9180 (N_9180,N_7722,N_7390);
nand U9181 (N_9181,N_8657,N_6728);
or U9182 (N_9182,N_8483,N_6413);
or U9183 (N_9183,N_7549,N_6235);
and U9184 (N_9184,N_8744,N_6263);
nor U9185 (N_9185,N_6262,N_7638);
nor U9186 (N_9186,N_6603,N_8293);
or U9187 (N_9187,N_7935,N_8314);
xor U9188 (N_9188,N_6098,N_7493);
nor U9189 (N_9189,N_7388,N_8140);
nand U9190 (N_9190,N_7113,N_6691);
or U9191 (N_9191,N_7913,N_8577);
nor U9192 (N_9192,N_8153,N_8456);
xnor U9193 (N_9193,N_8259,N_8977);
xor U9194 (N_9194,N_6519,N_6796);
or U9195 (N_9195,N_8423,N_7211);
and U9196 (N_9196,N_8637,N_8407);
or U9197 (N_9197,N_7589,N_8399);
xnor U9198 (N_9198,N_7715,N_8573);
nor U9199 (N_9199,N_7789,N_8373);
and U9200 (N_9200,N_7126,N_6473);
xnor U9201 (N_9201,N_7341,N_8895);
xor U9202 (N_9202,N_6754,N_6635);
nor U9203 (N_9203,N_7543,N_7175);
nor U9204 (N_9204,N_8422,N_6447);
xor U9205 (N_9205,N_6459,N_7533);
nand U9206 (N_9206,N_6799,N_8531);
nor U9207 (N_9207,N_6095,N_7433);
xnor U9208 (N_9208,N_7298,N_7453);
nand U9209 (N_9209,N_7417,N_7490);
nand U9210 (N_9210,N_8299,N_7301);
nor U9211 (N_9211,N_6813,N_8026);
nor U9212 (N_9212,N_8283,N_8431);
and U9213 (N_9213,N_6063,N_6848);
or U9214 (N_9214,N_8086,N_7069);
nand U9215 (N_9215,N_7346,N_7352);
or U9216 (N_9216,N_6256,N_6174);
or U9217 (N_9217,N_7675,N_8941);
or U9218 (N_9218,N_7320,N_7360);
and U9219 (N_9219,N_7398,N_8561);
or U9220 (N_9220,N_6905,N_8164);
nand U9221 (N_9221,N_7840,N_7925);
and U9222 (N_9222,N_7228,N_7619);
nand U9223 (N_9223,N_6082,N_6397);
nor U9224 (N_9224,N_8724,N_7457);
and U9225 (N_9225,N_7272,N_6362);
or U9226 (N_9226,N_7459,N_6797);
nor U9227 (N_9227,N_8978,N_8473);
xor U9228 (N_9228,N_8353,N_8235);
or U9229 (N_9229,N_6807,N_6199);
nand U9230 (N_9230,N_8011,N_8324);
nand U9231 (N_9231,N_6720,N_7233);
nand U9232 (N_9232,N_7519,N_7107);
nor U9233 (N_9233,N_6240,N_6066);
nor U9234 (N_9234,N_8552,N_8842);
nand U9235 (N_9235,N_8700,N_7027);
xnor U9236 (N_9236,N_7698,N_6683);
nand U9237 (N_9237,N_8951,N_6841);
nand U9238 (N_9238,N_6880,N_8956);
and U9239 (N_9239,N_7004,N_7844);
nor U9240 (N_9240,N_7528,N_7251);
xor U9241 (N_9241,N_7594,N_7034);
nor U9242 (N_9242,N_7595,N_6103);
nand U9243 (N_9243,N_7368,N_8496);
and U9244 (N_9244,N_6218,N_7328);
and U9245 (N_9245,N_7167,N_8535);
or U9246 (N_9246,N_8232,N_6215);
and U9247 (N_9247,N_6036,N_7745);
nand U9248 (N_9248,N_6146,N_6300);
or U9249 (N_9249,N_8718,N_6304);
or U9250 (N_9250,N_8570,N_7506);
nor U9251 (N_9251,N_8511,N_6793);
nor U9252 (N_9252,N_6417,N_7917);
nand U9253 (N_9253,N_8447,N_7355);
nor U9254 (N_9254,N_8667,N_6673);
or U9255 (N_9255,N_7879,N_7029);
nor U9256 (N_9256,N_6752,N_7764);
or U9257 (N_9257,N_8200,N_6775);
or U9258 (N_9258,N_6784,N_7887);
and U9259 (N_9259,N_7248,N_6709);
nand U9260 (N_9260,N_7023,N_8954);
nand U9261 (N_9261,N_8666,N_8845);
and U9262 (N_9262,N_7447,N_8626);
and U9263 (N_9263,N_6456,N_7747);
xor U9264 (N_9264,N_6941,N_7452);
xor U9265 (N_9265,N_6724,N_8928);
nand U9266 (N_9266,N_7356,N_6002);
nor U9267 (N_9267,N_6867,N_8474);
nor U9268 (N_9268,N_6606,N_6698);
xnor U9269 (N_9269,N_6557,N_7074);
nor U9270 (N_9270,N_6402,N_8081);
nand U9271 (N_9271,N_7596,N_6521);
nor U9272 (N_9272,N_8405,N_6287);
nand U9273 (N_9273,N_6408,N_6538);
and U9274 (N_9274,N_7362,N_8120);
or U9275 (N_9275,N_7504,N_6041);
nand U9276 (N_9276,N_7405,N_7739);
xnor U9277 (N_9277,N_7889,N_7870);
nand U9278 (N_9278,N_8880,N_6190);
or U9279 (N_9279,N_8618,N_7534);
and U9280 (N_9280,N_8523,N_8946);
or U9281 (N_9281,N_8778,N_8679);
nor U9282 (N_9282,N_8776,N_8791);
or U9283 (N_9283,N_8909,N_8891);
nand U9284 (N_9284,N_6530,N_7026);
nand U9285 (N_9285,N_8544,N_8428);
or U9286 (N_9286,N_8406,N_7202);
nand U9287 (N_9287,N_7031,N_7461);
nor U9288 (N_9288,N_7636,N_6320);
xor U9289 (N_9289,N_6248,N_6761);
or U9290 (N_9290,N_8115,N_8747);
xor U9291 (N_9291,N_7309,N_8837);
or U9292 (N_9292,N_8914,N_6672);
nor U9293 (N_9293,N_7989,N_6249);
nand U9294 (N_9294,N_7230,N_8182);
or U9295 (N_9295,N_7769,N_7915);
nand U9296 (N_9296,N_8057,N_7232);
xor U9297 (N_9297,N_8284,N_8814);
nand U9298 (N_9298,N_7827,N_7633);
and U9299 (N_9299,N_6135,N_7953);
nand U9300 (N_9300,N_7970,N_7622);
and U9301 (N_9301,N_8229,N_7671);
nor U9302 (N_9302,N_6515,N_6427);
xnor U9303 (N_9303,N_6733,N_6141);
or U9304 (N_9304,N_6699,N_8409);
and U9305 (N_9305,N_6520,N_8245);
or U9306 (N_9306,N_8001,N_6684);
nand U9307 (N_9307,N_7885,N_7868);
nand U9308 (N_9308,N_6667,N_7430);
nand U9309 (N_9309,N_7526,N_8034);
and U9310 (N_9310,N_6184,N_8824);
or U9311 (N_9311,N_6040,N_6495);
nor U9312 (N_9312,N_6979,N_6332);
or U9313 (N_9313,N_8264,N_8239);
or U9314 (N_9314,N_8247,N_6335);
xnor U9315 (N_9315,N_7402,N_7273);
xnor U9316 (N_9316,N_6821,N_7896);
xor U9317 (N_9317,N_8147,N_6242);
xor U9318 (N_9318,N_7466,N_7944);
and U9319 (N_9319,N_7383,N_6605);
and U9320 (N_9320,N_8472,N_6115);
nand U9321 (N_9321,N_6480,N_7801);
xor U9322 (N_9322,N_7322,N_8160);
or U9323 (N_9323,N_8952,N_7832);
nand U9324 (N_9324,N_7738,N_6171);
or U9325 (N_9325,N_7691,N_6640);
or U9326 (N_9326,N_6008,N_6465);
nor U9327 (N_9327,N_7413,N_6133);
nand U9328 (N_9328,N_7077,N_7237);
or U9329 (N_9329,N_6221,N_6537);
nor U9330 (N_9330,N_8884,N_8122);
and U9331 (N_9331,N_8782,N_7267);
nor U9332 (N_9332,N_7608,N_8713);
and U9333 (N_9333,N_8033,N_8634);
and U9334 (N_9334,N_7128,N_6766);
nand U9335 (N_9335,N_7078,N_6442);
xor U9336 (N_9336,N_6844,N_7373);
or U9337 (N_9337,N_6354,N_8823);
nor U9338 (N_9338,N_7743,N_6678);
xnor U9339 (N_9339,N_7520,N_8248);
nand U9340 (N_9340,N_6284,N_7959);
nor U9341 (N_9341,N_6461,N_8252);
nand U9342 (N_9342,N_8549,N_6018);
nand U9343 (N_9343,N_7685,N_8900);
xnor U9344 (N_9344,N_8003,N_6971);
xor U9345 (N_9345,N_7264,N_7851);
xnor U9346 (N_9346,N_6158,N_7900);
nand U9347 (N_9347,N_8671,N_8642);
nand U9348 (N_9348,N_6675,N_7278);
and U9349 (N_9349,N_6360,N_6628);
nor U9350 (N_9350,N_8996,N_8878);
nand U9351 (N_9351,N_6293,N_6876);
nand U9352 (N_9352,N_8189,N_7583);
or U9353 (N_9353,N_7414,N_8855);
and U9354 (N_9354,N_7838,N_6346);
nor U9355 (N_9355,N_8568,N_8822);
xnor U9356 (N_9356,N_8693,N_7940);
nand U9357 (N_9357,N_7367,N_6729);
or U9358 (N_9358,N_8112,N_6504);
nor U9359 (N_9359,N_6357,N_8425);
nor U9360 (N_9360,N_7877,N_6765);
or U9361 (N_9361,N_8118,N_7363);
nor U9362 (N_9362,N_8087,N_6028);
or U9363 (N_9363,N_7510,N_6118);
or U9364 (N_9364,N_6917,N_7756);
xnor U9365 (N_9365,N_7774,N_6400);
xnor U9366 (N_9366,N_7209,N_6358);
and U9367 (N_9367,N_6774,N_7311);
and U9368 (N_9368,N_7701,N_8206);
xor U9369 (N_9369,N_6076,N_8282);
or U9370 (N_9370,N_8722,N_8799);
xor U9371 (N_9371,N_6411,N_7239);
nor U9372 (N_9372,N_6366,N_8466);
nand U9373 (N_9373,N_6038,N_7656);
xor U9374 (N_9374,N_7195,N_8432);
or U9375 (N_9375,N_7499,N_6802);
or U9376 (N_9376,N_8124,N_6918);
xnor U9377 (N_9377,N_8685,N_6409);
xnor U9378 (N_9378,N_8408,N_8785);
nand U9379 (N_9379,N_8997,N_8683);
nand U9380 (N_9380,N_6420,N_6652);
or U9381 (N_9381,N_8365,N_8254);
and U9382 (N_9382,N_7802,N_6216);
or U9383 (N_9383,N_8534,N_8680);
nor U9384 (N_9384,N_8717,N_6987);
xor U9385 (N_9385,N_6993,N_6431);
nor U9386 (N_9386,N_7937,N_7750);
nor U9387 (N_9387,N_6381,N_6283);
nand U9388 (N_9388,N_7295,N_8832);
nand U9389 (N_9389,N_6608,N_7725);
xnor U9390 (N_9390,N_7302,N_7455);
or U9391 (N_9391,N_6159,N_7793);
xnor U9392 (N_9392,N_8519,N_7090);
xnor U9393 (N_9393,N_7216,N_8876);
or U9394 (N_9394,N_7842,N_7681);
and U9395 (N_9395,N_8144,N_8751);
and U9396 (N_9396,N_6999,N_8351);
nand U9397 (N_9397,N_8737,N_6496);
nor U9398 (N_9398,N_8482,N_7263);
xor U9399 (N_9399,N_6541,N_6554);
or U9400 (N_9400,N_7210,N_7791);
nand U9401 (N_9401,N_7162,N_7330);
nand U9402 (N_9402,N_8261,N_6827);
nand U9403 (N_9403,N_6165,N_6134);
nor U9404 (N_9404,N_8225,N_6730);
or U9405 (N_9405,N_7041,N_8735);
xnor U9406 (N_9406,N_7498,N_6143);
nand U9407 (N_9407,N_8304,N_8461);
or U9408 (N_9408,N_7689,N_6142);
and U9409 (N_9409,N_6859,N_8103);
nand U9410 (N_9410,N_8014,N_6580);
and U9411 (N_9411,N_7399,N_6561);
or U9412 (N_9412,N_8187,N_6015);
and U9413 (N_9413,N_8902,N_8805);
nor U9414 (N_9414,N_8224,N_7001);
nand U9415 (N_9415,N_7872,N_8165);
nor U9416 (N_9416,N_6960,N_6888);
nand U9417 (N_9417,N_8953,N_8234);
xnor U9418 (N_9418,N_7584,N_6763);
or U9419 (N_9419,N_6747,N_8540);
nor U9420 (N_9420,N_7871,N_6758);
nand U9421 (N_9421,N_8775,N_6081);
xnor U9422 (N_9422,N_6012,N_7255);
and U9423 (N_9423,N_7515,N_6663);
and U9424 (N_9424,N_8563,N_8621);
or U9425 (N_9425,N_7821,N_6980);
and U9426 (N_9426,N_6919,N_8883);
xor U9427 (N_9427,N_6885,N_7882);
and U9428 (N_9428,N_7540,N_6210);
or U9429 (N_9429,N_8355,N_7629);
nor U9430 (N_9430,N_8760,N_6487);
nand U9431 (N_9431,N_8027,N_6433);
nand U9432 (N_9432,N_8806,N_8463);
and U9433 (N_9433,N_8451,N_7512);
nand U9434 (N_9434,N_6011,N_6889);
and U9435 (N_9435,N_7907,N_7157);
xor U9436 (N_9436,N_7257,N_7037);
nand U9437 (N_9437,N_7283,N_7567);
and U9438 (N_9438,N_6624,N_6227);
xnor U9439 (N_9439,N_8396,N_7960);
or U9440 (N_9440,N_6745,N_8602);
and U9441 (N_9441,N_7581,N_8376);
nand U9442 (N_9442,N_8925,N_8919);
nand U9443 (N_9443,N_8127,N_7350);
xor U9444 (N_9444,N_8865,N_8692);
nand U9445 (N_9445,N_6855,N_6772);
xnor U9446 (N_9446,N_8615,N_6735);
and U9447 (N_9447,N_6246,N_6901);
or U9448 (N_9448,N_8201,N_8728);
and U9449 (N_9449,N_7866,N_8128);
or U9450 (N_9450,N_8643,N_6636);
xnor U9451 (N_9451,N_7978,N_7101);
or U9452 (N_9452,N_6890,N_6595);
nor U9453 (N_9453,N_7770,N_7203);
nor U9454 (N_9454,N_7538,N_6950);
or U9455 (N_9455,N_6617,N_8356);
and U9456 (N_9456,N_8767,N_6453);
nor U9457 (N_9457,N_7843,N_6599);
and U9458 (N_9458,N_7699,N_8998);
and U9459 (N_9459,N_8636,N_6152);
nor U9460 (N_9460,N_8508,N_8071);
nor U9461 (N_9461,N_6083,N_7163);
or U9462 (N_9462,N_7196,N_7946);
nand U9463 (N_9463,N_8278,N_7758);
nand U9464 (N_9464,N_8917,N_6666);
nand U9465 (N_9465,N_8709,N_8999);
xor U9466 (N_9466,N_8125,N_8106);
xnor U9467 (N_9467,N_8196,N_6156);
or U9468 (N_9468,N_8339,N_7703);
and U9469 (N_9469,N_7613,N_8745);
nor U9470 (N_9470,N_8868,N_7550);
and U9471 (N_9471,N_6313,N_7955);
nand U9472 (N_9472,N_6978,N_8397);
and U9473 (N_9473,N_6484,N_7062);
xor U9474 (N_9474,N_6488,N_7788);
and U9475 (N_9475,N_7936,N_8558);
and U9476 (N_9476,N_8326,N_7942);
xnor U9477 (N_9477,N_8858,N_8054);
xnor U9478 (N_9478,N_6025,N_6167);
nor U9479 (N_9479,N_7274,N_6601);
nand U9480 (N_9480,N_8440,N_8485);
and U9481 (N_9481,N_6655,N_7199);
nor U9482 (N_9482,N_8484,N_6042);
nor U9483 (N_9483,N_8812,N_8241);
nor U9484 (N_9484,N_7249,N_7687);
nand U9485 (N_9485,N_8268,N_6904);
xor U9486 (N_9486,N_7305,N_8789);
xnor U9487 (N_9487,N_6422,N_8673);
or U9488 (N_9488,N_8894,N_8959);
and U9489 (N_9489,N_8886,N_6329);
nand U9490 (N_9490,N_8911,N_6713);
xor U9491 (N_9491,N_6516,N_6205);
or U9492 (N_9492,N_8749,N_8231);
xnor U9493 (N_9493,N_8179,N_6860);
xnor U9494 (N_9494,N_8191,N_8594);
xnor U9495 (N_9495,N_6070,N_8236);
nor U9496 (N_9496,N_8530,N_6089);
and U9497 (N_9497,N_7135,N_8796);
or U9498 (N_9498,N_8627,N_6840);
nor U9499 (N_9499,N_8571,N_7856);
nand U9500 (N_9500,N_6153,N_8738);
nor U9501 (N_9501,N_8754,N_7614);
xor U9502 (N_9502,N_7857,N_6468);
xnor U9503 (N_9503,N_7035,N_7880);
nand U9504 (N_9504,N_8302,N_6870);
xor U9505 (N_9505,N_6107,N_7396);
nand U9506 (N_9506,N_8569,N_8340);
and U9507 (N_9507,N_7741,N_8238);
nor U9508 (N_9508,N_8926,N_8273);
nor U9509 (N_9509,N_7442,N_8426);
nand U9510 (N_9510,N_8813,N_8133);
or U9511 (N_9511,N_6985,N_8699);
nor U9512 (N_9512,N_8242,N_6230);
xor U9513 (N_9513,N_6085,N_6787);
or U9514 (N_9514,N_6250,N_7206);
or U9515 (N_9515,N_8433,N_6726);
and U9516 (N_9516,N_6176,N_7700);
or U9517 (N_9517,N_7658,N_6446);
xnor U9518 (N_9518,N_6755,N_8444);
nand U9519 (N_9519,N_8228,N_8318);
or U9520 (N_9520,N_6285,N_8263);
or U9521 (N_9521,N_6647,N_6239);
nor U9522 (N_9522,N_8040,N_7759);
xor U9523 (N_9523,N_6117,N_7487);
nand U9524 (N_9524,N_6150,N_6891);
or U9525 (N_9525,N_7746,N_6268);
and U9526 (N_9526,N_6255,N_8194);
nand U9527 (N_9527,N_7439,N_8458);
nor U9528 (N_9528,N_8350,N_8415);
and U9529 (N_9529,N_7223,N_7749);
or U9530 (N_9530,N_7713,N_8435);
nand U9531 (N_9531,N_7475,N_7296);
or U9532 (N_9532,N_7717,N_7993);
and U9533 (N_9533,N_8870,N_8869);
and U9534 (N_9534,N_8616,N_7655);
nor U9535 (N_9535,N_8743,N_6983);
and U9536 (N_9536,N_6933,N_7431);
nor U9537 (N_9537,N_8452,N_6671);
or U9538 (N_9538,N_8964,N_8295);
nand U9539 (N_9539,N_7799,N_7468);
nor U9540 (N_9540,N_8676,N_6507);
nand U9541 (N_9541,N_8184,N_6013);
nand U9542 (N_9542,N_8430,N_8345);
or U9543 (N_9543,N_7867,N_8898);
xor U9544 (N_9544,N_8515,N_6212);
xnor U9545 (N_9545,N_7033,N_6099);
and U9546 (N_9546,N_8607,N_6493);
or U9547 (N_9547,N_6315,N_7066);
and U9548 (N_9548,N_8732,N_8547);
nand U9549 (N_9549,N_7009,N_7820);
and U9550 (N_9550,N_7916,N_7256);
xnor U9551 (N_9551,N_6651,N_8073);
nor U9552 (N_9552,N_6305,N_6370);
xor U9553 (N_9553,N_6926,N_8062);
xor U9554 (N_9554,N_7094,N_6676);
and U9555 (N_9555,N_8137,N_8267);
and U9556 (N_9556,N_6031,N_8640);
nand U9557 (N_9557,N_6892,N_8475);
or U9558 (N_9558,N_7708,N_8000);
nand U9559 (N_9559,N_7537,N_6800);
nor U9560 (N_9560,N_8779,N_7491);
nand U9561 (N_9561,N_8536,N_7964);
nand U9562 (N_9562,N_8116,N_8593);
xnor U9563 (N_9563,N_8597,N_8157);
nor U9564 (N_9564,N_6543,N_8464);
nand U9565 (N_9565,N_7304,N_7648);
and U9566 (N_9566,N_7932,N_6794);
and U9567 (N_9567,N_8938,N_8459);
nand U9568 (N_9568,N_6836,N_7425);
xor U9569 (N_9569,N_6448,N_6386);
and U9570 (N_9570,N_8036,N_7377);
nand U9571 (N_9571,N_7834,N_8149);
or U9572 (N_9572,N_8258,N_8336);
or U9573 (N_9573,N_6097,N_8291);
xor U9574 (N_9574,N_8298,N_8096);
and U9575 (N_9575,N_8686,N_6322);
xnor U9576 (N_9576,N_7400,N_6703);
and U9577 (N_9577,N_7893,N_6646);
nand U9578 (N_9578,N_6204,N_7729);
or U9579 (N_9579,N_6570,N_7043);
or U9580 (N_9580,N_8631,N_6469);
and U9581 (N_9581,N_8927,N_7914);
and U9582 (N_9582,N_7354,N_7634);
xor U9583 (N_9583,N_8768,N_8053);
nand U9584 (N_9584,N_7451,N_8342);
nor U9585 (N_9585,N_7476,N_8847);
and U9586 (N_9586,N_8006,N_7019);
and U9587 (N_9587,N_7340,N_7170);
nor U9588 (N_9588,N_6177,N_7219);
xor U9589 (N_9589,N_8018,N_6077);
or U9590 (N_9590,N_7992,N_8513);
nand U9591 (N_9591,N_6924,N_6219);
or U9592 (N_9592,N_8253,N_8795);
nand U9593 (N_9593,N_7985,N_6186);
xor U9594 (N_9594,N_7226,N_6112);
nand U9595 (N_9595,N_8294,N_7424);
or U9596 (N_9596,N_7968,N_8987);
nor U9597 (N_9597,N_6045,N_6485);
nand U9598 (N_9598,N_6128,N_7768);
xor U9599 (N_9599,N_6047,N_7365);
and U9600 (N_9600,N_6470,N_6091);
nand U9601 (N_9601,N_7876,N_6307);
or U9602 (N_9602,N_8942,N_7548);
nand U9603 (N_9603,N_7945,N_8652);
or U9604 (N_9604,N_6589,N_6414);
and U9605 (N_9605,N_8382,N_8815);
nor U9606 (N_9606,N_6207,N_6653);
xor U9607 (N_9607,N_6705,N_8539);
and U9608 (N_9608,N_7883,N_6547);
nand U9609 (N_9609,N_6549,N_7579);
or U9610 (N_9610,N_7161,N_8333);
and U9611 (N_9611,N_8797,N_7229);
and U9612 (N_9612,N_7771,N_6030);
and U9613 (N_9613,N_8246,N_8672);
xor U9614 (N_9614,N_8857,N_8596);
or U9615 (N_9615,N_6622,N_6929);
nand U9616 (N_9616,N_6566,N_6016);
or U9617 (N_9617,N_8420,N_7963);
nor U9618 (N_9618,N_8969,N_8777);
xor U9619 (N_9619,N_8761,N_7332);
or U9620 (N_9620,N_8784,N_8590);
and U9621 (N_9621,N_8610,N_8470);
xor U9622 (N_9622,N_6364,N_8119);
nand U9623 (N_9623,N_8874,N_8579);
nand U9624 (N_9624,N_6818,N_8504);
xor U9625 (N_9625,N_8835,N_8527);
nand U9626 (N_9626,N_8109,N_8706);
xor U9627 (N_9627,N_7575,N_8532);
nand U9628 (N_9628,N_6782,N_7259);
nand U9629 (N_9629,N_6670,N_7809);
and U9630 (N_9630,N_8155,N_8514);
xor U9631 (N_9631,N_7145,N_7067);
xnor U9632 (N_9632,N_6795,N_6824);
or U9633 (N_9633,N_6556,N_8963);
nand U9634 (N_9634,N_7438,N_6764);
or U9635 (N_9635,N_7327,N_8185);
and U9636 (N_9636,N_6513,N_6524);
xnor U9637 (N_9637,N_8654,N_7086);
and U9638 (N_9638,N_6271,N_7334);
xor U9639 (N_9639,N_7102,N_7212);
and U9640 (N_9640,N_6991,N_7732);
xnor U9641 (N_9641,N_6518,N_8765);
and U9642 (N_9642,N_7449,N_7007);
xnor U9643 (N_9643,N_6548,N_7265);
xor U9644 (N_9644,N_8170,N_7118);
nand U9645 (N_9645,N_8479,N_7928);
and U9646 (N_9646,N_6994,N_8462);
and U9647 (N_9647,N_8811,N_8445);
and U9648 (N_9648,N_6877,N_6591);
or U9649 (N_9649,N_6384,N_8617);
or U9650 (N_9650,N_8720,N_7401);
nor U9651 (N_9651,N_8622,N_7994);
or U9652 (N_9652,N_6792,N_8852);
or U9653 (N_9653,N_7524,N_6887);
and U9654 (N_9654,N_6321,N_7939);
xor U9655 (N_9655,N_7122,N_8844);
xnor U9656 (N_9656,N_8820,N_7986);
xnor U9657 (N_9657,N_8988,N_8390);
xnor U9658 (N_9658,N_6111,N_6644);
and U9659 (N_9659,N_6349,N_7409);
nor U9660 (N_9660,N_7483,N_6149);
or U9661 (N_9661,N_6693,N_8825);
nand U9662 (N_9662,N_6491,N_6854);
xor U9663 (N_9663,N_6274,N_8150);
nand U9664 (N_9664,N_7064,N_7574);
and U9665 (N_9665,N_8551,N_6551);
and U9666 (N_9666,N_7003,N_7395);
nand U9667 (N_9667,N_7597,N_8305);
nor U9668 (N_9668,N_7785,N_8061);
or U9669 (N_9669,N_7342,N_8279);
xnor U9670 (N_9670,N_7751,N_8658);
xor U9671 (N_9671,N_8846,N_7384);
and U9672 (N_9672,N_6367,N_8383);
nor U9673 (N_9673,N_7280,N_7063);
nor U9674 (N_9674,N_8506,N_6306);
xnor U9675 (N_9675,N_6195,N_7181);
and U9676 (N_9676,N_7542,N_6482);
and U9677 (N_9677,N_7657,N_6394);
nand U9678 (N_9678,N_7080,N_6896);
xnor U9679 (N_9679,N_7927,N_6120);
xor U9680 (N_9680,N_7763,N_6110);
nor U9681 (N_9681,N_8439,N_6679);
nor U9682 (N_9682,N_6731,N_7492);
nand U9683 (N_9683,N_8611,N_7173);
and U9684 (N_9684,N_7270,N_7709);
xor U9685 (N_9685,N_6365,N_7214);
and U9686 (N_9686,N_8696,N_6734);
nor U9687 (N_9687,N_8924,N_7641);
and U9688 (N_9688,N_8792,N_8770);
or U9689 (N_9689,N_6736,N_7300);
nand U9690 (N_9690,N_7253,N_8682);
nand U9691 (N_9691,N_6244,N_8675);
xor U9692 (N_9692,N_6805,N_6259);
xnor U9693 (N_9693,N_7720,N_7039);
or U9694 (N_9694,N_8017,N_7324);
nand U9695 (N_9695,N_6690,N_7947);
nor U9696 (N_9696,N_8028,N_8041);
xor U9697 (N_9697,N_8138,N_6390);
xor U9698 (N_9698,N_7950,N_6209);
nand U9699 (N_9699,N_8421,N_6410);
xor U9700 (N_9700,N_8562,N_6127);
nor U9701 (N_9701,N_8205,N_6475);
nor U9702 (N_9702,N_6299,N_8887);
nor U9703 (N_9703,N_8901,N_7250);
or U9704 (N_9704,N_6737,N_8154);
xnor U9705 (N_9705,N_8967,N_8572);
nor U9706 (N_9706,N_8199,N_7910);
and U9707 (N_9707,N_8807,N_8152);
xnor U9708 (N_9708,N_8598,N_7923);
nor U9709 (N_9709,N_6785,N_7507);
nand U9710 (N_9710,N_6668,N_6455);
nand U9711 (N_9711,N_6027,N_8024);
nand U9712 (N_9712,N_8468,N_6371);
nor U9713 (N_9713,N_7318,N_8378);
xor U9714 (N_9714,N_6743,N_6862);
nor U9715 (N_9715,N_6952,N_7516);
and U9716 (N_9716,N_6101,N_6940);
nand U9717 (N_9717,N_8970,N_7030);
and U9718 (N_9718,N_8639,N_7038);
xor U9719 (N_9719,N_8221,N_7938);
nor U9720 (N_9720,N_8429,N_6812);
and U9721 (N_9721,N_7200,N_6178);
or U9722 (N_9722,N_6779,N_6829);
or U9723 (N_9723,N_6817,N_6884);
nor U9724 (N_9724,N_8721,N_7141);
nor U9725 (N_9725,N_8840,N_6464);
nor U9726 (N_9726,N_6798,N_7154);
nor U9727 (N_9727,N_7082,N_6192);
nand U9728 (N_9728,N_6757,N_8574);
xor U9729 (N_9729,N_8695,N_7615);
nor U9730 (N_9730,N_7563,N_7786);
or U9731 (N_9731,N_6816,N_7544);
and U9732 (N_9732,N_8972,N_6451);
xnor U9733 (N_9733,N_8107,N_7016);
and U9734 (N_9734,N_6925,N_6681);
or U9735 (N_9735,N_7664,N_8892);
xnor U9736 (N_9736,N_6777,N_6476);
and U9737 (N_9737,N_6404,N_6695);
and U9738 (N_9738,N_6514,N_8661);
nor U9739 (N_9739,N_6863,N_6938);
or U9740 (N_9740,N_8322,N_7804);
nor U9741 (N_9741,N_7227,N_7678);
nor U9742 (N_9742,N_8808,N_6363);
nand U9743 (N_9743,N_7535,N_7149);
or U9744 (N_9744,N_8038,N_7482);
nand U9745 (N_9745,N_7158,N_6791);
and U9746 (N_9746,N_7177,N_6550);
xnor U9747 (N_9747,N_8301,N_8489);
xor U9748 (N_9748,N_8156,N_8148);
or U9749 (N_9749,N_8044,N_6522);
nor U9750 (N_9750,N_8297,N_7443);
or U9751 (N_9751,N_7418,N_8851);
nor U9752 (N_9752,N_8763,N_6206);
nor U9753 (N_9753,N_6944,N_8843);
xnor U9754 (N_9754,N_7055,N_8162);
or U9755 (N_9755,N_8084,N_8604);
or U9756 (N_9756,N_8600,N_8899);
or U9757 (N_9757,N_6688,N_6939);
xor U9758 (N_9758,N_7266,N_6727);
nor U9759 (N_9759,N_7830,N_6783);
xnor U9760 (N_9760,N_8635,N_6869);
nand U9761 (N_9761,N_7582,N_7702);
xnor U9762 (N_9762,N_6474,N_6443);
and U9763 (N_9763,N_7855,N_8888);
nor U9764 (N_9764,N_7726,N_8346);
nand U9765 (N_9765,N_8402,N_7660);
and U9766 (N_9766,N_6631,N_7784);
nor U9767 (N_9767,N_8736,N_8538);
xnor U9768 (N_9768,N_7190,N_8528);
and U9769 (N_9769,N_7869,N_6341);
xnor U9770 (N_9770,N_6194,N_7823);
nand U9771 (N_9771,N_6879,N_8077);
xor U9772 (N_9772,N_6418,N_7022);
xor U9773 (N_9773,N_8209,N_7796);
xnor U9774 (N_9774,N_8986,N_8244);
nand U9775 (N_9775,N_8599,N_8650);
xnor U9776 (N_9776,N_7555,N_7920);
nor U9777 (N_9777,N_8861,N_7521);
or U9778 (N_9778,N_7040,N_6756);
nand U9779 (N_9779,N_8051,N_6886);
and U9780 (N_9780,N_8412,N_8949);
and U9781 (N_9781,N_8980,N_7464);
and U9782 (N_9782,N_8035,N_6990);
or U9783 (N_9783,N_6718,N_8121);
or U9784 (N_9784,N_6500,N_6711);
xnor U9785 (N_9785,N_8948,N_8031);
and U9786 (N_9786,N_7081,N_8930);
nor U9787 (N_9787,N_6510,N_8662);
or U9788 (N_9788,N_8113,N_7434);
nor U9789 (N_9789,N_7472,N_7906);
and U9790 (N_9790,N_6907,N_7448);
or U9791 (N_9791,N_6163,N_7625);
and U9792 (N_9792,N_6539,N_7805);
xnor U9793 (N_9793,N_7513,N_8691);
nor U9794 (N_9794,N_8380,N_6751);
nor U9795 (N_9795,N_7606,N_8875);
and U9796 (N_9796,N_6022,N_6913);
nand U9797 (N_9797,N_8168,N_8411);
nand U9798 (N_9798,N_6582,N_8507);
xor U9799 (N_9799,N_7683,N_7343);
xor U9800 (N_9800,N_6324,N_7221);
nand U9801 (N_9801,N_6290,N_7112);
or U9802 (N_9802,N_8005,N_6961);
nor U9803 (N_9803,N_6895,N_7716);
nor U9804 (N_9804,N_7337,N_6497);
xnor U9805 (N_9805,N_8860,N_7114);
xnor U9806 (N_9806,N_8771,N_6630);
or U9807 (N_9807,N_7299,N_8962);
and U9808 (N_9808,N_6694,N_7497);
and U9809 (N_9809,N_8730,N_8099);
or U9810 (N_9810,N_6273,N_8576);
nor U9811 (N_9811,N_6842,N_6035);
or U9812 (N_9812,N_7909,N_8764);
xor U9813 (N_9813,N_8067,N_8856);
or U9814 (N_9814,N_7471,N_8816);
nor U9815 (N_9815,N_6308,N_6102);
or U9816 (N_9816,N_6093,N_8467);
xnor U9817 (N_9817,N_7653,N_8794);
nor U9818 (N_9818,N_8498,N_7593);
or U9819 (N_9819,N_8366,N_6575);
nand U9820 (N_9820,N_6725,N_7983);
and U9821 (N_9821,N_7262,N_6723);
nand U9822 (N_9822,N_8029,N_6406);
or U9823 (N_9823,N_7197,N_7980);
xor U9824 (N_9824,N_7712,N_7735);
or U9825 (N_9825,N_7972,N_7560);
nand U9826 (N_9826,N_6680,N_8066);
and U9827 (N_9827,N_6881,N_7165);
nand U9828 (N_9828,N_6336,N_8275);
nand U9829 (N_9829,N_8015,N_6339);
or U9830 (N_9830,N_6157,N_6424);
nand U9831 (N_9831,N_6257,N_8774);
nand U9832 (N_9832,N_7024,N_8296);
nand U9833 (N_9833,N_7287,N_6056);
and U9834 (N_9834,N_7509,N_8180);
nand U9835 (N_9835,N_6625,N_6612);
xnor U9836 (N_9836,N_6770,N_6656);
and U9837 (N_9837,N_7775,N_6552);
or U9838 (N_9838,N_7426,N_7495);
nor U9839 (N_9839,N_7446,N_6626);
nand U9840 (N_9840,N_6191,N_7677);
and U9841 (N_9841,N_6545,N_6922);
or U9842 (N_9842,N_6838,N_7941);
xor U9843 (N_9843,N_8896,N_7238);
nand U9844 (N_9844,N_7598,N_6769);
or U9845 (N_9845,N_7545,N_8553);
and U9846 (N_9846,N_7949,N_7873);
nor U9847 (N_9847,N_8443,N_8100);
nand U9848 (N_9848,N_6949,N_6579);
nor U9849 (N_9849,N_7178,N_8525);
nand U9850 (N_9850,N_8704,N_6108);
xnor U9851 (N_9851,N_8516,N_8007);
nand U9852 (N_9852,N_6428,N_8937);
nor U9853 (N_9853,N_6309,N_7224);
or U9854 (N_9854,N_7234,N_8833);
nor U9855 (N_9855,N_8055,N_7990);
and U9856 (N_9856,N_7147,N_7602);
and U9857 (N_9857,N_7603,N_7111);
and U9858 (N_9858,N_6995,N_6071);
or U9859 (N_9859,N_6185,N_6387);
xor U9860 (N_9860,N_8933,N_6396);
nand U9861 (N_9861,N_6883,N_6074);
or U9862 (N_9862,N_6984,N_6170);
nand U9863 (N_9863,N_8453,N_8798);
or U9864 (N_9864,N_6075,N_8564);
nand U9865 (N_9865,N_6915,N_7132);
xor U9866 (N_9866,N_7737,N_7591);
and U9867 (N_9867,N_7361,N_7684);
xnor U9868 (N_9868,N_8804,N_7246);
and U9869 (N_9869,N_7166,N_8352);
nor U9870 (N_9870,N_8188,N_7370);
nor U9871 (N_9871,N_7119,N_6689);
and U9872 (N_9872,N_6963,N_7294);
nor U9873 (N_9873,N_7693,N_6203);
or U9874 (N_9874,N_8176,N_8939);
xnor U9875 (N_9875,N_7096,N_7293);
or U9876 (N_9876,N_7271,N_6437);
and U9877 (N_9877,N_6168,N_7954);
nor U9878 (N_9878,N_8134,N_7623);
nor U9879 (N_9879,N_6584,N_7961);
and U9880 (N_9880,N_7643,N_7586);
nand U9881 (N_9881,N_6369,N_6634);
and U9882 (N_9882,N_6826,N_8393);
nor U9883 (N_9883,N_8920,N_6900);
xor U9884 (N_9884,N_8379,N_8315);
or U9885 (N_9885,N_7480,N_7569);
and U9886 (N_9886,N_6182,N_6910);
nand U9887 (N_9887,N_8368,N_7474);
xnor U9888 (N_9888,N_7672,N_7312);
xor U9889 (N_9889,N_8829,N_8882);
nor U9890 (N_9890,N_8372,N_6162);
nand U9891 (N_9891,N_7998,N_7635);
nor U9892 (N_9892,N_7757,N_8110);
or U9893 (N_9893,N_7436,N_8853);
xor U9894 (N_9894,N_6615,N_8500);
or U9895 (N_9895,N_7284,N_6278);
nand U9896 (N_9896,N_6645,N_7728);
nor U9897 (N_9897,N_6325,N_6921);
xnor U9898 (N_9898,N_8971,N_7588);
or U9899 (N_9899,N_7473,N_8177);
and U9900 (N_9900,N_7839,N_6289);
xnor U9901 (N_9901,N_8694,N_7848);
nand U9902 (N_9902,N_6389,N_6405);
nor U9903 (N_9903,N_8233,N_8800);
nand U9904 (N_9904,N_7220,N_7639);
nor U9905 (N_9905,N_8879,N_7231);
or U9906 (N_9906,N_7665,N_7667);
nand U9907 (N_9907,N_7205,N_7815);
or U9908 (N_9908,N_8418,N_6226);
or U9909 (N_9909,N_6238,N_6555);
nand U9910 (N_9910,N_8381,N_7002);
xnor U9911 (N_9911,N_7704,N_7798);
nor U9912 (N_9912,N_8332,N_6048);
nor U9913 (N_9913,N_8688,N_7810);
or U9914 (N_9914,N_6505,N_6234);
nor U9915 (N_9915,N_7172,N_7884);
and U9916 (N_9916,N_7411,N_8603);
and U9917 (N_9917,N_6658,N_6032);
nor U9918 (N_9918,N_6220,N_7527);
or U9919 (N_9919,N_8614,N_8841);
and U9920 (N_9920,N_8687,N_8943);
nand U9921 (N_9921,N_8401,N_8524);
nor U9922 (N_9922,N_7776,N_8950);
or U9923 (N_9923,N_7243,N_8375);
xor U9924 (N_9924,N_8306,N_6222);
or U9925 (N_9925,N_6122,N_7140);
nor U9926 (N_9926,N_6148,N_6498);
and U9927 (N_9927,N_8400,N_7463);
or U9928 (N_9928,N_7841,N_7500);
xor U9929 (N_9929,N_8222,N_6739);
nor U9930 (N_9930,N_6738,N_8104);
nor U9931 (N_9931,N_6865,N_6340);
nor U9932 (N_9932,N_6853,N_7612);
nand U9933 (N_9933,N_7616,N_6017);
nor U9934 (N_9934,N_7092,N_6264);
or U9935 (N_9935,N_8126,N_7794);
or U9936 (N_9936,N_7015,N_6281);
nand U9937 (N_9937,N_8132,N_6350);
or U9938 (N_9938,N_8819,N_6090);
nor U9939 (N_9939,N_8348,N_8788);
nor U9940 (N_9940,N_8300,N_7973);
xnor U9941 (N_9941,N_8748,N_8554);
nand U9942 (N_9942,N_6121,N_8276);
or U9943 (N_9943,N_7957,N_8605);
or U9944 (N_9944,N_7012,N_6964);
nor U9945 (N_9945,N_7348,N_6432);
xnor U9946 (N_9946,N_6003,N_7744);
xnor U9947 (N_9947,N_7780,N_8756);
nor U9948 (N_9948,N_7692,N_8111);
or U9949 (N_9949,N_7668,N_6380);
nand U9950 (N_9950,N_7133,N_7098);
and U9951 (N_9951,N_6965,N_7247);
and U9952 (N_9952,N_7021,N_8520);
nor U9953 (N_9953,N_8337,N_6426);
and U9954 (N_9954,N_6708,N_8414);
or U9955 (N_9955,N_6132,N_7621);
and U9956 (N_9956,N_6311,N_8320);
nand U9957 (N_9957,N_6835,N_8338);
and U9958 (N_9958,N_7714,N_6781);
and U9959 (N_9959,N_7637,N_7000);
nand U9960 (N_9960,N_6124,N_8413);
xor U9961 (N_9961,N_8915,N_8936);
nor U9962 (N_9962,N_7710,N_7899);
or U9963 (N_9963,N_6856,N_7919);
nand U9964 (N_9964,N_6275,N_7321);
or U9965 (N_9965,N_8992,N_6292);
nor U9966 (N_9966,N_6169,N_7347);
and U9967 (N_9967,N_6109,N_8091);
nand U9968 (N_9968,N_8495,N_8834);
or U9969 (N_9969,N_8198,N_6338);
nor U9970 (N_9970,N_8714,N_6619);
nand U9971 (N_9971,N_7849,N_6164);
and U9972 (N_9972,N_7127,N_6189);
nand U9973 (N_9973,N_8043,N_7036);
nor U9974 (N_9974,N_7428,N_8102);
and U9975 (N_9975,N_7460,N_8958);
or U9976 (N_9976,N_6479,N_8499);
nor U9977 (N_9977,N_6581,N_7532);
xnor U9978 (N_9978,N_7921,N_7557);
and U9979 (N_9979,N_7164,N_8481);
nor U9980 (N_9980,N_7891,N_6512);
xor U9981 (N_9981,N_7967,N_7289);
and U9982 (N_9982,N_7673,N_7393);
xor U9983 (N_9983,N_6270,N_8512);
xnor U9984 (N_9984,N_8710,N_6223);
and U9985 (N_9985,N_8973,N_8114);
nor U9986 (N_9986,N_6014,N_7817);
or U9987 (N_9987,N_8862,N_6819);
and U9988 (N_9988,N_8074,N_8906);
xnor U9989 (N_9989,N_7319,N_8580);
nand U9990 (N_9990,N_6294,N_8173);
nor U9991 (N_9991,N_7878,N_6832);
nand U9992 (N_9992,N_8904,N_8923);
nor U9993 (N_9993,N_8910,N_6481);
nor U9994 (N_9994,N_7008,N_6225);
xor U9995 (N_9995,N_8509,N_6055);
or U9996 (N_9996,N_7138,N_6140);
nor U9997 (N_9997,N_7072,N_8219);
nand U9998 (N_9998,N_7682,N_7601);
nand U9999 (N_9999,N_8828,N_6179);
xnor U10000 (N_10000,N_7136,N_6379);
nand U10001 (N_10001,N_8701,N_7706);
xnor U10002 (N_10002,N_7807,N_7670);
nand U10003 (N_10003,N_8947,N_6654);
or U10004 (N_10004,N_6996,N_8139);
nor U10005 (N_10005,N_6621,N_6837);
and U10006 (N_10006,N_6419,N_8037);
and U10007 (N_10007,N_7285,N_8817);
xor U10008 (N_10008,N_7427,N_7364);
or U10009 (N_10009,N_6506,N_7217);
or U10010 (N_10010,N_6740,N_8668);
and U10011 (N_10011,N_7326,N_8908);
nand U10012 (N_10012,N_8490,N_7429);
or U10013 (N_10013,N_7349,N_7193);
xnor U10014 (N_10014,N_8982,N_7846);
or U10015 (N_10015,N_7279,N_7816);
or U10016 (N_10016,N_6657,N_8364);
and U10017 (N_10017,N_7088,N_6536);
or U10018 (N_10018,N_8961,N_8934);
and U10019 (N_10019,N_6574,N_8427);
nor U10020 (N_10020,N_6642,N_8070);
xnor U10021 (N_10021,N_7901,N_7982);
and U10022 (N_10022,N_7505,N_6353);
nand U10023 (N_10023,N_6198,N_8357);
or U10024 (N_10024,N_7371,N_8893);
nor U10025 (N_10025,N_7587,N_8588);
and U10026 (N_10026,N_6833,N_8646);
nand U10027 (N_10027,N_7423,N_6600);
or U10028 (N_10028,N_7686,N_6096);
or U10029 (N_10029,N_7014,N_8257);
or U10030 (N_10030,N_7093,N_7976);
and U10031 (N_10031,N_8012,N_6068);
or U10032 (N_10032,N_7911,N_7852);
nand U10033 (N_10033,N_8945,N_6272);
xor U10034 (N_10034,N_6741,N_6388);
nor U10035 (N_10035,N_6661,N_8719);
xor U10036 (N_10036,N_8592,N_8131);
xnor U10037 (N_10037,N_8867,N_7339);
nor U10038 (N_10038,N_8787,N_7477);
or U10039 (N_10039,N_7525,N_7198);
or U10040 (N_10040,N_6342,N_8935);
nand U10041 (N_10041,N_6197,N_7828);
nand U10042 (N_10042,N_6576,N_7194);
nand U10043 (N_10043,N_6874,N_7696);
or U10044 (N_10044,N_6104,N_7898);
nor U10045 (N_10045,N_7456,N_6586);
or U10046 (N_10046,N_6803,N_6649);
and U10047 (N_10047,N_6247,N_6607);
and U10048 (N_10048,N_6061,N_7862);
and U10049 (N_10049,N_6981,N_6228);
nand U10050 (N_10050,N_6943,N_7558);
nand U10051 (N_10051,N_8048,N_6231);
xnor U10052 (N_10052,N_7308,N_6049);
or U10053 (N_10053,N_8394,N_7536);
xor U10054 (N_10054,N_6558,N_8526);
nor U10055 (N_10055,N_7627,N_8557);
nand U10056 (N_10056,N_8595,N_7778);
and U10057 (N_10057,N_8994,N_8781);
or U10058 (N_10058,N_6778,N_6508);
and U10059 (N_10059,N_6125,N_8064);
xor U10060 (N_10060,N_6810,N_8873);
xnor U10061 (N_10061,N_7811,N_7011);
nor U10062 (N_10062,N_7730,N_7592);
or U10063 (N_10063,N_6503,N_8361);
nor U10064 (N_10064,N_6253,N_8759);
nand U10065 (N_10065,N_8663,N_8955);
and U10066 (N_10066,N_6771,N_7252);
nand U10067 (N_10067,N_6650,N_6788);
or U10068 (N_10068,N_7288,N_7169);
and U10069 (N_10069,N_8872,N_7462);
and U10070 (N_10070,N_8790,N_6878);
or U10071 (N_10071,N_7381,N_7631);
and U10072 (N_10072,N_8566,N_7508);
nand U10073 (N_10073,N_6563,N_7924);
or U10074 (N_10074,N_6078,N_6801);
nand U10075 (N_10075,N_7912,N_6452);
or U10076 (N_10076,N_6334,N_7046);
or U10077 (N_10077,N_7131,N_8183);
xor U10078 (N_10078,N_8172,N_6858);
xnor U10079 (N_10079,N_7060,N_6544);
and U10080 (N_10080,N_6843,N_6587);
nor U10081 (N_10081,N_6147,N_6613);
nand U10082 (N_10082,N_7782,N_8537);
nand U10083 (N_10083,N_6834,N_7573);
xnor U10084 (N_10084,N_7144,N_6986);
or U10085 (N_10085,N_6590,N_7523);
xor U10086 (N_10086,N_6052,N_6392);
and U10087 (N_10087,N_6585,N_8989);
xnor U10088 (N_10088,N_8521,N_8698);
nor U10089 (N_10089,N_7892,N_8065);
or U10090 (N_10090,N_6020,N_6845);
xor U10091 (N_10091,N_8285,N_8163);
xor U10092 (N_10092,N_8786,N_7766);
and U10093 (N_10093,N_6026,N_7895);
or U10094 (N_10094,N_8913,N_6955);
nand U10095 (N_10095,N_8159,N_6831);
or U10096 (N_10096,N_8123,N_8493);
or U10097 (N_10097,N_7416,N_8976);
and U10098 (N_10098,N_7754,N_8529);
or U10099 (N_10099,N_8494,N_8985);
xor U10100 (N_10100,N_7724,N_7378);
or U10101 (N_10101,N_6857,N_8249);
nor U10102 (N_10102,N_6151,N_6806);
nand U10103 (N_10103,N_7864,N_6004);
and U10104 (N_10104,N_8151,N_8308);
and U10105 (N_10105,N_7568,N_8307);
xnor U10106 (N_10106,N_6415,N_8210);
and U10107 (N_10107,N_8649,N_6664);
and U10108 (N_10108,N_6356,N_8343);
nand U10109 (N_10109,N_7357,N_6295);
and U10110 (N_10110,N_8117,N_8312);
xnor U10111 (N_10111,N_7422,N_8349);
nor U10112 (N_10112,N_6105,N_6997);
xor U10113 (N_10113,N_8289,N_8727);
or U10114 (N_10114,N_6438,N_7314);
and U10115 (N_10115,N_7661,N_6345);
or U10116 (N_10116,N_6188,N_8359);
nor U10117 (N_10117,N_6137,N_6361);
xor U10118 (N_10118,N_7282,N_8742);
nand U10119 (N_10119,N_8533,N_7333);
xor U10120 (N_10120,N_6942,N_8705);
or U10121 (N_10121,N_6069,N_6973);
or U10122 (N_10122,N_6202,N_6155);
xor U10123 (N_10123,N_7818,N_6893);
or U10124 (N_10124,N_6609,N_8341);
nand U10125 (N_10125,N_8921,N_7374);
nor U10126 (N_10126,N_6906,N_7191);
nand U10127 (N_10127,N_6043,N_7501);
nand U10128 (N_10128,N_6126,N_8905);
nor U10129 (N_10129,N_7387,N_7335);
nand U10130 (N_10130,N_6648,N_8330);
or U10131 (N_10131,N_8766,N_6967);
nor U10132 (N_10132,N_8503,N_7160);
nand U10133 (N_10133,N_6511,N_7005);
and U10134 (N_10134,N_8450,N_8080);
or U10135 (N_10135,N_6059,N_6395);
and U10136 (N_10136,N_7079,N_6374);
xor U10137 (N_10137,N_6347,N_8922);
xnor U10138 (N_10138,N_8290,N_8619);
xor U10139 (N_10139,N_7918,N_6687);
xor U10140 (N_10140,N_6749,N_8292);
or U10141 (N_10141,N_7556,N_6618);
and U10142 (N_10142,N_6903,N_6611);
or U10143 (N_10143,N_7105,N_7642);
nand U10144 (N_10144,N_6483,N_6337);
nor U10145 (N_10145,N_7109,N_7787);
nand U10146 (N_10146,N_7688,N_7707);
or U10147 (N_10147,N_8327,N_7013);
nor U10148 (N_10148,N_8681,N_6567);
or U10149 (N_10149,N_6578,N_8556);
and U10150 (N_10150,N_6677,N_6773);
or U10151 (N_10151,N_8362,N_8092);
nor U10152 (N_10152,N_7075,N_6931);
or U10153 (N_10153,N_8638,N_8655);
nand U10154 (N_10154,N_7761,N_6282);
nor U10155 (N_10155,N_7984,N_6828);
or U10156 (N_10156,N_8213,N_7125);
and U10157 (N_10157,N_6007,N_6266);
or U10158 (N_10158,N_8993,N_8010);
nor U10159 (N_10159,N_7546,N_7999);
nor U10160 (N_10160,N_7723,N_8587);
or U10161 (N_10161,N_6450,N_7790);
and U10162 (N_10162,N_8866,N_8347);
and U10163 (N_10163,N_7244,N_8130);
nand U10164 (N_10164,N_8193,N_8095);
xor U10165 (N_10165,N_7991,N_6458);
xnor U10166 (N_10166,N_7626,N_6119);
xnor U10167 (N_10167,N_7467,N_7511);
and U10168 (N_10168,N_8212,N_8750);
xnor U10169 (N_10169,N_6021,N_7329);
and U10170 (N_10170,N_7174,N_7344);
nand U10171 (N_10171,N_7171,N_6286);
nor U10172 (N_10172,N_8974,N_8223);
and U10173 (N_10173,N_8319,N_7752);
xor U10174 (N_10174,N_7156,N_6692);
nand U10175 (N_10175,N_7930,N_6462);
nand U10176 (N_10176,N_6492,N_8437);
nor U10177 (N_10177,N_7530,N_6211);
and U10178 (N_10178,N_6968,N_8586);
xnor U10179 (N_10179,N_6808,N_6001);
nand U10180 (N_10180,N_8449,N_7819);
xnor U10181 (N_10181,N_7087,N_7772);
or U10182 (N_10182,N_6123,N_7176);
nor U10183 (N_10183,N_7694,N_6160);
or U10184 (N_10184,N_6912,N_6559);
xnor U10185 (N_10185,N_6660,N_6882);
nor U10186 (N_10186,N_6762,N_7048);
nor U10187 (N_10187,N_6172,N_7089);
or U10188 (N_10188,N_6065,N_7676);
and U10189 (N_10189,N_6208,N_8589);
and U10190 (N_10190,N_6310,N_6909);
and U10191 (N_10191,N_8478,N_8046);
xnor U10192 (N_10192,N_8220,N_7554);
xor U10193 (N_10193,N_7420,N_6136);
nand U10194 (N_10194,N_8864,N_7571);
or U10195 (N_10195,N_7808,N_6750);
nand U10196 (N_10196,N_6830,N_8002);
xnor U10197 (N_10197,N_6368,N_8442);
or U10198 (N_10198,N_7006,N_6988);
or U10199 (N_10199,N_8575,N_6697);
or U10200 (N_10200,N_6977,N_8502);
nor U10201 (N_10201,N_8424,N_6825);
and U10202 (N_10202,N_8344,N_8190);
nand U10203 (N_10203,N_6145,N_6449);
xor U10204 (N_10204,N_7669,N_7032);
nand U10205 (N_10205,N_7208,N_7847);
xnor U10206 (N_10206,N_6954,N_8262);
and U10207 (N_10207,N_7740,N_6265);
nand U10208 (N_10208,N_6872,N_6927);
or U10209 (N_10209,N_8105,N_8830);
and U10210 (N_10210,N_6138,N_8146);
nand U10211 (N_10211,N_8089,N_8550);
nand U10212 (N_10212,N_7290,N_8871);
xnor U10213 (N_10213,N_7061,N_8020);
or U10214 (N_10214,N_8323,N_6316);
nor U10215 (N_10215,N_7489,N_8984);
nand U10216 (N_10216,N_7018,N_8217);
and U10217 (N_10217,N_7965,N_6669);
xor U10218 (N_10218,N_6116,N_6489);
nor U10219 (N_10219,N_6201,N_8310);
and U10220 (N_10220,N_6236,N_6224);
xor U10221 (N_10221,N_8849,N_7068);
and U10222 (N_10222,N_8388,N_8702);
xor U10223 (N_10223,N_8108,N_8623);
xor U10224 (N_10224,N_8256,N_7108);
nor U10225 (N_10225,N_6060,N_8505);
nor U10226 (N_10226,N_8826,N_6434);
nor U10227 (N_10227,N_6214,N_7599);
and U10228 (N_10228,N_8175,N_8358);
nand U10229 (N_10229,N_7159,N_8501);
or U10230 (N_10230,N_7137,N_8545);
or U10231 (N_10231,N_6531,N_7813);
and U10232 (N_10232,N_8455,N_6527);
nor U10233 (N_10233,N_7375,N_6560);
and U10234 (N_10234,N_6704,N_7073);
or U10235 (N_10235,N_8049,N_8335);
xor U10236 (N_10236,N_7189,N_7733);
or U10237 (N_10237,N_8758,N_7222);
or U10238 (N_10238,N_6269,N_8403);
nor U10239 (N_10239,N_6333,N_6084);
nand U10240 (N_10240,N_7561,N_8810);
or U10241 (N_10241,N_6460,N_6385);
and U10242 (N_10242,N_6087,N_7099);
nand U10243 (N_10243,N_7050,N_8030);
xor U10244 (N_10244,N_8803,N_8601);
and U10245 (N_10245,N_7366,N_6355);
and U10246 (N_10246,N_6391,N_6243);
or U10247 (N_10247,N_7721,N_7609);
and U10248 (N_10248,N_8434,N_6682);
xnor U10249 (N_10249,N_7268,N_6057);
xor U10250 (N_10250,N_8047,N_6352);
or U10251 (N_10251,N_6989,N_7797);
and U10252 (N_10252,N_6553,N_6526);
or U10253 (N_10253,N_8645,N_7139);
or U10254 (N_10254,N_8983,N_7380);
and U10255 (N_10255,N_8517,N_6328);
nand U10256 (N_10256,N_6445,N_7042);
xnor U10257 (N_10257,N_8316,N_8746);
xnor U10258 (N_10258,N_6540,N_6348);
nor U10259 (N_10259,N_6598,N_6839);
or U10260 (N_10260,N_6529,N_8325);
xor U10261 (N_10261,N_7213,N_6588);
xnor U10262 (N_10262,N_6959,N_7245);
or U10263 (N_10263,N_6196,N_6814);
nor U10264 (N_10264,N_6051,N_8633);
nor U10265 (N_10265,N_7792,N_6528);
or U10266 (N_10266,N_7719,N_6403);
nor U10267 (N_10267,N_6962,N_6261);
xor U10268 (N_10268,N_7974,N_8329);
and U10269 (N_10269,N_6846,N_6716);
or U10270 (N_10270,N_7045,N_6478);
nor U10271 (N_10271,N_8542,N_6953);
and U10272 (N_10272,N_7996,N_7762);
nor U10273 (N_10273,N_7890,N_7277);
and U10274 (N_10274,N_6372,N_8881);
nand U10275 (N_10275,N_6494,N_8733);
and U10276 (N_10276,N_6722,N_7415);
nor U10277 (N_10277,N_8266,N_6454);
xor U10278 (N_10278,N_7773,N_7539);
nand U10279 (N_10279,N_8226,N_6976);
and U10280 (N_10280,N_6706,N_6044);
nand U10281 (N_10281,N_7059,N_7650);
nand U10282 (N_10282,N_8145,N_7618);
xor U10283 (N_10283,N_6982,N_8186);
nor U10284 (N_10284,N_7406,N_6232);
nor U10285 (N_10285,N_8260,N_8334);
or U10286 (N_10286,N_8416,N_6318);
nand U10287 (N_10287,N_7731,N_6753);
or U10288 (N_10288,N_7372,N_6517);
or U10289 (N_10289,N_8313,N_7394);
xnor U10290 (N_10290,N_8755,N_6245);
or U10291 (N_10291,N_8286,N_8142);
and U10292 (N_10292,N_7454,N_7440);
nor U10293 (N_10293,N_7389,N_6094);
and U10294 (N_10294,N_8360,N_7386);
xor U10295 (N_10295,N_7152,N_7652);
nor U10296 (N_10296,N_8659,N_7829);
nand U10297 (N_10297,N_8918,N_8739);
nor U10298 (N_10298,N_8762,N_8204);
and U10299 (N_10299,N_8058,N_8583);
or U10300 (N_10300,N_7651,N_6714);
and U10301 (N_10301,N_8098,N_7958);
or U10302 (N_10302,N_8581,N_7552);
or U10303 (N_10303,N_7047,N_6298);
xor U10304 (N_10304,N_6312,N_6181);
and U10305 (N_10305,N_8648,N_8831);
nand U10306 (N_10306,N_8063,N_8052);
nor U10307 (N_10307,N_8966,N_7338);
nand U10308 (N_10308,N_6742,N_7421);
and U10309 (N_10309,N_6086,N_8731);
or U10310 (N_10310,N_8250,N_8890);
xor U10311 (N_10311,N_7541,N_8678);
and U10312 (N_10312,N_7484,N_6767);
xnor U10313 (N_10313,N_7734,N_8960);
nand U10314 (N_10314,N_8630,N_6130);
or U10315 (N_10315,N_6577,N_8136);
xor U10316 (N_10316,N_6934,N_7481);
or U10317 (N_10317,N_6760,N_8859);
xnor U10318 (N_10318,N_8083,N_8398);
or U10319 (N_10319,N_7905,N_8838);
nor U10320 (N_10320,N_7218,N_8715);
or U10321 (N_10321,N_7115,N_7860);
xor U10322 (N_10322,N_7779,N_6572);
xnor U10323 (N_10323,N_8560,N_7853);
nor U10324 (N_10324,N_7369,N_6019);
nand U10325 (N_10325,N_7076,N_8009);
and U10326 (N_10326,N_8281,N_6533);
or U10327 (N_10327,N_7767,N_8632);
and U10328 (N_10328,N_6873,N_6849);
or U10329 (N_10329,N_7085,N_7874);
nand U10330 (N_10330,N_8912,N_7566);
nand U10331 (N_10331,N_7183,N_8669);
nand U10332 (N_10332,N_8477,N_7680);
nand U10333 (N_10333,N_6662,N_6564);
and U10334 (N_10334,N_7103,N_8207);
nand U10335 (N_10335,N_8480,N_6399);
nand U10336 (N_10336,N_6039,N_7240);
xor U10337 (N_10337,N_7760,N_8697);
xor U10338 (N_10338,N_6441,N_8076);
and U10339 (N_10339,N_6106,N_6430);
nand U10340 (N_10340,N_8404,N_7494);
or U10341 (N_10341,N_8644,N_6490);
nor U10342 (N_10342,N_8821,N_6161);
or U10343 (N_10343,N_8202,N_8143);
nor U10344 (N_10344,N_6139,N_7260);
xor U10345 (N_10345,N_7863,N_6383);
xor U10346 (N_10346,N_6597,N_7044);
and U10347 (N_10347,N_7316,N_6998);
or U10348 (N_10348,N_7966,N_6951);
nand U10349 (N_10349,N_6701,N_7888);
xnor U10350 (N_10350,N_6710,N_7276);
or U10351 (N_10351,N_6412,N_7865);
nand U10352 (N_10352,N_6712,N_7803);
or U10353 (N_10353,N_7188,N_7777);
nand U10354 (N_10354,N_8641,N_8608);
nand U10355 (N_10355,N_6920,N_8280);
xnor U10356 (N_10356,N_7814,N_8167);
nand U10357 (N_10357,N_6252,N_8707);
nand U10358 (N_10358,N_8216,N_6958);
nand U10359 (N_10359,N_6440,N_6429);
nor U10360 (N_10360,N_7854,N_8078);
or U10361 (N_10361,N_7397,N_8469);
nand U10362 (N_10362,N_7408,N_6604);
and U10363 (N_10363,N_8438,N_6875);
nand U10364 (N_10364,N_8585,N_8460);
nand U10365 (N_10365,N_6780,N_7485);
or U10366 (N_10366,N_7323,N_6072);
and U10367 (N_10367,N_8476,N_7025);
nand U10368 (N_10368,N_8854,N_7151);
xnor U10369 (N_10369,N_8072,N_7281);
nand U10370 (N_10370,N_8897,N_7020);
nor U10371 (N_10371,N_8690,N_8101);
nand U10372 (N_10372,N_8624,N_6277);
nor U10373 (N_10373,N_8386,N_7922);
xor U10374 (N_10374,N_8419,N_6079);
nor U10375 (N_10375,N_7186,N_8620);
nand U10376 (N_10376,N_7674,N_8848);
or U10377 (N_10377,N_6894,N_7313);
nor U10378 (N_10378,N_7315,N_8725);
and U10379 (N_10379,N_8240,N_7663);
nor U10380 (N_10380,N_8265,N_6899);
and U10381 (N_10381,N_8023,N_6659);
nand U10382 (N_10382,N_8656,N_6323);
or U10383 (N_10383,N_7908,N_8753);
and U10384 (N_10384,N_6330,N_7204);
and U10385 (N_10385,N_7407,N_8488);
and U10386 (N_10386,N_6486,N_7083);
and U10387 (N_10387,N_7765,N_6296);
nand U10388 (N_10388,N_7934,N_6351);
xor U10389 (N_10389,N_8417,N_8965);
and U10390 (N_10390,N_6034,N_8158);
nand U10391 (N_10391,N_7410,N_7201);
nand U10392 (N_10392,N_8555,N_6776);
xor U10393 (N_10393,N_8171,N_6596);
nand U10394 (N_10394,N_8726,N_6421);
nand U10395 (N_10395,N_8723,N_8021);
or U10396 (N_10396,N_8068,N_7659);
nor U10397 (N_10397,N_7053,N_7502);
xnor U10398 (N_10398,N_8042,N_7580);
and U10399 (N_10399,N_7010,N_6852);
nand U10400 (N_10400,N_7929,N_6326);
xnor U10401 (N_10401,N_6936,N_8651);
and U10402 (N_10402,N_8317,N_6546);
or U10403 (N_10403,N_6129,N_8711);
nand U10404 (N_10404,N_6058,N_7736);
xor U10405 (N_10405,N_8628,N_7185);
nand U10406 (N_10406,N_7977,N_8757);
xnor U10407 (N_10407,N_7120,N_6700);
or U10408 (N_10408,N_6786,N_8446);
nand U10409 (N_10409,N_6966,N_7391);
nand U10410 (N_10410,N_8548,N_6301);
or U10411 (N_10411,N_7605,N_6935);
and U10412 (N_10412,N_6525,N_6956);
xnor U10413 (N_10413,N_6542,N_8995);
nand U10414 (N_10414,N_7705,N_7458);
and U10415 (N_10415,N_8827,N_7578);
nor U10416 (N_10416,N_6023,N_8932);
xor U10417 (N_10417,N_7353,N_7727);
nor U10418 (N_10418,N_8565,N_7610);
nor U10419 (N_10419,N_8772,N_7861);
and U10420 (N_10420,N_7858,N_7948);
nand U10421 (N_10421,N_8818,N_8436);
xor U10422 (N_10422,N_7071,N_7645);
xor U10423 (N_10423,N_7179,N_6113);
nor U10424 (N_10424,N_6276,N_8169);
nor U10425 (N_10425,N_8752,N_7577);
xor U10426 (N_10426,N_8272,N_7091);
xor U10427 (N_10427,N_8395,N_6534);
and U10428 (N_10428,N_8374,N_7117);
xor U10429 (N_10429,N_8022,N_7376);
and U10430 (N_10430,N_7931,N_6258);
nor U10431 (N_10431,N_7695,N_6241);
nand U10432 (N_10432,N_7121,N_8367);
xor U10433 (N_10433,N_6928,N_6610);
nor U10434 (N_10434,N_6707,N_6768);
and U10435 (N_10435,N_8013,N_6820);
and U10436 (N_10436,N_7951,N_8082);
xor U10437 (N_10437,N_6173,N_6696);
xor U10438 (N_10438,N_8957,N_6748);
nor U10439 (N_10439,N_6811,N_6425);
and U10440 (N_10440,N_8677,N_6902);
nor U10441 (N_10441,N_8090,N_6114);
xor U10442 (N_10442,N_7254,N_6233);
nor U10443 (N_10443,N_6947,N_7236);
or U10444 (N_10444,N_7095,N_8181);
xor U10445 (N_10445,N_8377,N_7403);
nand U10446 (N_10446,N_6866,N_7522);
xnor U10447 (N_10447,N_7306,N_6183);
xor U10448 (N_10448,N_7124,N_7419);
xor U10449 (N_10449,N_7134,N_8385);
and U10450 (N_10450,N_8609,N_7600);
or U10451 (N_10451,N_7836,N_7518);
xnor U10452 (N_10452,N_8032,N_8448);
xor U10453 (N_10453,N_6010,N_6686);
or U10454 (N_10454,N_7933,N_7054);
or U10455 (N_10455,N_7620,N_7084);
nand U10456 (N_10456,N_8311,N_7275);
xor U10457 (N_10457,N_6100,N_8740);
and U10458 (N_10458,N_7359,N_7437);
or U10459 (N_10459,N_8578,N_8802);
nor U10460 (N_10460,N_7404,N_7106);
or U10461 (N_10461,N_7187,N_8195);
or U10462 (N_10462,N_8863,N_7057);
or U10463 (N_10463,N_8877,N_7351);
and U10464 (N_10464,N_7845,N_7711);
xnor U10465 (N_10465,N_8197,N_7559);
nor U10466 (N_10466,N_8211,N_6868);
nand U10467 (N_10467,N_7962,N_6267);
or U10468 (N_10468,N_7755,N_6073);
or U10469 (N_10469,N_8612,N_8389);
nor U10470 (N_10470,N_8208,N_6217);
and U10471 (N_10471,N_7310,N_6050);
xnor U10472 (N_10472,N_8288,N_6861);
nor U10473 (N_10473,N_8321,N_8689);
nand U10474 (N_10474,N_6499,N_7975);
xor U10475 (N_10475,N_7943,N_8457);
nor U10476 (N_10476,N_8215,N_6633);
nor U10477 (N_10477,N_6435,N_6573);
xnor U10478 (N_10478,N_6620,N_6974);
xor U10479 (N_10479,N_6213,N_8931);
xnor U10480 (N_10480,N_8274,N_7258);
or U10481 (N_10481,N_6847,N_7070);
and U10482 (N_10482,N_8979,N_6643);
nand U10483 (N_10483,N_6080,N_6851);
and U10484 (N_10484,N_8975,N_7051);
and U10485 (N_10485,N_7358,N_6024);
nand U10486 (N_10486,N_8793,N_7833);
xnor U10487 (N_10487,N_7753,N_7130);
or U10488 (N_10488,N_8441,N_7979);
nand U10489 (N_10489,N_7207,N_8491);
or U10490 (N_10490,N_7215,N_7182);
nand U10491 (N_10491,N_6166,N_8981);
nand U10492 (N_10492,N_8069,N_8929);
or U10493 (N_10493,N_7123,N_8625);
nand U10494 (N_10494,N_6279,N_6254);
xnor U10495 (N_10495,N_6037,N_6721);
nor U10496 (N_10496,N_8227,N_7812);
nor U10497 (N_10497,N_7331,N_8850);
or U10498 (N_10498,N_6685,N_6594);
or U10499 (N_10499,N_8016,N_6180);
xor U10500 (N_10500,N_7750,N_6444);
xor U10501 (N_10501,N_7457,N_7239);
nor U10502 (N_10502,N_7042,N_6329);
or U10503 (N_10503,N_7730,N_8489);
or U10504 (N_10504,N_7171,N_7715);
or U10505 (N_10505,N_8826,N_7535);
nand U10506 (N_10506,N_7486,N_8793);
nor U10507 (N_10507,N_8923,N_7886);
or U10508 (N_10508,N_8627,N_7190);
and U10509 (N_10509,N_6725,N_8880);
nor U10510 (N_10510,N_8419,N_7389);
xnor U10511 (N_10511,N_8847,N_7929);
and U10512 (N_10512,N_7765,N_6538);
nor U10513 (N_10513,N_7797,N_8496);
xor U10514 (N_10514,N_8682,N_7607);
and U10515 (N_10515,N_6336,N_6040);
nand U10516 (N_10516,N_7274,N_8237);
xor U10517 (N_10517,N_7681,N_7580);
or U10518 (N_10518,N_7476,N_7871);
nand U10519 (N_10519,N_8004,N_6714);
or U10520 (N_10520,N_8261,N_6122);
or U10521 (N_10521,N_8507,N_7773);
xnor U10522 (N_10522,N_7913,N_7869);
nand U10523 (N_10523,N_8702,N_8663);
xnor U10524 (N_10524,N_6945,N_8006);
and U10525 (N_10525,N_6102,N_8514);
xnor U10526 (N_10526,N_8844,N_7836);
nor U10527 (N_10527,N_8827,N_8864);
xnor U10528 (N_10528,N_6490,N_8425);
nand U10529 (N_10529,N_8101,N_6969);
or U10530 (N_10530,N_8871,N_7219);
or U10531 (N_10531,N_7352,N_8026);
nor U10532 (N_10532,N_7611,N_8916);
nor U10533 (N_10533,N_7848,N_8938);
and U10534 (N_10534,N_8710,N_8038);
nor U10535 (N_10535,N_8060,N_6594);
and U10536 (N_10536,N_7937,N_7542);
and U10537 (N_10537,N_7115,N_8046);
or U10538 (N_10538,N_7437,N_6983);
nand U10539 (N_10539,N_6535,N_7100);
nand U10540 (N_10540,N_6304,N_8625);
xnor U10541 (N_10541,N_8215,N_8127);
or U10542 (N_10542,N_7413,N_8772);
nand U10543 (N_10543,N_7951,N_6500);
nor U10544 (N_10544,N_7947,N_8799);
xor U10545 (N_10545,N_6283,N_7299);
nor U10546 (N_10546,N_8297,N_6325);
or U10547 (N_10547,N_7748,N_8333);
or U10548 (N_10548,N_6283,N_8313);
or U10549 (N_10549,N_7618,N_6102);
nor U10550 (N_10550,N_7070,N_8123);
xnor U10551 (N_10551,N_6714,N_7150);
xnor U10552 (N_10552,N_8601,N_8467);
nor U10553 (N_10553,N_7309,N_6162);
xor U10554 (N_10554,N_8651,N_7370);
xor U10555 (N_10555,N_6796,N_6988);
and U10556 (N_10556,N_8378,N_6223);
nand U10557 (N_10557,N_6917,N_8547);
nor U10558 (N_10558,N_7397,N_7317);
nand U10559 (N_10559,N_8600,N_8341);
and U10560 (N_10560,N_8339,N_7406);
and U10561 (N_10561,N_8562,N_7291);
and U10562 (N_10562,N_7423,N_7368);
or U10563 (N_10563,N_8629,N_7017);
or U10564 (N_10564,N_8683,N_6855);
and U10565 (N_10565,N_7624,N_7873);
or U10566 (N_10566,N_7964,N_7668);
and U10567 (N_10567,N_6835,N_8517);
nand U10568 (N_10568,N_8117,N_6816);
nand U10569 (N_10569,N_6415,N_6221);
nor U10570 (N_10570,N_8652,N_8762);
xor U10571 (N_10571,N_6651,N_6789);
xor U10572 (N_10572,N_8839,N_6926);
and U10573 (N_10573,N_6283,N_7291);
or U10574 (N_10574,N_8616,N_6517);
nand U10575 (N_10575,N_6486,N_6243);
and U10576 (N_10576,N_8073,N_6880);
nor U10577 (N_10577,N_8893,N_8974);
xor U10578 (N_10578,N_6199,N_8058);
xnor U10579 (N_10579,N_6236,N_8110);
and U10580 (N_10580,N_8185,N_7403);
and U10581 (N_10581,N_6440,N_6872);
and U10582 (N_10582,N_7360,N_8656);
and U10583 (N_10583,N_6604,N_7494);
nand U10584 (N_10584,N_8264,N_8635);
and U10585 (N_10585,N_8511,N_8135);
nor U10586 (N_10586,N_6129,N_7998);
and U10587 (N_10587,N_6712,N_8396);
and U10588 (N_10588,N_7419,N_6620);
nor U10589 (N_10589,N_6317,N_8802);
nand U10590 (N_10590,N_7797,N_7347);
nor U10591 (N_10591,N_7178,N_6942);
nand U10592 (N_10592,N_6473,N_8348);
or U10593 (N_10593,N_6595,N_7903);
nor U10594 (N_10594,N_6207,N_7019);
nand U10595 (N_10595,N_6919,N_7340);
nand U10596 (N_10596,N_6444,N_8370);
xnor U10597 (N_10597,N_8280,N_8119);
xor U10598 (N_10598,N_7091,N_6206);
xnor U10599 (N_10599,N_7042,N_7641);
or U10600 (N_10600,N_8430,N_8243);
nand U10601 (N_10601,N_8728,N_7455);
and U10602 (N_10602,N_8749,N_7899);
nor U10603 (N_10603,N_8655,N_7979);
and U10604 (N_10604,N_6024,N_6086);
nand U10605 (N_10605,N_7541,N_8395);
and U10606 (N_10606,N_8466,N_8705);
or U10607 (N_10607,N_7590,N_7726);
xnor U10608 (N_10608,N_7572,N_7873);
and U10609 (N_10609,N_8915,N_6920);
and U10610 (N_10610,N_7726,N_7340);
nand U10611 (N_10611,N_6140,N_7820);
nor U10612 (N_10612,N_6598,N_7272);
nand U10613 (N_10613,N_8567,N_8282);
xor U10614 (N_10614,N_7062,N_7338);
nor U10615 (N_10615,N_6248,N_7307);
or U10616 (N_10616,N_6343,N_8316);
nor U10617 (N_10617,N_8516,N_8687);
nor U10618 (N_10618,N_6349,N_6602);
nor U10619 (N_10619,N_8887,N_7076);
or U10620 (N_10620,N_6420,N_7807);
nor U10621 (N_10621,N_7122,N_7702);
nand U10622 (N_10622,N_6172,N_7806);
or U10623 (N_10623,N_8085,N_7531);
xnor U10624 (N_10624,N_7565,N_8622);
or U10625 (N_10625,N_8010,N_7787);
xor U10626 (N_10626,N_6728,N_6048);
xor U10627 (N_10627,N_6974,N_6135);
nor U10628 (N_10628,N_7296,N_8500);
nor U10629 (N_10629,N_7176,N_6088);
xor U10630 (N_10630,N_7632,N_7946);
nand U10631 (N_10631,N_7781,N_7935);
nor U10632 (N_10632,N_8679,N_6792);
xnor U10633 (N_10633,N_7601,N_6307);
xor U10634 (N_10634,N_8817,N_7585);
and U10635 (N_10635,N_7344,N_8857);
or U10636 (N_10636,N_7924,N_6634);
xor U10637 (N_10637,N_8838,N_8971);
nand U10638 (N_10638,N_7282,N_8050);
or U10639 (N_10639,N_8471,N_7328);
nor U10640 (N_10640,N_8478,N_7214);
nand U10641 (N_10641,N_6279,N_6957);
or U10642 (N_10642,N_7454,N_8452);
xnor U10643 (N_10643,N_6079,N_8718);
nand U10644 (N_10644,N_6706,N_7753);
nand U10645 (N_10645,N_8511,N_8286);
or U10646 (N_10646,N_7121,N_8956);
nor U10647 (N_10647,N_6406,N_6284);
or U10648 (N_10648,N_6081,N_7462);
or U10649 (N_10649,N_8378,N_7287);
or U10650 (N_10650,N_7897,N_8712);
xnor U10651 (N_10651,N_7704,N_8515);
nand U10652 (N_10652,N_8583,N_8179);
or U10653 (N_10653,N_8123,N_6217);
nand U10654 (N_10654,N_8920,N_6701);
and U10655 (N_10655,N_7086,N_8181);
or U10656 (N_10656,N_7717,N_6270);
nor U10657 (N_10657,N_8337,N_6378);
nand U10658 (N_10658,N_8491,N_8885);
xor U10659 (N_10659,N_7512,N_6451);
and U10660 (N_10660,N_7085,N_8467);
nand U10661 (N_10661,N_7581,N_6170);
xnor U10662 (N_10662,N_8288,N_8350);
xnor U10663 (N_10663,N_7796,N_6412);
nand U10664 (N_10664,N_6428,N_7422);
or U10665 (N_10665,N_8647,N_7286);
nor U10666 (N_10666,N_7330,N_7739);
xor U10667 (N_10667,N_7536,N_8518);
nand U10668 (N_10668,N_7557,N_8422);
nor U10669 (N_10669,N_8934,N_7969);
xor U10670 (N_10670,N_8426,N_8491);
nor U10671 (N_10671,N_7428,N_6483);
xnor U10672 (N_10672,N_6831,N_6286);
and U10673 (N_10673,N_7588,N_8788);
or U10674 (N_10674,N_8240,N_7825);
xnor U10675 (N_10675,N_8512,N_7357);
and U10676 (N_10676,N_6364,N_7124);
or U10677 (N_10677,N_8676,N_8862);
or U10678 (N_10678,N_6983,N_6972);
and U10679 (N_10679,N_6234,N_6377);
or U10680 (N_10680,N_6990,N_8670);
xor U10681 (N_10681,N_8749,N_8212);
nand U10682 (N_10682,N_8879,N_7907);
xnor U10683 (N_10683,N_7777,N_6365);
nand U10684 (N_10684,N_8943,N_6226);
and U10685 (N_10685,N_6290,N_6938);
or U10686 (N_10686,N_6630,N_8911);
and U10687 (N_10687,N_6335,N_7155);
and U10688 (N_10688,N_6148,N_8474);
xnor U10689 (N_10689,N_8532,N_7341);
or U10690 (N_10690,N_6422,N_6080);
and U10691 (N_10691,N_7552,N_8578);
xnor U10692 (N_10692,N_7683,N_7092);
and U10693 (N_10693,N_8547,N_8586);
nor U10694 (N_10694,N_6913,N_8087);
nor U10695 (N_10695,N_7017,N_6667);
nand U10696 (N_10696,N_7195,N_8361);
nor U10697 (N_10697,N_8374,N_7832);
or U10698 (N_10698,N_6512,N_7869);
or U10699 (N_10699,N_7484,N_6051);
nand U10700 (N_10700,N_8663,N_8690);
and U10701 (N_10701,N_6584,N_7492);
and U10702 (N_10702,N_7010,N_7531);
and U10703 (N_10703,N_8008,N_6265);
or U10704 (N_10704,N_6824,N_7993);
or U10705 (N_10705,N_7633,N_6764);
nor U10706 (N_10706,N_6002,N_6524);
nor U10707 (N_10707,N_8614,N_7738);
and U10708 (N_10708,N_6438,N_8396);
nor U10709 (N_10709,N_6717,N_8165);
nand U10710 (N_10710,N_8180,N_8538);
xor U10711 (N_10711,N_6076,N_7887);
and U10712 (N_10712,N_7488,N_8898);
or U10713 (N_10713,N_6729,N_6063);
nand U10714 (N_10714,N_8440,N_7995);
nand U10715 (N_10715,N_6145,N_6381);
nor U10716 (N_10716,N_6681,N_7691);
nor U10717 (N_10717,N_6814,N_8932);
xor U10718 (N_10718,N_6971,N_6414);
xor U10719 (N_10719,N_6200,N_7532);
xnor U10720 (N_10720,N_8054,N_6734);
and U10721 (N_10721,N_8358,N_6723);
and U10722 (N_10722,N_6041,N_7516);
or U10723 (N_10723,N_6976,N_8924);
nand U10724 (N_10724,N_8913,N_8177);
or U10725 (N_10725,N_8286,N_7313);
or U10726 (N_10726,N_6514,N_6654);
or U10727 (N_10727,N_6254,N_7156);
xor U10728 (N_10728,N_6131,N_6099);
and U10729 (N_10729,N_6970,N_6162);
xor U10730 (N_10730,N_6748,N_8844);
nor U10731 (N_10731,N_7607,N_6564);
or U10732 (N_10732,N_6827,N_6539);
nor U10733 (N_10733,N_7649,N_8803);
nor U10734 (N_10734,N_6230,N_7142);
or U10735 (N_10735,N_8266,N_8548);
nor U10736 (N_10736,N_7952,N_8568);
xnor U10737 (N_10737,N_6173,N_8775);
or U10738 (N_10738,N_6063,N_8703);
or U10739 (N_10739,N_6904,N_8454);
xnor U10740 (N_10740,N_6589,N_7885);
or U10741 (N_10741,N_6778,N_6677);
nor U10742 (N_10742,N_8299,N_7601);
nand U10743 (N_10743,N_7087,N_8049);
xor U10744 (N_10744,N_6656,N_6173);
nor U10745 (N_10745,N_6096,N_8679);
or U10746 (N_10746,N_8484,N_8488);
and U10747 (N_10747,N_7509,N_6120);
nor U10748 (N_10748,N_6593,N_8650);
xnor U10749 (N_10749,N_7380,N_8180);
and U10750 (N_10750,N_7382,N_8900);
nor U10751 (N_10751,N_8905,N_8927);
xnor U10752 (N_10752,N_6521,N_6613);
or U10753 (N_10753,N_7687,N_6076);
xor U10754 (N_10754,N_8644,N_7686);
nand U10755 (N_10755,N_6129,N_6919);
nand U10756 (N_10756,N_6146,N_7863);
and U10757 (N_10757,N_8583,N_6990);
and U10758 (N_10758,N_8100,N_8624);
nand U10759 (N_10759,N_8562,N_6107);
and U10760 (N_10760,N_7105,N_7796);
or U10761 (N_10761,N_7736,N_6659);
xnor U10762 (N_10762,N_7231,N_7666);
or U10763 (N_10763,N_8092,N_6745);
or U10764 (N_10764,N_7847,N_6432);
xor U10765 (N_10765,N_6603,N_7681);
and U10766 (N_10766,N_7601,N_6841);
xor U10767 (N_10767,N_8430,N_8614);
nand U10768 (N_10768,N_6140,N_6305);
nor U10769 (N_10769,N_6031,N_8611);
nand U10770 (N_10770,N_6743,N_6939);
and U10771 (N_10771,N_6062,N_7407);
nand U10772 (N_10772,N_7082,N_6281);
xnor U10773 (N_10773,N_6766,N_7152);
nor U10774 (N_10774,N_8205,N_7802);
nand U10775 (N_10775,N_6557,N_6288);
nand U10776 (N_10776,N_6760,N_8493);
nor U10777 (N_10777,N_7041,N_6422);
and U10778 (N_10778,N_6896,N_7042);
xnor U10779 (N_10779,N_8981,N_8628);
nand U10780 (N_10780,N_6395,N_8794);
xnor U10781 (N_10781,N_7073,N_6801);
and U10782 (N_10782,N_7372,N_8800);
or U10783 (N_10783,N_6067,N_8102);
nor U10784 (N_10784,N_6932,N_6617);
nor U10785 (N_10785,N_6765,N_6646);
or U10786 (N_10786,N_8251,N_6432);
nand U10787 (N_10787,N_7721,N_7764);
nor U10788 (N_10788,N_6751,N_8016);
nand U10789 (N_10789,N_6403,N_8313);
xor U10790 (N_10790,N_8981,N_6640);
and U10791 (N_10791,N_8305,N_8190);
xnor U10792 (N_10792,N_6571,N_6453);
or U10793 (N_10793,N_6848,N_6935);
nor U10794 (N_10794,N_7624,N_7239);
or U10795 (N_10795,N_7652,N_7183);
nand U10796 (N_10796,N_8993,N_7815);
and U10797 (N_10797,N_8082,N_7144);
or U10798 (N_10798,N_6068,N_6751);
or U10799 (N_10799,N_7121,N_8662);
nor U10800 (N_10800,N_6660,N_8085);
nor U10801 (N_10801,N_6919,N_8573);
nor U10802 (N_10802,N_7112,N_7403);
or U10803 (N_10803,N_6066,N_6346);
and U10804 (N_10804,N_7191,N_6499);
nor U10805 (N_10805,N_8629,N_7574);
nor U10806 (N_10806,N_7869,N_6963);
nand U10807 (N_10807,N_6605,N_6549);
and U10808 (N_10808,N_6866,N_8165);
nand U10809 (N_10809,N_6868,N_7375);
nor U10810 (N_10810,N_7053,N_8878);
nand U10811 (N_10811,N_7592,N_6191);
nand U10812 (N_10812,N_8700,N_6743);
and U10813 (N_10813,N_7741,N_7510);
and U10814 (N_10814,N_8415,N_6714);
or U10815 (N_10815,N_7175,N_8669);
or U10816 (N_10816,N_6405,N_8064);
xnor U10817 (N_10817,N_7243,N_7563);
xor U10818 (N_10818,N_8471,N_6295);
xnor U10819 (N_10819,N_7915,N_6205);
xor U10820 (N_10820,N_6858,N_8356);
xor U10821 (N_10821,N_6396,N_7471);
and U10822 (N_10822,N_6776,N_7277);
nand U10823 (N_10823,N_6452,N_8318);
nand U10824 (N_10824,N_6591,N_6521);
nor U10825 (N_10825,N_6643,N_8377);
nand U10826 (N_10826,N_8315,N_7302);
or U10827 (N_10827,N_8919,N_6137);
and U10828 (N_10828,N_8814,N_8715);
nand U10829 (N_10829,N_7874,N_7855);
or U10830 (N_10830,N_8300,N_8514);
nor U10831 (N_10831,N_6230,N_6749);
or U10832 (N_10832,N_7223,N_8697);
nand U10833 (N_10833,N_6884,N_6072);
nor U10834 (N_10834,N_8457,N_8922);
xor U10835 (N_10835,N_8054,N_6762);
nor U10836 (N_10836,N_6024,N_7876);
and U10837 (N_10837,N_6291,N_7273);
and U10838 (N_10838,N_6804,N_6529);
or U10839 (N_10839,N_6977,N_6632);
or U10840 (N_10840,N_8423,N_8524);
and U10841 (N_10841,N_6007,N_6249);
xnor U10842 (N_10842,N_6013,N_8861);
nor U10843 (N_10843,N_7327,N_6842);
and U10844 (N_10844,N_6519,N_7133);
nor U10845 (N_10845,N_6106,N_8221);
nor U10846 (N_10846,N_7821,N_7643);
and U10847 (N_10847,N_7345,N_7481);
or U10848 (N_10848,N_8675,N_6806);
nor U10849 (N_10849,N_7680,N_7314);
or U10850 (N_10850,N_6373,N_7896);
or U10851 (N_10851,N_6790,N_8231);
nand U10852 (N_10852,N_7548,N_7994);
nor U10853 (N_10853,N_8080,N_7946);
xnor U10854 (N_10854,N_8565,N_8544);
and U10855 (N_10855,N_7090,N_8157);
and U10856 (N_10856,N_6852,N_7849);
xor U10857 (N_10857,N_6677,N_8947);
nand U10858 (N_10858,N_6192,N_6457);
and U10859 (N_10859,N_7078,N_8555);
and U10860 (N_10860,N_7082,N_7747);
nand U10861 (N_10861,N_6944,N_6939);
nand U10862 (N_10862,N_6998,N_8346);
nand U10863 (N_10863,N_8134,N_7060);
xnor U10864 (N_10864,N_8615,N_7133);
or U10865 (N_10865,N_8943,N_6533);
and U10866 (N_10866,N_6419,N_8431);
nor U10867 (N_10867,N_6410,N_6275);
nor U10868 (N_10868,N_7665,N_6358);
xor U10869 (N_10869,N_7046,N_7161);
and U10870 (N_10870,N_8571,N_6535);
nor U10871 (N_10871,N_8070,N_8899);
or U10872 (N_10872,N_6111,N_7937);
nor U10873 (N_10873,N_6710,N_6911);
nor U10874 (N_10874,N_6433,N_7247);
and U10875 (N_10875,N_8947,N_7717);
xnor U10876 (N_10876,N_6163,N_6472);
nor U10877 (N_10877,N_7091,N_7678);
or U10878 (N_10878,N_6381,N_7814);
nor U10879 (N_10879,N_7517,N_8861);
or U10880 (N_10880,N_8055,N_8490);
and U10881 (N_10881,N_6138,N_7319);
and U10882 (N_10882,N_6070,N_8503);
nor U10883 (N_10883,N_8287,N_8516);
nand U10884 (N_10884,N_7612,N_7582);
xnor U10885 (N_10885,N_7044,N_8600);
nor U10886 (N_10886,N_6057,N_6738);
nor U10887 (N_10887,N_6856,N_7658);
nand U10888 (N_10888,N_7091,N_6856);
and U10889 (N_10889,N_6140,N_6360);
nand U10890 (N_10890,N_8420,N_7733);
and U10891 (N_10891,N_8170,N_8644);
nand U10892 (N_10892,N_6345,N_7613);
or U10893 (N_10893,N_7769,N_7822);
or U10894 (N_10894,N_7267,N_8862);
nor U10895 (N_10895,N_7086,N_7153);
nand U10896 (N_10896,N_7081,N_8793);
and U10897 (N_10897,N_6241,N_8517);
xor U10898 (N_10898,N_6489,N_8632);
or U10899 (N_10899,N_6605,N_8136);
nand U10900 (N_10900,N_8549,N_8315);
nand U10901 (N_10901,N_8286,N_7809);
or U10902 (N_10902,N_8259,N_7958);
xor U10903 (N_10903,N_6119,N_7037);
nor U10904 (N_10904,N_6664,N_6633);
or U10905 (N_10905,N_6299,N_6603);
nand U10906 (N_10906,N_8447,N_8810);
or U10907 (N_10907,N_8654,N_6887);
nor U10908 (N_10908,N_6658,N_8511);
nand U10909 (N_10909,N_7378,N_6964);
or U10910 (N_10910,N_7021,N_7767);
and U10911 (N_10911,N_8960,N_6674);
and U10912 (N_10912,N_8198,N_8665);
and U10913 (N_10913,N_7848,N_6436);
xor U10914 (N_10914,N_6225,N_6369);
nand U10915 (N_10915,N_6847,N_8118);
and U10916 (N_10916,N_6660,N_6567);
and U10917 (N_10917,N_6712,N_8953);
nor U10918 (N_10918,N_7655,N_8085);
and U10919 (N_10919,N_7543,N_7366);
xor U10920 (N_10920,N_7766,N_6097);
nand U10921 (N_10921,N_6245,N_6159);
xnor U10922 (N_10922,N_7306,N_8463);
xnor U10923 (N_10923,N_8142,N_8726);
nand U10924 (N_10924,N_6505,N_6419);
nor U10925 (N_10925,N_6553,N_6559);
and U10926 (N_10926,N_6540,N_7539);
and U10927 (N_10927,N_8469,N_7673);
or U10928 (N_10928,N_8135,N_7035);
and U10929 (N_10929,N_8063,N_6652);
xnor U10930 (N_10930,N_8226,N_6141);
nor U10931 (N_10931,N_7320,N_6705);
and U10932 (N_10932,N_8959,N_7366);
or U10933 (N_10933,N_8916,N_7678);
nor U10934 (N_10934,N_6699,N_8026);
or U10935 (N_10935,N_7288,N_8269);
nand U10936 (N_10936,N_8357,N_7026);
or U10937 (N_10937,N_8745,N_6855);
nor U10938 (N_10938,N_8507,N_8478);
nor U10939 (N_10939,N_6509,N_7436);
and U10940 (N_10940,N_8983,N_7130);
xnor U10941 (N_10941,N_6893,N_6322);
nor U10942 (N_10942,N_7188,N_7698);
and U10943 (N_10943,N_8221,N_6363);
nor U10944 (N_10944,N_6548,N_8980);
xor U10945 (N_10945,N_7135,N_6687);
or U10946 (N_10946,N_8829,N_8001);
nand U10947 (N_10947,N_7768,N_6314);
xor U10948 (N_10948,N_6059,N_8629);
nor U10949 (N_10949,N_7923,N_7988);
xor U10950 (N_10950,N_6379,N_6715);
and U10951 (N_10951,N_6401,N_8073);
nor U10952 (N_10952,N_7759,N_6151);
nand U10953 (N_10953,N_8911,N_6267);
nand U10954 (N_10954,N_7368,N_6408);
nand U10955 (N_10955,N_6510,N_6529);
nor U10956 (N_10956,N_8511,N_7242);
nor U10957 (N_10957,N_8496,N_6522);
xnor U10958 (N_10958,N_8717,N_7243);
nor U10959 (N_10959,N_8554,N_8879);
nand U10960 (N_10960,N_7298,N_7430);
xor U10961 (N_10961,N_7809,N_6889);
nand U10962 (N_10962,N_6370,N_7367);
nand U10963 (N_10963,N_6676,N_6869);
and U10964 (N_10964,N_8504,N_7637);
and U10965 (N_10965,N_7602,N_8331);
and U10966 (N_10966,N_6409,N_8910);
xnor U10967 (N_10967,N_7883,N_8521);
and U10968 (N_10968,N_8984,N_7379);
nand U10969 (N_10969,N_7076,N_6282);
nor U10970 (N_10970,N_8561,N_7191);
xor U10971 (N_10971,N_8026,N_7858);
or U10972 (N_10972,N_7870,N_6408);
or U10973 (N_10973,N_7759,N_7327);
xor U10974 (N_10974,N_7971,N_7919);
nor U10975 (N_10975,N_6843,N_8901);
nand U10976 (N_10976,N_6988,N_8321);
nor U10977 (N_10977,N_7752,N_6646);
xor U10978 (N_10978,N_6450,N_7342);
nor U10979 (N_10979,N_8087,N_6940);
nor U10980 (N_10980,N_7779,N_7392);
nor U10981 (N_10981,N_7352,N_6412);
nand U10982 (N_10982,N_7644,N_8447);
and U10983 (N_10983,N_6473,N_6379);
xor U10984 (N_10984,N_8070,N_8328);
xnor U10985 (N_10985,N_8485,N_6609);
or U10986 (N_10986,N_8850,N_6379);
or U10987 (N_10987,N_6193,N_6534);
nor U10988 (N_10988,N_6116,N_7616);
or U10989 (N_10989,N_6692,N_6197);
xor U10990 (N_10990,N_7168,N_6922);
nor U10991 (N_10991,N_7984,N_7410);
nor U10992 (N_10992,N_8624,N_8927);
xnor U10993 (N_10993,N_8676,N_6236);
or U10994 (N_10994,N_7823,N_7277);
and U10995 (N_10995,N_8762,N_6128);
or U10996 (N_10996,N_6773,N_8042);
nand U10997 (N_10997,N_8781,N_6041);
nand U10998 (N_10998,N_7506,N_7162);
nand U10999 (N_10999,N_6591,N_7921);
nand U11000 (N_11000,N_8515,N_8220);
xnor U11001 (N_11001,N_8684,N_6888);
xor U11002 (N_11002,N_8292,N_7617);
nand U11003 (N_11003,N_7861,N_8766);
or U11004 (N_11004,N_6554,N_7733);
nand U11005 (N_11005,N_8755,N_8996);
or U11006 (N_11006,N_6323,N_6435);
and U11007 (N_11007,N_7712,N_7964);
xnor U11008 (N_11008,N_6943,N_8249);
nor U11009 (N_11009,N_6149,N_6463);
or U11010 (N_11010,N_8498,N_7500);
nor U11011 (N_11011,N_7777,N_6806);
nand U11012 (N_11012,N_6538,N_7826);
and U11013 (N_11013,N_6439,N_8316);
nor U11014 (N_11014,N_8678,N_8599);
or U11015 (N_11015,N_6845,N_8970);
or U11016 (N_11016,N_7788,N_8945);
or U11017 (N_11017,N_7132,N_8254);
xnor U11018 (N_11018,N_8069,N_7443);
nand U11019 (N_11019,N_7584,N_8501);
nand U11020 (N_11020,N_6821,N_7208);
and U11021 (N_11021,N_7844,N_8813);
and U11022 (N_11022,N_6434,N_7602);
nor U11023 (N_11023,N_6335,N_8497);
and U11024 (N_11024,N_6877,N_7320);
nand U11025 (N_11025,N_6733,N_8051);
nor U11026 (N_11026,N_6186,N_7152);
nand U11027 (N_11027,N_8575,N_6093);
or U11028 (N_11028,N_7248,N_6392);
or U11029 (N_11029,N_7546,N_6058);
xnor U11030 (N_11030,N_6460,N_7736);
nor U11031 (N_11031,N_6146,N_6228);
xor U11032 (N_11032,N_6730,N_6076);
or U11033 (N_11033,N_8772,N_8895);
and U11034 (N_11034,N_8124,N_6160);
xor U11035 (N_11035,N_7637,N_8659);
nor U11036 (N_11036,N_8611,N_7656);
nor U11037 (N_11037,N_8145,N_7562);
or U11038 (N_11038,N_6987,N_6712);
or U11039 (N_11039,N_6070,N_6406);
xnor U11040 (N_11040,N_6863,N_8865);
or U11041 (N_11041,N_7555,N_6418);
or U11042 (N_11042,N_8477,N_6943);
and U11043 (N_11043,N_7663,N_7767);
nor U11044 (N_11044,N_8331,N_6582);
or U11045 (N_11045,N_7684,N_6355);
or U11046 (N_11046,N_6371,N_7274);
or U11047 (N_11047,N_8050,N_6670);
xor U11048 (N_11048,N_7649,N_7905);
xnor U11049 (N_11049,N_8499,N_6138);
nand U11050 (N_11050,N_7327,N_6377);
or U11051 (N_11051,N_6158,N_7495);
nand U11052 (N_11052,N_7425,N_7782);
nor U11053 (N_11053,N_7688,N_7631);
nand U11054 (N_11054,N_7658,N_6596);
or U11055 (N_11055,N_8575,N_8909);
and U11056 (N_11056,N_7303,N_8691);
nand U11057 (N_11057,N_6532,N_8671);
xor U11058 (N_11058,N_8337,N_8295);
and U11059 (N_11059,N_8381,N_6029);
xnor U11060 (N_11060,N_8499,N_7205);
or U11061 (N_11061,N_8528,N_8589);
xor U11062 (N_11062,N_6150,N_6831);
or U11063 (N_11063,N_7928,N_7483);
and U11064 (N_11064,N_7639,N_6238);
and U11065 (N_11065,N_6481,N_6633);
nand U11066 (N_11066,N_6139,N_7073);
nor U11067 (N_11067,N_8693,N_8913);
nor U11068 (N_11068,N_8896,N_6600);
nand U11069 (N_11069,N_8195,N_6064);
or U11070 (N_11070,N_8493,N_7016);
and U11071 (N_11071,N_7076,N_8509);
nand U11072 (N_11072,N_7655,N_7145);
xor U11073 (N_11073,N_8646,N_7126);
nor U11074 (N_11074,N_7289,N_6470);
or U11075 (N_11075,N_8870,N_8506);
and U11076 (N_11076,N_8228,N_8007);
nor U11077 (N_11077,N_6537,N_6568);
or U11078 (N_11078,N_7511,N_6306);
xnor U11079 (N_11079,N_6226,N_7591);
nor U11080 (N_11080,N_6933,N_6871);
nand U11081 (N_11081,N_6866,N_6043);
or U11082 (N_11082,N_6861,N_6002);
nand U11083 (N_11083,N_7024,N_6045);
or U11084 (N_11084,N_6689,N_7202);
nor U11085 (N_11085,N_6034,N_7246);
xnor U11086 (N_11086,N_8839,N_7162);
xor U11087 (N_11087,N_7895,N_6554);
and U11088 (N_11088,N_6349,N_6245);
or U11089 (N_11089,N_7545,N_8735);
nand U11090 (N_11090,N_7271,N_6550);
xnor U11091 (N_11091,N_7977,N_8853);
and U11092 (N_11092,N_7559,N_6258);
or U11093 (N_11093,N_6733,N_6488);
or U11094 (N_11094,N_7752,N_6038);
nor U11095 (N_11095,N_8559,N_7008);
xor U11096 (N_11096,N_6720,N_6500);
xnor U11097 (N_11097,N_6886,N_8894);
nand U11098 (N_11098,N_6356,N_8005);
nand U11099 (N_11099,N_8108,N_6800);
nor U11100 (N_11100,N_8240,N_7617);
or U11101 (N_11101,N_8679,N_6149);
and U11102 (N_11102,N_8902,N_6817);
nor U11103 (N_11103,N_8818,N_8988);
and U11104 (N_11104,N_6974,N_8266);
and U11105 (N_11105,N_7419,N_6509);
xor U11106 (N_11106,N_6449,N_8169);
or U11107 (N_11107,N_7403,N_7357);
nor U11108 (N_11108,N_8219,N_6058);
or U11109 (N_11109,N_6426,N_6537);
nor U11110 (N_11110,N_7167,N_6571);
xnor U11111 (N_11111,N_7803,N_7814);
and U11112 (N_11112,N_7612,N_8390);
nand U11113 (N_11113,N_8759,N_6503);
nand U11114 (N_11114,N_8964,N_8920);
nand U11115 (N_11115,N_7336,N_8059);
and U11116 (N_11116,N_8510,N_8999);
or U11117 (N_11117,N_7044,N_6910);
nand U11118 (N_11118,N_8998,N_7999);
and U11119 (N_11119,N_7555,N_7941);
and U11120 (N_11120,N_6089,N_7141);
and U11121 (N_11121,N_6796,N_6497);
nor U11122 (N_11122,N_8255,N_8648);
or U11123 (N_11123,N_8158,N_6284);
and U11124 (N_11124,N_6099,N_7393);
or U11125 (N_11125,N_8937,N_8489);
nor U11126 (N_11126,N_8381,N_8363);
and U11127 (N_11127,N_7715,N_6686);
nor U11128 (N_11128,N_7289,N_8277);
or U11129 (N_11129,N_7354,N_8835);
nor U11130 (N_11130,N_6240,N_8834);
and U11131 (N_11131,N_8044,N_6936);
xnor U11132 (N_11132,N_7638,N_8478);
nand U11133 (N_11133,N_8105,N_6382);
xor U11134 (N_11134,N_7768,N_8947);
nand U11135 (N_11135,N_7036,N_6820);
nor U11136 (N_11136,N_8710,N_6888);
nor U11137 (N_11137,N_8585,N_6678);
or U11138 (N_11138,N_6501,N_6849);
and U11139 (N_11139,N_7051,N_8357);
nand U11140 (N_11140,N_7345,N_7850);
xor U11141 (N_11141,N_6184,N_8228);
and U11142 (N_11142,N_6470,N_7076);
and U11143 (N_11143,N_8578,N_8368);
or U11144 (N_11144,N_7517,N_8868);
nor U11145 (N_11145,N_7791,N_8398);
and U11146 (N_11146,N_7456,N_6285);
xor U11147 (N_11147,N_7724,N_8208);
or U11148 (N_11148,N_7754,N_8950);
nand U11149 (N_11149,N_7644,N_8519);
and U11150 (N_11150,N_8712,N_8865);
or U11151 (N_11151,N_6135,N_8220);
or U11152 (N_11152,N_7803,N_6678);
and U11153 (N_11153,N_7340,N_7134);
and U11154 (N_11154,N_8416,N_7052);
xor U11155 (N_11155,N_6943,N_8620);
and U11156 (N_11156,N_7504,N_6580);
and U11157 (N_11157,N_6534,N_6303);
nand U11158 (N_11158,N_6731,N_7520);
and U11159 (N_11159,N_7748,N_7993);
xor U11160 (N_11160,N_8390,N_6766);
xor U11161 (N_11161,N_8476,N_7543);
nand U11162 (N_11162,N_8099,N_7706);
xnor U11163 (N_11163,N_7114,N_8424);
xor U11164 (N_11164,N_8530,N_7335);
xnor U11165 (N_11165,N_6990,N_6895);
nor U11166 (N_11166,N_8917,N_8563);
xor U11167 (N_11167,N_6022,N_8597);
nand U11168 (N_11168,N_8632,N_6754);
and U11169 (N_11169,N_7118,N_7737);
and U11170 (N_11170,N_6755,N_6496);
nand U11171 (N_11171,N_6885,N_7665);
or U11172 (N_11172,N_7141,N_6080);
nor U11173 (N_11173,N_8510,N_6361);
and U11174 (N_11174,N_7634,N_8447);
or U11175 (N_11175,N_7404,N_7891);
and U11176 (N_11176,N_7962,N_6864);
xor U11177 (N_11177,N_7702,N_7515);
or U11178 (N_11178,N_8700,N_7733);
xor U11179 (N_11179,N_6697,N_8004);
and U11180 (N_11180,N_7876,N_7400);
xor U11181 (N_11181,N_8285,N_8612);
and U11182 (N_11182,N_6853,N_7530);
nand U11183 (N_11183,N_8257,N_7331);
or U11184 (N_11184,N_8875,N_6847);
xor U11185 (N_11185,N_6446,N_8434);
nand U11186 (N_11186,N_6921,N_6939);
nor U11187 (N_11187,N_7443,N_8642);
nand U11188 (N_11188,N_6777,N_8206);
or U11189 (N_11189,N_6774,N_8565);
xnor U11190 (N_11190,N_6522,N_6356);
or U11191 (N_11191,N_6831,N_8004);
nand U11192 (N_11192,N_6869,N_7126);
nor U11193 (N_11193,N_7786,N_6627);
and U11194 (N_11194,N_6976,N_7610);
nand U11195 (N_11195,N_6226,N_7624);
and U11196 (N_11196,N_7782,N_8876);
nand U11197 (N_11197,N_6082,N_7652);
xor U11198 (N_11198,N_8552,N_6924);
xnor U11199 (N_11199,N_8866,N_6205);
nand U11200 (N_11200,N_6310,N_7389);
xnor U11201 (N_11201,N_7392,N_6102);
xnor U11202 (N_11202,N_7966,N_6077);
xor U11203 (N_11203,N_8037,N_8647);
nand U11204 (N_11204,N_7610,N_7780);
nand U11205 (N_11205,N_8764,N_6757);
xnor U11206 (N_11206,N_7068,N_6382);
nor U11207 (N_11207,N_6603,N_6186);
or U11208 (N_11208,N_7525,N_7812);
nor U11209 (N_11209,N_8113,N_6166);
nand U11210 (N_11210,N_8429,N_7300);
and U11211 (N_11211,N_8779,N_6587);
and U11212 (N_11212,N_7547,N_8752);
nand U11213 (N_11213,N_7798,N_8714);
xnor U11214 (N_11214,N_7511,N_6173);
or U11215 (N_11215,N_7376,N_8708);
xor U11216 (N_11216,N_7701,N_7472);
xor U11217 (N_11217,N_7166,N_6207);
nor U11218 (N_11218,N_6504,N_8009);
or U11219 (N_11219,N_6016,N_7920);
nand U11220 (N_11220,N_6923,N_7882);
nor U11221 (N_11221,N_7941,N_7663);
xnor U11222 (N_11222,N_8951,N_6448);
and U11223 (N_11223,N_6747,N_8527);
nand U11224 (N_11224,N_6200,N_6711);
nand U11225 (N_11225,N_6997,N_8660);
or U11226 (N_11226,N_8279,N_7305);
nor U11227 (N_11227,N_8402,N_8215);
and U11228 (N_11228,N_8424,N_8934);
nor U11229 (N_11229,N_6406,N_7291);
nand U11230 (N_11230,N_7030,N_7186);
nand U11231 (N_11231,N_6337,N_6514);
xor U11232 (N_11232,N_7081,N_6246);
nor U11233 (N_11233,N_8785,N_7865);
xor U11234 (N_11234,N_8224,N_7596);
xor U11235 (N_11235,N_7001,N_8913);
nor U11236 (N_11236,N_7307,N_7396);
nor U11237 (N_11237,N_6918,N_8945);
and U11238 (N_11238,N_8634,N_6407);
or U11239 (N_11239,N_7727,N_8668);
nand U11240 (N_11240,N_8058,N_6867);
xor U11241 (N_11241,N_6762,N_6537);
nor U11242 (N_11242,N_7327,N_6239);
xnor U11243 (N_11243,N_8579,N_6839);
xor U11244 (N_11244,N_8710,N_7754);
xor U11245 (N_11245,N_6160,N_6288);
nand U11246 (N_11246,N_6103,N_6166);
and U11247 (N_11247,N_7920,N_8530);
nor U11248 (N_11248,N_7839,N_7622);
nand U11249 (N_11249,N_7390,N_7428);
and U11250 (N_11250,N_7153,N_6059);
nand U11251 (N_11251,N_6763,N_8904);
nor U11252 (N_11252,N_6210,N_7819);
and U11253 (N_11253,N_8991,N_6079);
or U11254 (N_11254,N_8917,N_7402);
nand U11255 (N_11255,N_6659,N_8075);
nor U11256 (N_11256,N_7653,N_7057);
or U11257 (N_11257,N_6194,N_6708);
and U11258 (N_11258,N_7384,N_6003);
xor U11259 (N_11259,N_6968,N_6446);
nand U11260 (N_11260,N_8017,N_7802);
xnor U11261 (N_11261,N_7041,N_7633);
and U11262 (N_11262,N_6245,N_7795);
nor U11263 (N_11263,N_7225,N_6580);
nor U11264 (N_11264,N_8039,N_6526);
nor U11265 (N_11265,N_7640,N_7606);
nor U11266 (N_11266,N_8567,N_8051);
and U11267 (N_11267,N_8515,N_8692);
nor U11268 (N_11268,N_8912,N_8943);
or U11269 (N_11269,N_8879,N_8705);
nand U11270 (N_11270,N_8573,N_8899);
nand U11271 (N_11271,N_7651,N_8934);
xor U11272 (N_11272,N_6397,N_8952);
nand U11273 (N_11273,N_8547,N_6628);
or U11274 (N_11274,N_7565,N_7172);
xor U11275 (N_11275,N_8336,N_8427);
nor U11276 (N_11276,N_7017,N_7848);
nand U11277 (N_11277,N_7109,N_6739);
and U11278 (N_11278,N_7962,N_6803);
nand U11279 (N_11279,N_8668,N_6111);
nand U11280 (N_11280,N_6916,N_7043);
xnor U11281 (N_11281,N_8596,N_8493);
nor U11282 (N_11282,N_6131,N_8751);
and U11283 (N_11283,N_6068,N_7342);
nand U11284 (N_11284,N_7974,N_7559);
nand U11285 (N_11285,N_6504,N_8021);
and U11286 (N_11286,N_6885,N_6916);
nor U11287 (N_11287,N_7800,N_6754);
xor U11288 (N_11288,N_8787,N_7884);
and U11289 (N_11289,N_8664,N_7431);
and U11290 (N_11290,N_8239,N_6465);
nor U11291 (N_11291,N_7876,N_7435);
and U11292 (N_11292,N_8166,N_7256);
nand U11293 (N_11293,N_7875,N_7513);
nor U11294 (N_11294,N_6168,N_7467);
xor U11295 (N_11295,N_6350,N_8171);
and U11296 (N_11296,N_8158,N_8571);
or U11297 (N_11297,N_7317,N_7855);
or U11298 (N_11298,N_7868,N_8493);
xor U11299 (N_11299,N_8891,N_7258);
nand U11300 (N_11300,N_6563,N_6086);
and U11301 (N_11301,N_6874,N_8381);
nor U11302 (N_11302,N_8630,N_6183);
nand U11303 (N_11303,N_6904,N_8384);
and U11304 (N_11304,N_8152,N_8368);
xor U11305 (N_11305,N_6773,N_6172);
nor U11306 (N_11306,N_7780,N_8619);
nor U11307 (N_11307,N_6648,N_6402);
and U11308 (N_11308,N_8096,N_7521);
nand U11309 (N_11309,N_8081,N_6907);
xor U11310 (N_11310,N_8746,N_8281);
nor U11311 (N_11311,N_7961,N_6901);
or U11312 (N_11312,N_7725,N_7971);
and U11313 (N_11313,N_7659,N_7403);
nor U11314 (N_11314,N_8423,N_7637);
nor U11315 (N_11315,N_6989,N_7459);
nor U11316 (N_11316,N_8851,N_6267);
nand U11317 (N_11317,N_6961,N_8371);
nand U11318 (N_11318,N_7261,N_7087);
nand U11319 (N_11319,N_6917,N_8326);
or U11320 (N_11320,N_6039,N_8422);
or U11321 (N_11321,N_8596,N_7746);
xnor U11322 (N_11322,N_7818,N_6900);
nand U11323 (N_11323,N_6104,N_7355);
or U11324 (N_11324,N_8499,N_7753);
nand U11325 (N_11325,N_7362,N_7937);
nor U11326 (N_11326,N_6836,N_6766);
nor U11327 (N_11327,N_6724,N_6899);
nor U11328 (N_11328,N_8879,N_6834);
nor U11329 (N_11329,N_6452,N_8278);
nand U11330 (N_11330,N_8154,N_7978);
or U11331 (N_11331,N_8693,N_8659);
xor U11332 (N_11332,N_6886,N_8399);
or U11333 (N_11333,N_6809,N_6978);
nor U11334 (N_11334,N_8410,N_8544);
xnor U11335 (N_11335,N_6012,N_8639);
and U11336 (N_11336,N_8182,N_8036);
nand U11337 (N_11337,N_8714,N_8872);
and U11338 (N_11338,N_6703,N_8869);
or U11339 (N_11339,N_6546,N_6742);
nand U11340 (N_11340,N_8492,N_8592);
nand U11341 (N_11341,N_7375,N_6862);
nor U11342 (N_11342,N_6248,N_6500);
or U11343 (N_11343,N_7035,N_6184);
nand U11344 (N_11344,N_8055,N_7673);
xor U11345 (N_11345,N_8303,N_7064);
xor U11346 (N_11346,N_6021,N_7468);
or U11347 (N_11347,N_6215,N_6530);
and U11348 (N_11348,N_6114,N_8677);
or U11349 (N_11349,N_7614,N_8210);
xor U11350 (N_11350,N_6087,N_8017);
nor U11351 (N_11351,N_8934,N_7636);
nand U11352 (N_11352,N_7013,N_8733);
nor U11353 (N_11353,N_8310,N_6034);
or U11354 (N_11354,N_7723,N_7435);
nand U11355 (N_11355,N_8762,N_6421);
nand U11356 (N_11356,N_7555,N_6997);
nand U11357 (N_11357,N_6291,N_7034);
nand U11358 (N_11358,N_6120,N_8132);
nor U11359 (N_11359,N_7257,N_6742);
or U11360 (N_11360,N_8617,N_6195);
or U11361 (N_11361,N_6728,N_7050);
nor U11362 (N_11362,N_7621,N_6461);
and U11363 (N_11363,N_6286,N_7012);
nand U11364 (N_11364,N_7839,N_7233);
xor U11365 (N_11365,N_8371,N_8128);
nand U11366 (N_11366,N_7776,N_7345);
nor U11367 (N_11367,N_6143,N_8311);
nor U11368 (N_11368,N_7894,N_7431);
and U11369 (N_11369,N_8653,N_6558);
nand U11370 (N_11370,N_8942,N_6287);
nor U11371 (N_11371,N_7394,N_7073);
nand U11372 (N_11372,N_6947,N_6916);
nor U11373 (N_11373,N_7018,N_7616);
xor U11374 (N_11374,N_6689,N_6198);
or U11375 (N_11375,N_7971,N_6233);
nand U11376 (N_11376,N_6777,N_6427);
nand U11377 (N_11377,N_8297,N_6682);
nor U11378 (N_11378,N_6859,N_7481);
nand U11379 (N_11379,N_6834,N_7822);
xor U11380 (N_11380,N_6491,N_7964);
xor U11381 (N_11381,N_8146,N_8888);
nand U11382 (N_11382,N_6078,N_8080);
or U11383 (N_11383,N_8591,N_8894);
nor U11384 (N_11384,N_8356,N_8838);
and U11385 (N_11385,N_8026,N_8551);
or U11386 (N_11386,N_7222,N_8048);
or U11387 (N_11387,N_6141,N_6153);
and U11388 (N_11388,N_8225,N_7841);
nor U11389 (N_11389,N_7200,N_7673);
xnor U11390 (N_11390,N_7964,N_6114);
or U11391 (N_11391,N_8471,N_8304);
nor U11392 (N_11392,N_6546,N_7726);
xnor U11393 (N_11393,N_8677,N_7516);
nand U11394 (N_11394,N_8831,N_8198);
or U11395 (N_11395,N_8663,N_8749);
nand U11396 (N_11396,N_8761,N_8846);
xnor U11397 (N_11397,N_6451,N_8530);
nand U11398 (N_11398,N_6768,N_7891);
xor U11399 (N_11399,N_6239,N_7722);
xor U11400 (N_11400,N_7233,N_7044);
or U11401 (N_11401,N_6989,N_8890);
nor U11402 (N_11402,N_7387,N_6061);
and U11403 (N_11403,N_7008,N_7436);
nand U11404 (N_11404,N_6437,N_8924);
nor U11405 (N_11405,N_8212,N_6102);
and U11406 (N_11406,N_8150,N_8666);
nand U11407 (N_11407,N_7481,N_7040);
nand U11408 (N_11408,N_6817,N_7918);
nor U11409 (N_11409,N_7891,N_7915);
xnor U11410 (N_11410,N_7927,N_7453);
and U11411 (N_11411,N_7269,N_6769);
and U11412 (N_11412,N_8912,N_7989);
nand U11413 (N_11413,N_6999,N_6774);
and U11414 (N_11414,N_6882,N_7830);
and U11415 (N_11415,N_8253,N_6837);
and U11416 (N_11416,N_7848,N_7790);
nand U11417 (N_11417,N_6511,N_6612);
nor U11418 (N_11418,N_8941,N_6275);
nand U11419 (N_11419,N_6157,N_8619);
xor U11420 (N_11420,N_6997,N_6901);
xnor U11421 (N_11421,N_8597,N_8158);
and U11422 (N_11422,N_8571,N_7431);
xor U11423 (N_11423,N_6500,N_6437);
nand U11424 (N_11424,N_8530,N_7736);
nand U11425 (N_11425,N_6713,N_6975);
xnor U11426 (N_11426,N_7818,N_6688);
or U11427 (N_11427,N_6906,N_6960);
nand U11428 (N_11428,N_7446,N_7550);
xor U11429 (N_11429,N_7770,N_6242);
xor U11430 (N_11430,N_6005,N_8361);
and U11431 (N_11431,N_7906,N_7255);
or U11432 (N_11432,N_7096,N_8695);
nand U11433 (N_11433,N_7148,N_6771);
nor U11434 (N_11434,N_6790,N_7553);
or U11435 (N_11435,N_8241,N_6159);
and U11436 (N_11436,N_6502,N_7159);
xor U11437 (N_11437,N_7610,N_8325);
xnor U11438 (N_11438,N_8628,N_7021);
and U11439 (N_11439,N_7479,N_6208);
nand U11440 (N_11440,N_6212,N_8602);
and U11441 (N_11441,N_7655,N_6367);
and U11442 (N_11442,N_6113,N_8181);
nor U11443 (N_11443,N_8431,N_8472);
xnor U11444 (N_11444,N_6926,N_8285);
nand U11445 (N_11445,N_7466,N_7311);
nor U11446 (N_11446,N_6317,N_7781);
or U11447 (N_11447,N_7535,N_8874);
and U11448 (N_11448,N_7821,N_6957);
or U11449 (N_11449,N_7464,N_8206);
xor U11450 (N_11450,N_8195,N_6154);
or U11451 (N_11451,N_6338,N_7961);
and U11452 (N_11452,N_8317,N_6444);
xnor U11453 (N_11453,N_7618,N_7294);
nand U11454 (N_11454,N_8671,N_8936);
xor U11455 (N_11455,N_8977,N_6375);
or U11456 (N_11456,N_6858,N_8465);
nor U11457 (N_11457,N_8067,N_8883);
nand U11458 (N_11458,N_6039,N_6804);
and U11459 (N_11459,N_8189,N_8776);
and U11460 (N_11460,N_7817,N_7291);
nor U11461 (N_11461,N_6282,N_7746);
and U11462 (N_11462,N_7679,N_8199);
or U11463 (N_11463,N_8483,N_8459);
nor U11464 (N_11464,N_8868,N_8951);
nand U11465 (N_11465,N_6553,N_6271);
or U11466 (N_11466,N_8683,N_6576);
nand U11467 (N_11467,N_8887,N_7940);
xor U11468 (N_11468,N_6598,N_8258);
or U11469 (N_11469,N_7596,N_7277);
and U11470 (N_11470,N_6049,N_6918);
nor U11471 (N_11471,N_8591,N_8598);
nor U11472 (N_11472,N_7521,N_6229);
xnor U11473 (N_11473,N_6445,N_7920);
xnor U11474 (N_11474,N_6081,N_7137);
nor U11475 (N_11475,N_8544,N_8436);
nand U11476 (N_11476,N_6992,N_7891);
nand U11477 (N_11477,N_7430,N_7960);
and U11478 (N_11478,N_6255,N_6202);
or U11479 (N_11479,N_8943,N_6831);
and U11480 (N_11480,N_6060,N_6660);
or U11481 (N_11481,N_8845,N_7047);
and U11482 (N_11482,N_8413,N_6513);
or U11483 (N_11483,N_8720,N_7778);
and U11484 (N_11484,N_8226,N_7464);
or U11485 (N_11485,N_7096,N_7665);
nor U11486 (N_11486,N_6725,N_7322);
nor U11487 (N_11487,N_8356,N_7353);
and U11488 (N_11488,N_7600,N_8714);
nor U11489 (N_11489,N_6142,N_6166);
and U11490 (N_11490,N_8822,N_7752);
nand U11491 (N_11491,N_6821,N_8685);
and U11492 (N_11492,N_7154,N_7738);
and U11493 (N_11493,N_7437,N_7950);
or U11494 (N_11494,N_7499,N_7830);
and U11495 (N_11495,N_8198,N_7901);
nand U11496 (N_11496,N_8831,N_6829);
xor U11497 (N_11497,N_6360,N_8844);
xor U11498 (N_11498,N_7978,N_7990);
and U11499 (N_11499,N_6152,N_8010);
xnor U11500 (N_11500,N_8400,N_8594);
xor U11501 (N_11501,N_8814,N_7897);
nor U11502 (N_11502,N_8922,N_8239);
xor U11503 (N_11503,N_6538,N_6747);
nor U11504 (N_11504,N_6034,N_7364);
or U11505 (N_11505,N_8627,N_6023);
or U11506 (N_11506,N_7044,N_6061);
nor U11507 (N_11507,N_6202,N_8997);
nor U11508 (N_11508,N_8668,N_6089);
nor U11509 (N_11509,N_7407,N_7901);
nor U11510 (N_11510,N_6971,N_8395);
or U11511 (N_11511,N_7897,N_8643);
and U11512 (N_11512,N_7132,N_8510);
xnor U11513 (N_11513,N_6970,N_7758);
xnor U11514 (N_11514,N_6270,N_7659);
xnor U11515 (N_11515,N_6090,N_6287);
and U11516 (N_11516,N_6649,N_7104);
nand U11517 (N_11517,N_7969,N_6403);
nor U11518 (N_11518,N_8933,N_8808);
or U11519 (N_11519,N_8181,N_7250);
and U11520 (N_11520,N_6165,N_8291);
or U11521 (N_11521,N_7642,N_6760);
or U11522 (N_11522,N_6236,N_6037);
or U11523 (N_11523,N_6836,N_7858);
or U11524 (N_11524,N_7844,N_6314);
xor U11525 (N_11525,N_6273,N_6428);
or U11526 (N_11526,N_8304,N_6192);
or U11527 (N_11527,N_6075,N_7835);
nor U11528 (N_11528,N_8081,N_6788);
or U11529 (N_11529,N_8691,N_7558);
and U11530 (N_11530,N_8340,N_7995);
nor U11531 (N_11531,N_7338,N_6254);
xnor U11532 (N_11532,N_8079,N_6689);
nor U11533 (N_11533,N_6316,N_7160);
nor U11534 (N_11534,N_8546,N_6510);
or U11535 (N_11535,N_6338,N_7008);
nor U11536 (N_11536,N_8368,N_8968);
nand U11537 (N_11537,N_7069,N_7445);
and U11538 (N_11538,N_8058,N_7665);
xor U11539 (N_11539,N_8371,N_8049);
xor U11540 (N_11540,N_7037,N_8482);
xor U11541 (N_11541,N_7009,N_6482);
nor U11542 (N_11542,N_8970,N_7442);
xnor U11543 (N_11543,N_6626,N_7062);
or U11544 (N_11544,N_7623,N_6688);
xnor U11545 (N_11545,N_7142,N_6787);
nor U11546 (N_11546,N_7919,N_8481);
xnor U11547 (N_11547,N_7840,N_6436);
and U11548 (N_11548,N_6152,N_7337);
and U11549 (N_11549,N_7102,N_7602);
or U11550 (N_11550,N_7899,N_8145);
nand U11551 (N_11551,N_8603,N_6992);
nor U11552 (N_11552,N_7910,N_7185);
or U11553 (N_11553,N_7040,N_8866);
nand U11554 (N_11554,N_7414,N_8913);
or U11555 (N_11555,N_8957,N_7343);
xor U11556 (N_11556,N_6513,N_6941);
nand U11557 (N_11557,N_7914,N_6321);
xnor U11558 (N_11558,N_6790,N_8720);
xnor U11559 (N_11559,N_6085,N_8065);
nor U11560 (N_11560,N_7706,N_8971);
xor U11561 (N_11561,N_6991,N_7140);
or U11562 (N_11562,N_6687,N_8822);
xor U11563 (N_11563,N_8495,N_8242);
or U11564 (N_11564,N_6158,N_6667);
nand U11565 (N_11565,N_7516,N_6402);
xnor U11566 (N_11566,N_6786,N_6374);
nand U11567 (N_11567,N_7240,N_8637);
or U11568 (N_11568,N_6081,N_7999);
nand U11569 (N_11569,N_8334,N_8176);
nand U11570 (N_11570,N_7758,N_8551);
xor U11571 (N_11571,N_8349,N_7047);
nand U11572 (N_11572,N_7264,N_6338);
or U11573 (N_11573,N_6995,N_8292);
nand U11574 (N_11574,N_6105,N_6520);
xor U11575 (N_11575,N_6673,N_7715);
and U11576 (N_11576,N_7634,N_6681);
nand U11577 (N_11577,N_7100,N_7653);
or U11578 (N_11578,N_6491,N_7588);
and U11579 (N_11579,N_8540,N_8839);
nand U11580 (N_11580,N_8058,N_6599);
nand U11581 (N_11581,N_8741,N_8545);
or U11582 (N_11582,N_8829,N_6126);
or U11583 (N_11583,N_7058,N_7032);
nand U11584 (N_11584,N_7812,N_7848);
nor U11585 (N_11585,N_7362,N_8710);
nand U11586 (N_11586,N_6413,N_6521);
or U11587 (N_11587,N_7141,N_8729);
or U11588 (N_11588,N_7037,N_7241);
or U11589 (N_11589,N_7407,N_6813);
nor U11590 (N_11590,N_7694,N_6862);
and U11591 (N_11591,N_7346,N_6836);
nor U11592 (N_11592,N_7267,N_8828);
and U11593 (N_11593,N_8752,N_8337);
nor U11594 (N_11594,N_7558,N_6760);
nand U11595 (N_11595,N_7777,N_6222);
nand U11596 (N_11596,N_6789,N_7228);
nand U11597 (N_11597,N_8476,N_8243);
nand U11598 (N_11598,N_8762,N_6561);
nand U11599 (N_11599,N_6486,N_8931);
and U11600 (N_11600,N_6935,N_8076);
or U11601 (N_11601,N_6480,N_6111);
nand U11602 (N_11602,N_8866,N_6380);
nor U11603 (N_11603,N_7464,N_8295);
nor U11604 (N_11604,N_7732,N_6674);
xor U11605 (N_11605,N_8573,N_7182);
or U11606 (N_11606,N_6838,N_6408);
and U11607 (N_11607,N_8245,N_7090);
nand U11608 (N_11608,N_7387,N_8486);
nor U11609 (N_11609,N_8001,N_7122);
nand U11610 (N_11610,N_7231,N_8765);
nor U11611 (N_11611,N_6584,N_6055);
nand U11612 (N_11612,N_8252,N_7241);
nor U11613 (N_11613,N_6178,N_6080);
nand U11614 (N_11614,N_7273,N_7878);
or U11615 (N_11615,N_8817,N_8603);
nor U11616 (N_11616,N_7170,N_7184);
and U11617 (N_11617,N_7043,N_7027);
xor U11618 (N_11618,N_8091,N_8679);
nor U11619 (N_11619,N_7606,N_8919);
nor U11620 (N_11620,N_6951,N_7245);
xor U11621 (N_11621,N_6966,N_7296);
and U11622 (N_11622,N_8717,N_6964);
xor U11623 (N_11623,N_8865,N_6391);
or U11624 (N_11624,N_7315,N_7014);
nand U11625 (N_11625,N_7302,N_8897);
nor U11626 (N_11626,N_8207,N_7799);
and U11627 (N_11627,N_6205,N_8341);
and U11628 (N_11628,N_8009,N_8178);
nand U11629 (N_11629,N_8468,N_8287);
nor U11630 (N_11630,N_6438,N_8220);
xor U11631 (N_11631,N_7098,N_7607);
xor U11632 (N_11632,N_8133,N_7773);
and U11633 (N_11633,N_6477,N_7369);
nand U11634 (N_11634,N_7662,N_7527);
or U11635 (N_11635,N_8938,N_6961);
nand U11636 (N_11636,N_8609,N_7854);
nor U11637 (N_11637,N_6377,N_6637);
or U11638 (N_11638,N_8169,N_8545);
and U11639 (N_11639,N_8668,N_8275);
or U11640 (N_11640,N_8040,N_7366);
or U11641 (N_11641,N_6973,N_6224);
xnor U11642 (N_11642,N_6315,N_6881);
nand U11643 (N_11643,N_7037,N_7176);
or U11644 (N_11644,N_6671,N_8450);
nand U11645 (N_11645,N_8715,N_6953);
and U11646 (N_11646,N_7635,N_6036);
or U11647 (N_11647,N_7881,N_7230);
or U11648 (N_11648,N_6722,N_7209);
xnor U11649 (N_11649,N_6295,N_7259);
nor U11650 (N_11650,N_6362,N_7196);
nand U11651 (N_11651,N_6022,N_8667);
nor U11652 (N_11652,N_6463,N_6309);
nand U11653 (N_11653,N_8540,N_8673);
nor U11654 (N_11654,N_8950,N_6794);
and U11655 (N_11655,N_7636,N_7090);
nor U11656 (N_11656,N_7727,N_6981);
xor U11657 (N_11657,N_8082,N_6233);
or U11658 (N_11658,N_8839,N_7149);
or U11659 (N_11659,N_7051,N_7701);
or U11660 (N_11660,N_8841,N_8809);
or U11661 (N_11661,N_6340,N_8269);
xnor U11662 (N_11662,N_6938,N_6358);
or U11663 (N_11663,N_8158,N_7404);
or U11664 (N_11664,N_6010,N_6190);
xor U11665 (N_11665,N_7992,N_7292);
xnor U11666 (N_11666,N_7572,N_8317);
or U11667 (N_11667,N_8746,N_6100);
or U11668 (N_11668,N_6550,N_8182);
xor U11669 (N_11669,N_7300,N_8891);
and U11670 (N_11670,N_6637,N_6834);
and U11671 (N_11671,N_8885,N_7354);
and U11672 (N_11672,N_7420,N_8043);
xnor U11673 (N_11673,N_6541,N_8959);
xor U11674 (N_11674,N_8238,N_7179);
nand U11675 (N_11675,N_7215,N_6058);
nor U11676 (N_11676,N_7694,N_8742);
xor U11677 (N_11677,N_6959,N_8891);
or U11678 (N_11678,N_6116,N_7460);
nand U11679 (N_11679,N_6840,N_8598);
nand U11680 (N_11680,N_7669,N_8915);
and U11681 (N_11681,N_8376,N_7170);
nor U11682 (N_11682,N_8641,N_8842);
or U11683 (N_11683,N_6434,N_7765);
nor U11684 (N_11684,N_7932,N_7686);
and U11685 (N_11685,N_8160,N_8417);
or U11686 (N_11686,N_8365,N_8479);
xnor U11687 (N_11687,N_6590,N_7118);
or U11688 (N_11688,N_7059,N_7746);
nand U11689 (N_11689,N_8759,N_6243);
or U11690 (N_11690,N_7287,N_6891);
nand U11691 (N_11691,N_7607,N_8935);
or U11692 (N_11692,N_7059,N_6375);
or U11693 (N_11693,N_7240,N_6842);
nand U11694 (N_11694,N_8557,N_6025);
nand U11695 (N_11695,N_8396,N_8351);
xor U11696 (N_11696,N_8282,N_6268);
nor U11697 (N_11697,N_6577,N_8110);
nor U11698 (N_11698,N_6396,N_6373);
and U11699 (N_11699,N_8697,N_6673);
nor U11700 (N_11700,N_6450,N_7621);
nand U11701 (N_11701,N_8242,N_6141);
nand U11702 (N_11702,N_6805,N_8566);
and U11703 (N_11703,N_7151,N_8808);
or U11704 (N_11704,N_8217,N_6662);
or U11705 (N_11705,N_8476,N_7260);
nand U11706 (N_11706,N_6869,N_7181);
and U11707 (N_11707,N_7889,N_7676);
and U11708 (N_11708,N_6011,N_7881);
or U11709 (N_11709,N_8274,N_7498);
nor U11710 (N_11710,N_7559,N_6136);
nand U11711 (N_11711,N_7028,N_8168);
nor U11712 (N_11712,N_6064,N_6368);
and U11713 (N_11713,N_8211,N_6724);
xnor U11714 (N_11714,N_8423,N_7303);
xor U11715 (N_11715,N_8737,N_8340);
xnor U11716 (N_11716,N_8115,N_6323);
and U11717 (N_11717,N_8495,N_7197);
or U11718 (N_11718,N_7907,N_7788);
or U11719 (N_11719,N_6289,N_7250);
or U11720 (N_11720,N_7897,N_8802);
and U11721 (N_11721,N_6899,N_7900);
and U11722 (N_11722,N_8381,N_8229);
xor U11723 (N_11723,N_7559,N_6668);
and U11724 (N_11724,N_6879,N_7961);
or U11725 (N_11725,N_7145,N_7717);
nand U11726 (N_11726,N_7043,N_6494);
and U11727 (N_11727,N_8807,N_6043);
nand U11728 (N_11728,N_6391,N_6941);
nor U11729 (N_11729,N_8522,N_6826);
xor U11730 (N_11730,N_7685,N_7995);
or U11731 (N_11731,N_8047,N_8643);
nand U11732 (N_11732,N_8950,N_6733);
xor U11733 (N_11733,N_8627,N_7763);
nand U11734 (N_11734,N_6186,N_8698);
or U11735 (N_11735,N_8674,N_8190);
xnor U11736 (N_11736,N_8573,N_6560);
nor U11737 (N_11737,N_8932,N_6453);
nand U11738 (N_11738,N_6136,N_8205);
nor U11739 (N_11739,N_6887,N_8926);
or U11740 (N_11740,N_8480,N_6587);
and U11741 (N_11741,N_8585,N_7574);
xor U11742 (N_11742,N_8217,N_8095);
xnor U11743 (N_11743,N_7120,N_6326);
xor U11744 (N_11744,N_8540,N_7308);
nand U11745 (N_11745,N_6725,N_8988);
nand U11746 (N_11746,N_8933,N_7878);
nand U11747 (N_11747,N_7810,N_8222);
and U11748 (N_11748,N_7246,N_8601);
xnor U11749 (N_11749,N_8315,N_7465);
nor U11750 (N_11750,N_7055,N_7183);
or U11751 (N_11751,N_7690,N_8332);
xnor U11752 (N_11752,N_6180,N_6884);
and U11753 (N_11753,N_7260,N_6653);
or U11754 (N_11754,N_6980,N_8293);
or U11755 (N_11755,N_8613,N_8802);
nand U11756 (N_11756,N_8553,N_7364);
and U11757 (N_11757,N_6641,N_7565);
and U11758 (N_11758,N_7303,N_6997);
xnor U11759 (N_11759,N_8419,N_7992);
nand U11760 (N_11760,N_6472,N_7259);
nor U11761 (N_11761,N_6012,N_7963);
nor U11762 (N_11762,N_8284,N_7196);
xor U11763 (N_11763,N_7524,N_8451);
and U11764 (N_11764,N_8013,N_7248);
and U11765 (N_11765,N_7438,N_8670);
and U11766 (N_11766,N_6760,N_8535);
and U11767 (N_11767,N_8493,N_8418);
and U11768 (N_11768,N_7008,N_8649);
and U11769 (N_11769,N_8088,N_7205);
nand U11770 (N_11770,N_8944,N_8357);
xor U11771 (N_11771,N_7589,N_7907);
or U11772 (N_11772,N_8389,N_6448);
nand U11773 (N_11773,N_6841,N_7810);
nand U11774 (N_11774,N_8111,N_6085);
nand U11775 (N_11775,N_6912,N_8131);
and U11776 (N_11776,N_7554,N_7969);
xnor U11777 (N_11777,N_7870,N_7059);
or U11778 (N_11778,N_7195,N_8023);
and U11779 (N_11779,N_6506,N_6018);
xnor U11780 (N_11780,N_6279,N_6240);
and U11781 (N_11781,N_6033,N_6704);
nor U11782 (N_11782,N_8191,N_8831);
and U11783 (N_11783,N_6654,N_7659);
nand U11784 (N_11784,N_7204,N_8175);
nor U11785 (N_11785,N_6103,N_8882);
nand U11786 (N_11786,N_6834,N_6377);
or U11787 (N_11787,N_7902,N_7560);
xnor U11788 (N_11788,N_7541,N_6782);
xnor U11789 (N_11789,N_8048,N_8383);
and U11790 (N_11790,N_7966,N_7403);
xor U11791 (N_11791,N_8168,N_8258);
xnor U11792 (N_11792,N_8475,N_6311);
and U11793 (N_11793,N_8149,N_6102);
and U11794 (N_11794,N_7339,N_7251);
or U11795 (N_11795,N_8243,N_6867);
nor U11796 (N_11796,N_8203,N_7235);
xor U11797 (N_11797,N_6017,N_6524);
xnor U11798 (N_11798,N_6239,N_7966);
xnor U11799 (N_11799,N_8230,N_6171);
and U11800 (N_11800,N_8609,N_7680);
and U11801 (N_11801,N_8012,N_8860);
nand U11802 (N_11802,N_6120,N_8633);
nand U11803 (N_11803,N_6413,N_8860);
and U11804 (N_11804,N_6851,N_8846);
and U11805 (N_11805,N_8346,N_8101);
nor U11806 (N_11806,N_7599,N_6652);
and U11807 (N_11807,N_7365,N_6186);
and U11808 (N_11808,N_8224,N_8344);
nor U11809 (N_11809,N_7240,N_7964);
or U11810 (N_11810,N_7996,N_7611);
nand U11811 (N_11811,N_8138,N_6339);
nor U11812 (N_11812,N_6887,N_7219);
nor U11813 (N_11813,N_7857,N_6209);
nor U11814 (N_11814,N_6143,N_7706);
and U11815 (N_11815,N_6784,N_8412);
xor U11816 (N_11816,N_8072,N_6484);
or U11817 (N_11817,N_7350,N_6861);
nor U11818 (N_11818,N_8130,N_8751);
xnor U11819 (N_11819,N_8799,N_8218);
nor U11820 (N_11820,N_6634,N_8860);
nand U11821 (N_11821,N_8029,N_6451);
nor U11822 (N_11822,N_8810,N_6811);
nor U11823 (N_11823,N_7859,N_8817);
xnor U11824 (N_11824,N_7199,N_8836);
and U11825 (N_11825,N_6639,N_6032);
nor U11826 (N_11826,N_6017,N_8393);
nand U11827 (N_11827,N_6665,N_8444);
and U11828 (N_11828,N_6722,N_7324);
nand U11829 (N_11829,N_7482,N_6563);
nand U11830 (N_11830,N_8238,N_8433);
nand U11831 (N_11831,N_7588,N_8355);
or U11832 (N_11832,N_8747,N_7761);
nand U11833 (N_11833,N_8249,N_7384);
xnor U11834 (N_11834,N_7229,N_6708);
nand U11835 (N_11835,N_6872,N_8071);
or U11836 (N_11836,N_8778,N_8402);
and U11837 (N_11837,N_7967,N_8188);
or U11838 (N_11838,N_8717,N_8579);
or U11839 (N_11839,N_6506,N_6686);
and U11840 (N_11840,N_8382,N_6734);
or U11841 (N_11841,N_8422,N_6921);
xnor U11842 (N_11842,N_8638,N_6823);
nand U11843 (N_11843,N_7336,N_8256);
and U11844 (N_11844,N_8268,N_7628);
or U11845 (N_11845,N_8422,N_6610);
and U11846 (N_11846,N_8872,N_6294);
xor U11847 (N_11847,N_8642,N_8907);
nand U11848 (N_11848,N_8402,N_7923);
nand U11849 (N_11849,N_6771,N_8304);
or U11850 (N_11850,N_7928,N_7192);
and U11851 (N_11851,N_8785,N_6641);
or U11852 (N_11852,N_6773,N_7057);
nand U11853 (N_11853,N_8858,N_7360);
and U11854 (N_11854,N_7618,N_7955);
or U11855 (N_11855,N_7390,N_7332);
and U11856 (N_11856,N_8056,N_7132);
nand U11857 (N_11857,N_6948,N_8409);
nand U11858 (N_11858,N_8621,N_8932);
or U11859 (N_11859,N_8022,N_6557);
xor U11860 (N_11860,N_7021,N_8533);
nand U11861 (N_11861,N_7687,N_6561);
and U11862 (N_11862,N_6329,N_8789);
xnor U11863 (N_11863,N_6315,N_8402);
nand U11864 (N_11864,N_8327,N_7118);
or U11865 (N_11865,N_6345,N_8705);
or U11866 (N_11866,N_6439,N_8329);
or U11867 (N_11867,N_6238,N_8655);
or U11868 (N_11868,N_8357,N_7196);
or U11869 (N_11869,N_8455,N_7726);
nor U11870 (N_11870,N_6705,N_8428);
and U11871 (N_11871,N_8988,N_8368);
xor U11872 (N_11872,N_7591,N_7174);
nor U11873 (N_11873,N_8188,N_7137);
or U11874 (N_11874,N_7316,N_7259);
xor U11875 (N_11875,N_6546,N_6739);
and U11876 (N_11876,N_6827,N_8713);
or U11877 (N_11877,N_6647,N_8770);
nand U11878 (N_11878,N_7693,N_8811);
nor U11879 (N_11879,N_6723,N_7936);
or U11880 (N_11880,N_6455,N_7436);
or U11881 (N_11881,N_7403,N_8146);
nand U11882 (N_11882,N_7533,N_6295);
nand U11883 (N_11883,N_6536,N_7586);
xnor U11884 (N_11884,N_6844,N_8387);
nor U11885 (N_11885,N_8531,N_6791);
nand U11886 (N_11886,N_6800,N_7199);
xor U11887 (N_11887,N_7073,N_6028);
and U11888 (N_11888,N_8814,N_8248);
and U11889 (N_11889,N_8786,N_7994);
nor U11890 (N_11890,N_6941,N_6893);
xor U11891 (N_11891,N_8777,N_8362);
or U11892 (N_11892,N_8777,N_8949);
nor U11893 (N_11893,N_7238,N_7968);
and U11894 (N_11894,N_8800,N_8020);
xnor U11895 (N_11895,N_6295,N_6301);
and U11896 (N_11896,N_8104,N_7099);
and U11897 (N_11897,N_8141,N_6855);
or U11898 (N_11898,N_6330,N_6254);
or U11899 (N_11899,N_8468,N_8465);
nand U11900 (N_11900,N_7044,N_6229);
or U11901 (N_11901,N_8329,N_7716);
xor U11902 (N_11902,N_6118,N_6919);
nand U11903 (N_11903,N_7229,N_8120);
nor U11904 (N_11904,N_7532,N_8322);
xor U11905 (N_11905,N_7335,N_8926);
nor U11906 (N_11906,N_7444,N_7584);
xor U11907 (N_11907,N_7878,N_6842);
nand U11908 (N_11908,N_7690,N_8804);
or U11909 (N_11909,N_7433,N_7122);
or U11910 (N_11910,N_8150,N_6549);
and U11911 (N_11911,N_7506,N_8321);
or U11912 (N_11912,N_8641,N_8572);
nor U11913 (N_11913,N_7374,N_6394);
xnor U11914 (N_11914,N_7072,N_7952);
and U11915 (N_11915,N_8722,N_7127);
nand U11916 (N_11916,N_7297,N_6156);
xnor U11917 (N_11917,N_8087,N_7693);
xor U11918 (N_11918,N_6735,N_8129);
nor U11919 (N_11919,N_7434,N_6469);
nor U11920 (N_11920,N_8311,N_8927);
nor U11921 (N_11921,N_7258,N_8028);
xor U11922 (N_11922,N_7689,N_7039);
xnor U11923 (N_11923,N_6491,N_7759);
or U11924 (N_11924,N_8608,N_6050);
nor U11925 (N_11925,N_8882,N_7264);
and U11926 (N_11926,N_8889,N_7630);
nor U11927 (N_11927,N_6219,N_7274);
xor U11928 (N_11928,N_7864,N_8342);
or U11929 (N_11929,N_6336,N_6528);
nor U11930 (N_11930,N_8529,N_8343);
or U11931 (N_11931,N_6753,N_6196);
nor U11932 (N_11932,N_8930,N_7616);
xnor U11933 (N_11933,N_6852,N_8687);
xor U11934 (N_11934,N_8483,N_7650);
or U11935 (N_11935,N_6288,N_8574);
or U11936 (N_11936,N_7319,N_7991);
and U11937 (N_11937,N_7763,N_8303);
or U11938 (N_11938,N_6215,N_7086);
or U11939 (N_11939,N_6845,N_7866);
and U11940 (N_11940,N_7495,N_7089);
or U11941 (N_11941,N_7651,N_6416);
nor U11942 (N_11942,N_8795,N_8389);
xnor U11943 (N_11943,N_7234,N_7570);
xnor U11944 (N_11944,N_7475,N_8934);
nand U11945 (N_11945,N_8945,N_6505);
nor U11946 (N_11946,N_8224,N_7820);
nand U11947 (N_11947,N_8926,N_7121);
nand U11948 (N_11948,N_8722,N_8261);
nand U11949 (N_11949,N_6905,N_7215);
nor U11950 (N_11950,N_6969,N_7997);
or U11951 (N_11951,N_7252,N_6817);
or U11952 (N_11952,N_7785,N_8184);
and U11953 (N_11953,N_8199,N_7076);
xnor U11954 (N_11954,N_8116,N_8261);
xnor U11955 (N_11955,N_7983,N_7367);
nor U11956 (N_11956,N_8084,N_8333);
nor U11957 (N_11957,N_6553,N_7288);
or U11958 (N_11958,N_7536,N_8933);
xnor U11959 (N_11959,N_8053,N_7939);
nand U11960 (N_11960,N_8640,N_7759);
xnor U11961 (N_11961,N_7844,N_7054);
and U11962 (N_11962,N_6629,N_7240);
nand U11963 (N_11963,N_8914,N_7834);
xnor U11964 (N_11964,N_8887,N_8230);
and U11965 (N_11965,N_8973,N_6924);
nand U11966 (N_11966,N_8869,N_7213);
nor U11967 (N_11967,N_7023,N_6704);
nand U11968 (N_11968,N_6678,N_8331);
nand U11969 (N_11969,N_8996,N_7087);
nand U11970 (N_11970,N_8267,N_8829);
nand U11971 (N_11971,N_6192,N_7802);
nand U11972 (N_11972,N_6005,N_7623);
and U11973 (N_11973,N_6925,N_6207);
xor U11974 (N_11974,N_7086,N_7433);
nor U11975 (N_11975,N_6277,N_6145);
xor U11976 (N_11976,N_7128,N_8070);
or U11977 (N_11977,N_8862,N_7708);
nand U11978 (N_11978,N_7995,N_8642);
xnor U11979 (N_11979,N_6923,N_8264);
nor U11980 (N_11980,N_8818,N_7349);
and U11981 (N_11981,N_8277,N_6275);
or U11982 (N_11982,N_6005,N_7776);
nand U11983 (N_11983,N_7795,N_6899);
nor U11984 (N_11984,N_6039,N_6607);
and U11985 (N_11985,N_6643,N_6285);
nor U11986 (N_11986,N_7321,N_8043);
nand U11987 (N_11987,N_6153,N_8043);
nand U11988 (N_11988,N_6648,N_7103);
xor U11989 (N_11989,N_8128,N_6694);
nor U11990 (N_11990,N_7970,N_7608);
nand U11991 (N_11991,N_6785,N_8904);
nand U11992 (N_11992,N_6313,N_8006);
xnor U11993 (N_11993,N_8200,N_8504);
xor U11994 (N_11994,N_7898,N_8661);
or U11995 (N_11995,N_8218,N_6801);
or U11996 (N_11996,N_7239,N_8160);
nand U11997 (N_11997,N_6313,N_7135);
nand U11998 (N_11998,N_6890,N_6716);
or U11999 (N_11999,N_7193,N_8697);
and U12000 (N_12000,N_9953,N_11731);
nand U12001 (N_12001,N_11930,N_10139);
nor U12002 (N_12002,N_9656,N_9360);
nor U12003 (N_12003,N_10142,N_10656);
nor U12004 (N_12004,N_11815,N_10507);
and U12005 (N_12005,N_9281,N_11092);
xor U12006 (N_12006,N_11929,N_9423);
nand U12007 (N_12007,N_11106,N_10104);
xor U12008 (N_12008,N_10683,N_9615);
xor U12009 (N_12009,N_11486,N_11042);
and U12010 (N_12010,N_10266,N_9301);
or U12011 (N_12011,N_10216,N_11728);
nor U12012 (N_12012,N_11420,N_10382);
nand U12013 (N_12013,N_9456,N_11666);
xor U12014 (N_12014,N_10843,N_10990);
or U12015 (N_12015,N_9106,N_11889);
xnor U12016 (N_12016,N_9708,N_9262);
xnor U12017 (N_12017,N_9088,N_9922);
xor U12018 (N_12018,N_9357,N_10762);
nor U12019 (N_12019,N_11047,N_9839);
nand U12020 (N_12020,N_10998,N_11747);
nor U12021 (N_12021,N_10985,N_10178);
nor U12022 (N_12022,N_9529,N_11090);
or U12023 (N_12023,N_11248,N_9381);
nand U12024 (N_12024,N_11607,N_11387);
or U12025 (N_12025,N_10637,N_9745);
or U12026 (N_12026,N_9721,N_9532);
nand U12027 (N_12027,N_9134,N_10514);
or U12028 (N_12028,N_11934,N_9858);
xnor U12029 (N_12029,N_9407,N_9069);
xnor U12030 (N_12030,N_10007,N_10112);
xnor U12031 (N_12031,N_11292,N_9831);
nor U12032 (N_12032,N_10881,N_10156);
nand U12033 (N_12033,N_10176,N_10483);
nand U12034 (N_12034,N_9097,N_11300);
xnor U12035 (N_12035,N_11673,N_9189);
xor U12036 (N_12036,N_11215,N_10133);
and U12037 (N_12037,N_9994,N_10753);
and U12038 (N_12038,N_9062,N_10123);
xnor U12039 (N_12039,N_9011,N_9022);
nand U12040 (N_12040,N_9241,N_11743);
or U12041 (N_12041,N_10220,N_9180);
nand U12042 (N_12042,N_10891,N_11030);
or U12043 (N_12043,N_10935,N_10061);
or U12044 (N_12044,N_10287,N_9815);
xnor U12045 (N_12045,N_9494,N_10849);
nor U12046 (N_12046,N_9890,N_11640);
nand U12047 (N_12047,N_9130,N_9761);
nor U12048 (N_12048,N_9206,N_10475);
nand U12049 (N_12049,N_11327,N_9782);
and U12050 (N_12050,N_9386,N_11115);
nand U12051 (N_12051,N_11739,N_10513);
nand U12052 (N_12052,N_11288,N_10032);
and U12053 (N_12053,N_10413,N_11459);
xnor U12054 (N_12054,N_9557,N_10207);
and U12055 (N_12055,N_11928,N_9682);
xnor U12056 (N_12056,N_11391,N_11571);
xnor U12057 (N_12057,N_10542,N_11053);
or U12058 (N_12058,N_9989,N_9033);
nor U12059 (N_12059,N_10950,N_10294);
xor U12060 (N_12060,N_9499,N_9065);
and U12061 (N_12061,N_10960,N_9050);
nand U12062 (N_12062,N_11500,N_10244);
xnor U12063 (N_12063,N_9644,N_9693);
nor U12064 (N_12064,N_10400,N_9163);
and U12065 (N_12065,N_9982,N_10047);
nand U12066 (N_12066,N_9034,N_11901);
or U12067 (N_12067,N_10128,N_11503);
nor U12068 (N_12068,N_10141,N_10800);
xnor U12069 (N_12069,N_10798,N_9877);
or U12070 (N_12070,N_11455,N_11360);
nor U12071 (N_12071,N_9916,N_10505);
nor U12072 (N_12072,N_11179,N_11907);
and U12073 (N_12073,N_9412,N_9370);
and U12074 (N_12074,N_9049,N_9201);
nor U12075 (N_12075,N_11301,N_11644);
nor U12076 (N_12076,N_9710,N_9876);
nor U12077 (N_12077,N_9125,N_11809);
or U12078 (N_12078,N_10841,N_9430);
or U12079 (N_12079,N_10541,N_10395);
and U12080 (N_12080,N_9726,N_11104);
and U12081 (N_12081,N_10968,N_9236);
nand U12082 (N_12082,N_9283,N_9316);
nor U12083 (N_12083,N_10371,N_11043);
or U12084 (N_12084,N_11745,N_10770);
or U12085 (N_12085,N_11594,N_9739);
nand U12086 (N_12086,N_11433,N_9508);
or U12087 (N_12087,N_9764,N_9903);
xor U12088 (N_12088,N_9152,N_10684);
or U12089 (N_12089,N_10794,N_10408);
and U12090 (N_12090,N_11130,N_10097);
nand U12091 (N_12091,N_11583,N_9830);
and U12092 (N_12092,N_10587,N_11397);
or U12093 (N_12093,N_10717,N_10819);
and U12094 (N_12094,N_11177,N_10042);
and U12095 (N_12095,N_9136,N_9471);
nand U12096 (N_12096,N_10389,N_9632);
nand U12097 (N_12097,N_9600,N_11938);
xor U12098 (N_12098,N_9758,N_9148);
nor U12099 (N_12099,N_9238,N_9874);
nand U12100 (N_12100,N_11997,N_10987);
nor U12101 (N_12101,N_9377,N_9649);
nand U12102 (N_12102,N_11328,N_11176);
nand U12103 (N_12103,N_10706,N_9829);
xnor U12104 (N_12104,N_10902,N_10373);
or U12105 (N_12105,N_11409,N_10551);
and U12106 (N_12106,N_9822,N_9654);
xnor U12107 (N_12107,N_9610,N_10461);
xnor U12108 (N_12108,N_9611,N_9379);
or U12109 (N_12109,N_9707,N_9571);
and U12110 (N_12110,N_11544,N_9437);
nor U12111 (N_12111,N_10642,N_11089);
nand U12112 (N_12112,N_11237,N_9017);
nand U12113 (N_12113,N_11070,N_10401);
xnor U12114 (N_12114,N_10409,N_9119);
xor U12115 (N_12115,N_10729,N_9185);
nor U12116 (N_12116,N_9555,N_9567);
xor U12117 (N_12117,N_9742,N_9757);
nand U12118 (N_12118,N_11556,N_9438);
or U12119 (N_12119,N_11192,N_9135);
or U12120 (N_12120,N_9162,N_9326);
nand U12121 (N_12121,N_11977,N_9419);
or U12122 (N_12122,N_10643,N_9380);
or U12123 (N_12123,N_10057,N_11353);
xnor U12124 (N_12124,N_11765,N_10058);
xnor U12125 (N_12125,N_9302,N_10816);
and U12126 (N_12126,N_10585,N_9123);
nand U12127 (N_12127,N_9714,N_9900);
and U12128 (N_12128,N_10926,N_10438);
nand U12129 (N_12129,N_11001,N_10424);
and U12130 (N_12130,N_9875,N_10808);
xnor U12131 (N_12131,N_9473,N_11870);
or U12132 (N_12132,N_9513,N_9428);
nand U12133 (N_12133,N_9651,N_11474);
xor U12134 (N_12134,N_9199,N_9952);
and U12135 (N_12135,N_11851,N_10972);
nand U12136 (N_12136,N_10658,N_9399);
or U12137 (N_12137,N_11082,N_11592);
xnor U12138 (N_12138,N_9333,N_10282);
and U12139 (N_12139,N_9595,N_10783);
xnor U12140 (N_12140,N_11406,N_9368);
xnor U12141 (N_12141,N_10710,N_11156);
and U12142 (N_12142,N_9583,N_10013);
nor U12143 (N_12143,N_11533,N_9871);
or U12144 (N_12144,N_11316,N_11935);
nor U12145 (N_12145,N_9814,N_11314);
and U12146 (N_12146,N_11591,N_9848);
nor U12147 (N_12147,N_11603,N_9717);
nor U12148 (N_12148,N_11998,N_11504);
or U12149 (N_12149,N_10928,N_10666);
or U12150 (N_12150,N_9582,N_11820);
and U12151 (N_12151,N_11638,N_9638);
or U12152 (N_12152,N_9665,N_10189);
nand U12153 (N_12153,N_11780,N_10754);
xnor U12154 (N_12154,N_11627,N_11491);
or U12155 (N_12155,N_9784,N_10495);
nand U12156 (N_12156,N_9663,N_11676);
xor U12157 (N_12157,N_11036,N_11727);
nor U12158 (N_12158,N_9558,N_11808);
nor U12159 (N_12159,N_9292,N_9608);
xnor U12160 (N_12160,N_9970,N_9934);
nand U12161 (N_12161,N_9156,N_10246);
or U12162 (N_12162,N_11402,N_9124);
nand U12163 (N_12163,N_9285,N_11847);
or U12164 (N_12164,N_10386,N_11733);
nand U12165 (N_12165,N_10259,N_9564);
nand U12166 (N_12166,N_9165,N_9451);
and U12167 (N_12167,N_11094,N_10027);
or U12168 (N_12168,N_10700,N_9485);
nand U12169 (N_12169,N_10722,N_10325);
xor U12170 (N_12170,N_10309,N_9841);
xnor U12171 (N_12171,N_9008,N_11667);
and U12172 (N_12172,N_9418,N_10043);
and U12173 (N_12173,N_9853,N_9643);
nor U12174 (N_12174,N_10641,N_10268);
nor U12175 (N_12175,N_11554,N_11172);
or U12176 (N_12176,N_11134,N_10512);
or U12177 (N_12177,N_11857,N_9237);
nor U12178 (N_12178,N_10975,N_9070);
or U12179 (N_12179,N_10035,N_11493);
nor U12180 (N_12180,N_11333,N_9667);
and U12181 (N_12181,N_10344,N_11978);
nand U12182 (N_12182,N_11914,N_10749);
xor U12183 (N_12183,N_9342,N_10671);
nor U12184 (N_12184,N_11118,N_9927);
and U12185 (N_12185,N_10117,N_11688);
nor U12186 (N_12186,N_9932,N_11983);
and U12187 (N_12187,N_11032,N_11212);
xnor U12188 (N_12188,N_10883,N_9224);
xor U12189 (N_12189,N_10872,N_11273);
or U12190 (N_12190,N_11852,N_10225);
nor U12191 (N_12191,N_9552,N_10138);
nor U12192 (N_12192,N_10378,N_10354);
nor U12193 (N_12193,N_11611,N_11700);
nor U12194 (N_12194,N_9480,N_10267);
and U12195 (N_12195,N_10312,N_10605);
nor U12196 (N_12196,N_10876,N_10110);
and U12197 (N_12197,N_10162,N_9700);
and U12198 (N_12198,N_10357,N_10126);
xnor U12199 (N_12199,N_10965,N_11169);
and U12200 (N_12200,N_11034,N_11323);
nand U12201 (N_12201,N_11136,N_11757);
and U12202 (N_12202,N_9099,N_11752);
or U12203 (N_12203,N_9543,N_10989);
xor U12204 (N_12204,N_10191,N_10233);
xor U12205 (N_12205,N_10650,N_11494);
nor U12206 (N_12206,N_11012,N_9760);
nand U12207 (N_12207,N_10780,N_10101);
nand U12208 (N_12208,N_9012,N_10583);
and U12209 (N_12209,N_9751,N_10860);
xnor U12210 (N_12210,N_9335,N_11619);
nand U12211 (N_12211,N_10439,N_9636);
nor U12212 (N_12212,N_10687,N_9055);
nand U12213 (N_12213,N_10689,N_10861);
nand U12214 (N_12214,N_11654,N_10611);
nor U12215 (N_12215,N_9196,N_10918);
nand U12216 (N_12216,N_10537,N_9730);
nand U12217 (N_12217,N_10526,N_11916);
or U12218 (N_12218,N_11536,N_11581);
nor U12219 (N_12219,N_10554,N_9735);
and U12220 (N_12220,N_10326,N_10823);
or U12221 (N_12221,N_10565,N_11840);
xor U12222 (N_12222,N_11343,N_10547);
xor U12223 (N_12223,N_9773,N_11223);
nand U12224 (N_12224,N_11527,N_10221);
nand U12225 (N_12225,N_11324,N_10202);
nand U12226 (N_12226,N_11797,N_9867);
or U12227 (N_12227,N_10083,N_9299);
and U12228 (N_12228,N_9104,N_9074);
xnor U12229 (N_12229,N_9043,N_10634);
or U12230 (N_12230,N_9391,N_9198);
or U12231 (N_12231,N_9512,N_11650);
xnor U12232 (N_12232,N_10925,N_10295);
nor U12233 (N_12233,N_11810,N_9576);
nor U12234 (N_12234,N_11423,N_10305);
and U12235 (N_12235,N_9680,N_9396);
and U12236 (N_12236,N_11199,N_10290);
nor U12237 (N_12237,N_11606,N_9996);
xnor U12238 (N_12238,N_9117,N_11718);
nand U12239 (N_12239,N_11959,N_9704);
xor U12240 (N_12240,N_11233,N_11087);
and U12241 (N_12241,N_10827,N_10089);
or U12242 (N_12242,N_10580,N_10517);
or U12243 (N_12243,N_10329,N_10405);
nor U12244 (N_12244,N_11129,N_9790);
xor U12245 (N_12245,N_11120,N_10361);
nand U12246 (N_12246,N_10053,N_11194);
nand U12247 (N_12247,N_11871,N_10343);
nand U12248 (N_12248,N_11645,N_10346);
nor U12249 (N_12249,N_9898,N_9369);
and U12250 (N_12250,N_11488,N_9039);
nor U12251 (N_12251,N_9294,N_10919);
nand U12252 (N_12252,N_11828,N_11767);
or U12253 (N_12253,N_11738,N_9015);
nand U12254 (N_12254,N_11213,N_9936);
xor U12255 (N_12255,N_10060,N_11970);
and U12256 (N_12256,N_11252,N_11967);
nand U12257 (N_12257,N_10723,N_11944);
or U12258 (N_12258,N_9647,N_9270);
nand U12259 (N_12259,N_9716,N_11760);
nand U12260 (N_12260,N_9140,N_10579);
nor U12261 (N_12261,N_9881,N_10468);
or U12262 (N_12262,N_9109,N_11270);
nand U12263 (N_12263,N_10536,N_11593);
xnor U12264 (N_12264,N_11203,N_9631);
nand U12265 (N_12265,N_10492,N_10278);
nor U12266 (N_12266,N_9635,N_11175);
and U12267 (N_12267,N_10734,N_10592);
nand U12268 (N_12268,N_11943,N_10347);
nor U12269 (N_12269,N_11712,N_9242);
and U12270 (N_12270,N_9247,N_10167);
nand U12271 (N_12271,N_9942,N_11263);
xnor U12272 (N_12272,N_9550,N_9303);
nor U12273 (N_12273,N_9882,N_10261);
and U12274 (N_12274,N_10423,N_10168);
nand U12275 (N_12275,N_10694,N_11547);
nand U12276 (N_12276,N_9522,N_10486);
nand U12277 (N_12277,N_10721,N_10442);
and U12278 (N_12278,N_10310,N_9448);
nand U12279 (N_12279,N_10429,N_10855);
nor U12280 (N_12280,N_10769,N_11296);
nand U12281 (N_12281,N_10792,N_11009);
xnor U12282 (N_12282,N_9265,N_11528);
and U12283 (N_12283,N_10284,N_11874);
and U12284 (N_12284,N_11584,N_11447);
xor U12285 (N_12285,N_10118,N_9534);
nand U12286 (N_12286,N_10021,N_9094);
nand U12287 (N_12287,N_10399,N_10654);
xnor U12288 (N_12288,N_10606,N_11701);
nor U12289 (N_12289,N_11643,N_11799);
and U12290 (N_12290,N_10328,N_11099);
or U12291 (N_12291,N_10196,N_11144);
and U12292 (N_12292,N_9346,N_10504);
nor U12293 (N_12293,N_9037,N_11677);
or U12294 (N_12294,N_9010,N_11893);
or U12295 (N_12295,N_10915,N_10655);
xnor U12296 (N_12296,N_11601,N_9744);
nor U12297 (N_12297,N_9483,N_9873);
and U12298 (N_12298,N_11839,N_9112);
nand U12299 (N_12299,N_9239,N_11431);
nand U12300 (N_12300,N_9071,N_11011);
and U12301 (N_12301,N_11347,N_10669);
nor U12302 (N_12302,N_9523,N_11329);
and U12303 (N_12303,N_10835,N_11499);
nor U12304 (N_12304,N_9808,N_9068);
xor U12305 (N_12305,N_10066,N_10924);
or U12306 (N_12306,N_10612,N_11853);
or U12307 (N_12307,N_10306,N_9753);
xnor U12308 (N_12308,N_11095,N_11725);
nand U12309 (N_12309,N_9329,N_11740);
nor U12310 (N_12310,N_10766,N_11662);
or U12311 (N_12311,N_9306,N_9233);
xor U12312 (N_12312,N_11386,N_11999);
xnor U12313 (N_12313,N_9161,N_10015);
or U12314 (N_12314,N_9249,N_9689);
or U12315 (N_12315,N_10026,N_10622);
or U12316 (N_12316,N_9819,N_11456);
nand U12317 (N_12317,N_9535,N_10488);
nand U12318 (N_12318,N_10456,N_9031);
nand U12319 (N_12319,N_11816,N_9215);
or U12320 (N_12320,N_11990,N_9332);
and U12321 (N_12321,N_11846,N_10943);
and U12322 (N_12322,N_11838,N_9536);
or U12323 (N_12323,N_11251,N_9517);
nor U12324 (N_12324,N_9177,N_9435);
or U12325 (N_12325,N_11337,N_10624);
or U12326 (N_12326,N_11180,N_11201);
and U12327 (N_12327,N_9669,N_11514);
nor U12328 (N_12328,N_9221,N_11649);
or U12329 (N_12329,N_9016,N_9063);
and U12330 (N_12330,N_10847,N_10828);
nor U12331 (N_12331,N_10750,N_10231);
or U12332 (N_12332,N_11535,N_11171);
and U12333 (N_12333,N_9209,N_11523);
xnor U12334 (N_12334,N_11559,N_10130);
and U12335 (N_12335,N_10010,N_11784);
xor U12336 (N_12336,N_11579,N_11404);
and U12337 (N_12337,N_11417,N_9677);
xor U12338 (N_12338,N_9083,N_10252);
and U12339 (N_12339,N_11257,N_11680);
or U12340 (N_12340,N_11265,N_9843);
nor U12341 (N_12341,N_9105,N_11598);
xnor U12342 (N_12342,N_11778,N_9759);
nor U12343 (N_12343,N_9729,N_9304);
or U12344 (N_12344,N_9780,N_10175);
or U12345 (N_12345,N_9400,N_11150);
nor U12346 (N_12346,N_9311,N_11102);
xnor U12347 (N_12347,N_9317,N_11178);
nor U12348 (N_12348,N_9637,N_10736);
nand U12349 (N_12349,N_11415,N_9405);
and U12350 (N_12350,N_9268,N_11256);
nand U12351 (N_12351,N_9639,N_10147);
nand U12352 (N_12352,N_10498,N_11278);
or U12353 (N_12353,N_11232,N_9443);
xor U12354 (N_12354,N_9577,N_11985);
and U12355 (N_12355,N_9051,N_9849);
or U12356 (N_12356,N_10795,N_9911);
nor U12357 (N_12357,N_9254,N_10867);
nand U12358 (N_12358,N_10682,N_11735);
and U12359 (N_12359,N_10374,N_10377);
and U12360 (N_12360,N_9336,N_9493);
xnor U12361 (N_12361,N_10834,N_10550);
and U12362 (N_12362,N_9089,N_9339);
nand U12363 (N_12363,N_9314,N_9851);
and U12364 (N_12364,N_9981,N_11989);
and U12365 (N_12365,N_9913,N_9605);
nand U12366 (N_12366,N_11621,N_10359);
or U12367 (N_12367,N_9439,N_9279);
xnor U12368 (N_12368,N_11298,N_11127);
nand U12369 (N_12369,N_10745,N_9211);
nor U12370 (N_12370,N_10190,N_11147);
nor U12371 (N_12371,N_9059,N_11158);
xor U12372 (N_12372,N_11345,N_10815);
xnor U12373 (N_12373,N_11761,N_11910);
xor U12374 (N_12374,N_10920,N_10322);
or U12375 (N_12375,N_11195,N_10760);
and U12376 (N_12376,N_9417,N_11793);
nand U12377 (N_12377,N_9171,N_10791);
nor U12378 (N_12378,N_10064,N_10940);
or U12379 (N_12379,N_11358,N_11413);
or U12380 (N_12380,N_11939,N_9793);
xor U12381 (N_12381,N_11782,N_11966);
or U12382 (N_12382,N_10124,N_9155);
and U12383 (N_12383,N_10255,N_11860);
and U12384 (N_12384,N_9521,N_9628);
and U12385 (N_12385,N_9698,N_10148);
xnor U12386 (N_12386,N_11585,N_9277);
or U12387 (N_12387,N_9118,N_9991);
and U12388 (N_12388,N_9406,N_10292);
nor U12389 (N_12389,N_11575,N_10997);
and U12390 (N_12390,N_9949,N_9393);
nand U12391 (N_12391,N_10906,N_10398);
nor U12392 (N_12392,N_9328,N_11497);
or U12393 (N_12393,N_10434,N_11240);
nand U12394 (N_12394,N_9217,N_10983);
nor U12395 (N_12395,N_11900,N_11421);
and U12396 (N_12396,N_9694,N_11121);
nand U12397 (N_12397,N_11781,N_11408);
and U12398 (N_12398,N_10868,N_9115);
or U12399 (N_12399,N_11084,N_9574);
and U12400 (N_12400,N_11786,N_10994);
nand U12401 (N_12401,N_11165,N_11798);
nand U12402 (N_12402,N_10562,N_11390);
and U12403 (N_12403,N_9581,N_9432);
or U12404 (N_12404,N_9044,N_10185);
xor U12405 (N_12405,N_11000,N_9640);
xnor U12406 (N_12406,N_10115,N_9609);
or U12407 (N_12407,N_11691,N_11365);
or U12408 (N_12408,N_10857,N_9786);
nor U12409 (N_12409,N_9347,N_11689);
xnor U12410 (N_12410,N_11166,N_10071);
xnor U12411 (N_12411,N_9081,N_10822);
and U12412 (N_12412,N_10809,N_9754);
nand U12413 (N_12413,N_9695,N_11829);
nand U12414 (N_12414,N_9442,N_10446);
or U12415 (N_12415,N_10376,N_9601);
xnor U12416 (N_12416,N_10515,N_11429);
nor U12417 (N_12417,N_11716,N_9652);
or U12418 (N_12418,N_9052,N_10738);
or U12419 (N_12419,N_9359,N_10052);
nor U12420 (N_12420,N_9169,N_10971);
nor U12421 (N_12421,N_11453,N_11438);
nand U12422 (N_12422,N_10151,N_9559);
or U12423 (N_12423,N_10356,N_9617);
xor U12424 (N_12424,N_10113,N_10544);
nand U12425 (N_12425,N_10991,N_11382);
or U12426 (N_12426,N_10197,N_9110);
nand U12427 (N_12427,N_9907,N_11200);
nand U12428 (N_12428,N_10023,N_11416);
xor U12429 (N_12429,N_10237,N_9312);
and U12430 (N_12430,N_10977,N_9519);
nand U12431 (N_12431,N_9572,N_9972);
nor U12432 (N_12432,N_11373,N_10132);
nor U12433 (N_12433,N_11831,N_11219);
nor U12434 (N_12434,N_10680,N_10457);
nand U12435 (N_12435,N_11018,N_11612);
nand U12436 (N_12436,N_10856,N_10672);
xor U12437 (N_12437,N_11834,N_9382);
or U12438 (N_12438,N_9846,N_11708);
nor U12439 (N_12439,N_9706,N_10892);
xor U12440 (N_12440,N_10315,N_10836);
xnor U12441 (N_12441,N_11958,N_10516);
nor U12442 (N_12442,N_9046,N_11792);
xnor U12443 (N_12443,N_11508,N_9421);
and U12444 (N_12444,N_9193,N_11440);
nand U12445 (N_12445,N_11015,N_11330);
nor U12446 (N_12446,N_11813,N_9928);
and U12447 (N_12447,N_11885,N_9768);
nand U12448 (N_12448,N_10718,N_10180);
nor U12449 (N_12449,N_10392,N_9959);
nand U12450 (N_12450,N_11254,N_10239);
or U12451 (N_12451,N_10415,N_9309);
nand U12452 (N_12452,N_11568,N_11833);
nand U12453 (N_12453,N_11126,N_11430);
or U12454 (N_12454,N_11204,N_10615);
xnor U12455 (N_12455,N_11564,N_11191);
xnor U12456 (N_12456,N_11826,N_10609);
nand U12457 (N_12457,N_10910,N_9660);
or U12458 (N_12458,N_11231,N_11529);
xor U12459 (N_12459,N_9666,N_9018);
or U12460 (N_12460,N_10430,N_9461);
xnor U12461 (N_12461,N_9733,N_10789);
nor U12462 (N_12462,N_11470,N_11209);
nand U12463 (N_12463,N_11214,N_10119);
nor U12464 (N_12464,N_9859,N_11613);
and U12465 (N_12465,N_11538,N_9533);
nand U12466 (N_12466,N_9833,N_9496);
nand U12467 (N_12467,N_11891,N_9240);
nand U12468 (N_12468,N_9527,N_11899);
and U12469 (N_12469,N_9073,N_9232);
nor U12470 (N_12470,N_10081,N_11908);
nor U12471 (N_12471,N_9894,N_10358);
nor U12472 (N_12472,N_9202,N_11909);
nor U12473 (N_12473,N_10425,N_10570);
nand U12474 (N_12474,N_11884,N_9918);
nand U12475 (N_12475,N_11143,N_11626);
or U12476 (N_12476,N_10257,N_11850);
and U12477 (N_12477,N_9672,N_9133);
nand U12478 (N_12478,N_11044,N_10801);
nand U12479 (N_12479,N_10209,N_9434);
and U12480 (N_12480,N_10603,N_9072);
and U12481 (N_12481,N_11291,N_11507);
nor U12482 (N_12482,N_10630,N_11887);
nand U12483 (N_12483,N_9464,N_10201);
and U12484 (N_12484,N_11450,N_10556);
and U12485 (N_12485,N_9093,N_10787);
or U12486 (N_12486,N_10441,N_9818);
and U12487 (N_12487,N_10616,N_10187);
or U12488 (N_12488,N_11525,N_11867);
nor U12489 (N_12489,N_11849,N_9899);
xnor U12490 (N_12490,N_10705,N_10355);
xor U12491 (N_12491,N_11753,N_11294);
and U12492 (N_12492,N_10059,N_10804);
nor U12493 (N_12493,N_11974,N_10796);
and U12494 (N_12494,N_9910,N_11803);
xnor U12495 (N_12495,N_10519,N_11726);
nor U12496 (N_12496,N_11790,N_9766);
xnor U12497 (N_12497,N_10317,N_11091);
or U12498 (N_12498,N_9909,N_9348);
nand U12499 (N_12499,N_11374,N_11577);
nand U12500 (N_12500,N_11751,N_10489);
or U12501 (N_12501,N_9486,N_9957);
or U12502 (N_12502,N_10487,N_11618);
or U12503 (N_12503,N_11141,N_10280);
nor U12504 (N_12504,N_9426,N_9560);
or U12505 (N_12505,N_11542,N_9884);
or U12506 (N_12506,N_10125,N_11196);
and U12507 (N_12507,N_9474,N_11925);
nor U12508 (N_12508,N_10170,N_10470);
and U12509 (N_12509,N_9186,N_9892);
nor U12510 (N_12510,N_9151,N_11758);
and U12511 (N_12511,N_10648,N_10548);
or U12512 (N_12512,N_11882,N_10896);
nor U12513 (N_12513,N_9102,N_10907);
and U12514 (N_12514,N_10385,N_9650);
nand U12515 (N_12515,N_10036,N_10079);
nand U12516 (N_12516,N_11377,N_9179);
and U12517 (N_12517,N_9886,N_11917);
nand U12518 (N_12518,N_10733,N_11635);
nand U12519 (N_12519,N_10589,N_10120);
nor U12520 (N_12520,N_10418,N_11325);
nor U12521 (N_12521,N_10407,N_10720);
xor U12522 (N_12522,N_9879,N_9344);
or U12523 (N_12523,N_11261,N_10393);
and U12524 (N_12524,N_10477,N_10406);
nand U12525 (N_12525,N_10116,N_11805);
xor U12526 (N_12526,N_10103,N_9095);
or U12527 (N_12527,N_11950,N_10039);
or U12528 (N_12528,N_11972,N_11634);
nor U12529 (N_12529,N_9436,N_10742);
xnor U12530 (N_12530,N_11424,N_11336);
nor U12531 (N_12531,N_11823,N_11512);
nand U12532 (N_12532,N_11439,N_11520);
nor U12533 (N_12533,N_11578,N_10955);
xnor U12534 (N_12534,N_9047,N_11551);
or U12535 (N_12535,N_10040,N_9844);
and U12536 (N_12536,N_9862,N_9541);
or U12537 (N_12537,N_9673,N_10664);
or U12538 (N_12538,N_11652,N_11137);
nand U12539 (N_12539,N_9845,N_11442);
and U12540 (N_12540,N_10024,N_9477);
nand U12541 (N_12541,N_10108,N_10397);
and U12542 (N_12542,N_11266,N_10959);
or U12543 (N_12543,N_9997,N_11351);
and U12544 (N_12544,N_11407,N_10333);
and U12545 (N_12545,N_10999,N_10069);
or U12546 (N_12546,N_10203,N_10254);
nor U12547 (N_12547,N_10524,N_9305);
or U12548 (N_12548,N_9816,N_10707);
xor U12549 (N_12549,N_9431,N_10695);
xnor U12550 (N_12550,N_10882,N_9961);
nor U12551 (N_12551,N_10049,N_11432);
nor U12552 (N_12552,N_10812,N_9681);
nor U12553 (N_12553,N_9925,N_10788);
xor U12554 (N_12554,N_10349,N_9860);
and U12555 (N_12555,N_11344,N_11865);
and U12556 (N_12556,N_10491,N_10600);
nor U12557 (N_12557,N_9116,N_10286);
nor U12558 (N_12558,N_11987,N_9834);
or U12559 (N_12559,N_11110,N_11088);
nand U12560 (N_12560,N_10618,N_10422);
nand U12561 (N_12561,N_11190,N_9999);
xnor U12562 (N_12562,N_10635,N_9863);
or U12563 (N_12563,N_9353,N_9491);
or U12564 (N_12564,N_11631,N_11703);
and U12565 (N_12565,N_11061,N_10062);
and U12566 (N_12566,N_10068,N_9150);
xor U12567 (N_12567,N_9902,N_9606);
and U12568 (N_12568,N_9678,N_10155);
nor U12569 (N_12569,N_10673,N_10414);
or U12570 (N_12570,N_11375,N_9274);
nor U12571 (N_12571,N_10417,N_11595);
or U12572 (N_12572,N_9103,N_10247);
nor U12573 (N_12573,N_10586,N_9087);
nand U12574 (N_12574,N_10150,N_10364);
and U12575 (N_12575,N_9979,N_10667);
and U12576 (N_12576,N_10253,N_11412);
xor U12577 (N_12577,N_9264,N_9207);
xor U12578 (N_12578,N_10888,N_10563);
xor U12579 (N_12579,N_9244,N_11124);
or U12580 (N_12580,N_9258,N_11228);
or U12581 (N_12581,N_10873,N_11821);
xnor U12582 (N_12582,N_9444,N_10370);
xnor U12583 (N_12583,N_10372,N_9250);
nor U12584 (N_12584,N_11020,N_11364);
xnor U12585 (N_12585,N_10779,N_11945);
and U12586 (N_12586,N_10552,N_9727);
and U12587 (N_12587,N_11004,N_10198);
and U12588 (N_12588,N_10394,N_9272);
or U12589 (N_12589,N_11817,N_10786);
nand U12590 (N_12590,N_10428,N_10232);
xor U12591 (N_12591,N_11617,N_11449);
nand U12592 (N_12592,N_9723,N_9544);
nor U12593 (N_12593,N_11289,N_11225);
xnor U12594 (N_12594,N_11267,N_9697);
or U12595 (N_12595,N_9414,N_11283);
and U12596 (N_12596,N_11825,N_11487);
and U12597 (N_12597,N_11246,N_9718);
nand U12598 (N_12598,N_11641,N_10432);
nand U12599 (N_12599,N_10445,N_9842);
nand U12600 (N_12600,N_10502,N_11932);
and U12601 (N_12601,N_11905,N_11276);
xnor U12602 (N_12602,N_11818,N_10362);
or U12603 (N_12603,N_9420,N_10012);
and U12604 (N_12604,N_10797,N_10345);
nand U12605 (N_12605,N_10838,N_11586);
or U12606 (N_12606,N_11660,N_10864);
xor U12607 (N_12607,N_11475,N_11019);
and U12608 (N_12608,N_11463,N_9515);
nand U12609 (N_12609,N_11844,N_9809);
or U12610 (N_12610,N_11182,N_10206);
xnor U12611 (N_12611,N_11992,N_9498);
and U12612 (N_12612,N_9481,N_11524);
nand U12613 (N_12613,N_9058,N_9187);
nand U12614 (N_12614,N_11842,N_11007);
nand U12615 (N_12615,N_10301,N_10452);
or U12616 (N_12616,N_10105,N_11713);
nor U12617 (N_12617,N_11081,N_10416);
or U12618 (N_12618,N_11969,N_11346);
nand U12619 (N_12619,N_11775,N_9865);
nor U12620 (N_12620,N_10623,N_10620);
nor U12621 (N_12621,N_9252,N_11736);
nor U12622 (N_12622,N_10837,N_11253);
or U12623 (N_12623,N_9804,N_10981);
or U12624 (N_12624,N_11651,N_10530);
and U12625 (N_12625,N_9067,N_10020);
nand U12626 (N_12626,N_10080,N_11444);
or U12627 (N_12627,N_10575,N_11545);
nor U12628 (N_12628,N_9253,N_11341);
nand U12629 (N_12629,N_11064,N_9630);
nand U12630 (N_12630,N_11894,N_9191);
or U12631 (N_12631,N_10258,N_10051);
and U12632 (N_12632,N_11706,N_9887);
and U12633 (N_12633,N_9944,N_11403);
nand U12634 (N_12634,N_9401,N_11509);
and U12635 (N_12635,N_9629,N_9463);
and U12636 (N_12636,N_10651,N_9824);
or U12637 (N_12637,N_11334,N_10588);
and U12638 (N_12638,N_11674,N_11675);
and U12639 (N_12639,N_11002,N_11458);
nor U12640 (N_12640,N_11112,N_11073);
and U12641 (N_12641,N_9158,N_10369);
or U12642 (N_12642,N_11451,N_9506);
nand U12643 (N_12643,N_9933,N_9256);
nand U12644 (N_12644,N_11160,N_9756);
xnor U12645 (N_12645,N_11303,N_10223);
nand U12646 (N_12646,N_10894,N_9947);
xor U12647 (N_12647,N_10473,N_11446);
nand U12648 (N_12648,N_10340,N_11518);
xor U12649 (N_12649,N_9554,N_11655);
nor U12650 (N_12650,N_9675,N_9798);
and U12651 (N_12651,N_11138,N_10916);
nand U12652 (N_12652,N_10929,N_11789);
nand U12653 (N_12653,N_10179,N_10805);
nor U12654 (N_12654,N_10462,N_9835);
xnor U12655 (N_12655,N_11227,N_11242);
and U12656 (N_12656,N_10599,N_9929);
nand U12657 (N_12657,N_11321,N_11913);
nand U12658 (N_12658,N_10852,N_11067);
or U12659 (N_12659,N_9866,N_11897);
nand U12660 (N_12660,N_10109,N_10352);
nor U12661 (N_12661,N_10067,N_10978);
nand U12662 (N_12662,N_10824,N_10245);
or U12663 (N_12663,N_10404,N_11472);
and U12664 (N_12664,N_10055,N_9930);
nor U12665 (N_12665,N_9287,N_9295);
or U12666 (N_12666,N_11744,N_11025);
and U12667 (N_12667,N_9785,N_10482);
nor U12668 (N_12668,N_11685,N_9230);
xor U12669 (N_12669,N_9223,N_9662);
or U12670 (N_12670,N_11021,N_11478);
nand U12671 (N_12671,N_9777,N_9338);
and U12672 (N_12672,N_10534,N_9561);
nor U12673 (N_12673,N_9752,N_9738);
nor U12674 (N_12674,N_9748,N_10958);
or U12675 (N_12675,N_11117,N_11841);
nor U12676 (N_12676,N_10321,N_10182);
xor U12677 (N_12677,N_11605,N_10213);
nor U12678 (N_12678,N_10183,N_10764);
nand U12679 (N_12679,N_11948,N_9322);
nand U12680 (N_12680,N_9164,N_10763);
xor U12681 (N_12681,N_9192,N_11320);
nand U12682 (N_12682,N_9243,N_10072);
or U12683 (N_12683,N_10540,N_11479);
or U12684 (N_12684,N_10711,N_11159);
or U12685 (N_12685,N_11773,N_11131);
nand U12686 (N_12686,N_11103,N_10158);
or U12687 (N_12687,N_9144,N_9946);
or U12688 (N_12688,N_11755,N_11275);
xnor U12689 (N_12689,N_9257,N_11065);
xor U12690 (N_12690,N_9114,N_9175);
nand U12691 (N_12691,N_11961,N_9183);
nand U12692 (N_12692,N_10004,N_10226);
nor U12693 (N_12693,N_9905,N_9409);
xor U12694 (N_12694,N_10793,N_10419);
xor U12695 (N_12695,N_11471,N_11097);
xnor U12696 (N_12696,N_9127,N_11921);
xor U12697 (N_12697,N_11123,N_10660);
and U12698 (N_12698,N_11060,N_10821);
or U12699 (N_12699,N_9734,N_10440);
and U12700 (N_12700,N_9983,N_10617);
nand U12701 (N_12701,N_10714,N_10017);
and U12702 (N_12702,N_10030,N_11548);
xnor U12703 (N_12703,N_11079,N_10289);
nor U12704 (N_12704,N_9378,N_11596);
nor U12705 (N_12705,N_9107,N_11732);
or U12706 (N_12706,N_10474,N_9159);
nor U12707 (N_12707,N_11604,N_11696);
xor U12708 (N_12708,N_9452,N_11582);
nor U12709 (N_12709,N_10308,N_11873);
and U12710 (N_12710,N_10165,N_9026);
xnor U12711 (N_12711,N_9658,N_11041);
or U12712 (N_12712,N_11530,N_11748);
nor U12713 (N_12713,N_10576,N_10879);
xor U12714 (N_12714,N_10200,N_9075);
nand U12715 (N_12715,N_9538,N_9872);
or U12716 (N_12716,N_11268,N_9562);
or U12717 (N_12717,N_10777,N_10677);
or U12718 (N_12718,N_11859,N_11863);
and U12719 (N_12719,N_10979,N_9064);
and U12720 (N_12720,N_11369,N_11574);
nand U12721 (N_12721,N_10005,N_9014);
or U12722 (N_12722,N_11173,N_9864);
nor U12723 (N_12723,N_10996,N_9318);
and U12724 (N_12724,N_9613,N_10647);
xnor U12725 (N_12725,N_9280,N_9313);
nor U12726 (N_12726,N_10549,N_10186);
nand U12727 (N_12727,N_9194,N_11947);
and U12728 (N_12728,N_10693,N_10045);
or U12729 (N_12729,N_11953,N_11567);
nor U12730 (N_12730,N_11342,N_11140);
or U12731 (N_12731,N_10316,N_10219);
nand U12732 (N_12732,N_11904,N_11653);
or U12733 (N_12733,N_11366,N_11274);
xor U12734 (N_12734,N_10192,N_10895);
nor U12735 (N_12735,N_9607,N_11170);
and U12736 (N_12736,N_11332,N_11226);
or U12737 (N_12737,N_9234,N_11720);
and U12738 (N_12738,N_9531,N_10063);
nand U12739 (N_12739,N_11188,N_10947);
or U12740 (N_12740,N_11981,N_9282);
and U12741 (N_12741,N_10503,N_11872);
and U12742 (N_12742,N_11384,N_9079);
xor U12743 (N_12743,N_9850,N_9950);
xnor U12744 (N_12744,N_11211,N_9692);
or U12745 (N_12745,N_11100,N_11794);
or U12746 (N_12746,N_11546,N_9980);
xnor U12747 (N_12747,N_9082,N_10134);
nand U12748 (N_12748,N_11210,N_11902);
and U12749 (N_12749,N_9614,N_11647);
nor U12750 (N_12750,N_11045,N_9904);
nor U12751 (N_12751,N_10210,N_9776);
or U12752 (N_12752,N_10702,N_9897);
nand U12753 (N_12753,N_11965,N_11774);
nand U12754 (N_12754,N_10511,N_10107);
nor U12755 (N_12755,N_11464,N_9131);
or U12756 (N_12756,N_10194,N_9968);
and U12757 (N_12757,N_9516,N_11050);
or U12758 (N_12758,N_11243,N_10001);
or U12759 (N_12759,N_9267,N_10136);
xnor U12760 (N_12760,N_9896,N_9108);
and U12761 (N_12761,N_11184,N_9091);
nand U12762 (N_12762,N_10966,N_11146);
xnor U12763 (N_12763,N_9168,N_10436);
xor U12764 (N_12764,N_10771,N_9990);
and U12765 (N_12765,N_11880,N_9006);
nor U12766 (N_12766,N_11926,N_9460);
nor U12767 (N_12767,N_11051,N_10993);
or U12768 (N_12768,N_11359,N_10022);
or U12769 (N_12769,N_11348,N_10785);
nor U12770 (N_12770,N_10140,N_11162);
nor U12771 (N_12771,N_10435,N_9747);
xor U12772 (N_12772,N_9926,N_10177);
and U12773 (N_12773,N_10988,N_11501);
and U12774 (N_12774,N_10731,N_11490);
or U12775 (N_12775,N_11796,N_9009);
xor U12776 (N_12776,N_9167,N_9172);
and U12777 (N_12777,N_11814,N_10521);
and U12778 (N_12778,N_10607,N_9984);
or U12779 (N_12779,N_9390,N_10256);
xnor U12780 (N_12780,N_11646,N_9501);
nand U12781 (N_12781,N_10845,N_10814);
nand U12782 (N_12782,N_9030,N_11602);
nand U12783 (N_12783,N_11915,N_10336);
or U12784 (N_12784,N_10041,N_11489);
xnor U12785 (N_12785,N_11105,N_11704);
nor U12786 (N_12786,N_11541,N_9288);
and U12787 (N_12787,N_11768,N_10494);
xor U12788 (N_12788,N_9085,N_9300);
nor U12789 (N_12789,N_11623,N_10555);
or U12790 (N_12790,N_9132,N_9066);
or U12791 (N_12791,N_10154,N_11496);
and U12792 (N_12792,N_10318,N_11202);
and U12793 (N_12793,N_9343,N_9603);
or U12794 (N_12794,N_11984,N_11637);
and U12795 (N_12795,N_9803,N_9702);
nand U12796 (N_12796,N_11622,N_9077);
nor U12797 (N_12797,N_11322,N_9113);
nor U12798 (N_12798,N_9424,N_9385);
xnor U12799 (N_12799,N_11505,N_10601);
nand U12800 (N_12800,N_11690,N_11772);
or U12801 (N_12801,N_11305,N_11993);
and U12802 (N_12802,N_10217,N_10135);
and U12803 (N_12803,N_11590,N_9324);
and U12804 (N_12804,N_10662,N_10782);
and U12805 (N_12805,N_10199,N_11624);
or U12806 (N_12806,N_11517,N_10222);
nor U12807 (N_12807,N_11466,N_10248);
nor U12808 (N_12808,N_11771,N_9284);
xor U12809 (N_12809,N_11918,N_10826);
or U12810 (N_12810,N_9251,N_11271);
nor U12811 (N_12811,N_10029,N_11671);
nand U12812 (N_12812,N_11107,N_9076);
and U12813 (N_12813,N_9553,N_10337);
xnor U12814 (N_12814,N_9255,N_9002);
nor U12815 (N_12815,N_10086,N_10597);
or U12816 (N_12816,N_9355,N_9184);
xnor U12817 (N_12817,N_11028,N_11888);
nand U12818 (N_12818,N_11832,N_11630);
nand U12819 (N_12819,N_10639,N_11443);
nor U12820 (N_12820,N_10751,N_10765);
and U12821 (N_12821,N_9634,N_11971);
and U12822 (N_12822,N_10802,N_11845);
xor U12823 (N_12823,N_9674,N_9810);
xnor U12824 (N_12824,N_9004,N_9290);
and U12825 (N_12825,N_9788,N_10778);
nand U12826 (N_12826,N_9963,N_10054);
nor U12827 (N_12827,N_10431,N_10636);
nand U12828 (N_12828,N_9563,N_9041);
nor U12829 (N_12829,N_10205,N_10848);
and U12830 (N_12830,N_11113,N_11457);
nor U12831 (N_12831,N_11356,N_9821);
nand U12832 (N_12832,N_11295,N_11040);
nor U12833 (N_12833,N_10887,N_11862);
and U12834 (N_12834,N_11588,N_11864);
xnor U12835 (N_12835,N_11371,N_10853);
or U12836 (N_12836,N_9885,N_9771);
and U12837 (N_12837,N_10214,N_11318);
or U12838 (N_12838,N_10341,N_9276);
xor U12839 (N_12839,N_11511,N_10961);
nor U12840 (N_12840,N_10529,N_10018);
nor U12841 (N_12841,N_10567,N_10293);
nor U12842 (N_12842,N_9731,N_11539);
nand U12843 (N_12843,N_10803,N_9213);
and U12844 (N_12844,N_10366,N_9732);
nand U12845 (N_12845,N_10901,N_10215);
xor U12846 (N_12846,N_10509,N_11010);
or U12847 (N_12847,N_11419,N_10313);
nor U12848 (N_12848,N_11665,N_9503);
or U12849 (N_12849,N_10884,N_11678);
xor U12850 (N_12850,N_9671,N_10320);
nand U12851 (N_12851,N_9408,N_9361);
nand U12852 (N_12852,N_10074,N_10003);
nor U12853 (N_12853,N_9955,N_9817);
nand U12854 (N_12854,N_10917,N_10087);
or U12855 (N_12855,N_11599,N_9286);
nand U12856 (N_12856,N_9373,N_11155);
or U12857 (N_12857,N_11848,N_9769);
or U12858 (N_12858,N_10368,N_10302);
nand U12859 (N_12859,N_11174,N_9228);
xor U12860 (N_12860,N_9743,N_9888);
nor U12861 (N_12861,N_11340,N_10970);
and U12862 (N_12862,N_9293,N_9278);
or U12863 (N_12863,N_10974,N_9546);
or U12864 (N_12864,N_9799,N_11264);
nor U12865 (N_12865,N_10332,N_9139);
or U12866 (N_12866,N_9826,N_10527);
xor U12867 (N_12867,N_9548,N_9259);
xor U12868 (N_12868,N_10840,N_9145);
nor U12869 (N_12869,N_10964,N_11394);
and U12870 (N_12870,N_10444,N_11052);
xor U12871 (N_12871,N_9319,N_10427);
and U12872 (N_12872,N_10810,N_10893);
xnor U12873 (N_12873,N_10874,N_10934);
or U12874 (N_12874,N_9027,N_9749);
nor U12875 (N_12875,N_11540,N_11954);
nor U12876 (N_12876,N_11080,N_11707);
nand U12877 (N_12877,N_11866,N_11759);
nand U12878 (N_12878,N_9720,N_10877);
nand U12879 (N_12879,N_11217,N_9837);
xnor U12880 (N_12880,N_11721,N_11093);
and U12881 (N_12881,N_10942,N_9870);
nand U12882 (N_12882,N_9551,N_9962);
nor U12883 (N_12883,N_11519,N_9021);
and U12884 (N_12884,N_9762,N_10743);
nand U12885 (N_12885,N_11385,N_9231);
nor U12886 (N_12886,N_10594,N_11230);
nand U12887 (N_12887,N_10476,N_10709);
nor U12888 (N_12888,N_10009,N_9993);
nand U12889 (N_12889,N_9547,N_11017);
or U12890 (N_12890,N_11198,N_11260);
and U12891 (N_12891,N_11742,N_11005);
and U12892 (N_12892,N_11657,N_11537);
nand U12893 (N_12893,N_10626,N_9641);
nand U12894 (N_12894,N_10016,N_9323);
nor U12895 (N_12895,N_10830,N_9204);
nor U12896 (N_12896,N_11920,N_11754);
nand U12897 (N_12897,N_11309,N_11506);
and U12898 (N_12898,N_10048,N_11686);
and U12899 (N_12899,N_9740,N_9197);
nor U12900 (N_12900,N_9479,N_11565);
and U12901 (N_12901,N_11572,N_11250);
nand U12902 (N_12902,N_10396,N_9147);
nor U12903 (N_12903,N_10466,N_9007);
xor U12904 (N_12904,N_9812,N_10277);
nand U12905 (N_12905,N_9525,N_10610);
or U12906 (N_12906,N_11310,N_11968);
nor U12907 (N_12907,N_9823,N_11620);
or U12908 (N_12908,N_10665,N_11795);
xnor U12909 (N_12909,N_11994,N_9320);
nor U12910 (N_12910,N_11694,N_10077);
or U12911 (N_12911,N_10229,N_11698);
nand U12912 (N_12912,N_10311,N_9956);
xor U12913 (N_12913,N_10932,N_9713);
xor U12914 (N_12914,N_9188,N_11668);
nor U12915 (N_12915,N_11566,N_11218);
xor U12916 (N_12916,N_11164,N_9584);
xor U12917 (N_12917,N_11378,N_10608);
and U12918 (N_12918,N_10732,N_10218);
nand U12919 (N_12919,N_11222,N_9797);
or U12920 (N_12920,N_9354,N_10264);
nand U12921 (N_12921,N_10335,N_11770);
or U12922 (N_12922,N_10716,N_9120);
xnor U12923 (N_12923,N_11957,N_10756);
or U12924 (N_12924,N_10034,N_10094);
or U12925 (N_12925,N_10211,N_10085);
or U12926 (N_12926,N_10172,N_9394);
nor U12927 (N_12927,N_9375,N_10652);
xnor U12928 (N_12928,N_9433,N_10545);
or U12929 (N_12929,N_11663,N_9441);
nor U12930 (N_12930,N_10161,N_11142);
nor U12931 (N_12931,N_10297,N_11980);
xor U12932 (N_12932,N_11379,N_9488);
or U12933 (N_12933,N_9664,N_11861);
nor U12934 (N_12934,N_10912,N_11317);
and U12935 (N_12935,N_11550,N_10727);
or U12936 (N_12936,N_9940,N_9931);
nand U12937 (N_12937,N_10092,N_11670);
nand U12938 (N_12938,N_10076,N_9969);
nor U12939 (N_12939,N_11033,N_9315);
nand U12940 (N_12940,N_9100,N_11062);
nor U12941 (N_12941,N_9703,N_11868);
or U12942 (N_12942,N_10595,N_11282);
and U12943 (N_12943,N_10921,N_9565);
nand U12944 (N_12944,N_9820,N_10739);
xor U12945 (N_12945,N_10342,N_9403);
or U12946 (N_12946,N_11687,N_9789);
nand U12947 (N_12947,N_11560,N_9340);
xor U12948 (N_12948,N_9964,N_9454);
xor U12949 (N_12949,N_11719,N_11858);
and U12950 (N_12950,N_10479,N_11608);
xor U12951 (N_12951,N_10806,N_10898);
or U12952 (N_12952,N_10460,N_9967);
nor U12953 (N_12953,N_9915,N_10152);
nand U12954 (N_12954,N_11682,N_9889);
nor U12955 (N_12955,N_10037,N_10890);
xnor U12956 (N_12956,N_9504,N_9349);
or U12957 (N_12957,N_11435,N_11843);
and U12958 (N_12958,N_10334,N_10508);
nor U12959 (N_12959,N_9923,N_11656);
nor U12960 (N_12960,N_10144,N_11824);
nand U12961 (N_12961,N_10908,N_9458);
and U12962 (N_12962,N_11710,N_10025);
and U12963 (N_12963,N_10799,N_9308);
or U12964 (N_12964,N_11370,N_10426);
and U12965 (N_12965,N_11023,N_11014);
xor U12966 (N_12966,N_9149,N_9868);
nand U12967 (N_12967,N_9042,N_10188);
nand U12968 (N_12968,N_11054,N_10686);
nor U12969 (N_12969,N_11259,N_9410);
xnor U12970 (N_12970,N_11462,N_10685);
and U12971 (N_12971,N_9101,N_11304);
xor U12972 (N_12972,N_9878,N_9805);
xnor U12973 (N_12973,N_10767,N_10388);
nand U12974 (N_12974,N_10692,N_10230);
and U12975 (N_12975,N_10558,N_9178);
and U12976 (N_12976,N_9618,N_11563);
nand U12977 (N_12977,N_9061,N_9387);
xnor U12978 (N_12978,N_11461,N_10568);
xor U12979 (N_12979,N_10360,N_10469);
and U12980 (N_12980,N_9170,N_11425);
nand U12981 (N_12981,N_11933,N_11411);
and U12982 (N_12982,N_10817,N_11128);
or U12983 (N_12983,N_9791,N_9901);
nand U12984 (N_12984,N_9668,N_9374);
and U12985 (N_12985,N_10453,N_9321);
nor U12986 (N_12986,N_11145,N_9054);
nand U12987 (N_12987,N_9832,N_9128);
xor U12988 (N_12988,N_10291,N_9966);
nor U12989 (N_12989,N_10288,N_11633);
and U12990 (N_12990,N_11193,N_10499);
and U12991 (N_12991,N_10954,N_10447);
or U12992 (N_12992,N_9141,N_11911);
nor U12993 (N_12993,N_11783,N_11361);
nand U12994 (N_12994,N_10455,N_11085);
and U12995 (N_12995,N_9450,N_9920);
or U12996 (N_12996,N_10327,N_10463);
and U12997 (N_12997,N_9783,N_11881);
nand U12998 (N_12998,N_10166,N_10296);
xnor U12999 (N_12999,N_11434,N_9998);
nor U13000 (N_13000,N_9003,N_11428);
nand U13001 (N_13001,N_10992,N_10271);
nor U13002 (N_13002,N_11116,N_10909);
and U13003 (N_13003,N_10272,N_10708);
nand U13004 (N_13004,N_11628,N_11395);
nor U13005 (N_13005,N_9469,N_11912);
nor U13006 (N_13006,N_11299,N_10986);
xnor U13007 (N_13007,N_11066,N_10520);
xor U13008 (N_13008,N_10299,N_10773);
nor U13009 (N_13009,N_11255,N_10688);
nand U13010 (N_13010,N_9205,N_11702);
or U13011 (N_13011,N_10633,N_9040);
nand U13012 (N_13012,N_9530,N_10383);
or U13013 (N_13013,N_10829,N_9086);
xor U13014 (N_13014,N_10353,N_11737);
or U13015 (N_13015,N_11426,N_11705);
nand U13016 (N_13016,N_9709,N_10644);
and U13017 (N_13017,N_10725,N_10056);
or U13018 (N_13018,N_9154,N_11277);
nor U13019 (N_13019,N_9182,N_9297);
nand U13020 (N_13020,N_9157,N_11122);
or U13021 (N_13021,N_11982,N_9919);
xor U13022 (N_13022,N_11437,N_10543);
nor U13023 (N_13023,N_9446,N_9856);
nor U13024 (N_13024,N_11549,N_11148);
and U13025 (N_13025,N_9599,N_9917);
or U13026 (N_13026,N_10236,N_9507);
nand U13027 (N_13027,N_11078,N_11580);
xnor U13028 (N_13028,N_9078,N_10839);
and U13029 (N_13029,N_11247,N_9514);
nor U13030 (N_13030,N_10948,N_11502);
and U13031 (N_13031,N_9445,N_11207);
nand U13032 (N_13032,N_10038,N_11272);
nand U13033 (N_13033,N_10561,N_10866);
and U13034 (N_13034,N_10875,N_10904);
or U13035 (N_13035,N_11454,N_10075);
nand U13036 (N_13036,N_9080,N_11238);
nand U13037 (N_13037,N_10050,N_9594);
and U13038 (N_13038,N_11923,N_11049);
nor U13039 (N_13039,N_11951,N_9219);
nor U13040 (N_13040,N_10820,N_9371);
nor U13041 (N_13041,N_9129,N_9976);
nand U13042 (N_13042,N_11483,N_10629);
nor U13043 (N_13043,N_10746,N_11306);
or U13044 (N_13044,N_11350,N_10591);
xor U13045 (N_13045,N_11096,N_9580);
nor U13046 (N_13046,N_9356,N_9415);
xnor U13047 (N_13047,N_10995,N_10412);
nand U13048 (N_13048,N_9440,N_10863);
nand U13049 (N_13049,N_10204,N_9852);
xor U13050 (N_13050,N_9813,N_11553);
nor U13051 (N_13051,N_9212,N_10250);
and U13052 (N_13052,N_10842,N_11422);
or U13053 (N_13053,N_11284,N_9362);
nor U13054 (N_13054,N_11477,N_10833);
and U13055 (N_13055,N_9457,N_10307);
or U13056 (N_13056,N_11349,N_10121);
or U13057 (N_13057,N_11764,N_10106);
xor U13058 (N_13058,N_11515,N_11035);
nand U13059 (N_13059,N_9096,N_11940);
nor U13060 (N_13060,N_11777,N_10102);
nand U13061 (N_13061,N_11995,N_9376);
nand U13062 (N_13062,N_9914,N_10846);
xnor U13063 (N_13063,N_10281,N_10235);
nor U13064 (N_13064,N_10367,N_9121);
nand U13065 (N_13065,N_10531,N_9225);
nor U13066 (N_13066,N_11157,N_11236);
xnor U13067 (N_13067,N_10065,N_11955);
nand U13068 (N_13068,N_9539,N_9985);
xnor U13069 (N_13069,N_11287,N_11639);
and U13070 (N_13070,N_11558,N_9200);
or U13071 (N_13071,N_11185,N_9598);
or U13072 (N_13072,N_10865,N_11986);
nand U13073 (N_13073,N_11521,N_11642);
and U13074 (N_13074,N_10577,N_9542);
or U13075 (N_13075,N_11281,N_9528);
and U13076 (N_13076,N_10927,N_10678);
nand U13077 (N_13077,N_10690,N_10973);
xnor U13078 (N_13078,N_11573,N_11279);
nor U13079 (N_13079,N_11187,N_11681);
and U13080 (N_13080,N_10471,N_11717);
or U13081 (N_13081,N_9470,N_11836);
nand U13082 (N_13082,N_10314,N_10696);
nor U13083 (N_13083,N_9684,N_9620);
xor U13084 (N_13084,N_9160,N_9719);
xor U13085 (N_13085,N_9388,N_11855);
and U13086 (N_13086,N_11892,N_9427);
nor U13087 (N_13087,N_11239,N_11109);
xnor U13088 (N_13088,N_10472,N_9263);
and U13089 (N_13089,N_10033,N_10234);
nor U13090 (N_13090,N_10645,N_9273);
xnor U13091 (N_13091,N_11039,N_11769);
nor U13092 (N_13092,N_10480,N_9587);
nor U13093 (N_13093,N_11380,N_9489);
and U13094 (N_13094,N_10465,N_11059);
or U13095 (N_13095,N_9948,N_9573);
or U13096 (N_13096,N_10748,N_9778);
nand U13097 (N_13097,N_11445,N_10880);
nor U13098 (N_13098,N_9468,N_10619);
and U13099 (N_13099,N_10251,N_9781);
and U13100 (N_13100,N_11679,N_10726);
nor U13101 (N_13101,N_9642,N_11835);
nor U13102 (N_13102,N_11869,N_9035);
nor U13103 (N_13103,N_9590,N_11363);
nand U13104 (N_13104,N_11569,N_11037);
or U13105 (N_13105,N_11302,N_11896);
xnor U13106 (N_13106,N_10967,N_11837);
and U13107 (N_13107,N_10933,N_11151);
nor U13108 (N_13108,N_10670,N_9505);
nor U13109 (N_13109,N_10911,N_9372);
xnor U13110 (N_13110,N_10174,N_9389);
nand U13111 (N_13111,N_10279,N_9023);
or U13112 (N_13112,N_11074,N_10443);
and U13113 (N_13113,N_11153,N_10844);
xor U13114 (N_13114,N_9722,N_10653);
nor U13115 (N_13115,N_9350,N_9455);
nand U13116 (N_13116,N_9053,N_11741);
or U13117 (N_13117,N_9210,N_10351);
or U13118 (N_13118,N_9974,N_11616);
and U13119 (N_13119,N_11749,N_11510);
or U13120 (N_13120,N_9724,N_9604);
nor U13121 (N_13121,N_10127,N_10338);
and U13122 (N_13122,N_10381,N_9337);
nand U13123 (N_13123,N_10625,N_10878);
and U13124 (N_13124,N_11086,N_9912);
or U13125 (N_13125,N_10631,N_10464);
xor U13126 (N_13126,N_10858,N_11355);
nand U13127 (N_13127,N_11132,N_10807);
and U13128 (N_13128,N_11075,N_10365);
nand U13129 (N_13129,N_10493,N_10273);
or U13130 (N_13130,N_11262,N_11072);
nand U13131 (N_13131,N_11636,N_11315);
or U13132 (N_13132,N_10324,N_11335);
nand U13133 (N_13133,N_11468,N_9482);
nand U13134 (N_13134,N_11946,N_9459);
nand U13135 (N_13135,N_9646,N_9174);
nor U13136 (N_13136,N_9765,N_10114);
and U13137 (N_13137,N_9422,N_9958);
nand U13138 (N_13138,N_11338,N_11672);
and U13139 (N_13139,N_11245,N_9478);
or U13140 (N_13140,N_9248,N_11936);
nand U13141 (N_13141,N_9869,N_10143);
nand U13142 (N_13142,N_10870,N_9838);
nand U13143 (N_13143,N_10938,N_9484);
nor U13144 (N_13144,N_10410,N_9945);
and U13145 (N_13145,N_11658,N_10028);
xor U13146 (N_13146,N_9825,N_10283);
and U13147 (N_13147,N_11555,N_9472);
or U13148 (N_13148,N_10523,N_9246);
and U13149 (N_13149,N_11258,N_10082);
xor U13150 (N_13150,N_9057,N_10402);
and U13151 (N_13151,N_11026,N_9275);
or U13152 (N_13152,N_9090,N_9975);
and U13153 (N_13153,N_11875,N_9402);
nor U13154 (N_13154,N_10679,N_11381);
nand U13155 (N_13155,N_11800,N_11807);
xor U13156 (N_13156,N_9404,N_11730);
nor U13157 (N_13157,N_10701,N_9951);
or U13158 (N_13158,N_11167,N_11711);
nor U13159 (N_13159,N_10095,N_11498);
or U13160 (N_13160,N_11919,N_11659);
or U13161 (N_13161,N_9511,N_10319);
nor U13162 (N_13162,N_10704,N_11988);
nor U13163 (N_13163,N_10730,N_11557);
nor U13164 (N_13164,N_10249,N_11922);
nor U13165 (N_13165,N_10070,N_11467);
or U13166 (N_13166,N_10712,N_11714);
nor U13167 (N_13167,N_10157,N_10478);
nor U13168 (N_13168,N_9384,N_9855);
and U13169 (N_13169,N_10621,N_10122);
nor U13170 (N_13170,N_11779,N_11220);
nor U13171 (N_13171,N_11038,N_10939);
nand U13172 (N_13172,N_10969,N_9593);
xor U13173 (N_13173,N_10862,N_10160);
nor U13174 (N_13174,N_9854,N_10238);
nor U13175 (N_13175,N_9173,N_10854);
or U13176 (N_13176,N_9366,N_10184);
xnor U13177 (N_13177,N_9029,N_10008);
or U13178 (N_13178,N_9895,N_11729);
xnor U13179 (N_13179,N_9020,N_10265);
nand U13180 (N_13180,N_9556,N_11648);
xor U13181 (N_13181,N_11561,N_11229);
or U13182 (N_13182,N_11952,N_9578);
or U13183 (N_13183,N_9537,N_10757);
xor U13184 (N_13184,N_9395,N_9220);
xnor U13185 (N_13185,N_9518,N_9619);
or U13186 (N_13186,N_9203,N_10775);
or U13187 (N_13187,N_10467,N_10241);
nand U13188 (N_13188,N_9190,N_10566);
or U13189 (N_13189,N_11063,N_9741);
nand U13190 (N_13190,N_9001,N_10433);
xnor U13191 (N_13191,N_9465,N_9943);
nor U13192 (N_13192,N_10582,N_10044);
xnor U13193 (N_13193,N_10091,N_10953);
nand U13194 (N_13194,N_10276,N_9216);
or U13195 (N_13195,N_11465,N_11206);
nand U13196 (N_13196,N_9492,N_9269);
nor U13197 (N_13197,N_11664,N_9623);
or U13198 (N_13198,N_9453,N_10945);
nor U13199 (N_13199,N_9291,N_11224);
or U13200 (N_13200,N_11452,N_9569);
nor U13201 (N_13201,N_9487,N_9019);
nand U13202 (N_13202,N_9995,N_10632);
nor U13203 (N_13203,N_10195,N_9737);
xnor U13204 (N_13204,N_10613,N_9659);
or U13205 (N_13205,N_11221,N_10535);
or U13206 (N_13206,N_10506,N_11629);
xor U13207 (N_13207,N_9038,N_11614);
or U13208 (N_13208,N_9891,N_9973);
xnor U13209 (N_13209,N_9307,N_9987);
xnor U13210 (N_13210,N_11941,N_11058);
and U13211 (N_13211,N_9143,N_10905);
nand U13212 (N_13212,N_9500,N_10006);
nor U13213 (N_13213,N_9736,N_10031);
xor U13214 (N_13214,N_11405,N_10899);
nor U13215 (N_13215,N_10573,N_11625);
xnor U13216 (N_13216,N_9626,N_11854);
nand U13217 (N_13217,N_11996,N_9334);
nor U13218 (N_13218,N_10533,N_9549);
or U13219 (N_13219,N_11576,N_11006);
nor U13220 (N_13220,N_9711,N_10951);
and U13221 (N_13221,N_11307,N_9310);
and U13222 (N_13222,N_10818,N_9938);
nand U13223 (N_13223,N_10640,N_11077);
nor U13224 (N_13224,N_9331,N_10752);
or U13225 (N_13225,N_9836,N_11308);
and U13226 (N_13226,N_11766,N_9060);
nor U13227 (N_13227,N_9545,N_10375);
and U13228 (N_13228,N_11234,N_9670);
nor U13229 (N_13229,N_9597,N_9772);
or U13230 (N_13230,N_11976,N_11285);
and U13231 (N_13231,N_9755,N_11290);
xnor U13232 (N_13232,N_10593,N_10496);
nor U13233 (N_13233,N_10298,N_10976);
xnor U13234 (N_13234,N_9126,N_11008);
nor U13235 (N_13235,N_11802,N_10638);
nor U13236 (N_13236,N_10581,N_11024);
nand U13237 (N_13237,N_9296,N_9490);
or U13238 (N_13238,N_11400,N_10946);
or U13239 (N_13239,N_11937,N_10900);
nand U13240 (N_13240,N_9806,N_9000);
xnor U13241 (N_13241,N_9327,N_11722);
nor U13242 (N_13242,N_9767,N_10173);
nand U13243 (N_13243,N_9775,N_10790);
xnor U13244 (N_13244,N_10501,N_11684);
or U13245 (N_13245,N_11964,N_9028);
or U13246 (N_13246,N_9345,N_10886);
nand U13247 (N_13247,N_10781,N_10153);
nand U13248 (N_13248,N_11297,N_10459);
nand U13249 (N_13249,N_9383,N_10099);
and U13250 (N_13250,N_9466,N_9425);
nor U13251 (N_13251,N_11027,N_11293);
or U13252 (N_13252,N_10871,N_11609);
nor U13253 (N_13253,N_10111,N_10242);
and U13254 (N_13254,N_10149,N_9449);
or U13255 (N_13255,N_9705,N_9679);
xor U13256 (N_13256,N_11280,N_10914);
nor U13257 (N_13257,N_11476,N_11482);
nor U13258 (N_13258,N_11393,N_11715);
and U13259 (N_13259,N_9750,N_11695);
or U13260 (N_13260,N_9495,N_9098);
and U13261 (N_13261,N_10832,N_11216);
xor U13262 (N_13262,N_9591,N_10137);
nor U13263 (N_13263,N_10604,N_10663);
xor U13264 (N_13264,N_11029,N_11522);
nand U13265 (N_13265,N_10772,N_10262);
nor U13266 (N_13266,N_9025,N_9971);
or U13267 (N_13267,N_9661,N_10661);
xor U13268 (N_13268,N_10596,N_10944);
nor U13269 (N_13269,N_11189,N_11133);
and U13270 (N_13270,N_10962,N_9687);
nor U13271 (N_13271,N_11763,N_9045);
or U13272 (N_13272,N_9166,N_10569);
and U13273 (N_13273,N_9712,N_10454);
nand U13274 (N_13274,N_11055,N_11979);
nand U13275 (N_13275,N_10510,N_11819);
or U13276 (N_13276,N_11975,N_10243);
nand U13277 (N_13277,N_9624,N_9792);
or U13278 (N_13278,N_11205,N_11788);
or U13279 (N_13279,N_11806,N_9588);
nor U13280 (N_13280,N_10146,N_11154);
nor U13281 (N_13281,N_11492,N_9111);
or U13282 (N_13282,N_9351,N_9992);
and U13283 (N_13283,N_11313,N_10403);
and U13284 (N_13284,N_11312,N_11181);
nand U13285 (N_13285,N_9794,N_11723);
nand U13286 (N_13286,N_9540,N_9032);
and U13287 (N_13287,N_9358,N_10614);
nand U13288 (N_13288,N_10285,N_11526);
and U13289 (N_13289,N_9622,N_9596);
xor U13290 (N_13290,N_9939,N_11822);
and U13291 (N_13291,N_11068,N_11016);
xnor U13292 (N_13292,N_9570,N_11878);
or U13293 (N_13293,N_10963,N_9056);
or U13294 (N_13294,N_11168,N_9586);
and U13295 (N_13295,N_9612,N_9245);
nor U13296 (N_13296,N_10602,N_9266);
nand U13297 (N_13297,N_10538,N_9092);
and U13298 (N_13298,N_11031,N_10572);
xnor U13299 (N_13299,N_9986,N_10741);
or U13300 (N_13300,N_9977,N_10703);
nor U13301 (N_13301,N_9467,N_10957);
xnor U13302 (N_13302,N_11108,N_9289);
and U13303 (N_13303,N_10098,N_11589);
and U13304 (N_13304,N_11372,N_10411);
or U13305 (N_13305,N_11269,N_10000);
or U13306 (N_13306,N_11311,N_11879);
nand U13307 (N_13307,N_10260,N_9728);
nor U13308 (N_13308,N_11516,N_10093);
or U13309 (N_13309,N_9941,N_9462);
nand U13310 (N_13310,N_9013,N_10813);
xor U13311 (N_13311,N_10952,N_9840);
nand U13312 (N_13312,N_9763,N_11183);
or U13313 (N_13313,N_11427,N_9411);
xnor U13314 (N_13314,N_11890,N_10546);
nand U13315 (N_13315,N_11697,N_11352);
nor U13316 (N_13316,N_9893,N_11367);
xor U13317 (N_13317,N_11208,N_10719);
nand U13318 (N_13318,N_11241,N_11801);
and U13319 (N_13319,N_10715,N_11197);
nand U13320 (N_13320,N_11410,N_11076);
nand U13321 (N_13321,N_11812,N_10956);
nand U13322 (N_13322,N_9341,N_10387);
xnor U13323 (N_13323,N_9222,N_9036);
or U13324 (N_13324,N_9847,N_11552);
and U13325 (N_13325,N_11804,N_9566);
or U13326 (N_13326,N_10628,N_11811);
and U13327 (N_13327,N_10303,N_11669);
and U13328 (N_13328,N_10761,N_10088);
nor U13329 (N_13329,N_10002,N_9330);
nor U13330 (N_13330,N_10421,N_9978);
nand U13331 (N_13331,N_11046,N_11362);
xnor U13332 (N_13332,N_11895,N_9024);
nand U13333 (N_13333,N_11973,N_9429);
nor U13334 (N_13334,N_11661,N_10096);
xnor U13335 (N_13335,N_11750,N_11481);
and U13336 (N_13336,N_11830,N_10212);
xor U13337 (N_13337,N_11587,N_10484);
or U13338 (N_13338,N_11249,N_11119);
xnor U13339 (N_13339,N_11469,N_11244);
nand U13340 (N_13340,N_11495,N_11139);
xnor U13341 (N_13341,N_9520,N_9510);
xor U13342 (N_13342,N_11963,N_10735);
nor U13343 (N_13343,N_11331,N_9795);
nor U13344 (N_13344,N_10913,N_10697);
nor U13345 (N_13345,N_9937,N_10449);
nor U13346 (N_13346,N_9616,N_11319);
nand U13347 (N_13347,N_9699,N_9214);
nand U13348 (N_13348,N_9226,N_10078);
nand U13349 (N_13349,N_10724,N_9857);
xnor U13350 (N_13350,N_9579,N_10522);
or U13351 (N_13351,N_9602,N_10949);
xor U13352 (N_13352,N_9475,N_11114);
nor U13353 (N_13353,N_9509,N_9625);
nand U13354 (N_13354,N_9627,N_11135);
and U13355 (N_13355,N_9690,N_10450);
xor U13356 (N_13356,N_9271,N_10747);
nor U13357 (N_13357,N_10363,N_9235);
xor U13358 (N_13358,N_10936,N_11056);
and U13359 (N_13359,N_9153,N_11098);
xor U13360 (N_13360,N_11401,N_9811);
or U13361 (N_13361,N_9364,N_11756);
xnor U13362 (N_13362,N_9122,N_11069);
nand U13363 (N_13363,N_10525,N_9048);
xor U13364 (N_13364,N_11484,N_11531);
and U13365 (N_13365,N_10559,N_11906);
or U13366 (N_13366,N_10379,N_10391);
and U13367 (N_13367,N_9725,N_9779);
nand U13368 (N_13368,N_9676,N_10627);
or U13369 (N_13369,N_11460,N_10274);
and U13370 (N_13370,N_11111,N_10451);
nand U13371 (N_13371,N_11152,N_9648);
nand U13372 (N_13372,N_11886,N_10181);
or U13373 (N_13373,N_9921,N_9416);
nand U13374 (N_13374,N_10941,N_10171);
nand U13375 (N_13375,N_9800,N_10676);
or U13376 (N_13376,N_9575,N_10657);
and U13377 (N_13377,N_10553,N_9657);
or U13378 (N_13378,N_10980,N_9954);
and U13379 (N_13379,N_10532,N_10649);
or U13380 (N_13380,N_10574,N_10193);
xnor U13381 (N_13381,N_11441,N_11543);
nor U13382 (N_13382,N_11931,N_11436);
nor U13383 (N_13383,N_9715,N_9828);
nand U13384 (N_13384,N_11856,N_10755);
nor U13385 (N_13385,N_11785,N_11762);
nor U13386 (N_13386,N_9827,N_10224);
nand U13387 (N_13387,N_9176,N_11013);
nor U13388 (N_13388,N_9397,N_10578);
and U13389 (N_13389,N_11692,N_10208);
or U13390 (N_13390,N_10758,N_9988);
xnor U13391 (N_13391,N_11791,N_9633);
or U13392 (N_13392,N_9701,N_11827);
or U13393 (N_13393,N_9796,N_11693);
xnor U13394 (N_13394,N_9365,N_10304);
nor U13395 (N_13395,N_10164,N_9653);
nor U13396 (N_13396,N_11746,N_11101);
or U13397 (N_13397,N_10269,N_10490);
and U13398 (N_13398,N_10691,N_9908);
nor U13399 (N_13399,N_10737,N_10339);
or U13400 (N_13400,N_9686,N_10922);
or U13401 (N_13401,N_9880,N_11388);
xor U13402 (N_13402,N_10560,N_10931);
and U13403 (N_13403,N_10163,N_9367);
nor U13404 (N_13404,N_11683,N_10889);
nor U13405 (N_13405,N_9688,N_11903);
or U13406 (N_13406,N_10159,N_11383);
xor U13407 (N_13407,N_9208,N_9787);
xor U13408 (N_13408,N_11534,N_9142);
nand U13409 (N_13409,N_11414,N_10448);
nor U13410 (N_13410,N_9861,N_11163);
and U13411 (N_13411,N_10698,N_11161);
and U13412 (N_13412,N_11898,N_9965);
nor U13413 (N_13413,N_11286,N_10046);
and U13414 (N_13414,N_11924,N_10350);
and U13415 (N_13415,N_9801,N_10923);
nor U13416 (N_13416,N_11927,N_10659);
xnor U13417 (N_13417,N_10458,N_10014);
or U13418 (N_13418,N_10675,N_10937);
or U13419 (N_13419,N_9746,N_11048);
and U13420 (N_13420,N_10584,N_10129);
nor U13421 (N_13421,N_10699,N_11392);
xnor U13422 (N_13422,N_10740,N_9526);
xor U13423 (N_13423,N_10759,N_9502);
or U13424 (N_13424,N_9363,N_11960);
or U13425 (N_13425,N_11235,N_9476);
and U13426 (N_13426,N_11071,N_9685);
and U13427 (N_13427,N_9802,N_10869);
and U13428 (N_13428,N_10713,N_9621);
nand U13429 (N_13429,N_11485,N_11877);
or U13430 (N_13430,N_9585,N_11326);
nor U13431 (N_13431,N_10390,N_10885);
xnor U13432 (N_13432,N_10598,N_11570);
xnor U13433 (N_13433,N_11149,N_9218);
nor U13434 (N_13434,N_9261,N_11991);
and U13435 (N_13435,N_11776,N_11339);
xnor U13436 (N_13436,N_9592,N_10300);
xnor U13437 (N_13437,N_11562,N_9137);
or U13438 (N_13438,N_11787,N_11083);
nor U13439 (N_13439,N_9883,N_9227);
nand U13440 (N_13440,N_10380,N_10263);
or U13441 (N_13441,N_10331,N_10784);
nor U13442 (N_13442,N_9906,N_10100);
and U13443 (N_13443,N_10348,N_10019);
nand U13444 (N_13444,N_9413,N_10227);
and U13445 (N_13445,N_11883,N_11389);
and U13446 (N_13446,N_11354,N_9084);
xnor U13447 (N_13447,N_10323,N_10851);
xnor U13448 (N_13448,N_10728,N_10859);
or U13449 (N_13449,N_11734,N_11600);
or U13450 (N_13450,N_10275,N_10982);
nand U13451 (N_13451,N_10073,N_9260);
xor U13452 (N_13452,N_9935,N_11699);
nand U13453 (N_13453,N_11003,N_10228);
nor U13454 (N_13454,N_11610,N_11632);
and U13455 (N_13455,N_10681,N_11448);
nor U13456 (N_13456,N_10497,N_10384);
xnor U13457 (N_13457,N_11480,N_9645);
xor U13458 (N_13458,N_11376,N_9352);
or U13459 (N_13459,N_11396,N_11597);
nand U13460 (N_13460,N_11876,N_10897);
xnor U13461 (N_13461,N_10557,N_11418);
or U13462 (N_13462,N_10646,N_10084);
or U13463 (N_13463,N_11724,N_9298);
nand U13464 (N_13464,N_10131,N_11956);
nand U13465 (N_13465,N_10437,N_10270);
xnor U13466 (N_13466,N_10984,N_11615);
or U13467 (N_13467,N_11962,N_10776);
nor U13468 (N_13468,N_9181,N_11513);
or U13469 (N_13469,N_10831,N_10145);
nor U13470 (N_13470,N_11186,N_11942);
xor U13471 (N_13471,N_11949,N_10668);
or U13472 (N_13472,N_9392,N_9589);
xnor U13473 (N_13473,N_11368,N_9924);
and U13474 (N_13474,N_9770,N_10930);
xnor U13475 (N_13475,N_9683,N_11532);
nor U13476 (N_13476,N_10571,N_11398);
or U13477 (N_13477,N_9774,N_10330);
xnor U13478 (N_13478,N_11125,N_10825);
nor U13479 (N_13479,N_9146,N_10744);
or U13480 (N_13480,N_10774,N_10500);
xor U13481 (N_13481,N_11022,N_9398);
nand U13482 (N_13482,N_11057,N_9807);
or U13483 (N_13483,N_9655,N_11709);
or U13484 (N_13484,N_10420,N_9524);
xnor U13485 (N_13485,N_9497,N_11399);
nand U13486 (N_13486,N_10011,N_9195);
or U13487 (N_13487,N_10528,N_10169);
nor U13488 (N_13488,N_9005,N_9229);
nor U13489 (N_13489,N_9696,N_10811);
xnor U13490 (N_13490,N_10768,N_9447);
nand U13491 (N_13491,N_10903,N_9960);
xnor U13492 (N_13492,N_10518,N_10674);
nand U13493 (N_13493,N_9325,N_11357);
nand U13494 (N_13494,N_11473,N_10481);
and U13495 (N_13495,N_10564,N_10240);
nand U13496 (N_13496,N_10539,N_10485);
nand U13497 (N_13497,N_10590,N_9568);
nand U13498 (N_13498,N_10090,N_10850);
and U13499 (N_13499,N_9138,N_9691);
nor U13500 (N_13500,N_9730,N_10378);
nor U13501 (N_13501,N_10028,N_10852);
xnor U13502 (N_13502,N_10464,N_9207);
nor U13503 (N_13503,N_9114,N_10330);
or U13504 (N_13504,N_10936,N_10138);
nor U13505 (N_13505,N_10541,N_11385);
and U13506 (N_13506,N_9382,N_9968);
xor U13507 (N_13507,N_9775,N_11383);
nand U13508 (N_13508,N_11543,N_11531);
or U13509 (N_13509,N_10250,N_10070);
and U13510 (N_13510,N_11114,N_11784);
nor U13511 (N_13511,N_10230,N_10396);
nand U13512 (N_13512,N_10839,N_9619);
xor U13513 (N_13513,N_11994,N_9137);
xnor U13514 (N_13514,N_9533,N_11652);
or U13515 (N_13515,N_10735,N_9108);
nand U13516 (N_13516,N_10384,N_10475);
or U13517 (N_13517,N_10083,N_9140);
or U13518 (N_13518,N_10138,N_9159);
or U13519 (N_13519,N_10123,N_10179);
nor U13520 (N_13520,N_11074,N_11099);
nor U13521 (N_13521,N_10737,N_9604);
nor U13522 (N_13522,N_11955,N_11012);
and U13523 (N_13523,N_10171,N_10694);
nand U13524 (N_13524,N_11432,N_9968);
nand U13525 (N_13525,N_11255,N_11159);
xnor U13526 (N_13526,N_9756,N_9128);
nor U13527 (N_13527,N_9055,N_10715);
nand U13528 (N_13528,N_10631,N_9374);
nand U13529 (N_13529,N_10883,N_11080);
and U13530 (N_13530,N_11468,N_9077);
and U13531 (N_13531,N_9918,N_11591);
nand U13532 (N_13532,N_9210,N_9720);
nor U13533 (N_13533,N_10815,N_11798);
or U13534 (N_13534,N_11925,N_9860);
nor U13535 (N_13535,N_11545,N_10224);
nor U13536 (N_13536,N_10690,N_9298);
xnor U13537 (N_13537,N_10382,N_10096);
or U13538 (N_13538,N_10218,N_10601);
nor U13539 (N_13539,N_9419,N_9926);
and U13540 (N_13540,N_10999,N_9884);
and U13541 (N_13541,N_10477,N_11248);
nor U13542 (N_13542,N_9387,N_10045);
and U13543 (N_13543,N_11414,N_11876);
or U13544 (N_13544,N_9809,N_9326);
and U13545 (N_13545,N_9426,N_9303);
xnor U13546 (N_13546,N_11885,N_9934);
xor U13547 (N_13547,N_9285,N_11112);
or U13548 (N_13548,N_11496,N_10046);
or U13549 (N_13549,N_10253,N_9590);
xor U13550 (N_13550,N_11208,N_11206);
xnor U13551 (N_13551,N_9270,N_9327);
nor U13552 (N_13552,N_10183,N_11689);
xor U13553 (N_13553,N_11652,N_9636);
nand U13554 (N_13554,N_10451,N_10658);
nor U13555 (N_13555,N_10257,N_10813);
or U13556 (N_13556,N_10159,N_10388);
xor U13557 (N_13557,N_10509,N_10544);
xnor U13558 (N_13558,N_11504,N_9336);
and U13559 (N_13559,N_10857,N_10684);
or U13560 (N_13560,N_10888,N_11940);
and U13561 (N_13561,N_9239,N_9702);
xnor U13562 (N_13562,N_11262,N_10004);
nor U13563 (N_13563,N_10755,N_9931);
nor U13564 (N_13564,N_10613,N_9095);
nor U13565 (N_13565,N_9332,N_11881);
xnor U13566 (N_13566,N_11055,N_11719);
xnor U13567 (N_13567,N_10080,N_10113);
and U13568 (N_13568,N_9333,N_10749);
or U13569 (N_13569,N_10789,N_9957);
nor U13570 (N_13570,N_11208,N_10321);
xor U13571 (N_13571,N_9370,N_10309);
xnor U13572 (N_13572,N_10524,N_11707);
nor U13573 (N_13573,N_10331,N_11004);
and U13574 (N_13574,N_9055,N_11283);
nor U13575 (N_13575,N_11283,N_11332);
or U13576 (N_13576,N_10912,N_11770);
xor U13577 (N_13577,N_9755,N_11722);
nor U13578 (N_13578,N_9288,N_9000);
nor U13579 (N_13579,N_9673,N_11768);
nand U13580 (N_13580,N_11313,N_11706);
and U13581 (N_13581,N_9800,N_11831);
nand U13582 (N_13582,N_11358,N_10275);
nor U13583 (N_13583,N_9714,N_10902);
nand U13584 (N_13584,N_10434,N_11503);
xnor U13585 (N_13585,N_9476,N_9561);
or U13586 (N_13586,N_10388,N_9097);
nand U13587 (N_13587,N_9787,N_11132);
xnor U13588 (N_13588,N_10319,N_10099);
or U13589 (N_13589,N_10997,N_9079);
nand U13590 (N_13590,N_9518,N_10954);
and U13591 (N_13591,N_9791,N_11080);
xor U13592 (N_13592,N_10530,N_9178);
or U13593 (N_13593,N_10938,N_10430);
or U13594 (N_13594,N_9434,N_9958);
or U13595 (N_13595,N_10363,N_11902);
or U13596 (N_13596,N_11289,N_11374);
xnor U13597 (N_13597,N_10388,N_9308);
nor U13598 (N_13598,N_9330,N_9850);
nand U13599 (N_13599,N_11060,N_10932);
nand U13600 (N_13600,N_11098,N_10801);
xnor U13601 (N_13601,N_9627,N_9465);
nand U13602 (N_13602,N_10414,N_9596);
xnor U13603 (N_13603,N_11552,N_9734);
xor U13604 (N_13604,N_9839,N_10205);
xnor U13605 (N_13605,N_11126,N_9539);
or U13606 (N_13606,N_9003,N_10769);
and U13607 (N_13607,N_9119,N_9278);
nand U13608 (N_13608,N_11945,N_10313);
xor U13609 (N_13609,N_10579,N_11769);
xor U13610 (N_13610,N_10104,N_9342);
and U13611 (N_13611,N_10801,N_9239);
nand U13612 (N_13612,N_10381,N_9156);
nor U13613 (N_13613,N_11441,N_10886);
or U13614 (N_13614,N_11677,N_11369);
xnor U13615 (N_13615,N_10131,N_9989);
xor U13616 (N_13616,N_9495,N_9053);
nand U13617 (N_13617,N_10320,N_10363);
and U13618 (N_13618,N_9575,N_11026);
and U13619 (N_13619,N_11031,N_10900);
and U13620 (N_13620,N_10054,N_9954);
or U13621 (N_13621,N_10911,N_11558);
or U13622 (N_13622,N_9174,N_10123);
and U13623 (N_13623,N_9158,N_11725);
nor U13624 (N_13624,N_9574,N_9756);
nor U13625 (N_13625,N_10213,N_11116);
and U13626 (N_13626,N_11268,N_11831);
or U13627 (N_13627,N_11706,N_9094);
xnor U13628 (N_13628,N_10076,N_10097);
and U13629 (N_13629,N_9571,N_11491);
and U13630 (N_13630,N_11355,N_9538);
and U13631 (N_13631,N_9041,N_11387);
nor U13632 (N_13632,N_9626,N_9282);
and U13633 (N_13633,N_9009,N_11037);
xnor U13634 (N_13634,N_10984,N_9683);
nand U13635 (N_13635,N_9216,N_11991);
nor U13636 (N_13636,N_9732,N_11820);
nand U13637 (N_13637,N_9903,N_11081);
or U13638 (N_13638,N_9322,N_10372);
or U13639 (N_13639,N_10171,N_10708);
xor U13640 (N_13640,N_9069,N_11841);
nor U13641 (N_13641,N_10878,N_10340);
xnor U13642 (N_13642,N_9599,N_9582);
nor U13643 (N_13643,N_11529,N_10780);
nand U13644 (N_13644,N_9739,N_11420);
or U13645 (N_13645,N_11378,N_10300);
or U13646 (N_13646,N_10425,N_10764);
or U13647 (N_13647,N_9085,N_9284);
and U13648 (N_13648,N_11080,N_9122);
nand U13649 (N_13649,N_10135,N_10943);
xnor U13650 (N_13650,N_10169,N_10447);
nor U13651 (N_13651,N_10995,N_10296);
nor U13652 (N_13652,N_10873,N_10072);
xor U13653 (N_13653,N_10989,N_10185);
nor U13654 (N_13654,N_11940,N_9298);
and U13655 (N_13655,N_9023,N_11576);
nand U13656 (N_13656,N_10718,N_10327);
xnor U13657 (N_13657,N_9148,N_9091);
xor U13658 (N_13658,N_9069,N_10738);
or U13659 (N_13659,N_9253,N_9357);
xnor U13660 (N_13660,N_9786,N_10980);
or U13661 (N_13661,N_11653,N_9799);
or U13662 (N_13662,N_9195,N_9166);
nor U13663 (N_13663,N_9785,N_10655);
nand U13664 (N_13664,N_11363,N_11941);
or U13665 (N_13665,N_11197,N_10443);
nand U13666 (N_13666,N_11572,N_10910);
xnor U13667 (N_13667,N_9027,N_11371);
and U13668 (N_13668,N_11299,N_9942);
nor U13669 (N_13669,N_9540,N_11362);
and U13670 (N_13670,N_10444,N_11106);
or U13671 (N_13671,N_11886,N_9549);
nand U13672 (N_13672,N_11066,N_11234);
nor U13673 (N_13673,N_11087,N_11012);
or U13674 (N_13674,N_11217,N_9617);
nand U13675 (N_13675,N_11178,N_9741);
or U13676 (N_13676,N_9833,N_9888);
nand U13677 (N_13677,N_11367,N_9085);
and U13678 (N_13678,N_9556,N_10850);
nor U13679 (N_13679,N_11712,N_10576);
xor U13680 (N_13680,N_10165,N_9790);
nand U13681 (N_13681,N_11085,N_9000);
and U13682 (N_13682,N_10892,N_9569);
or U13683 (N_13683,N_9672,N_10771);
nor U13684 (N_13684,N_9695,N_9872);
nand U13685 (N_13685,N_10949,N_9513);
nor U13686 (N_13686,N_11797,N_10023);
nor U13687 (N_13687,N_10988,N_11279);
or U13688 (N_13688,N_10241,N_10629);
nor U13689 (N_13689,N_9940,N_9101);
and U13690 (N_13690,N_10630,N_11259);
or U13691 (N_13691,N_10260,N_11152);
nand U13692 (N_13692,N_11857,N_11447);
xnor U13693 (N_13693,N_11834,N_10956);
nand U13694 (N_13694,N_9001,N_11637);
xor U13695 (N_13695,N_9426,N_11521);
nor U13696 (N_13696,N_9779,N_11238);
or U13697 (N_13697,N_10064,N_10239);
nor U13698 (N_13698,N_9857,N_9998);
or U13699 (N_13699,N_10769,N_10773);
nor U13700 (N_13700,N_9439,N_10627);
or U13701 (N_13701,N_9055,N_10288);
nor U13702 (N_13702,N_11376,N_11439);
or U13703 (N_13703,N_9053,N_10621);
nand U13704 (N_13704,N_11788,N_10019);
xor U13705 (N_13705,N_10820,N_9881);
or U13706 (N_13706,N_11738,N_9576);
nand U13707 (N_13707,N_9808,N_9925);
and U13708 (N_13708,N_10620,N_9418);
nor U13709 (N_13709,N_9556,N_11579);
nand U13710 (N_13710,N_10833,N_11303);
nor U13711 (N_13711,N_9334,N_11814);
nor U13712 (N_13712,N_11299,N_11955);
or U13713 (N_13713,N_9254,N_11748);
nand U13714 (N_13714,N_9966,N_9051);
nand U13715 (N_13715,N_9417,N_11969);
nor U13716 (N_13716,N_11852,N_11946);
xor U13717 (N_13717,N_9789,N_9278);
nor U13718 (N_13718,N_11547,N_9534);
nor U13719 (N_13719,N_9636,N_10811);
nor U13720 (N_13720,N_9890,N_9439);
and U13721 (N_13721,N_9009,N_11613);
nor U13722 (N_13722,N_9027,N_9656);
xnor U13723 (N_13723,N_9975,N_9265);
or U13724 (N_13724,N_11239,N_11999);
nor U13725 (N_13725,N_9387,N_11644);
and U13726 (N_13726,N_11755,N_10579);
nor U13727 (N_13727,N_11175,N_11342);
xnor U13728 (N_13728,N_10084,N_10205);
nor U13729 (N_13729,N_9061,N_11538);
xnor U13730 (N_13730,N_11339,N_9528);
nor U13731 (N_13731,N_10105,N_9794);
xor U13732 (N_13732,N_11740,N_10732);
nand U13733 (N_13733,N_11451,N_11053);
or U13734 (N_13734,N_9502,N_11024);
or U13735 (N_13735,N_9158,N_10299);
nor U13736 (N_13736,N_10426,N_9180);
or U13737 (N_13737,N_11859,N_11785);
or U13738 (N_13738,N_11803,N_11197);
nor U13739 (N_13739,N_10761,N_9281);
nand U13740 (N_13740,N_11921,N_10008);
and U13741 (N_13741,N_11456,N_9337);
and U13742 (N_13742,N_9568,N_11282);
nand U13743 (N_13743,N_11403,N_9221);
nor U13744 (N_13744,N_11622,N_10836);
nor U13745 (N_13745,N_11492,N_11085);
or U13746 (N_13746,N_10818,N_11187);
and U13747 (N_13747,N_9565,N_10200);
xnor U13748 (N_13748,N_9343,N_11359);
or U13749 (N_13749,N_10679,N_10853);
nor U13750 (N_13750,N_10738,N_9378);
nand U13751 (N_13751,N_10862,N_11557);
nor U13752 (N_13752,N_11476,N_10066);
and U13753 (N_13753,N_9190,N_9768);
and U13754 (N_13754,N_10109,N_9800);
or U13755 (N_13755,N_9155,N_10375);
nand U13756 (N_13756,N_10721,N_9065);
or U13757 (N_13757,N_11058,N_11024);
nor U13758 (N_13758,N_10580,N_9437);
nand U13759 (N_13759,N_9421,N_11436);
or U13760 (N_13760,N_11303,N_11109);
nand U13761 (N_13761,N_10879,N_10612);
nand U13762 (N_13762,N_9098,N_10754);
xor U13763 (N_13763,N_11476,N_9919);
and U13764 (N_13764,N_9327,N_10360);
and U13765 (N_13765,N_11467,N_9999);
xnor U13766 (N_13766,N_9376,N_10558);
or U13767 (N_13767,N_9557,N_11686);
xnor U13768 (N_13768,N_10679,N_10450);
nand U13769 (N_13769,N_11792,N_9604);
xnor U13770 (N_13770,N_11481,N_9573);
xor U13771 (N_13771,N_11565,N_10844);
and U13772 (N_13772,N_11616,N_9446);
or U13773 (N_13773,N_11152,N_9353);
and U13774 (N_13774,N_9787,N_9762);
or U13775 (N_13775,N_11661,N_9779);
nor U13776 (N_13776,N_9859,N_9226);
or U13777 (N_13777,N_9160,N_10243);
xor U13778 (N_13778,N_11698,N_9919);
or U13779 (N_13779,N_10278,N_9561);
and U13780 (N_13780,N_9848,N_10993);
xor U13781 (N_13781,N_9229,N_11951);
nand U13782 (N_13782,N_11118,N_10490);
nand U13783 (N_13783,N_10716,N_9803);
and U13784 (N_13784,N_11672,N_11127);
xor U13785 (N_13785,N_11351,N_9176);
and U13786 (N_13786,N_10859,N_11846);
nand U13787 (N_13787,N_11911,N_11364);
nand U13788 (N_13788,N_9930,N_11597);
and U13789 (N_13789,N_11232,N_10962);
or U13790 (N_13790,N_10144,N_10989);
or U13791 (N_13791,N_10273,N_11315);
xor U13792 (N_13792,N_11668,N_11204);
nand U13793 (N_13793,N_11516,N_11285);
nand U13794 (N_13794,N_10199,N_10032);
nor U13795 (N_13795,N_11322,N_10331);
and U13796 (N_13796,N_11598,N_10322);
and U13797 (N_13797,N_9346,N_9807);
or U13798 (N_13798,N_10874,N_10929);
and U13799 (N_13799,N_10023,N_11000);
xor U13800 (N_13800,N_9129,N_9769);
or U13801 (N_13801,N_10297,N_9144);
or U13802 (N_13802,N_11537,N_10812);
nor U13803 (N_13803,N_10590,N_10195);
or U13804 (N_13804,N_11143,N_11168);
xor U13805 (N_13805,N_10938,N_9517);
or U13806 (N_13806,N_11398,N_11493);
nand U13807 (N_13807,N_10808,N_11585);
and U13808 (N_13808,N_11280,N_11426);
nand U13809 (N_13809,N_9618,N_10023);
nor U13810 (N_13810,N_10154,N_9123);
nor U13811 (N_13811,N_10124,N_10075);
nand U13812 (N_13812,N_10710,N_9634);
and U13813 (N_13813,N_10181,N_10840);
nand U13814 (N_13814,N_11485,N_10350);
or U13815 (N_13815,N_11518,N_11046);
nor U13816 (N_13816,N_11733,N_11719);
and U13817 (N_13817,N_10743,N_9610);
nor U13818 (N_13818,N_10939,N_11927);
nand U13819 (N_13819,N_10672,N_11882);
or U13820 (N_13820,N_9666,N_11476);
nor U13821 (N_13821,N_10488,N_10931);
xor U13822 (N_13822,N_9289,N_10109);
and U13823 (N_13823,N_11177,N_9990);
nand U13824 (N_13824,N_10830,N_9684);
or U13825 (N_13825,N_10737,N_10298);
and U13826 (N_13826,N_10784,N_9551);
nor U13827 (N_13827,N_11259,N_9942);
xor U13828 (N_13828,N_9219,N_9649);
nor U13829 (N_13829,N_10653,N_9920);
nor U13830 (N_13830,N_11942,N_9134);
xnor U13831 (N_13831,N_9148,N_10883);
xor U13832 (N_13832,N_11466,N_10863);
nor U13833 (N_13833,N_11678,N_10989);
nor U13834 (N_13834,N_10272,N_11793);
and U13835 (N_13835,N_9582,N_11991);
nand U13836 (N_13836,N_11621,N_10443);
xnor U13837 (N_13837,N_10826,N_11236);
nand U13838 (N_13838,N_10010,N_9817);
nor U13839 (N_13839,N_10600,N_9368);
and U13840 (N_13840,N_11865,N_10106);
and U13841 (N_13841,N_9573,N_11116);
and U13842 (N_13842,N_9578,N_11038);
nor U13843 (N_13843,N_10090,N_11974);
and U13844 (N_13844,N_11815,N_11675);
nand U13845 (N_13845,N_9790,N_9803);
xor U13846 (N_13846,N_11145,N_10028);
xnor U13847 (N_13847,N_9490,N_9426);
nor U13848 (N_13848,N_9386,N_10286);
xor U13849 (N_13849,N_9801,N_9107);
or U13850 (N_13850,N_10833,N_11017);
or U13851 (N_13851,N_9194,N_9001);
nor U13852 (N_13852,N_11105,N_10867);
nor U13853 (N_13853,N_11136,N_9463);
and U13854 (N_13854,N_9294,N_10853);
nor U13855 (N_13855,N_11055,N_11829);
and U13856 (N_13856,N_10033,N_11255);
or U13857 (N_13857,N_11978,N_9632);
nand U13858 (N_13858,N_9249,N_10800);
nor U13859 (N_13859,N_9689,N_10913);
and U13860 (N_13860,N_10721,N_10574);
nor U13861 (N_13861,N_10401,N_11531);
xor U13862 (N_13862,N_10924,N_10363);
and U13863 (N_13863,N_11740,N_9975);
or U13864 (N_13864,N_11687,N_10410);
and U13865 (N_13865,N_10343,N_9287);
or U13866 (N_13866,N_10026,N_11661);
or U13867 (N_13867,N_10810,N_9627);
nor U13868 (N_13868,N_9425,N_10328);
xor U13869 (N_13869,N_9770,N_10321);
nor U13870 (N_13870,N_11433,N_9123);
nor U13871 (N_13871,N_11979,N_11222);
xor U13872 (N_13872,N_11373,N_10058);
xnor U13873 (N_13873,N_9404,N_10155);
xor U13874 (N_13874,N_11910,N_9051);
nor U13875 (N_13875,N_10704,N_9186);
nand U13876 (N_13876,N_10398,N_10968);
and U13877 (N_13877,N_9681,N_10797);
nor U13878 (N_13878,N_9416,N_9851);
and U13879 (N_13879,N_11985,N_10251);
nand U13880 (N_13880,N_10254,N_11223);
and U13881 (N_13881,N_11672,N_9203);
nand U13882 (N_13882,N_11080,N_10973);
and U13883 (N_13883,N_9727,N_9038);
xor U13884 (N_13884,N_10202,N_10967);
and U13885 (N_13885,N_11762,N_9035);
or U13886 (N_13886,N_11138,N_9477);
nor U13887 (N_13887,N_11641,N_11251);
nand U13888 (N_13888,N_9150,N_11042);
nor U13889 (N_13889,N_9281,N_9925);
and U13890 (N_13890,N_10242,N_11236);
xnor U13891 (N_13891,N_11203,N_9743);
or U13892 (N_13892,N_11018,N_10379);
nor U13893 (N_13893,N_9172,N_10214);
or U13894 (N_13894,N_10807,N_9692);
or U13895 (N_13895,N_10043,N_10039);
nand U13896 (N_13896,N_11765,N_11299);
xor U13897 (N_13897,N_9077,N_9818);
nand U13898 (N_13898,N_9112,N_9374);
and U13899 (N_13899,N_11039,N_10594);
or U13900 (N_13900,N_11161,N_9176);
nand U13901 (N_13901,N_10098,N_10316);
nor U13902 (N_13902,N_10598,N_9441);
and U13903 (N_13903,N_9335,N_10522);
and U13904 (N_13904,N_10366,N_9115);
nand U13905 (N_13905,N_9744,N_10450);
xnor U13906 (N_13906,N_10094,N_9365);
and U13907 (N_13907,N_9274,N_11733);
and U13908 (N_13908,N_11762,N_9295);
or U13909 (N_13909,N_10027,N_9943);
or U13910 (N_13910,N_11905,N_11086);
and U13911 (N_13911,N_9203,N_10273);
nor U13912 (N_13912,N_10460,N_9654);
or U13913 (N_13913,N_10161,N_10411);
xor U13914 (N_13914,N_11047,N_9008);
and U13915 (N_13915,N_10707,N_11869);
nand U13916 (N_13916,N_9718,N_10936);
nor U13917 (N_13917,N_11413,N_10201);
nand U13918 (N_13918,N_11339,N_9498);
or U13919 (N_13919,N_9701,N_9859);
xnor U13920 (N_13920,N_9077,N_10501);
or U13921 (N_13921,N_10951,N_11186);
xnor U13922 (N_13922,N_11206,N_11666);
xor U13923 (N_13923,N_10423,N_11215);
xnor U13924 (N_13924,N_9311,N_9148);
and U13925 (N_13925,N_9904,N_9181);
xor U13926 (N_13926,N_11417,N_11502);
xor U13927 (N_13927,N_9095,N_11859);
or U13928 (N_13928,N_10648,N_10479);
xnor U13929 (N_13929,N_9101,N_9108);
nand U13930 (N_13930,N_9365,N_11217);
nand U13931 (N_13931,N_9445,N_11361);
nand U13932 (N_13932,N_11707,N_11876);
nand U13933 (N_13933,N_9806,N_10803);
nor U13934 (N_13934,N_10798,N_10765);
or U13935 (N_13935,N_9566,N_11937);
nand U13936 (N_13936,N_10565,N_10817);
nand U13937 (N_13937,N_9189,N_10926);
or U13938 (N_13938,N_11645,N_10969);
and U13939 (N_13939,N_11895,N_10485);
nor U13940 (N_13940,N_9264,N_11865);
nor U13941 (N_13941,N_9345,N_11724);
and U13942 (N_13942,N_9786,N_9868);
or U13943 (N_13943,N_10153,N_9262);
nor U13944 (N_13944,N_10783,N_9220);
nand U13945 (N_13945,N_9199,N_10278);
nand U13946 (N_13946,N_11655,N_9783);
or U13947 (N_13947,N_9893,N_10034);
and U13948 (N_13948,N_9933,N_11637);
and U13949 (N_13949,N_10219,N_10194);
xnor U13950 (N_13950,N_11222,N_10770);
nor U13951 (N_13951,N_10368,N_11698);
and U13952 (N_13952,N_10395,N_10363);
nand U13953 (N_13953,N_10831,N_9422);
nor U13954 (N_13954,N_11630,N_9902);
and U13955 (N_13955,N_10888,N_11905);
nand U13956 (N_13956,N_9377,N_10277);
or U13957 (N_13957,N_10895,N_10839);
or U13958 (N_13958,N_9766,N_9558);
and U13959 (N_13959,N_9904,N_11940);
xor U13960 (N_13960,N_9893,N_9724);
xnor U13961 (N_13961,N_10828,N_11188);
xnor U13962 (N_13962,N_10750,N_11847);
xnor U13963 (N_13963,N_10900,N_11752);
xnor U13964 (N_13964,N_9291,N_10748);
nor U13965 (N_13965,N_9413,N_10114);
nor U13966 (N_13966,N_10671,N_11567);
nor U13967 (N_13967,N_10883,N_10859);
xor U13968 (N_13968,N_11773,N_11517);
and U13969 (N_13969,N_9255,N_10587);
nand U13970 (N_13970,N_10794,N_10895);
nor U13971 (N_13971,N_10234,N_10873);
and U13972 (N_13972,N_11551,N_11309);
nand U13973 (N_13973,N_10656,N_9872);
and U13974 (N_13974,N_9086,N_10760);
and U13975 (N_13975,N_9232,N_9477);
nand U13976 (N_13976,N_10327,N_9910);
nand U13977 (N_13977,N_11967,N_11876);
xnor U13978 (N_13978,N_9863,N_9018);
and U13979 (N_13979,N_9689,N_9264);
nand U13980 (N_13980,N_10181,N_10144);
nor U13981 (N_13981,N_9182,N_11051);
and U13982 (N_13982,N_9091,N_10336);
or U13983 (N_13983,N_9324,N_11529);
or U13984 (N_13984,N_9199,N_11519);
or U13985 (N_13985,N_9680,N_11735);
nand U13986 (N_13986,N_10802,N_10814);
nor U13987 (N_13987,N_10974,N_11097);
and U13988 (N_13988,N_11493,N_11967);
or U13989 (N_13989,N_9275,N_9855);
or U13990 (N_13990,N_10870,N_10424);
and U13991 (N_13991,N_11420,N_9412);
nor U13992 (N_13992,N_10714,N_9742);
nor U13993 (N_13993,N_11064,N_11818);
and U13994 (N_13994,N_10764,N_10464);
nor U13995 (N_13995,N_10075,N_10313);
nor U13996 (N_13996,N_11522,N_11280);
nand U13997 (N_13997,N_11320,N_10309);
xnor U13998 (N_13998,N_10507,N_9522);
or U13999 (N_13999,N_10398,N_10418);
nor U14000 (N_14000,N_11812,N_9689);
or U14001 (N_14001,N_10756,N_9570);
nor U14002 (N_14002,N_9201,N_10238);
nand U14003 (N_14003,N_10485,N_10295);
and U14004 (N_14004,N_9715,N_11883);
nor U14005 (N_14005,N_9262,N_11274);
xnor U14006 (N_14006,N_11123,N_9593);
nor U14007 (N_14007,N_10614,N_11104);
or U14008 (N_14008,N_11495,N_9336);
or U14009 (N_14009,N_11894,N_11730);
nor U14010 (N_14010,N_11882,N_9046);
or U14011 (N_14011,N_9772,N_9542);
nor U14012 (N_14012,N_9453,N_9112);
nor U14013 (N_14013,N_10928,N_10151);
xor U14014 (N_14014,N_11798,N_10971);
or U14015 (N_14015,N_9915,N_11413);
xnor U14016 (N_14016,N_11370,N_11274);
or U14017 (N_14017,N_9372,N_11306);
or U14018 (N_14018,N_11677,N_9470);
nor U14019 (N_14019,N_10752,N_9715);
and U14020 (N_14020,N_9163,N_10964);
nor U14021 (N_14021,N_11891,N_9241);
nor U14022 (N_14022,N_10813,N_10262);
nor U14023 (N_14023,N_11476,N_11648);
xnor U14024 (N_14024,N_10469,N_9168);
or U14025 (N_14025,N_9919,N_10407);
nor U14026 (N_14026,N_11582,N_11336);
and U14027 (N_14027,N_9047,N_10013);
or U14028 (N_14028,N_9230,N_11765);
nand U14029 (N_14029,N_9525,N_10990);
nand U14030 (N_14030,N_10643,N_11804);
nor U14031 (N_14031,N_9580,N_9886);
nand U14032 (N_14032,N_10793,N_10370);
xnor U14033 (N_14033,N_9895,N_11215);
or U14034 (N_14034,N_10046,N_10189);
nand U14035 (N_14035,N_11843,N_10690);
or U14036 (N_14036,N_10863,N_10299);
and U14037 (N_14037,N_10112,N_11881);
and U14038 (N_14038,N_9420,N_11364);
xnor U14039 (N_14039,N_10347,N_9003);
nor U14040 (N_14040,N_9682,N_10880);
or U14041 (N_14041,N_11962,N_11867);
or U14042 (N_14042,N_11597,N_11084);
or U14043 (N_14043,N_10561,N_11852);
or U14044 (N_14044,N_10138,N_10106);
or U14045 (N_14045,N_11506,N_10468);
nand U14046 (N_14046,N_11853,N_10834);
nand U14047 (N_14047,N_11714,N_10815);
xnor U14048 (N_14048,N_11379,N_9894);
nor U14049 (N_14049,N_11764,N_10455);
xor U14050 (N_14050,N_10716,N_10975);
xor U14051 (N_14051,N_11299,N_11784);
and U14052 (N_14052,N_9619,N_9974);
nor U14053 (N_14053,N_10970,N_11949);
xnor U14054 (N_14054,N_9725,N_10977);
and U14055 (N_14055,N_10686,N_9337);
or U14056 (N_14056,N_10167,N_11417);
and U14057 (N_14057,N_11753,N_9483);
or U14058 (N_14058,N_10541,N_9303);
nand U14059 (N_14059,N_9486,N_10488);
and U14060 (N_14060,N_11585,N_9047);
or U14061 (N_14061,N_11351,N_10613);
xor U14062 (N_14062,N_11474,N_11247);
nand U14063 (N_14063,N_9481,N_10831);
or U14064 (N_14064,N_9337,N_9340);
nor U14065 (N_14065,N_9818,N_9501);
and U14066 (N_14066,N_11768,N_10118);
xor U14067 (N_14067,N_9382,N_11245);
nand U14068 (N_14068,N_9145,N_9740);
or U14069 (N_14069,N_11286,N_9684);
and U14070 (N_14070,N_9349,N_9575);
or U14071 (N_14071,N_10775,N_11696);
xnor U14072 (N_14072,N_10780,N_11507);
nand U14073 (N_14073,N_11962,N_11726);
nor U14074 (N_14074,N_10232,N_9957);
or U14075 (N_14075,N_10738,N_10826);
nor U14076 (N_14076,N_11421,N_11499);
nand U14077 (N_14077,N_11157,N_9420);
xor U14078 (N_14078,N_11969,N_9720);
and U14079 (N_14079,N_10217,N_11028);
and U14080 (N_14080,N_11300,N_11582);
xnor U14081 (N_14081,N_11601,N_11911);
nand U14082 (N_14082,N_9357,N_9150);
xnor U14083 (N_14083,N_10723,N_11613);
xnor U14084 (N_14084,N_11897,N_9574);
or U14085 (N_14085,N_10695,N_11954);
and U14086 (N_14086,N_10509,N_10094);
nor U14087 (N_14087,N_10814,N_10627);
nand U14088 (N_14088,N_10722,N_10983);
or U14089 (N_14089,N_9089,N_11335);
and U14090 (N_14090,N_10620,N_11762);
nor U14091 (N_14091,N_11738,N_9607);
nand U14092 (N_14092,N_10971,N_11373);
nor U14093 (N_14093,N_11233,N_10489);
xnor U14094 (N_14094,N_9751,N_11938);
or U14095 (N_14095,N_9555,N_10348);
nand U14096 (N_14096,N_9237,N_10161);
and U14097 (N_14097,N_9236,N_11822);
nor U14098 (N_14098,N_11972,N_11598);
or U14099 (N_14099,N_9240,N_11772);
nor U14100 (N_14100,N_9882,N_11527);
nand U14101 (N_14101,N_11082,N_10416);
nor U14102 (N_14102,N_11097,N_11239);
or U14103 (N_14103,N_10408,N_10489);
or U14104 (N_14104,N_9091,N_11808);
and U14105 (N_14105,N_11931,N_9326);
nand U14106 (N_14106,N_10928,N_11235);
or U14107 (N_14107,N_10821,N_10314);
nor U14108 (N_14108,N_11647,N_9600);
nor U14109 (N_14109,N_10479,N_11108);
and U14110 (N_14110,N_10997,N_11590);
or U14111 (N_14111,N_10527,N_11795);
nor U14112 (N_14112,N_10599,N_9222);
nand U14113 (N_14113,N_9567,N_11158);
and U14114 (N_14114,N_10057,N_10531);
xnor U14115 (N_14115,N_11165,N_10448);
nand U14116 (N_14116,N_11148,N_10176);
or U14117 (N_14117,N_9318,N_10128);
and U14118 (N_14118,N_10697,N_9969);
nor U14119 (N_14119,N_9840,N_11445);
nor U14120 (N_14120,N_9722,N_9008);
nor U14121 (N_14121,N_10426,N_9044);
xor U14122 (N_14122,N_9938,N_10784);
or U14123 (N_14123,N_11808,N_9745);
and U14124 (N_14124,N_11503,N_11629);
and U14125 (N_14125,N_11265,N_9905);
and U14126 (N_14126,N_9712,N_9393);
xor U14127 (N_14127,N_10172,N_11822);
nor U14128 (N_14128,N_10899,N_9106);
or U14129 (N_14129,N_9607,N_10236);
xor U14130 (N_14130,N_11769,N_9546);
nand U14131 (N_14131,N_9099,N_11486);
nand U14132 (N_14132,N_9420,N_10803);
nand U14133 (N_14133,N_11725,N_10311);
nand U14134 (N_14134,N_11519,N_11701);
nand U14135 (N_14135,N_11241,N_11280);
xnor U14136 (N_14136,N_10030,N_10973);
and U14137 (N_14137,N_9114,N_9456);
nand U14138 (N_14138,N_10349,N_9796);
nand U14139 (N_14139,N_11887,N_9102);
nor U14140 (N_14140,N_10511,N_11231);
xnor U14141 (N_14141,N_11531,N_9093);
or U14142 (N_14142,N_11975,N_11332);
or U14143 (N_14143,N_10281,N_11425);
or U14144 (N_14144,N_9981,N_10015);
and U14145 (N_14145,N_9746,N_11126);
nand U14146 (N_14146,N_9144,N_9218);
xnor U14147 (N_14147,N_9913,N_10080);
and U14148 (N_14148,N_9401,N_10953);
nand U14149 (N_14149,N_11442,N_10877);
or U14150 (N_14150,N_9012,N_10616);
nor U14151 (N_14151,N_10783,N_9025);
or U14152 (N_14152,N_9931,N_9303);
or U14153 (N_14153,N_9063,N_9788);
nor U14154 (N_14154,N_10646,N_10864);
xor U14155 (N_14155,N_9384,N_10196);
nor U14156 (N_14156,N_9351,N_11382);
and U14157 (N_14157,N_11893,N_11303);
and U14158 (N_14158,N_11188,N_10595);
or U14159 (N_14159,N_9654,N_10658);
or U14160 (N_14160,N_10495,N_11424);
nor U14161 (N_14161,N_10511,N_9012);
or U14162 (N_14162,N_10627,N_10660);
or U14163 (N_14163,N_10687,N_10966);
xor U14164 (N_14164,N_10822,N_10476);
nand U14165 (N_14165,N_9959,N_9211);
and U14166 (N_14166,N_10352,N_9172);
nand U14167 (N_14167,N_10311,N_10532);
and U14168 (N_14168,N_10898,N_10853);
and U14169 (N_14169,N_9953,N_9221);
xnor U14170 (N_14170,N_9804,N_9840);
xnor U14171 (N_14171,N_9465,N_9749);
and U14172 (N_14172,N_9544,N_10325);
and U14173 (N_14173,N_10114,N_10783);
and U14174 (N_14174,N_11447,N_10702);
xor U14175 (N_14175,N_10081,N_9806);
nand U14176 (N_14176,N_11055,N_11809);
and U14177 (N_14177,N_11634,N_9576);
or U14178 (N_14178,N_10712,N_10170);
and U14179 (N_14179,N_11834,N_10068);
or U14180 (N_14180,N_9810,N_10582);
xnor U14181 (N_14181,N_11433,N_11567);
nand U14182 (N_14182,N_11408,N_11935);
nor U14183 (N_14183,N_11090,N_10588);
nor U14184 (N_14184,N_11823,N_11678);
or U14185 (N_14185,N_9867,N_10420);
nand U14186 (N_14186,N_9391,N_10806);
nand U14187 (N_14187,N_9452,N_10396);
nand U14188 (N_14188,N_10121,N_9042);
nand U14189 (N_14189,N_11139,N_11745);
or U14190 (N_14190,N_10653,N_9931);
nand U14191 (N_14191,N_11747,N_9664);
or U14192 (N_14192,N_11429,N_9786);
xor U14193 (N_14193,N_11749,N_10260);
nand U14194 (N_14194,N_11070,N_9783);
xor U14195 (N_14195,N_10844,N_9766);
or U14196 (N_14196,N_9513,N_9842);
or U14197 (N_14197,N_10736,N_9111);
xnor U14198 (N_14198,N_11099,N_10852);
nor U14199 (N_14199,N_11565,N_11176);
and U14200 (N_14200,N_9785,N_11944);
nand U14201 (N_14201,N_10748,N_9023);
nand U14202 (N_14202,N_9525,N_9920);
or U14203 (N_14203,N_11141,N_11210);
nor U14204 (N_14204,N_10844,N_9763);
nor U14205 (N_14205,N_11521,N_9371);
nand U14206 (N_14206,N_10422,N_11841);
and U14207 (N_14207,N_10110,N_10979);
and U14208 (N_14208,N_9283,N_10366);
and U14209 (N_14209,N_11835,N_10772);
xor U14210 (N_14210,N_11742,N_10149);
xor U14211 (N_14211,N_9827,N_11897);
or U14212 (N_14212,N_9647,N_11615);
nor U14213 (N_14213,N_11042,N_10672);
xor U14214 (N_14214,N_11057,N_9201);
and U14215 (N_14215,N_11359,N_10065);
nor U14216 (N_14216,N_10371,N_9170);
nand U14217 (N_14217,N_11534,N_10678);
nor U14218 (N_14218,N_9424,N_9777);
nor U14219 (N_14219,N_10562,N_10451);
and U14220 (N_14220,N_10833,N_9956);
and U14221 (N_14221,N_9369,N_9756);
nor U14222 (N_14222,N_9940,N_9950);
xor U14223 (N_14223,N_10477,N_11036);
xor U14224 (N_14224,N_9391,N_9471);
nor U14225 (N_14225,N_10373,N_9682);
and U14226 (N_14226,N_11698,N_10791);
nor U14227 (N_14227,N_9174,N_9965);
and U14228 (N_14228,N_10510,N_9098);
nor U14229 (N_14229,N_10932,N_9482);
and U14230 (N_14230,N_10498,N_9239);
and U14231 (N_14231,N_10686,N_10482);
xnor U14232 (N_14232,N_9758,N_11665);
and U14233 (N_14233,N_9741,N_11920);
and U14234 (N_14234,N_9608,N_10451);
xor U14235 (N_14235,N_11148,N_9493);
nor U14236 (N_14236,N_11012,N_10836);
xor U14237 (N_14237,N_11779,N_10206);
nor U14238 (N_14238,N_9903,N_11523);
or U14239 (N_14239,N_9376,N_10461);
nand U14240 (N_14240,N_11626,N_10718);
nand U14241 (N_14241,N_9548,N_11556);
nor U14242 (N_14242,N_9633,N_10701);
nor U14243 (N_14243,N_10495,N_10760);
nand U14244 (N_14244,N_9061,N_9751);
nor U14245 (N_14245,N_10560,N_9580);
nor U14246 (N_14246,N_9622,N_9640);
xor U14247 (N_14247,N_9310,N_11990);
nand U14248 (N_14248,N_10342,N_11054);
nand U14249 (N_14249,N_11782,N_11703);
and U14250 (N_14250,N_9298,N_9226);
and U14251 (N_14251,N_10333,N_10109);
and U14252 (N_14252,N_11191,N_11257);
nor U14253 (N_14253,N_10856,N_10801);
nor U14254 (N_14254,N_10765,N_9357);
nand U14255 (N_14255,N_11539,N_10780);
or U14256 (N_14256,N_10674,N_11137);
and U14257 (N_14257,N_9368,N_11311);
and U14258 (N_14258,N_11116,N_11054);
or U14259 (N_14259,N_9400,N_9025);
nand U14260 (N_14260,N_11460,N_9465);
or U14261 (N_14261,N_9836,N_11386);
xor U14262 (N_14262,N_10294,N_10212);
nor U14263 (N_14263,N_10174,N_11932);
xor U14264 (N_14264,N_10042,N_11863);
nor U14265 (N_14265,N_11624,N_9733);
nor U14266 (N_14266,N_10329,N_9161);
xor U14267 (N_14267,N_10543,N_11063);
or U14268 (N_14268,N_9644,N_11664);
nor U14269 (N_14269,N_9829,N_9891);
xor U14270 (N_14270,N_9821,N_10941);
and U14271 (N_14271,N_11904,N_11606);
or U14272 (N_14272,N_11077,N_10421);
nand U14273 (N_14273,N_11501,N_10841);
nor U14274 (N_14274,N_9379,N_11843);
and U14275 (N_14275,N_9631,N_10440);
or U14276 (N_14276,N_10284,N_9827);
or U14277 (N_14277,N_9883,N_9432);
and U14278 (N_14278,N_10351,N_9791);
xnor U14279 (N_14279,N_9712,N_10598);
and U14280 (N_14280,N_10850,N_9442);
xor U14281 (N_14281,N_10321,N_9028);
nand U14282 (N_14282,N_11300,N_11158);
or U14283 (N_14283,N_10587,N_11720);
or U14284 (N_14284,N_11628,N_11794);
and U14285 (N_14285,N_9381,N_10516);
nor U14286 (N_14286,N_11101,N_9203);
and U14287 (N_14287,N_10272,N_10879);
nand U14288 (N_14288,N_9987,N_10612);
or U14289 (N_14289,N_10685,N_11117);
nor U14290 (N_14290,N_9878,N_11070);
nand U14291 (N_14291,N_11041,N_9574);
nand U14292 (N_14292,N_11453,N_10846);
nor U14293 (N_14293,N_9591,N_10230);
xor U14294 (N_14294,N_9849,N_11270);
or U14295 (N_14295,N_11910,N_11684);
nand U14296 (N_14296,N_9415,N_10950);
xnor U14297 (N_14297,N_9065,N_11307);
nor U14298 (N_14298,N_9316,N_11672);
or U14299 (N_14299,N_9110,N_10028);
or U14300 (N_14300,N_10698,N_10996);
or U14301 (N_14301,N_9873,N_11121);
nor U14302 (N_14302,N_9180,N_11745);
nand U14303 (N_14303,N_11206,N_11048);
nand U14304 (N_14304,N_11998,N_10314);
xnor U14305 (N_14305,N_11408,N_9835);
or U14306 (N_14306,N_10001,N_9000);
nor U14307 (N_14307,N_10427,N_10330);
nand U14308 (N_14308,N_11838,N_11050);
and U14309 (N_14309,N_9410,N_11907);
xor U14310 (N_14310,N_9976,N_11179);
or U14311 (N_14311,N_11000,N_9789);
xor U14312 (N_14312,N_10051,N_9147);
xnor U14313 (N_14313,N_9881,N_10689);
or U14314 (N_14314,N_11797,N_9770);
and U14315 (N_14315,N_10056,N_9198);
xor U14316 (N_14316,N_10542,N_10194);
or U14317 (N_14317,N_9630,N_10727);
and U14318 (N_14318,N_11373,N_11219);
nand U14319 (N_14319,N_11997,N_10940);
nor U14320 (N_14320,N_9221,N_10292);
and U14321 (N_14321,N_10697,N_9807);
nand U14322 (N_14322,N_10292,N_9612);
nand U14323 (N_14323,N_10840,N_9446);
nand U14324 (N_14324,N_10728,N_10643);
or U14325 (N_14325,N_11569,N_11482);
nand U14326 (N_14326,N_11383,N_9650);
nor U14327 (N_14327,N_11951,N_11470);
or U14328 (N_14328,N_9813,N_11722);
or U14329 (N_14329,N_10417,N_9130);
or U14330 (N_14330,N_10414,N_9384);
nor U14331 (N_14331,N_11014,N_9798);
nand U14332 (N_14332,N_9050,N_9267);
nand U14333 (N_14333,N_10534,N_10589);
or U14334 (N_14334,N_9447,N_9835);
nor U14335 (N_14335,N_9776,N_11726);
xnor U14336 (N_14336,N_11543,N_11691);
nor U14337 (N_14337,N_11445,N_9241);
and U14338 (N_14338,N_10232,N_10850);
and U14339 (N_14339,N_10062,N_10582);
nor U14340 (N_14340,N_10607,N_9153);
nor U14341 (N_14341,N_11683,N_9702);
nand U14342 (N_14342,N_9047,N_11361);
and U14343 (N_14343,N_10092,N_11017);
or U14344 (N_14344,N_9263,N_10019);
or U14345 (N_14345,N_9402,N_10882);
nor U14346 (N_14346,N_9630,N_11921);
and U14347 (N_14347,N_9710,N_9662);
or U14348 (N_14348,N_11335,N_9425);
nand U14349 (N_14349,N_11297,N_10926);
xnor U14350 (N_14350,N_11859,N_9672);
or U14351 (N_14351,N_10416,N_10610);
xnor U14352 (N_14352,N_11564,N_11544);
or U14353 (N_14353,N_11650,N_9807);
nand U14354 (N_14354,N_11277,N_11424);
nor U14355 (N_14355,N_10181,N_9143);
xor U14356 (N_14356,N_9315,N_9202);
nand U14357 (N_14357,N_11732,N_10958);
nand U14358 (N_14358,N_11570,N_9203);
and U14359 (N_14359,N_10588,N_10044);
or U14360 (N_14360,N_9541,N_9906);
xnor U14361 (N_14361,N_11858,N_9865);
nand U14362 (N_14362,N_9242,N_11013);
nor U14363 (N_14363,N_9389,N_11943);
xnor U14364 (N_14364,N_10283,N_10127);
xor U14365 (N_14365,N_11931,N_10835);
nand U14366 (N_14366,N_9974,N_9609);
nand U14367 (N_14367,N_9227,N_10358);
nand U14368 (N_14368,N_11041,N_10209);
and U14369 (N_14369,N_11208,N_9558);
nor U14370 (N_14370,N_10592,N_11437);
or U14371 (N_14371,N_11259,N_11421);
nand U14372 (N_14372,N_11264,N_9679);
or U14373 (N_14373,N_11530,N_9567);
nand U14374 (N_14374,N_10180,N_10583);
xor U14375 (N_14375,N_10946,N_10623);
xor U14376 (N_14376,N_10338,N_9065);
or U14377 (N_14377,N_11827,N_9918);
xnor U14378 (N_14378,N_11786,N_9513);
xnor U14379 (N_14379,N_10492,N_9941);
and U14380 (N_14380,N_10124,N_11385);
xnor U14381 (N_14381,N_9990,N_9141);
or U14382 (N_14382,N_11189,N_11163);
nor U14383 (N_14383,N_10748,N_11965);
nand U14384 (N_14384,N_11812,N_10863);
nor U14385 (N_14385,N_9501,N_9865);
nand U14386 (N_14386,N_11374,N_9170);
nand U14387 (N_14387,N_9574,N_9980);
nand U14388 (N_14388,N_9715,N_11540);
nand U14389 (N_14389,N_9258,N_9737);
or U14390 (N_14390,N_11281,N_9262);
nor U14391 (N_14391,N_11338,N_10460);
nor U14392 (N_14392,N_9832,N_9450);
and U14393 (N_14393,N_9503,N_10960);
or U14394 (N_14394,N_10376,N_10676);
xnor U14395 (N_14395,N_9807,N_9867);
xnor U14396 (N_14396,N_10653,N_10537);
nand U14397 (N_14397,N_9246,N_10983);
or U14398 (N_14398,N_11404,N_11197);
xnor U14399 (N_14399,N_10698,N_11215);
nand U14400 (N_14400,N_11552,N_11764);
nor U14401 (N_14401,N_11794,N_9786);
nor U14402 (N_14402,N_10915,N_11503);
nand U14403 (N_14403,N_9723,N_10437);
nand U14404 (N_14404,N_9555,N_11021);
xor U14405 (N_14405,N_11451,N_11572);
nor U14406 (N_14406,N_11609,N_9116);
nand U14407 (N_14407,N_9452,N_9911);
xor U14408 (N_14408,N_9086,N_10436);
or U14409 (N_14409,N_11753,N_9269);
and U14410 (N_14410,N_9034,N_10401);
nor U14411 (N_14411,N_10370,N_9408);
and U14412 (N_14412,N_11273,N_9283);
xor U14413 (N_14413,N_9411,N_10987);
nor U14414 (N_14414,N_9974,N_9283);
nor U14415 (N_14415,N_11654,N_9748);
nor U14416 (N_14416,N_11465,N_11069);
nor U14417 (N_14417,N_11091,N_10337);
xnor U14418 (N_14418,N_11361,N_10883);
nor U14419 (N_14419,N_10641,N_9474);
nand U14420 (N_14420,N_10401,N_9996);
or U14421 (N_14421,N_10748,N_11791);
or U14422 (N_14422,N_11569,N_9562);
or U14423 (N_14423,N_10087,N_10592);
and U14424 (N_14424,N_10115,N_11537);
or U14425 (N_14425,N_10148,N_11900);
xor U14426 (N_14426,N_9037,N_9595);
nor U14427 (N_14427,N_9697,N_11439);
and U14428 (N_14428,N_10014,N_11487);
nand U14429 (N_14429,N_10111,N_9457);
xor U14430 (N_14430,N_11761,N_10016);
xor U14431 (N_14431,N_10769,N_11200);
and U14432 (N_14432,N_9503,N_10709);
xnor U14433 (N_14433,N_10856,N_11763);
nor U14434 (N_14434,N_10305,N_11040);
and U14435 (N_14435,N_9022,N_9311);
xor U14436 (N_14436,N_11385,N_11962);
and U14437 (N_14437,N_11668,N_10307);
or U14438 (N_14438,N_10104,N_10126);
xor U14439 (N_14439,N_9796,N_10482);
or U14440 (N_14440,N_10350,N_11778);
and U14441 (N_14441,N_10481,N_11178);
nor U14442 (N_14442,N_10941,N_9254);
or U14443 (N_14443,N_9670,N_10169);
or U14444 (N_14444,N_11052,N_10235);
nor U14445 (N_14445,N_10314,N_9228);
nand U14446 (N_14446,N_9362,N_10302);
and U14447 (N_14447,N_9690,N_10534);
xnor U14448 (N_14448,N_11230,N_9464);
or U14449 (N_14449,N_11116,N_10306);
nor U14450 (N_14450,N_9973,N_11095);
or U14451 (N_14451,N_9772,N_9712);
nand U14452 (N_14452,N_10266,N_10022);
or U14453 (N_14453,N_10947,N_9005);
xor U14454 (N_14454,N_10939,N_10325);
nor U14455 (N_14455,N_11234,N_10567);
nand U14456 (N_14456,N_10027,N_10102);
nor U14457 (N_14457,N_10454,N_10910);
and U14458 (N_14458,N_10926,N_9578);
and U14459 (N_14459,N_9846,N_11613);
nand U14460 (N_14460,N_9469,N_11507);
or U14461 (N_14461,N_10868,N_11980);
xor U14462 (N_14462,N_10558,N_11666);
and U14463 (N_14463,N_11177,N_11702);
and U14464 (N_14464,N_9489,N_11634);
and U14465 (N_14465,N_11860,N_9941);
nor U14466 (N_14466,N_9167,N_11165);
nand U14467 (N_14467,N_9299,N_9304);
or U14468 (N_14468,N_10422,N_10065);
and U14469 (N_14469,N_11799,N_10929);
xnor U14470 (N_14470,N_10018,N_10450);
nand U14471 (N_14471,N_10460,N_9394);
nor U14472 (N_14472,N_11063,N_9042);
and U14473 (N_14473,N_11550,N_11162);
and U14474 (N_14474,N_9850,N_10293);
or U14475 (N_14475,N_10430,N_10194);
nor U14476 (N_14476,N_10127,N_11504);
or U14477 (N_14477,N_11990,N_11886);
and U14478 (N_14478,N_11407,N_10778);
nand U14479 (N_14479,N_10187,N_9414);
xnor U14480 (N_14480,N_9147,N_9770);
and U14481 (N_14481,N_11118,N_10512);
and U14482 (N_14482,N_11503,N_10275);
nand U14483 (N_14483,N_11111,N_11438);
or U14484 (N_14484,N_11087,N_9791);
or U14485 (N_14485,N_11684,N_9261);
and U14486 (N_14486,N_11088,N_11191);
nand U14487 (N_14487,N_10026,N_9555);
or U14488 (N_14488,N_11960,N_11077);
nor U14489 (N_14489,N_9261,N_9836);
or U14490 (N_14490,N_11870,N_9282);
or U14491 (N_14491,N_9075,N_10569);
and U14492 (N_14492,N_10417,N_11395);
nand U14493 (N_14493,N_11923,N_11730);
nor U14494 (N_14494,N_11979,N_9957);
nand U14495 (N_14495,N_10418,N_9028);
xor U14496 (N_14496,N_10141,N_9627);
nand U14497 (N_14497,N_9654,N_9117);
and U14498 (N_14498,N_11851,N_9407);
xor U14499 (N_14499,N_11237,N_11520);
nand U14500 (N_14500,N_10108,N_9235);
and U14501 (N_14501,N_9387,N_9518);
nor U14502 (N_14502,N_11643,N_11620);
nand U14503 (N_14503,N_9416,N_10762);
xor U14504 (N_14504,N_11564,N_11462);
and U14505 (N_14505,N_10763,N_10674);
xor U14506 (N_14506,N_11792,N_9071);
nor U14507 (N_14507,N_10568,N_9841);
nand U14508 (N_14508,N_10557,N_11514);
xor U14509 (N_14509,N_9847,N_11739);
nor U14510 (N_14510,N_10266,N_9402);
nand U14511 (N_14511,N_9564,N_9290);
nor U14512 (N_14512,N_10737,N_10638);
xnor U14513 (N_14513,N_10989,N_10529);
and U14514 (N_14514,N_10006,N_11854);
nand U14515 (N_14515,N_9985,N_11567);
xor U14516 (N_14516,N_10476,N_9389);
xnor U14517 (N_14517,N_9629,N_11435);
or U14518 (N_14518,N_11971,N_10608);
nand U14519 (N_14519,N_9643,N_10834);
or U14520 (N_14520,N_10453,N_9179);
nor U14521 (N_14521,N_10112,N_10066);
nand U14522 (N_14522,N_11645,N_10229);
nand U14523 (N_14523,N_11149,N_11041);
nor U14524 (N_14524,N_10236,N_9705);
nand U14525 (N_14525,N_11798,N_10750);
and U14526 (N_14526,N_9453,N_10976);
xor U14527 (N_14527,N_10032,N_11399);
nor U14528 (N_14528,N_11042,N_10758);
or U14529 (N_14529,N_10096,N_10365);
and U14530 (N_14530,N_11479,N_9985);
xnor U14531 (N_14531,N_11559,N_9894);
xnor U14532 (N_14532,N_10620,N_9261);
xor U14533 (N_14533,N_11933,N_10517);
nand U14534 (N_14534,N_10484,N_11401);
xnor U14535 (N_14535,N_11582,N_9458);
or U14536 (N_14536,N_9177,N_10703);
and U14537 (N_14537,N_11998,N_11858);
xor U14538 (N_14538,N_10425,N_9205);
nand U14539 (N_14539,N_11591,N_11350);
or U14540 (N_14540,N_10963,N_10123);
and U14541 (N_14541,N_10750,N_9326);
and U14542 (N_14542,N_11640,N_11227);
and U14543 (N_14543,N_10952,N_11637);
nand U14544 (N_14544,N_9948,N_11843);
nor U14545 (N_14545,N_9297,N_10951);
and U14546 (N_14546,N_11612,N_9931);
and U14547 (N_14547,N_11735,N_9240);
nor U14548 (N_14548,N_9929,N_11610);
nand U14549 (N_14549,N_10690,N_9147);
nor U14550 (N_14550,N_9887,N_10746);
xnor U14551 (N_14551,N_11317,N_9282);
xor U14552 (N_14552,N_9459,N_10802);
xnor U14553 (N_14553,N_9227,N_9644);
nor U14554 (N_14554,N_11307,N_9772);
or U14555 (N_14555,N_10416,N_10866);
nand U14556 (N_14556,N_10256,N_9162);
and U14557 (N_14557,N_11074,N_9719);
nand U14558 (N_14558,N_11793,N_10180);
xor U14559 (N_14559,N_11965,N_9591);
or U14560 (N_14560,N_10845,N_11053);
and U14561 (N_14561,N_11885,N_10575);
xnor U14562 (N_14562,N_10358,N_10958);
nand U14563 (N_14563,N_10433,N_10786);
nor U14564 (N_14564,N_9428,N_10634);
xnor U14565 (N_14565,N_10275,N_10173);
xnor U14566 (N_14566,N_11445,N_9689);
or U14567 (N_14567,N_10837,N_10454);
nor U14568 (N_14568,N_9621,N_11639);
or U14569 (N_14569,N_9497,N_9125);
nand U14570 (N_14570,N_10761,N_11627);
nor U14571 (N_14571,N_10268,N_11585);
xor U14572 (N_14572,N_11260,N_10402);
or U14573 (N_14573,N_10388,N_9164);
and U14574 (N_14574,N_10441,N_9354);
nor U14575 (N_14575,N_11967,N_10715);
or U14576 (N_14576,N_11308,N_11496);
nand U14577 (N_14577,N_11527,N_9610);
or U14578 (N_14578,N_11074,N_9762);
xor U14579 (N_14579,N_11431,N_10188);
nand U14580 (N_14580,N_11182,N_10375);
or U14581 (N_14581,N_10363,N_11671);
and U14582 (N_14582,N_11558,N_9592);
nor U14583 (N_14583,N_9123,N_11703);
and U14584 (N_14584,N_9602,N_9426);
xnor U14585 (N_14585,N_9098,N_10093);
and U14586 (N_14586,N_9530,N_11034);
xnor U14587 (N_14587,N_10388,N_9701);
xnor U14588 (N_14588,N_10463,N_10211);
xor U14589 (N_14589,N_11833,N_10346);
nor U14590 (N_14590,N_10522,N_9412);
nand U14591 (N_14591,N_10141,N_11524);
and U14592 (N_14592,N_11639,N_11360);
or U14593 (N_14593,N_9955,N_9474);
and U14594 (N_14594,N_11432,N_10743);
nor U14595 (N_14595,N_10006,N_10543);
nor U14596 (N_14596,N_11803,N_9566);
nand U14597 (N_14597,N_10831,N_10709);
nand U14598 (N_14598,N_9127,N_9414);
and U14599 (N_14599,N_10768,N_9648);
nor U14600 (N_14600,N_10907,N_11235);
and U14601 (N_14601,N_11499,N_10041);
and U14602 (N_14602,N_11704,N_11968);
and U14603 (N_14603,N_9456,N_10823);
and U14604 (N_14604,N_11978,N_10844);
nor U14605 (N_14605,N_9845,N_11338);
or U14606 (N_14606,N_9493,N_11992);
nand U14607 (N_14607,N_11637,N_10028);
xnor U14608 (N_14608,N_9199,N_9360);
xor U14609 (N_14609,N_11978,N_9760);
or U14610 (N_14610,N_9092,N_9121);
nor U14611 (N_14611,N_11645,N_11734);
nor U14612 (N_14612,N_9757,N_10359);
or U14613 (N_14613,N_11280,N_9308);
or U14614 (N_14614,N_9627,N_10151);
nor U14615 (N_14615,N_10139,N_10545);
xor U14616 (N_14616,N_10487,N_11083);
xnor U14617 (N_14617,N_10792,N_9358);
or U14618 (N_14618,N_11269,N_9761);
nor U14619 (N_14619,N_9753,N_9421);
xor U14620 (N_14620,N_9116,N_9761);
nor U14621 (N_14621,N_9002,N_10273);
or U14622 (N_14622,N_10898,N_10193);
xor U14623 (N_14623,N_9592,N_10389);
nor U14624 (N_14624,N_9877,N_9032);
or U14625 (N_14625,N_9560,N_11355);
nand U14626 (N_14626,N_11945,N_11687);
or U14627 (N_14627,N_9285,N_11376);
xnor U14628 (N_14628,N_9440,N_9657);
nand U14629 (N_14629,N_11121,N_10371);
xor U14630 (N_14630,N_10322,N_10578);
nand U14631 (N_14631,N_11193,N_9533);
nor U14632 (N_14632,N_9679,N_10999);
nor U14633 (N_14633,N_9860,N_10696);
or U14634 (N_14634,N_10306,N_10126);
and U14635 (N_14635,N_9010,N_11728);
xnor U14636 (N_14636,N_10387,N_9531);
nor U14637 (N_14637,N_10253,N_11327);
nand U14638 (N_14638,N_9948,N_10259);
or U14639 (N_14639,N_9355,N_9594);
nor U14640 (N_14640,N_10849,N_11265);
nand U14641 (N_14641,N_9577,N_10554);
nor U14642 (N_14642,N_11892,N_9026);
nor U14643 (N_14643,N_11199,N_10962);
nand U14644 (N_14644,N_10471,N_11405);
nor U14645 (N_14645,N_10449,N_10371);
and U14646 (N_14646,N_10059,N_9458);
xnor U14647 (N_14647,N_9447,N_11554);
xor U14648 (N_14648,N_10982,N_11802);
or U14649 (N_14649,N_11446,N_9928);
nor U14650 (N_14650,N_9089,N_9388);
and U14651 (N_14651,N_10701,N_10688);
xnor U14652 (N_14652,N_9051,N_10571);
and U14653 (N_14653,N_11087,N_10447);
xnor U14654 (N_14654,N_10854,N_10152);
nand U14655 (N_14655,N_11197,N_10453);
or U14656 (N_14656,N_11804,N_11015);
and U14657 (N_14657,N_9947,N_10351);
xnor U14658 (N_14658,N_9435,N_9731);
nand U14659 (N_14659,N_10860,N_11070);
nand U14660 (N_14660,N_11427,N_10710);
xnor U14661 (N_14661,N_11037,N_10825);
nand U14662 (N_14662,N_9931,N_9654);
and U14663 (N_14663,N_10522,N_9770);
nand U14664 (N_14664,N_9609,N_10330);
or U14665 (N_14665,N_11739,N_10454);
nor U14666 (N_14666,N_9502,N_11546);
and U14667 (N_14667,N_11188,N_11052);
and U14668 (N_14668,N_9477,N_10489);
nor U14669 (N_14669,N_9976,N_9140);
nor U14670 (N_14670,N_11411,N_9072);
nor U14671 (N_14671,N_10213,N_9201);
and U14672 (N_14672,N_10215,N_9182);
nor U14673 (N_14673,N_9492,N_9413);
or U14674 (N_14674,N_11183,N_11111);
nand U14675 (N_14675,N_11612,N_11723);
or U14676 (N_14676,N_11123,N_9007);
and U14677 (N_14677,N_9280,N_9904);
xnor U14678 (N_14678,N_11448,N_10120);
nor U14679 (N_14679,N_9228,N_11995);
or U14680 (N_14680,N_9046,N_10568);
xnor U14681 (N_14681,N_10486,N_11683);
and U14682 (N_14682,N_11693,N_10125);
and U14683 (N_14683,N_10554,N_11582);
xor U14684 (N_14684,N_10293,N_9510);
xnor U14685 (N_14685,N_11435,N_9007);
nor U14686 (N_14686,N_10819,N_9245);
nand U14687 (N_14687,N_9709,N_10218);
xor U14688 (N_14688,N_9784,N_11821);
and U14689 (N_14689,N_11210,N_9666);
xnor U14690 (N_14690,N_11826,N_10147);
nor U14691 (N_14691,N_11456,N_10679);
and U14692 (N_14692,N_9076,N_11959);
or U14693 (N_14693,N_9461,N_11214);
nor U14694 (N_14694,N_11747,N_11592);
or U14695 (N_14695,N_11680,N_10740);
xnor U14696 (N_14696,N_10534,N_10616);
or U14697 (N_14697,N_11114,N_11414);
or U14698 (N_14698,N_9258,N_10704);
xor U14699 (N_14699,N_11491,N_9626);
and U14700 (N_14700,N_11397,N_9340);
and U14701 (N_14701,N_9802,N_11086);
and U14702 (N_14702,N_9847,N_9247);
and U14703 (N_14703,N_9136,N_11074);
nor U14704 (N_14704,N_11005,N_10237);
or U14705 (N_14705,N_11074,N_9674);
xnor U14706 (N_14706,N_11854,N_10620);
nand U14707 (N_14707,N_9804,N_9723);
or U14708 (N_14708,N_9288,N_9538);
and U14709 (N_14709,N_11705,N_9821);
nand U14710 (N_14710,N_10353,N_9126);
xnor U14711 (N_14711,N_9260,N_10067);
xnor U14712 (N_14712,N_9215,N_10913);
nand U14713 (N_14713,N_11664,N_10779);
nand U14714 (N_14714,N_10963,N_10927);
nor U14715 (N_14715,N_10920,N_10484);
nand U14716 (N_14716,N_11818,N_9267);
nand U14717 (N_14717,N_9389,N_11690);
xnor U14718 (N_14718,N_10375,N_10371);
xnor U14719 (N_14719,N_9267,N_10995);
nand U14720 (N_14720,N_11525,N_10884);
nor U14721 (N_14721,N_11513,N_11460);
xor U14722 (N_14722,N_9594,N_9589);
and U14723 (N_14723,N_11274,N_9600);
nand U14724 (N_14724,N_10441,N_10307);
and U14725 (N_14725,N_9236,N_11935);
and U14726 (N_14726,N_10090,N_10178);
xnor U14727 (N_14727,N_10843,N_9679);
nor U14728 (N_14728,N_9007,N_11641);
and U14729 (N_14729,N_11088,N_10278);
or U14730 (N_14730,N_10677,N_10810);
and U14731 (N_14731,N_9898,N_11439);
nand U14732 (N_14732,N_10246,N_10423);
or U14733 (N_14733,N_9098,N_11992);
nor U14734 (N_14734,N_11108,N_10735);
xnor U14735 (N_14735,N_9675,N_10116);
and U14736 (N_14736,N_11069,N_10078);
and U14737 (N_14737,N_10612,N_11336);
and U14738 (N_14738,N_9772,N_10093);
or U14739 (N_14739,N_11017,N_11310);
or U14740 (N_14740,N_11494,N_9012);
and U14741 (N_14741,N_9217,N_11088);
nand U14742 (N_14742,N_9621,N_9065);
xor U14743 (N_14743,N_9261,N_11298);
xnor U14744 (N_14744,N_11948,N_11723);
nand U14745 (N_14745,N_9471,N_10569);
nor U14746 (N_14746,N_10983,N_10584);
or U14747 (N_14747,N_9315,N_10957);
nor U14748 (N_14748,N_11745,N_11741);
nor U14749 (N_14749,N_9142,N_10780);
nor U14750 (N_14750,N_9131,N_9051);
and U14751 (N_14751,N_10769,N_11043);
and U14752 (N_14752,N_9414,N_9831);
xnor U14753 (N_14753,N_9017,N_11626);
nand U14754 (N_14754,N_10652,N_9069);
xor U14755 (N_14755,N_9248,N_11592);
xnor U14756 (N_14756,N_9859,N_11958);
or U14757 (N_14757,N_11179,N_11675);
and U14758 (N_14758,N_10038,N_9532);
and U14759 (N_14759,N_11180,N_11191);
xnor U14760 (N_14760,N_11520,N_9847);
nor U14761 (N_14761,N_11640,N_11202);
and U14762 (N_14762,N_11539,N_10910);
xor U14763 (N_14763,N_9581,N_10894);
xor U14764 (N_14764,N_10907,N_10396);
or U14765 (N_14765,N_10700,N_9523);
xor U14766 (N_14766,N_10471,N_10367);
xnor U14767 (N_14767,N_11431,N_11839);
and U14768 (N_14768,N_9963,N_10299);
nor U14769 (N_14769,N_10804,N_9719);
or U14770 (N_14770,N_9148,N_9452);
nor U14771 (N_14771,N_11255,N_9960);
nor U14772 (N_14772,N_11632,N_9746);
or U14773 (N_14773,N_10439,N_11104);
and U14774 (N_14774,N_10153,N_9548);
and U14775 (N_14775,N_11682,N_11020);
and U14776 (N_14776,N_11849,N_10072);
nor U14777 (N_14777,N_11189,N_10391);
or U14778 (N_14778,N_11252,N_11402);
and U14779 (N_14779,N_10380,N_10634);
nor U14780 (N_14780,N_11052,N_10229);
xor U14781 (N_14781,N_9829,N_10693);
nand U14782 (N_14782,N_9878,N_9006);
nor U14783 (N_14783,N_10189,N_9624);
nand U14784 (N_14784,N_11211,N_10045);
xnor U14785 (N_14785,N_10066,N_11356);
and U14786 (N_14786,N_10301,N_11049);
nor U14787 (N_14787,N_11748,N_9625);
or U14788 (N_14788,N_9386,N_9652);
and U14789 (N_14789,N_10632,N_9120);
or U14790 (N_14790,N_11302,N_10772);
nor U14791 (N_14791,N_11841,N_9686);
nor U14792 (N_14792,N_11592,N_10355);
nand U14793 (N_14793,N_9812,N_10088);
nand U14794 (N_14794,N_9568,N_9948);
xnor U14795 (N_14795,N_9394,N_9292);
nor U14796 (N_14796,N_9602,N_10142);
and U14797 (N_14797,N_11436,N_11094);
nand U14798 (N_14798,N_11419,N_10456);
or U14799 (N_14799,N_11583,N_11440);
nor U14800 (N_14800,N_9431,N_9381);
nand U14801 (N_14801,N_10923,N_11456);
and U14802 (N_14802,N_11808,N_10043);
and U14803 (N_14803,N_9943,N_11140);
xor U14804 (N_14804,N_10221,N_10447);
and U14805 (N_14805,N_11438,N_9727);
and U14806 (N_14806,N_10956,N_11863);
and U14807 (N_14807,N_10527,N_11702);
or U14808 (N_14808,N_11821,N_10673);
nor U14809 (N_14809,N_11139,N_11491);
xor U14810 (N_14810,N_9196,N_10281);
and U14811 (N_14811,N_11230,N_10695);
and U14812 (N_14812,N_10213,N_9657);
nor U14813 (N_14813,N_10671,N_11151);
and U14814 (N_14814,N_10608,N_9776);
and U14815 (N_14815,N_11642,N_11755);
or U14816 (N_14816,N_10208,N_9044);
or U14817 (N_14817,N_10305,N_11192);
and U14818 (N_14818,N_11445,N_10243);
or U14819 (N_14819,N_11205,N_11701);
and U14820 (N_14820,N_11996,N_11625);
xor U14821 (N_14821,N_10771,N_9688);
nor U14822 (N_14822,N_9364,N_10422);
and U14823 (N_14823,N_11389,N_11192);
and U14824 (N_14824,N_10075,N_11167);
nand U14825 (N_14825,N_10643,N_10770);
and U14826 (N_14826,N_11637,N_11851);
xnor U14827 (N_14827,N_10762,N_11503);
or U14828 (N_14828,N_11174,N_10369);
or U14829 (N_14829,N_11857,N_11183);
and U14830 (N_14830,N_10976,N_10926);
nor U14831 (N_14831,N_11859,N_9642);
or U14832 (N_14832,N_10209,N_11638);
or U14833 (N_14833,N_10338,N_10247);
xnor U14834 (N_14834,N_10106,N_9370);
xor U14835 (N_14835,N_11696,N_9383);
or U14836 (N_14836,N_9403,N_9950);
nor U14837 (N_14837,N_9444,N_9854);
and U14838 (N_14838,N_11567,N_9996);
nand U14839 (N_14839,N_10708,N_9505);
nand U14840 (N_14840,N_10290,N_11814);
xor U14841 (N_14841,N_9581,N_11172);
and U14842 (N_14842,N_10730,N_10856);
and U14843 (N_14843,N_10959,N_11972);
xnor U14844 (N_14844,N_10655,N_11781);
nand U14845 (N_14845,N_11377,N_10208);
and U14846 (N_14846,N_9077,N_11528);
or U14847 (N_14847,N_10551,N_9089);
and U14848 (N_14848,N_10295,N_10325);
nor U14849 (N_14849,N_9113,N_11898);
or U14850 (N_14850,N_9323,N_11925);
or U14851 (N_14851,N_11265,N_9143);
or U14852 (N_14852,N_9296,N_10766);
and U14853 (N_14853,N_10290,N_11083);
nor U14854 (N_14854,N_9652,N_10197);
xor U14855 (N_14855,N_10265,N_10586);
or U14856 (N_14856,N_9240,N_11332);
nand U14857 (N_14857,N_9585,N_11638);
and U14858 (N_14858,N_10115,N_10130);
or U14859 (N_14859,N_11820,N_10166);
nor U14860 (N_14860,N_9084,N_9892);
xnor U14861 (N_14861,N_11018,N_11056);
and U14862 (N_14862,N_11015,N_9072);
xor U14863 (N_14863,N_11474,N_10466);
or U14864 (N_14864,N_10535,N_10049);
nand U14865 (N_14865,N_11700,N_9778);
nor U14866 (N_14866,N_11819,N_9007);
nand U14867 (N_14867,N_9700,N_11587);
and U14868 (N_14868,N_11806,N_10196);
xnor U14869 (N_14869,N_11492,N_9874);
nand U14870 (N_14870,N_9072,N_11067);
nand U14871 (N_14871,N_11820,N_10605);
or U14872 (N_14872,N_11290,N_11232);
or U14873 (N_14873,N_10403,N_9707);
xnor U14874 (N_14874,N_10616,N_11639);
and U14875 (N_14875,N_11340,N_11448);
or U14876 (N_14876,N_9420,N_9238);
and U14877 (N_14877,N_10553,N_10643);
and U14878 (N_14878,N_10529,N_10727);
or U14879 (N_14879,N_10039,N_11358);
nand U14880 (N_14880,N_10682,N_10012);
nand U14881 (N_14881,N_9963,N_9393);
xor U14882 (N_14882,N_10841,N_10859);
or U14883 (N_14883,N_9814,N_10015);
or U14884 (N_14884,N_9886,N_11399);
and U14885 (N_14885,N_11028,N_9926);
xor U14886 (N_14886,N_10614,N_11986);
nor U14887 (N_14887,N_10676,N_10015);
xnor U14888 (N_14888,N_9851,N_10917);
xor U14889 (N_14889,N_9855,N_10090);
xor U14890 (N_14890,N_11316,N_11577);
nor U14891 (N_14891,N_11289,N_10744);
nand U14892 (N_14892,N_9201,N_10517);
nor U14893 (N_14893,N_9127,N_9797);
and U14894 (N_14894,N_9583,N_11564);
nor U14895 (N_14895,N_9721,N_9369);
and U14896 (N_14896,N_10073,N_10377);
xor U14897 (N_14897,N_10537,N_10268);
nand U14898 (N_14898,N_9944,N_9537);
nor U14899 (N_14899,N_10863,N_11938);
and U14900 (N_14900,N_11173,N_11071);
xnor U14901 (N_14901,N_11540,N_11512);
nand U14902 (N_14902,N_10190,N_9142);
or U14903 (N_14903,N_9532,N_10381);
and U14904 (N_14904,N_11142,N_10441);
or U14905 (N_14905,N_9522,N_10746);
or U14906 (N_14906,N_11537,N_10353);
xor U14907 (N_14907,N_9465,N_9307);
or U14908 (N_14908,N_9105,N_10847);
nand U14909 (N_14909,N_9424,N_11089);
xnor U14910 (N_14910,N_11559,N_9204);
and U14911 (N_14911,N_11848,N_10499);
xor U14912 (N_14912,N_11197,N_11158);
and U14913 (N_14913,N_11112,N_10913);
or U14914 (N_14914,N_11199,N_9374);
nand U14915 (N_14915,N_11514,N_11745);
and U14916 (N_14916,N_9834,N_10800);
nand U14917 (N_14917,N_10324,N_10628);
nor U14918 (N_14918,N_9193,N_11453);
nor U14919 (N_14919,N_11196,N_10318);
xnor U14920 (N_14920,N_11343,N_10294);
or U14921 (N_14921,N_10443,N_10015);
and U14922 (N_14922,N_9267,N_10302);
xnor U14923 (N_14923,N_10856,N_9769);
and U14924 (N_14924,N_11973,N_10308);
nor U14925 (N_14925,N_11021,N_10710);
nand U14926 (N_14926,N_9246,N_9265);
and U14927 (N_14927,N_11594,N_10878);
and U14928 (N_14928,N_11802,N_10346);
and U14929 (N_14929,N_10784,N_9718);
xnor U14930 (N_14930,N_11206,N_11813);
nor U14931 (N_14931,N_10015,N_9884);
nand U14932 (N_14932,N_10258,N_11178);
nor U14933 (N_14933,N_11777,N_10081);
nand U14934 (N_14934,N_11060,N_11667);
nand U14935 (N_14935,N_10816,N_11715);
nor U14936 (N_14936,N_10647,N_10596);
nand U14937 (N_14937,N_10057,N_10640);
xnor U14938 (N_14938,N_9699,N_11577);
xor U14939 (N_14939,N_11330,N_9064);
xnor U14940 (N_14940,N_9798,N_10837);
and U14941 (N_14941,N_11069,N_11542);
or U14942 (N_14942,N_11369,N_11541);
xor U14943 (N_14943,N_9418,N_11792);
nand U14944 (N_14944,N_11343,N_11544);
and U14945 (N_14945,N_11892,N_11087);
and U14946 (N_14946,N_11033,N_9241);
nor U14947 (N_14947,N_10183,N_9506);
nor U14948 (N_14948,N_9201,N_9362);
nand U14949 (N_14949,N_9242,N_9695);
and U14950 (N_14950,N_10146,N_9447);
or U14951 (N_14951,N_9028,N_9052);
nor U14952 (N_14952,N_10159,N_10493);
nand U14953 (N_14953,N_10413,N_9885);
nand U14954 (N_14954,N_9174,N_11278);
or U14955 (N_14955,N_10255,N_10144);
xor U14956 (N_14956,N_10644,N_11240);
xnor U14957 (N_14957,N_11856,N_9521);
xnor U14958 (N_14958,N_10277,N_9570);
nor U14959 (N_14959,N_10447,N_10131);
and U14960 (N_14960,N_10450,N_11166);
and U14961 (N_14961,N_11262,N_10779);
or U14962 (N_14962,N_10718,N_10810);
or U14963 (N_14963,N_11606,N_11965);
xnor U14964 (N_14964,N_11444,N_11682);
and U14965 (N_14965,N_9972,N_9811);
or U14966 (N_14966,N_10897,N_9687);
xnor U14967 (N_14967,N_11353,N_11071);
or U14968 (N_14968,N_11867,N_9367);
or U14969 (N_14969,N_9853,N_11817);
xor U14970 (N_14970,N_10883,N_9575);
and U14971 (N_14971,N_9774,N_9912);
xor U14972 (N_14972,N_10818,N_9519);
xor U14973 (N_14973,N_9514,N_10139);
or U14974 (N_14974,N_10660,N_9836);
xor U14975 (N_14975,N_9674,N_10945);
nand U14976 (N_14976,N_9341,N_10536);
nand U14977 (N_14977,N_10669,N_9510);
or U14978 (N_14978,N_10958,N_10471);
or U14979 (N_14979,N_11373,N_9536);
or U14980 (N_14980,N_9889,N_9075);
nor U14981 (N_14981,N_9480,N_10528);
or U14982 (N_14982,N_11075,N_11339);
xnor U14983 (N_14983,N_10117,N_10429);
or U14984 (N_14984,N_11260,N_9317);
nand U14985 (N_14985,N_9512,N_9329);
nand U14986 (N_14986,N_9616,N_11815);
nor U14987 (N_14987,N_9006,N_9606);
nand U14988 (N_14988,N_11266,N_10205);
nand U14989 (N_14989,N_11588,N_9261);
nand U14990 (N_14990,N_9993,N_9806);
and U14991 (N_14991,N_11505,N_10172);
xor U14992 (N_14992,N_11601,N_9584);
or U14993 (N_14993,N_10109,N_9294);
xor U14994 (N_14994,N_10304,N_11894);
nand U14995 (N_14995,N_9076,N_11278);
xnor U14996 (N_14996,N_11192,N_9323);
xnor U14997 (N_14997,N_9183,N_10504);
and U14998 (N_14998,N_10278,N_10181);
xor U14999 (N_14999,N_9942,N_11249);
or U15000 (N_15000,N_13205,N_12439);
nor U15001 (N_15001,N_13678,N_13174);
and U15002 (N_15002,N_13418,N_13777);
or U15003 (N_15003,N_13364,N_13389);
or U15004 (N_15004,N_12584,N_14996);
and U15005 (N_15005,N_13889,N_13791);
nor U15006 (N_15006,N_13692,N_13453);
or U15007 (N_15007,N_12437,N_13977);
nand U15008 (N_15008,N_14689,N_13461);
nor U15009 (N_15009,N_14869,N_12246);
nand U15010 (N_15010,N_12065,N_12184);
or U15011 (N_15011,N_14659,N_13387);
nand U15012 (N_15012,N_14178,N_13535);
or U15013 (N_15013,N_12374,N_13481);
nor U15014 (N_15014,N_14862,N_14025);
and U15015 (N_15015,N_12064,N_12669);
nor U15016 (N_15016,N_13573,N_14077);
nor U15017 (N_15017,N_13542,N_14079);
xnor U15018 (N_15018,N_12705,N_13508);
nor U15019 (N_15019,N_13798,N_13486);
or U15020 (N_15020,N_12706,N_12476);
or U15021 (N_15021,N_14492,N_14523);
nor U15022 (N_15022,N_13820,N_14486);
nor U15023 (N_15023,N_13636,N_14738);
and U15024 (N_15024,N_14274,N_13865);
nor U15025 (N_15025,N_13496,N_13804);
xor U15026 (N_15026,N_12166,N_14095);
nor U15027 (N_15027,N_13328,N_13623);
nand U15028 (N_15028,N_12906,N_13843);
or U15029 (N_15029,N_14709,N_14962);
or U15030 (N_15030,N_14594,N_12487);
xor U15031 (N_15031,N_12051,N_13303);
nor U15032 (N_15032,N_13849,N_13994);
nand U15033 (N_15033,N_12574,N_13634);
nor U15034 (N_15034,N_13464,N_14515);
xor U15035 (N_15035,N_14699,N_12638);
and U15036 (N_15036,N_13909,N_12348);
xnor U15037 (N_15037,N_12308,N_12038);
and U15038 (N_15038,N_13579,N_13908);
nor U15039 (N_15039,N_13093,N_13781);
nand U15040 (N_15040,N_13503,N_12471);
and U15041 (N_15041,N_12355,N_14859);
nand U15042 (N_15042,N_12548,N_12769);
and U15043 (N_15043,N_13583,N_13322);
and U15044 (N_15044,N_13026,N_12729);
or U15045 (N_15045,N_12104,N_14624);
nor U15046 (N_15046,N_14401,N_12014);
nand U15047 (N_15047,N_13317,N_13152);
nor U15048 (N_15048,N_12561,N_12273);
nor U15049 (N_15049,N_12863,N_14987);
nor U15050 (N_15050,N_14972,N_13089);
nand U15051 (N_15051,N_12956,N_12389);
and U15052 (N_15052,N_13731,N_12525);
nor U15053 (N_15053,N_13880,N_12690);
nand U15054 (N_15054,N_14309,N_14468);
xor U15055 (N_15055,N_13680,N_12429);
nor U15056 (N_15056,N_14549,N_12187);
or U15057 (N_15057,N_13431,N_13578);
nand U15058 (N_15058,N_13287,N_13188);
and U15059 (N_15059,N_12327,N_13939);
nand U15060 (N_15060,N_13885,N_12028);
xor U15061 (N_15061,N_12054,N_14616);
nor U15062 (N_15062,N_12459,N_13073);
xnor U15063 (N_15063,N_12275,N_12245);
xnor U15064 (N_15064,N_14123,N_14392);
nand U15065 (N_15065,N_13710,N_14982);
and U15066 (N_15066,N_14342,N_12617);
xnor U15067 (N_15067,N_12891,N_14819);
and U15068 (N_15068,N_12042,N_12504);
and U15069 (N_15069,N_13297,N_13639);
and U15070 (N_15070,N_13851,N_12277);
nor U15071 (N_15071,N_14881,N_14787);
nand U15072 (N_15072,N_13752,N_12711);
and U15073 (N_15073,N_13513,N_12077);
xnor U15074 (N_15074,N_12281,N_14225);
xnor U15075 (N_15075,N_14924,N_12511);
and U15076 (N_15076,N_12017,N_12211);
xor U15077 (N_15077,N_14591,N_12122);
and U15078 (N_15078,N_13762,N_14473);
nor U15079 (N_15079,N_12222,N_13632);
xnor U15080 (N_15080,N_14165,N_13263);
xnor U15081 (N_15081,N_13950,N_14315);
nand U15082 (N_15082,N_14526,N_14648);
nand U15083 (N_15083,N_13940,N_13620);
xor U15084 (N_15084,N_14806,N_13423);
or U15085 (N_15085,N_12328,N_13009);
or U15086 (N_15086,N_12960,N_12342);
nor U15087 (N_15087,N_13782,N_13608);
and U15088 (N_15088,N_12718,N_12571);
xor U15089 (N_15089,N_13109,N_14021);
and U15090 (N_15090,N_14730,N_13458);
and U15091 (N_15091,N_13022,N_12860);
or U15092 (N_15092,N_13404,N_12782);
nor U15093 (N_15093,N_14511,N_14109);
nand U15094 (N_15094,N_13320,N_12312);
xnor U15095 (N_15095,N_12259,N_13071);
xor U15096 (N_15096,N_12820,N_13310);
and U15097 (N_15097,N_12131,N_14443);
nand U15098 (N_15098,N_14821,N_12916);
nand U15099 (N_15099,N_12385,N_14833);
nand U15100 (N_15100,N_12864,N_14329);
nand U15101 (N_15101,N_14138,N_13243);
xor U15102 (N_15102,N_14965,N_14969);
xor U15103 (N_15103,N_13914,N_12047);
xnor U15104 (N_15104,N_14409,N_14192);
nand U15105 (N_15105,N_14425,N_12242);
and U15106 (N_15106,N_14502,N_13469);
or U15107 (N_15107,N_12905,N_14155);
nand U15108 (N_15108,N_12272,N_12917);
xor U15109 (N_15109,N_14817,N_12430);
or U15110 (N_15110,N_13403,N_12432);
or U15111 (N_15111,N_13748,N_12347);
nand U15112 (N_15112,N_14453,N_14105);
nor U15113 (N_15113,N_12133,N_13377);
and U15114 (N_15114,N_14610,N_14866);
or U15115 (N_15115,N_12999,N_14430);
or U15116 (N_15116,N_12514,N_12610);
nand U15117 (N_15117,N_14927,N_12417);
xor U15118 (N_15118,N_13457,N_13277);
and U15119 (N_15119,N_13478,N_13475);
nor U15120 (N_15120,N_14286,N_14220);
nor U15121 (N_15121,N_13334,N_14100);
nand U15122 (N_15122,N_13241,N_12697);
or U15123 (N_15123,N_13135,N_13086);
or U15124 (N_15124,N_14579,N_12084);
nand U15125 (N_15125,N_14121,N_13681);
nand U15126 (N_15126,N_14846,N_14068);
nand U15127 (N_15127,N_13144,N_14688);
or U15128 (N_15128,N_14215,N_13380);
and U15129 (N_15129,N_13696,N_12526);
xnor U15130 (N_15130,N_13569,N_12013);
and U15131 (N_15131,N_14568,N_12323);
nand U15132 (N_15132,N_14400,N_12679);
and U15133 (N_15133,N_13284,N_13252);
or U15134 (N_15134,N_14200,N_14134);
nand U15135 (N_15135,N_12087,N_12837);
nor U15136 (N_15136,N_13755,N_14887);
nand U15137 (N_15137,N_13424,N_14532);
nor U15138 (N_15138,N_13980,N_14487);
nand U15139 (N_15139,N_12807,N_13041);
or U15140 (N_15140,N_12735,N_12070);
nor U15141 (N_15141,N_14459,N_13153);
or U15142 (N_15142,N_12689,N_13861);
xor U15143 (N_15143,N_12321,N_14991);
or U15144 (N_15144,N_12416,N_12591);
and U15145 (N_15145,N_14693,N_12340);
and U15146 (N_15146,N_13723,N_14349);
xnor U15147 (N_15147,N_12800,N_14623);
xor U15148 (N_15148,N_13878,N_13839);
or U15149 (N_15149,N_14089,N_13197);
nand U15150 (N_15150,N_12377,N_13233);
xnor U15151 (N_15151,N_14886,N_12227);
xor U15152 (N_15152,N_12298,N_14574);
and U15153 (N_15153,N_13495,N_12151);
or U15154 (N_15154,N_14615,N_12564);
or U15155 (N_15155,N_13606,N_13417);
nor U15156 (N_15156,N_12886,N_12537);
nand U15157 (N_15157,N_12111,N_12176);
or U15158 (N_15158,N_12112,N_13039);
xnor U15159 (N_15159,N_13212,N_14046);
and U15160 (N_15160,N_14986,N_13788);
nor U15161 (N_15161,N_14446,N_12360);
nor U15162 (N_15162,N_14554,N_13485);
nor U15163 (N_15163,N_13747,N_14754);
or U15164 (N_15164,N_13042,N_14348);
nor U15165 (N_15165,N_12616,N_13765);
nor U15166 (N_15166,N_13619,N_14950);
nor U15167 (N_15167,N_14582,N_12760);
or U15168 (N_15168,N_14577,N_13090);
and U15169 (N_15169,N_12806,N_12710);
nand U15170 (N_15170,N_14153,N_12634);
nor U15171 (N_15171,N_12164,N_12319);
and U15172 (N_15172,N_14282,N_14935);
nor U15173 (N_15173,N_13560,N_14792);
or U15174 (N_15174,N_13142,N_13941);
and U15175 (N_15175,N_14781,N_12894);
nand U15176 (N_15176,N_13548,N_13740);
nor U15177 (N_15177,N_14474,N_14889);
nand U15178 (N_15178,N_13500,N_12027);
and U15179 (N_15179,N_14654,N_12269);
or U15180 (N_15180,N_13821,N_13528);
or U15181 (N_15181,N_12542,N_14545);
nand U15182 (N_15182,N_14107,N_14757);
xor U15183 (N_15183,N_13828,N_14370);
xnor U15184 (N_15184,N_13733,N_13444);
or U15185 (N_15185,N_12543,N_14227);
and U15186 (N_15186,N_12440,N_12513);
and U15187 (N_15187,N_14544,N_14120);
or U15188 (N_15188,N_14137,N_13575);
and U15189 (N_15189,N_14313,N_12761);
xnor U15190 (N_15190,N_14670,N_13506);
or U15191 (N_15191,N_12334,N_13553);
or U15192 (N_15192,N_13562,N_14396);
and U15193 (N_15193,N_13164,N_14876);
nand U15194 (N_15194,N_12892,N_13306);
nor U15195 (N_15195,N_12436,N_14060);
and U15196 (N_15196,N_14696,N_14675);
xor U15197 (N_15197,N_12431,N_13667);
xor U15198 (N_15198,N_12032,N_12506);
nand U15199 (N_15199,N_13649,N_14235);
or U15200 (N_15200,N_13177,N_13996);
nor U15201 (N_15201,N_13015,N_14219);
or U15202 (N_15202,N_13393,N_12503);
nand U15203 (N_15203,N_14669,N_14339);
nor U15204 (N_15204,N_13343,N_12908);
xnor U15205 (N_15205,N_13602,N_12502);
xnor U15206 (N_15206,N_14356,N_14359);
xnor U15207 (N_15207,N_13666,N_14237);
xor U15208 (N_15208,N_13884,N_13095);
and U15209 (N_15209,N_13329,N_13780);
nand U15210 (N_15210,N_13149,N_13346);
and U15211 (N_15211,N_13892,N_13075);
or U15212 (N_15212,N_12462,N_13055);
xor U15213 (N_15213,N_14457,N_14489);
or U15214 (N_15214,N_12376,N_13106);
nand U15215 (N_15215,N_12709,N_12927);
or U15216 (N_15216,N_14382,N_14032);
nand U15217 (N_15217,N_12873,N_13502);
xor U15218 (N_15218,N_12593,N_13442);
or U15219 (N_15219,N_13509,N_13260);
nor U15220 (N_15220,N_14510,N_12563);
and U15221 (N_15221,N_13871,N_13092);
xor U15222 (N_15222,N_13439,N_14531);
or U15223 (N_15223,N_14565,N_12068);
and U15224 (N_15224,N_13167,N_12508);
nor U15225 (N_15225,N_12658,N_13318);
nand U15226 (N_15226,N_14575,N_14625);
or U15227 (N_15227,N_12378,N_12030);
and U15228 (N_15228,N_12392,N_12985);
and U15229 (N_15229,N_14206,N_13436);
nor U15230 (N_15230,N_14395,N_13063);
and U15231 (N_15231,N_14980,N_12234);
nand U15232 (N_15232,N_12364,N_13081);
xnor U15233 (N_15233,N_13406,N_13652);
xor U15234 (N_15234,N_13120,N_14930);
nand U15235 (N_15235,N_13143,N_12991);
or U15236 (N_15236,N_13546,N_13557);
nor U15237 (N_15237,N_14783,N_13927);
or U15238 (N_15238,N_14805,N_14041);
xor U15239 (N_15239,N_14205,N_13217);
nor U15240 (N_15240,N_13807,N_14125);
or U15241 (N_15241,N_13414,N_12190);
nor U15242 (N_15242,N_12758,N_13072);
xor U15243 (N_15243,N_12824,N_12725);
and U15244 (N_15244,N_13450,N_14305);
and U15245 (N_15245,N_13048,N_13640);
xnor U15246 (N_15246,N_12520,N_14904);
nand U15247 (N_15247,N_13686,N_12799);
and U15248 (N_15248,N_12691,N_14891);
nor U15249 (N_15249,N_13510,N_14588);
or U15250 (N_15250,N_12583,N_13126);
or U15251 (N_15251,N_14649,N_14976);
or U15252 (N_15252,N_14288,N_14188);
and U15253 (N_15253,N_12393,N_13408);
and U15254 (N_15254,N_13915,N_12207);
nor U15255 (N_15255,N_14132,N_12781);
nor U15256 (N_15256,N_14199,N_12236);
and U15257 (N_15257,N_12081,N_14269);
nand U15258 (N_15258,N_12872,N_13805);
xnor U15259 (N_15259,N_13245,N_12589);
nor U15260 (N_15260,N_13311,N_14031);
and U15261 (N_15261,N_12839,N_13539);
xnor U15262 (N_15262,N_14147,N_14334);
nand U15263 (N_15263,N_12884,N_14708);
xnor U15264 (N_15264,N_13309,N_12156);
or U15265 (N_15265,N_14905,N_12674);
or U15266 (N_15266,N_13216,N_13848);
nand U15267 (N_15267,N_13743,N_12522);
and U15268 (N_15268,N_14190,N_12286);
xor U15269 (N_15269,N_13294,N_13151);
or U15270 (N_15270,N_12138,N_13845);
nor U15271 (N_15271,N_12912,N_13175);
or U15272 (N_15272,N_13677,N_13405);
xnor U15273 (N_15273,N_13957,N_14452);
and U15274 (N_15274,N_13267,N_13961);
nor U15275 (N_15275,N_13460,N_13066);
and U15276 (N_15276,N_12103,N_14431);
or U15277 (N_15277,N_14075,N_13314);
and U15278 (N_15278,N_13999,N_12980);
nor U15279 (N_15279,N_13498,N_12946);
and U15280 (N_15280,N_14426,N_13021);
xnor U15281 (N_15281,N_12663,N_14566);
or U15282 (N_15282,N_12859,N_12740);
or U15283 (N_15283,N_12359,N_14860);
nor U15284 (N_15284,N_14262,N_14010);
or U15285 (N_15285,N_14222,N_13159);
xor U15286 (N_15286,N_14715,N_14994);
xnor U15287 (N_15287,N_14844,N_12467);
nand U15288 (N_15288,N_14733,N_14530);
nor U15289 (N_15289,N_13069,N_12445);
nor U15290 (N_15290,N_12938,N_12410);
and U15291 (N_15291,N_14970,N_12909);
and U15292 (N_15292,N_13028,N_14083);
or U15293 (N_15293,N_14157,N_14778);
or U15294 (N_15294,N_12626,N_14364);
or U15295 (N_15295,N_14943,N_14583);
nand U15296 (N_15296,N_14072,N_14302);
nor U15297 (N_15297,N_14735,N_14258);
or U15298 (N_15298,N_13758,N_12585);
xnor U15299 (N_15299,N_12466,N_13477);
nand U15300 (N_15300,N_12093,N_13778);
and U15301 (N_15301,N_13901,N_14865);
nand U15302 (N_15302,N_14847,N_12094);
nor U15303 (N_15303,N_14790,N_14820);
or U15304 (N_15304,N_13124,N_12994);
xor U15305 (N_15305,N_13627,N_12284);
nand U15306 (N_15306,N_12639,N_12383);
nand U15307 (N_15307,N_13532,N_12607);
nand U15308 (N_15308,N_13269,N_14477);
xor U15309 (N_15309,N_14354,N_14008);
and U15310 (N_15310,N_13262,N_13326);
xor U15311 (N_15311,N_14618,N_13354);
or U15312 (N_15312,N_13717,N_14183);
xnor U15313 (N_15313,N_13952,N_12659);
or U15314 (N_15314,N_12576,N_14595);
nand U15315 (N_15315,N_14488,N_13626);
xnor U15316 (N_15316,N_13822,N_12443);
xnor U15317 (N_15317,N_14208,N_12536);
and U15318 (N_15318,N_12743,N_12568);
or U15319 (N_15319,N_12721,N_13797);
nor U15320 (N_15320,N_12011,N_12204);
and U15321 (N_15321,N_12596,N_14917);
or U15322 (N_15322,N_13497,N_12768);
nand U15323 (N_15323,N_14056,N_14294);
and U15324 (N_15324,N_13004,N_12021);
and U15325 (N_15325,N_13989,N_13025);
or U15326 (N_15326,N_14902,N_14187);
and U15327 (N_15327,N_14540,N_14166);
nand U15328 (N_15328,N_12484,N_12106);
nand U15329 (N_15329,N_12086,N_14209);
or U15330 (N_15330,N_13349,N_14635);
nand U15331 (N_15331,N_14605,N_12015);
or U15332 (N_15332,N_14470,N_14261);
xor U15333 (N_15333,N_12813,N_14494);
xnor U15334 (N_15334,N_12586,N_13598);
nor U15335 (N_15335,N_12664,N_13720);
or U15336 (N_15336,N_12939,N_12618);
and U15337 (N_15337,N_12581,N_14389);
nor U15338 (N_15338,N_13016,N_12950);
xor U15339 (N_15339,N_14436,N_13970);
nor U15340 (N_15340,N_13315,N_12305);
and U15341 (N_15341,N_14882,N_12688);
nor U15342 (N_15342,N_12770,N_13114);
and U15343 (N_15343,N_14015,N_14217);
and U15344 (N_15344,N_14690,N_12324);
nand U15345 (N_15345,N_13646,N_13261);
nor U15346 (N_15346,N_12179,N_12716);
and U15347 (N_15347,N_13972,N_14516);
or U15348 (N_15348,N_14196,N_13559);
and U15349 (N_15349,N_12606,N_12333);
xnor U15350 (N_15350,N_14131,N_13507);
nor U15351 (N_15351,N_14275,N_13727);
xor U15352 (N_15352,N_14168,N_13370);
and U15353 (N_15353,N_13257,N_14058);
xnor U15354 (N_15354,N_14241,N_14267);
and U15355 (N_15355,N_12351,N_12895);
nor U15356 (N_15356,N_13766,N_13253);
or U15357 (N_15357,N_13467,N_13480);
and U15358 (N_15358,N_14630,N_14745);
nor U15359 (N_15359,N_13984,N_12302);
nor U15360 (N_15360,N_12066,N_13115);
or U15361 (N_15361,N_14112,N_14835);
and U15362 (N_15362,N_13964,N_13366);
xnor U15363 (N_15363,N_13869,N_12264);
or U15364 (N_15364,N_14122,N_14938);
or U15365 (N_15365,N_13292,N_13886);
or U15366 (N_15366,N_13978,N_14377);
or U15367 (N_15367,N_12413,N_14503);
nor U15368 (N_15368,N_14900,N_12239);
nor U15369 (N_15369,N_13255,N_14599);
xor U15370 (N_15370,N_12149,N_13432);
nor U15371 (N_15371,N_13355,N_13836);
nand U15372 (N_15372,N_13122,N_12088);
and U15373 (N_15373,N_12258,N_13701);
nand U15374 (N_15374,N_12386,N_13058);
nor U15375 (N_15375,N_12408,N_12923);
xnor U15376 (N_15376,N_12796,N_12136);
or U15377 (N_15377,N_13059,N_12694);
and U15378 (N_15378,N_13520,N_14760);
xnor U15379 (N_15379,N_14203,N_14660);
xor U15380 (N_15380,N_14550,N_13827);
nand U15381 (N_15381,N_13744,N_13541);
or U15382 (N_15382,N_14586,N_13169);
nor U15383 (N_15383,N_14084,N_14316);
and U15384 (N_15384,N_12350,N_13556);
xnor U15385 (N_15385,N_12095,N_12448);
nand U15386 (N_15386,N_14016,N_12137);
nand U15387 (N_15387,N_14793,N_14920);
nor U15388 (N_15388,N_12717,N_12488);
and U15389 (N_15389,N_12609,N_14508);
and U15390 (N_15390,N_14884,N_12457);
nor U15391 (N_15391,N_14268,N_13867);
nand U15392 (N_15392,N_13190,N_12661);
and U15393 (N_15393,N_13554,N_12155);
or U15394 (N_15394,N_14038,N_12826);
xor U15395 (N_15395,N_13847,N_12165);
nand U15396 (N_15396,N_13925,N_13829);
nor U15397 (N_15397,N_12671,N_13566);
nand U15398 (N_15398,N_13248,N_12836);
nand U15399 (N_15399,N_12684,N_14872);
nor U15400 (N_15400,N_12556,N_12318);
xnor U15401 (N_15401,N_12987,N_13576);
nand U15402 (N_15402,N_14677,N_14513);
nand U15403 (N_15403,N_14786,N_12026);
nand U15404 (N_15404,N_14928,N_12091);
xor U15405 (N_15405,N_12665,N_14758);
nor U15406 (N_15406,N_14971,N_13753);
nand U15407 (N_15407,N_13584,N_13816);
nand U15408 (N_15408,N_12708,N_12861);
or U15409 (N_15409,N_12240,N_12325);
or U15410 (N_15410,N_14818,N_12967);
nor U15411 (N_15411,N_13278,N_13279);
xor U15412 (N_15412,N_12161,N_12919);
xnor U15413 (N_15413,N_12797,N_12110);
or U15414 (N_15414,N_13375,N_12680);
xnor U15415 (N_15415,N_12741,N_12134);
nor U15416 (N_15416,N_13705,N_12644);
and U15417 (N_15417,N_13664,N_14749);
xor U15418 (N_15418,N_13376,N_13934);
or U15419 (N_15419,N_12592,N_12557);
nor U15420 (N_15420,N_13180,N_12267);
and U15421 (N_15421,N_13357,N_13813);
xnor U15422 (N_15422,N_14429,N_14386);
or U15423 (N_15423,N_13105,N_14771);
or U15424 (N_15424,N_12854,N_14945);
nor U15425 (N_15425,N_13775,N_14973);
or U15426 (N_15426,N_14049,N_13050);
nor U15427 (N_15427,N_13494,N_13256);
or U15428 (N_15428,N_14604,N_13258);
or U15429 (N_15429,N_14941,N_13268);
and U15430 (N_15430,N_14779,N_14561);
nor U15431 (N_15431,N_13764,N_13631);
or U15432 (N_15432,N_13770,N_13131);
nor U15433 (N_15433,N_14877,N_14691);
and U15434 (N_15434,N_14394,N_14376);
nand U15435 (N_15435,N_13415,N_14759);
nand U15436 (N_15436,N_12270,N_14674);
or U15437 (N_15437,N_12489,N_13942);
or U15438 (N_15438,N_13855,N_13789);
nor U15439 (N_15439,N_12982,N_13675);
and U15440 (N_15440,N_14054,N_13123);
nand U15441 (N_15441,N_13465,N_12446);
or U15442 (N_15442,N_13006,N_12887);
and U15443 (N_15443,N_13953,N_13907);
xor U15444 (N_15444,N_14139,N_13078);
nor U15445 (N_15445,N_14460,N_13020);
and U15446 (N_15446,N_14608,N_12000);
xor U15447 (N_15447,N_12889,N_12830);
and U15448 (N_15448,N_12268,N_12670);
or U15449 (N_15449,N_12363,N_14587);
or U15450 (N_15450,N_14556,N_14422);
or U15451 (N_15451,N_12117,N_14230);
xor U15452 (N_15452,N_14416,N_12810);
and U15453 (N_15453,N_13472,N_13854);
and U15454 (N_15454,N_12130,N_13319);
nand U15455 (N_15455,N_14874,N_12306);
or U15456 (N_15456,N_12499,N_13818);
xnor U15457 (N_15457,N_12185,N_13603);
nor U15458 (N_15458,N_13371,N_12468);
nor U15459 (N_15459,N_13335,N_14908);
nand U15460 (N_15460,N_14434,N_13484);
nor U15461 (N_15461,N_13386,N_14870);
or U15462 (N_15462,N_14590,N_13969);
nand U15463 (N_15463,N_14250,N_12888);
nor U15464 (N_15464,N_13017,N_14118);
nor U15465 (N_15465,N_12271,N_13991);
nor U15466 (N_15466,N_13285,N_14464);
xor U15467 (N_15467,N_13443,N_12235);
nor U15468 (N_15468,N_14910,N_14849);
nor U15469 (N_15469,N_14201,N_13132);
xnor U15470 (N_15470,N_14585,N_12056);
xor U15471 (N_15471,N_13630,N_14600);
xnor U15472 (N_15472,N_13754,N_14580);
and U15473 (N_15473,N_14816,N_14761);
nor U15474 (N_15474,N_14255,N_12783);
xor U15475 (N_15475,N_12738,N_14161);
nand U15476 (N_15476,N_14365,N_14310);
or U15477 (N_15477,N_13997,N_12831);
or U15478 (N_15478,N_12793,N_13635);
or U15479 (N_15479,N_14522,N_14420);
xor U15480 (N_15480,N_14993,N_12507);
and U15481 (N_15481,N_14384,N_13921);
xnor U15482 (N_15482,N_14716,N_14233);
nand U15483 (N_15483,N_12212,N_12695);
and U15484 (N_15484,N_12719,N_12395);
nand U15485 (N_15485,N_13010,N_14172);
xor U15486 (N_15486,N_13185,N_13037);
nand U15487 (N_15487,N_13840,N_12624);
nand U15488 (N_15488,N_13928,N_14471);
xor U15489 (N_15489,N_13447,N_12951);
nand U15490 (N_15490,N_12712,N_13617);
xnor U15491 (N_15491,N_13385,N_14798);
and U15492 (N_15492,N_14458,N_13283);
or U15493 (N_15493,N_14080,N_13176);
nor U15494 (N_15494,N_13529,N_13760);
nand U15495 (N_15495,N_13476,N_14271);
or U15496 (N_15496,N_14026,N_13505);
xnor U15497 (N_15497,N_12139,N_13519);
xor U15498 (N_15498,N_12678,N_13170);
or U15499 (N_15499,N_13837,N_12141);
or U15500 (N_15500,N_12675,N_14483);
xnor U15501 (N_15501,N_13591,N_13049);
and U15502 (N_15502,N_13721,N_12229);
nor U15503 (N_15503,N_12444,N_14636);
and U15504 (N_15504,N_14005,N_13711);
and U15505 (N_15505,N_13700,N_12681);
and U15506 (N_15506,N_13526,N_14799);
nor U15507 (N_15507,N_12375,N_14727);
nor U15508 (N_15508,N_14328,N_13321);
nor U15509 (N_15509,N_14180,N_14283);
or U15510 (N_15510,N_13862,N_12910);
nand U15511 (N_15511,N_13325,N_14086);
or U15512 (N_15512,N_13193,N_13838);
or U15513 (N_15513,N_14335,N_14296);
xnor U15514 (N_15514,N_13693,N_12217);
and U15515 (N_15515,N_13129,N_13276);
nor U15516 (N_15516,N_12963,N_14788);
xor U15517 (N_15517,N_13787,N_12874);
or U15518 (N_15518,N_14702,N_14955);
and U15519 (N_15519,N_14645,N_13091);
or U15520 (N_15520,N_14330,N_14601);
or U15521 (N_15521,N_13930,N_12075);
and U15522 (N_15522,N_13419,N_14528);
or U15523 (N_15523,N_14948,N_12765);
xnor U15524 (N_15524,N_13353,N_13706);
xnor U15525 (N_15525,N_12414,N_12309);
or U15526 (N_15526,N_14323,N_13536);
xor U15527 (N_15527,N_12604,N_12613);
or U15528 (N_15528,N_13750,N_14106);
xor U15529 (N_15529,N_13521,N_13084);
or U15530 (N_15530,N_14169,N_14764);
nor U15531 (N_15531,N_12730,N_13601);
or U15532 (N_15532,N_13097,N_13511);
or U15533 (N_15533,N_14150,N_14260);
nor U15534 (N_15534,N_14243,N_13819);
nor U15535 (N_15535,N_13308,N_13060);
and U15536 (N_15536,N_12252,N_14952);
or U15537 (N_15537,N_14002,N_12205);
nor U15538 (N_15538,N_12942,N_13013);
nand U15539 (N_15539,N_12085,N_13713);
xor U15540 (N_15540,N_14776,N_14345);
xor U15541 (N_15541,N_12737,N_14104);
nand U15542 (N_15542,N_12373,N_13641);
and U15543 (N_15543,N_12411,N_12686);
or U15544 (N_15544,N_12475,N_13407);
nor U15545 (N_15545,N_12713,N_14148);
or U15546 (N_15546,N_13077,N_13944);
or U15547 (N_15547,N_14415,N_14977);
nand U15548 (N_15548,N_14747,N_14856);
nor U15549 (N_15549,N_14885,N_14322);
nand U15550 (N_15550,N_14609,N_13201);
nand U15551 (N_15551,N_13218,N_14559);
and U15552 (N_15552,N_14279,N_12534);
xnor U15553 (N_15553,N_12808,N_13155);
nor U15554 (N_15554,N_12341,N_14221);
nand U15555 (N_15555,N_12390,N_13416);
nor U15556 (N_15556,N_12577,N_14292);
xor U15557 (N_15557,N_13196,N_13499);
or U15558 (N_15558,N_14461,N_12653);
and U15559 (N_15559,N_14808,N_14320);
and U15560 (N_15560,N_14369,N_12315);
xor U15561 (N_15561,N_12546,N_13345);
or U15562 (N_15562,N_13220,N_13449);
and U15563 (N_15563,N_14765,N_12162);
and U15564 (N_15564,N_14332,N_12549);
nand U15565 (N_15565,N_13012,N_12304);
nor U15566 (N_15566,N_14841,N_12656);
or U15567 (N_15567,N_12580,N_14293);
nor U15568 (N_15568,N_14410,N_13734);
nand U15569 (N_15569,N_12198,N_13286);
xor U15570 (N_15570,N_13492,N_13756);
or U15571 (N_15571,N_13655,N_14366);
xor U15572 (N_15572,N_14607,N_12477);
nand U15573 (N_15573,N_14207,N_13644);
xor U15574 (N_15574,N_14641,N_13098);
xnor U15575 (N_15575,N_14517,N_13986);
nor U15576 (N_15576,N_13868,N_12575);
xnor U15577 (N_15577,N_12224,N_14722);
nor U15578 (N_15578,N_13290,N_13007);
and U15579 (N_15579,N_14358,N_13544);
xor U15580 (N_15580,N_14428,N_13487);
or U15581 (N_15581,N_12301,N_14496);
nand U15582 (N_15582,N_12778,N_14867);
and U15583 (N_15583,N_14957,N_13203);
nor U15584 (N_15584,N_12154,N_12337);
nand U15585 (N_15585,N_13574,N_12747);
nand U15586 (N_15586,N_12330,N_14307);
nor U15587 (N_15587,N_12693,N_12600);
xnor U15588 (N_15588,N_13582,N_12256);
nand U15589 (N_15589,N_12673,N_12707);
nor U15590 (N_15590,N_14658,N_13186);
nor U15591 (N_15591,N_12244,N_14399);
or U15592 (N_15592,N_13215,N_14581);
and U15593 (N_15593,N_13577,N_13563);
and U15594 (N_15594,N_14481,N_13796);
or U15595 (N_15595,N_14562,N_14999);
nor U15596 (N_15596,N_14814,N_14449);
xnor U15597 (N_15597,N_14499,N_12171);
xnor U15598 (N_15598,N_12196,N_12623);
and U15599 (N_15599,N_13147,N_13440);
nor U15600 (N_15600,N_14181,N_13670);
xnor U15601 (N_15601,N_14809,N_12763);
nand U15602 (N_15602,N_13222,N_14062);
nand U15603 (N_15603,N_13168,N_12899);
nor U15604 (N_15604,N_14916,N_12174);
xor U15605 (N_15605,N_12636,N_14954);
and U15606 (N_15606,N_14333,N_12934);
or U15607 (N_15607,N_13749,N_14287);
nand U15608 (N_15608,N_14055,N_14519);
and U15609 (N_15609,N_12687,N_13338);
xor U15610 (N_15610,N_14167,N_14663);
nor U15611 (N_15611,N_14001,N_14883);
xnor U15612 (N_15612,N_14076,N_14110);
xor U15613 (N_15613,N_12357,N_13125);
nor U15614 (N_15614,N_14257,N_12611);
and U15615 (N_15615,N_13558,N_13817);
xnor U15616 (N_15616,N_13206,N_14944);
nor U15617 (N_15617,N_12108,N_14078);
nor U15618 (N_15618,N_13875,N_14878);
nor U15619 (N_15619,N_12755,N_12965);
xnor U15620 (N_15620,N_13157,N_12178);
nor U15621 (N_15621,N_13102,N_12460);
and U15622 (N_15622,N_13189,N_12599);
and U15623 (N_15623,N_12300,N_13876);
and U15624 (N_15624,N_12495,N_12057);
xnor U15625 (N_15625,N_12394,N_14289);
xor U15626 (N_15626,N_12749,N_13794);
nand U15627 (N_15627,N_12172,N_14525);
nand U15628 (N_15628,N_12973,N_12573);
nand U15629 (N_15629,N_12846,N_12280);
or U15630 (N_15630,N_14019,N_12441);
nor U15631 (N_15631,N_12771,N_13360);
and U15632 (N_15632,N_14381,N_13965);
xnor U15633 (N_15633,N_13266,N_13894);
nand U15634 (N_15634,N_12996,N_14476);
nor U15635 (N_15635,N_12516,N_14462);
nor U15636 (N_15636,N_12424,N_13966);
nand U15637 (N_15637,N_12045,N_13468);
nor U15638 (N_15638,N_12067,N_14113);
nor U15639 (N_15639,N_12022,N_14837);
and U15640 (N_15640,N_14152,N_12898);
and U15641 (N_15641,N_13451,N_14212);
and U15642 (N_15642,N_13896,N_12135);
xor U15643 (N_15643,N_14210,N_12628);
or U15644 (N_15644,N_14903,N_13763);
nor U15645 (N_15645,N_12296,N_14149);
nor U15646 (N_15646,N_12058,N_12866);
nand U15647 (N_15647,N_13130,N_14729);
xnor U15648 (N_15648,N_12251,N_14438);
nor U15649 (N_15649,N_12602,N_12331);
xor U15650 (N_15650,N_13399,N_12948);
xor U15651 (N_15651,N_12515,N_12819);
and U15652 (N_15652,N_13833,N_14558);
nand U15653 (N_15653,N_12109,N_13585);
nand U15654 (N_15654,N_13580,N_14154);
and U15655 (N_15655,N_12019,N_14514);
nor U15656 (N_15656,N_13172,N_12862);
nor U15657 (N_15657,N_14070,N_12089);
xnor U15658 (N_15658,N_12226,N_13184);
nor U15659 (N_15659,N_13282,N_14739);
and U15660 (N_15660,N_12907,N_12492);
and U15661 (N_15661,N_14141,N_14782);
xor U15662 (N_15662,N_14469,N_13340);
and U15663 (N_15663,N_14959,N_13213);
xnor U15664 (N_15664,N_14682,N_14933);
or U15665 (N_15665,N_12335,N_14484);
xnor U15666 (N_15666,N_13614,N_14362);
nand U15667 (N_15667,N_13958,N_12241);
nor U15668 (N_15668,N_14890,N_13305);
or U15669 (N_15669,N_13434,N_13738);
or U15670 (N_15670,N_12114,N_12995);
and U15671 (N_15671,N_13561,N_14832);
and U15672 (N_15672,N_12143,N_14651);
and U15673 (N_15673,N_14875,N_12344);
nand U15674 (N_15674,N_14114,N_13211);
and U15675 (N_15675,N_12098,N_13388);
xor U15676 (N_15676,N_13295,N_12307);
xnor U15677 (N_15677,N_12883,N_12785);
or U15678 (N_15678,N_12425,N_13668);
nor U15679 (N_15679,N_14546,N_12777);
and U15680 (N_15680,N_14418,N_13029);
or U15681 (N_15681,N_13687,N_14280);
or U15682 (N_15682,N_12701,N_12029);
and U15683 (N_15683,N_13005,N_14151);
or U15684 (N_15684,N_13100,N_13547);
and U15685 (N_15685,N_13905,N_12418);
nor U15686 (N_15686,N_13138,N_13929);
and U15687 (N_15687,N_14082,N_14017);
nor U15688 (N_15688,N_14242,N_13919);
and U15689 (N_15689,N_12964,N_12442);
and U15690 (N_15690,N_12901,N_13221);
xor U15691 (N_15691,N_12060,N_14732);
or U15692 (N_15692,N_14057,N_14069);
or U15693 (N_15693,N_14406,N_14855);
and U15694 (N_15694,N_14836,N_12423);
nand U15695 (N_15695,N_12336,N_12402);
xnor U15696 (N_15696,N_14216,N_13182);
xor U15697 (N_15697,N_14919,N_12001);
and U15698 (N_15698,N_12757,N_12002);
or U15699 (N_15699,N_12036,N_13570);
or U15700 (N_15700,N_13783,N_14085);
or U15701 (N_15701,N_13435,N_12317);
nand U15702 (N_15702,N_14050,N_13411);
and U15703 (N_15703,N_13014,N_12642);
or U15704 (N_15704,N_14807,N_12494);
nand U15705 (N_15705,N_13913,N_14584);
or U15706 (N_15706,N_14101,N_14251);
and U15707 (N_15707,N_13975,N_13359);
nor U15708 (N_15708,N_14043,N_14228);
xor U15709 (N_15709,N_12775,N_13002);
nor U15710 (N_15710,N_14762,N_13070);
xnor U15711 (N_15711,N_12595,N_14045);
nor U15712 (N_15712,N_12834,N_12338);
nand U15713 (N_15713,N_14824,N_12438);
xor U15714 (N_15714,N_14572,N_14035);
nor U15715 (N_15715,N_14796,N_14851);
xnor U15716 (N_15716,N_14124,N_14937);
or U15717 (N_15717,N_12144,N_12332);
xor U15718 (N_15718,N_14592,N_13235);
nand U15719 (N_15719,N_12779,N_12751);
nand U15720 (N_15720,N_14317,N_13757);
xnor U15721 (N_15721,N_12566,N_14661);
and U15722 (N_15722,N_13860,N_12666);
xor U15723 (N_15723,N_12024,N_12005);
or U15724 (N_15724,N_14918,N_14947);
and U15725 (N_15725,N_14379,N_14672);
or U15726 (N_15726,N_12545,N_12645);
or U15727 (N_15727,N_14570,N_12853);
nand U15728 (N_15728,N_12262,N_13515);
xnor U15729 (N_15729,N_12474,N_14656);
and U15730 (N_15730,N_14236,N_13381);
xnor U15731 (N_15731,N_12533,N_14352);
or U15732 (N_15732,N_13690,N_12535);
and U15733 (N_15733,N_12195,N_13654);
and U15734 (N_15734,N_14065,N_13242);
and U15735 (N_15735,N_13533,N_12698);
xnor U15736 (N_15736,N_12852,N_12287);
and U15737 (N_15737,N_13792,N_12230);
nand U15738 (N_15738,N_14066,N_14119);
xor U15739 (N_15739,N_13232,N_12754);
nor U15740 (N_15740,N_13708,N_14555);
and U15741 (N_15741,N_12789,N_13967);
nor U15742 (N_15742,N_13810,N_12210);
nand U15743 (N_15743,N_14295,N_14911);
or U15744 (N_15744,N_12218,N_14687);
and U15745 (N_15745,N_14939,N_13581);
xor U15746 (N_15746,N_12092,N_13104);
nor U15747 (N_15747,N_14052,N_12496);
or U15748 (N_15748,N_14006,N_14873);
nor U15749 (N_15749,N_14925,N_12434);
or U15750 (N_15750,N_13685,N_13730);
or U15751 (N_15751,N_14324,N_12216);
nor U15752 (N_15752,N_14003,N_14706);
nand U15753 (N_15753,N_13682,N_14432);
nand U15754 (N_15754,N_12608,N_12935);
nor U15755 (N_15755,N_12491,N_13985);
xor U15756 (N_15756,N_14639,N_13244);
xor U15757 (N_15757,N_12524,N_14553);
nor U15758 (N_15758,N_14281,N_13378);
nor U15759 (N_15759,N_12231,N_13525);
and U15760 (N_15760,N_13906,N_13935);
xnor U15761 (N_15761,N_13113,N_14845);
nand U15762 (N_15762,N_14447,N_12667);
xnor U15763 (N_15763,N_12290,N_12101);
and U15764 (N_15764,N_12622,N_12147);
and U15765 (N_15765,N_14603,N_13462);
nor U15766 (N_15766,N_13236,N_12750);
xor U15767 (N_15767,N_13704,N_14263);
nand U15768 (N_15768,N_12248,N_13616);
or U15769 (N_15769,N_14229,N_14022);
xor U15770 (N_15770,N_14533,N_12016);
and U15771 (N_15771,N_14197,N_13858);
nor U15772 (N_15772,N_12560,N_13924);
nand U15773 (N_15773,N_12510,N_12992);
and U15774 (N_15774,N_14158,N_12023);
nand U15775 (N_15775,N_13527,N_14129);
nor U15776 (N_15776,N_14951,N_13830);
and U15777 (N_15777,N_12794,N_14393);
xnor U15778 (N_15778,N_12952,N_14748);
or U15779 (N_15779,N_12255,N_14811);
and U15780 (N_15780,N_14171,N_12289);
xor U15781 (N_15781,N_13148,N_12043);
and U15782 (N_15782,N_12827,N_13074);
nor U15783 (N_15783,N_12465,N_14198);
xor U15784 (N_15784,N_13859,N_12920);
xor U15785 (N_15785,N_14627,N_13207);
xnor U15786 (N_15786,N_12294,N_12943);
nand U15787 (N_15787,N_13162,N_12700);
or U15788 (N_15788,N_13651,N_12311);
and U15789 (N_15789,N_13337,N_14697);
and U15790 (N_15790,N_14785,N_14685);
or U15791 (N_15791,N_12579,N_14071);
and U15792 (N_15792,N_12815,N_14300);
and U15793 (N_15793,N_14276,N_13983);
xor U15794 (N_15794,N_14854,N_12562);
and U15795 (N_15795,N_12970,N_12464);
nand U15796 (N_15796,N_14465,N_14567);
nand U15797 (N_15797,N_12798,N_13313);
nor U15798 (N_15798,N_12527,N_14160);
xor U15799 (N_15799,N_13910,N_12523);
and U15800 (N_15800,N_13951,N_13832);
xor U15801 (N_15801,N_12984,N_13293);
xor U15802 (N_15802,N_14705,N_14115);
nor U15803 (N_15803,N_14304,N_12362);
xor U15804 (N_15804,N_14979,N_14098);
or U15805 (N_15805,N_14763,N_13219);
nor U15806 (N_15806,N_13150,N_12989);
nor U15807 (N_15807,N_13181,N_13085);
or U15808 (N_15808,N_12867,N_12010);
xnor U15809 (N_15809,N_14812,N_13112);
nor U15810 (N_15810,N_14175,N_13596);
nor U15811 (N_15811,N_14463,N_14711);
xor U15812 (N_15812,N_12079,N_13192);
and U15813 (N_15813,N_13251,N_14321);
nand U15814 (N_15814,N_13427,N_14337);
and U15815 (N_15815,N_14848,N_14963);
xor U15816 (N_15816,N_12865,N_14405);
xnor U15817 (N_15817,N_13564,N_12182);
xor U15818 (N_15818,N_13956,N_13410);
or U15819 (N_15819,N_13288,N_12276);
or U15820 (N_15820,N_12742,N_12463);
nor U15821 (N_15821,N_13684,N_14224);
nor U15822 (N_15822,N_13920,N_12397);
and U15823 (N_15823,N_14036,N_12339);
or U15824 (N_15824,N_14427,N_12979);
nor U15825 (N_15825,N_14680,N_14946);
nor U15826 (N_15826,N_14325,N_13348);
or U15827 (N_15827,N_13809,N_12261);
xnor U15828 (N_15828,N_12052,N_13032);
and U15829 (N_15829,N_12435,N_12062);
xnor U15830 (N_15830,N_13772,N_12582);
nand U15831 (N_15831,N_13594,N_14926);
and U15832 (N_15832,N_12682,N_14456);
xnor U15833 (N_15833,N_14914,N_12643);
nand U15834 (N_15834,N_12219,N_14331);
nor U15835 (N_15835,N_13397,N_14202);
and U15836 (N_15836,N_12870,N_12090);
nand U15837 (N_15837,N_12672,N_13735);
xor U15838 (N_15838,N_13146,N_14810);
xnor U15839 (N_15839,N_12221,N_14634);
nor U15840 (N_15840,N_13514,N_14244);
or U15841 (N_15841,N_14968,N_14831);
or U15842 (N_15842,N_13082,N_13490);
nand U15843 (N_15843,N_13689,N_14701);
or U15844 (N_15844,N_12329,N_14737);
or U15845 (N_15845,N_13488,N_13745);
and U15846 (N_15846,N_14380,N_12292);
xnor U15847 (N_15847,N_12931,N_12791);
xnor U15848 (N_15848,N_12553,N_13802);
and U15849 (N_15849,N_14922,N_12063);
nand U15850 (N_15850,N_12649,N_12454);
xor U15851 (N_15851,N_13080,N_12152);
xor U15852 (N_15852,N_13065,N_13550);
nand U15853 (N_15853,N_14720,N_14543);
or U15854 (N_15854,N_13779,N_12404);
and U15855 (N_15855,N_14681,N_13531);
xnor U15856 (N_15856,N_14512,N_14238);
and U15857 (N_15857,N_14259,N_13904);
and U15858 (N_15858,N_12199,N_12400);
nand U15859 (N_15859,N_13629,N_14504);
or U15860 (N_15860,N_13815,N_14989);
nor U15861 (N_15861,N_14226,N_12125);
or U15862 (N_15862,N_12519,N_14774);
and U15863 (N_15863,N_14686,N_13466);
nor U15864 (N_15864,N_14126,N_13463);
xnor U15865 (N_15865,N_14074,N_13624);
nor U15866 (N_15866,N_14520,N_12175);
nor U15867 (N_15867,N_13296,N_14423);
xnor U15868 (N_15868,N_12025,N_13790);
and U15869 (N_15869,N_14185,N_13607);
nand U15870 (N_15870,N_12816,N_14291);
xnor U15871 (N_15871,N_13633,N_12406);
nor U15872 (N_15872,N_12677,N_13163);
nor U15873 (N_15873,N_13280,N_14319);
or U15874 (N_15874,N_14913,N_12521);
nor U15875 (N_15875,N_12483,N_13872);
xnor U15876 (N_15876,N_12817,N_13773);
xnor U15877 (N_15877,N_13834,N_14374);
and U15878 (N_15878,N_13491,N_13173);
or U15879 (N_15879,N_13718,N_13053);
or U15880 (N_15880,N_13895,N_13881);
or U15881 (N_15881,N_14547,N_13119);
nor U15882 (N_15882,N_13604,N_13271);
and U15883 (N_15883,N_14412,N_13699);
nand U15884 (N_15884,N_14838,N_14684);
nor U15885 (N_15885,N_14692,N_13116);
and U15886 (N_15886,N_12915,N_14033);
nor U15887 (N_15887,N_14524,N_13725);
nand U15888 (N_15888,N_12558,N_14578);
or U15889 (N_15889,N_12843,N_13538);
or U15890 (N_15890,N_13136,N_13831);
and U15891 (N_15891,N_14439,N_14521);
or U15892 (N_15892,N_14211,N_12640);
nand U15893 (N_15893,N_12073,N_12696);
nand U15894 (N_15894,N_13356,N_13363);
or U15895 (N_15895,N_14509,N_14385);
nand U15896 (N_15896,N_12099,N_14030);
nand U15897 (N_15897,N_13425,N_13703);
and U15898 (N_15898,N_12384,N_12928);
nor U15899 (N_15899,N_14048,N_14498);
xnor U15900 (N_15900,N_12006,N_12206);
nor U15901 (N_15901,N_13767,N_14096);
or U15902 (N_15902,N_13275,N_12214);
nand U15903 (N_15903,N_14879,N_12470);
or U15904 (N_15904,N_14194,N_13224);
xnor U15905 (N_15905,N_12620,N_12215);
and U15906 (N_15906,N_12993,N_13281);
nand U15907 (N_15907,N_14040,N_12715);
nor U15908 (N_15908,N_14839,N_12879);
or U15909 (N_15909,N_14239,N_12662);
nand U15910 (N_15910,N_12451,N_13540);
or U15911 (N_15911,N_14589,N_14273);
and U15912 (N_15912,N_13995,N_13336);
xor U15913 (N_15913,N_14731,N_12396);
nor U15914 (N_15914,N_13659,N_13240);
or U15915 (N_15915,N_13199,N_14000);
xnor U15916 (N_15916,N_14898,N_12050);
nor U15917 (N_15917,N_14703,N_13237);
and U15918 (N_15918,N_14746,N_14466);
or U15919 (N_15919,N_14407,N_14892);
nor U15920 (N_15920,N_14772,N_13452);
xnor U15921 (N_15921,N_12209,N_12961);
and U15922 (N_15922,N_13043,N_13595);
or U15923 (N_15923,N_13108,N_13339);
or U15924 (N_15924,N_14303,N_14357);
nand U15925 (N_15925,N_14051,N_13567);
nor U15926 (N_15926,N_12253,N_13545);
nand U15927 (N_15927,N_12787,N_13900);
or U15928 (N_15928,N_13549,N_12278);
and U15929 (N_15929,N_14864,N_14961);
nor U15930 (N_15930,N_13799,N_14435);
or U15931 (N_15931,N_14403,N_14893);
and U15932 (N_15932,N_12541,N_12655);
nand U15933 (N_15933,N_13128,N_13998);
or U15934 (N_15934,N_14563,N_13518);
or U15935 (N_15935,N_12774,N_13300);
and U15936 (N_15936,N_13800,N_12732);
nor U15937 (N_15937,N_12249,N_12159);
nand U15938 (N_15938,N_12578,N_14800);
xor U15939 (N_15939,N_13611,N_14090);
xor U15940 (N_15940,N_12812,N_12728);
or U15941 (N_15941,N_12932,N_13530);
xnor U15942 (N_15942,N_12121,N_14742);
xor U15943 (N_15943,N_13134,N_14146);
and U15944 (N_15944,N_13739,N_14355);
and U15945 (N_15945,N_12998,N_12254);
and U15946 (N_15946,N_13099,N_12726);
or U15947 (N_15947,N_12974,N_14784);
nand U15948 (N_15948,N_14341,N_13101);
nor U15949 (N_15949,N_12570,N_13483);
nand U15950 (N_15950,N_12949,N_12447);
nand U15951 (N_15951,N_14662,N_12180);
nor U15952 (N_15952,N_13990,N_13974);
or U15953 (N_15953,N_13918,N_12356);
or U15954 (N_15954,N_12203,N_13396);
nor U15955 (N_15955,N_13165,N_12766);
nor U15956 (N_15956,N_12552,N_12648);
nor U15957 (N_15957,N_14564,N_12293);
or U15958 (N_15958,N_13400,N_12983);
nor U15959 (N_15959,N_12792,N_12518);
nand U15960 (N_15960,N_13759,N_13716);
xor U15961 (N_15961,N_13394,N_14633);
or U15962 (N_15962,N_12353,N_14666);
xor U15963 (N_15963,N_14441,N_14551);
nand U15964 (N_15964,N_13590,N_12724);
nor U15965 (N_15965,N_13883,N_12193);
and U15966 (N_15966,N_12345,N_14482);
nand U15967 (N_15967,N_12840,N_13674);
nor U15968 (N_15968,N_13019,N_13482);
and U15969 (N_15969,N_14830,N_13145);
nand U15970 (N_15970,N_12569,N_12129);
and U15971 (N_15971,N_14725,N_14248);
xor U15972 (N_15972,N_13384,N_14655);
or U15973 (N_15973,N_14894,N_14053);
nand U15974 (N_15974,N_14679,N_14527);
xor U15975 (N_15975,N_12547,N_14475);
nor U15976 (N_15976,N_13054,N_12225);
nor U15977 (N_15977,N_13628,N_13589);
or U15978 (N_15978,N_14290,N_14995);
xor U15979 (N_15979,N_12421,N_13350);
nand U15980 (N_15980,N_13426,N_13272);
and U15981 (N_15981,N_14097,N_13852);
or U15982 (N_15982,N_14990,N_13534);
xor U15983 (N_15983,N_12428,N_14361);
nand U15984 (N_15984,N_13094,N_13052);
xor U15985 (N_15985,N_14536,N_12646);
or U15986 (N_15986,N_12072,N_14698);
xnor U15987 (N_15987,N_13489,N_12472);
nor U15988 (N_15988,N_12723,N_13902);
nand U15989 (N_15989,N_12955,N_13835);
or U15990 (N_15990,N_13367,N_13746);
nand U15991 (N_15991,N_13959,N_12896);
and U15992 (N_15992,N_14723,N_12880);
xnor U15993 (N_15993,N_13141,N_12285);
nand U15994 (N_15994,N_12981,N_13362);
nor U15995 (N_15995,N_13517,N_13769);
or U15996 (N_15996,N_13903,N_14773);
xnor U15997 (N_15997,N_12266,N_12399);
xnor U15998 (N_15998,N_12118,N_12126);
nand U15999 (N_15999,N_13341,N_12603);
nor U16000 (N_16000,N_14170,N_13968);
xnor U16001 (N_16001,N_13737,N_13874);
or U16002 (N_16002,N_13289,N_13422);
and U16003 (N_16003,N_13209,N_14858);
nor U16004 (N_16004,N_14245,N_12361);
or U16005 (N_16005,N_13712,N_13784);
and U16006 (N_16006,N_12061,N_14454);
and U16007 (N_16007,N_13493,N_14145);
and U16008 (N_16008,N_12780,N_14710);
and U16009 (N_16009,N_13587,N_14472);
and U16010 (N_16010,N_14326,N_12871);
xnor U16011 (N_16011,N_13736,N_14014);
or U16012 (N_16012,N_12764,N_12482);
or U16013 (N_16013,N_13793,N_13259);
nand U16014 (N_16014,N_13210,N_13312);
or U16015 (N_16015,N_13808,N_14813);
nand U16016 (N_16016,N_13683,N_12288);
xnor U16017 (N_16017,N_12274,N_12105);
or U16018 (N_16018,N_14039,N_13035);
xnor U16019 (N_16019,N_13096,N_14897);
and U16020 (N_16020,N_13945,N_13270);
and U16021 (N_16021,N_14391,N_12921);
nor U16022 (N_16022,N_13140,N_12107);
and U16023 (N_16023,N_14953,N_12263);
nor U16024 (N_16024,N_12183,N_13161);
nand U16025 (N_16025,N_12914,N_12784);
or U16026 (N_16026,N_14539,N_14614);
or U16027 (N_16027,N_14011,N_12297);
nand U16028 (N_16028,N_14936,N_12220);
xnor U16029 (N_16029,N_14988,N_14253);
nand U16030 (N_16030,N_12734,N_13121);
nor U16031 (N_16031,N_14707,N_14500);
xnor U16032 (N_16032,N_13785,N_13932);
or U16033 (N_16033,N_14992,N_14612);
xor U16034 (N_16034,N_12703,N_12976);
xor U16035 (N_16035,N_13771,N_14535);
nand U16036 (N_16036,N_14622,N_12473);
nor U16037 (N_16037,N_14770,N_12832);
xnor U16038 (N_16038,N_13948,N_14346);
and U16039 (N_16039,N_13154,N_12189);
xnor U16040 (N_16040,N_13067,N_13888);
nor U16041 (N_16041,N_13653,N_14801);
nand U16042 (N_16042,N_14350,N_13501);
and U16043 (N_16043,N_14606,N_14643);
nor U16044 (N_16044,N_12371,N_12657);
and U16045 (N_16045,N_14768,N_14284);
or U16046 (N_16046,N_13420,N_14347);
and U16047 (N_16047,N_14724,N_13943);
or U16048 (N_16048,N_12401,N_14034);
xnor U16049 (N_16049,N_12055,N_12132);
or U16050 (N_16050,N_14007,N_12720);
nor U16051 (N_16051,N_12926,N_12654);
and U16052 (N_16052,N_12668,N_14353);
nand U16053 (N_16053,N_12039,N_12903);
and U16054 (N_16054,N_14712,N_13413);
nand U16055 (N_16055,N_14534,N_13873);
and U16056 (N_16056,N_14736,N_13722);
and U16057 (N_16057,N_12858,N_14179);
or U16058 (N_16058,N_12615,N_13850);
xor U16059 (N_16059,N_13391,N_12612);
and U16060 (N_16060,N_12181,N_12044);
nand U16061 (N_16061,N_14029,N_13046);
and U16062 (N_16062,N_13642,N_12746);
nand U16063 (N_16063,N_14367,N_14223);
nor U16064 (N_16064,N_14628,N_14853);
and U16065 (N_16065,N_13471,N_14542);
nor U16066 (N_16066,N_12391,N_14193);
xor U16067 (N_16067,N_14299,N_12539);
nand U16068 (N_16068,N_13395,N_12968);
nor U16069 (N_16069,N_12773,N_14372);
nand U16070 (N_16070,N_13038,N_13373);
and U16071 (N_16071,N_14099,N_13342);
xnor U16072 (N_16072,N_12403,N_13806);
nor U16073 (N_16073,N_13433,N_14013);
nand U16074 (N_16074,N_14640,N_14344);
and U16075 (N_16075,N_12588,N_14974);
xor U16076 (N_16076,N_12877,N_14834);
and U16077 (N_16077,N_12605,N_14493);
xnor U16078 (N_16078,N_13298,N_12382);
and U16079 (N_16079,N_14895,N_14028);
nor U16080 (N_16080,N_14414,N_14189);
nand U16081 (N_16081,N_14673,N_14177);
nor U16082 (N_16082,N_14794,N_14108);
nand U16083 (N_16083,N_12997,N_12811);
and U16084 (N_16084,N_14306,N_13897);
nand U16085 (N_16085,N_12890,N_12485);
nand U16086 (N_16086,N_13893,N_13613);
xor U16087 (N_16087,N_12786,N_13931);
or U16088 (N_16088,N_14650,N_14750);
nor U16089 (N_16089,N_14133,N_12619);
xor U16090 (N_16090,N_13264,N_12453);
nor U16091 (N_16091,N_13988,N_12478);
nor U16092 (N_16092,N_12500,N_13473);
nand U16093 (N_16093,N_12127,N_13709);
nor U16094 (N_16094,N_14195,N_12531);
and U16095 (N_16095,N_14507,N_14896);
and U16096 (N_16096,N_13470,N_13001);
nand U16097 (N_16097,N_12805,N_12486);
or U16098 (N_16098,N_12838,N_14548);
nand U16099 (N_16099,N_12802,N_14751);
or U16100 (N_16100,N_14665,N_12814);
nand U16101 (N_16101,N_12882,N_14383);
and U16102 (N_16102,N_12594,N_14863);
nand U16103 (N_16103,N_14653,N_13522);
xnor U16104 (N_16104,N_12823,N_13369);
nor U16105 (N_16105,N_12481,N_12469);
xor U16106 (N_16106,N_12082,N_12148);
nand U16107 (N_16107,N_12201,N_14621);
and U16108 (N_16108,N_12512,N_14127);
nand U16109 (N_16109,N_12829,N_14485);
xor U16110 (N_16110,N_12601,N_12009);
or U16111 (N_16111,N_12407,N_13307);
nor U16112 (N_16112,N_14204,N_12049);
or U16113 (N_16113,N_13226,N_14718);
xor U16114 (N_16114,N_12146,N_12971);
xor U16115 (N_16115,N_13625,N_13368);
or U16116 (N_16116,N_13657,N_12913);
and U16117 (N_16117,N_13327,N_14042);
nor U16118 (N_16118,N_12041,N_13008);
xor U16119 (N_16119,N_13194,N_12257);
or U16120 (N_16120,N_12422,N_12878);
nand U16121 (N_16121,N_13571,N_12567);
nand U16122 (N_16122,N_14949,N_13811);
or U16123 (N_16123,N_12753,N_14646);
nand U16124 (N_16124,N_13938,N_13857);
nor U16125 (N_16125,N_13971,N_12739);
nand U16126 (N_16126,N_13474,N_13592);
or U16127 (N_16127,N_14312,N_14560);
and U16128 (N_16128,N_12933,N_14827);
or U16129 (N_16129,N_14629,N_12381);
xor U16130 (N_16130,N_14888,N_14802);
xnor U16131 (N_16131,N_14741,N_12449);
or U16132 (N_16132,N_12752,N_13926);
xor U16133 (N_16133,N_13412,N_14402);
xor U16134 (N_16134,N_12299,N_12322);
or U16135 (N_16135,N_13127,N_14631);
or U16136 (N_16136,N_13249,N_12498);
and U16137 (N_16137,N_14444,N_14934);
nand U16138 (N_16138,N_13698,N_13139);
xnor U16139 (N_16139,N_14249,N_14308);
or U16140 (N_16140,N_12857,N_14419);
xor U16141 (N_16141,N_14254,N_13572);
and U16142 (N_16142,N_13599,N_12365);
and U16143 (N_16143,N_13234,N_12420);
nand U16144 (N_16144,N_14940,N_13239);
nand U16145 (N_16145,N_12059,N_13302);
nor U16146 (N_16146,N_12804,N_13331);
and U16147 (N_16147,N_12529,N_12736);
nor U16148 (N_16148,N_14652,N_14387);
nand U16149 (N_16149,N_12426,N_14044);
nor U16150 (N_16150,N_12772,N_14752);
nor U16151 (N_16151,N_13156,N_14272);
and U16152 (N_16152,N_14012,N_12714);
nand U16153 (N_16153,N_14103,N_14421);
nand U16154 (N_16154,N_12007,N_14506);
nor U16155 (N_16155,N_12020,N_13937);
nor U16156 (N_16156,N_14967,N_12343);
xnor U16157 (N_16157,N_12745,N_12958);
xor U16158 (N_16158,N_14529,N_14388);
or U16159 (N_16159,N_12733,N_13398);
or U16160 (N_16160,N_14159,N_14162);
or U16161 (N_16161,N_12809,N_13776);
or U16162 (N_16162,N_14912,N_14117);
nor U16163 (N_16163,N_12096,N_14868);
and U16164 (N_16164,N_14978,N_14373);
nand U16165 (N_16165,N_12501,N_12405);
or U16166 (N_16166,N_14619,N_14907);
nand U16167 (N_16167,N_12821,N_13324);
nor U16168 (N_16168,N_13605,N_13648);
or U16169 (N_16169,N_14130,N_14632);
xor U16170 (N_16170,N_12160,N_12731);
nor U16171 (N_16171,N_12505,N_12692);
nand U16172 (N_16172,N_12683,N_14455);
or U16173 (N_16173,N_13660,N_12660);
nor U16174 (N_16174,N_13023,N_14932);
nand U16175 (N_16175,N_12629,N_14186);
nor U16176 (N_16176,N_12621,N_14440);
nand U16177 (N_16177,N_13729,N_14997);
xnor U16178 (N_16178,N_12232,N_12415);
or U16179 (N_16179,N_12631,N_12283);
xnor U16180 (N_16180,N_14136,N_14297);
or U16181 (N_16181,N_14232,N_12250);
nand U16182 (N_16182,N_14804,N_12904);
nor U16183 (N_16183,N_14823,N_12699);
and U16184 (N_16184,N_12833,N_12497);
nor U16185 (N_16185,N_13187,N_14901);
and U16186 (N_16186,N_12140,N_14027);
xor U16187 (N_16187,N_14644,N_13656);
and U16188 (N_16188,N_13588,N_12555);
and U16189 (N_16189,N_13825,N_14942);
xor U16190 (N_16190,N_12048,N_12123);
or U16191 (N_16191,N_12550,N_13933);
xnor U16192 (N_16192,N_13724,N_14909);
or U16193 (N_16193,N_14695,N_12115);
nor U16194 (N_16194,N_14518,N_13160);
and U16195 (N_16195,N_13728,N_14714);
nand U16196 (N_16196,N_12031,N_14067);
nand U16197 (N_16197,N_12937,N_13565);
nor U16198 (N_16198,N_13768,N_12885);
nor U16199 (N_16199,N_13430,N_12169);
or U16200 (N_16200,N_14378,N_14557);
and U16201 (N_16201,N_14537,N_14734);
nor U16202 (N_16202,N_13786,N_13714);
nor U16203 (N_16203,N_13803,N_14915);
xnor U16204 (N_16204,N_12930,N_12369);
nand U16205 (N_16205,N_14218,N_14491);
xor U16206 (N_16206,N_14116,N_13568);
and U16207 (N_16207,N_12849,N_13841);
xnor U16208 (N_16208,N_13061,N_14797);
nor U16209 (N_16209,N_12855,N_12379);
and U16210 (N_16210,N_14642,N_13993);
and U16211 (N_16211,N_13936,N_13223);
nor U16212 (N_16212,N_14740,N_12598);
xor U16213 (N_16213,N_14998,N_14073);
and U16214 (N_16214,N_13647,N_13643);
and U16215 (N_16215,N_12150,N_12953);
xor U16216 (N_16216,N_12076,N_13018);
and U16217 (N_16217,N_12767,N_14984);
nand U16218 (N_16218,N_12071,N_12213);
xor U16219 (N_16219,N_13863,N_12188);
xor U16220 (N_16220,N_14327,N_13679);
or U16221 (N_16221,N_13795,N_14213);
xnor U16222 (N_16222,N_14505,N_14480);
and U16223 (N_16223,N_12040,N_12978);
nand U16224 (N_16224,N_13719,N_13650);
nor U16225 (N_16225,N_13178,N_12003);
xor U16226 (N_16226,N_13171,N_13911);
or U16227 (N_16227,N_12551,N_12632);
or U16228 (N_16228,N_12388,N_13118);
nor U16229 (N_16229,N_14880,N_12200);
or U16230 (N_16230,N_13673,N_13707);
nand U16231 (N_16231,N_14191,N_12528);
xor U16232 (N_16232,N_14842,N_12303);
or U16233 (N_16233,N_12647,N_13246);
and U16234 (N_16234,N_14301,N_12370);
nand U16235 (N_16235,N_12828,N_12493);
nor U16236 (N_16236,N_13379,N_14024);
nor U16237 (N_16237,N_13665,N_14975);
nand U16238 (N_16238,N_14495,N_13372);
xor U16239 (N_16239,N_13000,N_14617);
nand U16240 (N_16240,N_12450,N_14576);
nor U16241 (N_16241,N_13676,N_13344);
and U16242 (N_16242,N_12387,N_12316);
or U16243 (N_16243,N_14664,N_14598);
nor U16244 (N_16244,N_12034,N_14613);
nor U16245 (N_16245,N_14803,N_14981);
and U16246 (N_16246,N_13250,N_12158);
nor U16247 (N_16247,N_13361,N_12940);
and U16248 (N_16248,N_13179,N_13428);
and U16249 (N_16249,N_13438,N_13323);
nor U16250 (N_16250,N_12233,N_13382);
or U16251 (N_16251,N_14964,N_12157);
nand U16252 (N_16252,N_14174,N_13158);
nand U16253 (N_16253,N_12776,N_14448);
and U16254 (N_16254,N_13917,N_14497);
xnor U16255 (N_16255,N_12988,N_12544);
nor U16256 (N_16256,N_13229,N_14091);
nor U16257 (N_16257,N_12969,N_13231);
or U16258 (N_16258,N_13695,N_13437);
and U16259 (N_16259,N_14637,N_12947);
xor U16260 (N_16260,N_14899,N_14789);
or U16261 (N_16261,N_14037,N_12223);
or U16262 (N_16262,N_13333,N_12902);
nand U16263 (N_16263,N_12897,N_14087);
and U16264 (N_16264,N_13034,N_12936);
xnor U16265 (N_16265,N_14164,N_12966);
xnor U16266 (N_16266,N_14694,N_14719);
xnor U16267 (N_16267,N_13761,N_14143);
or U16268 (N_16268,N_13036,N_12479);
nor U16269 (N_16269,N_13955,N_13027);
or U16270 (N_16270,N_13741,N_13669);
nand U16271 (N_16271,N_13516,N_12004);
and U16272 (N_16272,N_13600,N_13688);
and U16273 (N_16273,N_13068,N_13672);
nor U16274 (N_16274,N_13076,N_12651);
or U16275 (N_16275,N_14815,N_12279);
nand U16276 (N_16276,N_13697,N_12490);
nor U16277 (N_16277,N_12456,N_12119);
nand U16278 (N_16278,N_12168,N_13979);
xor U16279 (N_16279,N_12247,N_14573);
nor U16280 (N_16280,N_13062,N_14753);
and U16281 (N_16281,N_13949,N_14128);
nand U16282 (N_16282,N_12142,N_12722);
nor U16283 (N_16283,N_14442,N_13742);
xnor U16284 (N_16284,N_13612,N_12398);
xnor U16285 (N_16285,N_14411,N_12929);
nor U16286 (N_16286,N_12676,N_12650);
xor U16287 (N_16287,N_14404,N_12532);
or U16288 (N_16288,N_13137,N_13671);
or U16289 (N_16289,N_13992,N_13374);
and U16290 (N_16290,N_12975,N_14956);
or U16291 (N_16291,N_12850,N_14828);
or U16292 (N_16292,N_12959,N_13057);
or U16293 (N_16293,N_14676,N_12008);
and U16294 (N_16294,N_13087,N_14417);
and U16295 (N_16295,N_13543,N_14596);
nand U16296 (N_16296,N_14020,N_13455);
nand U16297 (N_16297,N_14569,N_12554);
nand U16298 (N_16298,N_13198,N_12835);
or U16299 (N_16299,N_13024,N_14231);
nor U16300 (N_16300,N_14163,N_12652);
or U16301 (N_16301,N_12881,N_12803);
and U16302 (N_16302,N_14501,N_14064);
and U16303 (N_16303,N_12228,N_13645);
nor U16304 (N_16304,N_12727,N_12326);
nand U16305 (N_16305,N_13454,N_13751);
xnor U16306 (N_16306,N_12762,N_14843);
xor U16307 (N_16307,N_13826,N_13409);
xor U16308 (N_16308,N_12238,N_14647);
or U16309 (N_16309,N_13962,N_12177);
nor U16310 (N_16310,N_13030,N_13044);
or U16311 (N_16311,N_12194,N_12173);
or U16312 (N_16312,N_12587,N_13110);
and U16313 (N_16313,N_13512,N_13230);
nor U16314 (N_16314,N_13459,N_14144);
nand U16315 (N_16315,N_12517,N_14363);
nor U16316 (N_16316,N_12458,N_14375);
nor U16317 (N_16317,N_13877,N_14478);
and U16318 (N_16318,N_13555,N_13047);
or U16319 (N_16319,N_12635,N_12868);
and U16320 (N_16320,N_13638,N_14252);
xnor U16321 (N_16321,N_12035,N_12145);
or U16322 (N_16322,N_14620,N_14490);
xor U16323 (N_16323,N_13981,N_12627);
or U16324 (N_16324,N_14351,N_14467);
xnor U16325 (N_16325,N_12208,N_12876);
and U16326 (N_16326,N_12197,N_14102);
xnor U16327 (N_16327,N_13973,N_14593);
nor U16328 (N_16328,N_13103,N_14777);
and U16329 (N_16329,N_14958,N_13774);
or U16330 (N_16330,N_13214,N_13661);
or U16331 (N_16331,N_13301,N_13446);
nor U16332 (N_16332,N_13732,N_14140);
xnor U16333 (N_16333,N_13923,N_13621);
and U16334 (N_16334,N_12124,N_13637);
xor U16335 (N_16335,N_14795,N_14826);
and U16336 (N_16336,N_13597,N_13390);
and U16337 (N_16337,N_14368,N_14852);
xor U16338 (N_16338,N_13916,N_13133);
and U16339 (N_16339,N_13274,N_14921);
or U16340 (N_16340,N_14657,N_14111);
nand U16341 (N_16341,N_12844,N_12053);
nor U16342 (N_16342,N_13523,N_14277);
and U16343 (N_16343,N_13982,N_13200);
xor U16344 (N_16344,N_14611,N_13351);
and U16345 (N_16345,N_13987,N_12366);
nand U16346 (N_16346,N_13191,N_12455);
nor U16347 (N_16347,N_12572,N_14775);
and U16348 (N_16348,N_12078,N_14857);
nand U16349 (N_16349,N_14059,N_14602);
xor U16350 (N_16350,N_14298,N_13402);
and U16351 (N_16351,N_13079,N_12074);
xor U16352 (N_16352,N_14756,N_13088);
and U16353 (N_16353,N_14960,N_14923);
nand U16354 (N_16354,N_13890,N_12295);
nand U16355 (N_16355,N_12590,N_14424);
or U16356 (N_16356,N_13045,N_12313);
or U16357 (N_16357,N_13011,N_13195);
and U16358 (N_16358,N_13448,N_13031);
nand U16359 (N_16359,N_14018,N_13166);
xnor U16360 (N_16360,N_14023,N_14343);
xor U16361 (N_16361,N_13227,N_12100);
and U16362 (N_16362,N_12922,N_13291);
and U16363 (N_16363,N_14479,N_12790);
or U16364 (N_16364,N_13960,N_12972);
xnor U16365 (N_16365,N_14081,N_14270);
nand U16366 (N_16366,N_13265,N_12538);
nand U16367 (N_16367,N_13429,N_14445);
nor U16368 (N_16368,N_13479,N_14906);
and U16369 (N_16369,N_14728,N_14173);
nor U16370 (N_16370,N_12320,N_12841);
nor U16371 (N_16371,N_12433,N_12625);
xnor U16372 (N_16372,N_13202,N_14004);
nor U16373 (N_16373,N_14966,N_12847);
or U16374 (N_16374,N_14822,N_13726);
and U16375 (N_16375,N_14713,N_13117);
nand U16376 (N_16376,N_12614,N_12801);
nand U16377 (N_16377,N_13183,N_14266);
or U16378 (N_16378,N_14717,N_12856);
and U16379 (N_16379,N_13445,N_13273);
or U16380 (N_16380,N_12352,N_13663);
or U16381 (N_16381,N_14234,N_14671);
nand U16382 (N_16382,N_14451,N_13702);
nor U16383 (N_16383,N_13912,N_14340);
and U16384 (N_16384,N_13844,N_14700);
nand U16385 (N_16385,N_12282,N_14214);
or U16386 (N_16386,N_14047,N_13593);
nand U16387 (N_16387,N_14142,N_12990);
nand U16388 (N_16388,N_12260,N_12291);
or U16389 (N_16389,N_14063,N_14871);
or U16390 (N_16390,N_12358,N_14861);
xnor U16391 (N_16391,N_14825,N_13228);
or U16392 (N_16392,N_13879,N_14780);
nand U16393 (N_16393,N_13856,N_13812);
or U16394 (N_16394,N_14371,N_13954);
nor U16395 (N_16395,N_12349,N_12795);
and U16396 (N_16396,N_12748,N_12957);
nand U16397 (N_16397,N_13107,N_12945);
and U16398 (N_16398,N_13401,N_13003);
nand U16399 (N_16399,N_13947,N_12046);
and U16400 (N_16400,N_12924,N_12069);
xor U16401 (N_16401,N_14840,N_14135);
nor U16402 (N_16402,N_12962,N_14285);
or U16403 (N_16403,N_14721,N_14433);
or U16404 (N_16404,N_12097,N_14247);
or U16405 (N_16405,N_14985,N_13111);
nor U16406 (N_16406,N_13552,N_12685);
xnor U16407 (N_16407,N_12243,N_14538);
xnor U16408 (N_16408,N_12744,N_13551);
nor U16409 (N_16409,N_14638,N_14318);
nand U16410 (N_16410,N_12633,N_14769);
nand U16411 (N_16411,N_12412,N_13247);
xor U16412 (N_16412,N_12080,N_12102);
or U16413 (N_16413,N_12163,N_12788);
or U16414 (N_16414,N_14766,N_14791);
nand U16415 (N_16415,N_14390,N_12848);
xor U16416 (N_16416,N_12944,N_14246);
nor U16417 (N_16417,N_12630,N_14626);
xor U16418 (N_16418,N_13609,N_14850);
or U16419 (N_16419,N_13421,N_13610);
or U16420 (N_16420,N_14176,N_13618);
nand U16421 (N_16421,N_12452,N_14184);
xor U16422 (N_16422,N_13853,N_13064);
xnor U16423 (N_16423,N_12368,N_13504);
or U16424 (N_16424,N_13864,N_12941);
nor U16425 (N_16425,N_13842,N_14397);
nor U16426 (N_16426,N_12986,N_13033);
xnor U16427 (N_16427,N_12419,N_13823);
nor U16428 (N_16428,N_14093,N_12116);
nand U16429 (N_16429,N_12530,N_12237);
or U16430 (N_16430,N_14278,N_14311);
and U16431 (N_16431,N_13715,N_13615);
and U16432 (N_16432,N_14743,N_12565);
nand U16433 (N_16433,N_12113,N_12153);
and U16434 (N_16434,N_14338,N_12037);
and U16435 (N_16435,N_12925,N_14265);
nor U16436 (N_16436,N_14156,N_13083);
or U16437 (N_16437,N_12012,N_13586);
and U16438 (N_16438,N_13870,N_12367);
or U16439 (N_16439,N_12120,N_13694);
nor U16440 (N_16440,N_12354,N_12918);
nor U16441 (N_16441,N_13524,N_13352);
nand U16442 (N_16442,N_14360,N_13299);
xnor U16443 (N_16443,N_14571,N_14931);
nand U16444 (N_16444,N_12825,N_14829);
nor U16445 (N_16445,N_14240,N_12845);
nand U16446 (N_16446,N_14726,N_12559);
and U16447 (N_16447,N_14678,N_13622);
and U16448 (N_16448,N_14088,N_14744);
nor U16449 (N_16449,N_13662,N_12875);
xnor U16450 (N_16450,N_12509,N_14983);
xor U16451 (N_16451,N_13922,N_12202);
nor U16452 (N_16452,N_14256,N_13316);
and U16453 (N_16453,N_12409,N_12704);
nor U16454 (N_16454,N_12191,N_12954);
or U16455 (N_16455,N_12842,N_14398);
nor U16456 (N_16456,N_12033,N_13887);
or U16457 (N_16457,N_12702,N_14667);
and U16458 (N_16458,N_14061,N_12192);
or U16459 (N_16459,N_13204,N_12167);
xnor U16460 (N_16460,N_12759,N_14767);
nand U16461 (N_16461,N_12540,N_12170);
nand U16462 (N_16462,N_14336,N_12480);
nand U16463 (N_16463,N_14541,N_13814);
or U16464 (N_16464,N_14182,N_14408);
nand U16465 (N_16465,N_14552,N_13225);
xor U16466 (N_16466,N_12900,N_12597);
nor U16467 (N_16467,N_14929,N_13963);
or U16468 (N_16468,N_13040,N_14314);
and U16469 (N_16469,N_12851,N_13304);
and U16470 (N_16470,N_12641,N_14264);
nor U16471 (N_16471,N_13332,N_12083);
nor U16472 (N_16472,N_12893,N_13898);
nand U16473 (N_16473,N_12186,N_13846);
or U16474 (N_16474,N_13238,N_13392);
xor U16475 (N_16475,N_14094,N_14450);
or U16476 (N_16476,N_13056,N_12128);
nand U16477 (N_16477,N_14413,N_14009);
and U16478 (N_16478,N_13976,N_12018);
nor U16479 (N_16479,N_12265,N_12427);
and U16480 (N_16480,N_12461,N_13358);
nand U16481 (N_16481,N_12380,N_13658);
nor U16482 (N_16482,N_13891,N_13208);
nand U16483 (N_16483,N_13946,N_13866);
nor U16484 (N_16484,N_13691,N_12911);
xor U16485 (N_16485,N_12637,N_14437);
nor U16486 (N_16486,N_13365,N_13254);
nor U16487 (N_16487,N_12977,N_13801);
nand U16488 (N_16488,N_13441,N_14755);
and U16489 (N_16489,N_12372,N_12869);
and U16490 (N_16490,N_12818,N_14092);
xnor U16491 (N_16491,N_13383,N_13456);
and U16492 (N_16492,N_13824,N_12346);
nand U16493 (N_16493,N_14683,N_12314);
and U16494 (N_16494,N_12310,N_13882);
nor U16495 (N_16495,N_13537,N_12756);
nand U16496 (N_16496,N_13330,N_14704);
or U16497 (N_16497,N_12822,N_14668);
and U16498 (N_16498,N_13347,N_14597);
or U16499 (N_16499,N_13899,N_13051);
xnor U16500 (N_16500,N_14544,N_14470);
or U16501 (N_16501,N_12646,N_12533);
nand U16502 (N_16502,N_14981,N_14460);
or U16503 (N_16503,N_12043,N_13253);
nor U16504 (N_16504,N_13477,N_13503);
and U16505 (N_16505,N_14557,N_13609);
and U16506 (N_16506,N_14736,N_13875);
xor U16507 (N_16507,N_12821,N_13134);
xnor U16508 (N_16508,N_14313,N_12369);
nand U16509 (N_16509,N_12750,N_13315);
or U16510 (N_16510,N_13682,N_12582);
nor U16511 (N_16511,N_12183,N_13741);
or U16512 (N_16512,N_13724,N_14960);
nand U16513 (N_16513,N_14362,N_14986);
and U16514 (N_16514,N_14149,N_14084);
or U16515 (N_16515,N_14805,N_14148);
and U16516 (N_16516,N_14915,N_13421);
nor U16517 (N_16517,N_14565,N_13583);
nand U16518 (N_16518,N_14135,N_12015);
and U16519 (N_16519,N_13230,N_14388);
nand U16520 (N_16520,N_13553,N_14978);
or U16521 (N_16521,N_13534,N_13590);
or U16522 (N_16522,N_14854,N_14463);
nor U16523 (N_16523,N_14975,N_13773);
nor U16524 (N_16524,N_12401,N_13553);
and U16525 (N_16525,N_14861,N_13733);
nor U16526 (N_16526,N_13970,N_14044);
and U16527 (N_16527,N_14794,N_13717);
and U16528 (N_16528,N_13488,N_14978);
nand U16529 (N_16529,N_12449,N_14798);
and U16530 (N_16530,N_14029,N_14243);
nor U16531 (N_16531,N_12837,N_13607);
or U16532 (N_16532,N_12081,N_13862);
xor U16533 (N_16533,N_13377,N_12577);
or U16534 (N_16534,N_12093,N_14391);
or U16535 (N_16535,N_12514,N_13883);
nand U16536 (N_16536,N_14456,N_14320);
or U16537 (N_16537,N_14217,N_12484);
xor U16538 (N_16538,N_14269,N_14521);
or U16539 (N_16539,N_14297,N_14670);
and U16540 (N_16540,N_12890,N_13844);
nor U16541 (N_16541,N_13487,N_14140);
nor U16542 (N_16542,N_13317,N_13835);
or U16543 (N_16543,N_12794,N_14167);
or U16544 (N_16544,N_13469,N_14859);
and U16545 (N_16545,N_12403,N_14755);
nand U16546 (N_16546,N_13856,N_12874);
or U16547 (N_16547,N_12386,N_14545);
nand U16548 (N_16548,N_13563,N_12542);
xnor U16549 (N_16549,N_12754,N_12660);
or U16550 (N_16550,N_14212,N_14919);
and U16551 (N_16551,N_13805,N_13344);
xor U16552 (N_16552,N_12650,N_14047);
nand U16553 (N_16553,N_12569,N_12173);
and U16554 (N_16554,N_12448,N_12026);
nand U16555 (N_16555,N_13733,N_14807);
nand U16556 (N_16556,N_14466,N_13572);
or U16557 (N_16557,N_14215,N_13872);
nand U16558 (N_16558,N_14433,N_14604);
or U16559 (N_16559,N_12286,N_12167);
xnor U16560 (N_16560,N_12835,N_14107);
or U16561 (N_16561,N_14417,N_13332);
and U16562 (N_16562,N_13165,N_14618);
or U16563 (N_16563,N_14449,N_12769);
xor U16564 (N_16564,N_14836,N_12013);
xnor U16565 (N_16565,N_12842,N_13745);
nand U16566 (N_16566,N_14888,N_13159);
nor U16567 (N_16567,N_13977,N_12361);
and U16568 (N_16568,N_13204,N_13134);
or U16569 (N_16569,N_13349,N_13686);
nand U16570 (N_16570,N_13844,N_14255);
and U16571 (N_16571,N_14925,N_14452);
nor U16572 (N_16572,N_14754,N_12919);
or U16573 (N_16573,N_14226,N_14283);
xor U16574 (N_16574,N_12565,N_14936);
xor U16575 (N_16575,N_13728,N_12575);
and U16576 (N_16576,N_12663,N_14069);
nor U16577 (N_16577,N_14053,N_12880);
and U16578 (N_16578,N_12466,N_12922);
or U16579 (N_16579,N_12488,N_12122);
and U16580 (N_16580,N_12602,N_14436);
nand U16581 (N_16581,N_14601,N_14652);
xor U16582 (N_16582,N_14046,N_13104);
nand U16583 (N_16583,N_14992,N_14960);
nand U16584 (N_16584,N_13620,N_12904);
and U16585 (N_16585,N_13456,N_13541);
or U16586 (N_16586,N_13427,N_13358);
nand U16587 (N_16587,N_14491,N_12451);
xor U16588 (N_16588,N_12967,N_12179);
and U16589 (N_16589,N_13837,N_12884);
nor U16590 (N_16590,N_12233,N_13504);
xor U16591 (N_16591,N_13666,N_12503);
nor U16592 (N_16592,N_13405,N_14350);
and U16593 (N_16593,N_13001,N_13646);
or U16594 (N_16594,N_13642,N_12055);
nor U16595 (N_16595,N_14452,N_14462);
nand U16596 (N_16596,N_12801,N_12369);
or U16597 (N_16597,N_13198,N_14355);
xnor U16598 (N_16598,N_12911,N_13264);
and U16599 (N_16599,N_14237,N_13249);
xnor U16600 (N_16600,N_14684,N_13594);
nor U16601 (N_16601,N_13771,N_14309);
and U16602 (N_16602,N_13435,N_12337);
nor U16603 (N_16603,N_12001,N_14292);
xnor U16604 (N_16604,N_12271,N_12823);
or U16605 (N_16605,N_13994,N_12325);
xor U16606 (N_16606,N_13830,N_12573);
xnor U16607 (N_16607,N_13951,N_13262);
nand U16608 (N_16608,N_12581,N_12210);
and U16609 (N_16609,N_14457,N_14146);
nor U16610 (N_16610,N_14168,N_14105);
nor U16611 (N_16611,N_13111,N_13667);
nor U16612 (N_16612,N_12359,N_12577);
xnor U16613 (N_16613,N_14555,N_12688);
xnor U16614 (N_16614,N_14399,N_14854);
nor U16615 (N_16615,N_13910,N_13965);
and U16616 (N_16616,N_13424,N_14808);
nand U16617 (N_16617,N_13903,N_12191);
nand U16618 (N_16618,N_13313,N_13651);
nand U16619 (N_16619,N_14670,N_14344);
nor U16620 (N_16620,N_14789,N_13193);
xor U16621 (N_16621,N_13535,N_14842);
nand U16622 (N_16622,N_12725,N_14915);
xnor U16623 (N_16623,N_12610,N_13248);
nand U16624 (N_16624,N_12246,N_14793);
or U16625 (N_16625,N_12146,N_12938);
nand U16626 (N_16626,N_13818,N_14929);
nor U16627 (N_16627,N_12425,N_14228);
nor U16628 (N_16628,N_14345,N_12751);
nand U16629 (N_16629,N_13503,N_13942);
and U16630 (N_16630,N_12786,N_13820);
or U16631 (N_16631,N_12628,N_14535);
nor U16632 (N_16632,N_12465,N_14224);
nor U16633 (N_16633,N_12708,N_12539);
or U16634 (N_16634,N_14335,N_12817);
or U16635 (N_16635,N_13598,N_14698);
nand U16636 (N_16636,N_12722,N_14038);
xnor U16637 (N_16637,N_13844,N_14605);
and U16638 (N_16638,N_14151,N_14180);
and U16639 (N_16639,N_13146,N_13123);
or U16640 (N_16640,N_12633,N_12231);
or U16641 (N_16641,N_13959,N_13262);
and U16642 (N_16642,N_14526,N_13753);
nand U16643 (N_16643,N_13084,N_14078);
or U16644 (N_16644,N_12783,N_12291);
xnor U16645 (N_16645,N_13030,N_14492);
and U16646 (N_16646,N_13519,N_14288);
or U16647 (N_16647,N_14077,N_13944);
or U16648 (N_16648,N_12202,N_13540);
and U16649 (N_16649,N_12451,N_12389);
and U16650 (N_16650,N_12235,N_14836);
and U16651 (N_16651,N_13949,N_12056);
nor U16652 (N_16652,N_13165,N_12281);
nand U16653 (N_16653,N_12599,N_13787);
nand U16654 (N_16654,N_14195,N_14628);
or U16655 (N_16655,N_13617,N_12382);
xor U16656 (N_16656,N_14302,N_14969);
xor U16657 (N_16657,N_14852,N_14329);
xor U16658 (N_16658,N_13298,N_12850);
and U16659 (N_16659,N_14874,N_14754);
xor U16660 (N_16660,N_12418,N_14808);
nor U16661 (N_16661,N_12487,N_13817);
nor U16662 (N_16662,N_12845,N_13353);
xnor U16663 (N_16663,N_13629,N_12543);
and U16664 (N_16664,N_12655,N_13831);
nor U16665 (N_16665,N_14150,N_13837);
xnor U16666 (N_16666,N_13292,N_12606);
or U16667 (N_16667,N_14620,N_13306);
or U16668 (N_16668,N_14167,N_13749);
nand U16669 (N_16669,N_12669,N_14122);
xor U16670 (N_16670,N_12202,N_13733);
nor U16671 (N_16671,N_14988,N_13904);
xor U16672 (N_16672,N_13378,N_14540);
and U16673 (N_16673,N_13411,N_14203);
or U16674 (N_16674,N_13030,N_14169);
or U16675 (N_16675,N_12260,N_12390);
nand U16676 (N_16676,N_13087,N_14183);
or U16677 (N_16677,N_12472,N_14168);
and U16678 (N_16678,N_12023,N_13616);
nand U16679 (N_16679,N_12305,N_13127);
or U16680 (N_16680,N_12985,N_12470);
xnor U16681 (N_16681,N_13833,N_14723);
nand U16682 (N_16682,N_14740,N_14072);
and U16683 (N_16683,N_13424,N_12681);
xor U16684 (N_16684,N_12600,N_12144);
or U16685 (N_16685,N_12792,N_14997);
xnor U16686 (N_16686,N_12129,N_12275);
or U16687 (N_16687,N_13989,N_14803);
and U16688 (N_16688,N_12226,N_13837);
or U16689 (N_16689,N_12237,N_14362);
and U16690 (N_16690,N_14132,N_13950);
xnor U16691 (N_16691,N_14449,N_13783);
nor U16692 (N_16692,N_14069,N_13677);
and U16693 (N_16693,N_14502,N_12158);
and U16694 (N_16694,N_13010,N_14030);
xnor U16695 (N_16695,N_12823,N_13421);
or U16696 (N_16696,N_12636,N_13509);
nand U16697 (N_16697,N_12305,N_12347);
xor U16698 (N_16698,N_12784,N_14252);
nand U16699 (N_16699,N_12890,N_12939);
or U16700 (N_16700,N_13560,N_14841);
or U16701 (N_16701,N_12186,N_13812);
or U16702 (N_16702,N_12767,N_14705);
nor U16703 (N_16703,N_13488,N_14148);
or U16704 (N_16704,N_14493,N_12048);
nand U16705 (N_16705,N_14429,N_12622);
or U16706 (N_16706,N_14587,N_13531);
nor U16707 (N_16707,N_14083,N_13044);
nor U16708 (N_16708,N_13786,N_12297);
xnor U16709 (N_16709,N_12838,N_12967);
nand U16710 (N_16710,N_14803,N_14261);
xnor U16711 (N_16711,N_14309,N_14495);
nand U16712 (N_16712,N_14525,N_14596);
and U16713 (N_16713,N_12055,N_12332);
or U16714 (N_16714,N_13203,N_13746);
or U16715 (N_16715,N_12446,N_13272);
and U16716 (N_16716,N_13344,N_14010);
and U16717 (N_16717,N_12954,N_13515);
nor U16718 (N_16718,N_12697,N_13736);
nand U16719 (N_16719,N_14233,N_14866);
nor U16720 (N_16720,N_14173,N_12552);
and U16721 (N_16721,N_13586,N_12358);
nand U16722 (N_16722,N_12224,N_13630);
and U16723 (N_16723,N_12547,N_14241);
nor U16724 (N_16724,N_13222,N_12423);
or U16725 (N_16725,N_14032,N_14557);
nor U16726 (N_16726,N_14428,N_12579);
nand U16727 (N_16727,N_14034,N_13053);
and U16728 (N_16728,N_13123,N_13700);
and U16729 (N_16729,N_14710,N_13630);
xor U16730 (N_16730,N_12714,N_14837);
xor U16731 (N_16731,N_13160,N_13547);
or U16732 (N_16732,N_13262,N_13364);
or U16733 (N_16733,N_14471,N_14425);
nand U16734 (N_16734,N_14600,N_14950);
nand U16735 (N_16735,N_12541,N_14410);
and U16736 (N_16736,N_12321,N_14490);
nor U16737 (N_16737,N_12279,N_12329);
and U16738 (N_16738,N_12998,N_13196);
xor U16739 (N_16739,N_14722,N_12864);
nor U16740 (N_16740,N_12265,N_12625);
xnor U16741 (N_16741,N_12323,N_12343);
nor U16742 (N_16742,N_14741,N_13796);
or U16743 (N_16743,N_14278,N_14196);
or U16744 (N_16744,N_13845,N_12860);
or U16745 (N_16745,N_14156,N_14712);
nor U16746 (N_16746,N_12820,N_12653);
or U16747 (N_16747,N_13240,N_14435);
nor U16748 (N_16748,N_13408,N_13134);
or U16749 (N_16749,N_13715,N_14363);
or U16750 (N_16750,N_13674,N_12485);
or U16751 (N_16751,N_12304,N_13433);
nor U16752 (N_16752,N_12876,N_13933);
and U16753 (N_16753,N_12521,N_12865);
or U16754 (N_16754,N_14909,N_14927);
nor U16755 (N_16755,N_13105,N_13280);
and U16756 (N_16756,N_12443,N_14036);
and U16757 (N_16757,N_13670,N_14071);
xnor U16758 (N_16758,N_12914,N_13381);
nor U16759 (N_16759,N_12605,N_14311);
nand U16760 (N_16760,N_12870,N_14226);
xor U16761 (N_16761,N_14949,N_13390);
xnor U16762 (N_16762,N_12393,N_13343);
xnor U16763 (N_16763,N_14442,N_12981);
xnor U16764 (N_16764,N_13377,N_12564);
and U16765 (N_16765,N_14228,N_12587);
xnor U16766 (N_16766,N_12812,N_14776);
and U16767 (N_16767,N_13438,N_13750);
nand U16768 (N_16768,N_13699,N_12513);
and U16769 (N_16769,N_12345,N_14824);
and U16770 (N_16770,N_14809,N_12196);
nand U16771 (N_16771,N_13989,N_13653);
or U16772 (N_16772,N_14594,N_12907);
xnor U16773 (N_16773,N_14229,N_14175);
nand U16774 (N_16774,N_14349,N_12008);
nand U16775 (N_16775,N_13158,N_12450);
xor U16776 (N_16776,N_13632,N_12469);
or U16777 (N_16777,N_14515,N_12422);
nor U16778 (N_16778,N_12340,N_13110);
xor U16779 (N_16779,N_13995,N_12392);
xor U16780 (N_16780,N_12796,N_14943);
xnor U16781 (N_16781,N_12558,N_13831);
xor U16782 (N_16782,N_14447,N_12435);
nand U16783 (N_16783,N_14704,N_13546);
and U16784 (N_16784,N_14687,N_13704);
nand U16785 (N_16785,N_12560,N_12833);
nand U16786 (N_16786,N_14580,N_13002);
or U16787 (N_16787,N_12997,N_14120);
and U16788 (N_16788,N_13438,N_12384);
nand U16789 (N_16789,N_13675,N_12523);
nor U16790 (N_16790,N_12967,N_14648);
and U16791 (N_16791,N_13493,N_13942);
and U16792 (N_16792,N_14655,N_14559);
nand U16793 (N_16793,N_13537,N_12290);
xor U16794 (N_16794,N_13048,N_12811);
nand U16795 (N_16795,N_14412,N_13709);
and U16796 (N_16796,N_13712,N_13620);
nand U16797 (N_16797,N_14364,N_12259);
xor U16798 (N_16798,N_12725,N_13117);
xor U16799 (N_16799,N_12609,N_13787);
nand U16800 (N_16800,N_12741,N_14651);
or U16801 (N_16801,N_12368,N_14320);
nand U16802 (N_16802,N_13226,N_12107);
or U16803 (N_16803,N_13870,N_14385);
xnor U16804 (N_16804,N_12308,N_14564);
xnor U16805 (N_16805,N_12664,N_14901);
nor U16806 (N_16806,N_13365,N_14169);
nor U16807 (N_16807,N_12091,N_13923);
and U16808 (N_16808,N_13498,N_13231);
xnor U16809 (N_16809,N_12324,N_13015);
or U16810 (N_16810,N_14082,N_12203);
xnor U16811 (N_16811,N_13401,N_13315);
and U16812 (N_16812,N_14452,N_13587);
and U16813 (N_16813,N_14124,N_14156);
nand U16814 (N_16814,N_13028,N_14004);
xnor U16815 (N_16815,N_12325,N_13138);
or U16816 (N_16816,N_12851,N_14188);
nor U16817 (N_16817,N_13511,N_14634);
nor U16818 (N_16818,N_12948,N_13890);
nand U16819 (N_16819,N_12760,N_13763);
or U16820 (N_16820,N_13569,N_13576);
nor U16821 (N_16821,N_13696,N_12901);
nor U16822 (N_16822,N_13401,N_14043);
nor U16823 (N_16823,N_13368,N_12019);
xor U16824 (N_16824,N_14402,N_13834);
xor U16825 (N_16825,N_14881,N_13803);
xnor U16826 (N_16826,N_12211,N_14862);
xor U16827 (N_16827,N_12892,N_13957);
nand U16828 (N_16828,N_12923,N_14984);
nor U16829 (N_16829,N_12628,N_14069);
nor U16830 (N_16830,N_12925,N_14870);
nor U16831 (N_16831,N_14358,N_13263);
nand U16832 (N_16832,N_13452,N_12433);
nand U16833 (N_16833,N_13976,N_13436);
xnor U16834 (N_16834,N_13134,N_12677);
nand U16835 (N_16835,N_14896,N_13302);
and U16836 (N_16836,N_12684,N_12918);
and U16837 (N_16837,N_14157,N_13872);
nand U16838 (N_16838,N_14121,N_14327);
xor U16839 (N_16839,N_13507,N_13803);
or U16840 (N_16840,N_13591,N_13313);
xor U16841 (N_16841,N_12436,N_12347);
or U16842 (N_16842,N_13912,N_13058);
or U16843 (N_16843,N_14027,N_14816);
nor U16844 (N_16844,N_13887,N_12072);
nand U16845 (N_16845,N_14580,N_13544);
xor U16846 (N_16846,N_12609,N_13913);
nand U16847 (N_16847,N_14001,N_13200);
or U16848 (N_16848,N_14861,N_14252);
and U16849 (N_16849,N_13789,N_14835);
or U16850 (N_16850,N_14578,N_13743);
or U16851 (N_16851,N_13025,N_14113);
or U16852 (N_16852,N_12252,N_14010);
nor U16853 (N_16853,N_12007,N_13775);
and U16854 (N_16854,N_14548,N_12499);
nand U16855 (N_16855,N_12682,N_12466);
xor U16856 (N_16856,N_14876,N_12005);
nor U16857 (N_16857,N_12360,N_14372);
xnor U16858 (N_16858,N_13482,N_12237);
nor U16859 (N_16859,N_13709,N_14862);
xnor U16860 (N_16860,N_13909,N_14654);
nand U16861 (N_16861,N_12799,N_13877);
or U16862 (N_16862,N_13524,N_14478);
or U16863 (N_16863,N_13981,N_14000);
nor U16864 (N_16864,N_13833,N_12548);
and U16865 (N_16865,N_13493,N_12769);
nand U16866 (N_16866,N_13473,N_13403);
and U16867 (N_16867,N_12183,N_12643);
and U16868 (N_16868,N_13206,N_12780);
nand U16869 (N_16869,N_13268,N_13270);
and U16870 (N_16870,N_13931,N_14905);
nor U16871 (N_16871,N_14425,N_13164);
nand U16872 (N_16872,N_13968,N_12351);
nor U16873 (N_16873,N_13869,N_13159);
nand U16874 (N_16874,N_14390,N_13991);
nand U16875 (N_16875,N_14521,N_14562);
or U16876 (N_16876,N_14597,N_13232);
nand U16877 (N_16877,N_12763,N_13805);
xor U16878 (N_16878,N_14871,N_14600);
or U16879 (N_16879,N_13504,N_13318);
xor U16880 (N_16880,N_14730,N_14946);
xnor U16881 (N_16881,N_13515,N_13935);
and U16882 (N_16882,N_14133,N_14661);
and U16883 (N_16883,N_14828,N_14047);
and U16884 (N_16884,N_13486,N_13237);
or U16885 (N_16885,N_12131,N_12598);
or U16886 (N_16886,N_14009,N_13743);
xnor U16887 (N_16887,N_14657,N_14149);
and U16888 (N_16888,N_14335,N_12850);
nor U16889 (N_16889,N_14979,N_14840);
and U16890 (N_16890,N_14261,N_14534);
and U16891 (N_16891,N_12849,N_12939);
nand U16892 (N_16892,N_12253,N_12311);
or U16893 (N_16893,N_14450,N_13447);
and U16894 (N_16894,N_12454,N_12033);
or U16895 (N_16895,N_14818,N_12508);
xnor U16896 (N_16896,N_14922,N_14565);
and U16897 (N_16897,N_14273,N_14926);
nor U16898 (N_16898,N_12962,N_12217);
nor U16899 (N_16899,N_12983,N_14245);
nand U16900 (N_16900,N_14571,N_14015);
nand U16901 (N_16901,N_12083,N_12006);
or U16902 (N_16902,N_13060,N_13269);
nor U16903 (N_16903,N_12386,N_14146);
nor U16904 (N_16904,N_12921,N_12547);
or U16905 (N_16905,N_12928,N_12030);
or U16906 (N_16906,N_12854,N_14915);
and U16907 (N_16907,N_12171,N_14742);
nor U16908 (N_16908,N_12344,N_14619);
nor U16909 (N_16909,N_13954,N_12023);
and U16910 (N_16910,N_12242,N_12980);
nor U16911 (N_16911,N_14635,N_13312);
xnor U16912 (N_16912,N_12732,N_14655);
nand U16913 (N_16913,N_12485,N_13284);
nor U16914 (N_16914,N_12145,N_13432);
and U16915 (N_16915,N_12172,N_13026);
nor U16916 (N_16916,N_12465,N_12498);
nand U16917 (N_16917,N_13288,N_13858);
nand U16918 (N_16918,N_14195,N_12749);
xnor U16919 (N_16919,N_12249,N_12650);
and U16920 (N_16920,N_12124,N_13690);
and U16921 (N_16921,N_14584,N_13426);
nor U16922 (N_16922,N_12833,N_14244);
or U16923 (N_16923,N_13960,N_14773);
nand U16924 (N_16924,N_13854,N_12529);
xnor U16925 (N_16925,N_13336,N_13579);
nand U16926 (N_16926,N_13137,N_13697);
and U16927 (N_16927,N_14323,N_12461);
and U16928 (N_16928,N_13397,N_12601);
or U16929 (N_16929,N_12191,N_12081);
or U16930 (N_16930,N_14516,N_14504);
and U16931 (N_16931,N_13043,N_13169);
nand U16932 (N_16932,N_12777,N_12497);
xnor U16933 (N_16933,N_14686,N_14988);
nand U16934 (N_16934,N_12546,N_14296);
and U16935 (N_16935,N_13797,N_12007);
and U16936 (N_16936,N_12531,N_13580);
or U16937 (N_16937,N_14810,N_12132);
or U16938 (N_16938,N_12028,N_12358);
xnor U16939 (N_16939,N_13123,N_13002);
xor U16940 (N_16940,N_14897,N_14407);
nor U16941 (N_16941,N_14519,N_13233);
nand U16942 (N_16942,N_12633,N_13271);
nand U16943 (N_16943,N_14564,N_12514);
nand U16944 (N_16944,N_12393,N_12017);
nor U16945 (N_16945,N_13285,N_12361);
and U16946 (N_16946,N_12424,N_13835);
nor U16947 (N_16947,N_12746,N_13464);
nor U16948 (N_16948,N_14599,N_14486);
or U16949 (N_16949,N_12884,N_13826);
nand U16950 (N_16950,N_13005,N_12309);
nor U16951 (N_16951,N_13651,N_13700);
nor U16952 (N_16952,N_14094,N_13109);
nor U16953 (N_16953,N_12802,N_13814);
xor U16954 (N_16954,N_12058,N_14626);
xor U16955 (N_16955,N_12005,N_14717);
xnor U16956 (N_16956,N_13277,N_12052);
xor U16957 (N_16957,N_12718,N_13876);
nor U16958 (N_16958,N_14359,N_14667);
nor U16959 (N_16959,N_12226,N_13107);
nor U16960 (N_16960,N_14247,N_14079);
and U16961 (N_16961,N_13522,N_14400);
nor U16962 (N_16962,N_13905,N_13181);
nand U16963 (N_16963,N_13843,N_13274);
xor U16964 (N_16964,N_12996,N_14816);
nor U16965 (N_16965,N_14395,N_12608);
nand U16966 (N_16966,N_12778,N_14301);
and U16967 (N_16967,N_13656,N_12334);
xnor U16968 (N_16968,N_12054,N_13313);
and U16969 (N_16969,N_13022,N_14262);
xor U16970 (N_16970,N_14540,N_14141);
nand U16971 (N_16971,N_14596,N_12693);
xnor U16972 (N_16972,N_12366,N_13143);
and U16973 (N_16973,N_12669,N_14828);
and U16974 (N_16974,N_13995,N_14262);
and U16975 (N_16975,N_12935,N_14454);
or U16976 (N_16976,N_12322,N_13095);
and U16977 (N_16977,N_14683,N_14858);
nor U16978 (N_16978,N_14767,N_12172);
or U16979 (N_16979,N_12707,N_13057);
and U16980 (N_16980,N_14819,N_12854);
or U16981 (N_16981,N_13896,N_12728);
xor U16982 (N_16982,N_12207,N_13004);
xor U16983 (N_16983,N_14583,N_14515);
nand U16984 (N_16984,N_12025,N_13692);
nor U16985 (N_16985,N_14842,N_12650);
and U16986 (N_16986,N_14336,N_13892);
and U16987 (N_16987,N_13635,N_12432);
or U16988 (N_16988,N_13541,N_12585);
xor U16989 (N_16989,N_14429,N_12435);
and U16990 (N_16990,N_13344,N_14365);
xor U16991 (N_16991,N_14432,N_13463);
nand U16992 (N_16992,N_12101,N_13788);
nand U16993 (N_16993,N_14783,N_13612);
or U16994 (N_16994,N_12392,N_13406);
and U16995 (N_16995,N_14019,N_14347);
or U16996 (N_16996,N_14823,N_14958);
nand U16997 (N_16997,N_13902,N_12750);
xor U16998 (N_16998,N_12236,N_12269);
nand U16999 (N_16999,N_13506,N_13360);
xor U17000 (N_17000,N_12056,N_13280);
or U17001 (N_17001,N_12569,N_13683);
nor U17002 (N_17002,N_12843,N_14956);
or U17003 (N_17003,N_12450,N_13407);
xnor U17004 (N_17004,N_13214,N_12866);
and U17005 (N_17005,N_14520,N_12256);
nor U17006 (N_17006,N_14517,N_14990);
or U17007 (N_17007,N_14898,N_13582);
nor U17008 (N_17008,N_13582,N_12729);
nor U17009 (N_17009,N_13265,N_14856);
nor U17010 (N_17010,N_14508,N_14820);
xnor U17011 (N_17011,N_14192,N_12040);
or U17012 (N_17012,N_12329,N_14790);
or U17013 (N_17013,N_12302,N_12702);
or U17014 (N_17014,N_13199,N_12842);
or U17015 (N_17015,N_13625,N_14597);
nor U17016 (N_17016,N_14705,N_13755);
and U17017 (N_17017,N_13774,N_12134);
or U17018 (N_17018,N_13675,N_13558);
xor U17019 (N_17019,N_13358,N_14862);
and U17020 (N_17020,N_13376,N_13446);
xor U17021 (N_17021,N_13991,N_13193);
nand U17022 (N_17022,N_14409,N_12431);
nand U17023 (N_17023,N_14362,N_14803);
xor U17024 (N_17024,N_12694,N_12330);
xor U17025 (N_17025,N_12073,N_13727);
nand U17026 (N_17026,N_14982,N_13387);
xnor U17027 (N_17027,N_13180,N_13087);
and U17028 (N_17028,N_12651,N_12455);
and U17029 (N_17029,N_14052,N_13428);
or U17030 (N_17030,N_12778,N_14784);
xor U17031 (N_17031,N_13887,N_12038);
xnor U17032 (N_17032,N_12170,N_13468);
or U17033 (N_17033,N_13598,N_12362);
and U17034 (N_17034,N_13127,N_13954);
or U17035 (N_17035,N_14585,N_13423);
nand U17036 (N_17036,N_12450,N_12569);
nor U17037 (N_17037,N_12090,N_14896);
nor U17038 (N_17038,N_13753,N_12409);
xnor U17039 (N_17039,N_13070,N_12022);
nor U17040 (N_17040,N_13000,N_12281);
xor U17041 (N_17041,N_12010,N_14745);
and U17042 (N_17042,N_14831,N_14340);
nor U17043 (N_17043,N_13154,N_14241);
or U17044 (N_17044,N_12201,N_14558);
nor U17045 (N_17045,N_12452,N_12705);
and U17046 (N_17046,N_14607,N_12107);
nor U17047 (N_17047,N_12504,N_14790);
nand U17048 (N_17048,N_13589,N_14081);
nand U17049 (N_17049,N_12659,N_13475);
xor U17050 (N_17050,N_14485,N_14733);
and U17051 (N_17051,N_12987,N_12479);
xor U17052 (N_17052,N_13001,N_14315);
and U17053 (N_17053,N_14142,N_13007);
and U17054 (N_17054,N_14784,N_14057);
nand U17055 (N_17055,N_12649,N_14654);
nor U17056 (N_17056,N_14928,N_12280);
nand U17057 (N_17057,N_12672,N_12070);
and U17058 (N_17058,N_14005,N_14127);
nor U17059 (N_17059,N_13967,N_12143);
or U17060 (N_17060,N_14908,N_12274);
or U17061 (N_17061,N_12320,N_12806);
nand U17062 (N_17062,N_12806,N_13598);
or U17063 (N_17063,N_13549,N_14060);
nand U17064 (N_17064,N_13314,N_13975);
xnor U17065 (N_17065,N_13907,N_12452);
xor U17066 (N_17066,N_13151,N_14755);
nor U17067 (N_17067,N_13417,N_12975);
nand U17068 (N_17068,N_13048,N_14390);
and U17069 (N_17069,N_14966,N_14822);
and U17070 (N_17070,N_14285,N_14253);
nor U17071 (N_17071,N_14374,N_14012);
nor U17072 (N_17072,N_13171,N_14188);
nor U17073 (N_17073,N_14316,N_13393);
nand U17074 (N_17074,N_12125,N_14577);
or U17075 (N_17075,N_12352,N_12317);
or U17076 (N_17076,N_13967,N_12653);
and U17077 (N_17077,N_14724,N_12555);
or U17078 (N_17078,N_14186,N_13451);
or U17079 (N_17079,N_12789,N_14868);
or U17080 (N_17080,N_12070,N_13774);
and U17081 (N_17081,N_12120,N_14476);
or U17082 (N_17082,N_13551,N_14798);
nand U17083 (N_17083,N_12262,N_14789);
nor U17084 (N_17084,N_12974,N_12692);
xnor U17085 (N_17085,N_14628,N_13189);
or U17086 (N_17086,N_13580,N_14933);
nand U17087 (N_17087,N_14626,N_12959);
xor U17088 (N_17088,N_13647,N_12939);
or U17089 (N_17089,N_12901,N_12427);
nand U17090 (N_17090,N_12201,N_12961);
nor U17091 (N_17091,N_14282,N_13058);
nor U17092 (N_17092,N_12274,N_12517);
nor U17093 (N_17093,N_14009,N_14550);
and U17094 (N_17094,N_14314,N_13421);
xor U17095 (N_17095,N_14865,N_12000);
or U17096 (N_17096,N_12371,N_14138);
xnor U17097 (N_17097,N_14559,N_14293);
or U17098 (N_17098,N_12055,N_12807);
and U17099 (N_17099,N_12403,N_12470);
nor U17100 (N_17100,N_14917,N_12432);
xnor U17101 (N_17101,N_13832,N_14548);
and U17102 (N_17102,N_12085,N_13359);
or U17103 (N_17103,N_13047,N_12282);
or U17104 (N_17104,N_14223,N_12320);
nor U17105 (N_17105,N_12543,N_12107);
nand U17106 (N_17106,N_12215,N_14855);
and U17107 (N_17107,N_14182,N_13390);
nand U17108 (N_17108,N_12103,N_14268);
or U17109 (N_17109,N_13631,N_14977);
and U17110 (N_17110,N_12036,N_13645);
or U17111 (N_17111,N_13548,N_13485);
and U17112 (N_17112,N_14239,N_13958);
nor U17113 (N_17113,N_13812,N_13838);
nor U17114 (N_17114,N_13459,N_13971);
nor U17115 (N_17115,N_12043,N_14351);
and U17116 (N_17116,N_12955,N_14623);
nor U17117 (N_17117,N_13147,N_14649);
or U17118 (N_17118,N_14770,N_13941);
nor U17119 (N_17119,N_14802,N_13734);
xnor U17120 (N_17120,N_12850,N_13105);
xnor U17121 (N_17121,N_14435,N_13413);
nor U17122 (N_17122,N_13900,N_12297);
nand U17123 (N_17123,N_14406,N_13069);
nor U17124 (N_17124,N_14976,N_12117);
nand U17125 (N_17125,N_13164,N_14575);
nor U17126 (N_17126,N_14482,N_13624);
and U17127 (N_17127,N_12428,N_13888);
and U17128 (N_17128,N_12722,N_12099);
nand U17129 (N_17129,N_12959,N_13905);
xor U17130 (N_17130,N_14572,N_14566);
xnor U17131 (N_17131,N_14383,N_14875);
xnor U17132 (N_17132,N_12442,N_13322);
nand U17133 (N_17133,N_13629,N_13543);
nand U17134 (N_17134,N_14167,N_14235);
or U17135 (N_17135,N_12439,N_14275);
xnor U17136 (N_17136,N_13201,N_14621);
nand U17137 (N_17137,N_14195,N_12071);
and U17138 (N_17138,N_14757,N_13687);
or U17139 (N_17139,N_13488,N_14751);
nand U17140 (N_17140,N_14858,N_14309);
or U17141 (N_17141,N_14720,N_13551);
xnor U17142 (N_17142,N_13217,N_14637);
nand U17143 (N_17143,N_14984,N_13714);
nor U17144 (N_17144,N_13428,N_12874);
and U17145 (N_17145,N_12045,N_12038);
xor U17146 (N_17146,N_12422,N_14847);
and U17147 (N_17147,N_12450,N_14532);
or U17148 (N_17148,N_14545,N_13019);
nand U17149 (N_17149,N_13923,N_14625);
nor U17150 (N_17150,N_14618,N_13781);
xnor U17151 (N_17151,N_12296,N_14132);
and U17152 (N_17152,N_14742,N_12282);
nand U17153 (N_17153,N_14839,N_12372);
and U17154 (N_17154,N_13847,N_12809);
and U17155 (N_17155,N_13455,N_13061);
and U17156 (N_17156,N_12508,N_12633);
nor U17157 (N_17157,N_13531,N_12479);
and U17158 (N_17158,N_14259,N_13998);
or U17159 (N_17159,N_12456,N_14967);
nor U17160 (N_17160,N_14405,N_13379);
nor U17161 (N_17161,N_14836,N_13973);
xor U17162 (N_17162,N_13665,N_12625);
xor U17163 (N_17163,N_14846,N_12908);
xor U17164 (N_17164,N_13965,N_13599);
or U17165 (N_17165,N_13463,N_13130);
nand U17166 (N_17166,N_12678,N_13659);
nor U17167 (N_17167,N_14308,N_13974);
and U17168 (N_17168,N_13471,N_12557);
nand U17169 (N_17169,N_12946,N_13666);
xnor U17170 (N_17170,N_14969,N_12129);
or U17171 (N_17171,N_14648,N_13977);
nor U17172 (N_17172,N_13476,N_13416);
xor U17173 (N_17173,N_12568,N_12023);
nor U17174 (N_17174,N_14452,N_14690);
nand U17175 (N_17175,N_13487,N_14285);
nor U17176 (N_17176,N_13768,N_12667);
xnor U17177 (N_17177,N_12481,N_14268);
xor U17178 (N_17178,N_12453,N_12683);
xnor U17179 (N_17179,N_14891,N_12950);
xor U17180 (N_17180,N_14608,N_12249);
nand U17181 (N_17181,N_14969,N_13197);
nand U17182 (N_17182,N_13238,N_12157);
nand U17183 (N_17183,N_12675,N_12118);
and U17184 (N_17184,N_12377,N_13140);
and U17185 (N_17185,N_12586,N_12341);
nor U17186 (N_17186,N_13289,N_13389);
nand U17187 (N_17187,N_14624,N_13513);
xnor U17188 (N_17188,N_14510,N_14759);
xor U17189 (N_17189,N_12450,N_12247);
nor U17190 (N_17190,N_12571,N_13355);
xnor U17191 (N_17191,N_12716,N_12243);
and U17192 (N_17192,N_13182,N_13968);
nand U17193 (N_17193,N_14860,N_13557);
nand U17194 (N_17194,N_12247,N_12953);
xnor U17195 (N_17195,N_14403,N_13731);
and U17196 (N_17196,N_14493,N_14131);
nor U17197 (N_17197,N_13096,N_12009);
xor U17198 (N_17198,N_14394,N_12847);
nor U17199 (N_17199,N_12550,N_14976);
nor U17200 (N_17200,N_12859,N_12987);
or U17201 (N_17201,N_13113,N_13813);
nor U17202 (N_17202,N_14939,N_14204);
and U17203 (N_17203,N_12391,N_14070);
nor U17204 (N_17204,N_13460,N_13637);
nand U17205 (N_17205,N_13300,N_13018);
or U17206 (N_17206,N_12277,N_12822);
or U17207 (N_17207,N_13011,N_13223);
nand U17208 (N_17208,N_14917,N_14955);
xor U17209 (N_17209,N_13292,N_14333);
xnor U17210 (N_17210,N_13119,N_12906);
nor U17211 (N_17211,N_14982,N_12167);
nand U17212 (N_17212,N_13940,N_13847);
nor U17213 (N_17213,N_14434,N_14068);
xnor U17214 (N_17214,N_14320,N_12577);
xor U17215 (N_17215,N_14064,N_13740);
nand U17216 (N_17216,N_13619,N_13968);
and U17217 (N_17217,N_14916,N_12980);
and U17218 (N_17218,N_14141,N_14954);
and U17219 (N_17219,N_13546,N_12070);
xor U17220 (N_17220,N_13652,N_12688);
xnor U17221 (N_17221,N_13017,N_12100);
nor U17222 (N_17222,N_12767,N_12452);
and U17223 (N_17223,N_13114,N_14014);
xor U17224 (N_17224,N_12381,N_13844);
nand U17225 (N_17225,N_12447,N_13275);
and U17226 (N_17226,N_12601,N_14325);
nand U17227 (N_17227,N_14316,N_12156);
or U17228 (N_17228,N_14144,N_12268);
nor U17229 (N_17229,N_14668,N_12447);
or U17230 (N_17230,N_14238,N_14742);
xor U17231 (N_17231,N_12572,N_13546);
nor U17232 (N_17232,N_12013,N_14239);
or U17233 (N_17233,N_13359,N_14482);
nand U17234 (N_17234,N_14416,N_12363);
nand U17235 (N_17235,N_14912,N_14944);
or U17236 (N_17236,N_14900,N_14321);
xor U17237 (N_17237,N_14893,N_13400);
nand U17238 (N_17238,N_12422,N_13236);
xor U17239 (N_17239,N_12169,N_13442);
nor U17240 (N_17240,N_12887,N_14951);
nor U17241 (N_17241,N_14580,N_14491);
or U17242 (N_17242,N_14329,N_14369);
and U17243 (N_17243,N_14901,N_14936);
nand U17244 (N_17244,N_13193,N_13079);
or U17245 (N_17245,N_13791,N_14862);
and U17246 (N_17246,N_14326,N_12738);
or U17247 (N_17247,N_14709,N_14619);
or U17248 (N_17248,N_12283,N_13592);
xnor U17249 (N_17249,N_14765,N_12542);
xor U17250 (N_17250,N_12536,N_12695);
nand U17251 (N_17251,N_12135,N_12632);
nor U17252 (N_17252,N_14754,N_12276);
xnor U17253 (N_17253,N_12558,N_14164);
nand U17254 (N_17254,N_12226,N_12789);
xor U17255 (N_17255,N_14475,N_13461);
xnor U17256 (N_17256,N_13121,N_13390);
or U17257 (N_17257,N_12747,N_14789);
xor U17258 (N_17258,N_13822,N_13813);
or U17259 (N_17259,N_13602,N_12054);
nor U17260 (N_17260,N_12077,N_13342);
or U17261 (N_17261,N_12423,N_13509);
xor U17262 (N_17262,N_12746,N_13365);
or U17263 (N_17263,N_13147,N_13295);
and U17264 (N_17264,N_12663,N_14468);
xnor U17265 (N_17265,N_13487,N_13516);
xnor U17266 (N_17266,N_14866,N_14806);
nand U17267 (N_17267,N_14425,N_12975);
and U17268 (N_17268,N_13690,N_14918);
and U17269 (N_17269,N_13668,N_13712);
nor U17270 (N_17270,N_12299,N_13712);
or U17271 (N_17271,N_12365,N_13452);
xnor U17272 (N_17272,N_14680,N_12514);
nand U17273 (N_17273,N_13288,N_14294);
and U17274 (N_17274,N_14412,N_14697);
nor U17275 (N_17275,N_12162,N_12023);
nor U17276 (N_17276,N_14563,N_13835);
xnor U17277 (N_17277,N_14154,N_13424);
nand U17278 (N_17278,N_13926,N_14627);
xnor U17279 (N_17279,N_14503,N_13445);
or U17280 (N_17280,N_14490,N_13910);
or U17281 (N_17281,N_14283,N_12166);
and U17282 (N_17282,N_13918,N_13059);
nor U17283 (N_17283,N_12143,N_14783);
xor U17284 (N_17284,N_12739,N_12116);
or U17285 (N_17285,N_14724,N_13385);
nor U17286 (N_17286,N_12753,N_13578);
and U17287 (N_17287,N_12559,N_12472);
and U17288 (N_17288,N_13376,N_12354);
nand U17289 (N_17289,N_12671,N_14607);
nand U17290 (N_17290,N_12332,N_13497);
or U17291 (N_17291,N_12050,N_14938);
and U17292 (N_17292,N_13174,N_14858);
and U17293 (N_17293,N_12380,N_13812);
and U17294 (N_17294,N_12154,N_13015);
nand U17295 (N_17295,N_14602,N_14729);
or U17296 (N_17296,N_12514,N_13677);
and U17297 (N_17297,N_14589,N_13590);
nor U17298 (N_17298,N_14628,N_12479);
or U17299 (N_17299,N_12373,N_14755);
nand U17300 (N_17300,N_13198,N_13402);
or U17301 (N_17301,N_13962,N_12644);
nand U17302 (N_17302,N_12271,N_14891);
or U17303 (N_17303,N_12131,N_13510);
or U17304 (N_17304,N_14601,N_13058);
and U17305 (N_17305,N_14338,N_12259);
nor U17306 (N_17306,N_13201,N_12311);
nor U17307 (N_17307,N_14923,N_13721);
nand U17308 (N_17308,N_13716,N_14040);
or U17309 (N_17309,N_14244,N_14419);
xor U17310 (N_17310,N_13356,N_14691);
nand U17311 (N_17311,N_12181,N_14879);
or U17312 (N_17312,N_14736,N_13225);
or U17313 (N_17313,N_14540,N_12960);
or U17314 (N_17314,N_14204,N_12806);
or U17315 (N_17315,N_14626,N_12138);
or U17316 (N_17316,N_13382,N_13698);
nor U17317 (N_17317,N_13518,N_14581);
nor U17318 (N_17318,N_12551,N_14421);
xor U17319 (N_17319,N_14233,N_14980);
and U17320 (N_17320,N_12181,N_12739);
xnor U17321 (N_17321,N_12991,N_14093);
or U17322 (N_17322,N_12866,N_14463);
nor U17323 (N_17323,N_12872,N_13518);
xnor U17324 (N_17324,N_13982,N_14043);
nor U17325 (N_17325,N_12874,N_14773);
nor U17326 (N_17326,N_13513,N_12914);
and U17327 (N_17327,N_14492,N_12340);
nand U17328 (N_17328,N_14849,N_12067);
or U17329 (N_17329,N_14816,N_14137);
xnor U17330 (N_17330,N_14421,N_14870);
or U17331 (N_17331,N_14502,N_13248);
or U17332 (N_17332,N_14858,N_14955);
nor U17333 (N_17333,N_14821,N_14261);
xor U17334 (N_17334,N_13837,N_12019);
nand U17335 (N_17335,N_14030,N_14258);
nor U17336 (N_17336,N_12204,N_12532);
or U17337 (N_17337,N_14725,N_13331);
xor U17338 (N_17338,N_12811,N_13211);
or U17339 (N_17339,N_12143,N_14300);
or U17340 (N_17340,N_14344,N_14302);
nor U17341 (N_17341,N_13467,N_12231);
and U17342 (N_17342,N_13862,N_14560);
or U17343 (N_17343,N_13074,N_12787);
xnor U17344 (N_17344,N_14983,N_13552);
nor U17345 (N_17345,N_12563,N_13860);
and U17346 (N_17346,N_14678,N_13763);
nand U17347 (N_17347,N_12499,N_13584);
nor U17348 (N_17348,N_13452,N_14825);
and U17349 (N_17349,N_14310,N_13178);
and U17350 (N_17350,N_13253,N_12868);
xor U17351 (N_17351,N_13452,N_14794);
or U17352 (N_17352,N_13761,N_12201);
or U17353 (N_17353,N_14978,N_14193);
and U17354 (N_17354,N_13449,N_12588);
nor U17355 (N_17355,N_12403,N_13183);
or U17356 (N_17356,N_13048,N_13686);
nand U17357 (N_17357,N_12956,N_12746);
nand U17358 (N_17358,N_12486,N_13341);
nor U17359 (N_17359,N_13303,N_13527);
or U17360 (N_17360,N_12420,N_14577);
nand U17361 (N_17361,N_14566,N_14495);
or U17362 (N_17362,N_13484,N_13324);
or U17363 (N_17363,N_14932,N_14429);
or U17364 (N_17364,N_13783,N_13748);
xor U17365 (N_17365,N_14266,N_12086);
nand U17366 (N_17366,N_12157,N_13086);
nand U17367 (N_17367,N_12159,N_12217);
and U17368 (N_17368,N_12755,N_13075);
nand U17369 (N_17369,N_13230,N_13244);
nor U17370 (N_17370,N_13193,N_13071);
nor U17371 (N_17371,N_14630,N_12096);
and U17372 (N_17372,N_14945,N_12303);
xnor U17373 (N_17373,N_14488,N_14479);
nor U17374 (N_17374,N_13322,N_12121);
and U17375 (N_17375,N_12269,N_13911);
or U17376 (N_17376,N_12270,N_14129);
or U17377 (N_17377,N_13172,N_12022);
nand U17378 (N_17378,N_14004,N_12807);
xor U17379 (N_17379,N_14478,N_13297);
xnor U17380 (N_17380,N_13224,N_12513);
nand U17381 (N_17381,N_13717,N_12989);
nand U17382 (N_17382,N_14276,N_12639);
and U17383 (N_17383,N_14926,N_13277);
or U17384 (N_17384,N_13921,N_12853);
xnor U17385 (N_17385,N_13757,N_12773);
nand U17386 (N_17386,N_14740,N_14187);
nand U17387 (N_17387,N_14249,N_13986);
and U17388 (N_17388,N_12700,N_12970);
xor U17389 (N_17389,N_12115,N_13490);
xor U17390 (N_17390,N_12802,N_14470);
nand U17391 (N_17391,N_13409,N_13599);
xor U17392 (N_17392,N_14706,N_12391);
nor U17393 (N_17393,N_14103,N_14017);
nor U17394 (N_17394,N_14939,N_12264);
nand U17395 (N_17395,N_14828,N_12468);
xnor U17396 (N_17396,N_12484,N_13750);
and U17397 (N_17397,N_12793,N_12380);
nor U17398 (N_17398,N_14791,N_14428);
or U17399 (N_17399,N_12628,N_12876);
nor U17400 (N_17400,N_14749,N_12524);
nand U17401 (N_17401,N_14784,N_14078);
nor U17402 (N_17402,N_14658,N_14881);
nand U17403 (N_17403,N_14471,N_14346);
and U17404 (N_17404,N_12841,N_12574);
nor U17405 (N_17405,N_13243,N_12096);
or U17406 (N_17406,N_13403,N_14562);
nor U17407 (N_17407,N_13759,N_13693);
xor U17408 (N_17408,N_12749,N_12414);
or U17409 (N_17409,N_12131,N_14501);
xnor U17410 (N_17410,N_12704,N_14770);
xor U17411 (N_17411,N_13702,N_14755);
xnor U17412 (N_17412,N_14034,N_12154);
xor U17413 (N_17413,N_13626,N_12720);
and U17414 (N_17414,N_13204,N_13173);
and U17415 (N_17415,N_12151,N_14255);
xor U17416 (N_17416,N_13823,N_14550);
or U17417 (N_17417,N_14084,N_12360);
nor U17418 (N_17418,N_12780,N_14719);
nand U17419 (N_17419,N_14237,N_14489);
and U17420 (N_17420,N_14440,N_14084);
and U17421 (N_17421,N_13425,N_12642);
or U17422 (N_17422,N_12403,N_14044);
nor U17423 (N_17423,N_14857,N_13523);
or U17424 (N_17424,N_14196,N_14486);
xor U17425 (N_17425,N_14212,N_13860);
xor U17426 (N_17426,N_12417,N_12153);
and U17427 (N_17427,N_12594,N_14665);
nand U17428 (N_17428,N_13835,N_13291);
nand U17429 (N_17429,N_14744,N_13179);
nand U17430 (N_17430,N_14844,N_14272);
xnor U17431 (N_17431,N_14203,N_12148);
or U17432 (N_17432,N_12620,N_14571);
nand U17433 (N_17433,N_14222,N_12105);
and U17434 (N_17434,N_14143,N_13030);
xor U17435 (N_17435,N_12547,N_14278);
nand U17436 (N_17436,N_13011,N_14016);
xor U17437 (N_17437,N_14467,N_12467);
and U17438 (N_17438,N_14965,N_14523);
or U17439 (N_17439,N_12840,N_13886);
nand U17440 (N_17440,N_12978,N_13718);
or U17441 (N_17441,N_12619,N_14738);
or U17442 (N_17442,N_12597,N_12208);
xor U17443 (N_17443,N_14265,N_13331);
or U17444 (N_17444,N_13976,N_12955);
or U17445 (N_17445,N_14154,N_12321);
or U17446 (N_17446,N_14033,N_14311);
xnor U17447 (N_17447,N_13417,N_13547);
xor U17448 (N_17448,N_14545,N_14990);
xnor U17449 (N_17449,N_12344,N_13024);
xnor U17450 (N_17450,N_14228,N_12307);
nand U17451 (N_17451,N_12536,N_12909);
or U17452 (N_17452,N_14631,N_12091);
nand U17453 (N_17453,N_14256,N_12455);
and U17454 (N_17454,N_14936,N_13541);
or U17455 (N_17455,N_13562,N_13638);
xor U17456 (N_17456,N_14285,N_13461);
or U17457 (N_17457,N_14149,N_12494);
nor U17458 (N_17458,N_14207,N_14222);
nand U17459 (N_17459,N_12968,N_14099);
nor U17460 (N_17460,N_14997,N_13753);
xor U17461 (N_17461,N_14685,N_14666);
xnor U17462 (N_17462,N_12319,N_13064);
xor U17463 (N_17463,N_13622,N_13535);
and U17464 (N_17464,N_12087,N_12184);
and U17465 (N_17465,N_12579,N_12922);
and U17466 (N_17466,N_14045,N_13121);
and U17467 (N_17467,N_12214,N_13704);
nor U17468 (N_17468,N_13151,N_12151);
nor U17469 (N_17469,N_12392,N_12409);
and U17470 (N_17470,N_12209,N_13091);
xor U17471 (N_17471,N_13771,N_14943);
nand U17472 (N_17472,N_13002,N_12580);
and U17473 (N_17473,N_12079,N_12304);
or U17474 (N_17474,N_14731,N_14655);
xor U17475 (N_17475,N_12210,N_14007);
or U17476 (N_17476,N_14864,N_14376);
nand U17477 (N_17477,N_12691,N_12084);
or U17478 (N_17478,N_14382,N_12030);
nor U17479 (N_17479,N_13910,N_14840);
xor U17480 (N_17480,N_12420,N_12594);
and U17481 (N_17481,N_14672,N_13619);
and U17482 (N_17482,N_14529,N_13966);
nand U17483 (N_17483,N_14438,N_12680);
nor U17484 (N_17484,N_13286,N_13772);
nand U17485 (N_17485,N_13647,N_12721);
and U17486 (N_17486,N_12096,N_14551);
xnor U17487 (N_17487,N_12165,N_14825);
or U17488 (N_17488,N_13406,N_12132);
xor U17489 (N_17489,N_14076,N_13470);
nand U17490 (N_17490,N_13135,N_12229);
nand U17491 (N_17491,N_14338,N_12948);
and U17492 (N_17492,N_13703,N_14261);
nor U17493 (N_17493,N_12170,N_14653);
nor U17494 (N_17494,N_12368,N_14098);
nor U17495 (N_17495,N_13609,N_13810);
and U17496 (N_17496,N_13769,N_12525);
or U17497 (N_17497,N_14663,N_13874);
and U17498 (N_17498,N_14964,N_14828);
nor U17499 (N_17499,N_14150,N_12218);
nand U17500 (N_17500,N_14615,N_13168);
xnor U17501 (N_17501,N_14832,N_13527);
nor U17502 (N_17502,N_14666,N_13839);
and U17503 (N_17503,N_12265,N_14779);
and U17504 (N_17504,N_13322,N_13562);
or U17505 (N_17505,N_14440,N_13413);
nor U17506 (N_17506,N_13308,N_13174);
or U17507 (N_17507,N_14359,N_12386);
or U17508 (N_17508,N_13616,N_14036);
nor U17509 (N_17509,N_13576,N_14796);
xor U17510 (N_17510,N_14645,N_14906);
and U17511 (N_17511,N_13014,N_14792);
and U17512 (N_17512,N_12242,N_14051);
xnor U17513 (N_17513,N_14686,N_13068);
xnor U17514 (N_17514,N_12750,N_13344);
and U17515 (N_17515,N_13647,N_13252);
xor U17516 (N_17516,N_13991,N_12198);
xor U17517 (N_17517,N_14897,N_13841);
and U17518 (N_17518,N_14120,N_12921);
nor U17519 (N_17519,N_12749,N_14235);
or U17520 (N_17520,N_12473,N_14592);
nor U17521 (N_17521,N_14714,N_13888);
nand U17522 (N_17522,N_13746,N_12271);
nand U17523 (N_17523,N_12008,N_14225);
and U17524 (N_17524,N_12678,N_12072);
and U17525 (N_17525,N_12015,N_12180);
xnor U17526 (N_17526,N_14883,N_13405);
nand U17527 (N_17527,N_13848,N_14897);
and U17528 (N_17528,N_12035,N_13910);
xor U17529 (N_17529,N_13989,N_14832);
nor U17530 (N_17530,N_12963,N_13578);
nor U17531 (N_17531,N_13790,N_12708);
nor U17532 (N_17532,N_12992,N_14312);
or U17533 (N_17533,N_12727,N_14905);
xor U17534 (N_17534,N_12008,N_12558);
and U17535 (N_17535,N_12859,N_12263);
and U17536 (N_17536,N_13682,N_12122);
xor U17537 (N_17537,N_12968,N_12606);
nor U17538 (N_17538,N_12923,N_14813);
or U17539 (N_17539,N_14818,N_12996);
and U17540 (N_17540,N_12570,N_13588);
nor U17541 (N_17541,N_12409,N_14350);
or U17542 (N_17542,N_14351,N_13650);
and U17543 (N_17543,N_12416,N_12606);
nand U17544 (N_17544,N_14338,N_13560);
nand U17545 (N_17545,N_12190,N_12040);
xnor U17546 (N_17546,N_14039,N_12879);
xor U17547 (N_17547,N_12266,N_12499);
xor U17548 (N_17548,N_14339,N_13157);
or U17549 (N_17549,N_13050,N_12046);
nor U17550 (N_17550,N_12994,N_12717);
or U17551 (N_17551,N_13505,N_14636);
or U17552 (N_17552,N_13601,N_13886);
xor U17553 (N_17553,N_13587,N_12796);
nor U17554 (N_17554,N_12054,N_12676);
or U17555 (N_17555,N_14863,N_13697);
nor U17556 (N_17556,N_12621,N_12446);
nand U17557 (N_17557,N_12152,N_12285);
and U17558 (N_17558,N_14481,N_12616);
nor U17559 (N_17559,N_13581,N_12930);
and U17560 (N_17560,N_12535,N_13287);
nand U17561 (N_17561,N_13689,N_14761);
nand U17562 (N_17562,N_12826,N_13560);
and U17563 (N_17563,N_12924,N_14798);
and U17564 (N_17564,N_13282,N_13324);
and U17565 (N_17565,N_12631,N_12624);
xor U17566 (N_17566,N_14680,N_14492);
nor U17567 (N_17567,N_13223,N_14550);
xnor U17568 (N_17568,N_12923,N_13492);
or U17569 (N_17569,N_14297,N_14254);
xnor U17570 (N_17570,N_13580,N_14329);
or U17571 (N_17571,N_12400,N_12097);
or U17572 (N_17572,N_13942,N_14686);
xnor U17573 (N_17573,N_14520,N_14531);
nand U17574 (N_17574,N_13510,N_12156);
nand U17575 (N_17575,N_12047,N_12458);
nor U17576 (N_17576,N_14730,N_13178);
or U17577 (N_17577,N_13940,N_13272);
and U17578 (N_17578,N_12691,N_12765);
and U17579 (N_17579,N_12124,N_13702);
and U17580 (N_17580,N_12891,N_13469);
xnor U17581 (N_17581,N_14859,N_14721);
or U17582 (N_17582,N_14486,N_13395);
nor U17583 (N_17583,N_12070,N_12868);
and U17584 (N_17584,N_12736,N_14933);
xnor U17585 (N_17585,N_13520,N_14611);
and U17586 (N_17586,N_12904,N_14324);
or U17587 (N_17587,N_12112,N_13519);
nand U17588 (N_17588,N_14007,N_13778);
xor U17589 (N_17589,N_14863,N_14525);
or U17590 (N_17590,N_12842,N_14481);
nand U17591 (N_17591,N_12323,N_14862);
or U17592 (N_17592,N_12496,N_13718);
or U17593 (N_17593,N_12173,N_14783);
nand U17594 (N_17594,N_13453,N_13216);
nor U17595 (N_17595,N_12450,N_12583);
and U17596 (N_17596,N_13338,N_14211);
nand U17597 (N_17597,N_13844,N_13564);
nor U17598 (N_17598,N_13062,N_12787);
and U17599 (N_17599,N_12896,N_14993);
nand U17600 (N_17600,N_12370,N_13310);
nor U17601 (N_17601,N_12088,N_14204);
nand U17602 (N_17602,N_14870,N_14048);
nor U17603 (N_17603,N_13608,N_14117);
xor U17604 (N_17604,N_13076,N_13190);
and U17605 (N_17605,N_12145,N_12109);
or U17606 (N_17606,N_14824,N_14337);
nor U17607 (N_17607,N_13820,N_12920);
or U17608 (N_17608,N_12036,N_13498);
nor U17609 (N_17609,N_13182,N_12930);
or U17610 (N_17610,N_12536,N_14199);
nor U17611 (N_17611,N_14252,N_14384);
and U17612 (N_17612,N_12025,N_13161);
and U17613 (N_17613,N_12532,N_13171);
or U17614 (N_17614,N_13732,N_12342);
or U17615 (N_17615,N_13346,N_12599);
or U17616 (N_17616,N_13850,N_14674);
or U17617 (N_17617,N_13681,N_14651);
or U17618 (N_17618,N_12103,N_14591);
nand U17619 (N_17619,N_14180,N_14970);
nor U17620 (N_17620,N_13455,N_12142);
nor U17621 (N_17621,N_13270,N_12722);
xor U17622 (N_17622,N_12079,N_12873);
nor U17623 (N_17623,N_13627,N_12699);
xnor U17624 (N_17624,N_13989,N_12831);
xor U17625 (N_17625,N_13453,N_13691);
and U17626 (N_17626,N_14222,N_14997);
xnor U17627 (N_17627,N_13499,N_13346);
and U17628 (N_17628,N_13368,N_12866);
nand U17629 (N_17629,N_12997,N_13376);
and U17630 (N_17630,N_14289,N_13813);
nand U17631 (N_17631,N_12190,N_13954);
nand U17632 (N_17632,N_14306,N_13381);
xor U17633 (N_17633,N_13955,N_14273);
nand U17634 (N_17634,N_12168,N_12544);
or U17635 (N_17635,N_13153,N_14156);
xnor U17636 (N_17636,N_13486,N_14379);
nand U17637 (N_17637,N_14209,N_13029);
and U17638 (N_17638,N_14851,N_13544);
or U17639 (N_17639,N_14097,N_14785);
and U17640 (N_17640,N_12754,N_12896);
xor U17641 (N_17641,N_14872,N_13342);
or U17642 (N_17642,N_12311,N_12528);
and U17643 (N_17643,N_12798,N_13354);
or U17644 (N_17644,N_12879,N_12562);
nand U17645 (N_17645,N_12017,N_13116);
xnor U17646 (N_17646,N_12230,N_12466);
and U17647 (N_17647,N_14322,N_12524);
and U17648 (N_17648,N_12690,N_13706);
nor U17649 (N_17649,N_12934,N_12953);
xor U17650 (N_17650,N_14259,N_13198);
xnor U17651 (N_17651,N_14474,N_13686);
nor U17652 (N_17652,N_14935,N_14744);
nand U17653 (N_17653,N_12213,N_13992);
nand U17654 (N_17654,N_14695,N_14335);
xnor U17655 (N_17655,N_14511,N_12968);
and U17656 (N_17656,N_12343,N_12543);
nand U17657 (N_17657,N_14890,N_13808);
nand U17658 (N_17658,N_13083,N_14790);
or U17659 (N_17659,N_14364,N_13780);
xnor U17660 (N_17660,N_12093,N_13238);
nand U17661 (N_17661,N_13156,N_14564);
nand U17662 (N_17662,N_13444,N_12089);
and U17663 (N_17663,N_13489,N_14562);
xnor U17664 (N_17664,N_13366,N_14452);
nor U17665 (N_17665,N_14762,N_13558);
nand U17666 (N_17666,N_13829,N_13109);
nor U17667 (N_17667,N_12929,N_13920);
nand U17668 (N_17668,N_12705,N_14001);
and U17669 (N_17669,N_12351,N_13643);
xor U17670 (N_17670,N_14038,N_13637);
xor U17671 (N_17671,N_13370,N_12378);
xnor U17672 (N_17672,N_14876,N_12885);
and U17673 (N_17673,N_12761,N_12339);
and U17674 (N_17674,N_12199,N_13476);
nor U17675 (N_17675,N_14794,N_14465);
xnor U17676 (N_17676,N_12299,N_13140);
nor U17677 (N_17677,N_14690,N_13275);
or U17678 (N_17678,N_12971,N_12949);
or U17679 (N_17679,N_13593,N_14470);
nor U17680 (N_17680,N_14038,N_14108);
nor U17681 (N_17681,N_12499,N_14991);
or U17682 (N_17682,N_14500,N_12215);
nor U17683 (N_17683,N_13186,N_13738);
nand U17684 (N_17684,N_13480,N_13045);
xnor U17685 (N_17685,N_14533,N_13314);
nand U17686 (N_17686,N_14806,N_14275);
and U17687 (N_17687,N_14432,N_12943);
nor U17688 (N_17688,N_13433,N_13636);
nand U17689 (N_17689,N_12208,N_12859);
and U17690 (N_17690,N_14177,N_13705);
xnor U17691 (N_17691,N_14692,N_13759);
or U17692 (N_17692,N_14821,N_13728);
xor U17693 (N_17693,N_13403,N_14730);
and U17694 (N_17694,N_14952,N_13628);
nand U17695 (N_17695,N_12797,N_13251);
nor U17696 (N_17696,N_12110,N_13202);
and U17697 (N_17697,N_14725,N_14420);
xor U17698 (N_17698,N_14477,N_14999);
or U17699 (N_17699,N_12668,N_14331);
nand U17700 (N_17700,N_14266,N_12480);
and U17701 (N_17701,N_14338,N_12332);
xnor U17702 (N_17702,N_13990,N_14609);
nor U17703 (N_17703,N_14818,N_12781);
and U17704 (N_17704,N_12129,N_12722);
and U17705 (N_17705,N_13543,N_14701);
and U17706 (N_17706,N_12659,N_12415);
and U17707 (N_17707,N_14172,N_13964);
and U17708 (N_17708,N_12432,N_12313);
and U17709 (N_17709,N_14526,N_14595);
and U17710 (N_17710,N_13013,N_13055);
or U17711 (N_17711,N_12424,N_12674);
or U17712 (N_17712,N_14150,N_13383);
and U17713 (N_17713,N_14570,N_13816);
xnor U17714 (N_17714,N_13479,N_13075);
nand U17715 (N_17715,N_12939,N_12093);
and U17716 (N_17716,N_14997,N_13824);
and U17717 (N_17717,N_13614,N_14302);
nor U17718 (N_17718,N_13082,N_12985);
or U17719 (N_17719,N_14097,N_12076);
nor U17720 (N_17720,N_12882,N_12427);
xnor U17721 (N_17721,N_13846,N_14166);
nor U17722 (N_17722,N_12030,N_13170);
nor U17723 (N_17723,N_12416,N_13512);
or U17724 (N_17724,N_12246,N_14538);
xnor U17725 (N_17725,N_14673,N_14941);
nand U17726 (N_17726,N_13465,N_14451);
nor U17727 (N_17727,N_14349,N_12621);
nand U17728 (N_17728,N_12967,N_13115);
nor U17729 (N_17729,N_14017,N_14213);
nand U17730 (N_17730,N_12212,N_14632);
or U17731 (N_17731,N_13984,N_13352);
nor U17732 (N_17732,N_14600,N_13137);
xnor U17733 (N_17733,N_13846,N_12727);
or U17734 (N_17734,N_13681,N_12713);
and U17735 (N_17735,N_13691,N_14031);
nor U17736 (N_17736,N_13345,N_12818);
xor U17737 (N_17737,N_12492,N_14577);
or U17738 (N_17738,N_14288,N_14485);
and U17739 (N_17739,N_12171,N_12503);
nand U17740 (N_17740,N_12877,N_13601);
nor U17741 (N_17741,N_13525,N_13603);
and U17742 (N_17742,N_13239,N_14046);
and U17743 (N_17743,N_13359,N_13923);
nand U17744 (N_17744,N_13890,N_13279);
xnor U17745 (N_17745,N_12178,N_13433);
nand U17746 (N_17746,N_13403,N_13110);
or U17747 (N_17747,N_14717,N_12520);
nand U17748 (N_17748,N_14582,N_12328);
and U17749 (N_17749,N_14649,N_13941);
and U17750 (N_17750,N_13133,N_12570);
nor U17751 (N_17751,N_13477,N_13706);
xor U17752 (N_17752,N_13597,N_14606);
and U17753 (N_17753,N_13578,N_13523);
and U17754 (N_17754,N_13451,N_13052);
nor U17755 (N_17755,N_13122,N_12926);
or U17756 (N_17756,N_13837,N_13609);
or U17757 (N_17757,N_14910,N_13702);
or U17758 (N_17758,N_14031,N_13233);
and U17759 (N_17759,N_12753,N_12062);
nand U17760 (N_17760,N_12527,N_13443);
xor U17761 (N_17761,N_13588,N_14624);
or U17762 (N_17762,N_13493,N_14708);
nor U17763 (N_17763,N_13093,N_13835);
and U17764 (N_17764,N_13723,N_13312);
nor U17765 (N_17765,N_12105,N_14111);
nor U17766 (N_17766,N_14914,N_13696);
or U17767 (N_17767,N_13687,N_12397);
and U17768 (N_17768,N_12596,N_14305);
and U17769 (N_17769,N_14253,N_12803);
nor U17770 (N_17770,N_12815,N_12898);
nor U17771 (N_17771,N_14440,N_14516);
nor U17772 (N_17772,N_12390,N_13107);
or U17773 (N_17773,N_14982,N_14003);
nor U17774 (N_17774,N_12527,N_12044);
nor U17775 (N_17775,N_12316,N_12723);
nor U17776 (N_17776,N_12300,N_14889);
or U17777 (N_17777,N_14737,N_13402);
nand U17778 (N_17778,N_12810,N_14844);
nand U17779 (N_17779,N_12553,N_12359);
xor U17780 (N_17780,N_13435,N_12249);
and U17781 (N_17781,N_13632,N_14992);
and U17782 (N_17782,N_14157,N_12768);
nor U17783 (N_17783,N_14991,N_12071);
nor U17784 (N_17784,N_12440,N_14173);
and U17785 (N_17785,N_14996,N_14008);
nand U17786 (N_17786,N_13943,N_12474);
nor U17787 (N_17787,N_12448,N_12497);
and U17788 (N_17788,N_14605,N_14188);
nand U17789 (N_17789,N_13366,N_13149);
or U17790 (N_17790,N_14501,N_12348);
xnor U17791 (N_17791,N_14828,N_14622);
or U17792 (N_17792,N_13158,N_14476);
xnor U17793 (N_17793,N_13294,N_12836);
or U17794 (N_17794,N_12962,N_13846);
nor U17795 (N_17795,N_14673,N_13334);
or U17796 (N_17796,N_13778,N_13686);
and U17797 (N_17797,N_13627,N_13509);
nor U17798 (N_17798,N_13350,N_13654);
nand U17799 (N_17799,N_13375,N_13027);
and U17800 (N_17800,N_12405,N_12420);
nand U17801 (N_17801,N_14872,N_14624);
and U17802 (N_17802,N_12904,N_13919);
and U17803 (N_17803,N_14711,N_12364);
or U17804 (N_17804,N_13650,N_14147);
nand U17805 (N_17805,N_13571,N_12545);
nor U17806 (N_17806,N_13302,N_12007);
xor U17807 (N_17807,N_14959,N_13432);
xnor U17808 (N_17808,N_14158,N_13934);
nor U17809 (N_17809,N_14000,N_12568);
or U17810 (N_17810,N_14085,N_12554);
nand U17811 (N_17811,N_13838,N_12721);
or U17812 (N_17812,N_12580,N_13292);
or U17813 (N_17813,N_12740,N_14646);
and U17814 (N_17814,N_13277,N_12947);
or U17815 (N_17815,N_12863,N_13793);
xnor U17816 (N_17816,N_13419,N_13228);
xor U17817 (N_17817,N_12169,N_14737);
and U17818 (N_17818,N_14323,N_13275);
and U17819 (N_17819,N_14500,N_14747);
and U17820 (N_17820,N_13654,N_13596);
xor U17821 (N_17821,N_12065,N_12441);
and U17822 (N_17822,N_12432,N_14527);
nand U17823 (N_17823,N_12122,N_13457);
or U17824 (N_17824,N_12079,N_14038);
nand U17825 (N_17825,N_13075,N_14419);
and U17826 (N_17826,N_14080,N_12301);
nand U17827 (N_17827,N_12894,N_13155);
nor U17828 (N_17828,N_13158,N_14637);
nor U17829 (N_17829,N_14039,N_14264);
xnor U17830 (N_17830,N_13392,N_13731);
or U17831 (N_17831,N_14504,N_14123);
xor U17832 (N_17832,N_14603,N_14381);
or U17833 (N_17833,N_12010,N_12345);
nor U17834 (N_17834,N_12137,N_12539);
nor U17835 (N_17835,N_13550,N_12122);
or U17836 (N_17836,N_12450,N_14330);
nor U17837 (N_17837,N_13438,N_12150);
and U17838 (N_17838,N_13975,N_12127);
nor U17839 (N_17839,N_14753,N_12952);
and U17840 (N_17840,N_14502,N_14177);
xnor U17841 (N_17841,N_14161,N_12724);
and U17842 (N_17842,N_13629,N_14949);
xor U17843 (N_17843,N_14773,N_14768);
nand U17844 (N_17844,N_13174,N_13423);
nor U17845 (N_17845,N_14904,N_13308);
and U17846 (N_17846,N_12538,N_12249);
xnor U17847 (N_17847,N_12103,N_13047);
and U17848 (N_17848,N_14669,N_12494);
nand U17849 (N_17849,N_14286,N_12999);
and U17850 (N_17850,N_14144,N_13330);
nor U17851 (N_17851,N_13926,N_12379);
nand U17852 (N_17852,N_14839,N_12265);
and U17853 (N_17853,N_14246,N_14841);
nand U17854 (N_17854,N_14733,N_13995);
nand U17855 (N_17855,N_13726,N_12013);
nor U17856 (N_17856,N_13792,N_12410);
xor U17857 (N_17857,N_14009,N_13864);
or U17858 (N_17858,N_13946,N_14564);
and U17859 (N_17859,N_12631,N_12138);
xor U17860 (N_17860,N_12750,N_12204);
xnor U17861 (N_17861,N_12824,N_12652);
and U17862 (N_17862,N_14191,N_12200);
and U17863 (N_17863,N_12536,N_13628);
nor U17864 (N_17864,N_13516,N_12795);
nor U17865 (N_17865,N_12068,N_13025);
xnor U17866 (N_17866,N_14047,N_14086);
nor U17867 (N_17867,N_13166,N_14223);
nor U17868 (N_17868,N_13911,N_14656);
and U17869 (N_17869,N_13420,N_12120);
nor U17870 (N_17870,N_14909,N_14145);
or U17871 (N_17871,N_13995,N_14198);
and U17872 (N_17872,N_13091,N_12753);
and U17873 (N_17873,N_13560,N_12303);
or U17874 (N_17874,N_14084,N_12065);
xor U17875 (N_17875,N_13905,N_12150);
nor U17876 (N_17876,N_13187,N_13741);
nor U17877 (N_17877,N_12035,N_12965);
xor U17878 (N_17878,N_14981,N_13132);
xnor U17879 (N_17879,N_12389,N_14830);
nand U17880 (N_17880,N_14652,N_14746);
xor U17881 (N_17881,N_12232,N_14711);
nor U17882 (N_17882,N_12057,N_12901);
and U17883 (N_17883,N_13780,N_13406);
xor U17884 (N_17884,N_12305,N_14160);
nor U17885 (N_17885,N_14189,N_13774);
nor U17886 (N_17886,N_13522,N_12210);
nor U17887 (N_17887,N_14622,N_13047);
and U17888 (N_17888,N_14486,N_13133);
nand U17889 (N_17889,N_14400,N_14439);
nand U17890 (N_17890,N_13483,N_13361);
or U17891 (N_17891,N_14445,N_12185);
nor U17892 (N_17892,N_14522,N_13274);
xor U17893 (N_17893,N_14908,N_13116);
nand U17894 (N_17894,N_12891,N_12110);
or U17895 (N_17895,N_13894,N_13343);
and U17896 (N_17896,N_14164,N_14642);
nand U17897 (N_17897,N_13154,N_12770);
xnor U17898 (N_17898,N_13393,N_12648);
xor U17899 (N_17899,N_13645,N_13610);
or U17900 (N_17900,N_12657,N_13901);
or U17901 (N_17901,N_14762,N_13678);
xnor U17902 (N_17902,N_13251,N_14272);
nand U17903 (N_17903,N_13484,N_12091);
nor U17904 (N_17904,N_14783,N_13184);
and U17905 (N_17905,N_14436,N_12846);
nor U17906 (N_17906,N_12503,N_14508);
and U17907 (N_17907,N_13188,N_14072);
and U17908 (N_17908,N_13913,N_14944);
and U17909 (N_17909,N_13221,N_13052);
and U17910 (N_17910,N_14507,N_13874);
nor U17911 (N_17911,N_14480,N_12054);
nor U17912 (N_17912,N_14535,N_12908);
nor U17913 (N_17913,N_14717,N_14617);
and U17914 (N_17914,N_13098,N_12954);
nor U17915 (N_17915,N_12964,N_13329);
xor U17916 (N_17916,N_12650,N_12041);
xor U17917 (N_17917,N_13614,N_12677);
and U17918 (N_17918,N_13034,N_12553);
and U17919 (N_17919,N_12212,N_13405);
and U17920 (N_17920,N_13298,N_12360);
xor U17921 (N_17921,N_13667,N_14819);
or U17922 (N_17922,N_12185,N_14585);
and U17923 (N_17923,N_12942,N_12804);
xor U17924 (N_17924,N_13617,N_14299);
xnor U17925 (N_17925,N_14997,N_14862);
nand U17926 (N_17926,N_13711,N_13094);
xor U17927 (N_17927,N_13387,N_14199);
nor U17928 (N_17928,N_14540,N_14717);
nor U17929 (N_17929,N_14849,N_13549);
nor U17930 (N_17930,N_14859,N_13184);
nand U17931 (N_17931,N_13824,N_12182);
nand U17932 (N_17932,N_12086,N_14796);
and U17933 (N_17933,N_14940,N_12403);
nand U17934 (N_17934,N_13295,N_13235);
nand U17935 (N_17935,N_12418,N_12336);
nand U17936 (N_17936,N_12158,N_12614);
nor U17937 (N_17937,N_12253,N_12121);
xnor U17938 (N_17938,N_13629,N_14144);
nand U17939 (N_17939,N_12559,N_12510);
xnor U17940 (N_17940,N_14925,N_12378);
or U17941 (N_17941,N_13892,N_13718);
nand U17942 (N_17942,N_12770,N_14458);
xor U17943 (N_17943,N_14215,N_13511);
nor U17944 (N_17944,N_12829,N_13020);
nor U17945 (N_17945,N_13102,N_13884);
and U17946 (N_17946,N_13149,N_14129);
xor U17947 (N_17947,N_12296,N_12830);
or U17948 (N_17948,N_12596,N_14185);
and U17949 (N_17949,N_13411,N_14611);
or U17950 (N_17950,N_13250,N_13107);
and U17951 (N_17951,N_14638,N_12761);
and U17952 (N_17952,N_12589,N_14850);
and U17953 (N_17953,N_12587,N_12144);
nor U17954 (N_17954,N_12079,N_12158);
or U17955 (N_17955,N_14581,N_13969);
xnor U17956 (N_17956,N_13163,N_14056);
xor U17957 (N_17957,N_14825,N_12114);
nand U17958 (N_17958,N_12173,N_13944);
xnor U17959 (N_17959,N_13526,N_13172);
nor U17960 (N_17960,N_12670,N_13176);
nor U17961 (N_17961,N_12683,N_13752);
xnor U17962 (N_17962,N_14684,N_12962);
xor U17963 (N_17963,N_12242,N_13113);
or U17964 (N_17964,N_13639,N_13807);
nand U17965 (N_17965,N_12108,N_14938);
nand U17966 (N_17966,N_12631,N_12232);
nand U17967 (N_17967,N_13025,N_12291);
nor U17968 (N_17968,N_12183,N_13878);
xor U17969 (N_17969,N_14267,N_13205);
and U17970 (N_17970,N_13453,N_14412);
nand U17971 (N_17971,N_13982,N_13250);
and U17972 (N_17972,N_13708,N_14603);
xnor U17973 (N_17973,N_14237,N_12892);
nor U17974 (N_17974,N_14022,N_13339);
and U17975 (N_17975,N_13135,N_12234);
nor U17976 (N_17976,N_13670,N_13074);
xor U17977 (N_17977,N_13656,N_14743);
nand U17978 (N_17978,N_14986,N_14229);
or U17979 (N_17979,N_13342,N_14079);
and U17980 (N_17980,N_13609,N_13576);
xnor U17981 (N_17981,N_14082,N_13079);
nand U17982 (N_17982,N_13036,N_14876);
nand U17983 (N_17983,N_13488,N_12119);
or U17984 (N_17984,N_14155,N_12093);
and U17985 (N_17985,N_14467,N_13021);
nor U17986 (N_17986,N_12178,N_12560);
nand U17987 (N_17987,N_13006,N_13974);
and U17988 (N_17988,N_12985,N_12570);
nor U17989 (N_17989,N_13387,N_12216);
nor U17990 (N_17990,N_12375,N_12046);
or U17991 (N_17991,N_14626,N_12180);
xor U17992 (N_17992,N_14504,N_12563);
and U17993 (N_17993,N_13712,N_12261);
xor U17994 (N_17994,N_12153,N_13860);
or U17995 (N_17995,N_12399,N_13323);
xor U17996 (N_17996,N_14090,N_14240);
and U17997 (N_17997,N_14213,N_12648);
nor U17998 (N_17998,N_13753,N_13524);
xor U17999 (N_17999,N_14294,N_13730);
nand U18000 (N_18000,N_17843,N_17682);
nor U18001 (N_18001,N_15127,N_16496);
nor U18002 (N_18002,N_16242,N_15161);
or U18003 (N_18003,N_17239,N_17007);
nor U18004 (N_18004,N_17791,N_17549);
xnor U18005 (N_18005,N_16798,N_17245);
xor U18006 (N_18006,N_17509,N_17743);
nor U18007 (N_18007,N_15007,N_16054);
xor U18008 (N_18008,N_15016,N_17209);
or U18009 (N_18009,N_17412,N_17808);
and U18010 (N_18010,N_17069,N_17680);
xor U18011 (N_18011,N_17347,N_16746);
nand U18012 (N_18012,N_17656,N_17301);
and U18013 (N_18013,N_17231,N_16953);
and U18014 (N_18014,N_17519,N_16246);
or U18015 (N_18015,N_16661,N_15238);
and U18016 (N_18016,N_17583,N_17824);
and U18017 (N_18017,N_16811,N_16702);
nor U18018 (N_18018,N_15629,N_17480);
or U18019 (N_18019,N_17880,N_16861);
or U18020 (N_18020,N_17015,N_16845);
nor U18021 (N_18021,N_17688,N_15447);
nor U18022 (N_18022,N_17841,N_17102);
nand U18023 (N_18023,N_15578,N_15549);
and U18024 (N_18024,N_16468,N_15683);
or U18025 (N_18025,N_16976,N_17278);
or U18026 (N_18026,N_15569,N_15178);
and U18027 (N_18027,N_16170,N_15732);
and U18028 (N_18028,N_17956,N_16166);
nor U18029 (N_18029,N_16247,N_15965);
xnor U18030 (N_18030,N_15148,N_16268);
and U18031 (N_18031,N_15292,N_15940);
or U18032 (N_18032,N_16175,N_17960);
and U18033 (N_18033,N_15232,N_17426);
nand U18034 (N_18034,N_15956,N_17834);
and U18035 (N_18035,N_15710,N_15809);
nor U18036 (N_18036,N_17451,N_17391);
nor U18037 (N_18037,N_17847,N_15457);
and U18038 (N_18038,N_16136,N_16872);
xor U18039 (N_18039,N_15900,N_16086);
and U18040 (N_18040,N_17001,N_17285);
or U18041 (N_18041,N_16668,N_15189);
xor U18042 (N_18042,N_16141,N_16847);
nand U18043 (N_18043,N_17244,N_15833);
and U18044 (N_18044,N_15023,N_17121);
or U18045 (N_18045,N_17675,N_15327);
nor U18046 (N_18046,N_16912,N_15626);
or U18047 (N_18047,N_16534,N_17101);
nand U18048 (N_18048,N_17579,N_17143);
or U18049 (N_18049,N_17421,N_15707);
and U18050 (N_18050,N_15342,N_15039);
nand U18051 (N_18051,N_17779,N_15307);
and U18052 (N_18052,N_16821,N_15879);
and U18053 (N_18053,N_16714,N_15403);
nor U18054 (N_18054,N_15181,N_15970);
nor U18055 (N_18055,N_16184,N_15767);
or U18056 (N_18056,N_16424,N_16177);
nor U18057 (N_18057,N_15377,N_16435);
and U18058 (N_18058,N_15860,N_16838);
and U18059 (N_18059,N_17352,N_16551);
and U18060 (N_18060,N_16905,N_17505);
nor U18061 (N_18061,N_15923,N_17157);
xnor U18062 (N_18062,N_15436,N_17870);
nor U18063 (N_18063,N_16282,N_17689);
or U18064 (N_18064,N_16783,N_16236);
nand U18065 (N_18065,N_17514,N_16999);
and U18066 (N_18066,N_16816,N_16671);
nand U18067 (N_18067,N_17765,N_16635);
xnor U18068 (N_18068,N_15702,N_15701);
xor U18069 (N_18069,N_15361,N_15777);
or U18070 (N_18070,N_16874,N_17544);
or U18071 (N_18071,N_16589,N_17623);
nor U18072 (N_18072,N_16127,N_15577);
nor U18073 (N_18073,N_17810,N_15160);
nand U18074 (N_18074,N_16176,N_15362);
xor U18075 (N_18075,N_17695,N_16367);
xor U18076 (N_18076,N_16214,N_15163);
nand U18077 (N_18077,N_17324,N_16998);
nand U18078 (N_18078,N_16139,N_17433);
xor U18079 (N_18079,N_17194,N_17261);
and U18080 (N_18080,N_15453,N_15284);
nor U18081 (N_18081,N_15653,N_16760);
and U18082 (N_18082,N_16725,N_15691);
xnor U18083 (N_18083,N_17279,N_17502);
xor U18084 (N_18084,N_17089,N_16736);
nand U18085 (N_18085,N_16737,N_17162);
nand U18086 (N_18086,N_17876,N_16590);
nand U18087 (N_18087,N_17465,N_17388);
and U18088 (N_18088,N_16074,N_16051);
nand U18089 (N_18089,N_17540,N_16539);
and U18090 (N_18090,N_16995,N_15205);
and U18091 (N_18091,N_16672,N_17972);
and U18092 (N_18092,N_17443,N_16449);
nor U18093 (N_18093,N_15846,N_16209);
xor U18094 (N_18094,N_15088,N_17446);
xor U18095 (N_18095,N_15842,N_17319);
and U18096 (N_18096,N_15925,N_15158);
or U18097 (N_18097,N_16562,N_16450);
nand U18098 (N_18098,N_15644,N_16690);
nand U18099 (N_18099,N_16526,N_16949);
xor U18100 (N_18100,N_17294,N_16126);
xnor U18101 (N_18101,N_15267,N_15674);
xnor U18102 (N_18102,N_16092,N_16490);
xnor U18103 (N_18103,N_16831,N_15726);
and U18104 (N_18104,N_16498,N_17633);
nand U18105 (N_18105,N_15346,N_16947);
nand U18106 (N_18106,N_17066,N_16875);
nand U18107 (N_18107,N_15311,N_17335);
and U18108 (N_18108,N_17235,N_15737);
and U18109 (N_18109,N_16160,N_16055);
and U18110 (N_18110,N_15031,N_15152);
and U18111 (N_18111,N_15109,N_16673);
or U18112 (N_18112,N_15926,N_16622);
and U18113 (N_18113,N_15456,N_16470);
and U18114 (N_18114,N_17067,N_17123);
or U18115 (N_18115,N_15547,N_16320);
nand U18116 (N_18116,N_16713,N_15613);
or U18117 (N_18117,N_16401,N_16115);
nand U18118 (N_18118,N_17306,N_15741);
nand U18119 (N_18119,N_16550,N_15123);
nand U18120 (N_18120,N_16730,N_15250);
xnor U18121 (N_18121,N_17440,N_15554);
nand U18122 (N_18122,N_17078,N_16586);
nand U18123 (N_18123,N_16790,N_16801);
nand U18124 (N_18124,N_15884,N_16917);
xor U18125 (N_18125,N_15545,N_16605);
and U18126 (N_18126,N_17223,N_16759);
and U18127 (N_18127,N_17251,N_16716);
nand U18128 (N_18128,N_15988,N_15459);
xnor U18129 (N_18129,N_15987,N_16818);
xor U18130 (N_18130,N_16323,N_16094);
nor U18131 (N_18131,N_15495,N_16570);
or U18132 (N_18132,N_15428,N_17707);
nand U18133 (N_18133,N_16738,N_15038);
nor U18134 (N_18134,N_17207,N_17813);
nand U18135 (N_18135,N_17287,N_16504);
nor U18136 (N_18136,N_15128,N_16846);
or U18137 (N_18137,N_16013,N_16777);
or U18138 (N_18138,N_15560,N_16147);
nand U18139 (N_18139,N_17558,N_16755);
nor U18140 (N_18140,N_15258,N_16198);
nand U18141 (N_18141,N_15841,N_15605);
xnor U18142 (N_18142,N_17337,N_17471);
xor U18143 (N_18143,N_17897,N_16399);
nor U18144 (N_18144,N_16497,N_15091);
nand U18145 (N_18145,N_17499,N_15948);
or U18146 (N_18146,N_17916,N_16856);
nor U18147 (N_18147,N_16105,N_17355);
nand U18148 (N_18148,N_15274,N_16767);
or U18149 (N_18149,N_17628,N_17243);
xor U18150 (N_18150,N_16945,N_17895);
or U18151 (N_18151,N_17706,N_17770);
or U18152 (N_18152,N_17037,N_17564);
xor U18153 (N_18153,N_17190,N_15045);
nand U18154 (N_18154,N_17871,N_15454);
xor U18155 (N_18155,N_16789,N_16220);
or U18156 (N_18156,N_16785,N_16321);
nor U18157 (N_18157,N_15015,N_16499);
nor U18158 (N_18158,N_17875,N_15681);
or U18159 (N_18159,N_17181,N_17635);
and U18160 (N_18160,N_16171,N_15348);
nand U18161 (N_18161,N_15591,N_17679);
or U18162 (N_18162,N_16108,N_16890);
nor U18163 (N_18163,N_16311,N_17602);
nor U18164 (N_18164,N_15551,N_15944);
xor U18165 (N_18165,N_15381,N_15680);
nand U18166 (N_18166,N_17864,N_16287);
nor U18167 (N_18167,N_17634,N_17299);
nand U18168 (N_18168,N_15721,N_17401);
xnor U18169 (N_18169,N_15515,N_17376);
or U18170 (N_18170,N_15920,N_15586);
nand U18171 (N_18171,N_16805,N_16229);
xnor U18172 (N_18172,N_17075,N_15073);
nand U18173 (N_18173,N_16135,N_16604);
nor U18174 (N_18174,N_17892,N_15355);
nor U18175 (N_18175,N_15142,N_16806);
nor U18176 (N_18176,N_15434,N_15749);
nand U18177 (N_18177,N_17988,N_17716);
xnor U18178 (N_18178,N_15787,N_15172);
or U18179 (N_18179,N_15937,N_17185);
xor U18180 (N_18180,N_17477,N_17009);
xor U18181 (N_18181,N_16536,N_15954);
and U18182 (N_18182,N_16207,N_17804);
nand U18183 (N_18183,N_16354,N_16727);
nor U18184 (N_18184,N_17850,N_15079);
or U18185 (N_18185,N_15801,N_17310);
and U18186 (N_18186,N_16081,N_16415);
and U18187 (N_18187,N_15761,N_16839);
and U18188 (N_18188,N_16355,N_16537);
nand U18189 (N_18189,N_17367,N_16840);
and U18190 (N_18190,N_17933,N_15933);
xnor U18191 (N_18191,N_16491,N_17043);
and U18192 (N_18192,N_15976,N_16775);
nand U18193 (N_18193,N_16882,N_16598);
nor U18194 (N_18194,N_17441,N_16578);
or U18195 (N_18195,N_15876,N_15055);
nand U18196 (N_18196,N_15449,N_17297);
and U18197 (N_18197,N_15938,N_17710);
or U18198 (N_18198,N_16483,N_17839);
nor U18199 (N_18199,N_17920,N_16603);
or U18200 (N_18200,N_15999,N_17565);
or U18201 (N_18201,N_17774,N_15217);
nor U18202 (N_18202,N_15173,N_17236);
or U18203 (N_18203,N_15193,N_17021);
or U18204 (N_18204,N_17270,N_15485);
or U18205 (N_18205,N_17837,N_16204);
and U18206 (N_18206,N_17885,N_17869);
or U18207 (N_18207,N_15351,N_15201);
xnor U18208 (N_18208,N_16380,N_17378);
nand U18209 (N_18209,N_15823,N_15229);
and U18210 (N_18210,N_17795,N_15411);
xnor U18211 (N_18211,N_17486,N_17184);
nand U18212 (N_18212,N_16773,N_15901);
xor U18213 (N_18213,N_15572,N_15345);
nand U18214 (N_18214,N_17842,N_16495);
nand U18215 (N_18215,N_15365,N_15089);
nor U18216 (N_18216,N_15743,N_17618);
or U18217 (N_18217,N_17913,N_16478);
xor U18218 (N_18218,N_17444,N_15593);
or U18219 (N_18219,N_15738,N_16476);
or U18220 (N_18220,N_16901,N_15730);
xnor U18221 (N_18221,N_15924,N_15783);
and U18222 (N_18222,N_16072,N_17690);
nand U18223 (N_18223,N_16117,N_17228);
nand U18224 (N_18224,N_16663,N_17148);
nand U18225 (N_18225,N_15100,N_15388);
xnor U18226 (N_18226,N_16111,N_15471);
nand U18227 (N_18227,N_16623,N_16288);
and U18228 (N_18228,N_17676,N_17823);
or U18229 (N_18229,N_15199,N_16233);
xor U18230 (N_18230,N_15343,N_16431);
xnor U18231 (N_18231,N_15029,N_17755);
nand U18232 (N_18232,N_16869,N_16196);
xor U18233 (N_18233,N_16008,N_16269);
nand U18234 (N_18234,N_16626,N_16968);
xnor U18235 (N_18235,N_15861,N_16064);
or U18236 (N_18236,N_16509,N_17780);
or U18237 (N_18237,N_15147,N_15636);
nor U18238 (N_18238,N_15950,N_17079);
and U18239 (N_18239,N_15305,N_17359);
and U18240 (N_18240,N_15996,N_15138);
nand U18241 (N_18241,N_15864,N_17063);
nor U18242 (N_18242,N_15918,N_15022);
xnor U18243 (N_18243,N_17491,N_15435);
xor U18244 (N_18244,N_16880,N_17608);
nor U18245 (N_18245,N_16909,N_16330);
and U18246 (N_18246,N_15005,N_16594);
nand U18247 (N_18247,N_17095,N_15106);
nand U18248 (N_18248,N_16150,N_16352);
xor U18249 (N_18249,N_16308,N_15755);
xnor U18250 (N_18250,N_16853,N_17398);
or U18251 (N_18251,N_17452,N_17149);
xnor U18252 (N_18252,N_17493,N_17516);
or U18253 (N_18253,N_16344,N_15706);
and U18254 (N_18254,N_17399,N_15501);
xnor U18255 (N_18255,N_17120,N_17183);
nor U18256 (N_18256,N_16152,N_17957);
and U18257 (N_18257,N_17986,N_17886);
and U18258 (N_18258,N_17664,N_17816);
nand U18259 (N_18259,N_16057,N_15117);
and U18260 (N_18260,N_15083,N_15579);
or U18261 (N_18261,N_15703,N_16595);
or U18262 (N_18262,N_17621,N_16296);
and U18263 (N_18263,N_15108,N_16651);
nor U18264 (N_18264,N_15081,N_15659);
xor U18265 (N_18265,N_16185,N_15899);
nand U18266 (N_18266,N_15746,N_15675);
xnor U18267 (N_18267,N_15122,N_16337);
and U18268 (N_18268,N_17025,N_16934);
nor U18269 (N_18269,N_16366,N_15019);
nor U18270 (N_18270,N_17993,N_16698);
xor U18271 (N_18271,N_15573,N_15678);
nand U18272 (N_18272,N_15625,N_15968);
xnor U18273 (N_18273,N_16422,N_15143);
nor U18274 (N_18274,N_16896,N_15672);
nand U18275 (N_18275,N_17304,N_16270);
xor U18276 (N_18276,N_17757,N_17980);
xor U18277 (N_18277,N_16278,N_17436);
and U18278 (N_18278,N_17476,N_15513);
and U18279 (N_18279,N_16987,N_17607);
and U18280 (N_18280,N_17174,N_16010);
or U18281 (N_18281,N_16700,N_17645);
nor U18282 (N_18282,N_15687,N_16900);
nor U18283 (N_18283,N_17172,N_16190);
or U18284 (N_18284,N_17482,N_16280);
nor U18285 (N_18285,N_16262,N_15025);
nand U18286 (N_18286,N_17784,N_17016);
nand U18287 (N_18287,N_15149,N_16692);
or U18288 (N_18288,N_15051,N_17703);
nor U18289 (N_18289,N_17935,N_16319);
or U18290 (N_18290,N_16217,N_17827);
xor U18291 (N_18291,N_16257,N_16427);
and U18292 (N_18292,N_15870,N_15409);
nor U18293 (N_18293,N_15308,N_17445);
xnor U18294 (N_18294,N_15306,N_16649);
nor U18295 (N_18295,N_17466,N_16647);
or U18296 (N_18296,N_15419,N_16819);
or U18297 (N_18297,N_15991,N_16492);
and U18298 (N_18298,N_15027,N_16002);
and U18299 (N_18299,N_16373,N_17830);
or U18300 (N_18300,N_15426,N_16774);
and U18301 (N_18301,N_17714,N_16012);
and U18302 (N_18302,N_16924,N_17365);
and U18303 (N_18303,N_17070,N_15961);
nor U18304 (N_18304,N_15341,N_17744);
and U18305 (N_18305,N_15734,N_16206);
and U18306 (N_18306,N_15408,N_15270);
nand U18307 (N_18307,N_15759,N_17825);
nor U18308 (N_18308,N_15074,N_16334);
xor U18309 (N_18309,N_15685,N_15442);
and U18310 (N_18310,N_15294,N_16708);
nor U18311 (N_18311,N_15155,N_15317);
and U18312 (N_18312,N_17967,N_16452);
nor U18313 (N_18313,N_16800,N_17595);
xor U18314 (N_18314,N_16787,N_16751);
nor U18315 (N_18315,N_17907,N_16519);
nor U18316 (N_18316,N_15104,N_16822);
nand U18317 (N_18317,N_15093,N_17400);
or U18318 (N_18318,N_15740,N_16275);
and U18319 (N_18319,N_15097,N_16593);
and U18320 (N_18320,N_15745,N_15883);
nor U18321 (N_18321,N_17150,N_15760);
nand U18322 (N_18322,N_16022,N_16103);
nor U18323 (N_18323,N_17735,N_16547);
and U18324 (N_18324,N_17991,N_17425);
or U18325 (N_18325,N_16471,N_15866);
or U18326 (N_18326,N_15309,N_16513);
nor U18327 (N_18327,N_17005,N_16560);
nor U18328 (N_18328,N_17921,N_17368);
nand U18329 (N_18329,N_15553,N_17230);
nor U18330 (N_18330,N_17545,N_15008);
nor U18331 (N_18331,N_15931,N_16408);
nand U18332 (N_18332,N_16089,N_16300);
nor U18333 (N_18333,N_15522,N_15224);
and U18334 (N_18334,N_17216,N_17622);
and U18335 (N_18335,N_15725,N_15978);
and U18336 (N_18336,N_17360,N_15048);
and U18337 (N_18337,N_15246,N_17073);
and U18338 (N_18338,N_15359,N_16637);
xnor U18339 (N_18339,N_16629,N_17662);
or U18340 (N_18340,N_16631,N_17132);
xnor U18341 (N_18341,N_17567,N_16091);
nor U18342 (N_18342,N_16503,N_15642);
or U18343 (N_18343,N_15479,N_15917);
or U18344 (N_18344,N_15095,N_17255);
xor U18345 (N_18345,N_16379,N_17926);
or U18346 (N_18346,N_17981,N_15855);
xnor U18347 (N_18347,N_17248,N_17587);
and U18348 (N_18348,N_15230,N_17220);
nand U18349 (N_18349,N_15692,N_16159);
xor U18350 (N_18350,N_15260,N_17857);
nand U18351 (N_18351,N_16075,N_17569);
and U18352 (N_18352,N_16895,N_16813);
nor U18353 (N_18353,N_17561,N_17550);
or U18354 (N_18354,N_16388,N_15332);
and U18355 (N_18355,N_15890,N_17867);
nand U18356 (N_18356,N_16535,N_17923);
xor U18357 (N_18357,N_15807,N_16019);
xnor U18358 (N_18358,N_17024,N_17585);
or U18359 (N_18359,N_16048,N_17568);
and U18360 (N_18360,N_16740,N_15592);
nand U18361 (N_18361,N_16243,N_17694);
and U18362 (N_18362,N_16829,N_15329);
nand U18363 (N_18363,N_16045,N_16733);
or U18364 (N_18364,N_16003,N_17848);
nand U18365 (N_18365,N_16414,N_15330);
xnor U18366 (N_18366,N_15829,N_16812);
and U18367 (N_18367,N_16963,N_16704);
xnor U18368 (N_18368,N_17211,N_17548);
nor U18369 (N_18369,N_17363,N_17574);
or U18370 (N_18370,N_17948,N_17702);
xor U18371 (N_18371,N_15429,N_15298);
or U18372 (N_18372,N_17592,N_16646);
nor U18373 (N_18373,N_15661,N_15788);
nand U18374 (N_18374,N_17214,N_16133);
nand U18375 (N_18375,N_15945,N_15257);
or U18376 (N_18376,N_16786,N_17670);
or U18377 (N_18377,N_16301,N_16416);
and U18378 (N_18378,N_17720,N_17543);
nand U18379 (N_18379,N_15384,N_16689);
nor U18380 (N_18380,N_17718,N_15655);
or U18381 (N_18381,N_17929,N_15324);
nand U18382 (N_18382,N_16753,N_15752);
nand U18383 (N_18383,N_17331,N_16557);
nand U18384 (N_18384,N_15877,N_17210);
xnor U18385 (N_18385,N_17658,N_16252);
or U18386 (N_18386,N_16883,N_16169);
xor U18387 (N_18387,N_16318,N_17512);
or U18388 (N_18388,N_17076,N_17275);
nor U18389 (N_18389,N_15443,N_15076);
or U18390 (N_18390,N_16488,N_16804);
nor U18391 (N_18391,N_17171,N_15563);
and U18392 (N_18392,N_17693,N_15012);
nor U18393 (N_18393,N_16797,N_16706);
or U18394 (N_18394,N_16916,N_16973);
xnor U18395 (N_18395,N_16132,N_16678);
nand U18396 (N_18396,N_17213,N_17039);
xnor U18397 (N_18397,N_17193,N_15607);
or U18398 (N_18398,N_15476,N_17344);
or U18399 (N_18399,N_16600,N_16387);
and U18400 (N_18400,N_17560,N_15962);
nor U18401 (N_18401,N_15881,N_16038);
nand U18402 (N_18402,N_15843,N_15719);
and U18403 (N_18403,N_15376,N_15758);
and U18404 (N_18404,N_16046,N_17019);
nand U18405 (N_18405,N_17276,N_17257);
nor U18406 (N_18406,N_17723,N_15998);
xnor U18407 (N_18407,N_15656,N_15111);
or U18408 (N_18408,N_15378,N_15770);
xnor U18409 (N_18409,N_16087,N_16140);
or U18410 (N_18410,N_17659,N_16529);
nand U18411 (N_18411,N_15590,N_15134);
nor U18412 (N_18412,N_16335,N_15380);
or U18413 (N_18413,N_15555,N_15312);
or U18414 (N_18414,N_17435,N_16011);
and U18415 (N_18415,N_15718,N_16212);
nor U18416 (N_18416,N_17525,N_17683);
and U18417 (N_18417,N_17717,N_16406);
or U18418 (N_18418,N_17328,N_17394);
xor U18419 (N_18419,N_16893,N_15915);
or U18420 (N_18420,N_17195,N_16848);
and U18421 (N_18421,N_17772,N_15124);
xor U18422 (N_18422,N_17722,N_17122);
nor U18423 (N_18423,N_17059,N_15922);
nand U18424 (N_18424,N_17312,N_17600);
xor U18425 (N_18425,N_15280,N_15196);
and U18426 (N_18426,N_16304,N_16205);
nor U18427 (N_18427,N_17384,N_17733);
nor U18428 (N_18428,N_15043,N_17822);
nor U18429 (N_18429,N_17253,N_15892);
xor U18430 (N_18430,N_16686,N_17308);
xor U18431 (N_18431,N_16265,N_15383);
or U18432 (N_18432,N_16640,N_15180);
or U18433 (N_18433,N_16419,N_15693);
nand U18434 (N_18434,N_17749,N_17814);
nand U18435 (N_18435,N_16735,N_17826);
xnor U18436 (N_18436,N_17307,N_15575);
nor U18437 (N_18437,N_16579,N_16614);
and U18438 (N_18438,N_16922,N_15118);
nand U18439 (N_18439,N_15873,N_16633);
or U18440 (N_18440,N_15253,N_15774);
nand U18441 (N_18441,N_16681,N_16540);
and U18442 (N_18442,N_15474,N_16660);
and U18443 (N_18443,N_17003,N_16613);
nand U18444 (N_18444,N_16879,N_15619);
or U18445 (N_18445,N_16107,N_16454);
nor U18446 (N_18446,N_17756,N_15354);
nor U18447 (N_18447,N_16960,N_15096);
or U18448 (N_18448,N_15032,N_15098);
nand U18449 (N_18449,N_16305,N_17673);
nand U18450 (N_18450,N_16511,N_15574);
xor U18451 (N_18451,N_16615,N_17958);
nor U18452 (N_18452,N_17336,N_16941);
xnor U18453 (N_18453,N_15798,N_16393);
nor U18454 (N_18454,N_16250,N_17087);
nand U18455 (N_18455,N_17013,N_16911);
nand U18456 (N_18456,N_15964,N_17802);
nor U18457 (N_18457,N_16514,N_16699);
or U18458 (N_18458,N_15465,N_16644);
or U18459 (N_18459,N_16061,N_15407);
or U18460 (N_18460,N_16860,N_17937);
nand U18461 (N_18461,N_15728,N_16238);
xor U18462 (N_18462,N_17942,N_16292);
and U18463 (N_18463,N_17353,N_16267);
nor U18464 (N_18464,N_16173,N_16104);
nor U18465 (N_18465,N_15265,N_16095);
or U18466 (N_18466,N_15498,N_17721);
and U18467 (N_18467,N_15042,N_15778);
and U18468 (N_18468,N_15050,N_17748);
nor U18469 (N_18469,N_15699,N_17273);
xor U18470 (N_18470,N_17318,N_16902);
nor U18471 (N_18471,N_16884,N_17590);
nor U18472 (N_18472,N_16101,N_15623);
nor U18473 (N_18473,N_16720,N_15713);
nand U18474 (N_18474,N_15357,N_17186);
and U18475 (N_18475,N_15413,N_16620);
and U18476 (N_18476,N_16863,N_15662);
nand U18477 (N_18477,N_17022,N_15018);
nand U18478 (N_18478,N_16522,N_15468);
and U18479 (N_18479,N_16581,N_15386);
xor U18480 (N_18480,N_17503,N_15139);
and U18481 (N_18481,N_15507,N_16469);
nor U18482 (N_18482,N_15137,N_16619);
nor U18483 (N_18483,N_17467,N_17277);
nor U18484 (N_18484,N_16193,N_15437);
or U18485 (N_18485,N_15190,N_15530);
or U18486 (N_18486,N_17072,N_17665);
nor U18487 (N_18487,N_17283,N_17573);
xnor U18488 (N_18488,N_17295,N_15234);
nor U18489 (N_18489,N_16442,N_17153);
nand U18490 (N_18490,N_16426,N_16202);
xor U18491 (N_18491,N_17685,N_17853);
xnor U18492 (N_18492,N_15067,N_17752);
xor U18493 (N_18493,N_15589,N_15742);
nor U18494 (N_18494,N_15064,N_16018);
nand U18495 (N_18495,N_15611,N_17768);
nor U18496 (N_18496,N_15159,N_17612);
xnor U18497 (N_18497,N_17541,N_15223);
xnor U18498 (N_18498,N_16906,N_15790);
nor U18499 (N_18499,N_15314,N_17687);
nand U18500 (N_18500,N_15504,N_16761);
or U18501 (N_18501,N_16076,N_17860);
xor U18502 (N_18502,N_17542,N_15844);
nor U18503 (N_18503,N_17807,N_17941);
nand U18504 (N_18504,N_16610,N_16188);
nand U18505 (N_18505,N_17846,N_15582);
xnor U18506 (N_18506,N_16157,N_15119);
nor U18507 (N_18507,N_17115,N_15677);
nand U18508 (N_18508,N_17146,N_15814);
nand U18509 (N_18509,N_15167,N_17639);
and U18510 (N_18510,N_17696,N_17197);
and U18511 (N_18511,N_15338,N_16213);
nand U18512 (N_18512,N_16124,N_17027);
xor U18513 (N_18513,N_17092,N_15630);
nor U18514 (N_18514,N_15496,N_16390);
nand U18515 (N_18515,N_17096,N_15269);
nand U18516 (N_18516,N_17922,N_17292);
and U18517 (N_18517,N_17356,N_15518);
nand U18518 (N_18518,N_16162,N_16093);
nor U18519 (N_18519,N_17293,N_15502);
and U18520 (N_18520,N_17586,N_15544);
and U18521 (N_18521,N_17650,N_16571);
and U18522 (N_18522,N_16742,N_15430);
xnor U18523 (N_18523,N_16588,N_17229);
nor U18524 (N_18524,N_15643,N_16515);
and U18525 (N_18525,N_17382,N_17177);
and U18526 (N_18526,N_16378,N_16062);
nand U18527 (N_18527,N_17427,N_16585);
and U18528 (N_18528,N_15276,N_17051);
and U18529 (N_18529,N_16142,N_16464);
nor U18530 (N_18530,N_16034,N_17652);
and U18531 (N_18531,N_17859,N_16763);
or U18532 (N_18532,N_16398,N_16943);
nor U18533 (N_18533,N_17699,N_15062);
or U18534 (N_18534,N_17636,N_15059);
or U18535 (N_18535,N_17487,N_17028);
or U18536 (N_18536,N_16685,N_17199);
xnor U18537 (N_18537,N_16794,N_15406);
or U18538 (N_18538,N_17303,N_17762);
nor U18539 (N_18539,N_16272,N_15851);
and U18540 (N_18540,N_16697,N_15869);
nor U18541 (N_18541,N_17547,N_17379);
nor U18542 (N_18542,N_15566,N_15092);
xor U18543 (N_18543,N_16687,N_15242);
and U18544 (N_18544,N_15525,N_16591);
nor U18545 (N_18545,N_16962,N_17701);
or U18546 (N_18546,N_15011,N_17141);
nand U18547 (N_18547,N_15135,N_15825);
xnor U18548 (N_18548,N_17820,N_17334);
nor U18549 (N_18549,N_15716,N_17077);
nand U18550 (N_18550,N_15766,N_16659);
nor U18551 (N_18551,N_15666,N_17517);
and U18552 (N_18552,N_17256,N_17361);
or U18553 (N_18553,N_17222,N_16376);
nand U18554 (N_18554,N_15371,N_15552);
nor U18555 (N_18555,N_17118,N_15094);
or U18556 (N_18556,N_17874,N_15398);
or U18557 (N_18557,N_15461,N_16721);
nand U18558 (N_18558,N_16501,N_16020);
nand U18559 (N_18559,N_17494,N_15303);
xnor U18560 (N_18560,N_17498,N_16402);
nand U18561 (N_18561,N_17818,N_15885);
or U18562 (N_18562,N_16211,N_16667);
or U18563 (N_18563,N_16625,N_15557);
nand U18564 (N_18564,N_17741,N_15444);
or U18565 (N_18565,N_16750,N_15791);
nand U18566 (N_18566,N_17062,N_15686);
nand U18567 (N_18567,N_17831,N_17397);
and U18568 (N_18568,N_15857,N_16458);
xor U18569 (N_18569,N_15705,N_15310);
xnor U18570 (N_18570,N_15992,N_15800);
or U18571 (N_18571,N_17649,N_17803);
and U18572 (N_18572,N_17672,N_15914);
nand U18573 (N_18573,N_16429,N_16024);
and U18574 (N_18574,N_16796,N_15299);
and U18575 (N_18575,N_16182,N_16556);
nand U18576 (N_18576,N_16778,N_17877);
or U18577 (N_18577,N_17761,N_17182);
or U18578 (N_18578,N_16164,N_16850);
or U18579 (N_18579,N_16374,N_15487);
xor U18580 (N_18580,N_17202,N_15913);
or U18581 (N_18581,N_16044,N_15906);
xnor U18582 (N_18582,N_17994,N_16682);
xnor U18583 (N_18583,N_17747,N_17206);
nor U18584 (N_18584,N_16059,N_15185);
and U18585 (N_18585,N_17326,N_15405);
or U18586 (N_18586,N_15867,N_16729);
and U18587 (N_18587,N_16291,N_17418);
xnor U18588 (N_18588,N_17970,N_17899);
nand U18589 (N_18589,N_16340,N_16920);
and U18590 (N_18590,N_17591,N_16596);
xnor U18591 (N_18591,N_15896,N_17521);
or U18592 (N_18592,N_16532,N_16085);
xor U18593 (N_18593,N_17806,N_16251);
or U18594 (N_18594,N_17862,N_15739);
and U18595 (N_18595,N_17908,N_17392);
nand U18596 (N_18596,N_16837,N_17068);
or U18597 (N_18597,N_16479,N_17460);
or U18598 (N_18598,N_16273,N_16719);
nand U18599 (N_18599,N_16445,N_17601);
nor U18600 (N_18600,N_17074,N_16636);
xor U18601 (N_18601,N_17201,N_17963);
and U18602 (N_18602,N_16149,N_15514);
nor U18603 (N_18603,N_17849,N_16350);
xnor U18604 (N_18604,N_15087,N_15290);
or U18605 (N_18605,N_15077,N_16192);
nand U18606 (N_18606,N_16709,N_16871);
nor U18607 (N_18607,N_15379,N_17983);
or U18608 (N_18608,N_16518,N_16563);
nor U18609 (N_18609,N_15875,N_15908);
nor U18610 (N_18610,N_17109,N_17532);
or U18611 (N_18611,N_17180,N_16628);
xnor U18612 (N_18612,N_16241,N_17495);
or U18613 (N_18613,N_16358,N_15500);
and U18614 (N_18614,N_16118,N_15980);
or U18615 (N_18615,N_16473,N_15894);
xnor U18616 (N_18616,N_15632,N_17357);
or U18617 (N_18617,N_15609,N_17992);
or U18618 (N_18618,N_15150,N_16710);
and U18619 (N_18619,N_15550,N_17314);
xor U18620 (N_18620,N_16717,N_17404);
nor U18621 (N_18621,N_17644,N_15862);
nor U18622 (N_18622,N_15568,N_16817);
nor U18623 (N_18623,N_15275,N_16032);
xor U18624 (N_18624,N_15392,N_16852);
nand U18625 (N_18625,N_16680,N_17006);
nor U18626 (N_18626,N_17797,N_17571);
xor U18627 (N_18627,N_17098,N_16723);
or U18628 (N_18628,N_16025,N_17126);
or U18629 (N_18629,N_16711,N_17136);
or U18630 (N_18630,N_16239,N_16232);
xor U18631 (N_18631,N_15819,N_15903);
nand U18632 (N_18632,N_17835,N_17055);
nand U18633 (N_18633,N_17354,N_15366);
nand U18634 (N_18634,N_17375,N_17035);
and U18635 (N_18635,N_17840,N_17555);
nand U18636 (N_18636,N_16494,N_16283);
nand U18637 (N_18637,N_16326,N_15285);
xnor U18638 (N_18638,N_17546,N_17526);
xnor U18639 (N_18639,N_15146,N_15300);
nand U18640 (N_18640,N_16502,N_16967);
xnor U18641 (N_18641,N_15969,N_15600);
nand U18642 (N_18642,N_17648,N_15744);
nand U18643 (N_18643,N_16052,N_17884);
and U18644 (N_18644,N_15188,N_16203);
and U18645 (N_18645,N_15928,N_17461);
nor U18646 (N_18646,N_16258,N_17041);
or U18647 (N_18647,N_16972,N_15848);
and U18648 (N_18648,N_15129,N_16574);
nor U18649 (N_18649,N_16277,N_17358);
xnor U18650 (N_18650,N_15233,N_17790);
or U18651 (N_18651,N_16191,N_15198);
nand U18652 (N_18652,N_17204,N_15711);
or U18653 (N_18653,N_15439,N_16263);
nand U18654 (N_18654,N_17224,N_16658);
and U18655 (N_18655,N_15326,N_16102);
nor U18656 (N_18656,N_15868,N_16153);
xor U18657 (N_18657,N_16339,N_17730);
nand U18658 (N_18658,N_15245,N_15904);
and U18659 (N_18659,N_15919,N_16438);
or U18660 (N_18660,N_16016,N_16279);
nor U18661 (N_18661,N_17289,N_17943);
nand U18662 (N_18662,N_15154,N_15367);
nor U18663 (N_18663,N_16886,N_15112);
or U18664 (N_18664,N_17712,N_15440);
nor U18665 (N_18665,N_15849,N_15893);
nand U18666 (N_18666,N_15986,N_16618);
nor U18667 (N_18667,N_15785,N_15640);
nand U18668 (N_18668,N_17815,N_15202);
or U18669 (N_18669,N_17212,N_15977);
and U18670 (N_18670,N_15352,N_17651);
and U18671 (N_18671,N_16849,N_16066);
nand U18672 (N_18672,N_16942,N_16297);
and U18673 (N_18673,N_16958,N_16226);
xnor U18674 (N_18674,N_16684,N_15168);
or U18675 (N_18675,N_16575,N_15423);
nand U18676 (N_18676,N_16395,N_16332);
nor U18677 (N_18677,N_15840,N_15400);
or U18678 (N_18678,N_15262,N_15531);
nand U18679 (N_18679,N_17854,N_16289);
nand U18680 (N_18680,N_16070,N_15821);
nor U18681 (N_18681,N_15497,N_16158);
nand U18682 (N_18682,N_15220,N_15803);
nor U18683 (N_18683,N_16940,N_16938);
or U18684 (N_18684,N_16855,N_17969);
and U18685 (N_18685,N_17898,N_16506);
and U18686 (N_18686,N_15897,N_16937);
or U18687 (N_18687,N_17033,N_16576);
or U18688 (N_18688,N_15529,N_17738);
nand U18689 (N_18689,N_15221,N_16754);
nor U18690 (N_18690,N_15293,N_15668);
nor U18691 (N_18691,N_16749,N_16361);
nand U18692 (N_18692,N_17655,N_17137);
and U18693 (N_18693,N_17169,N_16073);
xor U18694 (N_18694,N_15949,N_16747);
nand U18695 (N_18695,N_15105,N_16423);
and U18696 (N_18696,N_16083,N_17527);
xnor U18697 (N_18697,N_15524,N_16616);
nor U18698 (N_18698,N_16769,N_15415);
nor U18699 (N_18699,N_16343,N_16219);
xor U18700 (N_18700,N_15966,N_16873);
nand U18701 (N_18701,N_15622,N_15072);
or U18702 (N_18702,N_15567,N_15289);
and U18703 (N_18703,N_16240,N_15268);
xnor U18704 (N_18704,N_15131,N_16826);
and U18705 (N_18705,N_17341,N_16181);
and U18706 (N_18706,N_17754,N_16641);
nor U18707 (N_18707,N_16215,N_15006);
nand U18708 (N_18708,N_16695,N_17531);
nor U18709 (N_18709,N_15478,N_17160);
nand U18710 (N_18710,N_16961,N_16583);
nor U18711 (N_18711,N_17053,N_16180);
or U18712 (N_18712,N_16919,N_17758);
nor U18713 (N_18713,N_17483,N_16383);
or U18714 (N_18714,N_15697,N_16225);
or U18715 (N_18715,N_15916,N_17504);
or U18716 (N_18716,N_16523,N_15254);
xnor U18717 (N_18717,N_15078,N_16538);
nor U18718 (N_18718,N_15107,N_16525);
nand U18719 (N_18719,N_15694,N_15325);
nand U18720 (N_18720,N_16923,N_16119);
nand U18721 (N_18721,N_17520,N_15971);
xor U18722 (N_18722,N_16151,N_15789);
nor U18723 (N_18723,N_17472,N_15153);
and U18724 (N_18724,N_16768,N_15735);
xor U18725 (N_18725,N_17851,N_17798);
xor U18726 (N_18726,N_17377,N_16360);
xnor U18727 (N_18727,N_15571,N_17794);
or U18728 (N_18728,N_16007,N_17061);
and U18729 (N_18729,N_17522,N_16167);
nor U18730 (N_18730,N_16621,N_16098);
and U18731 (N_18731,N_17271,N_15360);
or U18732 (N_18732,N_17778,N_16572);
and U18733 (N_18733,N_16969,N_15066);
xor U18734 (N_18734,N_15037,N_17534);
and U18735 (N_18735,N_15665,N_15784);
nor U18736 (N_18736,N_17409,N_15509);
or U18737 (N_18737,N_15256,N_16227);
xnor U18738 (N_18738,N_15344,N_15882);
and U18739 (N_18739,N_17615,N_15364);
nor U18740 (N_18740,N_16650,N_16517);
nor U18741 (N_18741,N_17934,N_17708);
or U18742 (N_18742,N_16313,N_16546);
or U18743 (N_18743,N_16568,N_17247);
and U18744 (N_18744,N_17606,N_15214);
and U18745 (N_18745,N_17393,N_15559);
nor U18746 (N_18746,N_15664,N_17950);
nand U18747 (N_18747,N_16877,N_16138);
or U18748 (N_18748,N_17164,N_15433);
xor U18749 (N_18749,N_17878,N_16925);
nor U18750 (N_18750,N_17065,N_17781);
nand U18751 (N_18751,N_17249,N_15905);
and U18752 (N_18752,N_16047,N_17045);
or U18753 (N_18753,N_16521,N_16447);
nand U18754 (N_18754,N_16980,N_15641);
and U18755 (N_18755,N_17881,N_15266);
nor U18756 (N_18756,N_16807,N_16617);
and U18757 (N_18757,N_15192,N_16030);
or U18758 (N_18758,N_17438,N_16143);
and U18759 (N_18759,N_15084,N_15004);
nor U18760 (N_18760,N_17402,N_16828);
nand U18761 (N_18761,N_17677,N_15047);
or U18762 (N_18762,N_17173,N_16299);
or U18763 (N_18763,N_15000,N_17238);
nand U18764 (N_18764,N_16389,N_17745);
nand U18765 (N_18765,N_15492,N_15255);
and U18766 (N_18766,N_15817,N_16462);
nor U18767 (N_18767,N_17932,N_15826);
nor U18768 (N_18768,N_16417,N_17513);
or U18769 (N_18769,N_15115,N_17108);
and U18770 (N_18770,N_15141,N_15700);
or U18771 (N_18771,N_17448,N_16975);
nand U18772 (N_18772,N_17478,N_17221);
nand U18773 (N_18773,N_15211,N_16077);
nor U18774 (N_18774,N_16859,N_16231);
xor U18775 (N_18775,N_16489,N_17728);
xor U18776 (N_18776,N_16049,N_17732);
or U18777 (N_18777,N_16017,N_17771);
or U18778 (N_18778,N_16724,N_15200);
or U18779 (N_18779,N_15934,N_16780);
nand U18780 (N_18780,N_15957,N_16163);
nor U18781 (N_18781,N_16000,N_16481);
nand U18782 (N_18782,N_17654,N_17004);
or U18783 (N_18783,N_17232,N_15363);
and U18784 (N_18784,N_15564,N_16333);
xnor U18785 (N_18785,N_15690,N_15395);
nand U18786 (N_18786,N_16701,N_16109);
nand U18787 (N_18787,N_15608,N_17489);
and U18788 (N_18788,N_15832,N_17947);
nor U18789 (N_18789,N_16266,N_16336);
xor U18790 (N_18790,N_17538,N_15714);
nand U18791 (N_18791,N_16112,N_15506);
and U18792 (N_18792,N_17011,N_15717);
or U18793 (N_18793,N_15594,N_17036);
xor U18794 (N_18794,N_15239,N_16122);
xnor U18795 (N_18795,N_15170,N_16391);
or U18796 (N_18796,N_17812,N_17023);
xnor U18797 (N_18797,N_17642,N_17582);
nor U18798 (N_18798,N_15649,N_16979);
and U18799 (N_18799,N_16779,N_17767);
nand U18800 (N_18800,N_17014,N_16554);
or U18801 (N_18801,N_17288,N_16516);
nand U18802 (N_18802,N_15516,N_17405);
nor U18803 (N_18803,N_17364,N_15373);
nor U18804 (N_18804,N_16932,N_15259);
xnor U18805 (N_18805,N_16131,N_15780);
nand U18806 (N_18806,N_15633,N_15085);
xnor U18807 (N_18807,N_17459,N_17267);
nand U18808 (N_18808,N_15660,N_17386);
xnor U18809 (N_18809,N_15370,N_16531);
or U18810 (N_18810,N_15508,N_15963);
and U18811 (N_18811,N_17071,N_15769);
or U18812 (N_18812,N_15989,N_15930);
or U18813 (N_18813,N_15763,N_15035);
and U18814 (N_18814,N_15542,N_15421);
and U18815 (N_18815,N_17484,N_15473);
and U18816 (N_18816,N_17127,N_16463);
or U18817 (N_18817,N_16654,N_17903);
nand U18818 (N_18818,N_15136,N_17242);
xor U18819 (N_18819,N_15116,N_15898);
and U18820 (N_18820,N_16558,N_16178);
nand U18821 (N_18821,N_17653,N_15075);
or U18822 (N_18822,N_15852,N_16121);
nand U18823 (N_18823,N_15187,N_16889);
and U18824 (N_18824,N_17369,N_17763);
and U18825 (N_18825,N_15183,N_16475);
nor U18826 (N_18826,N_16643,N_17610);
and U18827 (N_18827,N_15806,N_15837);
or U18828 (N_18828,N_17637,N_17609);
nand U18829 (N_18829,N_15993,N_17390);
nor U18830 (N_18830,N_16888,N_16234);
nand U18831 (N_18831,N_15824,N_17029);
xnor U18832 (N_18832,N_17604,N_16810);
nand U18833 (N_18833,N_15397,N_15709);
nand U18834 (N_18834,N_15537,N_16984);
xor U18835 (N_18835,N_17896,N_17593);
nand U18836 (N_18836,N_16466,N_15236);
xor U18837 (N_18837,N_16666,N_17403);
or U18838 (N_18838,N_16741,N_17927);
and U18839 (N_18839,N_17829,N_17291);
nor U18840 (N_18840,N_17868,N_16461);
nand U18841 (N_18841,N_17588,N_17518);
xnor U18842 (N_18842,N_15287,N_17281);
or U18843 (N_18843,N_15080,N_15396);
and U18844 (N_18844,N_17939,N_15816);
or U18845 (N_18845,N_15279,N_16113);
or U18846 (N_18846,N_16833,N_15771);
and U18847 (N_18847,N_16123,N_17130);
nor U18848 (N_18848,N_15034,N_15570);
or U18849 (N_18849,N_15033,N_17152);
nand U18850 (N_18850,N_16249,N_17617);
and U18851 (N_18851,N_15865,N_16410);
nand U18852 (N_18852,N_15399,N_16448);
nand U18853 (N_18853,N_15511,N_16281);
nor U18854 (N_18854,N_16453,N_16029);
and U18855 (N_18855,N_16611,N_16441);
xor U18856 (N_18856,N_15779,N_17989);
or U18857 (N_18857,N_16597,N_16357);
and U18858 (N_18858,N_17952,N_15805);
and U18859 (N_18859,N_16549,N_15333);
xnor U18860 (N_18860,N_15368,N_15975);
nor U18861 (N_18861,N_16696,N_17114);
nor U18862 (N_18862,N_16342,N_15061);
xnor U18863 (N_18863,N_15639,N_17315);
nor U18864 (N_18864,N_15418,N_17883);
nor U18865 (N_18865,N_17134,N_17031);
nor U18866 (N_18866,N_17032,N_16808);
nor U18867 (N_18867,N_15762,N_16770);
nand U18868 (N_18868,N_17280,N_15887);
nor U18869 (N_18869,N_15682,N_15935);
xnor U18870 (N_18870,N_17082,N_16370);
nor U18871 (N_18871,N_17979,N_15316);
nand U18872 (N_18872,N_17594,N_17982);
nand U18873 (N_18873,N_15044,N_15204);
xor U18874 (N_18874,N_16474,N_17254);
nor U18875 (N_18875,N_17966,N_17894);
nor U18876 (N_18876,N_15727,N_16624);
nand U18877 (N_18877,N_16939,N_16559);
and U18878 (N_18878,N_16430,N_16040);
or U18879 (N_18879,N_15375,N_15472);
or U18880 (N_18880,N_16836,N_17581);
xnor U18881 (N_18881,N_16765,N_16601);
and U18882 (N_18882,N_16400,N_17506);
or U18883 (N_18883,N_16782,N_15244);
or U18884 (N_18884,N_17578,N_17380);
xor U18885 (N_18885,N_16974,N_17340);
and U18886 (N_18886,N_15994,N_16134);
nor U18887 (N_18887,N_17724,N_17845);
xor U18888 (N_18888,N_16885,N_16221);
nor U18889 (N_18889,N_16844,N_16455);
xnor U18890 (N_18890,N_15616,N_15458);
nand U18891 (N_18891,N_17012,N_17198);
or U18892 (N_18892,N_16876,N_17084);
or U18893 (N_18893,N_17961,N_16125);
or U18894 (N_18894,N_16428,N_17362);
nor U18895 (N_18895,N_17246,N_15247);
or U18896 (N_18896,N_15226,N_16110);
nand U18897 (N_18897,N_17613,N_17097);
nor U18898 (N_18898,N_17501,N_15297);
xnor U18899 (N_18899,N_17282,N_17428);
xnor U18900 (N_18900,N_17396,N_17559);
or U18901 (N_18901,N_17431,N_16156);
nand U18902 (N_18902,N_16580,N_17373);
and U18903 (N_18903,N_17686,N_15446);
or U18904 (N_18904,N_15114,N_17047);
xnor U18905 (N_18905,N_15455,N_17879);
or U18906 (N_18906,N_15750,N_15912);
nor U18907 (N_18907,N_17454,N_16707);
xnor U18908 (N_18908,N_16200,N_16752);
nor U18909 (N_18909,N_16444,N_15486);
nand U18910 (N_18910,N_17817,N_17551);
and U18911 (N_18911,N_16561,N_17161);
xor U18912 (N_18912,N_17112,N_15243);
and U18913 (N_18913,N_17530,N_17462);
nor U18914 (N_18914,N_17984,N_16553);
xnor U18915 (N_18915,N_15820,N_16993);
nor U18916 (N_18916,N_17985,N_16345);
xor U18917 (N_18917,N_15972,N_16630);
xor U18918 (N_18918,N_16675,N_17167);
nor U18919 (N_18919,N_17217,N_16803);
or U18920 (N_18920,N_15583,N_15889);
and U18921 (N_18921,N_16276,N_16255);
xnor U18922 (N_18922,N_17086,N_17227);
xor U18923 (N_18923,N_17138,N_17828);
and U18924 (N_18924,N_15412,N_15657);
xor U18925 (N_18925,N_16820,N_16792);
nor U18926 (N_18926,N_15009,N_15604);
nand U18927 (N_18927,N_17479,N_16936);
nor U18928 (N_18928,N_15947,N_17166);
or U18929 (N_18929,N_15603,N_17713);
xor U18930 (N_18930,N_16843,N_16552);
xor U18931 (N_18931,N_15491,N_16609);
and U18932 (N_18932,N_15385,N_17417);
xor U18933 (N_18933,N_16039,N_17666);
xor U18934 (N_18934,N_16413,N_15477);
nor U18935 (N_18935,N_16565,N_15688);
and U18936 (N_18936,N_16068,N_17060);
xnor U18937 (N_18937,N_16359,N_17080);
or U18938 (N_18938,N_17905,N_16168);
nor U18939 (N_18939,N_16088,N_17240);
nor U18940 (N_18940,N_16259,N_16009);
xor U18941 (N_18941,N_16290,N_17188);
or U18942 (N_18942,N_16187,N_15667);
nor U18943 (N_18943,N_15228,N_16996);
nor U18944 (N_18944,N_17269,N_17965);
nor U18945 (N_18945,N_15069,N_16744);
or U18946 (N_18946,N_15505,N_15060);
xor U18947 (N_18947,N_15878,N_17030);
or U18948 (N_18948,N_17647,N_17684);
nand U18949 (N_18949,N_15401,N_17836);
and U18950 (N_18950,N_16507,N_15470);
and U18951 (N_18951,N_15561,N_15990);
nand U18952 (N_18952,N_16363,N_16935);
or U18953 (N_18953,N_16542,N_17557);
and U18954 (N_18954,N_17809,N_17170);
or U18955 (N_18955,N_17562,N_15130);
nand U18956 (N_18956,N_17090,N_17889);
nand U18957 (N_18957,N_16533,N_17450);
and U18958 (N_18958,N_17233,N_17104);
and U18959 (N_18959,N_16084,N_15598);
nor U18960 (N_18960,N_15110,N_17949);
xor U18961 (N_18961,N_16375,N_15517);
nor U18962 (N_18962,N_16632,N_16802);
and U18963 (N_18963,N_17663,N_17187);
xor U18964 (N_18964,N_17576,N_16688);
or U18965 (N_18965,N_15264,N_15302);
nand U18966 (N_18966,N_16964,N_16210);
or U18967 (N_18967,N_17154,N_17196);
xor U18968 (N_18968,N_15391,N_15535);
xor U18969 (N_18969,N_17599,N_16530);
and U18970 (N_18970,N_17002,N_15858);
and U18971 (N_18971,N_16599,N_16043);
nor U18972 (N_18972,N_16824,N_16756);
nor U18973 (N_18973,N_17698,N_17389);
nand U18974 (N_18974,N_17681,N_15834);
or U18975 (N_18975,N_16394,N_17930);
or U18976 (N_18976,N_17131,N_17189);
xor U18977 (N_18977,N_17919,N_16329);
nand U18978 (N_18978,N_17833,N_15822);
nand U18979 (N_18979,N_16353,N_17856);
or U18980 (N_18980,N_17366,N_17974);
or U18981 (N_18981,N_16997,N_16512);
xor U18982 (N_18982,N_15651,N_16703);
xnor U18983 (N_18983,N_15144,N_17844);
or U18984 (N_18984,N_15546,N_17524);
nand U18985 (N_18985,N_16566,N_15347);
nand U18986 (N_18986,N_15216,N_15002);
and U18987 (N_18987,N_16731,N_15252);
nand U18988 (N_18988,N_15175,N_17704);
and U18989 (N_18989,N_15548,N_15628);
nand U18990 (N_18990,N_17773,N_16878);
or U18991 (N_18991,N_17040,N_17018);
xnor U18992 (N_18992,N_16665,N_16670);
and U18993 (N_18993,N_17338,N_16679);
nor U18994 (N_18994,N_15708,N_16256);
xnor U18995 (N_18995,N_16456,N_17736);
xor U18996 (N_18996,N_17103,N_17449);
nand U18997 (N_18997,N_16172,N_17423);
nor U18998 (N_18998,N_15646,N_17589);
or U18999 (N_18999,N_16351,N_15856);
nand U19000 (N_19000,N_15793,N_17788);
nand U19001 (N_19001,N_16060,N_17575);
and U19002 (N_19002,N_15133,N_16146);
xnor U19003 (N_19003,N_16951,N_17129);
xnor U19004 (N_19004,N_15480,N_17139);
and U19005 (N_19005,N_16793,N_15053);
xor U19006 (N_19006,N_15339,N_16317);
nor U19007 (N_19007,N_15936,N_15792);
nand U19008 (N_19008,N_17523,N_15983);
and U19009 (N_19009,N_15318,N_16508);
nor U19010 (N_19010,N_16933,N_16485);
nand U19011 (N_19011,N_15845,N_16781);
or U19012 (N_19012,N_17598,N_16099);
and U19013 (N_19013,N_16510,N_17485);
nand U19014 (N_19014,N_17777,N_17734);
nand U19015 (N_19015,N_17995,N_17882);
xnor U19016 (N_19016,N_17669,N_15231);
and U19017 (N_19017,N_16082,N_15499);
or U19018 (N_19018,N_16248,N_15538);
nor U19019 (N_19019,N_16904,N_17640);
nor U19020 (N_19020,N_16758,N_15939);
xnor U19021 (N_19021,N_15113,N_16197);
nor U19022 (N_19022,N_17107,N_17678);
xnor U19023 (N_19023,N_16254,N_16653);
xnor U19024 (N_19024,N_17918,N_15071);
xnor U19025 (N_19025,N_17901,N_17432);
nor U19026 (N_19026,N_15637,N_17800);
xnor U19027 (N_19027,N_16825,N_17629);
or U19028 (N_19028,N_17351,N_16520);
nor U19029 (N_19029,N_16921,N_17584);
nor U19030 (N_19030,N_17711,N_17106);
nor U19031 (N_19031,N_16548,N_17488);
and U19032 (N_19032,N_16505,N_16541);
nor U19033 (N_19033,N_17492,N_16814);
nand U19034 (N_19034,N_15921,N_17998);
nand U19035 (N_19035,N_15489,N_17962);
nor U19036 (N_19036,N_16892,N_16480);
nor U19037 (N_19037,N_17697,N_17219);
nor U19038 (N_19038,N_15652,N_15584);
nand U19039 (N_19039,N_16477,N_15828);
nor U19040 (N_19040,N_17264,N_15387);
or U19041 (N_19041,N_15847,N_17192);
nand U19042 (N_19042,N_15014,N_16881);
nand U19043 (N_19043,N_17085,N_15618);
xor U19044 (N_19044,N_16528,N_15768);
or U19045 (N_19045,N_15467,N_15208);
nor U19046 (N_19046,N_16420,N_16063);
or U19047 (N_19047,N_16487,N_16058);
nand U19048 (N_19048,N_15911,N_16851);
nor U19049 (N_19049,N_17116,N_17147);
or U19050 (N_19050,N_16460,N_15539);
nand U19051 (N_19051,N_15974,N_15874);
and U19052 (N_19052,N_16015,N_17165);
xor U19053 (N_19053,N_16451,N_17420);
nand U19054 (N_19054,N_16986,N_16365);
or U19055 (N_19055,N_15218,N_15715);
nand U19056 (N_19056,N_16199,N_16069);
xor U19057 (N_19057,N_16764,N_15827);
or U19058 (N_19058,N_15764,N_16914);
xnor U19059 (N_19059,N_15812,N_16981);
and U19060 (N_19060,N_15369,N_17049);
or U19061 (N_19061,N_17872,N_15057);
nand U19062 (N_19062,N_16307,N_15331);
nand U19063 (N_19063,N_17349,N_15058);
or U19064 (N_19064,N_15724,N_15164);
and U19065 (N_19065,N_17751,N_15017);
and U19066 (N_19066,N_15291,N_17959);
xnor U19067 (N_19067,N_15526,N_17997);
xnor U19068 (N_19068,N_15241,N_15796);
or U19069 (N_19069,N_15462,N_16683);
nor U19070 (N_19070,N_15295,N_15967);
and U19071 (N_19071,N_17641,N_17323);
nand U19072 (N_19072,N_17168,N_16757);
nand U19073 (N_19073,N_17925,N_16245);
nand U19074 (N_19074,N_17203,N_15040);
nand U19075 (N_19075,N_16195,N_15052);
nor U19076 (N_19076,N_15955,N_16582);
xor U19077 (N_19077,N_17348,N_15054);
nand U19078 (N_19078,N_17911,N_17215);
xnor U19079 (N_19079,N_17081,N_16385);
nand U19080 (N_19080,N_16795,N_17268);
nand U19081 (N_19081,N_15736,N_15794);
and U19082 (N_19082,N_16096,N_16864);
xor U19083 (N_19083,N_15503,N_17776);
or U19084 (N_19084,N_15647,N_15301);
and U19085 (N_19085,N_15140,N_16484);
xor U19086 (N_19086,N_15958,N_17832);
nor U19087 (N_19087,N_16284,N_16303);
nor U19088 (N_19088,N_15612,N_17178);
nand U19089 (N_19089,N_16745,N_17145);
xor U19090 (N_19090,N_16274,N_15041);
nor U19091 (N_19091,N_16657,N_17094);
or U19092 (N_19092,N_17999,N_17411);
xor U19093 (N_19093,N_16691,N_16260);
nand U19094 (N_19094,N_15585,N_16612);
or U19095 (N_19095,N_15404,N_17510);
nor U19096 (N_19096,N_16228,N_16114);
or U19097 (N_19097,N_17611,N_16457);
xor U19098 (N_19098,N_17631,N_15382);
or U19099 (N_19099,N_16957,N_15179);
nor U19100 (N_19100,N_15340,N_15946);
or U19101 (N_19101,N_17580,N_15212);
and U19102 (N_19102,N_17630,N_15215);
and U19103 (N_19103,N_16116,N_17124);
nor U19104 (N_19104,N_16001,N_16870);
or U19105 (N_19105,N_15165,N_15534);
nand U19106 (N_19106,N_15070,N_16694);
nand U19107 (N_19107,N_17442,N_16377);
nor U19108 (N_19108,N_15960,N_15854);
and U19109 (N_19109,N_15985,N_15872);
xor U19110 (N_19110,N_15460,N_17350);
or U19111 (N_19111,N_16693,N_17931);
or U19112 (N_19112,N_16349,N_17290);
nand U19113 (N_19113,N_16179,N_16772);
xor U19114 (N_19114,N_17343,N_16493);
nor U19115 (N_19115,N_17265,N_15536);
or U19116 (N_19116,N_17596,N_15624);
nor U19117 (N_19117,N_16314,N_17329);
xnor U19118 (N_19118,N_16161,N_17263);
and U19119 (N_19119,N_15510,N_15445);
or U19120 (N_19120,N_17888,N_17739);
or U19121 (N_19121,N_15673,N_15850);
nand U19122 (N_19122,N_15859,N_17430);
and U19123 (N_19123,N_17218,N_15620);
nand U19124 (N_19124,N_15251,N_15320);
xor U19125 (N_19125,N_17783,N_15024);
xnor U19126 (N_19126,N_16977,N_15670);
nand U19127 (N_19127,N_15169,N_17453);
xnor U19128 (N_19128,N_17046,N_17996);
or U19129 (N_19129,N_15540,N_15174);
or U19130 (N_19130,N_15103,N_15273);
or U19131 (N_19131,N_17691,N_15049);
or U19132 (N_19132,N_16985,N_17321);
nand U19133 (N_19133,N_15802,N_15995);
or U19134 (N_19134,N_15438,N_15880);
nand U19135 (N_19135,N_16050,N_17100);
nand U19136 (N_19136,N_15464,N_15156);
or U19137 (N_19137,N_16569,N_16715);
or U19138 (N_19138,N_15283,N_16954);
and U19139 (N_19139,N_15527,N_16926);
or U19140 (N_19140,N_15731,N_17572);
or U19141 (N_19141,N_17657,N_15063);
or U19142 (N_19142,N_16067,N_16652);
nor U19143 (N_19143,N_15520,N_15207);
and U19144 (N_19144,N_15853,N_16183);
xor U19145 (N_19145,N_15206,N_16784);
nor U19146 (N_19146,N_17159,N_15082);
nor U19147 (N_19147,N_17305,N_17056);
nand U19148 (N_19148,N_17556,N_16544);
or U19149 (N_19149,N_17563,N_16189);
nor U19150 (N_19150,N_17978,N_15635);
or U19151 (N_19151,N_16587,N_17044);
or U19152 (N_19152,N_16823,N_17330);
nor U19153 (N_19153,N_17407,N_15277);
and U19154 (N_19154,N_17345,N_17260);
nand U19155 (N_19155,N_17156,N_16705);
and U19156 (N_19156,N_17346,N_15621);
and U19157 (N_19157,N_17317,N_17936);
xor U19158 (N_19158,N_17387,N_16989);
and U19159 (N_19159,N_15811,N_15747);
nand U19160 (N_19160,N_15722,N_17381);
or U19161 (N_19161,N_17144,N_17789);
and U19162 (N_19162,N_17439,N_17890);
and U19163 (N_19163,N_15532,N_17861);
nand U19164 (N_19164,N_16809,N_15102);
nand U19165 (N_19165,N_15389,N_15815);
nand U19166 (N_19166,N_16910,N_16201);
or U19167 (N_19167,N_15929,N_15427);
xnor U19168 (N_19168,N_16648,N_15225);
xnor U19169 (N_19169,N_17142,N_15543);
xnor U19170 (N_19170,N_16036,N_16712);
and U19171 (N_19171,N_16865,N_16154);
nor U19172 (N_19172,N_15720,N_15838);
xnor U19173 (N_19173,N_15020,N_17455);
nor U19174 (N_19174,N_16835,N_16293);
xor U19175 (N_19175,N_16129,N_16261);
nand U19176 (N_19176,N_16037,N_17553);
and U19177 (N_19177,N_16392,N_17468);
xnor U19178 (N_19178,N_16899,N_15587);
and U19179 (N_19179,N_17515,N_16421);
xnor U19180 (N_19180,N_16722,N_15634);
and U19181 (N_19181,N_15046,N_16328);
xor U19182 (N_19182,N_15209,N_17753);
xor U19183 (N_19183,N_16857,N_15151);
nor U19184 (N_19184,N_15886,N_16325);
and U19185 (N_19185,N_17272,N_16371);
nor U19186 (N_19186,N_17643,N_16216);
nor U19187 (N_19187,N_16930,N_15723);
nand U19188 (N_19188,N_15712,N_17964);
or U19189 (N_19189,N_15606,N_17413);
nor U19190 (N_19190,N_17539,N_15562);
nand U19191 (N_19191,N_16545,N_15086);
nand U19192 (N_19192,N_15772,N_17322);
nor U19193 (N_19193,N_15781,N_16316);
or U19194 (N_19194,N_15927,N_17865);
nand U19195 (N_19195,N_17262,N_16500);
nand U19196 (N_19196,N_17944,N_15490);
and U19197 (N_19197,N_17110,N_17507);
or U19198 (N_19198,N_16381,N_17866);
or U19199 (N_19199,N_16918,N_16144);
nor U19200 (N_19200,N_15249,N_16748);
nand U19201 (N_19201,N_15488,N_17151);
nand U19202 (N_19202,N_17469,N_15533);
xnor U19203 (N_19203,N_17370,N_15475);
or U19204 (N_19204,N_16955,N_17597);
xor U19205 (N_19205,N_17953,N_15493);
or U19206 (N_19206,N_15410,N_17333);
or U19207 (N_19207,N_16006,N_17977);
nor U19208 (N_19208,N_15658,N_17048);
nor U19209 (N_19209,N_17766,N_17727);
and U19210 (N_19210,N_17497,N_16230);
xnor U19211 (N_19211,N_16434,N_17208);
nand U19212 (N_19212,N_17300,N_17990);
nand U19213 (N_19213,N_17863,N_16384);
and U19214 (N_19214,N_16403,N_15390);
nand U19215 (N_19215,N_17422,N_16867);
nand U19216 (N_19216,N_17900,N_17529);
nand U19217 (N_19217,N_17241,N_15288);
nor U19218 (N_19218,N_17093,N_15402);
nand U19219 (N_19219,N_15319,N_17909);
xor U19220 (N_19220,N_16425,N_15799);
or U19221 (N_19221,N_17912,N_17415);
nor U19222 (N_19222,N_16404,N_16295);
nand U19223 (N_19223,N_17891,N_17490);
nand U19224 (N_19224,N_16244,N_15831);
nor U19225 (N_19225,N_17395,N_15782);
or U19226 (N_19226,N_15349,N_15296);
and U19227 (N_19227,N_16799,N_16302);
nor U19228 (N_19228,N_16766,N_17286);
nand U19229 (N_19229,N_15203,N_15450);
nand U19230 (N_19230,N_17385,N_15240);
and U19231 (N_19231,N_15304,N_16543);
nor U19232 (N_19232,N_15556,N_16908);
nor U19233 (N_19233,N_16411,N_17928);
xor U19234 (N_19234,N_17975,N_17105);
and U19235 (N_19235,N_16041,N_16970);
and U19236 (N_19236,N_15810,N_15335);
nand U19237 (N_19237,N_15704,N_15191);
xnor U19238 (N_19238,N_16155,N_16965);
nor U19239 (N_19239,N_17671,N_15595);
nor U19240 (N_19240,N_16433,N_17414);
nand U19241 (N_19241,N_15519,N_17906);
nor U19242 (N_19242,N_17910,N_15959);
nor U19243 (N_19243,N_16341,N_17437);
or U19244 (N_19244,N_17458,N_17296);
and U19245 (N_19245,N_16858,N_16555);
and U19246 (N_19246,N_17760,N_16298);
xnor U19247 (N_19247,N_16656,N_16090);
nand U19248 (N_19248,N_17200,N_15219);
xnor U19249 (N_19249,N_15271,N_16669);
and U19250 (N_19250,N_15483,N_16223);
and U19251 (N_19251,N_17284,N_16224);
nor U19252 (N_19252,N_17266,N_16369);
nand U19253 (N_19253,N_17057,N_16915);
or U19254 (N_19254,N_15648,N_15602);
nor U19255 (N_19255,N_15654,N_17064);
and U19256 (N_19256,N_17456,N_17973);
xnor U19257 (N_19257,N_15451,N_15176);
and U19258 (N_19258,N_15813,N_17787);
or U19259 (N_19259,N_16306,N_16465);
or U19260 (N_19260,N_16868,N_17374);
nor U19261 (N_19261,N_17020,N_15775);
xor U19262 (N_19262,N_15358,N_15596);
nand U19263 (N_19263,N_15902,N_16397);
nor U19264 (N_19264,N_17821,N_17058);
xnor U19265 (N_19265,N_15162,N_15237);
or U19266 (N_19266,N_17463,N_16959);
nand U19267 (N_19267,N_16027,N_15895);
nand U19268 (N_19268,N_16988,N_15979);
and U19269 (N_19269,N_16971,N_16927);
xnor U19270 (N_19270,N_17746,N_17938);
and U19271 (N_19271,N_17038,N_17000);
or U19272 (N_19272,N_15432,N_16524);
or U19273 (N_19273,N_16194,N_16928);
or U19274 (N_19274,N_15614,N_15484);
and U19275 (N_19275,N_15839,N_16567);
nand U19276 (N_19276,N_17372,N_16638);
xnor U19277 (N_19277,N_16418,N_16791);
nor U19278 (N_19278,N_15393,N_15863);
and U19279 (N_19279,N_16982,N_16639);
nand U19280 (N_19280,N_16409,N_16573);
and U19281 (N_19281,N_15235,N_16662);
and U19282 (N_19282,N_15521,N_16891);
and U19283 (N_19283,N_17902,N_16956);
xnor U19284 (N_19284,N_17819,N_16286);
nor U19285 (N_19285,N_16437,N_17091);
nand U19286 (N_19286,N_15030,N_15469);
nand U19287 (N_19287,N_17508,N_15984);
xnor U19288 (N_19288,N_15729,N_16362);
nand U19289 (N_19289,N_17785,N_15322);
nor U19290 (N_19290,N_17987,N_15610);
or U19291 (N_19291,N_15558,N_15696);
and U19292 (N_19292,N_15941,N_17408);
and U19293 (N_19293,N_17050,N_17237);
and U19294 (N_19294,N_15597,N_16137);
xor U19295 (N_19295,N_16602,N_17313);
xnor U19296 (N_19296,N_17796,N_15448);
nor U19297 (N_19297,N_17325,N_15121);
xnor U19298 (N_19298,N_15337,N_15615);
nand U19299 (N_19299,N_16097,N_17552);
xor U19300 (N_19300,N_15797,N_17252);
and U19301 (N_19301,N_16676,N_16372);
nor U19302 (N_19302,N_17971,N_15425);
or U19303 (N_19303,N_15907,N_17158);
or U19304 (N_19304,N_17893,N_17715);
or U19305 (N_19305,N_16235,N_17339);
nand U19306 (N_19306,N_16966,N_17719);
and U19307 (N_19307,N_16990,N_16327);
and U19308 (N_19308,N_15374,N_16486);
or U19309 (N_19309,N_16412,N_17179);
nand U19310 (N_19310,N_17302,N_17052);
or U19311 (N_19311,N_17692,N_15065);
nand U19312 (N_19312,N_15588,N_15528);
nor U19313 (N_19313,N_16405,N_16862);
or U19314 (N_19314,N_17855,N_16023);
nand U19315 (N_19315,N_17133,N_15182);
or U19316 (N_19316,N_15733,N_17128);
nand U19317 (N_19317,N_17537,N_16655);
and U19318 (N_19318,N_17536,N_16271);
nor U19319 (N_19319,N_16866,N_15120);
or U19320 (N_19320,N_17705,N_15576);
nand U19321 (N_19321,N_17457,N_17764);
or U19322 (N_19322,N_15910,N_15021);
nand U19323 (N_19323,N_16042,N_16948);
or U19324 (N_19324,N_15213,N_17625);
and U19325 (N_19325,N_16174,N_16439);
nor U19326 (N_19326,N_16718,N_15195);
nand U19327 (N_19327,N_15943,N_15599);
or U19328 (N_19328,N_17042,N_15776);
nor U19329 (N_19329,N_16827,N_16080);
nand U19330 (N_19330,N_15565,N_15756);
nor U19331 (N_19331,N_17968,N_15871);
or U19332 (N_19332,N_15891,N_16776);
or U19333 (N_19333,N_17924,N_15431);
xnor U19334 (N_19334,N_17873,N_16382);
or U19335 (N_19335,N_16842,N_15068);
nand U19336 (N_19336,N_16208,N_17017);
or U19337 (N_19337,N_15909,N_15090);
nand U19338 (N_19338,N_16634,N_15101);
xor U19339 (N_19339,N_17099,N_17259);
xor U19340 (N_19340,N_15748,N_15669);
nand U19341 (N_19341,N_17619,N_17111);
and U19342 (N_19342,N_15452,N_17533);
and U19343 (N_19343,N_17083,N_17119);
or U19344 (N_19344,N_16728,N_16771);
and U19345 (N_19345,N_16071,N_17946);
xnor U19346 (N_19346,N_15466,N_16033);
nand U19347 (N_19347,N_15951,N_17316);
or U19348 (N_19348,N_15581,N_17470);
xor U19349 (N_19349,N_17383,N_16165);
nand U19350 (N_19350,N_17320,N_17668);
and U19351 (N_19351,N_15765,N_17750);
nor U19352 (N_19352,N_17805,N_16854);
xor U19353 (N_19353,N_17496,N_17406);
xor U19354 (N_19354,N_17782,N_17626);
nand U19355 (N_19355,N_15166,N_17742);
nor U19356 (N_19356,N_15888,N_15261);
nor U19357 (N_19357,N_16946,N_15353);
nor U19358 (N_19358,N_16446,N_17416);
xnor U19359 (N_19359,N_15194,N_16120);
nand U19360 (N_19360,N_16992,N_17135);
nor U19361 (N_19361,N_15222,N_16364);
and U19362 (N_19362,N_17725,N_15835);
nand U19363 (N_19363,N_17976,N_16338);
or U19364 (N_19364,N_15321,N_17175);
nor U19365 (N_19365,N_17951,N_17954);
or U19366 (N_19366,N_17620,N_15753);
xor U19367 (N_19367,N_16348,N_15010);
nand U19368 (N_19368,N_17475,N_17410);
or U19369 (N_19369,N_17419,N_16983);
and U19370 (N_19370,N_15171,N_16677);
nor U19371 (N_19371,N_16331,N_15313);
xnor U19372 (N_19372,N_17140,N_15482);
nand U19373 (N_19373,N_15424,N_17309);
xnor U19374 (N_19374,N_17554,N_16004);
xnor U19375 (N_19375,N_17205,N_17447);
nand U19376 (N_19376,N_17117,N_15997);
and U19377 (N_19377,N_17500,N_15315);
and U19378 (N_19378,N_15272,N_16145);
or U19379 (N_19379,N_17535,N_16762);
and U19380 (N_19380,N_15323,N_17945);
nand U19381 (N_19381,N_15512,N_17700);
or U19382 (N_19382,N_17474,N_16065);
xnor U19383 (N_19383,N_16324,N_16952);
xnor U19384 (N_19384,N_16312,N_17234);
or U19385 (N_19385,N_15056,N_15003);
and U19386 (N_19386,N_16903,N_16584);
or U19387 (N_19387,N_17786,N_17191);
or U19388 (N_19388,N_16148,N_17225);
nand U19389 (N_19389,N_16432,N_16929);
and U19390 (N_19390,N_15036,N_17627);
and U19391 (N_19391,N_15282,N_16407);
nor U19392 (N_19392,N_16396,N_15210);
nor U19393 (N_19393,N_17915,N_17737);
nor U19394 (N_19394,N_16079,N_17113);
xnor U19395 (N_19395,N_15757,N_17481);
xor U19396 (N_19396,N_15414,N_15281);
nor U19397 (N_19397,N_17852,N_16031);
xnor U19398 (N_19398,N_16368,N_16310);
and U19399 (N_19399,N_17667,N_16832);
nor U19400 (N_19400,N_15186,N_15627);
nor U19401 (N_19401,N_15248,N_16894);
nand U19402 (N_19402,N_17311,N_15286);
xnor U19403 (N_19403,N_16467,N_15689);
nand U19404 (N_19404,N_17726,N_16897);
xnor U19405 (N_19405,N_16898,N_15676);
xor U19406 (N_19406,N_15145,N_16443);
or U19407 (N_19407,N_17274,N_15650);
nand U19408 (N_19408,N_15953,N_15932);
or U19409 (N_19409,N_16788,N_15227);
and U19410 (N_19410,N_17759,N_16994);
nand U19411 (N_19411,N_17624,N_17258);
nor U19412 (N_19412,N_16607,N_16056);
or U19413 (N_19413,N_16739,N_15420);
xor U19414 (N_19414,N_15026,N_16592);
and U19415 (N_19415,N_15422,N_17298);
xor U19416 (N_19416,N_16264,N_16346);
or U19417 (N_19417,N_17473,N_15334);
and U19418 (N_19418,N_17034,N_16606);
xor U19419 (N_19419,N_16440,N_17792);
nand U19420 (N_19420,N_16285,N_17088);
nand U19421 (N_19421,N_15638,N_16944);
xor U19422 (N_19422,N_17603,N_15157);
nand U19423 (N_19423,N_17740,N_15197);
xor U19424 (N_19424,N_16218,N_15804);
and U19425 (N_19425,N_15795,N_16732);
and U19426 (N_19426,N_15580,N_16577);
or U19427 (N_19427,N_17054,N_16386);
or U19428 (N_19428,N_17799,N_16931);
nand U19429 (N_19429,N_16950,N_16482);
nor U19430 (N_19430,N_16815,N_16564);
xnor U19431 (N_19431,N_15463,N_16322);
or U19432 (N_19432,N_17342,N_16078);
or U19433 (N_19433,N_15973,N_15836);
and U19434 (N_19434,N_17226,N_16830);
and U19435 (N_19435,N_15336,N_15631);
xnor U19436 (N_19436,N_15981,N_15982);
xor U19437 (N_19437,N_15695,N_17955);
or U19438 (N_19438,N_16253,N_17940);
and U19439 (N_19439,N_16309,N_17155);
nand U19440 (N_19440,N_16913,N_15356);
and U19441 (N_19441,N_16106,N_17566);
nand U19442 (N_19442,N_15441,N_17674);
xnor U19443 (N_19443,N_15013,N_17464);
nand U19444 (N_19444,N_15679,N_16222);
or U19445 (N_19445,N_16053,N_17616);
or U19446 (N_19446,N_16035,N_16237);
nand U19447 (N_19447,N_15394,N_17614);
nor U19448 (N_19448,N_16841,N_17332);
nand U19449 (N_19449,N_15099,N_17528);
nand U19450 (N_19450,N_15372,N_16834);
or U19451 (N_19451,N_17775,N_15350);
nor U19452 (N_19452,N_16608,N_17176);
or U19453 (N_19453,N_15177,N_16026);
nand U19454 (N_19454,N_15494,N_17424);
and U19455 (N_19455,N_17914,N_16021);
xor U19456 (N_19456,N_17026,N_17709);
nand U19457 (N_19457,N_17434,N_16347);
nor U19458 (N_19458,N_15754,N_17917);
nor U19459 (N_19459,N_15698,N_17577);
xnor U19460 (N_19460,N_17570,N_16743);
and U19461 (N_19461,N_16907,N_16887);
nor U19462 (N_19462,N_15263,N_15684);
nand U19463 (N_19463,N_15773,N_16315);
or U19464 (N_19464,N_16674,N_16459);
and U19465 (N_19465,N_15952,N_17801);
nand U19466 (N_19466,N_15645,N_16734);
and U19467 (N_19467,N_15278,N_17632);
nor U19468 (N_19468,N_17327,N_16991);
and U19469 (N_19469,N_17858,N_17010);
or U19470 (N_19470,N_17638,N_16294);
or U19471 (N_19471,N_15126,N_15617);
nand U19472 (N_19472,N_15416,N_15942);
nand U19473 (N_19473,N_17646,N_16028);
and U19474 (N_19474,N_15751,N_15125);
nor U19475 (N_19475,N_15671,N_16527);
or U19476 (N_19476,N_16436,N_16100);
nand U19477 (N_19477,N_17729,N_17008);
xor U19478 (N_19478,N_17769,N_16978);
nor U19479 (N_19479,N_16627,N_15328);
and U19480 (N_19480,N_15132,N_17793);
nand U19481 (N_19481,N_15786,N_15523);
nor U19482 (N_19482,N_17887,N_17371);
or U19483 (N_19483,N_17660,N_15808);
or U19484 (N_19484,N_16664,N_17661);
nand U19485 (N_19485,N_16472,N_17838);
or U19486 (N_19486,N_16130,N_17250);
or U19487 (N_19487,N_16356,N_17811);
and U19488 (N_19488,N_17511,N_16186);
or U19489 (N_19489,N_15001,N_17429);
or U19490 (N_19490,N_17731,N_17904);
nor U19491 (N_19491,N_16005,N_17605);
or U19492 (N_19492,N_15541,N_17163);
nor U19493 (N_19493,N_16014,N_16726);
xor U19494 (N_19494,N_16645,N_16128);
xnor U19495 (N_19495,N_17125,N_15830);
nor U19496 (N_19496,N_15184,N_15028);
and U19497 (N_19497,N_16642,N_15601);
nand U19498 (N_19498,N_15417,N_15663);
nor U19499 (N_19499,N_15481,N_15818);
or U19500 (N_19500,N_17755,N_17273);
nand U19501 (N_19501,N_16058,N_15260);
nand U19502 (N_19502,N_17105,N_16578);
nand U19503 (N_19503,N_17462,N_17449);
nor U19504 (N_19504,N_15807,N_17410);
nand U19505 (N_19505,N_16547,N_15307);
nor U19506 (N_19506,N_16743,N_17951);
nand U19507 (N_19507,N_15996,N_15129);
or U19508 (N_19508,N_16803,N_16741);
or U19509 (N_19509,N_17313,N_15605);
nor U19510 (N_19510,N_15649,N_17076);
xnor U19511 (N_19511,N_17139,N_16648);
nand U19512 (N_19512,N_15007,N_17614);
and U19513 (N_19513,N_16535,N_16735);
or U19514 (N_19514,N_15223,N_16844);
or U19515 (N_19515,N_16751,N_16622);
nand U19516 (N_19516,N_16939,N_17422);
nand U19517 (N_19517,N_17595,N_17658);
nand U19518 (N_19518,N_15826,N_15305);
nor U19519 (N_19519,N_15219,N_16181);
nor U19520 (N_19520,N_15583,N_16928);
xor U19521 (N_19521,N_17666,N_16001);
xor U19522 (N_19522,N_17517,N_15424);
nand U19523 (N_19523,N_16260,N_17541);
nor U19524 (N_19524,N_16087,N_17750);
and U19525 (N_19525,N_16981,N_17996);
nand U19526 (N_19526,N_16270,N_15609);
xnor U19527 (N_19527,N_17060,N_17860);
nand U19528 (N_19528,N_15002,N_16804);
nor U19529 (N_19529,N_17162,N_16126);
nand U19530 (N_19530,N_16670,N_16409);
nor U19531 (N_19531,N_16911,N_17423);
or U19532 (N_19532,N_17901,N_17588);
nand U19533 (N_19533,N_16395,N_16634);
nor U19534 (N_19534,N_15628,N_17306);
nand U19535 (N_19535,N_15711,N_15355);
nor U19536 (N_19536,N_17947,N_15765);
xor U19537 (N_19537,N_16472,N_17674);
xnor U19538 (N_19538,N_16982,N_15386);
or U19539 (N_19539,N_17093,N_17990);
nor U19540 (N_19540,N_17494,N_16451);
xnor U19541 (N_19541,N_17503,N_17358);
nand U19542 (N_19542,N_16441,N_16963);
nor U19543 (N_19543,N_16789,N_17560);
or U19544 (N_19544,N_17313,N_15737);
xnor U19545 (N_19545,N_17910,N_15245);
xor U19546 (N_19546,N_16935,N_15659);
or U19547 (N_19547,N_16917,N_17905);
nand U19548 (N_19548,N_15138,N_16847);
xnor U19549 (N_19549,N_16026,N_15866);
or U19550 (N_19550,N_16172,N_17055);
and U19551 (N_19551,N_15422,N_16599);
nor U19552 (N_19552,N_16110,N_17467);
xor U19553 (N_19553,N_17995,N_16540);
and U19554 (N_19554,N_17107,N_17916);
or U19555 (N_19555,N_15425,N_15400);
nor U19556 (N_19556,N_15920,N_15508);
xor U19557 (N_19557,N_15107,N_16299);
and U19558 (N_19558,N_16972,N_17863);
nand U19559 (N_19559,N_16573,N_16073);
or U19560 (N_19560,N_15212,N_15225);
nor U19561 (N_19561,N_16823,N_16362);
or U19562 (N_19562,N_15639,N_17178);
nand U19563 (N_19563,N_16193,N_17624);
and U19564 (N_19564,N_16653,N_17786);
nand U19565 (N_19565,N_15860,N_17639);
or U19566 (N_19566,N_17408,N_16292);
xor U19567 (N_19567,N_17164,N_16901);
nand U19568 (N_19568,N_15838,N_15958);
and U19569 (N_19569,N_15548,N_15857);
nand U19570 (N_19570,N_16220,N_17101);
nand U19571 (N_19571,N_15218,N_17290);
nand U19572 (N_19572,N_15371,N_15614);
nor U19573 (N_19573,N_17759,N_15158);
nor U19574 (N_19574,N_17360,N_15908);
nand U19575 (N_19575,N_15507,N_15391);
xor U19576 (N_19576,N_17906,N_17558);
or U19577 (N_19577,N_15848,N_15686);
xor U19578 (N_19578,N_15112,N_17481);
nand U19579 (N_19579,N_15267,N_15158);
nand U19580 (N_19580,N_15018,N_16041);
or U19581 (N_19581,N_17422,N_16559);
xnor U19582 (N_19582,N_15882,N_16004);
and U19583 (N_19583,N_17602,N_16539);
and U19584 (N_19584,N_16248,N_17519);
or U19585 (N_19585,N_17070,N_17686);
and U19586 (N_19586,N_17582,N_17913);
and U19587 (N_19587,N_17020,N_17667);
and U19588 (N_19588,N_17685,N_16162);
xor U19589 (N_19589,N_17019,N_15701);
nor U19590 (N_19590,N_16544,N_15121);
nand U19591 (N_19591,N_16364,N_16771);
nand U19592 (N_19592,N_17939,N_15042);
or U19593 (N_19593,N_17540,N_15882);
nand U19594 (N_19594,N_16875,N_16200);
and U19595 (N_19595,N_16180,N_17380);
nand U19596 (N_19596,N_16105,N_15959);
nand U19597 (N_19597,N_16279,N_17365);
xnor U19598 (N_19598,N_15702,N_16992);
and U19599 (N_19599,N_17455,N_16108);
and U19600 (N_19600,N_15430,N_15864);
nor U19601 (N_19601,N_15105,N_16796);
nor U19602 (N_19602,N_16175,N_16931);
nand U19603 (N_19603,N_17424,N_16259);
or U19604 (N_19604,N_17682,N_15707);
nand U19605 (N_19605,N_15245,N_17631);
xnor U19606 (N_19606,N_17977,N_15451);
xor U19607 (N_19607,N_16243,N_15083);
and U19608 (N_19608,N_17495,N_15203);
xor U19609 (N_19609,N_17069,N_16877);
or U19610 (N_19610,N_17432,N_17548);
xor U19611 (N_19611,N_16832,N_16267);
and U19612 (N_19612,N_15268,N_17662);
xnor U19613 (N_19613,N_15709,N_15733);
and U19614 (N_19614,N_15521,N_16225);
or U19615 (N_19615,N_17311,N_17113);
or U19616 (N_19616,N_16851,N_15442);
or U19617 (N_19617,N_15829,N_15091);
nor U19618 (N_19618,N_16021,N_15293);
xnor U19619 (N_19619,N_16887,N_15201);
nand U19620 (N_19620,N_16044,N_17582);
xnor U19621 (N_19621,N_15956,N_17861);
or U19622 (N_19622,N_16674,N_17652);
and U19623 (N_19623,N_16135,N_16366);
nor U19624 (N_19624,N_15846,N_15733);
xnor U19625 (N_19625,N_17146,N_17108);
or U19626 (N_19626,N_17349,N_16414);
nand U19627 (N_19627,N_16374,N_17263);
or U19628 (N_19628,N_17512,N_15700);
xnor U19629 (N_19629,N_15315,N_16558);
xnor U19630 (N_19630,N_16802,N_15337);
and U19631 (N_19631,N_15108,N_17398);
nor U19632 (N_19632,N_16480,N_15679);
or U19633 (N_19633,N_17145,N_16590);
or U19634 (N_19634,N_17745,N_15963);
and U19635 (N_19635,N_16880,N_15913);
or U19636 (N_19636,N_16631,N_16989);
or U19637 (N_19637,N_17638,N_17356);
nor U19638 (N_19638,N_17367,N_17838);
and U19639 (N_19639,N_15024,N_16452);
nand U19640 (N_19640,N_17950,N_16301);
xor U19641 (N_19641,N_15017,N_16698);
xnor U19642 (N_19642,N_16645,N_17114);
or U19643 (N_19643,N_15995,N_16665);
and U19644 (N_19644,N_17904,N_16930);
xor U19645 (N_19645,N_17127,N_16724);
nand U19646 (N_19646,N_15749,N_15040);
xor U19647 (N_19647,N_16631,N_15647);
xnor U19648 (N_19648,N_16158,N_15533);
and U19649 (N_19649,N_17965,N_15455);
or U19650 (N_19650,N_17123,N_16016);
nor U19651 (N_19651,N_17206,N_15408);
and U19652 (N_19652,N_15750,N_17962);
nand U19653 (N_19653,N_17438,N_17338);
and U19654 (N_19654,N_15763,N_16706);
xnor U19655 (N_19655,N_15848,N_16538);
and U19656 (N_19656,N_16549,N_17517);
and U19657 (N_19657,N_17593,N_16545);
or U19658 (N_19658,N_16256,N_17544);
nand U19659 (N_19659,N_16034,N_16251);
and U19660 (N_19660,N_15305,N_15427);
xor U19661 (N_19661,N_17443,N_17378);
and U19662 (N_19662,N_15249,N_16202);
nand U19663 (N_19663,N_16909,N_15605);
xor U19664 (N_19664,N_15610,N_15339);
or U19665 (N_19665,N_15817,N_17395);
nor U19666 (N_19666,N_16211,N_16025);
xnor U19667 (N_19667,N_15146,N_17191);
or U19668 (N_19668,N_15797,N_16916);
or U19669 (N_19669,N_15097,N_15197);
nand U19670 (N_19670,N_16100,N_17300);
or U19671 (N_19671,N_17754,N_16826);
xor U19672 (N_19672,N_15628,N_16654);
and U19673 (N_19673,N_15460,N_16573);
or U19674 (N_19674,N_16952,N_15669);
and U19675 (N_19675,N_15145,N_17429);
nand U19676 (N_19676,N_17358,N_17496);
or U19677 (N_19677,N_16909,N_15698);
nand U19678 (N_19678,N_16693,N_16462);
or U19679 (N_19679,N_17879,N_17829);
nand U19680 (N_19680,N_16610,N_15472);
nand U19681 (N_19681,N_15316,N_16138);
or U19682 (N_19682,N_17929,N_15050);
or U19683 (N_19683,N_15713,N_15889);
and U19684 (N_19684,N_15284,N_15901);
or U19685 (N_19685,N_17020,N_16343);
xor U19686 (N_19686,N_17280,N_16508);
or U19687 (N_19687,N_15176,N_16692);
xnor U19688 (N_19688,N_17239,N_15656);
and U19689 (N_19689,N_17913,N_15655);
nand U19690 (N_19690,N_15822,N_16044);
or U19691 (N_19691,N_16506,N_16211);
xor U19692 (N_19692,N_15794,N_15791);
xnor U19693 (N_19693,N_17992,N_17303);
xor U19694 (N_19694,N_15225,N_17398);
or U19695 (N_19695,N_16677,N_17386);
xnor U19696 (N_19696,N_15437,N_15907);
nand U19697 (N_19697,N_15320,N_16814);
nor U19698 (N_19698,N_17918,N_17985);
nor U19699 (N_19699,N_16151,N_15321);
and U19700 (N_19700,N_15272,N_17228);
and U19701 (N_19701,N_16758,N_17839);
nor U19702 (N_19702,N_16973,N_17972);
nor U19703 (N_19703,N_17434,N_17010);
xor U19704 (N_19704,N_16585,N_17846);
or U19705 (N_19705,N_17084,N_17015);
and U19706 (N_19706,N_16608,N_15550);
and U19707 (N_19707,N_16515,N_17284);
nor U19708 (N_19708,N_17589,N_16424);
or U19709 (N_19709,N_16078,N_16877);
and U19710 (N_19710,N_17348,N_17766);
and U19711 (N_19711,N_15404,N_16034);
nor U19712 (N_19712,N_17743,N_16405);
and U19713 (N_19713,N_17004,N_17939);
and U19714 (N_19714,N_16777,N_17467);
xnor U19715 (N_19715,N_16818,N_17798);
nand U19716 (N_19716,N_16624,N_17080);
or U19717 (N_19717,N_17732,N_16275);
nand U19718 (N_19718,N_16040,N_16153);
nand U19719 (N_19719,N_16017,N_15700);
or U19720 (N_19720,N_15163,N_16741);
nand U19721 (N_19721,N_16043,N_16979);
nor U19722 (N_19722,N_17937,N_17625);
or U19723 (N_19723,N_15302,N_17981);
nor U19724 (N_19724,N_17099,N_17267);
nand U19725 (N_19725,N_17390,N_15179);
or U19726 (N_19726,N_17044,N_15893);
nor U19727 (N_19727,N_17675,N_16065);
or U19728 (N_19728,N_17164,N_17130);
xor U19729 (N_19729,N_17605,N_17566);
or U19730 (N_19730,N_17914,N_17398);
or U19731 (N_19731,N_16485,N_16206);
nand U19732 (N_19732,N_15842,N_15979);
nand U19733 (N_19733,N_17748,N_15878);
and U19734 (N_19734,N_16233,N_17337);
nand U19735 (N_19735,N_15006,N_15858);
or U19736 (N_19736,N_15558,N_16792);
and U19737 (N_19737,N_17362,N_15496);
nand U19738 (N_19738,N_15651,N_15652);
nand U19739 (N_19739,N_15460,N_15350);
xnor U19740 (N_19740,N_17892,N_17682);
or U19741 (N_19741,N_15680,N_15672);
nand U19742 (N_19742,N_16253,N_16813);
or U19743 (N_19743,N_15148,N_15753);
and U19744 (N_19744,N_17001,N_15075);
or U19745 (N_19745,N_17204,N_15760);
xor U19746 (N_19746,N_16873,N_15798);
nand U19747 (N_19747,N_15396,N_15529);
nand U19748 (N_19748,N_17001,N_15470);
nand U19749 (N_19749,N_17895,N_15253);
and U19750 (N_19750,N_16689,N_15988);
and U19751 (N_19751,N_16722,N_16870);
nand U19752 (N_19752,N_16708,N_17136);
xor U19753 (N_19753,N_15913,N_15531);
xnor U19754 (N_19754,N_17440,N_17359);
and U19755 (N_19755,N_16749,N_16798);
xor U19756 (N_19756,N_16680,N_15089);
xnor U19757 (N_19757,N_15045,N_15477);
nand U19758 (N_19758,N_15975,N_15663);
nor U19759 (N_19759,N_17859,N_16606);
nand U19760 (N_19760,N_17672,N_16653);
or U19761 (N_19761,N_15987,N_15520);
nand U19762 (N_19762,N_16187,N_17119);
or U19763 (N_19763,N_15984,N_17250);
or U19764 (N_19764,N_15607,N_15220);
or U19765 (N_19765,N_17245,N_16661);
or U19766 (N_19766,N_17473,N_17851);
or U19767 (N_19767,N_15865,N_16605);
nand U19768 (N_19768,N_15810,N_17920);
and U19769 (N_19769,N_17053,N_17860);
or U19770 (N_19770,N_17710,N_15940);
or U19771 (N_19771,N_16822,N_17845);
and U19772 (N_19772,N_15501,N_16382);
and U19773 (N_19773,N_16809,N_15393);
nor U19774 (N_19774,N_17366,N_15142);
nand U19775 (N_19775,N_17429,N_16593);
xor U19776 (N_19776,N_15062,N_16255);
or U19777 (N_19777,N_17234,N_17365);
xnor U19778 (N_19778,N_15411,N_16670);
and U19779 (N_19779,N_16128,N_17436);
nand U19780 (N_19780,N_15953,N_15533);
nor U19781 (N_19781,N_16981,N_15717);
xnor U19782 (N_19782,N_15442,N_15840);
xnor U19783 (N_19783,N_15031,N_17932);
or U19784 (N_19784,N_17384,N_17395);
or U19785 (N_19785,N_17274,N_17791);
and U19786 (N_19786,N_16811,N_15631);
nand U19787 (N_19787,N_16052,N_16944);
nor U19788 (N_19788,N_16305,N_17992);
or U19789 (N_19789,N_17342,N_15531);
nand U19790 (N_19790,N_15051,N_15474);
nor U19791 (N_19791,N_16579,N_17095);
and U19792 (N_19792,N_15042,N_17299);
and U19793 (N_19793,N_15026,N_17626);
nor U19794 (N_19794,N_15769,N_16263);
nand U19795 (N_19795,N_17225,N_17671);
xor U19796 (N_19796,N_17699,N_16254);
or U19797 (N_19797,N_17795,N_17757);
nor U19798 (N_19798,N_17277,N_15172);
nor U19799 (N_19799,N_17372,N_16556);
or U19800 (N_19800,N_15731,N_17317);
or U19801 (N_19801,N_16435,N_15444);
xnor U19802 (N_19802,N_17398,N_17154);
and U19803 (N_19803,N_16236,N_16307);
nor U19804 (N_19804,N_15185,N_17124);
and U19805 (N_19805,N_17926,N_15537);
or U19806 (N_19806,N_15792,N_17975);
nand U19807 (N_19807,N_17932,N_15046);
or U19808 (N_19808,N_17901,N_17553);
or U19809 (N_19809,N_17955,N_15073);
or U19810 (N_19810,N_16932,N_16469);
or U19811 (N_19811,N_17451,N_15567);
or U19812 (N_19812,N_16991,N_17227);
or U19813 (N_19813,N_17371,N_15149);
nor U19814 (N_19814,N_17471,N_16092);
xnor U19815 (N_19815,N_15593,N_15508);
nor U19816 (N_19816,N_15813,N_16916);
or U19817 (N_19817,N_15478,N_16437);
nor U19818 (N_19818,N_17910,N_17317);
xor U19819 (N_19819,N_16470,N_17557);
nor U19820 (N_19820,N_15730,N_17954);
nand U19821 (N_19821,N_15190,N_17475);
and U19822 (N_19822,N_15297,N_16094);
nand U19823 (N_19823,N_16770,N_15165);
nand U19824 (N_19824,N_15626,N_16765);
nand U19825 (N_19825,N_16133,N_16352);
nor U19826 (N_19826,N_16270,N_15977);
xor U19827 (N_19827,N_16660,N_16787);
or U19828 (N_19828,N_16159,N_15306);
or U19829 (N_19829,N_17093,N_16363);
and U19830 (N_19830,N_15885,N_15486);
and U19831 (N_19831,N_15985,N_16000);
and U19832 (N_19832,N_15340,N_17670);
or U19833 (N_19833,N_15759,N_17619);
and U19834 (N_19834,N_15502,N_17516);
nand U19835 (N_19835,N_16161,N_15094);
nor U19836 (N_19836,N_16202,N_16264);
or U19837 (N_19837,N_15512,N_16915);
nor U19838 (N_19838,N_17299,N_16355);
and U19839 (N_19839,N_17452,N_16274);
and U19840 (N_19840,N_15517,N_15014);
and U19841 (N_19841,N_16778,N_16448);
nor U19842 (N_19842,N_15239,N_17020);
xor U19843 (N_19843,N_17359,N_15297);
and U19844 (N_19844,N_15462,N_17093);
or U19845 (N_19845,N_15603,N_17128);
nor U19846 (N_19846,N_17049,N_15462);
nor U19847 (N_19847,N_16615,N_15250);
xor U19848 (N_19848,N_16136,N_15424);
and U19849 (N_19849,N_16877,N_15628);
and U19850 (N_19850,N_15918,N_16159);
or U19851 (N_19851,N_16190,N_17874);
nor U19852 (N_19852,N_17953,N_17992);
xor U19853 (N_19853,N_15911,N_15902);
or U19854 (N_19854,N_17600,N_16407);
or U19855 (N_19855,N_16769,N_15554);
nor U19856 (N_19856,N_16489,N_16797);
nor U19857 (N_19857,N_17910,N_16543);
nand U19858 (N_19858,N_16113,N_17495);
xor U19859 (N_19859,N_16155,N_17635);
nand U19860 (N_19860,N_15650,N_16913);
nand U19861 (N_19861,N_16803,N_15302);
nand U19862 (N_19862,N_17891,N_17715);
and U19863 (N_19863,N_15002,N_16253);
nor U19864 (N_19864,N_15675,N_15154);
nor U19865 (N_19865,N_17978,N_16574);
or U19866 (N_19866,N_15402,N_17175);
xor U19867 (N_19867,N_17011,N_15505);
or U19868 (N_19868,N_16813,N_17743);
xor U19869 (N_19869,N_15797,N_17699);
and U19870 (N_19870,N_16915,N_16868);
nand U19871 (N_19871,N_17986,N_17282);
nor U19872 (N_19872,N_17052,N_16379);
or U19873 (N_19873,N_16219,N_15337);
nor U19874 (N_19874,N_16392,N_15918);
or U19875 (N_19875,N_15523,N_16661);
and U19876 (N_19876,N_16519,N_17916);
nor U19877 (N_19877,N_17194,N_17945);
nand U19878 (N_19878,N_17713,N_15538);
xor U19879 (N_19879,N_15128,N_17104);
or U19880 (N_19880,N_15377,N_15520);
nand U19881 (N_19881,N_17489,N_15916);
and U19882 (N_19882,N_16784,N_16161);
or U19883 (N_19883,N_17409,N_15608);
and U19884 (N_19884,N_16447,N_15630);
xor U19885 (N_19885,N_15565,N_17715);
or U19886 (N_19886,N_16744,N_15243);
or U19887 (N_19887,N_16423,N_15146);
nor U19888 (N_19888,N_17986,N_15964);
or U19889 (N_19889,N_16485,N_16412);
nand U19890 (N_19890,N_17114,N_15920);
xor U19891 (N_19891,N_15115,N_16778);
xor U19892 (N_19892,N_17709,N_17595);
nor U19893 (N_19893,N_15773,N_16738);
xor U19894 (N_19894,N_15566,N_16507);
and U19895 (N_19895,N_16355,N_15198);
or U19896 (N_19896,N_17283,N_17850);
nand U19897 (N_19897,N_15835,N_16355);
nand U19898 (N_19898,N_15776,N_16854);
and U19899 (N_19899,N_16984,N_15746);
or U19900 (N_19900,N_15829,N_17717);
and U19901 (N_19901,N_15062,N_15853);
xnor U19902 (N_19902,N_15872,N_15907);
and U19903 (N_19903,N_16889,N_17828);
and U19904 (N_19904,N_16050,N_17310);
or U19905 (N_19905,N_15611,N_17423);
nand U19906 (N_19906,N_16796,N_17066);
nand U19907 (N_19907,N_17311,N_17760);
nand U19908 (N_19908,N_17388,N_17086);
and U19909 (N_19909,N_17918,N_17791);
and U19910 (N_19910,N_17232,N_15649);
nor U19911 (N_19911,N_16210,N_16396);
nand U19912 (N_19912,N_17820,N_15297);
or U19913 (N_19913,N_15459,N_17421);
and U19914 (N_19914,N_17308,N_17841);
and U19915 (N_19915,N_17520,N_15140);
nand U19916 (N_19916,N_17032,N_15818);
or U19917 (N_19917,N_17130,N_15689);
xor U19918 (N_19918,N_16823,N_15332);
xor U19919 (N_19919,N_16627,N_15162);
and U19920 (N_19920,N_16661,N_17128);
and U19921 (N_19921,N_17740,N_17615);
nand U19922 (N_19922,N_16416,N_16772);
nand U19923 (N_19923,N_17692,N_16692);
xor U19924 (N_19924,N_16923,N_16292);
and U19925 (N_19925,N_15459,N_16730);
nand U19926 (N_19926,N_15598,N_16829);
or U19927 (N_19927,N_15613,N_15258);
nand U19928 (N_19928,N_17798,N_15607);
and U19929 (N_19929,N_16289,N_15701);
nand U19930 (N_19930,N_15101,N_15458);
xnor U19931 (N_19931,N_17455,N_16844);
xnor U19932 (N_19932,N_17148,N_15964);
nand U19933 (N_19933,N_15129,N_17890);
nand U19934 (N_19934,N_17710,N_17685);
and U19935 (N_19935,N_17422,N_16094);
or U19936 (N_19936,N_15853,N_16380);
nor U19937 (N_19937,N_17282,N_17719);
and U19938 (N_19938,N_15567,N_17352);
and U19939 (N_19939,N_16294,N_16204);
nor U19940 (N_19940,N_16069,N_16864);
and U19941 (N_19941,N_16148,N_15540);
nor U19942 (N_19942,N_16292,N_17242);
or U19943 (N_19943,N_15595,N_16299);
nor U19944 (N_19944,N_15192,N_17939);
and U19945 (N_19945,N_17708,N_16801);
xor U19946 (N_19946,N_17430,N_15643);
nor U19947 (N_19947,N_15162,N_17664);
nor U19948 (N_19948,N_16330,N_17193);
nand U19949 (N_19949,N_16059,N_16017);
nor U19950 (N_19950,N_16875,N_16195);
xor U19951 (N_19951,N_17193,N_17423);
nor U19952 (N_19952,N_17682,N_16808);
xnor U19953 (N_19953,N_17843,N_15509);
xnor U19954 (N_19954,N_17649,N_15757);
and U19955 (N_19955,N_15891,N_17861);
and U19956 (N_19956,N_16427,N_15617);
and U19957 (N_19957,N_15459,N_17957);
nor U19958 (N_19958,N_17062,N_17939);
xor U19959 (N_19959,N_16937,N_16596);
xnor U19960 (N_19960,N_15996,N_17659);
nor U19961 (N_19961,N_15264,N_17143);
or U19962 (N_19962,N_15030,N_15161);
xnor U19963 (N_19963,N_15552,N_15415);
nor U19964 (N_19964,N_17658,N_15365);
or U19965 (N_19965,N_15243,N_15711);
xor U19966 (N_19966,N_16585,N_17693);
or U19967 (N_19967,N_16847,N_15149);
and U19968 (N_19968,N_15413,N_16022);
and U19969 (N_19969,N_16105,N_16290);
nor U19970 (N_19970,N_16171,N_17441);
nand U19971 (N_19971,N_16274,N_15684);
xnor U19972 (N_19972,N_17997,N_15566);
nor U19973 (N_19973,N_15661,N_17121);
or U19974 (N_19974,N_16959,N_17304);
nand U19975 (N_19975,N_16970,N_15398);
and U19976 (N_19976,N_17448,N_16137);
or U19977 (N_19977,N_16671,N_17783);
nand U19978 (N_19978,N_15647,N_15715);
nor U19979 (N_19979,N_16903,N_16280);
nor U19980 (N_19980,N_16014,N_16614);
xnor U19981 (N_19981,N_17444,N_17845);
and U19982 (N_19982,N_17913,N_17876);
or U19983 (N_19983,N_16285,N_16997);
xnor U19984 (N_19984,N_17950,N_15484);
xnor U19985 (N_19985,N_16043,N_16035);
nor U19986 (N_19986,N_16240,N_16560);
and U19987 (N_19987,N_17409,N_17945);
nor U19988 (N_19988,N_15505,N_16391);
nand U19989 (N_19989,N_16868,N_17452);
or U19990 (N_19990,N_15697,N_16096);
nor U19991 (N_19991,N_16188,N_15170);
or U19992 (N_19992,N_15673,N_15587);
or U19993 (N_19993,N_15496,N_17807);
nor U19994 (N_19994,N_16729,N_16273);
nor U19995 (N_19995,N_16544,N_17667);
nor U19996 (N_19996,N_16056,N_16066);
and U19997 (N_19997,N_15762,N_17650);
nor U19998 (N_19998,N_16937,N_15118);
or U19999 (N_19999,N_16338,N_15964);
or U20000 (N_20000,N_15715,N_16392);
nand U20001 (N_20001,N_15369,N_15034);
and U20002 (N_20002,N_17067,N_15865);
nand U20003 (N_20003,N_15880,N_15722);
xnor U20004 (N_20004,N_15803,N_15015);
nand U20005 (N_20005,N_16311,N_17783);
xor U20006 (N_20006,N_15988,N_17955);
nor U20007 (N_20007,N_17380,N_17624);
nand U20008 (N_20008,N_15491,N_15085);
and U20009 (N_20009,N_15914,N_17271);
or U20010 (N_20010,N_15019,N_15030);
and U20011 (N_20011,N_16076,N_16464);
nand U20012 (N_20012,N_17668,N_15917);
or U20013 (N_20013,N_15529,N_16381);
xnor U20014 (N_20014,N_17488,N_17881);
nand U20015 (N_20015,N_15794,N_16088);
and U20016 (N_20016,N_16149,N_17604);
or U20017 (N_20017,N_17752,N_16720);
xnor U20018 (N_20018,N_15960,N_16594);
and U20019 (N_20019,N_17960,N_15815);
nand U20020 (N_20020,N_17262,N_15309);
or U20021 (N_20021,N_15663,N_16175);
and U20022 (N_20022,N_16361,N_15213);
and U20023 (N_20023,N_17175,N_16746);
nor U20024 (N_20024,N_15271,N_16249);
and U20025 (N_20025,N_16548,N_16788);
nand U20026 (N_20026,N_16885,N_15899);
nor U20027 (N_20027,N_16018,N_17206);
or U20028 (N_20028,N_15875,N_16815);
nor U20029 (N_20029,N_16508,N_16400);
nand U20030 (N_20030,N_17535,N_16203);
nor U20031 (N_20031,N_15642,N_15754);
xnor U20032 (N_20032,N_16007,N_16803);
nor U20033 (N_20033,N_15373,N_17680);
or U20034 (N_20034,N_17016,N_15849);
xnor U20035 (N_20035,N_15422,N_16602);
xnor U20036 (N_20036,N_15151,N_17551);
xnor U20037 (N_20037,N_17682,N_15768);
nor U20038 (N_20038,N_17588,N_17438);
and U20039 (N_20039,N_16344,N_16541);
xor U20040 (N_20040,N_16880,N_17452);
xor U20041 (N_20041,N_17056,N_16141);
nor U20042 (N_20042,N_16959,N_16876);
nand U20043 (N_20043,N_17770,N_15893);
or U20044 (N_20044,N_15959,N_17309);
xor U20045 (N_20045,N_16100,N_16921);
nand U20046 (N_20046,N_16775,N_16495);
or U20047 (N_20047,N_15100,N_16875);
and U20048 (N_20048,N_15668,N_17179);
and U20049 (N_20049,N_17551,N_15216);
xnor U20050 (N_20050,N_16681,N_15533);
and U20051 (N_20051,N_16863,N_15515);
nand U20052 (N_20052,N_15340,N_16645);
nor U20053 (N_20053,N_15924,N_16570);
or U20054 (N_20054,N_15184,N_17911);
nand U20055 (N_20055,N_17104,N_16361);
and U20056 (N_20056,N_15057,N_17750);
and U20057 (N_20057,N_17811,N_16093);
and U20058 (N_20058,N_15537,N_16200);
nand U20059 (N_20059,N_17844,N_16975);
nand U20060 (N_20060,N_15691,N_16918);
nand U20061 (N_20061,N_16748,N_15292);
nand U20062 (N_20062,N_15382,N_17571);
nor U20063 (N_20063,N_15309,N_17416);
nand U20064 (N_20064,N_15636,N_17914);
xor U20065 (N_20065,N_15299,N_16663);
nor U20066 (N_20066,N_15018,N_16882);
and U20067 (N_20067,N_16594,N_15382);
or U20068 (N_20068,N_16933,N_17437);
nor U20069 (N_20069,N_15941,N_16634);
or U20070 (N_20070,N_17917,N_15305);
or U20071 (N_20071,N_16188,N_17102);
nor U20072 (N_20072,N_16831,N_17898);
and U20073 (N_20073,N_16983,N_17898);
xor U20074 (N_20074,N_16093,N_17349);
nor U20075 (N_20075,N_15199,N_17136);
and U20076 (N_20076,N_16256,N_17210);
nand U20077 (N_20077,N_17838,N_15016);
or U20078 (N_20078,N_15891,N_16936);
nor U20079 (N_20079,N_15681,N_15277);
nor U20080 (N_20080,N_15544,N_16479);
and U20081 (N_20081,N_15131,N_16113);
nand U20082 (N_20082,N_17020,N_16372);
or U20083 (N_20083,N_16372,N_15841);
xnor U20084 (N_20084,N_16310,N_15968);
and U20085 (N_20085,N_16949,N_17935);
nand U20086 (N_20086,N_17622,N_16425);
or U20087 (N_20087,N_15617,N_15571);
or U20088 (N_20088,N_17870,N_17321);
or U20089 (N_20089,N_17804,N_16765);
and U20090 (N_20090,N_15746,N_17686);
or U20091 (N_20091,N_15051,N_16681);
nor U20092 (N_20092,N_15699,N_15865);
nor U20093 (N_20093,N_16950,N_17117);
and U20094 (N_20094,N_17829,N_17885);
and U20095 (N_20095,N_15584,N_16650);
and U20096 (N_20096,N_16408,N_17536);
nor U20097 (N_20097,N_16238,N_15616);
nor U20098 (N_20098,N_17556,N_15253);
and U20099 (N_20099,N_15807,N_17865);
nand U20100 (N_20100,N_16319,N_15862);
or U20101 (N_20101,N_16997,N_15290);
xor U20102 (N_20102,N_16636,N_16117);
nor U20103 (N_20103,N_15193,N_17545);
nor U20104 (N_20104,N_17192,N_16025);
or U20105 (N_20105,N_15552,N_15078);
xor U20106 (N_20106,N_15021,N_17384);
nor U20107 (N_20107,N_16057,N_17155);
xor U20108 (N_20108,N_15110,N_17061);
nand U20109 (N_20109,N_15823,N_15921);
xnor U20110 (N_20110,N_15584,N_16942);
nor U20111 (N_20111,N_15299,N_17610);
nor U20112 (N_20112,N_16139,N_16613);
xnor U20113 (N_20113,N_16047,N_16862);
nand U20114 (N_20114,N_17528,N_15179);
xor U20115 (N_20115,N_16120,N_17776);
and U20116 (N_20116,N_15401,N_17426);
xnor U20117 (N_20117,N_17089,N_15014);
or U20118 (N_20118,N_15143,N_17903);
and U20119 (N_20119,N_16412,N_15360);
or U20120 (N_20120,N_16646,N_16273);
xnor U20121 (N_20121,N_15148,N_16398);
and U20122 (N_20122,N_16432,N_17246);
and U20123 (N_20123,N_17952,N_17726);
or U20124 (N_20124,N_16289,N_17326);
and U20125 (N_20125,N_15977,N_17303);
nand U20126 (N_20126,N_16821,N_16219);
nor U20127 (N_20127,N_17942,N_15863);
nand U20128 (N_20128,N_17122,N_17312);
xor U20129 (N_20129,N_16712,N_16648);
nand U20130 (N_20130,N_15550,N_16551);
nor U20131 (N_20131,N_15915,N_15963);
nor U20132 (N_20132,N_15995,N_16428);
nor U20133 (N_20133,N_17930,N_16559);
or U20134 (N_20134,N_17569,N_16566);
nand U20135 (N_20135,N_16000,N_16960);
nand U20136 (N_20136,N_15564,N_15514);
nand U20137 (N_20137,N_17454,N_15076);
nor U20138 (N_20138,N_15970,N_16581);
nor U20139 (N_20139,N_15965,N_15558);
or U20140 (N_20140,N_17566,N_17465);
nor U20141 (N_20141,N_16004,N_15150);
xnor U20142 (N_20142,N_17126,N_16471);
xnor U20143 (N_20143,N_15819,N_16206);
nor U20144 (N_20144,N_17653,N_16374);
and U20145 (N_20145,N_17510,N_16089);
or U20146 (N_20146,N_16951,N_15088);
or U20147 (N_20147,N_16345,N_16618);
or U20148 (N_20148,N_15857,N_17032);
nor U20149 (N_20149,N_17954,N_16685);
xor U20150 (N_20150,N_17633,N_17270);
or U20151 (N_20151,N_16261,N_17381);
nor U20152 (N_20152,N_17745,N_16222);
nand U20153 (N_20153,N_16438,N_15241);
xor U20154 (N_20154,N_15636,N_16208);
and U20155 (N_20155,N_15352,N_17951);
or U20156 (N_20156,N_15745,N_15413);
nand U20157 (N_20157,N_15083,N_16339);
nand U20158 (N_20158,N_16519,N_17340);
nor U20159 (N_20159,N_16176,N_16716);
nand U20160 (N_20160,N_15136,N_15961);
nor U20161 (N_20161,N_17410,N_17173);
nor U20162 (N_20162,N_16263,N_17761);
nand U20163 (N_20163,N_15717,N_15928);
or U20164 (N_20164,N_15275,N_15457);
or U20165 (N_20165,N_15717,N_16968);
nand U20166 (N_20166,N_16741,N_15194);
nor U20167 (N_20167,N_16363,N_16928);
xnor U20168 (N_20168,N_16070,N_17104);
xor U20169 (N_20169,N_17740,N_16554);
nor U20170 (N_20170,N_15857,N_17527);
nor U20171 (N_20171,N_15150,N_15020);
nor U20172 (N_20172,N_15165,N_16871);
and U20173 (N_20173,N_17074,N_17040);
xnor U20174 (N_20174,N_17339,N_16622);
or U20175 (N_20175,N_17844,N_16724);
nor U20176 (N_20176,N_16955,N_17254);
nand U20177 (N_20177,N_15033,N_17085);
nor U20178 (N_20178,N_16808,N_15842);
or U20179 (N_20179,N_17156,N_15784);
and U20180 (N_20180,N_16655,N_17452);
or U20181 (N_20181,N_17776,N_17101);
xnor U20182 (N_20182,N_17895,N_17333);
xor U20183 (N_20183,N_17122,N_17242);
nand U20184 (N_20184,N_17284,N_15504);
or U20185 (N_20185,N_15011,N_17494);
and U20186 (N_20186,N_17741,N_17067);
nand U20187 (N_20187,N_17059,N_15212);
nand U20188 (N_20188,N_15977,N_17107);
nand U20189 (N_20189,N_16778,N_15431);
nor U20190 (N_20190,N_16583,N_15492);
nor U20191 (N_20191,N_15299,N_15194);
xnor U20192 (N_20192,N_16672,N_17879);
nor U20193 (N_20193,N_15766,N_15584);
xor U20194 (N_20194,N_15581,N_15015);
nand U20195 (N_20195,N_15001,N_15788);
nand U20196 (N_20196,N_16930,N_17960);
nor U20197 (N_20197,N_17343,N_17353);
xor U20198 (N_20198,N_17137,N_15649);
xor U20199 (N_20199,N_16372,N_15839);
and U20200 (N_20200,N_16435,N_15227);
xor U20201 (N_20201,N_16118,N_16102);
nand U20202 (N_20202,N_15397,N_16802);
and U20203 (N_20203,N_15429,N_16939);
nor U20204 (N_20204,N_15062,N_15469);
nand U20205 (N_20205,N_16960,N_17720);
or U20206 (N_20206,N_16013,N_17266);
or U20207 (N_20207,N_15793,N_16353);
and U20208 (N_20208,N_17317,N_16585);
xor U20209 (N_20209,N_17080,N_15476);
and U20210 (N_20210,N_15301,N_15582);
or U20211 (N_20211,N_17920,N_17111);
nor U20212 (N_20212,N_17802,N_15518);
xor U20213 (N_20213,N_16570,N_17173);
and U20214 (N_20214,N_16473,N_17805);
nand U20215 (N_20215,N_16052,N_15843);
nor U20216 (N_20216,N_15841,N_16381);
or U20217 (N_20217,N_16673,N_15878);
nor U20218 (N_20218,N_17522,N_15147);
nor U20219 (N_20219,N_17584,N_15149);
nor U20220 (N_20220,N_17657,N_15568);
and U20221 (N_20221,N_16332,N_17658);
xnor U20222 (N_20222,N_15622,N_16930);
nor U20223 (N_20223,N_15457,N_16325);
or U20224 (N_20224,N_15870,N_15415);
nand U20225 (N_20225,N_16946,N_15203);
xnor U20226 (N_20226,N_17015,N_15198);
nor U20227 (N_20227,N_15467,N_16322);
xnor U20228 (N_20228,N_16368,N_17468);
xnor U20229 (N_20229,N_16289,N_17379);
nor U20230 (N_20230,N_17886,N_15564);
and U20231 (N_20231,N_17976,N_15802);
nand U20232 (N_20232,N_16313,N_16766);
xnor U20233 (N_20233,N_16274,N_15969);
nand U20234 (N_20234,N_16168,N_17810);
xnor U20235 (N_20235,N_16598,N_16488);
nor U20236 (N_20236,N_15135,N_17266);
or U20237 (N_20237,N_17044,N_15608);
or U20238 (N_20238,N_15562,N_15588);
or U20239 (N_20239,N_16169,N_17477);
nand U20240 (N_20240,N_15858,N_15021);
nor U20241 (N_20241,N_17008,N_15991);
and U20242 (N_20242,N_15166,N_15576);
xnor U20243 (N_20243,N_16660,N_16079);
or U20244 (N_20244,N_15294,N_17042);
and U20245 (N_20245,N_15238,N_16758);
nor U20246 (N_20246,N_15141,N_15688);
nand U20247 (N_20247,N_15069,N_17230);
nand U20248 (N_20248,N_17963,N_17849);
or U20249 (N_20249,N_17069,N_17723);
nand U20250 (N_20250,N_15813,N_16210);
xnor U20251 (N_20251,N_17896,N_17157);
or U20252 (N_20252,N_16792,N_17197);
xor U20253 (N_20253,N_17362,N_16702);
nand U20254 (N_20254,N_16592,N_16034);
xor U20255 (N_20255,N_15256,N_15470);
or U20256 (N_20256,N_16309,N_17399);
nor U20257 (N_20257,N_15153,N_16358);
nor U20258 (N_20258,N_17020,N_17802);
or U20259 (N_20259,N_15111,N_16914);
or U20260 (N_20260,N_15056,N_15219);
xnor U20261 (N_20261,N_17829,N_17781);
or U20262 (N_20262,N_17999,N_17709);
and U20263 (N_20263,N_15230,N_17637);
or U20264 (N_20264,N_15640,N_16234);
and U20265 (N_20265,N_16265,N_15541);
nor U20266 (N_20266,N_15364,N_16452);
and U20267 (N_20267,N_16874,N_16602);
or U20268 (N_20268,N_15941,N_15768);
nand U20269 (N_20269,N_15138,N_15014);
xor U20270 (N_20270,N_15735,N_16507);
and U20271 (N_20271,N_16627,N_17134);
nand U20272 (N_20272,N_15059,N_16495);
and U20273 (N_20273,N_15949,N_16536);
and U20274 (N_20274,N_17755,N_16230);
and U20275 (N_20275,N_16446,N_17726);
nand U20276 (N_20276,N_15616,N_15906);
or U20277 (N_20277,N_17594,N_15768);
nand U20278 (N_20278,N_16653,N_16143);
and U20279 (N_20279,N_17606,N_15076);
and U20280 (N_20280,N_16991,N_16558);
nor U20281 (N_20281,N_17423,N_15780);
nand U20282 (N_20282,N_16602,N_15437);
and U20283 (N_20283,N_15619,N_15972);
and U20284 (N_20284,N_17019,N_17412);
or U20285 (N_20285,N_16728,N_15680);
nand U20286 (N_20286,N_16309,N_17430);
or U20287 (N_20287,N_17894,N_15568);
nor U20288 (N_20288,N_16732,N_16077);
nor U20289 (N_20289,N_15104,N_15478);
nor U20290 (N_20290,N_16047,N_16612);
nand U20291 (N_20291,N_17628,N_17877);
and U20292 (N_20292,N_15002,N_17434);
or U20293 (N_20293,N_16291,N_15254);
nor U20294 (N_20294,N_15167,N_15521);
or U20295 (N_20295,N_17685,N_16331);
and U20296 (N_20296,N_15222,N_16897);
nand U20297 (N_20297,N_15231,N_17911);
or U20298 (N_20298,N_15703,N_15871);
nor U20299 (N_20299,N_16176,N_16484);
or U20300 (N_20300,N_16440,N_17764);
and U20301 (N_20301,N_17493,N_15308);
xor U20302 (N_20302,N_17963,N_16647);
xor U20303 (N_20303,N_16273,N_17789);
and U20304 (N_20304,N_16789,N_16647);
and U20305 (N_20305,N_17615,N_16704);
nor U20306 (N_20306,N_16359,N_16287);
xnor U20307 (N_20307,N_17274,N_15005);
xnor U20308 (N_20308,N_15825,N_17120);
nand U20309 (N_20309,N_16017,N_15697);
nor U20310 (N_20310,N_16110,N_16124);
and U20311 (N_20311,N_15193,N_16770);
nand U20312 (N_20312,N_17093,N_16073);
nand U20313 (N_20313,N_17759,N_17174);
nor U20314 (N_20314,N_16715,N_17111);
nand U20315 (N_20315,N_17012,N_15408);
nor U20316 (N_20316,N_15568,N_16346);
and U20317 (N_20317,N_15911,N_17770);
or U20318 (N_20318,N_17244,N_15940);
and U20319 (N_20319,N_15774,N_16181);
or U20320 (N_20320,N_16690,N_16309);
xor U20321 (N_20321,N_16741,N_15620);
nand U20322 (N_20322,N_16473,N_17314);
xnor U20323 (N_20323,N_17461,N_16023);
or U20324 (N_20324,N_16176,N_15573);
or U20325 (N_20325,N_16147,N_16672);
and U20326 (N_20326,N_16861,N_16819);
or U20327 (N_20327,N_15750,N_16617);
xor U20328 (N_20328,N_16859,N_15488);
and U20329 (N_20329,N_15751,N_17046);
nor U20330 (N_20330,N_15463,N_16232);
xnor U20331 (N_20331,N_15436,N_16623);
nand U20332 (N_20332,N_15577,N_17564);
and U20333 (N_20333,N_16264,N_16645);
and U20334 (N_20334,N_17612,N_16483);
xnor U20335 (N_20335,N_17626,N_17073);
or U20336 (N_20336,N_17217,N_17429);
nor U20337 (N_20337,N_17107,N_15724);
nor U20338 (N_20338,N_17087,N_16927);
xor U20339 (N_20339,N_17222,N_16110);
nand U20340 (N_20340,N_17248,N_16136);
nand U20341 (N_20341,N_17194,N_16640);
or U20342 (N_20342,N_15079,N_15118);
and U20343 (N_20343,N_17181,N_16213);
nand U20344 (N_20344,N_17242,N_17197);
or U20345 (N_20345,N_17610,N_16613);
or U20346 (N_20346,N_17852,N_16235);
nand U20347 (N_20347,N_15980,N_17829);
xor U20348 (N_20348,N_15181,N_16131);
nor U20349 (N_20349,N_16030,N_17431);
xor U20350 (N_20350,N_16572,N_17099);
nor U20351 (N_20351,N_17805,N_16880);
and U20352 (N_20352,N_17701,N_17419);
xor U20353 (N_20353,N_16251,N_17678);
xnor U20354 (N_20354,N_16974,N_17007);
nand U20355 (N_20355,N_15031,N_15118);
or U20356 (N_20356,N_16808,N_15736);
or U20357 (N_20357,N_17974,N_17963);
xor U20358 (N_20358,N_16727,N_15090);
nand U20359 (N_20359,N_16913,N_15017);
or U20360 (N_20360,N_17482,N_16025);
and U20361 (N_20361,N_15497,N_15597);
nor U20362 (N_20362,N_16779,N_17237);
and U20363 (N_20363,N_17034,N_16984);
nor U20364 (N_20364,N_17663,N_17344);
nor U20365 (N_20365,N_17597,N_17106);
or U20366 (N_20366,N_16808,N_17959);
nand U20367 (N_20367,N_15355,N_15968);
nand U20368 (N_20368,N_16813,N_15759);
xnor U20369 (N_20369,N_15075,N_16503);
xnor U20370 (N_20370,N_16669,N_16523);
or U20371 (N_20371,N_15901,N_15960);
xnor U20372 (N_20372,N_16404,N_15868);
nor U20373 (N_20373,N_16321,N_16099);
nor U20374 (N_20374,N_16137,N_15591);
nand U20375 (N_20375,N_17226,N_16893);
and U20376 (N_20376,N_15829,N_16519);
nand U20377 (N_20377,N_15721,N_15417);
or U20378 (N_20378,N_17559,N_16508);
and U20379 (N_20379,N_16612,N_16964);
or U20380 (N_20380,N_15431,N_15504);
and U20381 (N_20381,N_15504,N_16605);
xor U20382 (N_20382,N_17634,N_15499);
nand U20383 (N_20383,N_17163,N_15097);
nor U20384 (N_20384,N_16617,N_15330);
and U20385 (N_20385,N_17657,N_15327);
and U20386 (N_20386,N_16521,N_17919);
xnor U20387 (N_20387,N_16630,N_16070);
xnor U20388 (N_20388,N_15241,N_16510);
or U20389 (N_20389,N_15956,N_16223);
and U20390 (N_20390,N_17432,N_16519);
and U20391 (N_20391,N_16118,N_15925);
or U20392 (N_20392,N_16600,N_15324);
and U20393 (N_20393,N_17572,N_15194);
nor U20394 (N_20394,N_16835,N_15684);
nor U20395 (N_20395,N_15034,N_16186);
and U20396 (N_20396,N_15892,N_15457);
xor U20397 (N_20397,N_15706,N_15031);
and U20398 (N_20398,N_15179,N_17913);
and U20399 (N_20399,N_15189,N_16751);
xnor U20400 (N_20400,N_16811,N_16338);
or U20401 (N_20401,N_15704,N_16207);
xor U20402 (N_20402,N_15733,N_16115);
nor U20403 (N_20403,N_16002,N_17979);
or U20404 (N_20404,N_16502,N_17188);
xnor U20405 (N_20405,N_15801,N_17444);
xor U20406 (N_20406,N_16481,N_17340);
and U20407 (N_20407,N_17384,N_17656);
and U20408 (N_20408,N_15915,N_15441);
and U20409 (N_20409,N_17083,N_15743);
nor U20410 (N_20410,N_17221,N_17540);
nor U20411 (N_20411,N_16895,N_15506);
or U20412 (N_20412,N_15873,N_16922);
nor U20413 (N_20413,N_16396,N_16037);
or U20414 (N_20414,N_16146,N_16974);
xor U20415 (N_20415,N_15132,N_16693);
nor U20416 (N_20416,N_15987,N_16852);
xor U20417 (N_20417,N_15880,N_15980);
or U20418 (N_20418,N_17573,N_17731);
and U20419 (N_20419,N_15867,N_17715);
nor U20420 (N_20420,N_16696,N_15755);
and U20421 (N_20421,N_15331,N_16950);
or U20422 (N_20422,N_17135,N_17258);
nand U20423 (N_20423,N_15291,N_15779);
and U20424 (N_20424,N_17518,N_15038);
and U20425 (N_20425,N_16071,N_15474);
or U20426 (N_20426,N_17029,N_16429);
and U20427 (N_20427,N_15181,N_17279);
xor U20428 (N_20428,N_16727,N_16611);
and U20429 (N_20429,N_17102,N_16743);
and U20430 (N_20430,N_17844,N_16334);
and U20431 (N_20431,N_16372,N_17619);
nand U20432 (N_20432,N_16941,N_15213);
and U20433 (N_20433,N_16581,N_16770);
or U20434 (N_20434,N_16715,N_17896);
nor U20435 (N_20435,N_15287,N_15066);
or U20436 (N_20436,N_16611,N_16448);
nand U20437 (N_20437,N_17430,N_17063);
and U20438 (N_20438,N_16200,N_17923);
and U20439 (N_20439,N_17654,N_17671);
xor U20440 (N_20440,N_17680,N_17066);
and U20441 (N_20441,N_17322,N_15800);
xor U20442 (N_20442,N_15943,N_15722);
xor U20443 (N_20443,N_17048,N_15745);
or U20444 (N_20444,N_16150,N_17082);
nor U20445 (N_20445,N_16382,N_16054);
nand U20446 (N_20446,N_16659,N_17807);
nor U20447 (N_20447,N_17176,N_15254);
nor U20448 (N_20448,N_17088,N_17653);
or U20449 (N_20449,N_17373,N_17923);
or U20450 (N_20450,N_15616,N_17285);
nand U20451 (N_20451,N_15260,N_17362);
or U20452 (N_20452,N_15128,N_17551);
nor U20453 (N_20453,N_16280,N_17772);
nor U20454 (N_20454,N_15833,N_17507);
and U20455 (N_20455,N_17748,N_15846);
or U20456 (N_20456,N_16906,N_17174);
or U20457 (N_20457,N_16208,N_17153);
nor U20458 (N_20458,N_15362,N_16975);
nor U20459 (N_20459,N_17127,N_15325);
and U20460 (N_20460,N_16114,N_16934);
xnor U20461 (N_20461,N_15511,N_15410);
nand U20462 (N_20462,N_15950,N_15530);
nor U20463 (N_20463,N_16104,N_15833);
xnor U20464 (N_20464,N_16089,N_16935);
nor U20465 (N_20465,N_15873,N_16247);
nand U20466 (N_20466,N_15005,N_15638);
nand U20467 (N_20467,N_15572,N_15874);
nand U20468 (N_20468,N_16233,N_16012);
xor U20469 (N_20469,N_15427,N_16920);
or U20470 (N_20470,N_17875,N_15820);
xor U20471 (N_20471,N_15431,N_15286);
xor U20472 (N_20472,N_15558,N_15487);
or U20473 (N_20473,N_16482,N_16048);
nor U20474 (N_20474,N_15408,N_16827);
nor U20475 (N_20475,N_17580,N_15047);
nand U20476 (N_20476,N_16451,N_17137);
or U20477 (N_20477,N_15090,N_15781);
xor U20478 (N_20478,N_16882,N_15026);
nand U20479 (N_20479,N_16304,N_15598);
nand U20480 (N_20480,N_17574,N_15088);
or U20481 (N_20481,N_15401,N_15233);
or U20482 (N_20482,N_15618,N_15191);
and U20483 (N_20483,N_15377,N_16112);
nand U20484 (N_20484,N_16638,N_17439);
xnor U20485 (N_20485,N_15944,N_15524);
xor U20486 (N_20486,N_15353,N_15514);
nor U20487 (N_20487,N_16832,N_17686);
or U20488 (N_20488,N_17371,N_16957);
nand U20489 (N_20489,N_15614,N_17245);
and U20490 (N_20490,N_17567,N_15287);
nand U20491 (N_20491,N_17727,N_15083);
or U20492 (N_20492,N_15158,N_15107);
nand U20493 (N_20493,N_16522,N_15982);
nand U20494 (N_20494,N_15751,N_16574);
nand U20495 (N_20495,N_15629,N_16949);
or U20496 (N_20496,N_15392,N_16995);
nand U20497 (N_20497,N_17050,N_16352);
nor U20498 (N_20498,N_17188,N_16976);
nor U20499 (N_20499,N_16742,N_17262);
and U20500 (N_20500,N_17601,N_17313);
nand U20501 (N_20501,N_15398,N_16628);
or U20502 (N_20502,N_16657,N_15788);
nand U20503 (N_20503,N_17010,N_15796);
or U20504 (N_20504,N_15694,N_16785);
xor U20505 (N_20505,N_15299,N_17317);
and U20506 (N_20506,N_17642,N_16296);
nor U20507 (N_20507,N_15523,N_17442);
and U20508 (N_20508,N_17534,N_15592);
nand U20509 (N_20509,N_15617,N_16541);
nand U20510 (N_20510,N_15329,N_17861);
nand U20511 (N_20511,N_16139,N_16080);
or U20512 (N_20512,N_16725,N_16213);
nand U20513 (N_20513,N_15838,N_15333);
xor U20514 (N_20514,N_15502,N_15910);
xnor U20515 (N_20515,N_17851,N_17668);
and U20516 (N_20516,N_15386,N_16729);
nor U20517 (N_20517,N_16428,N_17315);
nand U20518 (N_20518,N_15084,N_16611);
xor U20519 (N_20519,N_16195,N_16352);
nor U20520 (N_20520,N_17142,N_15424);
or U20521 (N_20521,N_17793,N_15838);
or U20522 (N_20522,N_16035,N_16450);
or U20523 (N_20523,N_17279,N_17834);
nand U20524 (N_20524,N_17250,N_15094);
and U20525 (N_20525,N_17975,N_15928);
or U20526 (N_20526,N_17546,N_17686);
and U20527 (N_20527,N_17876,N_17861);
and U20528 (N_20528,N_17338,N_15194);
and U20529 (N_20529,N_16525,N_15698);
nand U20530 (N_20530,N_17846,N_15865);
and U20531 (N_20531,N_16166,N_16358);
nand U20532 (N_20532,N_17665,N_17233);
nand U20533 (N_20533,N_17961,N_17061);
nand U20534 (N_20534,N_17412,N_15264);
nand U20535 (N_20535,N_16000,N_16081);
nor U20536 (N_20536,N_17518,N_15722);
or U20537 (N_20537,N_15231,N_15764);
or U20538 (N_20538,N_15239,N_15515);
and U20539 (N_20539,N_17100,N_17345);
nor U20540 (N_20540,N_16061,N_15354);
nor U20541 (N_20541,N_17760,N_16943);
xor U20542 (N_20542,N_16009,N_17452);
or U20543 (N_20543,N_15970,N_15264);
or U20544 (N_20544,N_17536,N_16022);
nand U20545 (N_20545,N_17716,N_17617);
xnor U20546 (N_20546,N_15657,N_16930);
and U20547 (N_20547,N_15609,N_15329);
and U20548 (N_20548,N_17925,N_17995);
xnor U20549 (N_20549,N_16596,N_15965);
xor U20550 (N_20550,N_15063,N_16541);
nor U20551 (N_20551,N_16709,N_16160);
nand U20552 (N_20552,N_17923,N_17219);
nand U20553 (N_20553,N_15780,N_17203);
or U20554 (N_20554,N_17498,N_17732);
nand U20555 (N_20555,N_17355,N_16922);
or U20556 (N_20556,N_16371,N_15335);
nand U20557 (N_20557,N_17171,N_17374);
nand U20558 (N_20558,N_15621,N_15702);
nand U20559 (N_20559,N_16881,N_17337);
and U20560 (N_20560,N_15953,N_15792);
or U20561 (N_20561,N_15122,N_16219);
nand U20562 (N_20562,N_16807,N_15335);
nand U20563 (N_20563,N_17012,N_17828);
xnor U20564 (N_20564,N_17640,N_16716);
xor U20565 (N_20565,N_15544,N_17152);
and U20566 (N_20566,N_15705,N_16688);
and U20567 (N_20567,N_15476,N_17343);
nor U20568 (N_20568,N_17726,N_17094);
and U20569 (N_20569,N_17621,N_17172);
nand U20570 (N_20570,N_17367,N_17033);
or U20571 (N_20571,N_15901,N_15620);
and U20572 (N_20572,N_15989,N_15454);
or U20573 (N_20573,N_16241,N_15863);
or U20574 (N_20574,N_15723,N_15260);
nor U20575 (N_20575,N_15167,N_15573);
xor U20576 (N_20576,N_16966,N_16764);
and U20577 (N_20577,N_17621,N_16181);
xor U20578 (N_20578,N_17681,N_15203);
or U20579 (N_20579,N_15482,N_17221);
nor U20580 (N_20580,N_17488,N_16411);
and U20581 (N_20581,N_17849,N_17728);
and U20582 (N_20582,N_15701,N_16487);
nand U20583 (N_20583,N_15007,N_17313);
nand U20584 (N_20584,N_17294,N_15145);
nand U20585 (N_20585,N_16464,N_15168);
xnor U20586 (N_20586,N_15626,N_16758);
nor U20587 (N_20587,N_17829,N_15223);
and U20588 (N_20588,N_16433,N_17499);
nor U20589 (N_20589,N_17241,N_17389);
xor U20590 (N_20590,N_17900,N_16866);
and U20591 (N_20591,N_17656,N_16886);
or U20592 (N_20592,N_17491,N_15730);
and U20593 (N_20593,N_17465,N_17881);
nand U20594 (N_20594,N_17238,N_15163);
or U20595 (N_20595,N_15182,N_16344);
and U20596 (N_20596,N_17036,N_17708);
nand U20597 (N_20597,N_17519,N_17429);
and U20598 (N_20598,N_17758,N_17369);
nor U20599 (N_20599,N_17004,N_17408);
or U20600 (N_20600,N_16502,N_17812);
nand U20601 (N_20601,N_17906,N_15170);
or U20602 (N_20602,N_16921,N_17603);
or U20603 (N_20603,N_17488,N_17714);
nor U20604 (N_20604,N_15049,N_17954);
xnor U20605 (N_20605,N_16431,N_16339);
and U20606 (N_20606,N_17371,N_17188);
and U20607 (N_20607,N_17355,N_16391);
or U20608 (N_20608,N_16527,N_15601);
xnor U20609 (N_20609,N_15079,N_17749);
or U20610 (N_20610,N_15838,N_16569);
nand U20611 (N_20611,N_15393,N_17251);
or U20612 (N_20612,N_15248,N_17624);
nor U20613 (N_20613,N_15159,N_17970);
and U20614 (N_20614,N_17831,N_15801);
xor U20615 (N_20615,N_15841,N_17866);
xnor U20616 (N_20616,N_15907,N_15017);
nand U20617 (N_20617,N_17556,N_16675);
or U20618 (N_20618,N_17355,N_16304);
xnor U20619 (N_20619,N_15611,N_16444);
nor U20620 (N_20620,N_16932,N_16117);
or U20621 (N_20621,N_16076,N_17152);
and U20622 (N_20622,N_15636,N_17429);
nor U20623 (N_20623,N_16731,N_16171);
nand U20624 (N_20624,N_17492,N_15339);
and U20625 (N_20625,N_16270,N_15962);
or U20626 (N_20626,N_17168,N_17979);
or U20627 (N_20627,N_16715,N_17227);
or U20628 (N_20628,N_15997,N_16283);
or U20629 (N_20629,N_15632,N_15835);
nand U20630 (N_20630,N_17925,N_17376);
xor U20631 (N_20631,N_15746,N_17892);
nor U20632 (N_20632,N_15433,N_17350);
and U20633 (N_20633,N_16059,N_17221);
or U20634 (N_20634,N_17709,N_16026);
nand U20635 (N_20635,N_15464,N_17668);
nor U20636 (N_20636,N_15368,N_15812);
xnor U20637 (N_20637,N_16894,N_17127);
and U20638 (N_20638,N_16697,N_15843);
or U20639 (N_20639,N_17866,N_15308);
xnor U20640 (N_20640,N_15059,N_16423);
nand U20641 (N_20641,N_15831,N_17329);
and U20642 (N_20642,N_17721,N_15769);
or U20643 (N_20643,N_15312,N_15845);
xor U20644 (N_20644,N_17087,N_15509);
xor U20645 (N_20645,N_17200,N_16762);
xor U20646 (N_20646,N_16806,N_16001);
nand U20647 (N_20647,N_17846,N_16668);
nand U20648 (N_20648,N_16784,N_17498);
xor U20649 (N_20649,N_17570,N_17126);
nand U20650 (N_20650,N_17802,N_17518);
nor U20651 (N_20651,N_17413,N_15784);
xor U20652 (N_20652,N_17738,N_17664);
nor U20653 (N_20653,N_17529,N_17623);
nor U20654 (N_20654,N_16673,N_16936);
and U20655 (N_20655,N_15523,N_15252);
xnor U20656 (N_20656,N_16541,N_15641);
nand U20657 (N_20657,N_16103,N_15873);
or U20658 (N_20658,N_15576,N_16523);
xnor U20659 (N_20659,N_15821,N_15562);
or U20660 (N_20660,N_16895,N_17772);
xor U20661 (N_20661,N_15326,N_16305);
xnor U20662 (N_20662,N_16630,N_15267);
xnor U20663 (N_20663,N_16000,N_15853);
nor U20664 (N_20664,N_16946,N_16238);
or U20665 (N_20665,N_15861,N_16836);
or U20666 (N_20666,N_16259,N_16930);
nand U20667 (N_20667,N_15900,N_17327);
or U20668 (N_20668,N_16371,N_16694);
xor U20669 (N_20669,N_17478,N_15832);
or U20670 (N_20670,N_16557,N_16608);
xnor U20671 (N_20671,N_17669,N_15968);
nor U20672 (N_20672,N_15657,N_17846);
or U20673 (N_20673,N_17856,N_15740);
or U20674 (N_20674,N_15193,N_16080);
nor U20675 (N_20675,N_17930,N_17265);
and U20676 (N_20676,N_15446,N_17278);
nand U20677 (N_20677,N_15584,N_17978);
or U20678 (N_20678,N_17233,N_16374);
nor U20679 (N_20679,N_15884,N_16124);
or U20680 (N_20680,N_15480,N_15692);
nand U20681 (N_20681,N_16918,N_17303);
or U20682 (N_20682,N_17962,N_17538);
and U20683 (N_20683,N_15210,N_15200);
xor U20684 (N_20684,N_16543,N_17879);
and U20685 (N_20685,N_15108,N_17302);
nand U20686 (N_20686,N_16027,N_16028);
and U20687 (N_20687,N_15398,N_16440);
and U20688 (N_20688,N_17168,N_16580);
and U20689 (N_20689,N_15538,N_15829);
or U20690 (N_20690,N_17262,N_15479);
xnor U20691 (N_20691,N_16804,N_17333);
and U20692 (N_20692,N_17152,N_15814);
nand U20693 (N_20693,N_15368,N_17685);
nor U20694 (N_20694,N_16706,N_17397);
or U20695 (N_20695,N_16813,N_15361);
and U20696 (N_20696,N_15177,N_15049);
or U20697 (N_20697,N_16589,N_15250);
and U20698 (N_20698,N_16529,N_16340);
xor U20699 (N_20699,N_16365,N_17072);
and U20700 (N_20700,N_15649,N_17223);
nand U20701 (N_20701,N_15911,N_15606);
nand U20702 (N_20702,N_16036,N_16057);
nand U20703 (N_20703,N_15654,N_17796);
or U20704 (N_20704,N_17430,N_17144);
and U20705 (N_20705,N_16959,N_15485);
or U20706 (N_20706,N_17150,N_15562);
or U20707 (N_20707,N_15486,N_17488);
nor U20708 (N_20708,N_16763,N_15564);
nand U20709 (N_20709,N_16218,N_15915);
xor U20710 (N_20710,N_17435,N_17309);
nor U20711 (N_20711,N_16446,N_16641);
and U20712 (N_20712,N_16211,N_17564);
nor U20713 (N_20713,N_16154,N_15090);
nor U20714 (N_20714,N_17535,N_15693);
nand U20715 (N_20715,N_16836,N_16573);
nor U20716 (N_20716,N_15653,N_16804);
nor U20717 (N_20717,N_17136,N_17811);
xnor U20718 (N_20718,N_17578,N_17729);
or U20719 (N_20719,N_16735,N_17337);
nand U20720 (N_20720,N_16090,N_16024);
nand U20721 (N_20721,N_16531,N_17200);
or U20722 (N_20722,N_16394,N_17178);
nor U20723 (N_20723,N_17969,N_15768);
xnor U20724 (N_20724,N_16311,N_16182);
nor U20725 (N_20725,N_15480,N_15964);
and U20726 (N_20726,N_16858,N_15527);
nor U20727 (N_20727,N_15352,N_15956);
or U20728 (N_20728,N_15646,N_17846);
nor U20729 (N_20729,N_15864,N_17992);
nand U20730 (N_20730,N_16711,N_17928);
xnor U20731 (N_20731,N_15632,N_15262);
and U20732 (N_20732,N_16853,N_15964);
and U20733 (N_20733,N_16963,N_15037);
nand U20734 (N_20734,N_16418,N_17769);
xnor U20735 (N_20735,N_17670,N_16857);
nor U20736 (N_20736,N_15325,N_17717);
xnor U20737 (N_20737,N_16844,N_16191);
xor U20738 (N_20738,N_16587,N_15133);
or U20739 (N_20739,N_15497,N_15170);
nand U20740 (N_20740,N_16918,N_16049);
xnor U20741 (N_20741,N_17973,N_16706);
xnor U20742 (N_20742,N_15885,N_16389);
nand U20743 (N_20743,N_15825,N_15958);
and U20744 (N_20744,N_15229,N_16186);
nor U20745 (N_20745,N_15575,N_16897);
nor U20746 (N_20746,N_16275,N_16722);
xnor U20747 (N_20747,N_17698,N_15975);
or U20748 (N_20748,N_16201,N_15634);
xnor U20749 (N_20749,N_16134,N_17802);
and U20750 (N_20750,N_16124,N_16931);
nor U20751 (N_20751,N_17474,N_17122);
nand U20752 (N_20752,N_15183,N_15739);
xnor U20753 (N_20753,N_15384,N_16425);
nor U20754 (N_20754,N_15660,N_15747);
xor U20755 (N_20755,N_17085,N_17179);
nor U20756 (N_20756,N_16644,N_15831);
nor U20757 (N_20757,N_15836,N_16622);
and U20758 (N_20758,N_15743,N_15676);
xor U20759 (N_20759,N_17717,N_16817);
nand U20760 (N_20760,N_15903,N_16427);
nor U20761 (N_20761,N_17692,N_17946);
xor U20762 (N_20762,N_17703,N_15893);
nand U20763 (N_20763,N_17324,N_17685);
nor U20764 (N_20764,N_17672,N_17234);
xor U20765 (N_20765,N_17899,N_15936);
or U20766 (N_20766,N_15273,N_15264);
xor U20767 (N_20767,N_15712,N_15692);
xnor U20768 (N_20768,N_16250,N_16010);
nand U20769 (N_20769,N_15391,N_15600);
and U20770 (N_20770,N_15762,N_15426);
nand U20771 (N_20771,N_16406,N_16664);
and U20772 (N_20772,N_17661,N_15355);
nor U20773 (N_20773,N_16766,N_16213);
and U20774 (N_20774,N_15849,N_16443);
and U20775 (N_20775,N_16147,N_17920);
or U20776 (N_20776,N_17672,N_17053);
or U20777 (N_20777,N_16912,N_15868);
nor U20778 (N_20778,N_15565,N_15313);
nor U20779 (N_20779,N_15699,N_15620);
xnor U20780 (N_20780,N_16789,N_16673);
nor U20781 (N_20781,N_17158,N_16456);
and U20782 (N_20782,N_15015,N_17783);
nor U20783 (N_20783,N_17528,N_16122);
nand U20784 (N_20784,N_17829,N_17438);
xor U20785 (N_20785,N_16474,N_15772);
and U20786 (N_20786,N_17003,N_15472);
or U20787 (N_20787,N_17269,N_16900);
xnor U20788 (N_20788,N_16300,N_15194);
nor U20789 (N_20789,N_17938,N_17740);
nor U20790 (N_20790,N_15711,N_17801);
and U20791 (N_20791,N_17689,N_17721);
xnor U20792 (N_20792,N_17118,N_17942);
or U20793 (N_20793,N_17619,N_15878);
nand U20794 (N_20794,N_17388,N_17176);
and U20795 (N_20795,N_16359,N_15844);
nor U20796 (N_20796,N_16255,N_17943);
nor U20797 (N_20797,N_17631,N_16781);
and U20798 (N_20798,N_15575,N_17232);
or U20799 (N_20799,N_16051,N_16493);
and U20800 (N_20800,N_17058,N_15538);
nor U20801 (N_20801,N_15808,N_15861);
and U20802 (N_20802,N_16611,N_16893);
nand U20803 (N_20803,N_16377,N_15859);
nor U20804 (N_20804,N_17837,N_15287);
xnor U20805 (N_20805,N_15159,N_15454);
and U20806 (N_20806,N_17823,N_15525);
xor U20807 (N_20807,N_17177,N_15317);
and U20808 (N_20808,N_15207,N_17016);
nor U20809 (N_20809,N_16524,N_17409);
xnor U20810 (N_20810,N_16913,N_15506);
nand U20811 (N_20811,N_16310,N_17601);
xor U20812 (N_20812,N_16188,N_17165);
and U20813 (N_20813,N_17032,N_15579);
nand U20814 (N_20814,N_15195,N_16634);
nand U20815 (N_20815,N_15546,N_16087);
or U20816 (N_20816,N_16030,N_15233);
and U20817 (N_20817,N_17994,N_17530);
nor U20818 (N_20818,N_15271,N_17323);
or U20819 (N_20819,N_15778,N_15379);
or U20820 (N_20820,N_16677,N_16964);
nor U20821 (N_20821,N_16944,N_17737);
nor U20822 (N_20822,N_15362,N_15083);
or U20823 (N_20823,N_17752,N_16660);
nor U20824 (N_20824,N_16343,N_16449);
nor U20825 (N_20825,N_15535,N_15323);
xnor U20826 (N_20826,N_17753,N_16435);
or U20827 (N_20827,N_16281,N_15376);
xor U20828 (N_20828,N_15062,N_15836);
nand U20829 (N_20829,N_15844,N_17311);
xor U20830 (N_20830,N_17473,N_16222);
nor U20831 (N_20831,N_15116,N_16321);
and U20832 (N_20832,N_15748,N_16302);
xnor U20833 (N_20833,N_15029,N_16971);
or U20834 (N_20834,N_15366,N_17562);
nor U20835 (N_20835,N_15661,N_17732);
nand U20836 (N_20836,N_15241,N_16835);
nand U20837 (N_20837,N_17723,N_16684);
xor U20838 (N_20838,N_16344,N_16678);
nor U20839 (N_20839,N_16071,N_17187);
nand U20840 (N_20840,N_17504,N_17493);
nand U20841 (N_20841,N_16113,N_17841);
xnor U20842 (N_20842,N_16527,N_17003);
or U20843 (N_20843,N_15629,N_15524);
or U20844 (N_20844,N_15276,N_16112);
and U20845 (N_20845,N_16586,N_15866);
or U20846 (N_20846,N_17659,N_15511);
xnor U20847 (N_20847,N_17479,N_17668);
nor U20848 (N_20848,N_15266,N_15066);
xnor U20849 (N_20849,N_16155,N_17280);
xnor U20850 (N_20850,N_17597,N_17232);
nor U20851 (N_20851,N_15645,N_16561);
nor U20852 (N_20852,N_15651,N_16971);
nor U20853 (N_20853,N_15464,N_15744);
nand U20854 (N_20854,N_17153,N_16729);
and U20855 (N_20855,N_16301,N_17759);
nand U20856 (N_20856,N_17000,N_15765);
xor U20857 (N_20857,N_17513,N_15658);
nand U20858 (N_20858,N_17203,N_17095);
and U20859 (N_20859,N_17413,N_17895);
nand U20860 (N_20860,N_15236,N_17876);
xnor U20861 (N_20861,N_17252,N_15834);
nand U20862 (N_20862,N_15739,N_16315);
xor U20863 (N_20863,N_15542,N_17045);
xor U20864 (N_20864,N_16516,N_16409);
nor U20865 (N_20865,N_15514,N_16457);
xnor U20866 (N_20866,N_16147,N_17420);
xor U20867 (N_20867,N_16895,N_16386);
nand U20868 (N_20868,N_16478,N_17077);
and U20869 (N_20869,N_15438,N_16026);
nor U20870 (N_20870,N_15776,N_17624);
and U20871 (N_20871,N_17814,N_17254);
nand U20872 (N_20872,N_15452,N_16295);
or U20873 (N_20873,N_17512,N_15606);
nor U20874 (N_20874,N_16450,N_15900);
or U20875 (N_20875,N_15387,N_17001);
and U20876 (N_20876,N_17548,N_15382);
and U20877 (N_20877,N_17197,N_15124);
nand U20878 (N_20878,N_17707,N_16623);
xnor U20879 (N_20879,N_17819,N_17436);
nor U20880 (N_20880,N_15092,N_15802);
and U20881 (N_20881,N_15989,N_16329);
or U20882 (N_20882,N_16826,N_17977);
nor U20883 (N_20883,N_17327,N_17411);
xor U20884 (N_20884,N_17379,N_17722);
nand U20885 (N_20885,N_17942,N_15589);
nand U20886 (N_20886,N_16261,N_16673);
or U20887 (N_20887,N_17773,N_15082);
xor U20888 (N_20888,N_16444,N_15813);
nand U20889 (N_20889,N_17502,N_17190);
xnor U20890 (N_20890,N_16481,N_16251);
and U20891 (N_20891,N_16104,N_17749);
nor U20892 (N_20892,N_17623,N_17429);
xnor U20893 (N_20893,N_15301,N_17544);
nor U20894 (N_20894,N_17023,N_15328);
and U20895 (N_20895,N_15771,N_15203);
nand U20896 (N_20896,N_16924,N_16205);
and U20897 (N_20897,N_16323,N_17358);
xnor U20898 (N_20898,N_16511,N_16449);
nand U20899 (N_20899,N_17602,N_16781);
xor U20900 (N_20900,N_17755,N_17093);
or U20901 (N_20901,N_15373,N_17815);
nand U20902 (N_20902,N_15922,N_16070);
xnor U20903 (N_20903,N_16320,N_16011);
xor U20904 (N_20904,N_17688,N_15464);
and U20905 (N_20905,N_17961,N_17689);
and U20906 (N_20906,N_17350,N_16166);
and U20907 (N_20907,N_16669,N_17833);
xnor U20908 (N_20908,N_15225,N_16518);
nor U20909 (N_20909,N_16266,N_16918);
and U20910 (N_20910,N_17449,N_15799);
or U20911 (N_20911,N_15853,N_17926);
or U20912 (N_20912,N_16899,N_15232);
nor U20913 (N_20913,N_15387,N_15303);
or U20914 (N_20914,N_16816,N_15521);
nand U20915 (N_20915,N_16774,N_16293);
and U20916 (N_20916,N_16974,N_16598);
or U20917 (N_20917,N_15822,N_15784);
xnor U20918 (N_20918,N_15071,N_17685);
or U20919 (N_20919,N_16667,N_16112);
nand U20920 (N_20920,N_16409,N_15587);
and U20921 (N_20921,N_16305,N_15812);
nand U20922 (N_20922,N_15459,N_17828);
xor U20923 (N_20923,N_15162,N_17312);
and U20924 (N_20924,N_15800,N_16722);
nor U20925 (N_20925,N_17743,N_16055);
nand U20926 (N_20926,N_17258,N_16794);
xnor U20927 (N_20927,N_17486,N_16608);
xor U20928 (N_20928,N_17600,N_15705);
or U20929 (N_20929,N_16062,N_17826);
and U20930 (N_20930,N_15825,N_17273);
and U20931 (N_20931,N_15514,N_17927);
and U20932 (N_20932,N_16873,N_15700);
nand U20933 (N_20933,N_16786,N_15098);
nor U20934 (N_20934,N_15696,N_16752);
or U20935 (N_20935,N_15220,N_17548);
nand U20936 (N_20936,N_17560,N_15828);
or U20937 (N_20937,N_15176,N_17950);
or U20938 (N_20938,N_16056,N_15355);
and U20939 (N_20939,N_17887,N_15751);
or U20940 (N_20940,N_16142,N_16598);
and U20941 (N_20941,N_15343,N_15945);
xor U20942 (N_20942,N_16902,N_16466);
or U20943 (N_20943,N_17060,N_15124);
xnor U20944 (N_20944,N_16032,N_15087);
and U20945 (N_20945,N_16197,N_15792);
nor U20946 (N_20946,N_17713,N_17436);
or U20947 (N_20947,N_16122,N_16867);
nand U20948 (N_20948,N_15038,N_15416);
or U20949 (N_20949,N_17346,N_15238);
nor U20950 (N_20950,N_17127,N_17641);
nor U20951 (N_20951,N_17919,N_15383);
or U20952 (N_20952,N_15081,N_17473);
nor U20953 (N_20953,N_15421,N_16700);
nand U20954 (N_20954,N_17335,N_17489);
nor U20955 (N_20955,N_15244,N_15473);
and U20956 (N_20956,N_17111,N_16532);
or U20957 (N_20957,N_17374,N_16843);
and U20958 (N_20958,N_16419,N_16772);
and U20959 (N_20959,N_16174,N_15302);
nand U20960 (N_20960,N_17053,N_17468);
xnor U20961 (N_20961,N_17704,N_17766);
and U20962 (N_20962,N_17489,N_15374);
xor U20963 (N_20963,N_17336,N_17472);
and U20964 (N_20964,N_15107,N_17022);
xor U20965 (N_20965,N_17090,N_15146);
nor U20966 (N_20966,N_15852,N_17848);
or U20967 (N_20967,N_16502,N_17077);
or U20968 (N_20968,N_17676,N_15998);
nand U20969 (N_20969,N_16829,N_16251);
xnor U20970 (N_20970,N_17962,N_17310);
xnor U20971 (N_20971,N_17479,N_16032);
nor U20972 (N_20972,N_15144,N_16355);
nor U20973 (N_20973,N_15097,N_15352);
and U20974 (N_20974,N_17858,N_15410);
and U20975 (N_20975,N_17449,N_17906);
or U20976 (N_20976,N_16091,N_15929);
nor U20977 (N_20977,N_16983,N_17820);
xor U20978 (N_20978,N_15267,N_15463);
and U20979 (N_20979,N_16289,N_15089);
or U20980 (N_20980,N_16537,N_15814);
nor U20981 (N_20981,N_17682,N_17109);
nand U20982 (N_20982,N_16558,N_17294);
and U20983 (N_20983,N_15519,N_15792);
nor U20984 (N_20984,N_15857,N_15127);
nand U20985 (N_20985,N_16962,N_16804);
nand U20986 (N_20986,N_16389,N_16004);
nor U20987 (N_20987,N_17438,N_16211);
or U20988 (N_20988,N_17206,N_15656);
and U20989 (N_20989,N_16645,N_15749);
or U20990 (N_20990,N_17610,N_16241);
xnor U20991 (N_20991,N_17731,N_17823);
nand U20992 (N_20992,N_16675,N_17042);
or U20993 (N_20993,N_15174,N_15099);
or U20994 (N_20994,N_15365,N_17669);
or U20995 (N_20995,N_16604,N_15462);
nand U20996 (N_20996,N_15257,N_17007);
xor U20997 (N_20997,N_17008,N_17159);
and U20998 (N_20998,N_15790,N_17520);
and U20999 (N_20999,N_15783,N_17451);
and U21000 (N_21000,N_18958,N_18200);
and U21001 (N_21001,N_18223,N_18161);
nor U21002 (N_21002,N_19975,N_19594);
or U21003 (N_21003,N_20831,N_19143);
nand U21004 (N_21004,N_18427,N_19201);
nor U21005 (N_21005,N_18904,N_20553);
xnor U21006 (N_21006,N_18253,N_18300);
nor U21007 (N_21007,N_20737,N_19878);
nand U21008 (N_21008,N_19586,N_20129);
nand U21009 (N_21009,N_18713,N_20182);
nor U21010 (N_21010,N_18746,N_19185);
nand U21011 (N_21011,N_20720,N_18421);
nor U21012 (N_21012,N_18864,N_19607);
xor U21013 (N_21013,N_20342,N_20391);
nor U21014 (N_21014,N_18263,N_19520);
or U21015 (N_21015,N_19826,N_19895);
xor U21016 (N_21016,N_20983,N_19401);
nand U21017 (N_21017,N_18224,N_18041);
xor U21018 (N_21018,N_19810,N_20603);
nand U21019 (N_21019,N_18109,N_18750);
nand U21020 (N_21020,N_18890,N_18052);
nor U21021 (N_21021,N_20407,N_20344);
xnor U21022 (N_21022,N_18553,N_19085);
or U21023 (N_21023,N_18025,N_19868);
and U21024 (N_21024,N_20476,N_18309);
nor U21025 (N_21025,N_19277,N_19126);
nor U21026 (N_21026,N_18800,N_19656);
xnor U21027 (N_21027,N_20313,N_19617);
nor U21028 (N_21028,N_18605,N_20232);
nor U21029 (N_21029,N_19339,N_18671);
or U21030 (N_21030,N_20125,N_19765);
nor U21031 (N_21031,N_18008,N_19273);
and U21032 (N_21032,N_19861,N_19553);
nand U21033 (N_21033,N_19396,N_19596);
xnor U21034 (N_21034,N_20994,N_20289);
xnor U21035 (N_21035,N_18388,N_20543);
xor U21036 (N_21036,N_19735,N_20634);
or U21037 (N_21037,N_20462,N_18521);
nand U21038 (N_21038,N_18554,N_19335);
nand U21039 (N_21039,N_19777,N_19441);
nor U21040 (N_21040,N_19511,N_19857);
and U21041 (N_21041,N_20447,N_20378);
and U21042 (N_21042,N_20417,N_18013);
and U21043 (N_21043,N_19489,N_18289);
xnor U21044 (N_21044,N_20796,N_20561);
nand U21045 (N_21045,N_19111,N_19963);
nand U21046 (N_21046,N_18432,N_18349);
nor U21047 (N_21047,N_20879,N_19039);
nand U21048 (N_21048,N_18422,N_20485);
or U21049 (N_21049,N_18797,N_20691);
xor U21050 (N_21050,N_19803,N_18192);
nand U21051 (N_21051,N_18218,N_20638);
nor U21052 (N_21052,N_20173,N_18941);
nor U21053 (N_21053,N_18456,N_20893);
nand U21054 (N_21054,N_20293,N_18697);
or U21055 (N_21055,N_20774,N_20949);
and U21056 (N_21056,N_20657,N_19147);
or U21057 (N_21057,N_20220,N_20936);
nand U21058 (N_21058,N_20705,N_20132);
or U21059 (N_21059,N_19634,N_18573);
xor U21060 (N_21060,N_19746,N_20702);
or U21061 (N_21061,N_19896,N_18510);
and U21062 (N_21062,N_19574,N_19303);
and U21063 (N_21063,N_20904,N_18947);
or U21064 (N_21064,N_20397,N_18793);
nor U21065 (N_21065,N_19707,N_18882);
nor U21066 (N_21066,N_19679,N_20057);
nand U21067 (N_21067,N_20430,N_18257);
xor U21068 (N_21068,N_18572,N_19812);
or U21069 (N_21069,N_18649,N_19595);
or U21070 (N_21070,N_19612,N_18806);
or U21071 (N_21071,N_18972,N_19301);
and U21072 (N_21072,N_18466,N_20744);
and U21073 (N_21073,N_19853,N_18031);
or U21074 (N_21074,N_18485,N_18443);
nor U21075 (N_21075,N_20756,N_18540);
and U21076 (N_21076,N_18894,N_20593);
or U21077 (N_21077,N_19157,N_18121);
xnor U21078 (N_21078,N_19722,N_20834);
or U21079 (N_21079,N_20510,N_20729);
or U21080 (N_21080,N_19808,N_19446);
nand U21081 (N_21081,N_20009,N_18526);
and U21082 (N_21082,N_19940,N_20497);
nand U21083 (N_21083,N_20590,N_19429);
nor U21084 (N_21084,N_20083,N_20078);
and U21085 (N_21085,N_20206,N_19032);
xnor U21086 (N_21086,N_19877,N_18560);
xnor U21087 (N_21087,N_19800,N_18475);
and U21088 (N_21088,N_18799,N_19205);
nand U21089 (N_21089,N_19824,N_19738);
xnor U21090 (N_21090,N_20086,N_18870);
nor U21091 (N_21091,N_18429,N_18562);
and U21092 (N_21092,N_19976,N_20771);
nand U21093 (N_21093,N_19272,N_19716);
xor U21094 (N_21094,N_19398,N_19908);
or U21095 (N_21095,N_18463,N_20183);
nand U21096 (N_21096,N_20130,N_20789);
nor U21097 (N_21097,N_18663,N_18624);
nor U21098 (N_21098,N_18019,N_19364);
or U21099 (N_21099,N_20303,N_18804);
or U21100 (N_21100,N_18928,N_18711);
or U21101 (N_21101,N_20887,N_18255);
nor U21102 (N_21102,N_19203,N_19843);
nand U21103 (N_21103,N_18665,N_18791);
nand U21104 (N_21104,N_18323,N_19115);
and U21105 (N_21105,N_20360,N_19180);
and U21106 (N_21106,N_18499,N_20586);
nor U21107 (N_21107,N_19996,N_18504);
nand U21108 (N_21108,N_19954,N_20808);
nor U21109 (N_21109,N_20519,N_18460);
or U21110 (N_21110,N_18126,N_20810);
nand U21111 (N_21111,N_20516,N_20653);
nor U21112 (N_21112,N_19320,N_18749);
or U21113 (N_21113,N_18637,N_20703);
or U21114 (N_21114,N_20168,N_18459);
xor U21115 (N_21115,N_18868,N_18285);
and U21116 (N_21116,N_19757,N_20885);
and U21117 (N_21117,N_20223,N_20048);
nand U21118 (N_21118,N_19033,N_18401);
xor U21119 (N_21119,N_18513,N_18819);
nand U21120 (N_21120,N_20514,N_19845);
nand U21121 (N_21121,N_19493,N_19183);
xnor U21122 (N_21122,N_20038,N_19353);
and U21123 (N_21123,N_18563,N_19282);
or U21124 (N_21124,N_19733,N_20861);
or U21125 (N_21125,N_20375,N_20148);
and U21126 (N_21126,N_18174,N_20572);
nor U21127 (N_21127,N_19099,N_18943);
xnor U21128 (N_21128,N_18351,N_18133);
xnor U21129 (N_21129,N_18853,N_19864);
or U21130 (N_21130,N_18375,N_20785);
nand U21131 (N_21131,N_19740,N_20860);
xnor U21132 (N_21132,N_19955,N_18875);
xnor U21133 (N_21133,N_19584,N_18970);
nor U21134 (N_21134,N_20929,N_19044);
nand U21135 (N_21135,N_19713,N_19342);
nor U21136 (N_21136,N_19967,N_19268);
or U21137 (N_21137,N_20570,N_18143);
nand U21138 (N_21138,N_18018,N_20413);
and U21139 (N_21139,N_19542,N_20560);
nor U21140 (N_21140,N_20311,N_19070);
and U21141 (N_21141,N_18311,N_20478);
nand U21142 (N_21142,N_20833,N_20601);
or U21143 (N_21143,N_20135,N_18036);
nor U21144 (N_21144,N_19223,N_18156);
or U21145 (N_21145,N_20911,N_18846);
and U21146 (N_21146,N_20169,N_20645);
nand U21147 (N_21147,N_19754,N_19762);
or U21148 (N_21148,N_20315,N_19181);
nand U21149 (N_21149,N_18215,N_20882);
nor U21150 (N_21150,N_19731,N_18211);
nor U21151 (N_21151,N_18337,N_19238);
or U21152 (N_21152,N_19726,N_18680);
and U21153 (N_21153,N_18887,N_19382);
nor U21154 (N_21154,N_18472,N_18653);
nor U21155 (N_21155,N_18145,N_19992);
nand U21156 (N_21156,N_18382,N_19890);
nor U21157 (N_21157,N_18395,N_19621);
xor U21158 (N_21158,N_19444,N_20990);
and U21159 (N_21159,N_18998,N_20963);
nand U21160 (N_21160,N_19755,N_18938);
xnor U21161 (N_21161,N_19240,N_18623);
xor U21162 (N_21162,N_19789,N_19776);
nor U21163 (N_21163,N_20002,N_19611);
nor U21164 (N_21164,N_20575,N_19072);
nand U21165 (N_21165,N_20946,N_18674);
and U21166 (N_21166,N_19415,N_19737);
and U21167 (N_21167,N_20512,N_18759);
nand U21168 (N_21168,N_18178,N_18157);
and U21169 (N_21169,N_19347,N_19197);
and U21170 (N_21170,N_18328,N_18493);
xnor U21171 (N_21171,N_20120,N_20938);
xnor U21172 (N_21172,N_19253,N_18542);
nand U21173 (N_21173,N_18641,N_19941);
or U21174 (N_21174,N_18181,N_20014);
xor U21175 (N_21175,N_18518,N_20773);
xnor U21176 (N_21176,N_19426,N_19051);
xnor U21177 (N_21177,N_19951,N_19291);
xor U21178 (N_21178,N_20186,N_18770);
nor U21179 (N_21179,N_20473,N_20174);
xnor U21180 (N_21180,N_20469,N_20905);
or U21181 (N_21181,N_18915,N_18616);
or U21182 (N_21182,N_19334,N_20386);
and U21183 (N_21183,N_18268,N_19948);
xor U21184 (N_21184,N_18079,N_20244);
xnor U21185 (N_21185,N_19552,N_19593);
or U21186 (N_21186,N_19189,N_19079);
nor U21187 (N_21187,N_18503,N_20082);
nor U21188 (N_21188,N_18301,N_20141);
xor U21189 (N_21189,N_18033,N_19094);
nand U21190 (N_21190,N_20827,N_20266);
and U21191 (N_21191,N_19781,N_19966);
xor U21192 (N_21192,N_19608,N_18940);
xnor U21193 (N_21193,N_20433,N_18247);
and U21194 (N_21194,N_18537,N_19406);
or U21195 (N_21195,N_20323,N_19638);
nand U21196 (N_21196,N_18000,N_19784);
or U21197 (N_21197,N_18840,N_19515);
or U21198 (N_21198,N_18108,N_19249);
and U21199 (N_21199,N_20448,N_20072);
xnor U21200 (N_21200,N_19131,N_20330);
and U21201 (N_21201,N_20114,N_18555);
nor U21202 (N_21202,N_19293,N_19388);
xnor U21203 (N_21203,N_18264,N_18015);
xor U21204 (N_21204,N_18815,N_20542);
nor U21205 (N_21205,N_19547,N_18135);
nand U21206 (N_21206,N_18372,N_20111);
nand U21207 (N_21207,N_19438,N_20506);
or U21208 (N_21208,N_18557,N_20370);
or U21209 (N_21209,N_19807,N_18104);
nand U21210 (N_21210,N_19215,N_20492);
and U21211 (N_21211,N_20380,N_19255);
or U21212 (N_21212,N_18269,N_19306);
or U21213 (N_21213,N_20919,N_20589);
xnor U21214 (N_21214,N_20405,N_19903);
nand U21215 (N_21215,N_18210,N_18613);
or U21216 (N_21216,N_20906,N_20611);
nor U21217 (N_21217,N_19770,N_18185);
or U21218 (N_21218,N_20346,N_18040);
and U21219 (N_21219,N_19121,N_19926);
or U21220 (N_21220,N_20486,N_20224);
and U21221 (N_21221,N_18974,N_19891);
nor U21222 (N_21222,N_18294,N_20468);
nand U21223 (N_21223,N_20364,N_18175);
and U21224 (N_21224,N_18619,N_20942);
nor U21225 (N_21225,N_19471,N_19299);
nand U21226 (N_21226,N_18968,N_18534);
or U21227 (N_21227,N_18775,N_18752);
nand U21228 (N_21228,N_20715,N_19312);
xnor U21229 (N_21229,N_20727,N_19905);
nor U21230 (N_21230,N_18198,N_19799);
nand U21231 (N_21231,N_19886,N_18646);
or U21232 (N_21232,N_19743,N_20193);
xor U21233 (N_21233,N_18760,N_18638);
nor U21234 (N_21234,N_18390,N_19164);
and U21235 (N_21235,N_20354,N_19508);
and U21236 (N_21236,N_20208,N_20353);
nor U21237 (N_21237,N_18709,N_18841);
nor U21238 (N_21238,N_19324,N_18001);
xnor U21239 (N_21239,N_19919,N_19610);
or U21240 (N_21240,N_20219,N_18107);
xor U21241 (N_21241,N_18457,N_18802);
or U21242 (N_21242,N_19606,N_20373);
or U21243 (N_21243,N_19927,N_20243);
or U21244 (N_21244,N_20445,N_18235);
xor U21245 (N_21245,N_20273,N_18384);
and U21246 (N_21246,N_18444,N_18072);
or U21247 (N_21247,N_18229,N_19822);
xor U21248 (N_21248,N_18676,N_18071);
and U21249 (N_21249,N_19972,N_18705);
or U21250 (N_21250,N_19912,N_19830);
and U21251 (N_21251,N_20803,N_19659);
nand U21252 (N_21252,N_19260,N_19866);
and U21253 (N_21253,N_18528,N_19235);
and U21254 (N_21254,N_20844,N_18441);
and U21255 (N_21255,N_20275,N_18524);
and U21256 (N_21256,N_18392,N_20846);
nand U21257 (N_21257,N_18789,N_19145);
nor U21258 (N_21258,N_20137,N_18159);
nor U21259 (N_21259,N_18176,N_20961);
or U21260 (N_21260,N_20976,N_18465);
nand U21261 (N_21261,N_20830,N_19880);
and U21262 (N_21262,N_18964,N_18533);
nor U21263 (N_21263,N_20240,N_18413);
xnor U21264 (N_21264,N_19624,N_19329);
nor U21265 (N_21265,N_20334,N_20369);
nand U21266 (N_21266,N_18902,N_20056);
xor U21267 (N_21267,N_20805,N_20187);
and U21268 (N_21268,N_19583,N_20922);
xor U21269 (N_21269,N_18276,N_20863);
nor U21270 (N_21270,N_19805,N_20063);
nand U21271 (N_21271,N_18796,N_20118);
and U21272 (N_21272,N_19297,N_19597);
nand U21273 (N_21273,N_20167,N_19958);
nand U21274 (N_21274,N_18618,N_18411);
xor U21275 (N_21275,N_19491,N_20680);
xnor U21276 (N_21276,N_19831,N_18827);
nand U21277 (N_21277,N_18244,N_19832);
nand U21278 (N_21278,N_18869,N_19988);
nand U21279 (N_21279,N_18230,N_19663);
nor U21280 (N_21280,N_19969,N_20857);
xor U21281 (N_21281,N_19113,N_19788);
and U21282 (N_21282,N_20787,N_18855);
or U21283 (N_21283,N_19809,N_19524);
nor U21284 (N_21284,N_18483,N_18895);
xor U21285 (N_21285,N_18569,N_19869);
nand U21286 (N_21286,N_20674,N_19474);
nand U21287 (N_21287,N_18381,N_20799);
and U21288 (N_21288,N_18509,N_18330);
nand U21289 (N_21289,N_19742,N_18719);
xor U21290 (N_21290,N_19821,N_18614);
xnor U21291 (N_21291,N_20161,N_20775);
xor U21292 (N_21292,N_19623,N_19437);
or U21293 (N_21293,N_19098,N_18380);
nor U21294 (N_21294,N_18822,N_19395);
xor U21295 (N_21295,N_19753,N_19495);
xor U21296 (N_21296,N_18609,N_18856);
and U21297 (N_21297,N_20035,N_19016);
nand U21298 (N_21298,N_19688,N_20006);
nand U21299 (N_21299,N_18452,N_18738);
nor U21300 (N_21300,N_19723,N_18197);
xor U21301 (N_21301,N_19206,N_19798);
xnor U21302 (N_21302,N_18782,N_18361);
or U21303 (N_21303,N_20227,N_19413);
nor U21304 (N_21304,N_18993,N_18847);
or U21305 (N_21305,N_20716,N_20097);
or U21306 (N_21306,N_18721,N_20900);
nand U21307 (N_21307,N_20849,N_20229);
or U21308 (N_21308,N_19355,N_20019);
and U21309 (N_21309,N_20113,N_20207);
xnor U21310 (N_21310,N_19137,N_18897);
nor U21311 (N_21311,N_20112,N_20203);
xor U21312 (N_21312,N_18730,N_18691);
nor U21313 (N_21313,N_18136,N_20614);
nor U21314 (N_21314,N_19778,N_19117);
xor U21315 (N_21315,N_20284,N_20644);
nor U21316 (N_21316,N_18669,N_19862);
and U21317 (N_21317,N_18281,N_20608);
nand U21318 (N_21318,N_18273,N_20088);
or U21319 (N_21319,N_20684,N_18843);
xor U21320 (N_21320,N_18881,N_20176);
xnor U21321 (N_21321,N_20084,N_19818);
xnor U21322 (N_21322,N_18470,N_20152);
or U21323 (N_21323,N_19641,N_19643);
and U21324 (N_21324,N_19374,N_18474);
xor U21325 (N_21325,N_20390,N_20046);
or U21326 (N_21326,N_19962,N_19785);
nor U21327 (N_21327,N_19747,N_18595);
and U21328 (N_21328,N_18580,N_20443);
or U21329 (N_21329,N_18559,N_19519);
xnor U21330 (N_21330,N_20673,N_18689);
nand U21331 (N_21331,N_20779,N_20962);
nand U21332 (N_21332,N_20957,N_20915);
xnor U21333 (N_21333,N_19626,N_19899);
or U21334 (N_21334,N_18462,N_20899);
and U21335 (N_21335,N_18758,N_18433);
and U21336 (N_21336,N_18944,N_19211);
xor U21337 (N_21337,N_18854,N_19184);
and U21338 (N_21338,N_18536,N_18310);
nor U21339 (N_21339,N_20274,N_18583);
or U21340 (N_21340,N_19834,N_20117);
or U21341 (N_21341,N_19448,N_18809);
or U21342 (N_21342,N_20842,N_18666);
xnor U21343 (N_21343,N_18383,N_18515);
or U21344 (N_21344,N_20852,N_18450);
nor U21345 (N_21345,N_18773,N_19013);
nand U21346 (N_21346,N_19363,N_18673);
xor U21347 (N_21347,N_19083,N_19420);
nor U21348 (N_21348,N_18836,N_18724);
and U21349 (N_21349,N_20459,N_18714);
nand U21350 (N_21350,N_19871,N_18756);
nor U21351 (N_21351,N_19207,N_18265);
nand U21352 (N_21352,N_19008,N_19337);
nand U21353 (N_21353,N_20299,N_18507);
nand U21354 (N_21354,N_19175,N_18453);
nand U21355 (N_21355,N_18657,N_18919);
nor U21356 (N_21356,N_20321,N_18949);
nor U21357 (N_21357,N_20965,N_20339);
nand U21358 (N_21358,N_19466,N_19771);
nand U21359 (N_21359,N_18908,N_20331);
nand U21360 (N_21360,N_18593,N_18857);
or U21361 (N_21361,N_19631,N_20625);
or U21362 (N_21362,N_18948,N_18322);
xor U21363 (N_21363,N_18929,N_20766);
nor U21364 (N_21364,N_19011,N_19526);
nor U21365 (N_21365,N_18408,N_20754);
or U21366 (N_21366,N_18339,N_18734);
nor U21367 (N_21367,N_19604,N_20429);
or U21368 (N_21368,N_20719,N_18530);
nand U21369 (N_21369,N_19950,N_18129);
nor U21370 (N_21370,N_19144,N_19528);
nand U21371 (N_21371,N_18007,N_19411);
nand U21372 (N_21372,N_18587,N_19484);
nand U21373 (N_21373,N_18042,N_20341);
nand U21374 (N_21374,N_20934,N_19691);
xnor U21375 (N_21375,N_18306,N_20730);
xnor U21376 (N_21376,N_18102,N_18122);
or U21377 (N_21377,N_18716,N_20633);
and U21378 (N_21378,N_20968,N_19535);
nand U21379 (N_21379,N_20947,N_19993);
or U21380 (N_21380,N_20242,N_20298);
nor U21381 (N_21381,N_18581,N_20616);
or U21382 (N_21382,N_20998,N_20986);
nor U21383 (N_21383,N_19436,N_18118);
nand U21384 (N_21384,N_19427,N_20277);
or U21385 (N_21385,N_19046,N_18704);
nand U21386 (N_21386,N_18766,N_19431);
nor U21387 (N_21387,N_18718,N_19501);
xnor U21388 (N_21388,N_18741,N_18514);
or U21389 (N_21389,N_20491,N_20425);
xor U21390 (N_21390,N_19561,N_18446);
nand U21391 (N_21391,N_20356,N_18893);
or U21392 (N_21392,N_18282,N_19412);
nor U21393 (N_21393,N_19182,N_20080);
or U21394 (N_21394,N_20432,N_18034);
nor U21395 (N_21395,N_20697,N_18952);
nor U21396 (N_21396,N_20000,N_19802);
nand U21397 (N_21397,N_18240,N_20689);
nand U21398 (N_21398,N_18021,N_20843);
nand U21399 (N_21399,N_18907,N_18014);
nor U21400 (N_21400,N_20073,N_18124);
or U21401 (N_21401,N_20108,N_19823);
xor U21402 (N_21402,N_19487,N_20527);
and U21403 (N_21403,N_19846,N_19579);
or U21404 (N_21404,N_20595,N_20454);
nand U21405 (N_21405,N_20982,N_20667);
xnor U21406 (N_21406,N_19024,N_20768);
xor U21407 (N_21407,N_18883,N_20579);
xnor U21408 (N_21408,N_20023,N_20622);
xnor U21409 (N_21409,N_20455,N_20412);
or U21410 (N_21410,N_19825,N_18055);
nand U21411 (N_21411,N_18763,N_20555);
xnor U21412 (N_21412,N_20932,N_19684);
xor U21413 (N_21413,N_18538,N_18226);
or U21414 (N_21414,N_18468,N_19275);
and U21415 (N_21415,N_19366,N_19479);
and U21416 (N_21416,N_20735,N_20672);
and U21417 (N_21417,N_20828,N_20870);
and U21418 (N_21418,N_20098,N_20956);
and U21419 (N_21419,N_20007,N_18873);
and U21420 (N_21420,N_19669,N_18821);
xor U21421 (N_21421,N_18279,N_20253);
nor U21422 (N_21422,N_18062,N_20204);
xnor U21423 (N_21423,N_19724,N_20191);
nand U21424 (N_21424,N_20003,N_19222);
nand U21425 (N_21425,N_19300,N_20794);
and U21426 (N_21426,N_18137,N_18017);
and U21427 (N_21427,N_20862,N_18978);
or U21428 (N_21428,N_19380,N_19763);
or U21429 (N_21429,N_20295,N_19461);
or U21430 (N_21430,N_20138,N_19739);
xor U21431 (N_21431,N_18410,N_20690);
xnor U21432 (N_21432,N_19425,N_19149);
xnor U21433 (N_21433,N_18527,N_18205);
or U21434 (N_21434,N_18199,N_20669);
nor U21435 (N_21435,N_20767,N_18561);
xnor U21436 (N_21436,N_20257,N_19835);
or U21437 (N_21437,N_19794,N_20874);
and U21438 (N_21438,N_20359,N_18078);
and U21439 (N_21439,N_18747,N_19344);
nor U21440 (N_21440,N_20145,N_20820);
xnor U21441 (N_21441,N_19901,N_20875);
nor U21442 (N_21442,N_18389,N_20126);
nor U21443 (N_21443,N_19158,N_19061);
xnor U21444 (N_21444,N_18083,N_18877);
nand U21445 (N_21445,N_19793,N_20267);
or U21446 (N_21446,N_18054,N_20461);
nand U21447 (N_21447,N_19680,N_18829);
nor U21448 (N_21448,N_19587,N_20192);
nand U21449 (N_21449,N_20308,N_18794);
nand U21450 (N_21450,N_19378,N_20881);
and U21451 (N_21451,N_18367,N_19708);
nor U21452 (N_21452,N_18428,N_19964);
and U21453 (N_21453,N_18622,N_20818);
nand U21454 (N_21454,N_18814,N_19327);
and U21455 (N_21455,N_20565,N_19360);
nor U21456 (N_21456,N_18757,N_20959);
xor U21457 (N_21457,N_18787,N_20095);
and U21458 (N_21458,N_20972,N_20571);
or U21459 (N_21459,N_19168,N_18725);
xnor U21460 (N_21460,N_20695,N_19837);
nor U21461 (N_21461,N_19959,N_19827);
nand U21462 (N_21462,N_20738,N_20851);
and U21463 (N_21463,N_18303,N_18731);
nand U21464 (N_21464,N_19994,N_18099);
and U21465 (N_21465,N_20474,N_20517);
nand U21466 (N_21466,N_20637,N_20508);
or U21467 (N_21467,N_19460,N_20610);
and U21468 (N_21468,N_19359,N_18011);
or U21469 (N_21469,N_19893,N_18818);
and U21470 (N_21470,N_19775,N_18082);
nor U21471 (N_21471,N_19585,N_20858);
nor U21472 (N_21472,N_20538,N_20952);
nand U21473 (N_21473,N_20939,N_19106);
nand U21474 (N_21474,N_18859,N_20646);
nand U21475 (N_21475,N_18440,N_19397);
nor U21476 (N_21476,N_19549,N_20066);
and U21477 (N_21477,N_20709,N_19923);
nor U21478 (N_21478,N_19577,N_20055);
xnor U21479 (N_21479,N_19256,N_18278);
and U21480 (N_21480,N_19251,N_20550);
xor U21481 (N_21481,N_19443,N_20530);
or U21482 (N_21482,N_20535,N_20248);
nor U21483 (N_21483,N_20978,N_20580);
or U21484 (N_21484,N_18584,N_20977);
or U21485 (N_21485,N_19555,N_18103);
nor U21486 (N_21486,N_20401,N_20150);
xor U21487 (N_21487,N_18251,N_19816);
or U21488 (N_21488,N_18291,N_20623);
nand U21489 (N_21489,N_18491,N_20398);
or U21490 (N_21490,N_19760,N_18329);
and U21491 (N_21491,N_20345,N_20792);
and U21492 (N_21492,N_18642,N_18308);
nand U21493 (N_21493,N_20013,N_19539);
nand U21494 (N_21494,N_20573,N_18274);
and U21495 (N_21495,N_20795,N_20696);
and U21496 (N_21496,N_19567,N_20418);
nand U21497 (N_21497,N_19404,N_19936);
nor U21498 (N_21498,N_18652,N_18032);
or U21499 (N_21499,N_18471,N_18973);
nand U21500 (N_21500,N_19125,N_18267);
nor U21501 (N_21501,N_20008,N_20935);
and U21502 (N_21502,N_20605,N_19410);
nand U21503 (N_21503,N_20707,N_18629);
nor U21504 (N_21504,N_20999,N_18636);
xor U21505 (N_21505,N_20297,N_20835);
or U21506 (N_21506,N_18213,N_18567);
xor U21507 (N_21507,N_20261,N_20062);
xor U21508 (N_21508,N_18312,N_18299);
and U21509 (N_21509,N_20711,N_18173);
xnor U21510 (N_21510,N_19408,N_18737);
xnor U21511 (N_21511,N_18350,N_19455);
nor U21512 (N_21512,N_19981,N_18073);
nor U21513 (N_21513,N_20399,N_20419);
nor U21514 (N_21514,N_19054,N_19889);
and U21515 (N_21515,N_19689,N_19195);
and U21516 (N_21516,N_19243,N_19178);
nor U21517 (N_21517,N_19224,N_20237);
xor U21518 (N_21518,N_19714,N_20495);
nor U21519 (N_21519,N_20172,N_18183);
nor U21520 (N_21520,N_18356,N_18458);
or U21521 (N_21521,N_20258,N_20597);
or U21522 (N_21522,N_18620,N_18611);
and U21523 (N_21523,N_20306,N_18110);
or U21524 (N_21524,N_20434,N_19409);
nand U21525 (N_21525,N_19968,N_19390);
xnor U21526 (N_21526,N_18551,N_18956);
xnor U21527 (N_21527,N_19002,N_20352);
or U21528 (N_21528,N_18900,N_20071);
and U21529 (N_21529,N_19109,N_19531);
or U21530 (N_21530,N_19541,N_20175);
or U21531 (N_21531,N_20903,N_18347);
xnor U21532 (N_21532,N_20499,N_19854);
and U21533 (N_21533,N_19108,N_20723);
nand U21534 (N_21534,N_19569,N_19063);
and U21535 (N_21535,N_20596,N_19190);
nand U21536 (N_21536,N_20181,N_19933);
xor U21537 (N_21537,N_20065,N_18736);
or U21538 (N_21538,N_18354,N_18830);
nand U21539 (N_21539,N_19169,N_18028);
or U21540 (N_21540,N_18270,N_19354);
or U21541 (N_21541,N_18597,N_18101);
or U21542 (N_21542,N_20093,N_18774);
xor U21543 (N_21543,N_20782,N_20943);
nand U21544 (N_21544,N_18848,N_19156);
xor U21545 (N_21545,N_18933,N_20357);
xnor U21546 (N_21546,N_18579,N_18795);
xor U21547 (N_21547,N_19122,N_20464);
nand U21548 (N_21548,N_18942,N_18425);
nand U21549 (N_21549,N_20416,N_19598);
and U21550 (N_21550,N_19118,N_20384);
and U21551 (N_21551,N_19451,N_20146);
nand U21552 (N_21552,N_20487,N_19176);
and U21553 (N_21553,N_18926,N_20800);
or U21554 (N_21554,N_20692,N_20250);
or U21555 (N_21555,N_18788,N_18955);
and U21556 (N_21556,N_19292,N_20609);
nor U21557 (N_21557,N_19730,N_20049);
nor U21558 (N_21558,N_19562,N_20739);
nor U21559 (N_21559,N_18068,N_20040);
nor U21560 (N_21560,N_20160,N_20995);
nor U21561 (N_21561,N_18729,N_18690);
nor U21562 (N_21562,N_20713,N_19309);
and U21563 (N_21563,N_19467,N_20896);
or U21564 (N_21564,N_20801,N_19841);
and U21565 (N_21565,N_19371,N_18243);
nor U21566 (N_21566,N_20490,N_19879);
nand U21567 (N_21567,N_18517,N_19850);
xnor U21568 (N_21568,N_19305,N_19219);
nand U21569 (N_21569,N_20195,N_18698);
and U21570 (N_21570,N_18828,N_20154);
or U21571 (N_21571,N_20850,N_18026);
nand U21572 (N_21572,N_20764,N_19314);
nor U21573 (N_21573,N_20470,N_18292);
nor U21574 (N_21574,N_18385,N_18767);
nand U21575 (N_21575,N_20873,N_20042);
or U21576 (N_21576,N_20740,N_19573);
nor U21577 (N_21577,N_20467,N_18761);
and U21578 (N_21578,N_18063,N_19081);
nor U21579 (N_21579,N_19720,N_18262);
or U21580 (N_21580,N_19946,N_20028);
nor U21581 (N_21581,N_18353,N_18575);
or U21582 (N_21582,N_20757,N_20089);
xor U21583 (N_21583,N_18832,N_18903);
nand U21584 (N_21584,N_20749,N_20194);
nand U21585 (N_21585,N_18190,N_18045);
and U21586 (N_21586,N_20090,N_20964);
or U21587 (N_21587,N_20650,N_18088);
and U21588 (N_21588,N_20515,N_20676);
and U21589 (N_21589,N_18650,N_18030);
nor U21590 (N_21590,N_19833,N_20276);
and U21591 (N_21591,N_19523,N_20269);
and U21592 (N_21592,N_20493,N_19613);
nand U21593 (N_21593,N_20142,N_18442);
nor U21594 (N_21594,N_19650,N_20246);
or U21595 (N_21595,N_18643,N_20780);
xnor U21596 (N_21596,N_20351,N_20980);
and U21597 (N_21597,N_18825,N_19661);
or U21598 (N_21598,N_20102,N_20675);
or U21599 (N_21599,N_20329,N_19038);
nand U21600 (N_21600,N_20200,N_18051);
nor U21601 (N_21601,N_19198,N_20688);
nor U21602 (N_21602,N_20414,N_20379);
nor U21603 (N_21603,N_19172,N_19407);
nor U21604 (N_21604,N_18860,N_19234);
xor U21605 (N_21605,N_18111,N_20128);
or U21606 (N_21606,N_18469,N_18820);
nand U21607 (N_21607,N_19450,N_18307);
nand U21608 (N_21608,N_20544,N_20921);
nor U21609 (N_21609,N_20325,N_18574);
xnor U21610 (N_21610,N_19086,N_19161);
xnor U21611 (N_21611,N_19322,N_19192);
nor U21612 (N_21612,N_19699,N_20950);
nand U21613 (N_21613,N_18152,N_18961);
or U21614 (N_21614,N_18925,N_20234);
nor U21615 (N_21615,N_20324,N_18723);
xnor U21616 (N_21616,N_19060,N_18971);
nand U21617 (N_21617,N_18505,N_20365);
or U21618 (N_21618,N_20436,N_19490);
or U21619 (N_21619,N_18128,N_19973);
nor U21620 (N_21620,N_18996,N_20296);
xnor U21621 (N_21621,N_20427,N_19852);
xnor U21622 (N_21622,N_20513,N_18187);
or U21623 (N_21623,N_19654,N_20180);
and U21624 (N_21624,N_19662,N_19296);
nor U21625 (N_21625,N_18043,N_20765);
nor U21626 (N_21626,N_20772,N_19998);
xor U21627 (N_21627,N_18430,N_19304);
nand U21628 (N_21628,N_18371,N_18639);
and U21629 (N_21629,N_19226,N_20725);
and U21630 (N_21630,N_18149,N_19073);
nor U21631 (N_21631,N_19751,N_19625);
and U21632 (N_21632,N_20326,N_20670);
nor U21633 (N_21633,N_18119,N_20291);
nor U21634 (N_21634,N_19261,N_19332);
xnor U21635 (N_21635,N_19375,N_20840);
xor U21636 (N_21636,N_20435,N_20123);
nor U21637 (N_21637,N_19855,N_18029);
xor U21638 (N_21638,N_19294,N_19422);
xor U21639 (N_21639,N_18997,N_19130);
xnor U21640 (N_21640,N_19673,N_19554);
or U21641 (N_21641,N_19154,N_20471);
nand U21642 (N_21642,N_19365,N_19048);
nand U21643 (N_21643,N_20721,N_18745);
or U21644 (N_21644,N_18061,N_20812);
nand U21645 (N_21645,N_20664,N_19434);
xnor U21646 (N_21646,N_18332,N_19924);
or U21647 (N_21647,N_19066,N_19120);
xor U21648 (N_21648,N_19875,N_20902);
xor U21649 (N_21649,N_19470,N_18113);
xor U21650 (N_21650,N_20845,N_20880);
nor U21651 (N_21651,N_18100,N_18748);
nand U21652 (N_21652,N_20559,N_19037);
xnor U21653 (N_21653,N_20958,N_20439);
and U21654 (N_21654,N_18193,N_20981);
xor U21655 (N_21655,N_18438,N_19942);
nor U21656 (N_21656,N_19019,N_19870);
nand U21657 (N_21657,N_19697,N_18212);
or U21658 (N_21658,N_19527,N_19346);
or U21659 (N_21659,N_19544,N_20635);
xnor U21660 (N_21660,N_20070,N_20472);
xor U21661 (N_21661,N_19637,N_20892);
nor U21662 (N_21662,N_20235,N_19482);
and U21663 (N_21663,N_18047,N_19828);
and U21664 (N_21664,N_18314,N_18345);
or U21665 (N_21665,N_20993,N_19307);
nor U21666 (N_21666,N_18246,N_20966);
xor U21667 (N_21667,N_18081,N_20005);
nand U21668 (N_21668,N_20388,N_20973);
and U21669 (N_21669,N_20358,N_18962);
xor U21670 (N_21670,N_18715,N_19208);
or U21671 (N_21671,N_20824,N_20221);
and U21672 (N_21672,N_20115,N_20338);
nor U21673 (N_21673,N_20037,N_19376);
xnor U21674 (N_21674,N_20525,N_18418);
xor U21675 (N_21675,N_19333,N_20829);
xor U21676 (N_21676,N_19931,N_18906);
nand U21677 (N_21677,N_20582,N_19863);
nor U21678 (N_21678,N_18685,N_20872);
and U21679 (N_21679,N_18975,N_19394);
nand U21680 (N_21680,N_18874,N_20316);
or U21681 (N_21681,N_20908,N_19295);
nor U21682 (N_21682,N_20975,N_20918);
nor U21683 (N_21683,N_20587,N_19909);
nor U21684 (N_21684,N_20494,N_19766);
or U21685 (N_21685,N_18365,N_20547);
or U21686 (N_21686,N_19683,N_19392);
nor U21687 (N_21687,N_20894,N_20163);
xnor U21688 (N_21688,N_18910,N_20811);
xnor U21689 (N_21689,N_19384,N_18377);
nor U21690 (N_21690,N_20626,N_19510);
nand U21691 (N_21691,N_18954,N_18409);
nand U21692 (N_21692,N_19664,N_20641);
or U21693 (N_21693,N_19814,N_18688);
and U21694 (N_21694,N_20778,N_19741);
and U21695 (N_21695,N_20233,N_20682);
nor U21696 (N_21696,N_18529,N_20157);
nor U21697 (N_21697,N_20604,N_20528);
xnor U21698 (N_21698,N_19475,N_18046);
xor U21699 (N_21699,N_18325,N_18654);
or U21700 (N_21700,N_19225,N_20997);
nor U21701 (N_21701,N_19907,N_20848);
nand U21702 (N_21702,N_20256,N_20821);
and U21703 (N_21703,N_18627,N_18436);
nand U21704 (N_21704,N_18899,N_19315);
or U21705 (N_21705,N_19635,N_20050);
or U21706 (N_21706,N_20534,N_20750);
nand U21707 (N_21707,N_19015,N_19774);
xor U21708 (N_21708,N_20970,N_18256);
and U21709 (N_21709,N_20985,N_18922);
xnor U21710 (N_21710,N_20030,N_19628);
and U21711 (N_21711,N_20155,N_19010);
nor U21712 (N_21712,N_19135,N_19900);
xnor U21713 (N_21713,N_18850,N_19045);
and U21714 (N_21714,N_18842,N_19012);
or U21715 (N_21715,N_19026,N_20909);
and U21716 (N_21716,N_18496,N_20826);
or U21717 (N_21717,N_18449,N_18640);
nor U21718 (N_21718,N_19265,N_18792);
xnor U21719 (N_21719,N_19499,N_20712);
nor U21720 (N_21720,N_19712,N_20283);
xnor U21721 (N_21721,N_19336,N_19050);
or U21722 (N_21722,N_19089,N_20133);
xor U21723 (N_21723,N_20091,N_18960);
nand U21724 (N_21724,N_19170,N_20131);
xnor U21725 (N_21725,N_19468,N_19417);
and U21726 (N_21726,N_19949,N_20300);
or U21727 (N_21727,N_19302,N_20521);
nand U21728 (N_21728,N_18556,N_18576);
nor U21729 (N_21729,N_18659,N_18437);
and U21730 (N_21730,N_19672,N_20629);
nand U21731 (N_21731,N_20558,N_18612);
xor U21732 (N_21732,N_18831,N_19529);
or U21733 (N_21733,N_18484,N_19564);
or U21734 (N_21734,N_19984,N_20483);
nand U21735 (N_21735,N_19883,N_18845);
xnor U21736 (N_21736,N_19744,N_19367);
and U21737 (N_21737,N_20698,N_20392);
and U21738 (N_21738,N_20280,N_20836);
and U21739 (N_21739,N_20322,N_18839);
or U21740 (N_21740,N_19402,N_18995);
and U21741 (N_21741,N_20226,N_18490);
xor U21742 (N_21742,N_20823,N_18523);
nor U21743 (N_21743,N_19982,N_18252);
and U21744 (N_21744,N_20683,N_20337);
and U21745 (N_21745,N_19980,N_18607);
nor U21746 (N_21746,N_18880,N_18675);
and U21747 (N_21747,N_20511,N_19452);
or U21748 (N_21748,N_19618,N_19736);
nor U21749 (N_21749,N_18805,N_19580);
and U21750 (N_21750,N_19653,N_18889);
nor U21751 (N_21751,N_19685,N_18865);
nand U21752 (N_21752,N_20798,N_19003);
xnor U21753 (N_21753,N_18498,N_20409);
or U21754 (N_21754,N_19362,N_18568);
nor U21755 (N_21755,N_19271,N_20211);
nand U21756 (N_21756,N_19262,N_18260);
nand U21757 (N_21757,N_19537,N_20318);
xor U21758 (N_21758,N_19480,N_18539);
xnor U21759 (N_21759,N_19352,N_18057);
nand U21760 (N_21760,N_19649,N_18006);
and U21761 (N_21761,N_20700,N_19811);
nor U21762 (N_21762,N_18403,N_19345);
nand U21763 (N_21763,N_19590,N_18258);
nand U21764 (N_21764,N_20212,N_19095);
nor U21765 (N_21765,N_18150,N_19377);
nor U21766 (N_21766,N_20940,N_18163);
nand U21767 (N_21767,N_20241,N_18242);
xor U21768 (N_21768,N_18097,N_19040);
and U21769 (N_21769,N_19732,N_20411);
and U21770 (N_21770,N_18357,N_18114);
or U21771 (N_21771,N_18398,N_18376);
or U21772 (N_21772,N_18976,N_19704);
xnor U21773 (N_21773,N_19551,N_20199);
or U21774 (N_21774,N_19357,N_20503);
nor U21775 (N_21775,N_20655,N_20190);
nand U21776 (N_21776,N_20876,N_18801);
xor U21777 (N_21777,N_19943,N_18044);
xor U21778 (N_21778,N_18535,N_19186);
or U21779 (N_21779,N_19840,N_18565);
nor U21780 (N_21780,N_19110,N_19018);
xor U21781 (N_21781,N_19343,N_20628);
and U21782 (N_21782,N_18070,N_20343);
nand U21783 (N_21783,N_18195,N_19386);
nand U21784 (N_21784,N_20282,N_18824);
and U21785 (N_21785,N_20198,N_18182);
nor U21786 (N_21786,N_18885,N_19571);
and U21787 (N_21787,N_18677,N_18950);
xor U21788 (N_21788,N_19906,N_19350);
or U21789 (N_21789,N_20403,N_20446);
nand U21790 (N_21790,N_19876,N_20426);
or U21791 (N_21791,N_20501,N_18790);
or U21792 (N_21792,N_19920,N_20658);
nor U21793 (N_21793,N_20489,N_20285);
nor U21794 (N_21794,N_20706,N_19488);
nand U21795 (N_21795,N_20656,N_20751);
nand U21796 (N_21796,N_19134,N_19560);
or U21797 (N_21797,N_19806,N_20526);
nand U21798 (N_21798,N_18153,N_19370);
nand U21799 (N_21799,N_18851,N_20562);
xnor U21800 (N_21800,N_19418,N_18399);
nor U21801 (N_21801,N_20475,N_19892);
and U21802 (N_21802,N_20753,N_18604);
nand U21803 (N_21803,N_19642,N_20171);
nor U21804 (N_21804,N_20577,N_18482);
and U21805 (N_21805,N_19543,N_19423);
nand U21806 (N_21806,N_20967,N_18672);
xor U21807 (N_21807,N_18402,N_19989);
and U21808 (N_21808,N_18872,N_19558);
or U21809 (N_21809,N_18155,N_20410);
or U21810 (N_21810,N_20336,N_20722);
nor U21811 (N_21811,N_18589,N_19280);
nand U21812 (N_21812,N_18939,N_19979);
nor U21813 (N_21813,N_20421,N_19167);
or U21814 (N_21814,N_20149,N_18086);
and U21815 (N_21815,N_19514,N_18203);
and U21816 (N_21816,N_19057,N_18977);
nor U21817 (N_21817,N_18570,N_19447);
nand U21818 (N_21818,N_19187,N_20907);
or U21819 (N_21819,N_19476,N_18981);
xnor U21820 (N_21820,N_20576,N_19267);
or U21821 (N_21821,N_20854,N_19559);
nand U21822 (N_21822,N_19006,N_18769);
nand U21823 (N_21823,N_18884,N_19644);
or U21824 (N_21824,N_20106,N_20231);
and U21825 (N_21825,N_18481,N_18115);
nor U21826 (N_21826,N_18983,N_20536);
and U21827 (N_21827,N_20500,N_18909);
xor U21828 (N_21828,N_18188,N_19419);
and U21829 (N_21829,N_20394,N_20039);
nand U21830 (N_21830,N_19053,N_20012);
or U21831 (N_21831,N_20731,N_20743);
xnor U21832 (N_21832,N_20518,N_19286);
or U21833 (N_21833,N_20660,N_18295);
and U21834 (N_21834,N_19938,N_18420);
nor U21835 (N_21835,N_20304,N_20926);
nand U21836 (N_21836,N_18379,N_19247);
xnor U21837 (N_21837,N_20745,N_18067);
or U21838 (N_21838,N_19331,N_18002);
or U21839 (N_21839,N_19165,N_18679);
nor U21840 (N_21840,N_20574,N_19759);
nor U21841 (N_21841,N_19605,N_18091);
and U21842 (N_21842,N_18577,N_18123);
xor U21843 (N_21843,N_20393,N_19087);
and U21844 (N_21844,N_20502,N_19056);
nand U21845 (N_21845,N_20910,N_18386);
or U21846 (N_21846,N_19783,N_20444);
xor U21847 (N_21847,N_18404,N_20081);
xnor U21848 (N_21848,N_19074,N_19014);
nand U21849 (N_21849,N_18066,N_20979);
and U21850 (N_21850,N_18867,N_20685);
nand U21851 (N_21851,N_20317,N_18991);
or U21852 (N_21852,N_20271,N_20217);
nor U21853 (N_21853,N_20551,N_18979);
nand U21854 (N_21854,N_18016,N_20917);
nand U21855 (N_21855,N_19849,N_20069);
nor U21856 (N_21856,N_18358,N_19709);
nand U21857 (N_21857,N_18823,N_19341);
nor U21858 (N_21858,N_18891,N_18117);
nand U21859 (N_21859,N_20928,N_18686);
or U21860 (N_21860,N_19281,N_19349);
xnor U21861 (N_21861,N_19278,N_18617);
or U21862 (N_21862,N_18967,N_19361);
or U21863 (N_21863,N_18317,N_20602);
xnor U21864 (N_21864,N_19518,N_18610);
or U21865 (N_21865,N_18833,N_18177);
nand U21866 (N_21866,N_19568,N_18670);
xnor U21867 (N_21867,N_18348,N_18953);
nor U21868 (N_21868,N_20328,N_18184);
or U21869 (N_21869,N_20777,N_19603);
nand U21870 (N_21870,N_19602,N_19191);
nand U21871 (N_21871,N_19140,N_20355);
xnor U21872 (N_21872,N_19403,N_19640);
or U21873 (N_21873,N_18056,N_19421);
and U21874 (N_21874,N_19695,N_18930);
and U21875 (N_21875,N_20699,N_18003);
or U21876 (N_21876,N_18010,N_18708);
nand U21877 (N_21877,N_18374,N_19387);
or U21878 (N_21878,N_20036,N_19525);
xnor U21879 (N_21879,N_19848,N_20933);
or U21880 (N_21880,N_20170,N_19123);
nand U21881 (N_21881,N_19405,N_19496);
nand U21882 (N_21882,N_18360,N_20817);
xor U21883 (N_21883,N_20566,N_20948);
or U21884 (N_21884,N_19160,N_18626);
and U21885 (N_21885,N_20011,N_18201);
nand U21886 (N_21886,N_19454,N_19681);
and U21887 (N_21887,N_20955,N_18492);
nand U21888 (N_21888,N_20498,N_20632);
nand U21889 (N_21889,N_19453,N_19067);
nor U21890 (N_21890,N_19701,N_18196);
and U21891 (N_21891,N_18106,N_18660);
or U21892 (N_21892,N_18985,N_18861);
nand U21893 (N_21893,N_18022,N_18603);
or U21894 (N_21894,N_18664,N_19449);
nor U21895 (N_21895,N_20053,N_20886);
or U21896 (N_21896,N_19241,N_19445);
nand U21897 (N_21897,N_18141,N_20607);
nand U21898 (N_21898,N_20760,N_18957);
or U21899 (N_21899,N_19358,N_20424);
xor U21900 (N_21900,N_18632,N_19096);
xnor U21901 (N_21901,N_19088,N_18248);
nor U21902 (N_21902,N_19270,N_18710);
xnor U21903 (N_21903,N_20793,N_18448);
xor U21904 (N_21904,N_18726,N_18844);
and U21905 (N_21905,N_18166,N_20287);
xnor U21906 (N_21906,N_18886,N_19430);
and U21907 (N_21907,N_20366,N_19600);
or U21908 (N_21908,N_19769,N_18324);
nand U21909 (N_21909,N_20599,N_20568);
nor U21910 (N_21910,N_18105,N_18546);
nand U21911 (N_21911,N_18781,N_18838);
nor U21912 (N_21912,N_20374,N_18578);
nor U21913 (N_21913,N_18712,N_18621);
nand U21914 (N_21914,N_20047,N_18778);
and U21915 (N_21915,N_18194,N_20096);
nor U21916 (N_21916,N_20941,N_18986);
nor U21917 (N_21917,N_20371,N_18602);
or U21918 (N_21918,N_20838,N_20668);
nand U21919 (N_21919,N_18651,N_18835);
or U21920 (N_21920,N_18239,N_19572);
and U21921 (N_21921,N_19945,N_19483);
or U21922 (N_21922,N_20540,N_18206);
or U21923 (N_21923,N_19188,N_18144);
nor U21924 (N_21924,N_20776,N_19502);
nand U21925 (N_21925,N_20877,N_18259);
xor U21926 (N_21926,N_18913,N_19498);
nand U21927 (N_21927,N_18502,N_19974);
and U21928 (N_21928,N_18035,N_20969);
and U21929 (N_21929,N_20819,N_19245);
nand U21930 (N_21930,N_18811,N_18232);
nand U21931 (N_21931,N_20652,N_20327);
xnor U21932 (N_21932,N_19310,N_18768);
xor U21933 (N_21933,N_18717,N_18720);
xor U21934 (N_21934,N_19874,N_20718);
or U21935 (N_21935,N_19700,N_19935);
nor U21936 (N_21936,N_18937,N_19636);
xnor U21937 (N_21937,N_19082,N_20815);
nor U21938 (N_21938,N_19791,N_20164);
or U21939 (N_21939,N_20914,N_20924);
xor U21940 (N_21940,N_19497,N_19252);
nor U21941 (N_21941,N_20710,N_20184);
nor U21942 (N_21942,N_19043,N_19632);
nand U21943 (N_21943,N_19171,N_19000);
and U21944 (N_21944,N_18984,N_19986);
nor U21945 (N_21945,N_18304,N_18658);
xnor U21946 (N_21946,N_18753,N_19677);
nor U21947 (N_21947,N_19204,N_19639);
or U21948 (N_21948,N_20453,N_20992);
nand U21949 (N_21949,N_18170,N_18959);
and U21950 (N_21950,N_20215,N_20239);
xor U21951 (N_21951,N_19727,N_20052);
nor U21952 (N_21952,N_19773,N_18684);
nand U21953 (N_21953,N_19004,N_19075);
or U21954 (N_21954,N_18120,N_20033);
nor U21955 (N_21955,N_20585,N_19373);
and U21956 (N_21956,N_19667,N_20479);
xnor U21957 (N_21957,N_19285,N_20856);
and U21958 (N_21958,N_20438,N_19212);
or U21959 (N_21959,N_18911,N_19034);
and U21960 (N_21960,N_19705,N_18473);
and U21961 (N_21961,N_18516,N_19244);
xor U21962 (N_21962,N_19721,N_20649);
and U21963 (N_21963,N_19492,N_19105);
and U21964 (N_21964,N_20925,N_20265);
xnor U21965 (N_21965,N_20752,N_20665);
nor U21966 (N_21966,N_18284,N_20804);
and U21967 (N_21967,N_19934,N_20621);
nor U21968 (N_21968,N_19504,N_18207);
xnor U21969 (N_21969,N_19507,N_20989);
or U21970 (N_21970,N_18849,N_20726);
nand U21971 (N_21971,N_19961,N_18549);
nor U21972 (N_21972,N_18134,N_20059);
xor U21973 (N_21973,N_19078,N_18588);
nand U21974 (N_21974,N_18520,N_19939);
and U21975 (N_21975,N_18249,N_19796);
or U21976 (N_21976,N_18005,N_18275);
and U21977 (N_21977,N_20441,N_18219);
xnor U21978 (N_21978,N_19399,N_19589);
nand U21979 (N_21979,N_20017,N_20020);
and U21980 (N_21980,N_20724,N_20758);
nor U21981 (N_21981,N_18283,N_19627);
xnor U21982 (N_21982,N_19666,N_18417);
and U21983 (N_21983,N_18740,N_18414);
nor U21984 (N_21984,N_20651,N_19231);
nor U21985 (N_21985,N_20895,N_19847);
nand U21986 (N_21986,N_20058,N_20064);
or U21987 (N_21987,N_18692,N_20100);
xor U21988 (N_21988,N_19199,N_20376);
nand U21989 (N_21989,N_20027,N_20539);
nand U21990 (N_21990,N_20122,N_19381);
nor U21991 (N_21991,N_18346,N_20404);
nor U21992 (N_21992,N_20477,N_20153);
nand U21993 (N_21993,N_20578,N_19792);
nor U21994 (N_21994,N_20546,N_19250);
nand U21995 (N_21995,N_18732,N_19462);
and U21996 (N_21996,N_19985,N_20381);
or U21997 (N_21997,N_19193,N_18591);
or U21998 (N_21998,N_18764,N_19575);
nor U21999 (N_21999,N_18245,N_19660);
and U22000 (N_22000,N_20103,N_18095);
nor U22001 (N_22001,N_18335,N_18455);
or U22002 (N_22002,N_19200,N_19856);
nand U22003 (N_22003,N_19609,N_20281);
xor U22004 (N_22004,N_20151,N_18992);
nor U22005 (N_22005,N_18898,N_20564);
and U22006 (N_22006,N_19128,N_20583);
nand U22007 (N_22007,N_18344,N_18431);
nand U22008 (N_22008,N_18585,N_18209);
and U22009 (N_22009,N_19022,N_18706);
or U22010 (N_22010,N_18318,N_19898);
nand U22011 (N_22011,N_18139,N_18238);
nor U22012 (N_22012,N_20484,N_18004);
nand U22013 (N_22013,N_20024,N_19991);
or U22014 (N_22014,N_19017,N_19977);
nand U22015 (N_22015,N_18340,N_19706);
nor U22016 (N_22016,N_20755,N_18138);
or U22017 (N_22017,N_18461,N_20788);
or U22018 (N_22018,N_18076,N_19916);
or U22019 (N_22019,N_20319,N_20654);
and U22020 (N_22020,N_18784,N_18334);
or U22021 (N_22021,N_19391,N_20251);
nor U22022 (N_22022,N_20320,N_18703);
or U22023 (N_22023,N_20717,N_18445);
nand U22024 (N_22024,N_19965,N_19686);
or U22025 (N_22025,N_18277,N_18980);
nor U22026 (N_22026,N_18287,N_19459);
nand U22027 (N_22027,N_19914,N_19888);
nand U22028 (N_22028,N_19601,N_20889);
nor U22029 (N_22029,N_18965,N_18631);
xor U22030 (N_22030,N_18634,N_19062);
xnor U22031 (N_22031,N_18234,N_18341);
xnor U22032 (N_22032,N_20901,N_19065);
or U22033 (N_22033,N_19433,N_19953);
nor U22034 (N_22034,N_20124,N_19718);
or U22035 (N_22035,N_20613,N_20913);
nand U22036 (N_22036,N_19059,N_19473);
xor U22037 (N_22037,N_19532,N_18116);
xnor U22038 (N_22038,N_18447,N_18148);
nand U22039 (N_22039,N_18012,N_18480);
or U22040 (N_22040,N_19970,N_19414);
nor U22041 (N_22041,N_19174,N_19290);
nor U22042 (N_22042,N_18500,N_19179);
nor U22043 (N_22043,N_19790,N_18048);
nand U22044 (N_22044,N_20504,N_18327);
or U22045 (N_22045,N_20734,N_18338);
or U22046 (N_22046,N_20783,N_19055);
or U22047 (N_22047,N_20624,N_19860);
xnor U22048 (N_22048,N_20268,N_18302);
nand U22049 (N_22049,N_19859,N_20119);
and U22050 (N_22050,N_18364,N_19071);
nor U22051 (N_22051,N_19209,N_19768);
nor U22052 (N_22052,N_18776,N_19092);
xor U22053 (N_22053,N_20189,N_20853);
xnor U22054 (N_22054,N_19242,N_19340);
xnor U22055 (N_22055,N_20026,N_19379);
and U22056 (N_22056,N_20620,N_20290);
nand U22057 (N_22057,N_20871,N_19540);
or U22058 (N_22058,N_20238,N_18655);
or U22059 (N_22059,N_18586,N_18092);
and U22060 (N_22060,N_20139,N_20837);
or U22061 (N_22061,N_20255,N_18932);
nand U22062 (N_22062,N_20807,N_18596);
xnor U22063 (N_22063,N_19795,N_18359);
xnor U22064 (N_22064,N_18084,N_19505);
nand U22065 (N_22065,N_20389,N_18216);
or U22066 (N_22066,N_18858,N_18142);
nor U22067 (N_22067,N_18087,N_20617);
nand U22068 (N_22068,N_18037,N_19839);
xnor U22069 (N_22069,N_18271,N_19670);
nand U22070 (N_22070,N_18416,N_20032);
xor U22071 (N_22071,N_20523,N_20288);
nor U22072 (N_22072,N_20701,N_19533);
and U22073 (N_22073,N_18647,N_19020);
or U22074 (N_22074,N_18582,N_18494);
and U22075 (N_22075,N_19592,N_19633);
xnor U22076 (N_22076,N_19076,N_19330);
or U22077 (N_22077,N_18648,N_18315);
or U22078 (N_22078,N_18221,N_19486);
or U22079 (N_22079,N_18476,N_18405);
and U22080 (N_22080,N_19915,N_20449);
and U22081 (N_22081,N_18225,N_20532);
and U22082 (N_22082,N_18543,N_18936);
and U22083 (N_22083,N_20930,N_19124);
and U22084 (N_22084,N_19782,N_20761);
and U22085 (N_22085,N_18892,N_20127);
xor U22086 (N_22086,N_18164,N_18934);
xnor U22087 (N_22087,N_20584,N_18297);
nand U22088 (N_22088,N_19521,N_18552);
or U22089 (N_22089,N_20524,N_20178);
xnor U22090 (N_22090,N_20143,N_19904);
or U22091 (N_22091,N_20890,N_19254);
or U22092 (N_22092,N_19902,N_18728);
and U22093 (N_22093,N_19978,N_19881);
xor U22094 (N_22094,N_20736,N_18606);
xor U22095 (N_22095,N_19932,N_19001);
xnor U22096 (N_22096,N_18296,N_19995);
or U22097 (N_22097,N_18286,N_19372);
and U22098 (N_22098,N_20482,N_20920);
nand U22099 (N_22099,N_19173,N_20883);
nor U22100 (N_22100,N_19102,N_18059);
xnor U22101 (N_22101,N_18167,N_20677);
xnor U22102 (N_22102,N_18931,N_19786);
xnor U22103 (N_22103,N_18131,N_19930);
nor U22104 (N_22104,N_19997,N_19581);
and U22105 (N_22105,N_19091,N_20797);
or U22106 (N_22106,N_18024,N_20302);
or U22107 (N_22107,N_20912,N_18969);
nand U22108 (N_22108,N_19308,N_20600);
xnor U22109 (N_22109,N_20465,N_19274);
nand U22110 (N_22110,N_19725,N_19318);
nor U22111 (N_22111,N_19690,N_19298);
or U22112 (N_22112,N_19440,N_19682);
nor U22113 (N_22113,N_20209,N_18320);
nor U22114 (N_22114,N_18594,N_19464);
and U22115 (N_22115,N_20382,N_19556);
or U22116 (N_22116,N_20802,N_19668);
or U22117 (N_22117,N_18488,N_20868);
and U22118 (N_22118,N_19546,N_20786);
nor U22119 (N_22119,N_19987,N_19166);
and U22120 (N_22120,N_19328,N_18369);
and U22121 (N_22121,N_20733,N_20110);
or U22122 (N_22122,N_18151,N_18982);
and U22123 (N_22123,N_20387,N_18707);
or U22124 (N_22124,N_19313,N_20545);
nor U22125 (N_22125,N_20385,N_20627);
and U22126 (N_22126,N_18918,N_20060);
xor U22127 (N_22127,N_20814,N_20648);
xnor U22128 (N_22128,N_18816,N_18293);
and U22129 (N_22129,N_18871,N_19107);
nand U22130 (N_22130,N_20681,N_20423);
and U22131 (N_22131,N_20061,N_19534);
xor U22132 (N_22132,N_18393,N_18601);
or U22133 (N_22133,N_18739,N_20666);
or U22134 (N_22134,N_20222,N_19494);
xnor U22135 (N_22135,N_20262,N_19356);
and U22136 (N_22136,N_19469,N_19321);
nor U22137 (N_22137,N_20422,N_19687);
and U22138 (N_22138,N_20270,N_18812);
or U22139 (N_22139,N_19481,N_18089);
nor U22140 (N_22140,N_20944,N_18656);
nor U22141 (N_22141,N_18233,N_20878);
or U22142 (N_22142,N_19041,N_20144);
xnor U22143 (N_22143,N_18125,N_20898);
xor U22144 (N_22144,N_20367,N_18093);
nor U22145 (N_22145,N_19228,N_20897);
nor U22146 (N_22146,N_19665,N_18807);
nor U22147 (N_22147,N_20451,N_18169);
or U22148 (N_22148,N_19952,N_20079);
nor U22149 (N_22149,N_20647,N_19136);
nand U22150 (N_22150,N_18727,N_19052);
nor U22151 (N_22151,N_19266,N_20639);
xor U22152 (N_22152,N_19084,N_19233);
xnor U22153 (N_22153,N_18179,N_19548);
xnor U22154 (N_22154,N_19646,N_18896);
xnor U22155 (N_22155,N_20041,N_20663);
xor U22156 (N_22156,N_18366,N_20264);
nor U22157 (N_22157,N_19146,N_18755);
nand U22158 (N_22158,N_19645,N_18863);
and U22159 (N_22159,N_20025,N_18434);
and U22160 (N_22160,N_19884,N_19517);
or U22161 (N_22161,N_18963,N_19007);
and U22162 (N_22162,N_18415,N_20162);
nor U22163 (N_22163,N_18406,N_20507);
xor U22164 (N_22164,N_18400,N_20105);
and U22165 (N_22165,N_20077,N_20631);
xor U22166 (N_22166,N_20252,N_20147);
and U22167 (N_22167,N_19651,N_20556);
or U22168 (N_22168,N_18467,N_19112);
and U22169 (N_22169,N_20984,N_20636);
and U22170 (N_22170,N_20770,N_20292);
and U22171 (N_22171,N_18548,N_18700);
and U22172 (N_22172,N_20107,N_19619);
nor U22173 (N_22173,N_19911,N_19957);
or U22174 (N_22174,N_20630,N_18945);
xor U22175 (N_22175,N_18290,N_20748);
or U22176 (N_22176,N_20864,N_20552);
xor U22177 (N_22177,N_19750,N_19289);
nand U22178 (N_22178,N_18058,N_18454);
nand U22179 (N_22179,N_20708,N_19283);
nand U22180 (N_22180,N_20569,N_19913);
nand U22181 (N_22181,N_20452,N_18412);
xor U22182 (N_22182,N_18486,N_20847);
xor U22183 (N_22183,N_19042,N_18592);
or U22184 (N_22184,N_19910,N_19944);
nand U22185 (N_22185,N_19264,N_18550);
and U22186 (N_22186,N_18701,N_19990);
and U22187 (N_22187,N_19400,N_20010);
xor U22188 (N_22188,N_19248,N_18343);
nand U22189 (N_22189,N_19867,N_20272);
or U22190 (N_22190,N_19947,N_19153);
or U22191 (N_22191,N_20791,N_19550);
xor U22192 (N_22192,N_19756,N_19432);
xor U22193 (N_22193,N_20312,N_18326);
nor U22194 (N_22194,N_19049,N_19615);
nor U22195 (N_22195,N_19027,N_20015);
nor U22196 (N_22196,N_18288,N_19530);
xor U22197 (N_22197,N_18541,N_19858);
nor U22198 (N_22198,N_18668,N_20450);
nor U22199 (N_22199,N_18879,N_20099);
xor U22200 (N_22200,N_18171,N_20396);
nor U22201 (N_22201,N_18754,N_20361);
nand U22202 (N_22202,N_20260,N_20567);
or U22203 (N_22203,N_19570,N_19035);
xor U22204 (N_22204,N_20742,N_19263);
xor U22205 (N_22205,N_19678,N_18319);
nor U22206 (N_22206,N_20185,N_18020);
or U22207 (N_22207,N_18826,N_20116);
nor U22208 (N_22208,N_18765,N_20054);
nand U22209 (N_22209,N_18250,N_18785);
nor U22210 (N_22210,N_19069,N_18316);
xor U22211 (N_22211,N_18920,N_19393);
or U22212 (N_22212,N_19021,N_19276);
or U22213 (N_22213,N_18571,N_19279);
nor U22214 (N_22214,N_19897,N_18060);
and U22215 (N_22215,N_18662,N_20101);
and U22216 (N_22216,N_20531,N_18935);
and U22217 (N_22217,N_20460,N_20594);
or U22218 (N_22218,N_19269,N_20606);
and U22219 (N_22219,N_19383,N_20085);
xnor U22220 (N_22220,N_18424,N_20166);
nand U22221 (N_22221,N_18075,N_18917);
nand U22222 (N_22222,N_19804,N_18921);
and U22223 (N_22223,N_18189,N_19133);
nor U22224 (N_22224,N_19311,N_20214);
and U22225 (N_22225,N_19236,N_19652);
and U22226 (N_22226,N_19710,N_19416);
nor U22227 (N_22227,N_19104,N_19820);
nor U22228 (N_22228,N_18464,N_20549);
and U22229 (N_22229,N_18228,N_19028);
nand U22230 (N_22230,N_18168,N_18333);
xor U22231 (N_22231,N_18678,N_18477);
xor U22232 (N_22232,N_20022,N_18777);
nor U22233 (N_22233,N_18387,N_18023);
and U22234 (N_22234,N_19458,N_20619);
or U22235 (N_22235,N_18501,N_20463);
nor U22236 (N_22236,N_18172,N_19093);
xnor U22237 (N_22237,N_19578,N_18876);
xor U22238 (N_22238,N_19323,N_18479);
and U22239 (N_22239,N_19917,N_19692);
nand U22240 (N_22240,N_18558,N_20732);
nand U22241 (N_22241,N_19703,N_19748);
and U22242 (N_22242,N_20988,N_20402);
nand U22243 (N_22243,N_18077,N_18532);
and U22244 (N_22244,N_19325,N_20044);
nand U22245 (N_22245,N_18423,N_20996);
xnor U22246 (N_22246,N_18220,N_18050);
or U22247 (N_22247,N_19338,N_18888);
xor U22248 (N_22248,N_20400,N_19865);
or U22249 (N_22249,N_19442,N_18038);
xnor U22250 (N_22250,N_19694,N_20953);
or U22251 (N_22251,N_19616,N_19068);
or U22252 (N_22252,N_20201,N_19138);
xor U22253 (N_22253,N_20420,N_19152);
xor U22254 (N_22254,N_19477,N_18236);
nor U22255 (N_22255,N_20951,N_18489);
or U22256 (N_22256,N_18519,N_19815);
or U22257 (N_22257,N_18162,N_18667);
nor U22258 (N_22258,N_20159,N_19457);
or U22259 (N_22259,N_19210,N_20520);
nor U22260 (N_22260,N_18681,N_19538);
nor U22261 (N_22261,N_18478,N_19513);
nand U22262 (N_22262,N_18987,N_19509);
nor U22263 (N_22263,N_18771,N_20529);
nand U22264 (N_22264,N_20813,N_18132);
or U22265 (N_22265,N_20591,N_20822);
xor U22266 (N_22266,N_20245,N_19918);
and U22267 (N_22267,N_19647,N_19090);
xnor U22268 (N_22268,N_19674,N_20333);
nor U22269 (N_22269,N_18762,N_18487);
xnor U22270 (N_22270,N_20016,N_20196);
nand U22271 (N_22271,N_18733,N_19385);
nand U22272 (N_22272,N_20855,N_18695);
xor U22273 (N_22273,N_18813,N_19536);
or U22274 (N_22274,N_20496,N_20121);
nor U22275 (N_22275,N_20671,N_18635);
xnor U22276 (N_22276,N_20307,N_18140);
nor U22277 (N_22277,N_18999,N_20762);
nand U22278 (N_22278,N_19557,N_19676);
and U22279 (N_22279,N_19671,N_18682);
nor U22280 (N_22280,N_20156,N_20937);
nor U22281 (N_22281,N_20362,N_19036);
and U22282 (N_22282,N_20884,N_19151);
xor U22283 (N_22283,N_19463,N_20714);
xor U22284 (N_22284,N_19202,N_20197);
nor U22285 (N_22285,N_19925,N_19129);
or U22286 (N_22286,N_20747,N_19284);
nor U22287 (N_22287,N_18508,N_19287);
or U22288 (N_22288,N_20916,N_20225);
or U22289 (N_22289,N_18694,N_18751);
nand U22290 (N_22290,N_19127,N_18661);
or U22291 (N_22291,N_19435,N_18495);
xor U22292 (N_22292,N_20563,N_20618);
nor U22293 (N_22293,N_20522,N_20839);
xnor U22294 (N_22294,N_18923,N_18608);
nand U22295 (N_22295,N_18191,N_20927);
nor U22296 (N_22296,N_20678,N_19319);
xor U22297 (N_22297,N_20442,N_18254);
or U22298 (N_22298,N_20888,N_19882);
xnor U22299 (N_22299,N_18074,N_18742);
nand U22300 (N_22300,N_20305,N_19080);
nand U22301 (N_22301,N_19999,N_20368);
or U22302 (N_22302,N_20431,N_19937);
nor U22303 (N_22303,N_18966,N_18599);
xor U22304 (N_22304,N_18564,N_18261);
and U22305 (N_22305,N_18362,N_18098);
nor U22306 (N_22306,N_18096,N_19838);
nor U22307 (N_22307,N_19844,N_19348);
and U22308 (N_22308,N_19693,N_19259);
or U22309 (N_22309,N_20859,N_19064);
xnor U22310 (N_22310,N_18878,N_19921);
nor U22311 (N_22311,N_18687,N_18511);
nor U22312 (N_22312,N_19030,N_18419);
nor U22313 (N_22313,N_19728,N_18154);
nor U22314 (N_22314,N_20408,N_18180);
nor U22315 (N_22315,N_18547,N_20350);
or U22316 (N_22316,N_20458,N_19717);
or U22317 (N_22317,N_18146,N_20548);
and U22318 (N_22318,N_20643,N_20335);
nor U22319 (N_22319,N_18394,N_19047);
xnor U22320 (N_22320,N_20971,N_19620);
and U22321 (N_22321,N_20067,N_18130);
nand U22322 (N_22322,N_18231,N_20769);
nor U22323 (N_22323,N_20301,N_20347);
and U22324 (N_22324,N_20687,N_19797);
and U22325 (N_22325,N_19214,N_19928);
or U22326 (N_22326,N_20437,N_18545);
or U22327 (N_22327,N_19031,N_18531);
and U22328 (N_22328,N_19657,N_18378);
xor U22329 (N_22329,N_20869,N_20279);
nor U22330 (N_22330,N_20034,N_19023);
or U22331 (N_22331,N_18165,N_20541);
or U22332 (N_22332,N_19229,N_18039);
and U22333 (N_22333,N_20781,N_19614);
and U22334 (N_22334,N_20340,N_19752);
and U22335 (N_22335,N_19960,N_20488);
xor U22336 (N_22336,N_20612,N_19369);
and U22337 (N_22337,N_18426,N_18342);
xor U22338 (N_22338,N_19761,N_20263);
or U22339 (N_22339,N_20165,N_20923);
and U22340 (N_22340,N_20076,N_20210);
or U22341 (N_22341,N_18810,N_19428);
or U22342 (N_22342,N_19159,N_19591);
nor U22343 (N_22343,N_20991,N_19232);
or U22344 (N_22344,N_20202,N_18202);
or U22345 (N_22345,N_19630,N_19101);
or U22346 (N_22346,N_18435,N_20314);
nand U22347 (N_22347,N_20865,N_20094);
xor U22348 (N_22348,N_20481,N_19230);
and U22349 (N_22349,N_19675,N_18397);
nand U22350 (N_22350,N_18506,N_18702);
or U22351 (N_22351,N_19142,N_19139);
or U22352 (N_22352,N_18065,N_18772);
nand U22353 (N_22353,N_18009,N_18914);
or U22354 (N_22354,N_18837,N_19801);
nand U22355 (N_22355,N_19516,N_20348);
or U22356 (N_22356,N_18186,N_18628);
and U22357 (N_22357,N_19500,N_19503);
or U22358 (N_22358,N_18266,N_18803);
nor U22359 (N_22359,N_20457,N_18916);
nand U22360 (N_22360,N_20179,N_18683);
xor U22361 (N_22361,N_18127,N_18313);
xor U22362 (N_22362,N_20259,N_18208);
xnor U22363 (N_22363,N_18988,N_18053);
nor U22364 (N_22364,N_20841,N_18590);
nand U22365 (N_22365,N_19894,N_20790);
and U22366 (N_22366,N_18852,N_19813);
nor U22367 (N_22367,N_20109,N_20554);
nor U22368 (N_22368,N_19005,N_19563);
nand U22369 (N_22369,N_20021,N_20945);
xor U22370 (N_22370,N_18085,N_20428);
or U22371 (N_22371,N_19077,N_19711);
or U22372 (N_22372,N_18696,N_19114);
xor U22373 (N_22373,N_18644,N_19512);
nand U22374 (N_22374,N_19829,N_20642);
nor U22375 (N_22375,N_19887,N_18783);
or U22376 (N_22376,N_19648,N_19132);
and U22377 (N_22377,N_18817,N_20784);
and U22378 (N_22378,N_18522,N_20809);
or U22379 (N_22379,N_18924,N_20480);
or U22380 (N_22380,N_18069,N_18946);
nand U22381 (N_22381,N_18331,N_20092);
and U22382 (N_22382,N_20960,N_20537);
xor U22383 (N_22383,N_20213,N_19116);
nor U22384 (N_22384,N_19658,N_18204);
xnor U22385 (N_22385,N_20987,N_20074);
and U22386 (N_22386,N_18439,N_20051);
or U22387 (N_22387,N_20087,N_20954);
or U22388 (N_22388,N_19971,N_20068);
nor U22389 (N_22389,N_20693,N_20236);
nand U22390 (N_22390,N_19148,N_20816);
nand U22391 (N_22391,N_18798,N_19227);
nand U22392 (N_22392,N_20759,N_20045);
nand U22393 (N_22393,N_19629,N_18158);
xnor U22394 (N_22394,N_18090,N_19424);
or U22395 (N_22395,N_20640,N_20031);
and U22396 (N_22396,N_18080,N_19194);
and U22397 (N_22397,N_19983,N_19779);
nor U22398 (N_22398,N_18352,N_20581);
nand U22399 (N_22399,N_18512,N_20134);
or U22400 (N_22400,N_20891,N_18912);
nand U22401 (N_22401,N_19885,N_19316);
and U22402 (N_22402,N_20247,N_20931);
nand U22403 (N_22403,N_18497,N_19582);
nor U22404 (N_22404,N_19119,N_20018);
and U22405 (N_22405,N_20588,N_19702);
nor U22406 (N_22406,N_19221,N_18989);
nand U22407 (N_22407,N_19622,N_18373);
xnor U22408 (N_22408,N_19472,N_18927);
or U22409 (N_22409,N_20825,N_19213);
nand U22410 (N_22410,N_19565,N_20177);
or U22411 (N_22411,N_18905,N_18027);
xnor U22412 (N_22412,N_19851,N_19141);
xnor U22413 (N_22413,N_20661,N_18808);
and U22414 (N_22414,N_20763,N_20029);
and U22415 (N_22415,N_18744,N_20158);
or U22416 (N_22416,N_20466,N_19956);
nor U22417 (N_22417,N_18407,N_20140);
and U22418 (N_22418,N_20505,N_20136);
nor U22419 (N_22419,N_18901,N_18214);
or U22420 (N_22420,N_18272,N_20383);
nor U22421 (N_22421,N_20746,N_18544);
and U22422 (N_22422,N_18722,N_18321);
nor U22423 (N_22423,N_20230,N_18625);
xnor U22424 (N_22424,N_20694,N_20395);
or U22425 (N_22425,N_18237,N_18336);
nor U22426 (N_22426,N_20867,N_20741);
xor U22427 (N_22427,N_18391,N_18862);
xnor U22428 (N_22428,N_20415,N_19545);
or U22429 (N_22429,N_18049,N_19220);
and U22430 (N_22430,N_19764,N_20332);
nand U22431 (N_22431,N_19576,N_20254);
and U22432 (N_22432,N_20205,N_20216);
nand U22433 (N_22433,N_19439,N_19787);
nand U22434 (N_22434,N_19655,N_19715);
nand U22435 (N_22435,N_19288,N_19100);
and U22436 (N_22436,N_19817,N_19749);
xor U22437 (N_22437,N_18786,N_19196);
or U22438 (N_22438,N_18645,N_18735);
xor U22439 (N_22439,N_18451,N_20456);
nor U22440 (N_22440,N_18160,N_18217);
nor U22441 (N_22441,N_18305,N_18064);
xor U22442 (N_22442,N_20001,N_18779);
nand U22443 (N_22443,N_19767,N_18227);
and U22444 (N_22444,N_20686,N_18866);
nor U22445 (N_22445,N_18222,N_18525);
and U22446 (N_22446,N_20662,N_19522);
xnor U22447 (N_22447,N_20372,N_20440);
or U22448 (N_22448,N_19103,N_18615);
or U22449 (N_22449,N_19029,N_19465);
or U22450 (N_22450,N_18112,N_19155);
and U22451 (N_22451,N_18396,N_19456);
or U22452 (N_22452,N_19873,N_18598);
or U22453 (N_22453,N_19326,N_18241);
nand U22454 (N_22454,N_19780,N_20363);
nor U22455 (N_22455,N_18147,N_19025);
or U22456 (N_22456,N_19150,N_20679);
or U22457 (N_22457,N_18693,N_18743);
nand U22458 (N_22458,N_19929,N_18566);
nor U22459 (N_22459,N_19058,N_20592);
nor U22460 (N_22460,N_19485,N_19599);
xnor U22461 (N_22461,N_18994,N_20188);
nand U22462 (N_22462,N_20866,N_19836);
nor U22463 (N_22463,N_20615,N_19566);
nor U22464 (N_22464,N_20228,N_19368);
or U22465 (N_22465,N_18094,N_20557);
or U22466 (N_22466,N_19588,N_20249);
nor U22467 (N_22467,N_18368,N_20832);
nor U22468 (N_22468,N_20659,N_19842);
xnor U22469 (N_22469,N_19478,N_18370);
or U22470 (N_22470,N_20806,N_20309);
xnor U22471 (N_22471,N_19506,N_19246);
or U22472 (N_22472,N_19177,N_18780);
and U22473 (N_22473,N_20533,N_18951);
nor U22474 (N_22474,N_20075,N_20377);
and U22475 (N_22475,N_18633,N_19009);
nand U22476 (N_22476,N_18355,N_20406);
or U22477 (N_22477,N_20278,N_18363);
nor U22478 (N_22478,N_20004,N_19389);
nor U22479 (N_22479,N_18990,N_20104);
xnor U22480 (N_22480,N_20598,N_19719);
and U22481 (N_22481,N_19097,N_19772);
nor U22482 (N_22482,N_20509,N_20286);
or U22483 (N_22483,N_19162,N_18834);
nand U22484 (N_22484,N_19218,N_19239);
or U22485 (N_22485,N_19351,N_19216);
nor U22486 (N_22486,N_20704,N_19257);
and U22487 (N_22487,N_18280,N_19872);
nor U22488 (N_22488,N_18699,N_19734);
nand U22489 (N_22489,N_18298,N_19217);
or U22490 (N_22490,N_19237,N_19163);
nand U22491 (N_22491,N_20728,N_19696);
xnor U22492 (N_22492,N_19758,N_19258);
or U22493 (N_22493,N_19922,N_20294);
and U22494 (N_22494,N_18600,N_20349);
nor U22495 (N_22495,N_19729,N_19698);
xnor U22496 (N_22496,N_20043,N_19745);
or U22497 (N_22497,N_19819,N_20310);
xnor U22498 (N_22498,N_19317,N_20974);
nand U22499 (N_22499,N_20218,N_18630);
xnor U22500 (N_22500,N_20144,N_20073);
nand U22501 (N_22501,N_19656,N_19052);
nor U22502 (N_22502,N_18561,N_20083);
and U22503 (N_22503,N_18224,N_19151);
xnor U22504 (N_22504,N_19159,N_20051);
nand U22505 (N_22505,N_19590,N_19967);
nor U22506 (N_22506,N_18585,N_20197);
and U22507 (N_22507,N_20259,N_19215);
or U22508 (N_22508,N_18351,N_20178);
and U22509 (N_22509,N_18845,N_20293);
and U22510 (N_22510,N_18933,N_19342);
or U22511 (N_22511,N_18527,N_19071);
or U22512 (N_22512,N_19247,N_18763);
and U22513 (N_22513,N_19670,N_19978);
nand U22514 (N_22514,N_18563,N_18117);
nor U22515 (N_22515,N_18641,N_18940);
and U22516 (N_22516,N_20584,N_19752);
or U22517 (N_22517,N_20157,N_19657);
nor U22518 (N_22518,N_20440,N_18859);
and U22519 (N_22519,N_20088,N_20823);
nor U22520 (N_22520,N_20768,N_18595);
xor U22521 (N_22521,N_18537,N_19788);
nor U22522 (N_22522,N_20855,N_18382);
or U22523 (N_22523,N_20502,N_20545);
nor U22524 (N_22524,N_18582,N_18007);
xor U22525 (N_22525,N_20332,N_20081);
or U22526 (N_22526,N_18141,N_19695);
and U22527 (N_22527,N_20130,N_19584);
nor U22528 (N_22528,N_19861,N_20401);
nand U22529 (N_22529,N_19547,N_18131);
nor U22530 (N_22530,N_20371,N_20408);
nor U22531 (N_22531,N_19153,N_19392);
and U22532 (N_22532,N_19337,N_19045);
nand U22533 (N_22533,N_19927,N_18670);
and U22534 (N_22534,N_19501,N_18249);
and U22535 (N_22535,N_20642,N_18995);
nand U22536 (N_22536,N_20814,N_20374);
xnor U22537 (N_22537,N_19573,N_20260);
nor U22538 (N_22538,N_20483,N_18968);
xor U22539 (N_22539,N_20788,N_20466);
nand U22540 (N_22540,N_19679,N_20776);
and U22541 (N_22541,N_20140,N_18692);
xnor U22542 (N_22542,N_20567,N_19091);
xor U22543 (N_22543,N_19542,N_19702);
or U22544 (N_22544,N_18832,N_20008);
or U22545 (N_22545,N_19444,N_18815);
or U22546 (N_22546,N_18545,N_19611);
or U22547 (N_22547,N_20072,N_18963);
and U22548 (N_22548,N_19041,N_20162);
or U22549 (N_22549,N_19481,N_18907);
nand U22550 (N_22550,N_19179,N_18568);
nor U22551 (N_22551,N_19148,N_19498);
and U22552 (N_22552,N_18242,N_20615);
nand U22553 (N_22553,N_19420,N_18703);
or U22554 (N_22554,N_20899,N_20401);
and U22555 (N_22555,N_19300,N_19509);
xnor U22556 (N_22556,N_19232,N_18555);
nand U22557 (N_22557,N_18141,N_20380);
nand U22558 (N_22558,N_19134,N_18671);
and U22559 (N_22559,N_18156,N_19480);
or U22560 (N_22560,N_19477,N_19341);
xnor U22561 (N_22561,N_19063,N_18438);
and U22562 (N_22562,N_19032,N_19215);
xnor U22563 (N_22563,N_19106,N_20466);
xor U22564 (N_22564,N_18876,N_19325);
and U22565 (N_22565,N_19761,N_20975);
or U22566 (N_22566,N_18235,N_20082);
and U22567 (N_22567,N_18186,N_18939);
and U22568 (N_22568,N_19813,N_19708);
and U22569 (N_22569,N_20032,N_19395);
nor U22570 (N_22570,N_20661,N_18880);
nand U22571 (N_22571,N_20762,N_20690);
xnor U22572 (N_22572,N_18728,N_18163);
nand U22573 (N_22573,N_18402,N_20918);
xor U22574 (N_22574,N_19374,N_20989);
nand U22575 (N_22575,N_18796,N_18303);
nand U22576 (N_22576,N_18422,N_20325);
nor U22577 (N_22577,N_20964,N_18914);
xnor U22578 (N_22578,N_18924,N_19805);
or U22579 (N_22579,N_19266,N_20345);
or U22580 (N_22580,N_20920,N_19495);
xor U22581 (N_22581,N_18662,N_20977);
and U22582 (N_22582,N_19062,N_20534);
or U22583 (N_22583,N_20208,N_20035);
nand U22584 (N_22584,N_19841,N_19477);
and U22585 (N_22585,N_19708,N_19886);
or U22586 (N_22586,N_19345,N_18363);
nand U22587 (N_22587,N_20999,N_18931);
nor U22588 (N_22588,N_19118,N_18561);
xor U22589 (N_22589,N_18471,N_19083);
or U22590 (N_22590,N_19747,N_18737);
nor U22591 (N_22591,N_20443,N_20968);
or U22592 (N_22592,N_20233,N_20728);
and U22593 (N_22593,N_20276,N_18722);
nor U22594 (N_22594,N_19114,N_19238);
and U22595 (N_22595,N_19886,N_18244);
nand U22596 (N_22596,N_19256,N_18891);
nor U22597 (N_22597,N_18687,N_19810);
xnor U22598 (N_22598,N_20347,N_18256);
xor U22599 (N_22599,N_18634,N_19602);
nand U22600 (N_22600,N_18493,N_19142);
and U22601 (N_22601,N_19762,N_18715);
or U22602 (N_22602,N_20162,N_20383);
nor U22603 (N_22603,N_18829,N_20159);
and U22604 (N_22604,N_18513,N_18485);
and U22605 (N_22605,N_19810,N_19159);
xor U22606 (N_22606,N_19032,N_18712);
xnor U22607 (N_22607,N_18733,N_19930);
nand U22608 (N_22608,N_18072,N_19560);
nor U22609 (N_22609,N_19577,N_19405);
nor U22610 (N_22610,N_19618,N_18059);
nand U22611 (N_22611,N_18718,N_20772);
or U22612 (N_22612,N_18907,N_19475);
and U22613 (N_22613,N_19151,N_19918);
or U22614 (N_22614,N_18130,N_18953);
xor U22615 (N_22615,N_19509,N_18158);
nor U22616 (N_22616,N_20232,N_19331);
nand U22617 (N_22617,N_20033,N_18123);
or U22618 (N_22618,N_18812,N_19148);
xor U22619 (N_22619,N_18700,N_19063);
xnor U22620 (N_22620,N_19340,N_19995);
nand U22621 (N_22621,N_19339,N_18941);
nor U22622 (N_22622,N_20540,N_19798);
nand U22623 (N_22623,N_20499,N_18541);
and U22624 (N_22624,N_20270,N_20265);
or U22625 (N_22625,N_20400,N_20874);
or U22626 (N_22626,N_20149,N_19011);
xnor U22627 (N_22627,N_19100,N_19032);
or U22628 (N_22628,N_20578,N_20841);
nand U22629 (N_22629,N_19155,N_19471);
xor U22630 (N_22630,N_19988,N_18842);
nor U22631 (N_22631,N_20041,N_20347);
and U22632 (N_22632,N_20848,N_18757);
nor U22633 (N_22633,N_19510,N_19766);
or U22634 (N_22634,N_18599,N_18116);
nand U22635 (N_22635,N_20718,N_19833);
or U22636 (N_22636,N_19048,N_18548);
xor U22637 (N_22637,N_20310,N_19838);
xor U22638 (N_22638,N_19113,N_18765);
xor U22639 (N_22639,N_18463,N_18468);
nand U22640 (N_22640,N_19221,N_18978);
and U22641 (N_22641,N_20636,N_18135);
or U22642 (N_22642,N_19595,N_19564);
or U22643 (N_22643,N_20356,N_20977);
or U22644 (N_22644,N_20365,N_20802);
nor U22645 (N_22645,N_19249,N_18622);
nor U22646 (N_22646,N_19917,N_18866);
nand U22647 (N_22647,N_20659,N_20853);
or U22648 (N_22648,N_19693,N_18761);
or U22649 (N_22649,N_20940,N_20382);
and U22650 (N_22650,N_18349,N_18710);
xor U22651 (N_22651,N_20526,N_18201);
nand U22652 (N_22652,N_19632,N_18833);
xnor U22653 (N_22653,N_18114,N_19342);
nand U22654 (N_22654,N_20955,N_18150);
or U22655 (N_22655,N_18770,N_19567);
and U22656 (N_22656,N_19423,N_20214);
nor U22657 (N_22657,N_19920,N_19564);
and U22658 (N_22658,N_20178,N_19936);
nand U22659 (N_22659,N_19158,N_19885);
or U22660 (N_22660,N_19747,N_20438);
nor U22661 (N_22661,N_19652,N_18594);
or U22662 (N_22662,N_19285,N_18501);
and U22663 (N_22663,N_19601,N_20835);
xor U22664 (N_22664,N_19397,N_20930);
nand U22665 (N_22665,N_18556,N_20986);
and U22666 (N_22666,N_20728,N_20008);
or U22667 (N_22667,N_18606,N_19913);
and U22668 (N_22668,N_20363,N_19218);
or U22669 (N_22669,N_20676,N_18598);
nor U22670 (N_22670,N_20543,N_18080);
and U22671 (N_22671,N_19878,N_19880);
and U22672 (N_22672,N_18178,N_18584);
and U22673 (N_22673,N_18535,N_19212);
nand U22674 (N_22674,N_18428,N_20044);
and U22675 (N_22675,N_18186,N_18950);
nand U22676 (N_22676,N_19704,N_19528);
or U22677 (N_22677,N_18193,N_19303);
nand U22678 (N_22678,N_18732,N_20406);
nor U22679 (N_22679,N_19418,N_18766);
xor U22680 (N_22680,N_20954,N_18922);
xnor U22681 (N_22681,N_20265,N_20908);
xor U22682 (N_22682,N_19406,N_18279);
nand U22683 (N_22683,N_19751,N_20362);
xnor U22684 (N_22684,N_18495,N_19496);
and U22685 (N_22685,N_18549,N_19274);
and U22686 (N_22686,N_19913,N_18521);
or U22687 (N_22687,N_19011,N_20256);
xnor U22688 (N_22688,N_19022,N_18541);
nor U22689 (N_22689,N_18668,N_19099);
and U22690 (N_22690,N_18335,N_18553);
or U22691 (N_22691,N_18804,N_19211);
nand U22692 (N_22692,N_20319,N_19147);
and U22693 (N_22693,N_20197,N_19716);
nand U22694 (N_22694,N_19095,N_20296);
nand U22695 (N_22695,N_18309,N_20709);
xor U22696 (N_22696,N_19483,N_20430);
and U22697 (N_22697,N_19714,N_20539);
xor U22698 (N_22698,N_18678,N_20254);
nor U22699 (N_22699,N_19366,N_19388);
nand U22700 (N_22700,N_20694,N_18093);
or U22701 (N_22701,N_19517,N_18518);
nand U22702 (N_22702,N_18629,N_18536);
and U22703 (N_22703,N_20953,N_20344);
xnor U22704 (N_22704,N_18196,N_18628);
xor U22705 (N_22705,N_18621,N_18562);
or U22706 (N_22706,N_20678,N_20075);
nor U22707 (N_22707,N_19078,N_18053);
xor U22708 (N_22708,N_18113,N_18858);
xnor U22709 (N_22709,N_20037,N_18726);
and U22710 (N_22710,N_20146,N_19079);
nor U22711 (N_22711,N_18602,N_19365);
or U22712 (N_22712,N_18570,N_20167);
xnor U22713 (N_22713,N_19672,N_18284);
xor U22714 (N_22714,N_18393,N_18860);
xnor U22715 (N_22715,N_19589,N_19179);
nor U22716 (N_22716,N_20455,N_18336);
or U22717 (N_22717,N_19172,N_19183);
and U22718 (N_22718,N_19437,N_18607);
xnor U22719 (N_22719,N_20988,N_18419);
nor U22720 (N_22720,N_19573,N_19823);
and U22721 (N_22721,N_20158,N_20065);
or U22722 (N_22722,N_20083,N_19961);
nor U22723 (N_22723,N_20303,N_19948);
nand U22724 (N_22724,N_18842,N_20903);
or U22725 (N_22725,N_18961,N_18223);
and U22726 (N_22726,N_18906,N_18077);
nand U22727 (N_22727,N_20081,N_19405);
nand U22728 (N_22728,N_20010,N_20136);
nor U22729 (N_22729,N_19393,N_20472);
or U22730 (N_22730,N_18346,N_19991);
xnor U22731 (N_22731,N_18273,N_19811);
xnor U22732 (N_22732,N_20426,N_20620);
or U22733 (N_22733,N_18952,N_20891);
and U22734 (N_22734,N_19210,N_18614);
xor U22735 (N_22735,N_18552,N_18272);
nor U22736 (N_22736,N_19016,N_20137);
and U22737 (N_22737,N_18240,N_19044);
and U22738 (N_22738,N_19997,N_18778);
and U22739 (N_22739,N_20581,N_19348);
nor U22740 (N_22740,N_18852,N_20067);
and U22741 (N_22741,N_20022,N_19324);
nor U22742 (N_22742,N_18564,N_18237);
and U22743 (N_22743,N_18141,N_18126);
nor U22744 (N_22744,N_19250,N_20848);
or U22745 (N_22745,N_18819,N_19554);
and U22746 (N_22746,N_18638,N_18296);
nor U22747 (N_22747,N_19730,N_18833);
or U22748 (N_22748,N_18903,N_19915);
and U22749 (N_22749,N_18939,N_18304);
and U22750 (N_22750,N_18188,N_18436);
nand U22751 (N_22751,N_19335,N_18910);
and U22752 (N_22752,N_19149,N_19070);
and U22753 (N_22753,N_19296,N_18395);
nand U22754 (N_22754,N_19457,N_19903);
and U22755 (N_22755,N_19459,N_20376);
nor U22756 (N_22756,N_18664,N_20303);
or U22757 (N_22757,N_19649,N_19895);
or U22758 (N_22758,N_18399,N_19400);
nand U22759 (N_22759,N_20845,N_18905);
or U22760 (N_22760,N_20681,N_18860);
nor U22761 (N_22761,N_20713,N_18563);
xor U22762 (N_22762,N_18234,N_18023);
and U22763 (N_22763,N_18165,N_18535);
or U22764 (N_22764,N_20876,N_18932);
and U22765 (N_22765,N_18361,N_20881);
and U22766 (N_22766,N_18012,N_18117);
and U22767 (N_22767,N_18067,N_19545);
xnor U22768 (N_22768,N_19523,N_20136);
xnor U22769 (N_22769,N_18390,N_18959);
nor U22770 (N_22770,N_18817,N_19534);
nand U22771 (N_22771,N_19460,N_19402);
nand U22772 (N_22772,N_20110,N_20345);
or U22773 (N_22773,N_20911,N_20612);
nor U22774 (N_22774,N_18817,N_18607);
and U22775 (N_22775,N_19130,N_19555);
nand U22776 (N_22776,N_18545,N_20602);
xnor U22777 (N_22777,N_18592,N_19792);
nor U22778 (N_22778,N_20676,N_18810);
nor U22779 (N_22779,N_19686,N_18679);
nand U22780 (N_22780,N_20704,N_18922);
nand U22781 (N_22781,N_18821,N_18863);
xnor U22782 (N_22782,N_19086,N_20210);
or U22783 (N_22783,N_19574,N_19414);
xnor U22784 (N_22784,N_20412,N_20827);
nor U22785 (N_22785,N_19817,N_18661);
xnor U22786 (N_22786,N_18032,N_20557);
or U22787 (N_22787,N_20617,N_20873);
nand U22788 (N_22788,N_18884,N_19128);
nand U22789 (N_22789,N_20260,N_19623);
or U22790 (N_22790,N_20189,N_19293);
nor U22791 (N_22791,N_19124,N_18219);
nand U22792 (N_22792,N_20589,N_18409);
or U22793 (N_22793,N_18010,N_19530);
and U22794 (N_22794,N_19896,N_18913);
xor U22795 (N_22795,N_20404,N_18359);
or U22796 (N_22796,N_20874,N_20562);
nand U22797 (N_22797,N_18734,N_19665);
nor U22798 (N_22798,N_18414,N_20666);
xnor U22799 (N_22799,N_18291,N_20295);
xnor U22800 (N_22800,N_19679,N_20437);
xor U22801 (N_22801,N_19267,N_18230);
or U22802 (N_22802,N_20199,N_20846);
nand U22803 (N_22803,N_18263,N_19100);
xnor U22804 (N_22804,N_20194,N_20481);
xor U22805 (N_22805,N_18189,N_20140);
nand U22806 (N_22806,N_20320,N_19997);
xor U22807 (N_22807,N_18727,N_18187);
xor U22808 (N_22808,N_18466,N_19461);
nand U22809 (N_22809,N_20295,N_18093);
and U22810 (N_22810,N_19181,N_20165);
nor U22811 (N_22811,N_18109,N_18953);
nor U22812 (N_22812,N_18588,N_18701);
nand U22813 (N_22813,N_20664,N_20363);
xnor U22814 (N_22814,N_20577,N_18798);
xnor U22815 (N_22815,N_19740,N_18881);
and U22816 (N_22816,N_19879,N_20736);
nand U22817 (N_22817,N_19179,N_19105);
xnor U22818 (N_22818,N_19938,N_18141);
nor U22819 (N_22819,N_19360,N_19419);
or U22820 (N_22820,N_18806,N_19237);
xor U22821 (N_22821,N_18360,N_18620);
nor U22822 (N_22822,N_19151,N_20527);
and U22823 (N_22823,N_19770,N_19293);
and U22824 (N_22824,N_20399,N_20727);
or U22825 (N_22825,N_19197,N_20974);
xor U22826 (N_22826,N_19893,N_19541);
nor U22827 (N_22827,N_19112,N_18355);
xnor U22828 (N_22828,N_18732,N_19478);
or U22829 (N_22829,N_19977,N_20178);
or U22830 (N_22830,N_19118,N_18842);
and U22831 (N_22831,N_18270,N_20634);
and U22832 (N_22832,N_18748,N_18475);
xor U22833 (N_22833,N_18245,N_19763);
nor U22834 (N_22834,N_19769,N_19989);
or U22835 (N_22835,N_20578,N_19669);
nor U22836 (N_22836,N_19952,N_18352);
and U22837 (N_22837,N_20235,N_18894);
or U22838 (N_22838,N_18801,N_19731);
nand U22839 (N_22839,N_19917,N_20642);
xor U22840 (N_22840,N_19067,N_20531);
xnor U22841 (N_22841,N_20092,N_18047);
and U22842 (N_22842,N_20537,N_20451);
nor U22843 (N_22843,N_20351,N_19014);
or U22844 (N_22844,N_18750,N_20244);
and U22845 (N_22845,N_19686,N_18071);
nor U22846 (N_22846,N_20442,N_19037);
nand U22847 (N_22847,N_19657,N_20788);
nand U22848 (N_22848,N_19567,N_20580);
xnor U22849 (N_22849,N_20148,N_19431);
or U22850 (N_22850,N_20639,N_20902);
xor U22851 (N_22851,N_18151,N_19605);
or U22852 (N_22852,N_20527,N_18761);
and U22853 (N_22853,N_20847,N_19341);
xor U22854 (N_22854,N_20386,N_18081);
nand U22855 (N_22855,N_18332,N_18245);
and U22856 (N_22856,N_19537,N_20418);
and U22857 (N_22857,N_20914,N_20758);
nor U22858 (N_22858,N_18329,N_18665);
and U22859 (N_22859,N_18092,N_18672);
xnor U22860 (N_22860,N_18261,N_20425);
and U22861 (N_22861,N_19379,N_18596);
nor U22862 (N_22862,N_18389,N_18409);
xnor U22863 (N_22863,N_19528,N_20192);
nand U22864 (N_22864,N_19746,N_19716);
or U22865 (N_22865,N_20446,N_18576);
and U22866 (N_22866,N_19607,N_20114);
nand U22867 (N_22867,N_18236,N_19424);
nand U22868 (N_22868,N_19691,N_18496);
nand U22869 (N_22869,N_20862,N_20680);
nand U22870 (N_22870,N_18988,N_18367);
nand U22871 (N_22871,N_19542,N_19044);
nand U22872 (N_22872,N_18403,N_20063);
xnor U22873 (N_22873,N_18537,N_19294);
and U22874 (N_22874,N_20090,N_20131);
nand U22875 (N_22875,N_18308,N_20424);
nand U22876 (N_22876,N_20076,N_19762);
nand U22877 (N_22877,N_18904,N_19694);
nor U22878 (N_22878,N_19902,N_18977);
nand U22879 (N_22879,N_19066,N_18543);
or U22880 (N_22880,N_20526,N_19155);
or U22881 (N_22881,N_20786,N_20237);
nor U22882 (N_22882,N_20573,N_18891);
and U22883 (N_22883,N_19765,N_20190);
xor U22884 (N_22884,N_20529,N_20464);
or U22885 (N_22885,N_18714,N_19752);
xnor U22886 (N_22886,N_19953,N_18894);
nor U22887 (N_22887,N_19662,N_18044);
xnor U22888 (N_22888,N_18477,N_19112);
nor U22889 (N_22889,N_18598,N_18234);
xor U22890 (N_22890,N_18770,N_19668);
nand U22891 (N_22891,N_19480,N_20467);
nor U22892 (N_22892,N_20522,N_20025);
nor U22893 (N_22893,N_20449,N_19905);
or U22894 (N_22894,N_19571,N_18940);
xnor U22895 (N_22895,N_18958,N_19825);
xnor U22896 (N_22896,N_20934,N_19972);
nor U22897 (N_22897,N_18432,N_20118);
and U22898 (N_22898,N_19485,N_18181);
nand U22899 (N_22899,N_20364,N_20543);
nor U22900 (N_22900,N_19678,N_18216);
and U22901 (N_22901,N_20778,N_18488);
or U22902 (N_22902,N_20491,N_18107);
nor U22903 (N_22903,N_20083,N_19644);
nor U22904 (N_22904,N_18406,N_19310);
and U22905 (N_22905,N_18380,N_19026);
nand U22906 (N_22906,N_20060,N_20654);
xnor U22907 (N_22907,N_18569,N_18760);
xor U22908 (N_22908,N_19969,N_19433);
nand U22909 (N_22909,N_19736,N_20109);
and U22910 (N_22910,N_19915,N_18825);
nand U22911 (N_22911,N_19907,N_18622);
xor U22912 (N_22912,N_18746,N_19641);
nor U22913 (N_22913,N_18252,N_19995);
and U22914 (N_22914,N_18961,N_18636);
and U22915 (N_22915,N_18711,N_18534);
nor U22916 (N_22916,N_20840,N_19562);
xnor U22917 (N_22917,N_19106,N_18658);
nor U22918 (N_22918,N_18629,N_18639);
nand U22919 (N_22919,N_19169,N_19586);
xnor U22920 (N_22920,N_18465,N_18026);
nor U22921 (N_22921,N_18149,N_20739);
or U22922 (N_22922,N_19832,N_20799);
or U22923 (N_22923,N_19791,N_19223);
nand U22924 (N_22924,N_20925,N_18188);
xor U22925 (N_22925,N_19056,N_19565);
xnor U22926 (N_22926,N_18036,N_20240);
nand U22927 (N_22927,N_19129,N_18984);
nor U22928 (N_22928,N_18333,N_18247);
xor U22929 (N_22929,N_20096,N_19066);
nand U22930 (N_22930,N_18416,N_20983);
xor U22931 (N_22931,N_18155,N_19691);
and U22932 (N_22932,N_20172,N_19839);
and U22933 (N_22933,N_18323,N_19574);
nand U22934 (N_22934,N_20882,N_20248);
xor U22935 (N_22935,N_20108,N_19916);
xor U22936 (N_22936,N_20938,N_18341);
nor U22937 (N_22937,N_20342,N_18237);
nand U22938 (N_22938,N_20849,N_20766);
nor U22939 (N_22939,N_19835,N_18472);
and U22940 (N_22940,N_19644,N_20071);
or U22941 (N_22941,N_20766,N_20866);
or U22942 (N_22942,N_18071,N_19309);
or U22943 (N_22943,N_20158,N_20929);
or U22944 (N_22944,N_19397,N_18927);
and U22945 (N_22945,N_19564,N_20467);
nor U22946 (N_22946,N_18194,N_20267);
and U22947 (N_22947,N_18393,N_18651);
or U22948 (N_22948,N_20451,N_19851);
xor U22949 (N_22949,N_20454,N_18196);
or U22950 (N_22950,N_20541,N_20043);
nor U22951 (N_22951,N_19489,N_18155);
nand U22952 (N_22952,N_19111,N_19348);
or U22953 (N_22953,N_20212,N_20926);
or U22954 (N_22954,N_18058,N_18576);
nor U22955 (N_22955,N_18763,N_19462);
and U22956 (N_22956,N_20944,N_20900);
nand U22957 (N_22957,N_19062,N_19794);
or U22958 (N_22958,N_19177,N_19002);
nand U22959 (N_22959,N_19451,N_20060);
or U22960 (N_22960,N_19332,N_19521);
xnor U22961 (N_22961,N_19774,N_18193);
nor U22962 (N_22962,N_19997,N_18925);
nand U22963 (N_22963,N_20122,N_19114);
nand U22964 (N_22964,N_19218,N_18389);
or U22965 (N_22965,N_20496,N_19296);
nand U22966 (N_22966,N_18520,N_20126);
and U22967 (N_22967,N_18230,N_19634);
nand U22968 (N_22968,N_18188,N_20896);
or U22969 (N_22969,N_19262,N_19243);
or U22970 (N_22970,N_18647,N_19791);
nand U22971 (N_22971,N_20581,N_18950);
or U22972 (N_22972,N_19417,N_20302);
xnor U22973 (N_22973,N_18705,N_18453);
xnor U22974 (N_22974,N_20672,N_20487);
nor U22975 (N_22975,N_18295,N_19230);
nor U22976 (N_22976,N_19745,N_18391);
xnor U22977 (N_22977,N_20208,N_18549);
xor U22978 (N_22978,N_18310,N_20116);
xnor U22979 (N_22979,N_20885,N_20642);
nand U22980 (N_22980,N_18081,N_19903);
nor U22981 (N_22981,N_20426,N_20918);
nor U22982 (N_22982,N_20351,N_19270);
xnor U22983 (N_22983,N_18412,N_20606);
nand U22984 (N_22984,N_20098,N_18903);
xor U22985 (N_22985,N_18496,N_20949);
nor U22986 (N_22986,N_18895,N_20164);
and U22987 (N_22987,N_20868,N_20710);
nand U22988 (N_22988,N_19628,N_19820);
and U22989 (N_22989,N_18615,N_19614);
and U22990 (N_22990,N_19781,N_20434);
and U22991 (N_22991,N_20541,N_19783);
and U22992 (N_22992,N_20725,N_20696);
nor U22993 (N_22993,N_18639,N_20650);
xnor U22994 (N_22994,N_19367,N_20652);
nand U22995 (N_22995,N_20676,N_19722);
or U22996 (N_22996,N_19969,N_20488);
nand U22997 (N_22997,N_19638,N_18294);
or U22998 (N_22998,N_19188,N_20240);
nor U22999 (N_22999,N_20644,N_18674);
nand U23000 (N_23000,N_20450,N_18317);
or U23001 (N_23001,N_19153,N_20262);
nand U23002 (N_23002,N_18702,N_18010);
nand U23003 (N_23003,N_20648,N_19461);
and U23004 (N_23004,N_18033,N_19021);
xor U23005 (N_23005,N_20768,N_18947);
or U23006 (N_23006,N_18636,N_20256);
nor U23007 (N_23007,N_18666,N_19640);
xor U23008 (N_23008,N_19834,N_18081);
and U23009 (N_23009,N_19336,N_20924);
or U23010 (N_23010,N_19413,N_19199);
nand U23011 (N_23011,N_19414,N_19222);
or U23012 (N_23012,N_18415,N_19856);
xnor U23013 (N_23013,N_19592,N_18446);
xnor U23014 (N_23014,N_20608,N_18237);
and U23015 (N_23015,N_19821,N_18114);
or U23016 (N_23016,N_19499,N_18415);
xnor U23017 (N_23017,N_20426,N_20272);
and U23018 (N_23018,N_18713,N_20079);
and U23019 (N_23019,N_20909,N_20150);
and U23020 (N_23020,N_19231,N_19462);
nor U23021 (N_23021,N_20347,N_19213);
and U23022 (N_23022,N_18353,N_19529);
nand U23023 (N_23023,N_18090,N_20092);
and U23024 (N_23024,N_19886,N_18267);
xor U23025 (N_23025,N_20908,N_19125);
nor U23026 (N_23026,N_19074,N_19488);
nor U23027 (N_23027,N_18732,N_19534);
or U23028 (N_23028,N_20919,N_18229);
or U23029 (N_23029,N_19328,N_19248);
or U23030 (N_23030,N_19830,N_18722);
nor U23031 (N_23031,N_18512,N_19648);
nor U23032 (N_23032,N_18608,N_18594);
and U23033 (N_23033,N_20695,N_20579);
or U23034 (N_23034,N_18999,N_20963);
nand U23035 (N_23035,N_20967,N_18138);
and U23036 (N_23036,N_19369,N_18763);
nor U23037 (N_23037,N_19329,N_20675);
nand U23038 (N_23038,N_18261,N_19194);
xnor U23039 (N_23039,N_18483,N_18346);
xor U23040 (N_23040,N_18047,N_20589);
and U23041 (N_23041,N_19196,N_19737);
or U23042 (N_23042,N_19891,N_20487);
and U23043 (N_23043,N_19725,N_18294);
or U23044 (N_23044,N_20260,N_19955);
nand U23045 (N_23045,N_20384,N_20164);
nor U23046 (N_23046,N_20526,N_20471);
nor U23047 (N_23047,N_18742,N_18245);
nand U23048 (N_23048,N_19499,N_19611);
nand U23049 (N_23049,N_20120,N_18279);
and U23050 (N_23050,N_18200,N_19654);
or U23051 (N_23051,N_20888,N_20044);
xor U23052 (N_23052,N_20275,N_18105);
or U23053 (N_23053,N_19146,N_20875);
or U23054 (N_23054,N_19590,N_19035);
nor U23055 (N_23055,N_19547,N_20882);
nand U23056 (N_23056,N_20904,N_20738);
xor U23057 (N_23057,N_18550,N_20295);
nor U23058 (N_23058,N_20596,N_19744);
or U23059 (N_23059,N_19135,N_19272);
or U23060 (N_23060,N_20501,N_20914);
nor U23061 (N_23061,N_18996,N_18824);
nand U23062 (N_23062,N_19129,N_20687);
xor U23063 (N_23063,N_18476,N_18725);
and U23064 (N_23064,N_18253,N_19130);
nor U23065 (N_23065,N_18256,N_20166);
xnor U23066 (N_23066,N_20712,N_19436);
nor U23067 (N_23067,N_19365,N_18463);
nand U23068 (N_23068,N_18734,N_19170);
and U23069 (N_23069,N_19948,N_18618);
nand U23070 (N_23070,N_19884,N_19855);
nor U23071 (N_23071,N_19821,N_20073);
nor U23072 (N_23072,N_20980,N_18218);
and U23073 (N_23073,N_20612,N_20589);
nor U23074 (N_23074,N_19486,N_18720);
nor U23075 (N_23075,N_18110,N_19590);
nand U23076 (N_23076,N_18041,N_18151);
and U23077 (N_23077,N_19692,N_18655);
and U23078 (N_23078,N_20258,N_19891);
nand U23079 (N_23079,N_20023,N_19458);
or U23080 (N_23080,N_19818,N_19298);
nor U23081 (N_23081,N_19010,N_18108);
nand U23082 (N_23082,N_19425,N_18135);
nand U23083 (N_23083,N_18423,N_20461);
or U23084 (N_23084,N_18877,N_19431);
xor U23085 (N_23085,N_19612,N_20709);
nand U23086 (N_23086,N_19372,N_20665);
and U23087 (N_23087,N_18458,N_20429);
or U23088 (N_23088,N_18794,N_20169);
or U23089 (N_23089,N_20732,N_20823);
nand U23090 (N_23090,N_18881,N_18326);
and U23091 (N_23091,N_18421,N_20265);
nand U23092 (N_23092,N_18280,N_19631);
and U23093 (N_23093,N_20711,N_20307);
nand U23094 (N_23094,N_20720,N_18235);
or U23095 (N_23095,N_18274,N_18854);
xnor U23096 (N_23096,N_18941,N_20722);
nand U23097 (N_23097,N_19858,N_19598);
nand U23098 (N_23098,N_18626,N_19553);
and U23099 (N_23099,N_19787,N_18610);
nor U23100 (N_23100,N_18228,N_18933);
nand U23101 (N_23101,N_19940,N_20691);
or U23102 (N_23102,N_19912,N_19258);
xnor U23103 (N_23103,N_20227,N_19538);
xnor U23104 (N_23104,N_20222,N_20630);
nand U23105 (N_23105,N_18319,N_19914);
and U23106 (N_23106,N_18707,N_18420);
nand U23107 (N_23107,N_20987,N_20233);
or U23108 (N_23108,N_19439,N_18181);
or U23109 (N_23109,N_19937,N_20030);
nor U23110 (N_23110,N_20701,N_18912);
or U23111 (N_23111,N_18119,N_19729);
or U23112 (N_23112,N_19849,N_20151);
or U23113 (N_23113,N_19230,N_18263);
and U23114 (N_23114,N_20909,N_19894);
and U23115 (N_23115,N_19016,N_20952);
nor U23116 (N_23116,N_20233,N_19256);
and U23117 (N_23117,N_18959,N_18783);
xnor U23118 (N_23118,N_18576,N_20255);
or U23119 (N_23119,N_20575,N_20401);
or U23120 (N_23120,N_19422,N_20796);
xnor U23121 (N_23121,N_19389,N_18677);
and U23122 (N_23122,N_18499,N_18161);
nand U23123 (N_23123,N_18137,N_20055);
and U23124 (N_23124,N_18886,N_19110);
or U23125 (N_23125,N_19207,N_20145);
xor U23126 (N_23126,N_20500,N_19414);
or U23127 (N_23127,N_18732,N_18356);
and U23128 (N_23128,N_20237,N_20611);
nand U23129 (N_23129,N_19164,N_18568);
or U23130 (N_23130,N_19491,N_18981);
xor U23131 (N_23131,N_20149,N_19706);
nand U23132 (N_23132,N_18164,N_18829);
nand U23133 (N_23133,N_18258,N_19776);
or U23134 (N_23134,N_19584,N_20494);
or U23135 (N_23135,N_20666,N_18751);
or U23136 (N_23136,N_18848,N_19416);
xnor U23137 (N_23137,N_18650,N_18145);
nand U23138 (N_23138,N_19927,N_19297);
nand U23139 (N_23139,N_19236,N_20033);
or U23140 (N_23140,N_18222,N_18004);
nand U23141 (N_23141,N_19431,N_18743);
xor U23142 (N_23142,N_18868,N_19406);
and U23143 (N_23143,N_19003,N_20953);
xor U23144 (N_23144,N_20390,N_20976);
or U23145 (N_23145,N_19600,N_20662);
nor U23146 (N_23146,N_19274,N_20331);
nor U23147 (N_23147,N_19725,N_20313);
xor U23148 (N_23148,N_18277,N_20069);
and U23149 (N_23149,N_19495,N_18325);
and U23150 (N_23150,N_19656,N_20977);
nand U23151 (N_23151,N_19745,N_20220);
or U23152 (N_23152,N_19246,N_20617);
nand U23153 (N_23153,N_18941,N_20134);
nand U23154 (N_23154,N_18232,N_19415);
nor U23155 (N_23155,N_18150,N_18002);
xnor U23156 (N_23156,N_19246,N_20454);
xnor U23157 (N_23157,N_20896,N_20730);
xor U23158 (N_23158,N_20018,N_18377);
nor U23159 (N_23159,N_19648,N_18474);
and U23160 (N_23160,N_19823,N_19983);
nor U23161 (N_23161,N_18996,N_18886);
or U23162 (N_23162,N_18916,N_20883);
or U23163 (N_23163,N_20283,N_19234);
and U23164 (N_23164,N_20356,N_18828);
nand U23165 (N_23165,N_19397,N_18402);
nand U23166 (N_23166,N_18615,N_19860);
xnor U23167 (N_23167,N_18560,N_20694);
nand U23168 (N_23168,N_18265,N_19293);
xor U23169 (N_23169,N_20394,N_18806);
or U23170 (N_23170,N_20102,N_20860);
or U23171 (N_23171,N_19702,N_18878);
or U23172 (N_23172,N_20648,N_20876);
or U23173 (N_23173,N_20035,N_18958);
and U23174 (N_23174,N_18529,N_20518);
or U23175 (N_23175,N_20489,N_19548);
xnor U23176 (N_23176,N_19802,N_20327);
nand U23177 (N_23177,N_20889,N_19505);
nand U23178 (N_23178,N_18657,N_20021);
or U23179 (N_23179,N_19004,N_20248);
nor U23180 (N_23180,N_20730,N_19747);
or U23181 (N_23181,N_18264,N_18583);
nand U23182 (N_23182,N_18875,N_19770);
or U23183 (N_23183,N_20958,N_20639);
nand U23184 (N_23184,N_18452,N_20303);
and U23185 (N_23185,N_18639,N_19008);
nor U23186 (N_23186,N_20278,N_19889);
nor U23187 (N_23187,N_19773,N_19152);
nand U23188 (N_23188,N_19503,N_20516);
or U23189 (N_23189,N_18861,N_18453);
or U23190 (N_23190,N_18526,N_19179);
nor U23191 (N_23191,N_19369,N_19884);
nand U23192 (N_23192,N_20088,N_18146);
xnor U23193 (N_23193,N_18461,N_18126);
nand U23194 (N_23194,N_20288,N_20603);
and U23195 (N_23195,N_19552,N_18220);
xor U23196 (N_23196,N_18415,N_18571);
xnor U23197 (N_23197,N_20888,N_18098);
nor U23198 (N_23198,N_18461,N_20655);
and U23199 (N_23199,N_20264,N_19402);
or U23200 (N_23200,N_19583,N_18981);
nor U23201 (N_23201,N_19940,N_18404);
xor U23202 (N_23202,N_18889,N_18933);
and U23203 (N_23203,N_20621,N_18862);
nor U23204 (N_23204,N_20436,N_19817);
or U23205 (N_23205,N_19215,N_19349);
or U23206 (N_23206,N_18859,N_19569);
nor U23207 (N_23207,N_20420,N_19711);
or U23208 (N_23208,N_19269,N_18097);
or U23209 (N_23209,N_18702,N_18785);
or U23210 (N_23210,N_19392,N_18444);
nor U23211 (N_23211,N_20571,N_19222);
xor U23212 (N_23212,N_20294,N_20767);
xor U23213 (N_23213,N_19632,N_18560);
and U23214 (N_23214,N_19395,N_20109);
nand U23215 (N_23215,N_18542,N_20716);
nand U23216 (N_23216,N_18223,N_19399);
nand U23217 (N_23217,N_18874,N_19558);
nand U23218 (N_23218,N_18983,N_19063);
or U23219 (N_23219,N_18664,N_18072);
and U23220 (N_23220,N_18362,N_18036);
xor U23221 (N_23221,N_18901,N_20748);
or U23222 (N_23222,N_18951,N_19631);
nor U23223 (N_23223,N_20476,N_18875);
or U23224 (N_23224,N_18531,N_18437);
or U23225 (N_23225,N_18051,N_18713);
or U23226 (N_23226,N_19753,N_20114);
and U23227 (N_23227,N_20180,N_18238);
or U23228 (N_23228,N_19579,N_19983);
nor U23229 (N_23229,N_18261,N_20199);
or U23230 (N_23230,N_18639,N_18331);
xor U23231 (N_23231,N_18847,N_20165);
and U23232 (N_23232,N_18715,N_19331);
xor U23233 (N_23233,N_19964,N_18957);
xor U23234 (N_23234,N_20769,N_19032);
and U23235 (N_23235,N_20129,N_20224);
and U23236 (N_23236,N_19930,N_18377);
and U23237 (N_23237,N_18083,N_19392);
and U23238 (N_23238,N_20288,N_18331);
nor U23239 (N_23239,N_19696,N_20486);
and U23240 (N_23240,N_20259,N_19836);
nand U23241 (N_23241,N_20179,N_20518);
or U23242 (N_23242,N_19564,N_19178);
nand U23243 (N_23243,N_20101,N_19192);
nand U23244 (N_23244,N_20029,N_18715);
or U23245 (N_23245,N_19036,N_19624);
nor U23246 (N_23246,N_20187,N_20208);
nor U23247 (N_23247,N_18685,N_18715);
nor U23248 (N_23248,N_18178,N_18891);
and U23249 (N_23249,N_20691,N_20080);
and U23250 (N_23250,N_18737,N_20366);
and U23251 (N_23251,N_18023,N_20446);
and U23252 (N_23252,N_18916,N_19324);
and U23253 (N_23253,N_19533,N_20904);
or U23254 (N_23254,N_18239,N_20835);
nor U23255 (N_23255,N_20443,N_20435);
or U23256 (N_23256,N_18401,N_19262);
nor U23257 (N_23257,N_18970,N_18199);
or U23258 (N_23258,N_18367,N_19353);
or U23259 (N_23259,N_19300,N_18735);
or U23260 (N_23260,N_20383,N_18160);
or U23261 (N_23261,N_18908,N_19259);
nand U23262 (N_23262,N_18817,N_18425);
xor U23263 (N_23263,N_19237,N_20062);
or U23264 (N_23264,N_20057,N_18082);
xor U23265 (N_23265,N_18521,N_20159);
nor U23266 (N_23266,N_19491,N_20242);
nand U23267 (N_23267,N_18926,N_19434);
and U23268 (N_23268,N_18429,N_18826);
xnor U23269 (N_23269,N_18496,N_19036);
or U23270 (N_23270,N_20761,N_20366);
nor U23271 (N_23271,N_20526,N_19128);
nor U23272 (N_23272,N_19654,N_20267);
xor U23273 (N_23273,N_18659,N_20978);
xor U23274 (N_23274,N_20746,N_18875);
and U23275 (N_23275,N_20649,N_19608);
nand U23276 (N_23276,N_19465,N_20612);
or U23277 (N_23277,N_19815,N_18625);
and U23278 (N_23278,N_19207,N_18898);
or U23279 (N_23279,N_18357,N_20772);
or U23280 (N_23280,N_20620,N_18163);
xnor U23281 (N_23281,N_19327,N_19012);
or U23282 (N_23282,N_18607,N_19979);
nor U23283 (N_23283,N_18174,N_20255);
or U23284 (N_23284,N_20746,N_19149);
and U23285 (N_23285,N_19209,N_19382);
or U23286 (N_23286,N_19801,N_20388);
nor U23287 (N_23287,N_20796,N_20108);
xor U23288 (N_23288,N_18707,N_19268);
and U23289 (N_23289,N_20014,N_18827);
nor U23290 (N_23290,N_19214,N_20610);
nor U23291 (N_23291,N_19844,N_18512);
xnor U23292 (N_23292,N_19251,N_20078);
nor U23293 (N_23293,N_19736,N_20061);
and U23294 (N_23294,N_19191,N_19512);
nand U23295 (N_23295,N_18573,N_18699);
xnor U23296 (N_23296,N_20872,N_20488);
xor U23297 (N_23297,N_20678,N_19228);
xor U23298 (N_23298,N_19348,N_18218);
nand U23299 (N_23299,N_18645,N_18210);
or U23300 (N_23300,N_20428,N_20106);
nand U23301 (N_23301,N_18186,N_19028);
or U23302 (N_23302,N_19818,N_18520);
or U23303 (N_23303,N_18444,N_19956);
or U23304 (N_23304,N_20709,N_20677);
xor U23305 (N_23305,N_18346,N_19868);
or U23306 (N_23306,N_18106,N_19027);
xor U23307 (N_23307,N_18273,N_20910);
nand U23308 (N_23308,N_20323,N_20270);
nor U23309 (N_23309,N_20517,N_19628);
xor U23310 (N_23310,N_18503,N_18810);
nand U23311 (N_23311,N_19232,N_20352);
nand U23312 (N_23312,N_19949,N_18880);
or U23313 (N_23313,N_18907,N_20415);
xnor U23314 (N_23314,N_19173,N_18895);
xnor U23315 (N_23315,N_19194,N_18783);
nand U23316 (N_23316,N_18656,N_20806);
and U23317 (N_23317,N_20909,N_18748);
or U23318 (N_23318,N_18007,N_20348);
or U23319 (N_23319,N_18582,N_19825);
nand U23320 (N_23320,N_19628,N_18604);
xor U23321 (N_23321,N_18947,N_18670);
nand U23322 (N_23322,N_20963,N_19231);
xor U23323 (N_23323,N_19058,N_20488);
xnor U23324 (N_23324,N_18195,N_19456);
and U23325 (N_23325,N_19484,N_20266);
and U23326 (N_23326,N_19470,N_19545);
nor U23327 (N_23327,N_19750,N_20955);
xnor U23328 (N_23328,N_20795,N_20132);
nand U23329 (N_23329,N_20672,N_19420);
xor U23330 (N_23330,N_19664,N_18327);
nor U23331 (N_23331,N_19696,N_20518);
nand U23332 (N_23332,N_20043,N_19129);
nor U23333 (N_23333,N_20523,N_19738);
xnor U23334 (N_23334,N_18177,N_20420);
and U23335 (N_23335,N_19222,N_19142);
or U23336 (N_23336,N_20502,N_19018);
nand U23337 (N_23337,N_20126,N_19334);
nor U23338 (N_23338,N_20220,N_19497);
and U23339 (N_23339,N_18816,N_20249);
or U23340 (N_23340,N_19998,N_19073);
nand U23341 (N_23341,N_20518,N_20608);
or U23342 (N_23342,N_20789,N_19573);
and U23343 (N_23343,N_18244,N_20714);
or U23344 (N_23344,N_19729,N_20089);
or U23345 (N_23345,N_19249,N_20805);
xor U23346 (N_23346,N_19283,N_20614);
xnor U23347 (N_23347,N_20441,N_19369);
or U23348 (N_23348,N_19600,N_19003);
xor U23349 (N_23349,N_18915,N_20957);
and U23350 (N_23350,N_18997,N_19280);
xnor U23351 (N_23351,N_20328,N_18041);
nor U23352 (N_23352,N_18178,N_20172);
or U23353 (N_23353,N_20260,N_19115);
nor U23354 (N_23354,N_20340,N_20087);
nor U23355 (N_23355,N_20486,N_18951);
nand U23356 (N_23356,N_18500,N_19146);
and U23357 (N_23357,N_18432,N_20838);
nand U23358 (N_23358,N_20872,N_18702);
and U23359 (N_23359,N_20417,N_19879);
and U23360 (N_23360,N_20195,N_20312);
xnor U23361 (N_23361,N_20210,N_20437);
and U23362 (N_23362,N_20283,N_19091);
nor U23363 (N_23363,N_20877,N_18180);
xor U23364 (N_23364,N_20470,N_19914);
nand U23365 (N_23365,N_18255,N_20461);
and U23366 (N_23366,N_18554,N_18754);
or U23367 (N_23367,N_18102,N_20354);
nor U23368 (N_23368,N_18597,N_19626);
xor U23369 (N_23369,N_20151,N_19206);
or U23370 (N_23370,N_19106,N_18429);
nand U23371 (N_23371,N_18721,N_19676);
xor U23372 (N_23372,N_19193,N_19400);
nand U23373 (N_23373,N_18174,N_19179);
nor U23374 (N_23374,N_20232,N_18661);
or U23375 (N_23375,N_19251,N_18481);
xnor U23376 (N_23376,N_20707,N_19888);
or U23377 (N_23377,N_20330,N_20704);
nor U23378 (N_23378,N_18399,N_19058);
and U23379 (N_23379,N_18589,N_18640);
or U23380 (N_23380,N_20066,N_18913);
nor U23381 (N_23381,N_19328,N_20574);
xor U23382 (N_23382,N_20025,N_20970);
xnor U23383 (N_23383,N_19124,N_20741);
or U23384 (N_23384,N_19211,N_18136);
xnor U23385 (N_23385,N_20199,N_19199);
nand U23386 (N_23386,N_19974,N_20942);
and U23387 (N_23387,N_18548,N_19029);
and U23388 (N_23388,N_20891,N_19903);
nor U23389 (N_23389,N_19176,N_19560);
nor U23390 (N_23390,N_20230,N_18575);
nand U23391 (N_23391,N_18986,N_20228);
nand U23392 (N_23392,N_18313,N_18012);
nor U23393 (N_23393,N_18800,N_19641);
xor U23394 (N_23394,N_18540,N_18608);
or U23395 (N_23395,N_18926,N_19043);
or U23396 (N_23396,N_18774,N_18885);
xnor U23397 (N_23397,N_18506,N_19294);
nand U23398 (N_23398,N_18127,N_18285);
nor U23399 (N_23399,N_18315,N_18380);
xnor U23400 (N_23400,N_19955,N_18320);
xor U23401 (N_23401,N_20504,N_20585);
nor U23402 (N_23402,N_19957,N_20079);
nand U23403 (N_23403,N_18287,N_20344);
nand U23404 (N_23404,N_19412,N_18298);
or U23405 (N_23405,N_18989,N_20031);
nor U23406 (N_23406,N_19383,N_20741);
and U23407 (N_23407,N_18567,N_20465);
and U23408 (N_23408,N_18734,N_18371);
or U23409 (N_23409,N_20242,N_19697);
nor U23410 (N_23410,N_18744,N_20542);
and U23411 (N_23411,N_18879,N_20471);
nor U23412 (N_23412,N_19653,N_18900);
nand U23413 (N_23413,N_19151,N_20236);
nand U23414 (N_23414,N_20559,N_18900);
nand U23415 (N_23415,N_19444,N_18028);
nand U23416 (N_23416,N_19864,N_20730);
xnor U23417 (N_23417,N_19790,N_20326);
or U23418 (N_23418,N_18995,N_19644);
nor U23419 (N_23419,N_20418,N_19648);
and U23420 (N_23420,N_19801,N_19301);
and U23421 (N_23421,N_18829,N_20959);
and U23422 (N_23422,N_18638,N_20451);
and U23423 (N_23423,N_20198,N_19462);
nor U23424 (N_23424,N_20285,N_18792);
and U23425 (N_23425,N_19011,N_18433);
or U23426 (N_23426,N_19450,N_19178);
nand U23427 (N_23427,N_20837,N_18431);
nand U23428 (N_23428,N_18975,N_20127);
nor U23429 (N_23429,N_19029,N_20054);
xnor U23430 (N_23430,N_18956,N_18919);
or U23431 (N_23431,N_20225,N_19407);
or U23432 (N_23432,N_20876,N_18239);
xnor U23433 (N_23433,N_18745,N_20624);
nand U23434 (N_23434,N_18042,N_18306);
nand U23435 (N_23435,N_18449,N_19145);
nand U23436 (N_23436,N_20428,N_18290);
xnor U23437 (N_23437,N_19763,N_18686);
nor U23438 (N_23438,N_19075,N_20591);
nor U23439 (N_23439,N_18999,N_19698);
xor U23440 (N_23440,N_20099,N_20283);
nor U23441 (N_23441,N_20332,N_18801);
nand U23442 (N_23442,N_19922,N_20961);
nor U23443 (N_23443,N_18248,N_19678);
nand U23444 (N_23444,N_20885,N_20409);
and U23445 (N_23445,N_18187,N_20183);
xor U23446 (N_23446,N_18047,N_19358);
and U23447 (N_23447,N_19226,N_20379);
xor U23448 (N_23448,N_20056,N_20832);
xor U23449 (N_23449,N_19411,N_19761);
nand U23450 (N_23450,N_18799,N_18994);
xnor U23451 (N_23451,N_19194,N_18028);
and U23452 (N_23452,N_18207,N_20756);
nand U23453 (N_23453,N_18612,N_20736);
or U23454 (N_23454,N_18887,N_20572);
or U23455 (N_23455,N_19904,N_19303);
nand U23456 (N_23456,N_18806,N_20523);
nand U23457 (N_23457,N_18465,N_18745);
nand U23458 (N_23458,N_19661,N_20434);
xnor U23459 (N_23459,N_18109,N_18441);
nor U23460 (N_23460,N_19559,N_18487);
and U23461 (N_23461,N_18977,N_18327);
or U23462 (N_23462,N_20637,N_19723);
nand U23463 (N_23463,N_20485,N_18107);
nor U23464 (N_23464,N_20864,N_18949);
nand U23465 (N_23465,N_18857,N_20156);
nor U23466 (N_23466,N_19062,N_19944);
nand U23467 (N_23467,N_18615,N_18168);
and U23468 (N_23468,N_20685,N_19552);
or U23469 (N_23469,N_20691,N_19012);
or U23470 (N_23470,N_20897,N_20056);
nor U23471 (N_23471,N_19169,N_18284);
xor U23472 (N_23472,N_18474,N_19682);
or U23473 (N_23473,N_20227,N_19305);
and U23474 (N_23474,N_18221,N_18318);
nand U23475 (N_23475,N_19302,N_18251);
and U23476 (N_23476,N_19374,N_19768);
xnor U23477 (N_23477,N_19482,N_20020);
and U23478 (N_23478,N_19244,N_20379);
nand U23479 (N_23479,N_20542,N_18495);
and U23480 (N_23480,N_19826,N_20977);
nor U23481 (N_23481,N_20315,N_20991);
xor U23482 (N_23482,N_20077,N_19000);
xor U23483 (N_23483,N_20268,N_19127);
and U23484 (N_23484,N_19583,N_19890);
or U23485 (N_23485,N_19452,N_18188);
nand U23486 (N_23486,N_20669,N_18701);
or U23487 (N_23487,N_19152,N_20147);
and U23488 (N_23488,N_19806,N_19412);
xnor U23489 (N_23489,N_20903,N_19822);
or U23490 (N_23490,N_18154,N_18594);
nand U23491 (N_23491,N_20810,N_20631);
nor U23492 (N_23492,N_20224,N_19021);
nand U23493 (N_23493,N_20310,N_18693);
nand U23494 (N_23494,N_18709,N_20373);
or U23495 (N_23495,N_18542,N_20944);
and U23496 (N_23496,N_18421,N_19618);
nand U23497 (N_23497,N_18291,N_18133);
and U23498 (N_23498,N_19656,N_19408);
nand U23499 (N_23499,N_18158,N_20895);
and U23500 (N_23500,N_18161,N_20423);
nor U23501 (N_23501,N_19456,N_19780);
xor U23502 (N_23502,N_18609,N_19928);
nor U23503 (N_23503,N_19546,N_19725);
and U23504 (N_23504,N_18530,N_20884);
or U23505 (N_23505,N_20064,N_18409);
and U23506 (N_23506,N_19147,N_18276);
or U23507 (N_23507,N_18319,N_19490);
and U23508 (N_23508,N_18414,N_18080);
nand U23509 (N_23509,N_18520,N_18644);
xnor U23510 (N_23510,N_19434,N_18112);
xor U23511 (N_23511,N_20390,N_20363);
nand U23512 (N_23512,N_20974,N_18504);
xor U23513 (N_23513,N_20782,N_18953);
and U23514 (N_23514,N_18196,N_19238);
nand U23515 (N_23515,N_19320,N_18120);
nor U23516 (N_23516,N_19755,N_19166);
nor U23517 (N_23517,N_18144,N_18407);
and U23518 (N_23518,N_20394,N_18796);
nand U23519 (N_23519,N_19365,N_19875);
nor U23520 (N_23520,N_20698,N_20447);
or U23521 (N_23521,N_19431,N_18734);
xor U23522 (N_23522,N_19665,N_18359);
nand U23523 (N_23523,N_20671,N_19245);
nor U23524 (N_23524,N_20861,N_18675);
nand U23525 (N_23525,N_18643,N_18610);
nor U23526 (N_23526,N_19880,N_19385);
nand U23527 (N_23527,N_18926,N_18443);
and U23528 (N_23528,N_19852,N_19675);
xnor U23529 (N_23529,N_18263,N_20737);
or U23530 (N_23530,N_19517,N_18000);
nor U23531 (N_23531,N_19774,N_18564);
or U23532 (N_23532,N_19828,N_18956);
and U23533 (N_23533,N_20615,N_20602);
or U23534 (N_23534,N_18230,N_19886);
nor U23535 (N_23535,N_20606,N_19137);
or U23536 (N_23536,N_20397,N_19752);
or U23537 (N_23537,N_20867,N_20303);
or U23538 (N_23538,N_19111,N_18848);
nor U23539 (N_23539,N_20361,N_18082);
nor U23540 (N_23540,N_19517,N_20679);
and U23541 (N_23541,N_19474,N_20641);
or U23542 (N_23542,N_19392,N_20877);
nor U23543 (N_23543,N_18235,N_19125);
nor U23544 (N_23544,N_18182,N_18175);
or U23545 (N_23545,N_19812,N_18992);
xnor U23546 (N_23546,N_19266,N_20397);
or U23547 (N_23547,N_19414,N_19076);
or U23548 (N_23548,N_18259,N_18126);
or U23549 (N_23549,N_20010,N_20646);
or U23550 (N_23550,N_18453,N_19049);
xnor U23551 (N_23551,N_19828,N_20482);
xor U23552 (N_23552,N_19733,N_20643);
nand U23553 (N_23553,N_18074,N_19539);
nor U23554 (N_23554,N_18423,N_20673);
and U23555 (N_23555,N_18293,N_18132);
or U23556 (N_23556,N_18796,N_19162);
and U23557 (N_23557,N_19115,N_18123);
and U23558 (N_23558,N_20746,N_19741);
nor U23559 (N_23559,N_20888,N_19535);
nand U23560 (N_23560,N_20424,N_19981);
nor U23561 (N_23561,N_19644,N_19472);
nand U23562 (N_23562,N_19328,N_19662);
or U23563 (N_23563,N_18882,N_20275);
and U23564 (N_23564,N_18572,N_18136);
and U23565 (N_23565,N_20976,N_19093);
and U23566 (N_23566,N_20863,N_19731);
or U23567 (N_23567,N_19440,N_18982);
nor U23568 (N_23568,N_19077,N_18772);
nor U23569 (N_23569,N_20670,N_19803);
nor U23570 (N_23570,N_18692,N_18372);
nor U23571 (N_23571,N_20984,N_18638);
or U23572 (N_23572,N_19225,N_19726);
nand U23573 (N_23573,N_18890,N_18891);
nor U23574 (N_23574,N_19791,N_18919);
xnor U23575 (N_23575,N_20321,N_19701);
nor U23576 (N_23576,N_20414,N_19273);
or U23577 (N_23577,N_20669,N_19730);
xor U23578 (N_23578,N_18685,N_19970);
nor U23579 (N_23579,N_20218,N_18651);
or U23580 (N_23580,N_18322,N_19050);
nor U23581 (N_23581,N_19793,N_18990);
and U23582 (N_23582,N_19357,N_18080);
nor U23583 (N_23583,N_20545,N_20522);
xor U23584 (N_23584,N_20858,N_20845);
nand U23585 (N_23585,N_19869,N_18327);
nor U23586 (N_23586,N_20916,N_20398);
xor U23587 (N_23587,N_20565,N_19155);
nor U23588 (N_23588,N_19175,N_20709);
nor U23589 (N_23589,N_18120,N_20470);
xor U23590 (N_23590,N_18868,N_20830);
and U23591 (N_23591,N_18140,N_18559);
or U23592 (N_23592,N_18809,N_20912);
and U23593 (N_23593,N_20902,N_20229);
xor U23594 (N_23594,N_18334,N_18848);
nor U23595 (N_23595,N_20642,N_20374);
xnor U23596 (N_23596,N_19345,N_18974);
xor U23597 (N_23597,N_19917,N_18454);
and U23598 (N_23598,N_20604,N_19158);
or U23599 (N_23599,N_20286,N_20717);
nor U23600 (N_23600,N_19255,N_20370);
or U23601 (N_23601,N_20147,N_18337);
or U23602 (N_23602,N_18366,N_19022);
xnor U23603 (N_23603,N_18069,N_20104);
or U23604 (N_23604,N_19621,N_20990);
and U23605 (N_23605,N_20943,N_19006);
or U23606 (N_23606,N_19716,N_19886);
nand U23607 (N_23607,N_18993,N_18756);
and U23608 (N_23608,N_20437,N_18133);
xnor U23609 (N_23609,N_20947,N_18399);
nor U23610 (N_23610,N_20688,N_19927);
xnor U23611 (N_23611,N_19836,N_19294);
xnor U23612 (N_23612,N_19916,N_18493);
or U23613 (N_23613,N_20272,N_19898);
nor U23614 (N_23614,N_19154,N_18280);
or U23615 (N_23615,N_20298,N_19370);
nand U23616 (N_23616,N_18855,N_18140);
and U23617 (N_23617,N_19428,N_18552);
nor U23618 (N_23618,N_19115,N_19442);
xor U23619 (N_23619,N_18903,N_19880);
xnor U23620 (N_23620,N_18384,N_19223);
xor U23621 (N_23621,N_19793,N_18769);
and U23622 (N_23622,N_19156,N_20511);
xor U23623 (N_23623,N_20711,N_20293);
xnor U23624 (N_23624,N_18445,N_20763);
nor U23625 (N_23625,N_20731,N_20770);
nand U23626 (N_23626,N_20692,N_20847);
or U23627 (N_23627,N_19087,N_20485);
xnor U23628 (N_23628,N_20589,N_20226);
nand U23629 (N_23629,N_19177,N_18228);
or U23630 (N_23630,N_20100,N_19423);
or U23631 (N_23631,N_18265,N_19208);
xnor U23632 (N_23632,N_18421,N_20313);
or U23633 (N_23633,N_19873,N_19946);
and U23634 (N_23634,N_18748,N_20834);
and U23635 (N_23635,N_20874,N_18982);
nor U23636 (N_23636,N_18207,N_18539);
nand U23637 (N_23637,N_19165,N_20384);
or U23638 (N_23638,N_20210,N_20830);
or U23639 (N_23639,N_19993,N_18317);
and U23640 (N_23640,N_18497,N_18958);
xnor U23641 (N_23641,N_19208,N_19183);
nor U23642 (N_23642,N_18840,N_20250);
and U23643 (N_23643,N_19281,N_20488);
xor U23644 (N_23644,N_18947,N_19045);
or U23645 (N_23645,N_18873,N_18197);
xnor U23646 (N_23646,N_20114,N_19685);
and U23647 (N_23647,N_18838,N_19583);
xor U23648 (N_23648,N_20326,N_18118);
nor U23649 (N_23649,N_19071,N_19562);
xor U23650 (N_23650,N_18314,N_18047);
nor U23651 (N_23651,N_18159,N_19550);
nor U23652 (N_23652,N_20220,N_18200);
and U23653 (N_23653,N_19142,N_20077);
xor U23654 (N_23654,N_20269,N_19515);
nand U23655 (N_23655,N_18263,N_19097);
nand U23656 (N_23656,N_20828,N_18106);
or U23657 (N_23657,N_19028,N_20911);
nor U23658 (N_23658,N_19238,N_18476);
nand U23659 (N_23659,N_19944,N_19198);
nand U23660 (N_23660,N_20774,N_19365);
nand U23661 (N_23661,N_20201,N_19340);
xnor U23662 (N_23662,N_18354,N_20366);
nor U23663 (N_23663,N_18003,N_19189);
nand U23664 (N_23664,N_19966,N_18487);
nand U23665 (N_23665,N_18661,N_18702);
and U23666 (N_23666,N_20812,N_20479);
xnor U23667 (N_23667,N_18818,N_20018);
nand U23668 (N_23668,N_18601,N_18917);
nand U23669 (N_23669,N_18122,N_19328);
nor U23670 (N_23670,N_18325,N_18759);
xor U23671 (N_23671,N_20106,N_18320);
nand U23672 (N_23672,N_18030,N_18727);
nor U23673 (N_23673,N_18451,N_20062);
xor U23674 (N_23674,N_19440,N_20690);
nand U23675 (N_23675,N_19806,N_19391);
and U23676 (N_23676,N_19657,N_20620);
nand U23677 (N_23677,N_19561,N_19227);
xnor U23678 (N_23678,N_19278,N_18806);
nor U23679 (N_23679,N_18213,N_18360);
xnor U23680 (N_23680,N_20546,N_20290);
and U23681 (N_23681,N_20429,N_18267);
nor U23682 (N_23682,N_19154,N_18479);
xnor U23683 (N_23683,N_20585,N_19790);
nand U23684 (N_23684,N_20055,N_19480);
nand U23685 (N_23685,N_18768,N_19635);
nor U23686 (N_23686,N_20840,N_20908);
and U23687 (N_23687,N_18411,N_20194);
xnor U23688 (N_23688,N_18469,N_18402);
xnor U23689 (N_23689,N_19147,N_18993);
or U23690 (N_23690,N_19242,N_20411);
nor U23691 (N_23691,N_18917,N_19454);
and U23692 (N_23692,N_18867,N_18100);
nand U23693 (N_23693,N_20125,N_18670);
nor U23694 (N_23694,N_18657,N_18165);
and U23695 (N_23695,N_20203,N_20120);
nor U23696 (N_23696,N_18229,N_19994);
and U23697 (N_23697,N_18961,N_18994);
xor U23698 (N_23698,N_19772,N_18684);
and U23699 (N_23699,N_18244,N_18295);
xor U23700 (N_23700,N_19950,N_19827);
nor U23701 (N_23701,N_18966,N_19592);
xnor U23702 (N_23702,N_20941,N_19967);
xor U23703 (N_23703,N_20364,N_19701);
xor U23704 (N_23704,N_20756,N_18990);
nand U23705 (N_23705,N_18732,N_19117);
xnor U23706 (N_23706,N_19720,N_18153);
nand U23707 (N_23707,N_18245,N_20354);
or U23708 (N_23708,N_18014,N_19615);
and U23709 (N_23709,N_19157,N_18039);
xnor U23710 (N_23710,N_18290,N_18621);
nand U23711 (N_23711,N_20887,N_19646);
xor U23712 (N_23712,N_20844,N_18767);
or U23713 (N_23713,N_20242,N_20423);
or U23714 (N_23714,N_19960,N_20757);
or U23715 (N_23715,N_20453,N_20377);
nor U23716 (N_23716,N_18476,N_18527);
or U23717 (N_23717,N_18719,N_19040);
nand U23718 (N_23718,N_19185,N_19411);
xor U23719 (N_23719,N_18959,N_19393);
xnor U23720 (N_23720,N_18818,N_18640);
or U23721 (N_23721,N_18770,N_20735);
nand U23722 (N_23722,N_18787,N_19486);
and U23723 (N_23723,N_18177,N_18012);
nor U23724 (N_23724,N_18558,N_18454);
nor U23725 (N_23725,N_18696,N_20306);
nand U23726 (N_23726,N_18761,N_19547);
nand U23727 (N_23727,N_19849,N_20057);
xnor U23728 (N_23728,N_18724,N_19111);
or U23729 (N_23729,N_20028,N_19396);
nor U23730 (N_23730,N_19786,N_20993);
and U23731 (N_23731,N_18706,N_19834);
nor U23732 (N_23732,N_19507,N_18497);
and U23733 (N_23733,N_20989,N_19481);
nand U23734 (N_23734,N_18893,N_19206);
and U23735 (N_23735,N_20977,N_20691);
nand U23736 (N_23736,N_20313,N_19929);
nor U23737 (N_23737,N_18336,N_18887);
and U23738 (N_23738,N_19331,N_19694);
nor U23739 (N_23739,N_18451,N_18565);
and U23740 (N_23740,N_19164,N_20255);
xnor U23741 (N_23741,N_20920,N_19382);
xnor U23742 (N_23742,N_18229,N_18572);
or U23743 (N_23743,N_18911,N_19694);
nor U23744 (N_23744,N_18635,N_19549);
or U23745 (N_23745,N_19067,N_20882);
nand U23746 (N_23746,N_18970,N_18376);
xor U23747 (N_23747,N_18984,N_19254);
and U23748 (N_23748,N_19963,N_18633);
nor U23749 (N_23749,N_20282,N_20610);
or U23750 (N_23750,N_20395,N_19043);
xnor U23751 (N_23751,N_18651,N_19365);
and U23752 (N_23752,N_18234,N_20903);
and U23753 (N_23753,N_20422,N_18456);
nor U23754 (N_23754,N_20522,N_20514);
nand U23755 (N_23755,N_19302,N_18300);
xor U23756 (N_23756,N_19509,N_20483);
xnor U23757 (N_23757,N_18879,N_20031);
or U23758 (N_23758,N_18928,N_19237);
nand U23759 (N_23759,N_19334,N_18586);
or U23760 (N_23760,N_19453,N_18274);
nand U23761 (N_23761,N_19827,N_19983);
nor U23762 (N_23762,N_20344,N_18586);
or U23763 (N_23763,N_18476,N_20941);
xnor U23764 (N_23764,N_19214,N_18027);
xor U23765 (N_23765,N_18876,N_19258);
nand U23766 (N_23766,N_18955,N_20361);
or U23767 (N_23767,N_20518,N_20243);
or U23768 (N_23768,N_20266,N_20499);
nor U23769 (N_23769,N_19569,N_18026);
xor U23770 (N_23770,N_20765,N_18195);
nor U23771 (N_23771,N_19897,N_20354);
and U23772 (N_23772,N_20101,N_20884);
and U23773 (N_23773,N_20405,N_18582);
nor U23774 (N_23774,N_20464,N_19161);
xnor U23775 (N_23775,N_20266,N_19360);
and U23776 (N_23776,N_20550,N_19774);
nand U23777 (N_23777,N_20563,N_18857);
xnor U23778 (N_23778,N_20884,N_19869);
nor U23779 (N_23779,N_19546,N_20988);
and U23780 (N_23780,N_18524,N_18240);
or U23781 (N_23781,N_18028,N_18586);
nand U23782 (N_23782,N_18745,N_19413);
or U23783 (N_23783,N_18066,N_20607);
and U23784 (N_23784,N_20960,N_19416);
nor U23785 (N_23785,N_20263,N_18235);
and U23786 (N_23786,N_20518,N_18469);
and U23787 (N_23787,N_20871,N_18446);
or U23788 (N_23788,N_20271,N_20942);
or U23789 (N_23789,N_19888,N_20179);
nand U23790 (N_23790,N_18223,N_20343);
and U23791 (N_23791,N_18838,N_18406);
and U23792 (N_23792,N_20072,N_18941);
nand U23793 (N_23793,N_18209,N_20091);
or U23794 (N_23794,N_18958,N_18923);
and U23795 (N_23795,N_18460,N_19327);
nand U23796 (N_23796,N_20094,N_18476);
nand U23797 (N_23797,N_18279,N_20112);
or U23798 (N_23798,N_18869,N_19421);
nand U23799 (N_23799,N_18934,N_18174);
or U23800 (N_23800,N_18086,N_20155);
xor U23801 (N_23801,N_19370,N_19591);
xor U23802 (N_23802,N_18542,N_20417);
xor U23803 (N_23803,N_20411,N_19562);
nor U23804 (N_23804,N_20812,N_20263);
nand U23805 (N_23805,N_19648,N_19007);
and U23806 (N_23806,N_18580,N_18910);
nand U23807 (N_23807,N_18307,N_19538);
and U23808 (N_23808,N_18711,N_20664);
nand U23809 (N_23809,N_20449,N_20376);
and U23810 (N_23810,N_19922,N_20019);
xnor U23811 (N_23811,N_18689,N_19497);
nor U23812 (N_23812,N_18615,N_20869);
and U23813 (N_23813,N_20438,N_19053);
or U23814 (N_23814,N_18176,N_18844);
xnor U23815 (N_23815,N_19411,N_18286);
and U23816 (N_23816,N_19346,N_20498);
or U23817 (N_23817,N_20494,N_19989);
nand U23818 (N_23818,N_20966,N_19598);
nand U23819 (N_23819,N_18448,N_18643);
or U23820 (N_23820,N_20066,N_19641);
or U23821 (N_23821,N_18931,N_18807);
nor U23822 (N_23822,N_20437,N_20816);
or U23823 (N_23823,N_18351,N_19741);
xor U23824 (N_23824,N_18043,N_20783);
or U23825 (N_23825,N_18873,N_20044);
and U23826 (N_23826,N_18609,N_19319);
and U23827 (N_23827,N_18167,N_18052);
xnor U23828 (N_23828,N_18425,N_20006);
and U23829 (N_23829,N_20345,N_20082);
nand U23830 (N_23830,N_19333,N_18088);
nand U23831 (N_23831,N_18876,N_19896);
nor U23832 (N_23832,N_18271,N_20014);
nor U23833 (N_23833,N_18275,N_20194);
nand U23834 (N_23834,N_20739,N_18497);
xor U23835 (N_23835,N_20467,N_18187);
nand U23836 (N_23836,N_19050,N_19470);
xnor U23837 (N_23837,N_20651,N_20761);
xnor U23838 (N_23838,N_18003,N_19959);
or U23839 (N_23839,N_20871,N_18632);
or U23840 (N_23840,N_19697,N_18959);
nand U23841 (N_23841,N_18228,N_20433);
nand U23842 (N_23842,N_19180,N_18113);
xnor U23843 (N_23843,N_19627,N_19545);
nor U23844 (N_23844,N_19940,N_19771);
or U23845 (N_23845,N_20114,N_19323);
nand U23846 (N_23846,N_20129,N_20994);
and U23847 (N_23847,N_19672,N_19360);
nand U23848 (N_23848,N_18958,N_18708);
or U23849 (N_23849,N_19964,N_18869);
nand U23850 (N_23850,N_18583,N_20148);
nor U23851 (N_23851,N_18085,N_18905);
nand U23852 (N_23852,N_19210,N_20440);
or U23853 (N_23853,N_20451,N_18880);
and U23854 (N_23854,N_19694,N_19263);
nand U23855 (N_23855,N_20127,N_18176);
or U23856 (N_23856,N_18706,N_18750);
xor U23857 (N_23857,N_18780,N_18885);
and U23858 (N_23858,N_20433,N_19449);
nor U23859 (N_23859,N_19891,N_20281);
nand U23860 (N_23860,N_20561,N_18737);
xnor U23861 (N_23861,N_18716,N_20076);
and U23862 (N_23862,N_18523,N_18786);
nand U23863 (N_23863,N_19681,N_19080);
nand U23864 (N_23864,N_18959,N_19993);
nor U23865 (N_23865,N_20464,N_20535);
or U23866 (N_23866,N_20718,N_19976);
and U23867 (N_23867,N_18402,N_19915);
nand U23868 (N_23868,N_18286,N_19718);
and U23869 (N_23869,N_20746,N_20876);
or U23870 (N_23870,N_20318,N_19725);
nor U23871 (N_23871,N_19545,N_20808);
or U23872 (N_23872,N_19385,N_19254);
and U23873 (N_23873,N_20532,N_19657);
xor U23874 (N_23874,N_20641,N_18530);
and U23875 (N_23875,N_20518,N_20265);
xnor U23876 (N_23876,N_19292,N_18762);
or U23877 (N_23877,N_19292,N_18435);
nor U23878 (N_23878,N_19685,N_19998);
and U23879 (N_23879,N_20157,N_19842);
nor U23880 (N_23880,N_19801,N_18528);
or U23881 (N_23881,N_18929,N_18159);
or U23882 (N_23882,N_19460,N_18290);
and U23883 (N_23883,N_19373,N_18606);
or U23884 (N_23884,N_18344,N_18992);
nor U23885 (N_23885,N_20178,N_19954);
xor U23886 (N_23886,N_20883,N_19372);
nor U23887 (N_23887,N_20849,N_20758);
xor U23888 (N_23888,N_19236,N_20294);
and U23889 (N_23889,N_19116,N_20604);
xor U23890 (N_23890,N_18185,N_20347);
nor U23891 (N_23891,N_19037,N_18858);
xnor U23892 (N_23892,N_18963,N_18931);
nor U23893 (N_23893,N_19800,N_18302);
nor U23894 (N_23894,N_18017,N_19458);
nand U23895 (N_23895,N_20564,N_18876);
and U23896 (N_23896,N_18534,N_19695);
nand U23897 (N_23897,N_18504,N_19542);
nor U23898 (N_23898,N_19579,N_19628);
and U23899 (N_23899,N_19159,N_18360);
nor U23900 (N_23900,N_19862,N_18401);
xnor U23901 (N_23901,N_18724,N_19018);
xor U23902 (N_23902,N_20141,N_18894);
nor U23903 (N_23903,N_20737,N_20311);
nor U23904 (N_23904,N_19606,N_19077);
xor U23905 (N_23905,N_19195,N_18638);
nor U23906 (N_23906,N_19517,N_19240);
or U23907 (N_23907,N_19314,N_20005);
nand U23908 (N_23908,N_19110,N_19971);
and U23909 (N_23909,N_19707,N_20314);
and U23910 (N_23910,N_19854,N_19475);
xnor U23911 (N_23911,N_20054,N_20412);
and U23912 (N_23912,N_20006,N_20881);
nand U23913 (N_23913,N_19464,N_19953);
nand U23914 (N_23914,N_19035,N_18358);
nor U23915 (N_23915,N_19896,N_18330);
and U23916 (N_23916,N_20111,N_20485);
or U23917 (N_23917,N_18676,N_19646);
xnor U23918 (N_23918,N_18930,N_20589);
nand U23919 (N_23919,N_18087,N_18841);
xnor U23920 (N_23920,N_20829,N_18569);
nor U23921 (N_23921,N_19480,N_19259);
nor U23922 (N_23922,N_18760,N_19258);
nand U23923 (N_23923,N_18412,N_18865);
nand U23924 (N_23924,N_19680,N_18898);
nor U23925 (N_23925,N_19246,N_20370);
and U23926 (N_23926,N_18301,N_20000);
nor U23927 (N_23927,N_18911,N_20720);
and U23928 (N_23928,N_19997,N_19474);
nand U23929 (N_23929,N_19355,N_18300);
nor U23930 (N_23930,N_20733,N_20346);
xor U23931 (N_23931,N_18181,N_19967);
nor U23932 (N_23932,N_19033,N_20931);
and U23933 (N_23933,N_20515,N_19661);
nand U23934 (N_23934,N_18717,N_18264);
or U23935 (N_23935,N_18049,N_19113);
and U23936 (N_23936,N_19654,N_20057);
or U23937 (N_23937,N_18394,N_19325);
and U23938 (N_23938,N_19048,N_19688);
xor U23939 (N_23939,N_19292,N_19063);
and U23940 (N_23940,N_20152,N_19705);
or U23941 (N_23941,N_20046,N_20806);
nand U23942 (N_23942,N_19500,N_18238);
xor U23943 (N_23943,N_19261,N_19688);
or U23944 (N_23944,N_19572,N_18233);
xnor U23945 (N_23945,N_19009,N_19379);
or U23946 (N_23946,N_18188,N_20458);
and U23947 (N_23947,N_20752,N_18821);
xor U23948 (N_23948,N_19609,N_18679);
and U23949 (N_23949,N_20373,N_20307);
and U23950 (N_23950,N_18835,N_18817);
and U23951 (N_23951,N_18635,N_19136);
xnor U23952 (N_23952,N_19699,N_19706);
or U23953 (N_23953,N_20086,N_18840);
nor U23954 (N_23954,N_19423,N_18233);
nand U23955 (N_23955,N_20417,N_20776);
xnor U23956 (N_23956,N_20437,N_19638);
nand U23957 (N_23957,N_20301,N_18749);
and U23958 (N_23958,N_18455,N_19637);
nand U23959 (N_23959,N_20159,N_19729);
nor U23960 (N_23960,N_19905,N_20839);
and U23961 (N_23961,N_18413,N_20002);
xnor U23962 (N_23962,N_20269,N_18289);
xor U23963 (N_23963,N_19817,N_20566);
and U23964 (N_23964,N_19293,N_19035);
nor U23965 (N_23965,N_18212,N_19241);
nand U23966 (N_23966,N_20001,N_20639);
nand U23967 (N_23967,N_19907,N_20268);
nand U23968 (N_23968,N_20035,N_18886);
nor U23969 (N_23969,N_18679,N_19210);
nor U23970 (N_23970,N_19242,N_19747);
and U23971 (N_23971,N_19583,N_20934);
nor U23972 (N_23972,N_20408,N_19224);
nor U23973 (N_23973,N_19599,N_19516);
nand U23974 (N_23974,N_20904,N_18918);
xor U23975 (N_23975,N_20419,N_18959);
xnor U23976 (N_23976,N_20076,N_19300);
and U23977 (N_23977,N_18881,N_20670);
xnor U23978 (N_23978,N_19206,N_18881);
nand U23979 (N_23979,N_20943,N_20463);
or U23980 (N_23980,N_20711,N_20166);
nor U23981 (N_23981,N_18072,N_19788);
nor U23982 (N_23982,N_18019,N_18980);
nor U23983 (N_23983,N_20958,N_20418);
nand U23984 (N_23984,N_19203,N_19160);
and U23985 (N_23985,N_19526,N_18780);
xnor U23986 (N_23986,N_20424,N_20884);
or U23987 (N_23987,N_19112,N_19543);
nor U23988 (N_23988,N_20060,N_18343);
nand U23989 (N_23989,N_20827,N_19756);
and U23990 (N_23990,N_19403,N_19095);
and U23991 (N_23991,N_20249,N_18876);
nand U23992 (N_23992,N_20350,N_19794);
nor U23993 (N_23993,N_19549,N_18178);
nand U23994 (N_23994,N_19516,N_18530);
xnor U23995 (N_23995,N_19948,N_18065);
and U23996 (N_23996,N_18738,N_19251);
nand U23997 (N_23997,N_19021,N_18115);
and U23998 (N_23998,N_18691,N_20816);
or U23999 (N_23999,N_19843,N_20980);
and U24000 (N_24000,N_21806,N_23509);
nor U24001 (N_24001,N_21537,N_21319);
nand U24002 (N_24002,N_21487,N_23914);
nor U24003 (N_24003,N_21950,N_23792);
xor U24004 (N_24004,N_21168,N_21101);
xor U24005 (N_24005,N_22502,N_22302);
nand U24006 (N_24006,N_21780,N_23584);
or U24007 (N_24007,N_23888,N_21332);
nor U24008 (N_24008,N_21540,N_22402);
nand U24009 (N_24009,N_21027,N_23678);
xor U24010 (N_24010,N_21561,N_22681);
nor U24011 (N_24011,N_23111,N_22359);
nor U24012 (N_24012,N_21461,N_21276);
nor U24013 (N_24013,N_22065,N_23169);
xor U24014 (N_24014,N_22441,N_21630);
xor U24015 (N_24015,N_21569,N_23104);
and U24016 (N_24016,N_22121,N_21883);
and U24017 (N_24017,N_21170,N_22588);
nand U24018 (N_24018,N_23322,N_23839);
or U24019 (N_24019,N_23347,N_23101);
and U24020 (N_24020,N_22711,N_23125);
nor U24021 (N_24021,N_23773,N_23410);
nand U24022 (N_24022,N_23036,N_21703);
or U24023 (N_24023,N_21909,N_21894);
xor U24024 (N_24024,N_22244,N_22025);
or U24025 (N_24025,N_21896,N_22089);
nand U24026 (N_24026,N_23966,N_21103);
nor U24027 (N_24027,N_21667,N_23129);
nand U24028 (N_24028,N_22592,N_22717);
nand U24029 (N_24029,N_21681,N_23687);
nand U24030 (N_24030,N_21543,N_22564);
or U24031 (N_24031,N_21545,N_23569);
xor U24032 (N_24032,N_22611,N_23699);
xnor U24033 (N_24033,N_22078,N_21732);
xnor U24034 (N_24034,N_22801,N_21824);
or U24035 (N_24035,N_22267,N_21660);
nor U24036 (N_24036,N_22428,N_23901);
and U24037 (N_24037,N_21081,N_21707);
and U24038 (N_24038,N_23124,N_21311);
nand U24039 (N_24039,N_22511,N_23818);
nor U24040 (N_24040,N_23988,N_23740);
or U24041 (N_24041,N_21893,N_22173);
nand U24042 (N_24042,N_23619,N_22756);
nor U24043 (N_24043,N_21375,N_23995);
and U24044 (N_24044,N_22882,N_22258);
nor U24045 (N_24045,N_22182,N_21699);
xnor U24046 (N_24046,N_23334,N_23644);
or U24047 (N_24047,N_22817,N_22016);
nor U24048 (N_24048,N_22687,N_21470);
nand U24049 (N_24049,N_23099,N_23607);
xnor U24050 (N_24050,N_23498,N_22480);
and U24051 (N_24051,N_21271,N_22532);
xnor U24052 (N_24052,N_22591,N_23365);
xnor U24053 (N_24053,N_23010,N_22674);
xnor U24054 (N_24054,N_21614,N_22630);
and U24055 (N_24055,N_23208,N_21078);
xor U24056 (N_24056,N_22038,N_22180);
and U24057 (N_24057,N_22160,N_23374);
nand U24058 (N_24058,N_21558,N_21826);
nand U24059 (N_24059,N_22238,N_22645);
or U24060 (N_24060,N_22922,N_22221);
nor U24061 (N_24061,N_23028,N_21257);
nand U24062 (N_24062,N_23952,N_22654);
nor U24063 (N_24063,N_23603,N_22587);
nor U24064 (N_24064,N_22789,N_21121);
nand U24065 (N_24065,N_21600,N_21258);
and U24066 (N_24066,N_21165,N_21798);
nor U24067 (N_24067,N_23331,N_21821);
nand U24068 (N_24068,N_21739,N_23568);
or U24069 (N_24069,N_22603,N_21546);
and U24070 (N_24070,N_23034,N_23395);
xnor U24071 (N_24071,N_23711,N_22014);
and U24072 (N_24072,N_22708,N_22570);
xnor U24073 (N_24073,N_22279,N_23944);
or U24074 (N_24074,N_21178,N_21035);
and U24075 (N_24075,N_21900,N_22100);
nand U24076 (N_24076,N_21716,N_23146);
xnor U24077 (N_24077,N_22518,N_21518);
and U24078 (N_24078,N_23704,N_21992);
nand U24079 (N_24079,N_23978,N_22757);
or U24080 (N_24080,N_23590,N_21326);
and U24081 (N_24081,N_22350,N_23192);
nor U24082 (N_24082,N_23795,N_21337);
and U24083 (N_24083,N_22577,N_23135);
and U24084 (N_24084,N_22977,N_22211);
nor U24085 (N_24085,N_23548,N_22522);
nand U24086 (N_24086,N_22585,N_22928);
or U24087 (N_24087,N_22019,N_23244);
and U24088 (N_24088,N_22872,N_23237);
or U24089 (N_24089,N_23726,N_22155);
nor U24090 (N_24090,N_21901,N_21683);
xnor U24091 (N_24091,N_23522,N_22675);
xor U24092 (N_24092,N_23179,N_22622);
nor U24093 (N_24093,N_22635,N_22933);
and U24094 (N_24094,N_21757,N_23817);
or U24095 (N_24095,N_22519,N_23758);
or U24096 (N_24096,N_22444,N_23965);
or U24097 (N_24097,N_21570,N_23381);
and U24098 (N_24098,N_22209,N_22356);
and U24099 (N_24099,N_21316,N_21512);
nor U24100 (N_24100,N_21046,N_22056);
xnor U24101 (N_24101,N_22462,N_22573);
or U24102 (N_24102,N_22252,N_21483);
nor U24103 (N_24103,N_23149,N_23656);
or U24104 (N_24104,N_23930,N_23318);
or U24105 (N_24105,N_22979,N_23187);
nor U24106 (N_24106,N_22669,N_23885);
and U24107 (N_24107,N_22305,N_22030);
xnor U24108 (N_24108,N_22138,N_22855);
nor U24109 (N_24109,N_23462,N_23132);
or U24110 (N_24110,N_23575,N_23855);
or U24111 (N_24111,N_22317,N_21008);
and U24112 (N_24112,N_21553,N_22994);
or U24113 (N_24113,N_22957,N_21188);
and U24114 (N_24114,N_21997,N_23642);
nand U24115 (N_24115,N_22796,N_23542);
nand U24116 (N_24116,N_21535,N_23653);
or U24117 (N_24117,N_23130,N_21669);
and U24118 (N_24118,N_22710,N_23892);
and U24119 (N_24119,N_21599,N_22720);
or U24120 (N_24120,N_22142,N_21364);
and U24121 (N_24121,N_21231,N_23880);
and U24122 (N_24122,N_21787,N_22364);
and U24123 (N_24123,N_21639,N_22501);
or U24124 (N_24124,N_22257,N_22672);
xnor U24125 (N_24125,N_21583,N_21576);
and U24126 (N_24126,N_21864,N_22561);
nand U24127 (N_24127,N_22046,N_21814);
xor U24128 (N_24128,N_21084,N_22240);
nand U24129 (N_24129,N_22540,N_23985);
nand U24130 (N_24130,N_23161,N_22090);
nand U24131 (N_24131,N_23730,N_22083);
and U24132 (N_24132,N_22960,N_23241);
nor U24133 (N_24133,N_23386,N_23434);
and U24134 (N_24134,N_21209,N_21175);
xor U24135 (N_24135,N_22490,N_21176);
nand U24136 (N_24136,N_23001,N_23211);
xor U24137 (N_24137,N_22133,N_22880);
nand U24138 (N_24138,N_22907,N_22772);
nor U24139 (N_24139,N_23765,N_23538);
nor U24140 (N_24140,N_23108,N_22651);
or U24141 (N_24141,N_23442,N_23634);
xor U24142 (N_24142,N_23706,N_21465);
or U24143 (N_24143,N_22066,N_21080);
or U24144 (N_24144,N_21056,N_21898);
nor U24145 (N_24145,N_22218,N_21714);
and U24146 (N_24146,N_21542,N_22311);
nor U24147 (N_24147,N_23759,N_22120);
nand U24148 (N_24148,N_21781,N_21376);
nand U24149 (N_24149,N_23513,N_21734);
nand U24150 (N_24150,N_21162,N_22321);
xnor U24151 (N_24151,N_21579,N_22262);
nor U24152 (N_24152,N_21194,N_21827);
xnor U24153 (N_24153,N_23891,N_21857);
nand U24154 (N_24154,N_22164,N_21264);
nand U24155 (N_24155,N_21142,N_22354);
or U24156 (N_24156,N_22981,N_22528);
xor U24157 (N_24157,N_21010,N_22600);
nor U24158 (N_24158,N_23763,N_23629);
nor U24159 (N_24159,N_21448,N_23025);
and U24160 (N_24160,N_21661,N_23646);
or U24161 (N_24161,N_23874,N_23554);
nand U24162 (N_24162,N_22068,N_23577);
nor U24163 (N_24163,N_21832,N_22741);
nand U24164 (N_24164,N_23037,N_23677);
xnor U24165 (N_24165,N_23981,N_23591);
nand U24166 (N_24166,N_22166,N_22470);
and U24167 (N_24167,N_21708,N_21947);
or U24168 (N_24168,N_22202,N_22483);
nand U24169 (N_24169,N_23326,N_21524);
xor U24170 (N_24170,N_21346,N_21575);
and U24171 (N_24171,N_21874,N_21335);
nand U24172 (N_24172,N_21801,N_23937);
xor U24173 (N_24173,N_22270,N_22963);
or U24174 (N_24174,N_22287,N_23731);
nand U24175 (N_24175,N_23357,N_22123);
and U24176 (N_24176,N_22639,N_23349);
xor U24177 (N_24177,N_23651,N_23540);
xor U24178 (N_24178,N_22558,N_23422);
nor U24179 (N_24179,N_22153,N_22316);
xnor U24180 (N_24180,N_23920,N_22198);
xnor U24181 (N_24181,N_23346,N_21320);
xnor U24182 (N_24182,N_23781,N_21492);
or U24183 (N_24183,N_21970,N_21885);
and U24184 (N_24184,N_22306,N_22011);
nor U24185 (N_24185,N_21899,N_21833);
nor U24186 (N_24186,N_22572,N_22769);
nand U24187 (N_24187,N_21634,N_23481);
nor U24188 (N_24188,N_22498,N_23123);
nor U24189 (N_24189,N_21815,N_21878);
and U24190 (N_24190,N_23964,N_22454);
nand U24191 (N_24191,N_23466,N_22181);
and U24192 (N_24192,N_22278,N_23317);
nor U24193 (N_24193,N_22329,N_22878);
nand U24194 (N_24194,N_21060,N_22831);
xor U24195 (N_24195,N_22952,N_22781);
and U24196 (N_24196,N_22931,N_22885);
or U24197 (N_24197,N_21638,N_22870);
nor U24198 (N_24198,N_21432,N_23243);
nor U24199 (N_24199,N_22103,N_21761);
xor U24200 (N_24200,N_22514,N_21235);
nand U24201 (N_24201,N_21972,N_23446);
and U24202 (N_24202,N_23717,N_21467);
and U24203 (N_24203,N_21534,N_23062);
or U24204 (N_24204,N_21499,N_21834);
nand U24205 (N_24205,N_23269,N_23685);
nand U24206 (N_24206,N_22055,N_23316);
or U24207 (N_24207,N_23040,N_21865);
nor U24208 (N_24208,N_23957,N_23833);
and U24209 (N_24209,N_23770,N_21382);
or U24210 (N_24210,N_21809,N_21582);
nor U24211 (N_24211,N_23048,N_21160);
and U24212 (N_24212,N_21091,N_22666);
or U24213 (N_24213,N_22313,N_23573);
nor U24214 (N_24214,N_23375,N_22367);
or U24215 (N_24215,N_21766,N_22704);
nor U24216 (N_24216,N_23471,N_21895);
nand U24217 (N_24217,N_23339,N_21476);
xnor U24218 (N_24218,N_23368,N_22750);
nand U24219 (N_24219,N_23152,N_22088);
xnor U24220 (N_24220,N_23014,N_22539);
or U24221 (N_24221,N_23093,N_23789);
nor U24222 (N_24222,N_21069,N_23449);
or U24223 (N_24223,N_23004,N_21505);
nor U24224 (N_24224,N_22344,N_23738);
nand U24225 (N_24225,N_22242,N_23098);
nor U24226 (N_24226,N_21184,N_23411);
nand U24227 (N_24227,N_23210,N_23635);
or U24228 (N_24228,N_21636,N_21549);
and U24229 (N_24229,N_23016,N_21632);
xor U24230 (N_24230,N_21641,N_22111);
xor U24231 (N_24231,N_22832,N_23610);
xnor U24232 (N_24232,N_21689,N_21270);
xor U24233 (N_24233,N_21195,N_22076);
xor U24234 (N_24234,N_21125,N_23417);
or U24235 (N_24235,N_21611,N_21064);
and U24236 (N_24236,N_22288,N_23117);
xor U24237 (N_24237,N_23786,N_21233);
and U24238 (N_24238,N_23173,N_22455);
xnor U24239 (N_24239,N_21598,N_21205);
or U24240 (N_24240,N_22226,N_22541);
and U24241 (N_24241,N_22736,N_21528);
nand U24242 (N_24242,N_23259,N_23013);
xor U24243 (N_24243,N_22308,N_23360);
or U24244 (N_24244,N_21890,N_21908);
xor U24245 (N_24245,N_22434,N_21710);
nand U24246 (N_24246,N_21758,N_23332);
nand U24247 (N_24247,N_21265,N_23217);
nand U24248 (N_24248,N_22535,N_23831);
xor U24249 (N_24249,N_22323,N_23068);
nand U24250 (N_24250,N_23131,N_21621);
nor U24251 (N_24251,N_22948,N_23521);
nor U24252 (N_24252,N_21650,N_23837);
and U24253 (N_24253,N_21737,N_21116);
and U24254 (N_24254,N_21665,N_23592);
xnor U24255 (N_24255,N_21808,N_22315);
xor U24256 (N_24256,N_23842,N_22604);
xnor U24257 (N_24257,N_23814,N_23063);
nor U24258 (N_24258,N_23572,N_22524);
xor U24259 (N_24259,N_21988,N_21215);
and U24260 (N_24260,N_23515,N_22951);
or U24261 (N_24261,N_21082,N_22059);
and U24262 (N_24262,N_23799,N_23707);
and U24263 (N_24263,N_21902,N_21007);
nand U24264 (N_24264,N_21656,N_23887);
nor U24265 (N_24265,N_23596,N_23967);
and U24266 (N_24266,N_21717,N_22170);
nor U24267 (N_24267,N_22684,N_22377);
nand U24268 (N_24268,N_23491,N_23444);
nor U24269 (N_24269,N_23119,N_23820);
nor U24270 (N_24270,N_23254,N_21753);
or U24271 (N_24271,N_21799,N_23121);
xor U24272 (N_24272,N_21321,N_23652);
and U24273 (N_24273,N_21419,N_23908);
nand U24274 (N_24274,N_23325,N_22440);
or U24275 (N_24275,N_23432,N_21052);
and U24276 (N_24276,N_23670,N_23497);
nor U24277 (N_24277,N_21214,N_21937);
or U24278 (N_24278,N_22760,N_21243);
and U24279 (N_24279,N_22900,N_23815);
and U24280 (N_24280,N_22326,N_23680);
nor U24281 (N_24281,N_21719,N_21323);
or U24282 (N_24282,N_22521,N_23055);
or U24283 (N_24283,N_23846,N_23045);
xnor U24284 (N_24284,N_23663,N_23660);
xnor U24285 (N_24285,N_22830,N_22447);
nor U24286 (N_24286,N_21230,N_22077);
nor U24287 (N_24287,N_22303,N_21208);
xnor U24288 (N_24288,N_22230,N_22833);
or U24289 (N_24289,N_22212,N_22613);
or U24290 (N_24290,N_22099,N_22340);
nor U24291 (N_24291,N_22775,N_22899);
nand U24292 (N_24292,N_21241,N_23585);
xnor U24293 (N_24293,N_23275,N_23777);
or U24294 (N_24294,N_21429,N_23682);
or U24295 (N_24295,N_23771,N_23945);
nor U24296 (N_24296,N_23485,N_21629);
xor U24297 (N_24297,N_21604,N_21458);
or U24298 (N_24298,N_23936,N_23774);
xor U24299 (N_24299,N_22399,N_21106);
and U24300 (N_24300,N_21526,N_21395);
and U24301 (N_24301,N_21880,N_22538);
or U24302 (N_24302,N_21314,N_23484);
nand U24303 (N_24303,N_22475,N_22752);
nand U24304 (N_24304,N_21502,N_23293);
nor U24305 (N_24305,N_22962,N_21450);
nand U24306 (N_24306,N_21481,N_21181);
or U24307 (N_24307,N_22877,N_21498);
and U24308 (N_24308,N_23746,N_23654);
nand U24309 (N_24309,N_21401,N_22837);
xor U24310 (N_24310,N_23595,N_21562);
or U24311 (N_24311,N_22840,N_23066);
nor U24312 (N_24312,N_22567,N_21519);
or U24313 (N_24313,N_21515,N_22274);
or U24314 (N_24314,N_22887,N_21559);
and U24315 (N_24315,N_22777,N_23718);
nand U24316 (N_24316,N_22964,N_22894);
xnor U24317 (N_24317,N_22730,N_21643);
and U24318 (N_24318,N_21507,N_23089);
or U24319 (N_24319,N_22466,N_23379);
or U24320 (N_24320,N_21642,N_22966);
xnor U24321 (N_24321,N_22512,N_23180);
xor U24322 (N_24322,N_23313,N_23396);
nand U24323 (N_24323,N_22488,N_23252);
nor U24324 (N_24324,N_22905,N_23693);
nor U24325 (N_24325,N_23665,N_22534);
or U24326 (N_24326,N_22788,N_22136);
nand U24327 (N_24327,N_22277,N_23401);
nor U24328 (N_24328,N_23069,N_22283);
xor U24329 (N_24329,N_22372,N_22643);
xnor U24330 (N_24330,N_21802,N_22683);
xnor U24331 (N_24331,N_23928,N_22219);
or U24332 (N_24332,N_21755,N_21917);
xor U24333 (N_24333,N_22879,N_22767);
nor U24334 (N_24334,N_22184,N_21097);
nand U24335 (N_24335,N_21313,N_22724);
nand U24336 (N_24336,N_21330,N_22379);
nand U24337 (N_24337,N_21385,N_22576);
xnor U24338 (N_24338,N_21236,N_23655);
xor U24339 (N_24339,N_23239,N_22268);
and U24340 (N_24340,N_22131,N_21613);
or U24341 (N_24341,N_22759,N_22382);
nand U24342 (N_24342,N_22874,N_23176);
and U24343 (N_24343,N_22820,N_21963);
xnor U24344 (N_24344,N_21939,N_22940);
nand U24345 (N_24345,N_21351,N_23947);
or U24346 (N_24346,N_23373,N_21620);
nand U24347 (N_24347,N_22481,N_22063);
and U24348 (N_24348,N_21751,N_22550);
or U24349 (N_24349,N_21594,N_22728);
and U24350 (N_24350,N_22688,N_23011);
xnor U24351 (N_24351,N_21394,N_23226);
nand U24352 (N_24352,N_22312,N_22050);
nand U24353 (N_24353,N_21431,N_22734);
xnor U24354 (N_24354,N_21793,N_21866);
or U24355 (N_24355,N_21501,N_21362);
and U24356 (N_24356,N_23630,N_23074);
and U24357 (N_24357,N_21151,N_22108);
xor U24358 (N_24358,N_23006,N_21436);
or U24359 (N_24359,N_22439,N_21285);
nor U24360 (N_24360,N_22537,N_23489);
or U24361 (N_24361,N_22914,N_21146);
xnor U24362 (N_24362,N_21031,N_21926);
and U24363 (N_24363,N_23263,N_21156);
nand U24364 (N_24364,N_23227,N_23112);
nor U24365 (N_24365,N_21509,N_21167);
nand U24366 (N_24366,N_21293,N_22568);
nor U24367 (N_24367,N_22918,N_23312);
nor U24368 (N_24368,N_23664,N_21810);
xnor U24369 (N_24369,N_23405,N_21527);
xnor U24370 (N_24370,N_21690,N_22069);
nand U24371 (N_24371,N_21722,N_22562);
or U24372 (N_24372,N_23953,N_23608);
nand U24373 (N_24373,N_23854,N_21847);
or U24374 (N_24374,N_22510,N_22873);
xnor U24375 (N_24375,N_22851,N_23571);
nor U24376 (N_24376,N_22582,N_23769);
and U24377 (N_24377,N_23950,N_22961);
nor U24378 (N_24378,N_21906,N_23715);
or U24379 (N_24379,N_22154,N_23804);
nand U24380 (N_24380,N_22429,N_22939);
xor U24381 (N_24381,N_23305,N_23990);
and U24382 (N_24382,N_22700,N_22006);
and U24383 (N_24383,N_23159,N_23235);
nor U24384 (N_24384,N_21872,N_22783);
and U24385 (N_24385,N_22616,N_23274);
and U24386 (N_24386,N_22906,N_23750);
xor U24387 (N_24387,N_21249,N_22546);
nor U24388 (N_24388,N_23836,N_23064);
or U24389 (N_24389,N_22052,N_22698);
nand U24390 (N_24390,N_21006,N_23470);
nand U24391 (N_24391,N_23206,N_23898);
nand U24392 (N_24392,N_22269,N_22169);
or U24393 (N_24393,N_22770,N_21676);
and U24394 (N_24394,N_21486,N_22886);
and U24395 (N_24395,N_21366,N_21100);
and U24396 (N_24396,N_22969,N_21514);
nand U24397 (N_24397,N_22332,N_23921);
nor U24398 (N_24398,N_21173,N_22468);
xor U24399 (N_24399,N_21563,N_23701);
xnor U24400 (N_24400,N_22040,N_23170);
xnor U24401 (N_24401,N_21943,N_23499);
nor U24402 (N_24402,N_21975,N_22509);
nand U24403 (N_24403,N_22156,N_23775);
xnor U24404 (N_24404,N_21731,N_22442);
nand U24405 (N_24405,N_21371,N_22930);
and U24406 (N_24406,N_23043,N_21094);
and U24407 (N_24407,N_21550,N_21666);
nor U24408 (N_24408,N_22690,N_21500);
and U24409 (N_24409,N_23376,N_21133);
xnor U24410 (N_24410,N_21618,N_21193);
nand U24411 (N_24411,N_23684,N_21459);
nand U24412 (N_24412,N_23207,N_22721);
nor U24413 (N_24413,N_22671,N_23397);
or U24414 (N_24414,N_22780,N_22469);
and U24415 (N_24415,N_22165,N_21662);
and U24416 (N_24416,N_22929,N_21029);
nand U24417 (N_24417,N_22822,N_21155);
nand U24418 (N_24418,N_21945,N_21554);
nor U24419 (N_24419,N_23683,N_21141);
nand U24420 (N_24420,N_22478,N_21427);
xnor U24421 (N_24421,N_22061,N_21132);
nor U24422 (N_24422,N_22755,N_22937);
or U24423 (N_24423,N_22002,N_21012);
xnor U24424 (N_24424,N_21196,N_23197);
or U24425 (N_24425,N_23155,N_22485);
xor U24426 (N_24426,N_23412,N_23918);
xor U24427 (N_24427,N_23157,N_23856);
xor U24428 (N_24428,N_21508,N_21308);
xnor U24429 (N_24429,N_23618,N_22443);
nor U24430 (N_24430,N_21875,N_23150);
or U24431 (N_24431,N_21406,N_21817);
nor U24432 (N_24432,N_23165,N_22857);
xor U24433 (N_24433,N_22102,N_23223);
or U24434 (N_24434,N_21174,N_22458);
nor U24435 (N_24435,N_23539,N_23338);
or U24436 (N_24436,N_21986,N_22908);
or U24437 (N_24437,N_22991,N_23810);
nor U24438 (N_24438,N_22207,N_21355);
nand U24439 (N_24439,N_22224,N_23559);
xor U24440 (N_24440,N_23492,N_22548);
and U24441 (N_24441,N_21255,N_23288);
xnor U24442 (N_24442,N_23761,N_23026);
and U24443 (N_24443,N_23118,N_21791);
and U24444 (N_24444,N_23361,N_22146);
or U24445 (N_24445,N_22999,N_21199);
and U24446 (N_24446,N_22593,N_23393);
and U24447 (N_24447,N_21804,N_21659);
nor U24448 (N_24448,N_21882,N_22460);
nor U24449 (N_24449,N_22495,N_22369);
nor U24450 (N_24450,N_21068,N_21727);
nor U24451 (N_24451,N_23268,N_21663);
and U24452 (N_24452,N_23824,N_22975);
nor U24453 (N_24453,N_21568,N_21334);
xor U24454 (N_24454,N_23336,N_22714);
nor U24455 (N_24455,N_23031,N_21770);
or U24456 (N_24456,N_23327,N_21224);
or U24457 (N_24457,N_23531,N_22608);
nor U24458 (N_24458,N_22685,N_23705);
and U24459 (N_24459,N_22265,N_21948);
and U24460 (N_24460,N_23020,N_22118);
or U24461 (N_24461,N_22841,N_21402);
or U24462 (N_24462,N_23348,N_22633);
xnor U24463 (N_24463,N_23175,N_22794);
and U24464 (N_24464,N_21548,N_22846);
nor U24465 (N_24465,N_21277,N_22208);
and U24466 (N_24466,N_23383,N_21887);
nand U24467 (N_24467,N_21748,N_21998);
nor U24468 (N_24468,N_21841,N_23232);
and U24469 (N_24469,N_21407,N_23437);
nor U24470 (N_24470,N_22174,N_23319);
or U24471 (N_24471,N_23504,N_21318);
and U24472 (N_24472,N_21981,N_22810);
nand U24473 (N_24473,N_23700,N_21735);
or U24474 (N_24474,N_21113,N_22217);
and U24475 (N_24475,N_22664,N_22575);
nor U24476 (N_24476,N_22113,N_21596);
or U24477 (N_24477,N_22946,N_23834);
and U24478 (N_24478,N_23760,N_22915);
nand U24479 (N_24479,N_22368,N_22526);
or U24480 (N_24480,N_22084,N_23469);
and U24481 (N_24481,N_22266,N_23983);
or U24482 (N_24482,N_22124,N_22686);
xor U24483 (N_24483,N_21016,N_23742);
or U24484 (N_24484,N_22871,N_22579);
or U24485 (N_24485,N_21163,N_22804);
nand U24486 (N_24486,N_23181,N_21304);
xnor U24487 (N_24487,N_22095,N_23975);
xnor U24488 (N_24488,N_22761,N_23436);
nor U24489 (N_24489,N_22875,N_23844);
nand U24490 (N_24490,N_23281,N_22586);
or U24491 (N_24491,N_21488,N_22927);
and U24492 (N_24492,N_21213,N_21434);
and U24493 (N_24493,N_22881,N_23056);
or U24494 (N_24494,N_21516,N_21138);
xnor U24495 (N_24495,N_22631,N_23343);
and U24496 (N_24496,N_22978,N_21679);
xnor U24497 (N_24497,N_21036,N_22974);
nand U24498 (N_24498,N_23895,N_21248);
nand U24499 (N_24499,N_22916,N_23574);
nand U24500 (N_24500,N_22427,N_23986);
nor U24501 (N_24501,N_23260,N_23935);
nor U24502 (N_24502,N_21698,N_23113);
nor U24503 (N_24503,N_22298,N_23023);
nand U24504 (N_24504,N_21740,N_22707);
nor U24505 (N_24505,N_22405,N_21372);
and U24506 (N_24506,N_22956,N_22281);
or U24507 (N_24507,N_22791,N_23675);
and U24508 (N_24508,N_22194,N_22413);
nor U24509 (N_24509,N_23218,N_21095);
nand U24510 (N_24510,N_22876,N_21686);
or U24511 (N_24511,N_22275,N_21587);
nor U24512 (N_24512,N_23586,N_22492);
and U24513 (N_24513,N_21021,N_23924);
nor U24514 (N_24514,N_21993,N_22727);
and U24515 (N_24515,N_22128,N_22012);
or U24516 (N_24516,N_22255,N_22706);
xnor U24517 (N_24517,N_22171,N_23507);
nor U24518 (N_24518,N_22091,N_23065);
or U24519 (N_24519,N_22338,N_23423);
nor U24520 (N_24520,N_23694,N_21433);
nor U24521 (N_24521,N_22234,N_22292);
nand U24522 (N_24522,N_23483,N_21622);
and U24523 (N_24523,N_21328,N_23264);
xnor U24524 (N_24524,N_22057,N_22895);
nor U24525 (N_24525,N_21261,N_22869);
xor U24526 (N_24526,N_22339,N_21298);
nand U24527 (N_24527,N_21991,N_22370);
nand U24528 (N_24528,N_21603,N_23440);
xnor U24529 (N_24529,N_22003,N_21794);
and U24530 (N_24530,N_23354,N_23794);
xnor U24531 (N_24531,N_21111,N_23782);
and U24532 (N_24532,N_23448,N_23151);
nor U24533 (N_24533,N_21278,N_21680);
or U24534 (N_24534,N_22722,N_22000);
and U24535 (N_24535,N_22667,N_23257);
nor U24536 (N_24536,N_23960,N_22758);
or U24537 (N_24537,N_23583,N_22607);
xor U24538 (N_24538,N_21736,N_23793);
and U24539 (N_24539,N_22723,N_23916);
nor U24540 (N_24540,N_21273,N_21564);
and U24541 (N_24541,N_23600,N_22264);
nor U24542 (N_24542,N_23353,N_23303);
and U24543 (N_24543,N_23735,N_21897);
nor U24544 (N_24544,N_22725,N_23852);
or U24545 (N_24545,N_23177,N_21705);
nand U24546 (N_24546,N_23903,N_21284);
nand U24547 (N_24547,N_23106,N_21557);
xor U24548 (N_24548,N_23472,N_23196);
and U24549 (N_24549,N_23005,N_21633);
nand U24550 (N_24550,N_23429,N_21860);
and U24551 (N_24551,N_23451,N_21222);
and U24552 (N_24552,N_23878,N_21921);
nor U24553 (N_24553,N_22404,N_21024);
and U24554 (N_24554,N_21837,N_22347);
xnor U24555 (N_24555,N_22987,N_21073);
nor U24556 (N_24556,N_21977,N_23306);
and U24557 (N_24557,N_23753,N_23096);
nand U24558 (N_24558,N_22231,N_23661);
or U24559 (N_24559,N_23768,N_22856);
and U24560 (N_24560,N_21119,N_21503);
nand U24561 (N_24561,N_21592,N_21390);
nor U24562 (N_24562,N_23039,N_21039);
xor U24563 (N_24563,N_22425,N_22477);
nand U24564 (N_24564,N_21154,N_23058);
nor U24565 (N_24565,N_21083,N_21469);
or U24566 (N_24566,N_22009,N_23503);
nand U24567 (N_24567,N_22744,N_22920);
nand U24568 (N_24568,N_22891,N_21159);
nand U24569 (N_24569,N_21760,N_21387);
nand U24570 (N_24570,N_21368,N_21670);
nand U24571 (N_24571,N_23358,N_22765);
and U24572 (N_24572,N_23077,N_23766);
xnor U24573 (N_24573,N_22319,N_22549);
nor U24574 (N_24574,N_22609,N_22190);
or U24575 (N_24575,N_21531,N_23091);
nand U24576 (N_24576,N_22449,N_21905);
nand U24577 (N_24577,N_22383,N_21397);
and U24578 (N_24578,N_21093,N_23917);
nor U24579 (N_24579,N_21924,N_23216);
or U24580 (N_24580,N_22973,N_21225);
or U24581 (N_24581,N_22612,N_23184);
nor U24582 (N_24582,N_21189,N_23289);
nor U24583 (N_24583,N_22792,N_22204);
or U24584 (N_24584,N_23454,N_22943);
nor U24585 (N_24585,N_22530,N_22807);
nand U24586 (N_24586,N_21315,N_22619);
nand U24587 (N_24587,N_23476,N_22574);
nor U24588 (N_24588,N_21043,N_22996);
and U24589 (N_24589,N_23482,N_21615);
and U24590 (N_24590,N_23723,N_23459);
nor U24591 (N_24591,N_21042,N_22293);
or U24592 (N_24592,N_22699,N_23341);
or U24593 (N_24593,N_21474,N_23416);
and U24594 (N_24594,N_22280,N_22893);
and U24595 (N_24595,N_23363,N_22680);
or U24596 (N_24596,N_21800,N_23617);
nor U24597 (N_24597,N_21691,N_21451);
nand U24598 (N_24598,N_23038,N_22349);
nand U24599 (N_24599,N_22597,N_22779);
nor U24600 (N_24600,N_22122,N_23490);
or U24601 (N_24601,N_22625,N_21358);
xnor U24602 (N_24602,N_22566,N_22678);
xnor U24603 (N_24603,N_21109,N_23413);
or U24604 (N_24604,N_22516,N_23183);
nand U24605 (N_24605,N_23578,N_21653);
nand U24606 (N_24606,N_21953,N_23905);
or U24607 (N_24607,N_22450,N_21070);
nand U24608 (N_24608,N_21694,N_22085);
nand U24609 (N_24609,N_21829,N_21171);
nor U24610 (N_24610,N_21797,N_23262);
or U24611 (N_24611,N_21033,N_22814);
and U24612 (N_24612,N_23639,N_23959);
and U24613 (N_24613,N_23246,N_21259);
and U24614 (N_24614,N_23547,N_22259);
xnor U24615 (N_24615,N_23291,N_23812);
nand U24616 (N_24616,N_22653,N_23080);
xnor U24617 (N_24617,N_23979,N_22733);
or U24618 (N_24618,N_23648,N_21729);
nor U24619 (N_24619,N_23602,N_21709);
nand U24620 (N_24620,N_21169,N_21657);
and U24621 (N_24621,N_23251,N_22330);
and U24622 (N_24622,N_21245,N_22074);
and U24623 (N_24623,N_21923,N_23452);
and U24624 (N_24624,N_22378,N_23597);
and U24625 (N_24625,N_23075,N_22494);
xnor U24626 (N_24626,N_23282,N_23072);
nor U24627 (N_24627,N_23713,N_21025);
and U24628 (N_24628,N_21437,N_21347);
and U24629 (N_24629,N_23550,N_23463);
xor U24630 (N_24630,N_21764,N_22150);
nand U24631 (N_24631,N_23962,N_23998);
or U24632 (N_24632,N_22452,N_22793);
or U24633 (N_24633,N_21307,N_21370);
or U24634 (N_24634,N_21336,N_21692);
nor U24635 (N_24635,N_21099,N_23832);
and U24636 (N_24636,N_23853,N_23984);
nand U24637 (N_24637,N_22261,N_23299);
nor U24638 (N_24638,N_23356,N_23876);
and U24639 (N_24639,N_21995,N_22029);
xor U24640 (N_24640,N_22416,N_23816);
xor U24641 (N_24641,N_21238,N_22112);
xor U24642 (N_24642,N_22529,N_22663);
or U24643 (N_24643,N_22027,N_23225);
nor U24644 (N_24644,N_21223,N_22971);
nand U24645 (N_24645,N_21718,N_22601);
xnor U24646 (N_24646,N_23879,N_23431);
nor U24647 (N_24647,N_22965,N_21685);
xor U24648 (N_24648,N_21200,N_23002);
or U24649 (N_24649,N_22145,N_23666);
nor U24650 (N_24650,N_21369,N_21957);
or U24651 (N_24651,N_21244,N_22245);
and U24652 (N_24652,N_23530,N_23494);
or U24653 (N_24653,N_22913,N_21616);
nand U24654 (N_24654,N_21379,N_23051);
nor U24655 (N_24655,N_23022,N_22191);
xnor U24656 (N_24656,N_21374,N_22754);
or U24657 (N_24657,N_22583,N_21135);
xnor U24658 (N_24658,N_23897,N_21365);
xor U24659 (N_24659,N_23755,N_21712);
and U24660 (N_24660,N_22045,N_22644);
or U24661 (N_24661,N_21888,N_23277);
nand U24662 (N_24662,N_22497,N_23193);
nor U24663 (N_24663,N_21654,N_21849);
nand U24664 (N_24664,N_23414,N_23479);
nand U24665 (N_24665,N_21157,N_21462);
nand U24666 (N_24666,N_22953,N_23860);
and U24667 (N_24667,N_22251,N_21702);
or U24668 (N_24668,N_22086,N_23946);
nor U24669 (N_24669,N_23667,N_23778);
xor U24670 (N_24670,N_23743,N_23579);
nand U24671 (N_24671,N_23127,N_21000);
nand U24672 (N_24672,N_23739,N_21706);
or U24673 (N_24673,N_21438,N_22921);
or U24674 (N_24674,N_21664,N_23620);
xor U24675 (N_24675,N_23047,N_22203);
or U24676 (N_24676,N_22105,N_23370);
xor U24677 (N_24677,N_21009,N_23893);
nor U24678 (N_24678,N_23078,N_22995);
and U24679 (N_24679,N_23601,N_22803);
xnor U24680 (N_24680,N_21966,N_22001);
nor U24681 (N_24681,N_21625,N_23546);
nand U24682 (N_24682,N_23567,N_23716);
and U24683 (N_24683,N_21851,N_23142);
or U24684 (N_24684,N_23194,N_23162);
nor U24685 (N_24685,N_22401,N_22420);
nand U24686 (N_24686,N_23433,N_22580);
nand U24687 (N_24687,N_22042,N_22314);
and U24688 (N_24688,N_23889,N_21274);
nand U24689 (N_24689,N_23736,N_23869);
nand U24690 (N_24690,N_21919,N_21449);
and U24691 (N_24691,N_22676,N_23071);
nand U24692 (N_24692,N_22013,N_22799);
and U24693 (N_24693,N_22243,N_23455);
nor U24694 (N_24694,N_23993,N_21086);
nand U24695 (N_24695,N_23565,N_21823);
nor U24696 (N_24696,N_22185,N_23017);
nand U24697 (N_24697,N_21357,N_23372);
nor U24698 (N_24698,N_21074,N_22361);
nand U24699 (N_24699,N_23367,N_21581);
nand U24700 (N_24700,N_23344,N_22944);
xor U24701 (N_24701,N_22589,N_23553);
nor U24702 (N_24702,N_22073,N_21836);
nor U24703 (N_24703,N_21842,N_23721);
and U24704 (N_24704,N_21775,N_22423);
or U24705 (N_24705,N_22697,N_22130);
xor U24706 (N_24706,N_21920,N_21960);
xor U24707 (N_24707,N_23202,N_23958);
xnor U24708 (N_24708,N_22192,N_22390);
and U24709 (N_24709,N_21969,N_23790);
and U24710 (N_24710,N_23858,N_23500);
and U24711 (N_24711,N_23532,N_23681);
nor U24712 (N_24712,N_23114,N_23606);
or U24713 (N_24713,N_23229,N_23866);
nor U24714 (N_24714,N_22163,N_21114);
and U24715 (N_24715,N_22571,N_23857);
or U24716 (N_24716,N_23609,N_23942);
and U24717 (N_24717,N_21124,N_21312);
or U24718 (N_24718,N_22022,N_22637);
or U24719 (N_24719,N_21058,N_22044);
or U24720 (N_24720,N_21941,N_21144);
nor U24721 (N_24721,N_23076,N_22092);
nand U24722 (N_24722,N_23390,N_22997);
nor U24723 (N_24723,N_23188,N_22408);
xor U24724 (N_24724,N_23863,N_21301);
xor U24725 (N_24725,N_23938,N_23487);
xnor U24726 (N_24726,N_21547,N_23948);
xor U24727 (N_24727,N_23633,N_21342);
nand U24728 (N_24728,N_21404,N_21066);
and U24729 (N_24729,N_23980,N_23829);
and U24730 (N_24730,N_21340,N_23209);
and U24731 (N_24731,N_21098,N_23838);
or U24732 (N_24732,N_22162,N_23972);
or U24733 (N_24733,N_23329,N_21322);
or U24734 (N_24734,N_23137,N_23110);
xnor U24735 (N_24735,N_21158,N_21854);
xnor U24736 (N_24736,N_23732,N_23594);
nor U24737 (N_24737,N_21417,N_22396);
nand U24738 (N_24738,N_21595,N_23402);
xnor U24739 (N_24739,N_22228,N_21946);
xor U24740 (N_24740,N_22419,N_21602);
or U24741 (N_24741,N_22551,N_22407);
or U24742 (N_24742,N_21037,N_22149);
nand U24743 (N_24743,N_22958,N_22461);
nand U24744 (N_24744,N_21938,N_23126);
nand U24745 (N_24745,N_21903,N_21813);
and U24746 (N_24746,N_22813,N_23690);
and U24747 (N_24747,N_23851,N_22071);
or U24748 (N_24748,N_22936,N_21034);
or U24749 (N_24749,N_21446,N_21750);
nand U24750 (N_24750,N_23779,N_23754);
xnor U24751 (N_24751,N_23018,N_22087);
xor U24752 (N_24752,N_21044,N_21305);
nand U24753 (N_24753,N_22638,N_22888);
and U24754 (N_24754,N_21183,N_21345);
and U24755 (N_24755,N_22954,N_21482);
nor U24756 (N_24756,N_22641,N_23556);
nor U24757 (N_24757,N_23148,N_21348);
xor U24758 (N_24758,N_23951,N_21517);
and U24759 (N_24759,N_21696,N_21164);
nand U24760 (N_24760,N_23662,N_23185);
and U24761 (N_24761,N_22167,N_21206);
nor U24762 (N_24762,N_23849,N_22229);
and U24763 (N_24763,N_23398,N_23371);
nand U24764 (N_24764,N_22499,N_23672);
xnor U24765 (N_24765,N_21004,N_21415);
and U24766 (N_24766,N_22866,N_22842);
nor U24767 (N_24767,N_22624,N_23278);
nand U24768 (N_24768,N_21868,N_23250);
or U24769 (N_24769,N_21789,N_23668);
xor U24770 (N_24770,N_22819,N_21746);
and U24771 (N_24771,N_22668,N_23286);
or U24772 (N_24772,N_23636,N_23989);
and U24773 (N_24773,N_23848,N_21782);
nor U24774 (N_24774,N_23797,N_22082);
nand U24775 (N_24775,N_22812,N_22035);
nor U24776 (N_24776,N_22718,N_21881);
xor U24777 (N_24777,N_23255,N_21424);
and U24778 (N_24778,N_22868,N_22426);
nor U24779 (N_24779,N_21090,N_22410);
nor U24780 (N_24780,N_21695,N_22227);
nor U24781 (N_24781,N_21936,N_23973);
nor U24782 (N_24782,N_22271,N_21771);
nand U24783 (N_24783,N_23377,N_22137);
nor U24784 (N_24784,N_21541,N_22865);
xor U24785 (N_24785,N_21935,N_22646);
and U24786 (N_24786,N_21493,N_22640);
xnor U24787 (N_24787,N_21983,N_23638);
and U24788 (N_24788,N_22890,N_21333);
nand U24789 (N_24789,N_23526,N_21460);
xor U24790 (N_24790,N_22041,N_22299);
nand U24791 (N_24791,N_22053,N_21018);
nor U24792 (N_24792,N_22861,N_21041);
nand U24793 (N_24793,N_23087,N_22621);
xnor U24794 (N_24794,N_23727,N_23906);
and U24795 (N_24795,N_21911,N_21013);
nand U24796 (N_24796,N_21844,N_22360);
nor U24797 (N_24797,N_22409,N_21915);
xor U24798 (N_24798,N_23201,N_21990);
or U24799 (N_24799,N_22847,N_23819);
and U24800 (N_24800,N_21521,N_23495);
and U24801 (N_24801,N_23267,N_23615);
nand U24802 (N_24802,N_21677,N_23136);
nor U24803 (N_24803,N_22358,N_23070);
or U24804 (N_24804,N_23439,N_23674);
nor U24805 (N_24805,N_23213,N_21682);
nor U24806 (N_24806,N_22036,N_23649);
and U24807 (N_24807,N_21658,N_23204);
nor U24808 (N_24808,N_23399,N_21555);
or U24809 (N_24809,N_22431,N_21971);
nand U24810 (N_24810,N_23249,N_21152);
or U24811 (N_24811,N_21848,N_23190);
nand U24812 (N_24812,N_21354,N_22691);
nand U24813 (N_24813,N_23450,N_22742);
nor U24814 (N_24814,N_22766,N_23722);
or U24815 (N_24815,N_21480,N_22864);
nor U24816 (N_24816,N_23109,N_21022);
xnor U24817 (N_24817,N_22594,N_23473);
or U24818 (N_24818,N_22557,N_21934);
nor U24819 (N_24819,N_22737,N_23896);
or U24820 (N_24820,N_22967,N_22605);
nand U24821 (N_24821,N_22862,N_22828);
nor U24822 (N_24822,N_23841,N_22309);
nand U24823 (N_24823,N_23107,N_22371);
and U24824 (N_24824,N_21715,N_23425);
and U24825 (N_24825,N_21356,N_21651);
xnor U24826 (N_24826,N_21085,N_21232);
xnor U24827 (N_24827,N_22422,N_22615);
or U24828 (N_24828,N_23659,N_22139);
nor U24829 (N_24829,N_22289,N_22062);
or U24830 (N_24830,N_21687,N_22385);
or U24831 (N_24831,N_21944,N_23421);
nand U24832 (N_24832,N_22626,N_22183);
and U24833 (N_24833,N_23640,N_21053);
xnor U24834 (N_24834,N_21092,N_22301);
and U24835 (N_24835,N_23147,N_21343);
xor U24836 (N_24836,N_21263,N_21968);
or U24837 (N_24837,N_22902,N_23221);
and U24838 (N_24838,N_21444,N_21769);
xnor U24839 (N_24839,N_22489,N_23555);
xor U24840 (N_24840,N_21015,N_22463);
or U24841 (N_24841,N_21982,N_22179);
nand U24842 (N_24842,N_21704,N_21339);
or U24843 (N_24843,N_21510,N_23141);
and U24844 (N_24844,N_21108,N_22451);
nor U24845 (N_24845,N_23276,N_21850);
and U24846 (N_24846,N_22197,N_23999);
nor U24847 (N_24847,N_23825,N_22768);
and U24848 (N_24848,N_22010,N_23787);
nor U24849 (N_24849,N_22188,N_23710);
xor U24850 (N_24850,N_23468,N_21272);
xor U24851 (N_24851,N_23186,N_22239);
and U24852 (N_24852,N_22388,N_22525);
xnor U24853 (N_24853,N_22634,N_22565);
or U24854 (N_24854,N_21186,N_23708);
nor U24855 (N_24855,N_23882,N_23516);
nand U24856 (N_24856,N_21795,N_21380);
or U24857 (N_24857,N_22135,N_22863);
and U24858 (N_24858,N_21752,N_23971);
nor U24859 (N_24859,N_21267,N_22273);
nor U24860 (N_24860,N_22655,N_21048);
or U24861 (N_24861,N_22983,N_21217);
nor U24862 (N_24862,N_22786,N_21839);
xnor U24863 (N_24863,N_23456,N_22161);
nand U24864 (N_24864,N_23611,N_22506);
and U24865 (N_24865,N_22661,N_21051);
nor U24866 (N_24866,N_22465,N_22376);
and U24867 (N_24867,N_23941,N_23899);
or U24868 (N_24868,N_23134,N_22453);
nor U24869 (N_24869,N_21471,N_22448);
xor U24870 (N_24870,N_21299,N_23156);
nand U24871 (N_24871,N_22556,N_21552);
nand U24872 (N_24872,N_22215,N_22998);
or U24873 (N_24873,N_23551,N_23140);
xnor U24874 (N_24874,N_22196,N_23032);
nand U24875 (N_24875,N_23776,N_21096);
xnor U24876 (N_24876,N_23909,N_22693);
and U24877 (N_24877,N_23007,N_21463);
xnor U24878 (N_24878,N_21023,N_23785);
xor U24879 (N_24879,N_22606,N_21644);
xnor U24880 (N_24880,N_23205,N_22250);
or U24881 (N_24881,N_22642,N_21627);
nand U24882 (N_24882,N_23926,N_21538);
or U24883 (N_24883,N_22295,N_22096);
nor U24884 (N_24884,N_21061,N_22858);
nor U24885 (N_24885,N_23612,N_23406);
and U24886 (N_24886,N_22026,N_22286);
xor U24887 (N_24887,N_23486,N_23695);
and U24888 (N_24888,N_21269,N_22101);
nand U24889 (N_24889,N_23877,N_23258);
xor U24890 (N_24890,N_23474,N_22235);
and U24891 (N_24891,N_21112,N_23380);
or U24892 (N_24892,N_23447,N_23292);
or U24893 (N_24893,N_23835,N_23534);
xnor U24894 (N_24894,N_21984,N_23290);
or U24895 (N_24895,N_22839,N_23525);
nor U24896 (N_24896,N_21478,N_23021);
xor U24897 (N_24897,N_23581,N_21589);
or U24898 (N_24898,N_21254,N_21913);
nand U24899 (N_24899,N_21745,N_22140);
and U24900 (N_24900,N_23932,N_22836);
nor U24901 (N_24901,N_21522,N_21028);
xnor U24902 (N_24902,N_21967,N_23524);
nand U24903 (N_24903,N_21453,N_23308);
nor U24904 (N_24904,N_22263,N_23933);
or U24905 (N_24905,N_21204,N_23426);
nor U24906 (N_24906,N_23566,N_23294);
nand U24907 (N_24907,N_21219,N_23757);
and U24908 (N_24908,N_23480,N_23593);
and U24909 (N_24909,N_22032,N_22692);
or U24910 (N_24910,N_22432,N_21220);
and U24911 (N_24911,N_21586,N_23283);
and U24912 (N_24912,N_23060,N_21341);
or U24913 (N_24913,N_22505,N_22713);
and U24914 (N_24914,N_23224,N_23762);
nand U24915 (N_24915,N_23923,N_22249);
nand U24916 (N_24916,N_23536,N_21118);
or U24917 (N_24917,N_21907,N_23315);
nand U24918 (N_24918,N_23900,N_23345);
xnor U24919 (N_24919,N_22942,N_22797);
or U24920 (N_24920,N_22848,N_23297);
or U24921 (N_24921,N_22610,N_22838);
or U24922 (N_24922,N_23987,N_21803);
nand U24923 (N_24923,N_22374,N_22152);
nor U24924 (N_24924,N_23219,N_22411);
or U24925 (N_24925,N_22620,N_22753);
xor U24926 (N_24926,N_22892,N_22884);
or U24927 (N_24927,N_21102,N_21405);
nand U24928 (N_24928,N_21930,N_22386);
nand U24929 (N_24929,N_22049,N_23019);
nand U24930 (N_24930,N_23982,N_23384);
or U24931 (N_24931,N_22362,N_21054);
xor U24932 (N_24932,N_21026,N_22346);
nand U24933 (N_24933,N_22923,N_23859);
or U24934 (N_24934,N_23756,N_21282);
nand U24935 (N_24935,N_23520,N_22950);
or U24936 (N_24936,N_22694,N_23955);
nand U24937 (N_24937,N_21306,N_21884);
nor U24938 (N_24938,N_22673,N_21425);
nand U24939 (N_24939,N_21645,N_23172);
and U24940 (N_24940,N_21190,N_23138);
nand U24941 (N_24941,N_23543,N_21378);
nand U24942 (N_24942,N_21593,N_23168);
xnor U24943 (N_24943,N_23913,N_22392);
nand U24944 (N_24944,N_21454,N_22670);
xnor U24945 (N_24945,N_21525,N_23576);
or U24946 (N_24946,N_22393,N_23418);
nand U24947 (N_24947,N_21588,N_21107);
nor U24948 (N_24948,N_22553,N_22531);
nor U24949 (N_24949,N_22784,N_21143);
and U24950 (N_24950,N_23919,N_22764);
xnor U24951 (N_24951,N_23350,N_23247);
nor U24952 (N_24952,N_21741,N_21940);
and U24953 (N_24953,N_21822,N_23845);
or U24954 (N_24954,N_21242,N_22177);
xnor U24955 (N_24955,N_22547,N_23231);
nor U24956 (N_24956,N_21001,N_21626);
or U24957 (N_24957,N_22980,N_22802);
xnor U24958 (N_24958,N_23865,N_23697);
or U24959 (N_24959,N_21038,N_22189);
xnor U24960 (N_24960,N_21916,N_22375);
xor U24961 (N_24961,N_23806,N_22187);
nor U24962 (N_24962,N_22487,N_22220);
or U24963 (N_24963,N_21128,N_23968);
and U24964 (N_24964,N_21129,N_21229);
xor U24965 (N_24965,N_23645,N_21198);
and U24966 (N_24966,N_23240,N_23974);
nand U24967 (N_24967,N_23904,N_22125);
nand U24968 (N_24968,N_23419,N_21765);
nor U24969 (N_24969,N_23042,N_22618);
nor U24970 (N_24970,N_23385,N_21497);
and U24971 (N_24971,N_21918,N_23800);
or U24972 (N_24972,N_23057,N_23287);
nand U24973 (N_24973,N_22745,N_22949);
or U24974 (N_24974,N_21005,N_23915);
xnor U24975 (N_24975,N_23061,N_22127);
or U24976 (N_24976,N_23588,N_21855);
and U24977 (N_24977,N_22336,N_22925);
xor U24978 (N_24978,N_22748,N_23698);
xor U24979 (N_24979,N_21951,N_23272);
or U24980 (N_24980,N_22325,N_21843);
or U24981 (N_24981,N_21819,N_21668);
nand U24982 (N_24982,N_21414,N_21439);
xor U24983 (N_24983,N_23940,N_22004);
or U24984 (N_24984,N_21830,N_23541);
nor U24985 (N_24985,N_21724,N_22195);
or U24986 (N_24986,N_23475,N_21647);
nor U24987 (N_24987,N_21728,N_23544);
or U24988 (N_24988,N_23364,N_21472);
nor U24989 (N_24989,N_22926,N_21253);
xnor U24990 (N_24990,N_22989,N_23008);
or U24991 (N_24991,N_22352,N_21566);
nand U24992 (N_24992,N_22028,N_23296);
xor U24993 (N_24993,N_23518,N_23323);
and U24994 (N_24994,N_22703,N_23931);
and U24995 (N_24995,N_22366,N_22705);
and U24996 (N_24996,N_23994,N_21959);
xor U24997 (N_24997,N_22232,N_21076);
nand U24998 (N_24998,N_23488,N_21688);
and U24999 (N_24999,N_21762,N_23545);
or U25000 (N_25000,N_21237,N_22896);
xor U25001 (N_25001,N_23658,N_21807);
nand U25002 (N_25002,N_23641,N_21597);
or U25003 (N_25003,N_22901,N_21327);
nor U25004 (N_25004,N_21182,N_23772);
or U25005 (N_25005,N_21288,N_22075);
xor U25006 (N_25006,N_21733,N_23605);
xor U25007 (N_25007,N_21291,N_23868);
or U25008 (N_25008,N_23265,N_22039);
nor U25009 (N_25009,N_21989,N_22484);
nand U25010 (N_25010,N_21996,N_22993);
nand U25011 (N_25011,N_22335,N_22513);
nor U25012 (N_25012,N_21377,N_21980);
nand U25013 (N_25013,N_22341,N_22808);
xor U25014 (N_25014,N_22992,N_21726);
or U25015 (N_25015,N_21773,N_22479);
nor U25016 (N_25016,N_22018,N_22406);
xor U25017 (N_25017,N_21294,N_21565);
or U25018 (N_25018,N_21544,N_21147);
nand U25019 (N_25019,N_22132,N_22829);
xor U25020 (N_25020,N_22072,N_22318);
and U25021 (N_25021,N_22732,N_23506);
nand U25022 (N_25022,N_21050,N_23352);
nor U25023 (N_25023,N_22193,N_23320);
nor U25024 (N_25024,N_23430,N_21495);
xnor U25025 (N_25025,N_23189,N_22776);
xnor U25026 (N_25026,N_22175,N_21631);
nand U25027 (N_25027,N_21796,N_23200);
or U25028 (N_25028,N_22749,N_21831);
nand U25029 (N_25029,N_21421,N_22774);
nor U25030 (N_25030,N_21475,N_21759);
xnor U25031 (N_25031,N_23084,N_23587);
and U25032 (N_25032,N_23558,N_23164);
xor U25033 (N_25033,N_22985,N_23604);
or U25034 (N_25034,N_21409,N_23163);
nand U25035 (N_25035,N_21300,N_23519);
and U25036 (N_25036,N_23059,N_22260);
nand U25037 (N_25037,N_23862,N_22144);
nor U25038 (N_25038,N_22932,N_21105);
or U25039 (N_25039,N_22104,N_22115);
nand U25040 (N_25040,N_22222,N_22496);
nor U25041 (N_25041,N_21410,N_23003);
nand U25042 (N_25042,N_21296,N_22782);
xor U25043 (N_25043,N_21423,N_23890);
nor U25044 (N_25044,N_21281,N_21349);
nor U25045 (N_25045,N_21649,N_22109);
nor U25046 (N_25046,N_23178,N_21331);
and U25047 (N_25047,N_21876,N_22380);
or U25048 (N_25048,N_23970,N_21873);
nand U25049 (N_25049,N_22689,N_22805);
nor U25050 (N_25050,N_23801,N_21556);
xor U25051 (N_25051,N_21671,N_22094);
nand U25052 (N_25052,N_23441,N_21958);
or U25053 (N_25053,N_21442,N_22544);
nor U25054 (N_25054,N_22253,N_21292);
xor U25055 (N_25055,N_23085,N_21513);
or U25056 (N_25056,N_23400,N_23528);
xnor U25057 (N_25057,N_21720,N_22126);
nor U25058 (N_25058,N_23788,N_22322);
and U25059 (N_25059,N_22067,N_21585);
and U25060 (N_25060,N_23822,N_21126);
and U25061 (N_25061,N_22435,N_21756);
and U25062 (N_25062,N_22297,N_23510);
or U25063 (N_25063,N_22581,N_23079);
xor U25064 (N_25064,N_21166,N_21088);
nor U25065 (N_25065,N_21352,N_22503);
and U25066 (N_25066,N_23477,N_22735);
xnor U25067 (N_25067,N_21353,N_23861);
or U25068 (N_25068,N_21725,N_21646);
or U25069 (N_25069,N_21927,N_23301);
nand U25070 (N_25070,N_22515,N_22024);
and U25071 (N_25071,N_21260,N_23686);
nor U25072 (N_25072,N_21573,N_23105);
or U25073 (N_25073,N_23737,N_22845);
xnor U25074 (N_25074,N_23000,N_22984);
nand U25075 (N_25075,N_21790,N_22859);
and U25076 (N_25076,N_21047,N_21678);
or U25077 (N_25077,N_23458,N_22342);
and U25078 (N_25078,N_21601,N_23387);
or U25079 (N_25079,N_22627,N_21045);
nand U25080 (N_25080,N_23807,N_22517);
nand U25081 (N_25081,N_21104,N_21049);
nor U25082 (N_25082,N_22731,N_22739);
nor U25083 (N_25083,N_22843,N_21137);
and U25084 (N_25084,N_23404,N_21360);
xor U25085 (N_25085,N_22348,N_21136);
nand U25086 (N_25086,N_22363,N_23741);
or U25087 (N_25087,N_23637,N_23115);
or U25088 (N_25088,N_21965,N_23464);
or U25089 (N_25089,N_21443,N_21933);
nor U25090 (N_25090,N_21684,N_21324);
or U25091 (N_25091,N_22430,N_22206);
and U25092 (N_25092,N_21999,N_21411);
xnor U25093 (N_25093,N_21250,N_23691);
xnor U25094 (N_25094,N_21673,N_21496);
or U25095 (N_25095,N_21367,N_22778);
nor U25096 (N_25096,N_22716,N_22623);
nor U25097 (N_25097,N_23692,N_21612);
nand U25098 (N_25098,N_21777,N_21252);
nor U25099 (N_25099,N_22134,N_21754);
or U25100 (N_25100,N_22762,N_22986);
or U25101 (N_25101,N_22047,N_21846);
and U25102 (N_25102,N_22826,N_22178);
nor U25103 (N_25103,N_22659,N_23378);
nand U25104 (N_25104,N_21289,N_21227);
nor U25105 (N_25105,N_22387,N_22563);
or U25106 (N_25106,N_22889,N_22414);
nand U25107 (N_25107,N_21494,N_21578);
nand U25108 (N_25108,N_23803,N_22233);
and U25109 (N_25109,N_23233,N_23335);
or U25110 (N_25110,N_23864,N_22486);
xor U25111 (N_25111,N_22291,N_21617);
nand U25112 (N_25112,N_23613,N_23709);
or U25113 (N_25113,N_21381,N_23871);
or U25114 (N_25114,N_23092,N_23408);
xnor U25115 (N_25115,N_22818,N_23333);
or U25116 (N_25116,N_22785,N_23647);
or U25117 (N_25117,N_22738,N_22394);
nand U25118 (N_25118,N_22464,N_22210);
nand U25119 (N_25119,N_22459,N_23929);
nor U25120 (N_25120,N_22437,N_22327);
nand U25121 (N_25121,N_23256,N_22353);
nand U25122 (N_25122,N_21479,N_21511);
nand U25123 (N_25123,N_22844,N_21490);
nand U25124 (N_25124,N_23214,N_23073);
nor U25125 (N_25125,N_21216,N_21418);
or U25126 (N_25126,N_21317,N_21122);
and U25127 (N_25127,N_23570,N_21979);
nand U25128 (N_25128,N_21361,N_21400);
xnor U25129 (N_25129,N_21059,N_23044);
nand U25130 (N_25130,N_21786,N_22080);
nand U25131 (N_25131,N_22064,N_21145);
and U25132 (N_25132,N_23300,N_21539);
nor U25133 (N_25133,N_21701,N_22021);
nand U25134 (N_25134,N_23403,N_22007);
nand U25135 (N_25135,N_21551,N_22559);
xor U25136 (N_25136,N_22493,N_22015);
xor U25137 (N_25137,N_23167,N_23501);
nor U25138 (N_25138,N_23883,N_22320);
nor U25139 (N_25139,N_22241,N_21290);
nand U25140 (N_25140,N_23409,N_23461);
nor U25141 (N_25141,N_22457,N_21134);
xnor U25142 (N_25142,N_21580,N_23453);
or U25143 (N_25143,N_23632,N_23052);
and U25144 (N_25144,N_21976,N_23496);
xor U25145 (N_25145,N_22500,N_22897);
or U25146 (N_25146,N_21140,N_23725);
nand U25147 (N_25147,N_21845,N_23631);
xor U25148 (N_25148,N_21925,N_21744);
xnor U25149 (N_25149,N_21303,N_21994);
and U25150 (N_25150,N_22912,N_22106);
nor U25151 (N_25151,N_22938,N_21838);
or U25152 (N_25152,N_22424,N_21914);
and U25153 (N_25153,N_22602,N_21877);
nand U25154 (N_25154,N_21075,N_21452);
nor U25155 (N_25155,N_23420,N_23562);
nand U25156 (N_25156,N_21325,N_22421);
or U25157 (N_25157,N_23719,N_23362);
and U25158 (N_25158,N_23465,N_21891);
and U25159 (N_25159,N_21422,N_23273);
nor U25160 (N_25160,N_23295,N_23867);
or U25161 (N_25161,N_22054,N_22048);
xnor U25162 (N_25162,N_23097,N_22119);
and U25163 (N_25163,N_23095,N_23266);
xor U25164 (N_25164,N_21130,N_21591);
or U25165 (N_25165,N_21210,N_23744);
xor U25166 (N_25166,N_23963,N_22709);
xor U25167 (N_25167,N_21389,N_21388);
or U25168 (N_25168,N_23523,N_23598);
and U25169 (N_25169,N_23088,N_21440);
and U25170 (N_25170,N_23212,N_22236);
xor U25171 (N_25171,N_22107,N_23512);
nor U25172 (N_25172,N_23625,N_22093);
nor U25173 (N_25173,N_23094,N_23203);
nand U25174 (N_25174,N_22473,N_23537);
and U25175 (N_25175,N_21161,N_23811);
or U25176 (N_25176,N_22290,N_21571);
nor U25177 (N_25177,N_22337,N_23751);
or U25178 (N_25178,N_23703,N_22924);
nand U25179 (N_25179,N_21825,N_23580);
nand U25180 (N_25180,N_22403,N_21456);
nand U25181 (N_25181,N_23813,N_22648);
nand U25182 (N_25182,N_22990,N_21283);
nand U25183 (N_25183,N_23388,N_21655);
nand U25184 (N_25184,N_22715,N_21115);
nand U25185 (N_25185,N_22660,N_21779);
nor U25186 (N_25186,N_22285,N_21506);
or U25187 (N_25187,N_21956,N_21445);
nand U25188 (N_25188,N_23041,N_22246);
nand U25189 (N_25189,N_22474,N_21120);
and U25190 (N_25190,N_23614,N_22116);
nand U25191 (N_25191,N_22070,N_21973);
nor U25192 (N_25192,N_21672,N_21457);
nor U25193 (N_25193,N_22904,N_21863);
or U25194 (N_25194,N_23527,N_23389);
nor U25195 (N_25195,N_22117,N_23171);
xor U25196 (N_25196,N_22147,N_23242);
nor U25197 (N_25197,N_23049,N_21087);
xnor U25198 (N_25198,N_21590,N_22058);
or U25199 (N_25199,N_21738,N_21955);
nand U25200 (N_25200,N_21922,N_23236);
nand U25201 (N_25201,N_22647,N_23153);
xnor U25202 (N_25202,N_23911,N_21491);
nor U25203 (N_25203,N_23894,N_23391);
and U25204 (N_25204,N_22333,N_23616);
nand U25205 (N_25205,N_21768,N_22827);
nand U25206 (N_25206,N_22151,N_22795);
nand U25207 (N_25207,N_23850,N_21403);
nor U25208 (N_25208,N_21275,N_22148);
nor U25209 (N_25209,N_21286,N_22304);
or U25210 (N_25210,N_22205,N_21187);
or U25211 (N_25211,N_23067,N_23884);
and U25212 (N_25212,N_21473,N_23870);
nand U25213 (N_25213,N_22560,N_22658);
nand U25214 (N_25214,N_23907,N_23166);
or U25215 (N_25215,N_21392,N_23342);
and U25216 (N_25216,N_23688,N_21040);
nor U25217 (N_25217,N_22213,N_22806);
nor U25218 (N_25218,N_23808,N_23443);
or U25219 (N_25219,N_21749,N_23657);
and U25220 (N_25220,N_22186,N_22199);
xnor U25221 (N_25221,N_22296,N_23791);
xor U25222 (N_25222,N_23696,N_21610);
or U25223 (N_25223,N_23144,N_22815);
nor U25224 (N_25224,N_22282,N_22712);
nand U25225 (N_25225,N_21785,N_21344);
nor U25226 (N_25226,N_23912,N_22043);
nor U25227 (N_25227,N_23445,N_21648);
nand U25228 (N_25228,N_22343,N_21886);
and U25229 (N_25229,N_22417,N_23033);
xor U25230 (N_25230,N_21567,N_22701);
nand U25231 (N_25231,N_21533,N_21778);
nor U25232 (N_25232,N_21426,N_23827);
or U25233 (N_25233,N_23643,N_22398);
nand U25234 (N_25234,N_22545,N_22237);
or U25235 (N_25235,N_23934,N_21386);
nand U25236 (N_25236,N_23366,N_22883);
and U25237 (N_25237,N_23712,N_23103);
nand U25238 (N_25238,N_22934,N_22223);
and U25239 (N_25239,N_21675,N_21110);
nand U25240 (N_25240,N_22389,N_23029);
and U25241 (N_25241,N_22276,N_23529);
nor U25242 (N_25242,N_23747,N_21089);
nand U25243 (N_25243,N_22005,N_23961);
nand U25244 (N_25244,N_22650,N_21468);
nand U25245 (N_25245,N_23828,N_23116);
and U25246 (N_25246,N_22400,N_22114);
nor U25247 (N_25247,N_21961,N_22214);
nand U25248 (N_25248,N_22536,N_22696);
xnor U25249 (N_25249,N_23174,N_21072);
xor U25250 (N_25250,N_23745,N_22176);
nor U25251 (N_25251,N_22652,N_23280);
xor U25252 (N_25252,N_23514,N_23424);
or U25253 (N_25253,N_21674,N_23143);
or U25254 (N_25254,N_22598,N_23012);
nand U25255 (N_25255,N_22853,N_21430);
nor U25256 (N_25256,N_21123,N_22898);
nor U25257 (N_25257,N_21520,N_23460);
nor U25258 (N_25258,N_21032,N_23086);
and U25259 (N_25259,N_23805,N_21859);
xor U25260 (N_25260,N_23627,N_21030);
or U25261 (N_25261,N_22365,N_21228);
xnor U25262 (N_25262,N_22790,N_23314);
nor U25263 (N_25263,N_21011,N_22482);
xnor U25264 (N_25264,N_21861,N_23493);
or U25265 (N_25265,N_22520,N_21234);
nand U25266 (N_25266,N_21466,N_23764);
and U25267 (N_25267,N_23328,N_22657);
and U25268 (N_25268,N_21867,N_22835);
xnor U25269 (N_25269,N_23102,N_22569);
and U25270 (N_25270,N_22256,N_21221);
xnor U25271 (N_25271,N_21399,N_22636);
nand U25272 (N_25272,N_22729,N_22060);
xor U25273 (N_25273,N_21607,N_22472);
or U25274 (N_25274,N_23285,N_23623);
and U25275 (N_25275,N_21784,N_23533);
nor U25276 (N_25276,N_23729,N_23478);
nor U25277 (N_25277,N_21852,N_23133);
xor U25278 (N_25278,N_21774,N_22307);
nor U25279 (N_25279,N_23939,N_23796);
xnor U25280 (N_25280,N_21150,N_21359);
nor U25281 (N_25281,N_21869,N_21077);
nand U25282 (N_25282,N_21577,N_21504);
or U25283 (N_25283,N_22695,N_23552);
xnor U25284 (N_25284,N_23798,N_22771);
or U25285 (N_25285,N_23875,N_23949);
xnor U25286 (N_25286,N_23270,N_22972);
nor U25287 (N_25287,N_21020,N_22020);
nand U25288 (N_25288,N_23100,N_23925);
nor U25289 (N_25289,N_22854,N_22945);
and U25290 (N_25290,N_23191,N_22617);
nor U25291 (N_25291,N_23847,N_23843);
xnor U25292 (N_25292,N_23809,N_21820);
nand U25293 (N_25293,N_22976,N_22008);
or U25294 (N_25294,N_21420,N_21952);
nor U25295 (N_25295,N_23840,N_21266);
or U25296 (N_25296,N_23160,N_22284);
nor U25297 (N_25297,N_23128,N_23826);
xor U25298 (N_25298,N_22037,N_21017);
nand U25299 (N_25299,N_23549,N_23027);
or U25300 (N_25300,N_22850,N_21929);
nand U25301 (N_25301,N_22157,N_21910);
xnor U25302 (N_25302,N_21153,N_23253);
nand U25303 (N_25303,N_23122,N_21435);
or U25304 (N_25304,N_21572,N_21384);
and U25305 (N_25305,N_23053,N_23050);
or U25306 (N_25306,N_23910,N_22629);
nor U25307 (N_25307,N_21247,N_22834);
and U25308 (N_25308,N_22159,N_22216);
nor U25309 (N_25309,N_22911,N_21428);
nand U25310 (N_25310,N_23589,N_22294);
or U25311 (N_25311,N_21117,N_22412);
xnor U25312 (N_25312,N_21623,N_21393);
and U25313 (N_25313,N_23956,N_23881);
or U25314 (N_25314,N_21721,N_22345);
nand U25315 (N_25315,N_21747,N_23324);
nor U25316 (N_25316,N_22800,N_23505);
xor U25317 (N_25317,N_21297,N_21987);
and U25318 (N_25318,N_22381,N_23238);
xor U25319 (N_25319,N_23311,N_23198);
xnor U25320 (N_25320,N_21149,N_21262);
nor U25321 (N_25321,N_23748,N_21350);
or U25322 (N_25322,N_21309,N_21606);
or U25323 (N_25323,N_23457,N_21700);
xor U25324 (N_25324,N_21723,N_22552);
and U25325 (N_25325,N_23030,N_21065);
or U25326 (N_25326,N_21239,N_23557);
or U25327 (N_25327,N_23298,N_21713);
xnor U25328 (N_25328,N_22034,N_21609);
or U25329 (N_25329,N_21310,N_22743);
nor U25330 (N_25330,N_21180,N_21079);
and U25331 (N_25331,N_21287,N_22051);
nor U25332 (N_25332,N_23245,N_23872);
nand U25333 (N_25333,N_23139,N_22357);
xor U25334 (N_25334,N_22097,N_23428);
xor U25335 (N_25335,N_23309,N_22272);
xnor U25336 (N_25336,N_23369,N_22555);
xor U25337 (N_25337,N_23669,N_23081);
xnor U25338 (N_25338,N_21148,N_21742);
or U25339 (N_25339,N_22373,N_23563);
xnor U25340 (N_25340,N_21931,N_23284);
xnor U25341 (N_25341,N_23230,N_22533);
xor U25342 (N_25342,N_23671,N_23024);
nand U25343 (N_25343,N_23054,N_21211);
xnor U25344 (N_25344,N_23009,N_22395);
and U25345 (N_25345,N_21871,N_22079);
xnor U25346 (N_25346,N_22665,N_21251);
nor U25347 (N_25347,N_22747,N_22632);
and U25348 (N_25348,N_21408,N_23438);
or U25349 (N_25349,N_21338,N_22849);
or U25350 (N_25350,N_23922,N_21240);
nor U25351 (N_25351,N_21816,N_21485);
or U25352 (N_25352,N_23407,N_23355);
nor U25353 (N_25353,N_21218,N_23996);
xor U25354 (N_25354,N_22491,N_22917);
nor U25355 (N_25355,N_21063,N_21828);
nand U25356 (N_25356,N_21711,N_21062);
and U25357 (N_25357,N_23714,N_23304);
nand U25358 (N_25358,N_21912,N_23991);
nor U25359 (N_25359,N_21652,N_23802);
xor U25360 (N_25360,N_21974,N_21560);
and U25361 (N_25361,N_22254,N_21892);
or U25362 (N_25362,N_22200,N_21391);
xor U25363 (N_25363,N_22143,N_22467);
nor U25364 (N_25364,N_21192,N_22433);
xor U25365 (N_25365,N_22773,N_22445);
or U25366 (N_25366,N_21942,N_21853);
and U25367 (N_25367,N_23261,N_21396);
or U25368 (N_25368,N_22023,N_22798);
xnor U25369 (N_25369,N_23234,N_22746);
nor U25370 (N_25370,N_21928,N_21730);
nand U25371 (N_25371,N_21879,N_23090);
or U25372 (N_25372,N_21256,N_21279);
xnor U25373 (N_25373,N_23351,N_21792);
xnor U25374 (N_25374,N_22959,N_21628);
or U25375 (N_25375,N_23415,N_21523);
and U25376 (N_25376,N_22507,N_22081);
xor U25377 (N_25377,N_23886,N_22719);
nand U25378 (N_25378,N_23427,N_21697);
and U25379 (N_25379,N_23321,N_21207);
nand U25380 (N_25380,N_21202,N_22110);
nor U25381 (N_25381,N_23083,N_22141);
and U25382 (N_25382,N_23902,N_21818);
and U25383 (N_25383,N_21484,N_22129);
and U25384 (N_25384,N_23154,N_23517);
nor U25385 (N_25385,N_21783,N_23599);
xor U25386 (N_25386,N_21619,N_22017);
or U25387 (N_25387,N_21477,N_23830);
or U25388 (N_25388,N_23976,N_22649);
or U25389 (N_25389,N_21529,N_22824);
and U25390 (N_25390,N_21226,N_21185);
and U25391 (N_25391,N_22823,N_21131);
nor U25392 (N_25392,N_21203,N_22816);
nand U25393 (N_25393,N_22504,N_21763);
and U25394 (N_25394,N_22554,N_23215);
and U25395 (N_25395,N_22941,N_22415);
or U25396 (N_25396,N_21019,N_22909);
xor U25397 (N_25397,N_21003,N_23673);
nor U25398 (N_25398,N_23535,N_22300);
and U25399 (N_25399,N_23435,N_21002);
or U25400 (N_25400,N_21536,N_23873);
nand U25401 (N_25401,N_22578,N_23977);
or U25402 (N_25402,N_23046,N_22763);
or U25403 (N_25403,N_22751,N_23734);
or U25404 (N_25404,N_23621,N_23676);
or U25405 (N_25405,N_23145,N_21605);
nand U25406 (N_25406,N_21624,N_23622);
nor U25407 (N_25407,N_22033,N_22310);
xnor U25408 (N_25408,N_22324,N_23310);
nor U25409 (N_25409,N_23823,N_22438);
nand U25410 (N_25410,N_21862,N_21840);
nand U25411 (N_25411,N_22355,N_23467);
or U25412 (N_25412,N_21295,N_23564);
nand U25413 (N_25413,N_23927,N_23767);
and U25414 (N_25414,N_23195,N_23228);
and U25415 (N_25415,N_23679,N_22543);
and U25416 (N_25416,N_21212,N_23382);
nor U25417 (N_25417,N_23943,N_22679);
and U25418 (N_25418,N_21949,N_23359);
xnor U25419 (N_25419,N_22860,N_21139);
or U25420 (N_25420,N_22628,N_21179);
nor U25421 (N_25421,N_22471,N_22682);
nand U25422 (N_25422,N_21441,N_22662);
xnor U25423 (N_25423,N_23307,N_22599);
nand U25424 (N_25424,N_22910,N_23783);
or U25425 (N_25425,N_23015,N_23702);
nor U25426 (N_25426,N_21373,N_23689);
nand U25427 (N_25427,N_21954,N_22935);
nand U25428 (N_25428,N_21280,N_22418);
and U25429 (N_25429,N_22821,N_22542);
nand U25430 (N_25430,N_21127,N_21856);
nor U25431 (N_25431,N_21172,N_22726);
xnor U25432 (N_25432,N_21246,N_23222);
xor U25433 (N_25433,N_22328,N_23330);
nor U25434 (N_25434,N_22677,N_22334);
xnor U25435 (N_25435,N_22523,N_22702);
xor U25436 (N_25436,N_21574,N_21268);
nor U25437 (N_25437,N_22787,N_22825);
or U25438 (N_25438,N_23035,N_22201);
nor U25439 (N_25439,N_22811,N_21383);
and U25440 (N_25440,N_21398,N_21788);
nor U25441 (N_25441,N_21532,N_23954);
and U25442 (N_25442,N_23337,N_23969);
or U25443 (N_25443,N_21743,N_21835);
nand U25444 (N_25444,N_22614,N_21455);
xnor U25445 (N_25445,N_23780,N_22247);
nor U25446 (N_25446,N_23720,N_21447);
nand U25447 (N_25447,N_21635,N_22955);
or U25448 (N_25448,N_22397,N_21811);
nor U25449 (N_25449,N_22595,N_23511);
xnor U25450 (N_25450,N_23279,N_22384);
nand U25451 (N_25451,N_23560,N_21197);
and U25452 (N_25452,N_23992,N_22970);
and U25453 (N_25453,N_21858,N_21489);
nand U25454 (N_25454,N_21191,N_21329);
xor U25455 (N_25455,N_22809,N_21177);
nand U25456 (N_25456,N_21302,N_23394);
nand U25457 (N_25457,N_23120,N_22968);
or U25458 (N_25458,N_23997,N_22158);
nand U25459 (N_25459,N_23158,N_21014);
nand U25460 (N_25460,N_21962,N_21071);
nor U25461 (N_25461,N_21805,N_21413);
nor U25462 (N_25462,N_21978,N_22456);
nand U25463 (N_25463,N_23392,N_21608);
nand U25464 (N_25464,N_22476,N_22168);
and U25465 (N_25465,N_23821,N_23784);
and U25466 (N_25466,N_22852,N_23302);
or U25467 (N_25467,N_21932,N_22740);
nor U25468 (N_25468,N_21640,N_22596);
and U25469 (N_25469,N_23340,N_22446);
or U25470 (N_25470,N_22508,N_21904);
nand U25471 (N_25471,N_23182,N_23271);
or U25472 (N_25472,N_22248,N_22903);
and U25473 (N_25473,N_22656,N_21363);
and U25474 (N_25474,N_23582,N_22098);
and U25475 (N_25475,N_21412,N_21057);
and U25476 (N_25476,N_23733,N_22031);
and U25477 (N_25477,N_21776,N_21812);
nand U25478 (N_25478,N_23220,N_23624);
and U25479 (N_25479,N_23724,N_22988);
and U25480 (N_25480,N_23248,N_22867);
xnor U25481 (N_25481,N_21693,N_22436);
or U25482 (N_25482,N_21767,N_23502);
nor U25483 (N_25483,N_21870,N_21637);
nand U25484 (N_25484,N_21201,N_23752);
nand U25485 (N_25485,N_22919,N_21530);
nand U25486 (N_25486,N_23626,N_23628);
or U25487 (N_25487,N_22527,N_23561);
xor U25488 (N_25488,N_21985,N_22584);
or U25489 (N_25489,N_23749,N_21964);
nor U25490 (N_25490,N_22331,N_23728);
xor U25491 (N_25491,N_22351,N_23082);
or U25492 (N_25492,N_21055,N_22947);
xnor U25493 (N_25493,N_21584,N_21464);
or U25494 (N_25494,N_21067,N_22225);
and U25495 (N_25495,N_22982,N_22172);
or U25496 (N_25496,N_22391,N_23199);
and U25497 (N_25497,N_21889,N_21772);
xnor U25498 (N_25498,N_23650,N_23508);
or U25499 (N_25499,N_21416,N_22590);
or U25500 (N_25500,N_22169,N_22581);
nand U25501 (N_25501,N_23260,N_21795);
nor U25502 (N_25502,N_21963,N_22608);
xnor U25503 (N_25503,N_23368,N_22489);
xor U25504 (N_25504,N_22854,N_22232);
nor U25505 (N_25505,N_23297,N_22641);
nor U25506 (N_25506,N_23563,N_21874);
and U25507 (N_25507,N_23252,N_21842);
xnor U25508 (N_25508,N_23531,N_23789);
nor U25509 (N_25509,N_21363,N_21255);
and U25510 (N_25510,N_23410,N_23110);
xor U25511 (N_25511,N_23622,N_21764);
nand U25512 (N_25512,N_23324,N_21275);
nand U25513 (N_25513,N_21156,N_23722);
nor U25514 (N_25514,N_23381,N_22877);
xnor U25515 (N_25515,N_22875,N_21196);
and U25516 (N_25516,N_21664,N_23125);
nor U25517 (N_25517,N_21727,N_23454);
nand U25518 (N_25518,N_23996,N_21289);
or U25519 (N_25519,N_21247,N_21975);
nand U25520 (N_25520,N_21541,N_21523);
xnor U25521 (N_25521,N_21311,N_21061);
xnor U25522 (N_25522,N_23627,N_21667);
xnor U25523 (N_25523,N_22682,N_22300);
or U25524 (N_25524,N_22650,N_22180);
xnor U25525 (N_25525,N_23320,N_21216);
nor U25526 (N_25526,N_22552,N_22476);
or U25527 (N_25527,N_22510,N_22667);
or U25528 (N_25528,N_23905,N_22272);
nor U25529 (N_25529,N_23448,N_22229);
or U25530 (N_25530,N_23211,N_21965);
and U25531 (N_25531,N_23311,N_23370);
nor U25532 (N_25532,N_23362,N_22968);
or U25533 (N_25533,N_22453,N_23214);
xor U25534 (N_25534,N_23923,N_21369);
or U25535 (N_25535,N_23256,N_23576);
and U25536 (N_25536,N_22940,N_23529);
xor U25537 (N_25537,N_21803,N_23005);
and U25538 (N_25538,N_22797,N_22827);
and U25539 (N_25539,N_22017,N_21261);
nor U25540 (N_25540,N_23150,N_23925);
or U25541 (N_25541,N_22595,N_22351);
or U25542 (N_25542,N_23943,N_21973);
nand U25543 (N_25543,N_22040,N_21760);
xor U25544 (N_25544,N_23106,N_23421);
nor U25545 (N_25545,N_21286,N_23529);
or U25546 (N_25546,N_23496,N_22456);
or U25547 (N_25547,N_22328,N_23877);
nor U25548 (N_25548,N_21600,N_21720);
nand U25549 (N_25549,N_22491,N_22067);
or U25550 (N_25550,N_22281,N_22752);
nor U25551 (N_25551,N_22863,N_23236);
nand U25552 (N_25552,N_22754,N_23000);
nand U25553 (N_25553,N_21882,N_23991);
nand U25554 (N_25554,N_21414,N_22450);
nor U25555 (N_25555,N_22191,N_22071);
or U25556 (N_25556,N_23924,N_23880);
nand U25557 (N_25557,N_22204,N_22029);
or U25558 (N_25558,N_21220,N_22753);
nand U25559 (N_25559,N_23447,N_23929);
nand U25560 (N_25560,N_22162,N_21225);
and U25561 (N_25561,N_21443,N_22948);
nor U25562 (N_25562,N_21705,N_21550);
and U25563 (N_25563,N_22157,N_22109);
nand U25564 (N_25564,N_21316,N_22134);
nand U25565 (N_25565,N_21654,N_22213);
nor U25566 (N_25566,N_21540,N_21922);
nand U25567 (N_25567,N_21891,N_21387);
nand U25568 (N_25568,N_23844,N_22653);
and U25569 (N_25569,N_22477,N_21357);
nor U25570 (N_25570,N_23414,N_21797);
and U25571 (N_25571,N_21784,N_23685);
and U25572 (N_25572,N_22756,N_21306);
xor U25573 (N_25573,N_22486,N_22823);
nand U25574 (N_25574,N_22918,N_23720);
or U25575 (N_25575,N_21552,N_23158);
xor U25576 (N_25576,N_21850,N_21375);
nor U25577 (N_25577,N_21707,N_23080);
nor U25578 (N_25578,N_22429,N_22948);
or U25579 (N_25579,N_22772,N_23902);
nor U25580 (N_25580,N_21364,N_23259);
nor U25581 (N_25581,N_23364,N_23341);
and U25582 (N_25582,N_21942,N_22206);
or U25583 (N_25583,N_23948,N_23011);
and U25584 (N_25584,N_22084,N_21000);
nand U25585 (N_25585,N_23050,N_22875);
and U25586 (N_25586,N_21558,N_21281);
or U25587 (N_25587,N_22748,N_23920);
and U25588 (N_25588,N_22464,N_21632);
nand U25589 (N_25589,N_21437,N_22584);
nand U25590 (N_25590,N_21440,N_21364);
nand U25591 (N_25591,N_23339,N_21388);
nor U25592 (N_25592,N_23083,N_22844);
xnor U25593 (N_25593,N_22604,N_21516);
or U25594 (N_25594,N_23134,N_23507);
or U25595 (N_25595,N_22404,N_22453);
or U25596 (N_25596,N_21872,N_22750);
nor U25597 (N_25597,N_22718,N_21303);
nor U25598 (N_25598,N_23807,N_23175);
xor U25599 (N_25599,N_22665,N_22498);
and U25600 (N_25600,N_22544,N_23006);
nor U25601 (N_25601,N_21991,N_23270);
xnor U25602 (N_25602,N_23695,N_21790);
and U25603 (N_25603,N_22792,N_22373);
or U25604 (N_25604,N_23767,N_22367);
nor U25605 (N_25605,N_23184,N_21601);
or U25606 (N_25606,N_22639,N_22187);
nand U25607 (N_25607,N_22616,N_22276);
and U25608 (N_25608,N_22716,N_23685);
and U25609 (N_25609,N_23186,N_21770);
or U25610 (N_25610,N_22233,N_22876);
xnor U25611 (N_25611,N_21933,N_21865);
and U25612 (N_25612,N_21168,N_21576);
or U25613 (N_25613,N_22974,N_23339);
and U25614 (N_25614,N_23565,N_22071);
or U25615 (N_25615,N_22025,N_22942);
and U25616 (N_25616,N_23803,N_23526);
or U25617 (N_25617,N_23035,N_21316);
nor U25618 (N_25618,N_23690,N_22603);
nor U25619 (N_25619,N_23524,N_23861);
or U25620 (N_25620,N_21981,N_22267);
nor U25621 (N_25621,N_23004,N_23256);
and U25622 (N_25622,N_22584,N_23145);
xor U25623 (N_25623,N_22300,N_21161);
nand U25624 (N_25624,N_22557,N_21875);
and U25625 (N_25625,N_23376,N_22287);
nor U25626 (N_25626,N_22336,N_23250);
nor U25627 (N_25627,N_23540,N_21394);
xnor U25628 (N_25628,N_22663,N_22286);
and U25629 (N_25629,N_22643,N_22742);
nor U25630 (N_25630,N_21879,N_22706);
or U25631 (N_25631,N_22735,N_23828);
and U25632 (N_25632,N_22208,N_22817);
and U25633 (N_25633,N_21019,N_22190);
and U25634 (N_25634,N_22919,N_23220);
nand U25635 (N_25635,N_21762,N_22054);
and U25636 (N_25636,N_23602,N_21861);
or U25637 (N_25637,N_21950,N_22556);
or U25638 (N_25638,N_22142,N_21056);
nor U25639 (N_25639,N_21245,N_22976);
and U25640 (N_25640,N_23927,N_21848);
nor U25641 (N_25641,N_23183,N_22601);
xnor U25642 (N_25642,N_22882,N_21746);
xor U25643 (N_25643,N_22403,N_23633);
nor U25644 (N_25644,N_23060,N_22046);
and U25645 (N_25645,N_22594,N_22567);
and U25646 (N_25646,N_22657,N_21132);
nor U25647 (N_25647,N_23447,N_22965);
or U25648 (N_25648,N_22884,N_21336);
or U25649 (N_25649,N_23699,N_22975);
nor U25650 (N_25650,N_21732,N_22330);
or U25651 (N_25651,N_23135,N_23641);
nor U25652 (N_25652,N_23053,N_23834);
and U25653 (N_25653,N_23275,N_22464);
xor U25654 (N_25654,N_21585,N_21214);
and U25655 (N_25655,N_22655,N_22970);
nand U25656 (N_25656,N_23217,N_23508);
nand U25657 (N_25657,N_22223,N_23987);
and U25658 (N_25658,N_21033,N_21805);
xnor U25659 (N_25659,N_22189,N_22703);
and U25660 (N_25660,N_21327,N_22482);
xor U25661 (N_25661,N_21694,N_23284);
xor U25662 (N_25662,N_21561,N_22338);
and U25663 (N_25663,N_21608,N_23568);
nor U25664 (N_25664,N_23581,N_23962);
nor U25665 (N_25665,N_21569,N_21649);
nand U25666 (N_25666,N_22926,N_21192);
nor U25667 (N_25667,N_21034,N_21769);
xnor U25668 (N_25668,N_21384,N_23504);
and U25669 (N_25669,N_23297,N_21003);
or U25670 (N_25670,N_23890,N_23438);
nand U25671 (N_25671,N_21199,N_21251);
or U25672 (N_25672,N_22237,N_23090);
and U25673 (N_25673,N_22242,N_23715);
and U25674 (N_25674,N_21249,N_21277);
or U25675 (N_25675,N_22301,N_21118);
nand U25676 (N_25676,N_22459,N_22754);
xor U25677 (N_25677,N_23197,N_23834);
xnor U25678 (N_25678,N_23132,N_21419);
xnor U25679 (N_25679,N_23089,N_21954);
xor U25680 (N_25680,N_23175,N_21387);
xnor U25681 (N_25681,N_21572,N_23323);
xnor U25682 (N_25682,N_23767,N_22322);
xor U25683 (N_25683,N_23938,N_22509);
nor U25684 (N_25684,N_22460,N_22970);
nand U25685 (N_25685,N_23086,N_22082);
and U25686 (N_25686,N_22413,N_22492);
nor U25687 (N_25687,N_21134,N_21257);
or U25688 (N_25688,N_22961,N_22997);
xnor U25689 (N_25689,N_23943,N_22771);
or U25690 (N_25690,N_23972,N_21164);
nand U25691 (N_25691,N_23066,N_21950);
xor U25692 (N_25692,N_21305,N_21253);
and U25693 (N_25693,N_23248,N_23059);
or U25694 (N_25694,N_22230,N_22650);
or U25695 (N_25695,N_22301,N_21721);
nand U25696 (N_25696,N_23615,N_22317);
or U25697 (N_25697,N_21944,N_23173);
nor U25698 (N_25698,N_21798,N_21299);
xnor U25699 (N_25699,N_23931,N_21372);
xnor U25700 (N_25700,N_21419,N_22646);
nor U25701 (N_25701,N_23472,N_22107);
and U25702 (N_25702,N_22528,N_23866);
or U25703 (N_25703,N_23460,N_22606);
nor U25704 (N_25704,N_23486,N_21485);
nand U25705 (N_25705,N_23716,N_23213);
and U25706 (N_25706,N_21974,N_23723);
and U25707 (N_25707,N_21256,N_23799);
nor U25708 (N_25708,N_23582,N_22082);
and U25709 (N_25709,N_21332,N_23424);
xor U25710 (N_25710,N_21788,N_21477);
nand U25711 (N_25711,N_21704,N_22247);
nand U25712 (N_25712,N_21204,N_22294);
xor U25713 (N_25713,N_22249,N_21462);
nand U25714 (N_25714,N_21321,N_22910);
nor U25715 (N_25715,N_21859,N_22410);
nand U25716 (N_25716,N_23078,N_21630);
nand U25717 (N_25717,N_23257,N_21372);
nand U25718 (N_25718,N_21553,N_23358);
and U25719 (N_25719,N_21321,N_21160);
or U25720 (N_25720,N_21158,N_22655);
nand U25721 (N_25721,N_22223,N_22040);
nand U25722 (N_25722,N_22378,N_23873);
and U25723 (N_25723,N_21920,N_21178);
or U25724 (N_25724,N_21043,N_21808);
or U25725 (N_25725,N_23943,N_21234);
and U25726 (N_25726,N_21113,N_23788);
xor U25727 (N_25727,N_23398,N_23496);
nor U25728 (N_25728,N_21860,N_21483);
nor U25729 (N_25729,N_23648,N_21775);
and U25730 (N_25730,N_23865,N_23453);
xor U25731 (N_25731,N_23607,N_23306);
and U25732 (N_25732,N_22431,N_22837);
or U25733 (N_25733,N_22752,N_23759);
nand U25734 (N_25734,N_23515,N_23300);
or U25735 (N_25735,N_22977,N_21012);
nor U25736 (N_25736,N_23564,N_23812);
or U25737 (N_25737,N_22209,N_21057);
nand U25738 (N_25738,N_21839,N_22971);
or U25739 (N_25739,N_22322,N_21391);
nand U25740 (N_25740,N_21547,N_22772);
nor U25741 (N_25741,N_22480,N_21839);
or U25742 (N_25742,N_21587,N_22797);
or U25743 (N_25743,N_22329,N_22079);
nor U25744 (N_25744,N_22241,N_21301);
nor U25745 (N_25745,N_23471,N_23902);
and U25746 (N_25746,N_22262,N_21050);
nand U25747 (N_25747,N_23144,N_22476);
and U25748 (N_25748,N_23923,N_23443);
and U25749 (N_25749,N_23613,N_21387);
nor U25750 (N_25750,N_21803,N_21819);
xnor U25751 (N_25751,N_21389,N_22723);
or U25752 (N_25752,N_21235,N_21897);
nor U25753 (N_25753,N_23774,N_22359);
nand U25754 (N_25754,N_21274,N_22587);
or U25755 (N_25755,N_22409,N_22374);
nand U25756 (N_25756,N_21881,N_22706);
nand U25757 (N_25757,N_23289,N_22871);
and U25758 (N_25758,N_23970,N_22053);
or U25759 (N_25759,N_21837,N_23862);
or U25760 (N_25760,N_23687,N_21771);
xnor U25761 (N_25761,N_21720,N_22158);
nand U25762 (N_25762,N_23392,N_23391);
nor U25763 (N_25763,N_21119,N_23619);
nand U25764 (N_25764,N_23317,N_22190);
xnor U25765 (N_25765,N_23815,N_21012);
xor U25766 (N_25766,N_21275,N_22186);
or U25767 (N_25767,N_21444,N_22762);
and U25768 (N_25768,N_21425,N_22274);
xor U25769 (N_25769,N_21226,N_23012);
nand U25770 (N_25770,N_21997,N_21992);
nor U25771 (N_25771,N_21349,N_23308);
xor U25772 (N_25772,N_21715,N_22278);
and U25773 (N_25773,N_22888,N_21020);
and U25774 (N_25774,N_21740,N_22394);
xnor U25775 (N_25775,N_22167,N_23742);
nor U25776 (N_25776,N_21814,N_21869);
xnor U25777 (N_25777,N_23357,N_21345);
and U25778 (N_25778,N_22429,N_22669);
nor U25779 (N_25779,N_21023,N_22532);
nor U25780 (N_25780,N_22243,N_22284);
nand U25781 (N_25781,N_21672,N_21483);
and U25782 (N_25782,N_22723,N_21914);
xor U25783 (N_25783,N_22403,N_21732);
or U25784 (N_25784,N_22383,N_23849);
nor U25785 (N_25785,N_23309,N_21883);
and U25786 (N_25786,N_21781,N_23043);
or U25787 (N_25787,N_23027,N_22138);
and U25788 (N_25788,N_22566,N_21420);
or U25789 (N_25789,N_22462,N_23020);
xnor U25790 (N_25790,N_23554,N_23838);
nor U25791 (N_25791,N_21612,N_21768);
and U25792 (N_25792,N_23440,N_21222);
xnor U25793 (N_25793,N_22908,N_21263);
nor U25794 (N_25794,N_23267,N_21715);
nand U25795 (N_25795,N_23591,N_22904);
nand U25796 (N_25796,N_22660,N_23527);
nor U25797 (N_25797,N_23537,N_23553);
nand U25798 (N_25798,N_22607,N_23710);
nor U25799 (N_25799,N_23362,N_23103);
or U25800 (N_25800,N_22008,N_23448);
or U25801 (N_25801,N_22077,N_22372);
nand U25802 (N_25802,N_21844,N_21262);
nor U25803 (N_25803,N_23387,N_21353);
nor U25804 (N_25804,N_22491,N_22924);
and U25805 (N_25805,N_21396,N_23829);
or U25806 (N_25806,N_21400,N_23771);
and U25807 (N_25807,N_23155,N_21191);
or U25808 (N_25808,N_22748,N_21287);
nand U25809 (N_25809,N_23558,N_23512);
xor U25810 (N_25810,N_22995,N_22192);
nor U25811 (N_25811,N_22579,N_22185);
nand U25812 (N_25812,N_23778,N_22012);
nand U25813 (N_25813,N_21345,N_21967);
xor U25814 (N_25814,N_23151,N_22598);
nor U25815 (N_25815,N_22008,N_23481);
and U25816 (N_25816,N_23815,N_23716);
nor U25817 (N_25817,N_23727,N_21805);
or U25818 (N_25818,N_23791,N_23641);
or U25819 (N_25819,N_23265,N_23552);
nor U25820 (N_25820,N_21191,N_21177);
and U25821 (N_25821,N_23845,N_22417);
and U25822 (N_25822,N_21574,N_23208);
and U25823 (N_25823,N_23815,N_23635);
nand U25824 (N_25824,N_21123,N_22377);
or U25825 (N_25825,N_22141,N_22609);
nand U25826 (N_25826,N_21087,N_23510);
or U25827 (N_25827,N_22238,N_21812);
nand U25828 (N_25828,N_22020,N_22653);
nor U25829 (N_25829,N_21389,N_22267);
xnor U25830 (N_25830,N_22022,N_22285);
and U25831 (N_25831,N_23844,N_23955);
xor U25832 (N_25832,N_22302,N_23777);
or U25833 (N_25833,N_22127,N_23907);
xor U25834 (N_25834,N_23854,N_22806);
and U25835 (N_25835,N_23842,N_23805);
xor U25836 (N_25836,N_23681,N_21482);
or U25837 (N_25837,N_23004,N_23035);
nand U25838 (N_25838,N_22008,N_22860);
nand U25839 (N_25839,N_22227,N_22051);
and U25840 (N_25840,N_22511,N_21494);
nand U25841 (N_25841,N_21437,N_21132);
and U25842 (N_25842,N_23780,N_21094);
nor U25843 (N_25843,N_21238,N_23266);
nor U25844 (N_25844,N_22385,N_23601);
xnor U25845 (N_25845,N_22269,N_23023);
nor U25846 (N_25846,N_22632,N_21451);
nand U25847 (N_25847,N_22548,N_21159);
and U25848 (N_25848,N_21609,N_23823);
nor U25849 (N_25849,N_21427,N_21423);
nand U25850 (N_25850,N_21325,N_22882);
nor U25851 (N_25851,N_23676,N_22940);
and U25852 (N_25852,N_21890,N_22535);
nor U25853 (N_25853,N_23648,N_23810);
nand U25854 (N_25854,N_22067,N_21170);
or U25855 (N_25855,N_22908,N_23913);
and U25856 (N_25856,N_23235,N_23247);
or U25857 (N_25857,N_21758,N_22872);
and U25858 (N_25858,N_23600,N_22167);
nand U25859 (N_25859,N_23086,N_22284);
or U25860 (N_25860,N_23622,N_23165);
xnor U25861 (N_25861,N_23697,N_22143);
and U25862 (N_25862,N_22321,N_22245);
xnor U25863 (N_25863,N_21081,N_21360);
nor U25864 (N_25864,N_21768,N_21301);
xnor U25865 (N_25865,N_22578,N_23312);
or U25866 (N_25866,N_21902,N_21549);
xnor U25867 (N_25867,N_23981,N_22159);
or U25868 (N_25868,N_23528,N_22690);
and U25869 (N_25869,N_23852,N_21313);
xor U25870 (N_25870,N_23054,N_22949);
and U25871 (N_25871,N_22606,N_22682);
or U25872 (N_25872,N_21773,N_22238);
nand U25873 (N_25873,N_21290,N_23279);
and U25874 (N_25874,N_22504,N_23663);
or U25875 (N_25875,N_21764,N_21338);
or U25876 (N_25876,N_22049,N_22045);
nor U25877 (N_25877,N_22062,N_22679);
or U25878 (N_25878,N_22916,N_23128);
and U25879 (N_25879,N_21810,N_22828);
or U25880 (N_25880,N_23128,N_23646);
or U25881 (N_25881,N_22085,N_21693);
nand U25882 (N_25882,N_21889,N_22827);
nor U25883 (N_25883,N_23635,N_23439);
nand U25884 (N_25884,N_22596,N_23039);
nor U25885 (N_25885,N_23776,N_22233);
or U25886 (N_25886,N_21385,N_21673);
nand U25887 (N_25887,N_22505,N_21506);
or U25888 (N_25888,N_23591,N_23103);
nand U25889 (N_25889,N_23767,N_21648);
nand U25890 (N_25890,N_21912,N_21298);
or U25891 (N_25891,N_22143,N_23709);
and U25892 (N_25892,N_23028,N_23725);
and U25893 (N_25893,N_22184,N_21004);
and U25894 (N_25894,N_23932,N_22802);
or U25895 (N_25895,N_21313,N_21208);
and U25896 (N_25896,N_22476,N_23449);
nor U25897 (N_25897,N_21982,N_22388);
nand U25898 (N_25898,N_22885,N_22235);
or U25899 (N_25899,N_21056,N_21315);
nor U25900 (N_25900,N_23301,N_22446);
or U25901 (N_25901,N_23027,N_23899);
xnor U25902 (N_25902,N_22437,N_22265);
and U25903 (N_25903,N_21965,N_21630);
and U25904 (N_25904,N_23265,N_22995);
or U25905 (N_25905,N_21630,N_23576);
nand U25906 (N_25906,N_21656,N_22359);
xor U25907 (N_25907,N_22607,N_21561);
and U25908 (N_25908,N_21429,N_22866);
nand U25909 (N_25909,N_23728,N_22528);
and U25910 (N_25910,N_22135,N_22680);
nand U25911 (N_25911,N_23285,N_21590);
and U25912 (N_25912,N_21508,N_22443);
nand U25913 (N_25913,N_23072,N_21927);
nor U25914 (N_25914,N_23709,N_21555);
and U25915 (N_25915,N_22881,N_21402);
and U25916 (N_25916,N_23979,N_21751);
or U25917 (N_25917,N_21475,N_21314);
nor U25918 (N_25918,N_23775,N_23488);
xnor U25919 (N_25919,N_22911,N_23038);
nand U25920 (N_25920,N_23285,N_22594);
nor U25921 (N_25921,N_23399,N_23682);
nor U25922 (N_25922,N_22235,N_21553);
nand U25923 (N_25923,N_22864,N_23610);
nor U25924 (N_25924,N_22463,N_21446);
or U25925 (N_25925,N_23070,N_21277);
and U25926 (N_25926,N_23851,N_22192);
or U25927 (N_25927,N_22266,N_22381);
xor U25928 (N_25928,N_21055,N_23423);
or U25929 (N_25929,N_23262,N_23737);
nor U25930 (N_25930,N_22949,N_21240);
or U25931 (N_25931,N_21880,N_21556);
xnor U25932 (N_25932,N_23943,N_22705);
or U25933 (N_25933,N_21527,N_22482);
nor U25934 (N_25934,N_22183,N_23552);
nor U25935 (N_25935,N_23895,N_23928);
and U25936 (N_25936,N_21137,N_23581);
or U25937 (N_25937,N_23769,N_23863);
xnor U25938 (N_25938,N_23429,N_23866);
nor U25939 (N_25939,N_21432,N_21278);
xor U25940 (N_25940,N_23374,N_22849);
or U25941 (N_25941,N_22095,N_21182);
nor U25942 (N_25942,N_21308,N_23497);
nand U25943 (N_25943,N_22685,N_22073);
nand U25944 (N_25944,N_21899,N_21506);
and U25945 (N_25945,N_21178,N_22809);
or U25946 (N_25946,N_23651,N_23822);
xnor U25947 (N_25947,N_21770,N_22097);
nor U25948 (N_25948,N_21382,N_21718);
nor U25949 (N_25949,N_23595,N_21875);
or U25950 (N_25950,N_21726,N_23615);
xnor U25951 (N_25951,N_22076,N_22763);
nor U25952 (N_25952,N_22207,N_22251);
xor U25953 (N_25953,N_22076,N_22374);
or U25954 (N_25954,N_21871,N_22162);
or U25955 (N_25955,N_22750,N_23008);
and U25956 (N_25956,N_21114,N_23231);
nor U25957 (N_25957,N_23161,N_22576);
nand U25958 (N_25958,N_23837,N_21353);
nand U25959 (N_25959,N_23859,N_22907);
xnor U25960 (N_25960,N_21688,N_23234);
nand U25961 (N_25961,N_22251,N_22735);
and U25962 (N_25962,N_23691,N_22037);
nor U25963 (N_25963,N_21070,N_22466);
xnor U25964 (N_25964,N_23796,N_21463);
or U25965 (N_25965,N_21813,N_22727);
and U25966 (N_25966,N_23636,N_22149);
nor U25967 (N_25967,N_23770,N_21796);
nand U25968 (N_25968,N_22187,N_21976);
nor U25969 (N_25969,N_22944,N_21502);
or U25970 (N_25970,N_23525,N_22579);
xor U25971 (N_25971,N_21480,N_23060);
nand U25972 (N_25972,N_22920,N_21745);
nor U25973 (N_25973,N_21926,N_23504);
nand U25974 (N_25974,N_23471,N_23835);
nand U25975 (N_25975,N_22295,N_23516);
and U25976 (N_25976,N_22580,N_23959);
and U25977 (N_25977,N_23250,N_22474);
and U25978 (N_25978,N_21700,N_22433);
or U25979 (N_25979,N_22915,N_22652);
nand U25980 (N_25980,N_23494,N_21152);
or U25981 (N_25981,N_21965,N_22127);
nand U25982 (N_25982,N_23102,N_22953);
nand U25983 (N_25983,N_23012,N_23597);
nor U25984 (N_25984,N_21310,N_21512);
and U25985 (N_25985,N_23256,N_22224);
and U25986 (N_25986,N_22769,N_22123);
and U25987 (N_25987,N_22427,N_22398);
nand U25988 (N_25988,N_21554,N_21023);
and U25989 (N_25989,N_21546,N_22711);
and U25990 (N_25990,N_23919,N_23130);
or U25991 (N_25991,N_23850,N_23431);
nor U25992 (N_25992,N_22808,N_22121);
xnor U25993 (N_25993,N_21346,N_23030);
or U25994 (N_25994,N_23903,N_23791);
xnor U25995 (N_25995,N_21519,N_21611);
nand U25996 (N_25996,N_21133,N_22265);
or U25997 (N_25997,N_22500,N_21488);
nand U25998 (N_25998,N_21147,N_22955);
nor U25999 (N_25999,N_23273,N_22105);
nor U26000 (N_26000,N_22925,N_21884);
nand U26001 (N_26001,N_22360,N_23762);
xor U26002 (N_26002,N_21853,N_23244);
or U26003 (N_26003,N_23783,N_21156);
and U26004 (N_26004,N_22631,N_23316);
xnor U26005 (N_26005,N_21948,N_21338);
nand U26006 (N_26006,N_21767,N_22749);
nor U26007 (N_26007,N_22866,N_23546);
xnor U26008 (N_26008,N_21637,N_22491);
and U26009 (N_26009,N_23269,N_21524);
nor U26010 (N_26010,N_21720,N_21947);
nand U26011 (N_26011,N_21090,N_23963);
and U26012 (N_26012,N_21885,N_22122);
and U26013 (N_26013,N_21854,N_22977);
and U26014 (N_26014,N_23632,N_21831);
and U26015 (N_26015,N_21887,N_22194);
or U26016 (N_26016,N_23508,N_23923);
nand U26017 (N_26017,N_21835,N_22515);
nand U26018 (N_26018,N_22435,N_22164);
and U26019 (N_26019,N_21696,N_22126);
and U26020 (N_26020,N_23944,N_23151);
xnor U26021 (N_26021,N_23836,N_22952);
xnor U26022 (N_26022,N_22039,N_21293);
xor U26023 (N_26023,N_21424,N_23793);
or U26024 (N_26024,N_22374,N_21928);
nand U26025 (N_26025,N_22394,N_22539);
or U26026 (N_26026,N_22415,N_22129);
nand U26027 (N_26027,N_21598,N_22840);
or U26028 (N_26028,N_21905,N_23172);
or U26029 (N_26029,N_23377,N_22246);
nor U26030 (N_26030,N_22345,N_21951);
xnor U26031 (N_26031,N_21818,N_23443);
and U26032 (N_26032,N_22005,N_22965);
nor U26033 (N_26033,N_23271,N_21438);
nor U26034 (N_26034,N_22492,N_22581);
nor U26035 (N_26035,N_22217,N_23288);
nand U26036 (N_26036,N_23113,N_23177);
nand U26037 (N_26037,N_22141,N_23214);
or U26038 (N_26038,N_22443,N_22721);
and U26039 (N_26039,N_21306,N_21204);
xnor U26040 (N_26040,N_23368,N_22931);
or U26041 (N_26041,N_22801,N_23109);
nor U26042 (N_26042,N_23428,N_22844);
xor U26043 (N_26043,N_23844,N_21149);
nand U26044 (N_26044,N_23336,N_23407);
nand U26045 (N_26045,N_23765,N_22514);
and U26046 (N_26046,N_21780,N_23191);
nand U26047 (N_26047,N_23563,N_23613);
and U26048 (N_26048,N_21428,N_23643);
and U26049 (N_26049,N_23537,N_21399);
and U26050 (N_26050,N_22557,N_22989);
xor U26051 (N_26051,N_22716,N_21909);
or U26052 (N_26052,N_21541,N_21322);
xor U26053 (N_26053,N_22499,N_22105);
xnor U26054 (N_26054,N_22201,N_22448);
and U26055 (N_26055,N_21328,N_22274);
nand U26056 (N_26056,N_21991,N_22288);
or U26057 (N_26057,N_22026,N_23670);
nor U26058 (N_26058,N_21535,N_23151);
xor U26059 (N_26059,N_21189,N_21411);
and U26060 (N_26060,N_21370,N_23391);
nor U26061 (N_26061,N_23434,N_21484);
or U26062 (N_26062,N_23782,N_23818);
or U26063 (N_26063,N_21483,N_22082);
xor U26064 (N_26064,N_23873,N_21051);
nand U26065 (N_26065,N_21429,N_22351);
nor U26066 (N_26066,N_22688,N_23288);
xor U26067 (N_26067,N_23112,N_22586);
nor U26068 (N_26068,N_21283,N_21867);
or U26069 (N_26069,N_22199,N_23606);
or U26070 (N_26070,N_22996,N_23331);
xor U26071 (N_26071,N_21986,N_23374);
nand U26072 (N_26072,N_22327,N_22947);
xnor U26073 (N_26073,N_23866,N_21164);
or U26074 (N_26074,N_21218,N_21578);
xnor U26075 (N_26075,N_21757,N_21834);
nand U26076 (N_26076,N_22536,N_21068);
and U26077 (N_26077,N_23583,N_21757);
xnor U26078 (N_26078,N_22198,N_21933);
or U26079 (N_26079,N_21513,N_21354);
or U26080 (N_26080,N_23464,N_22143);
nand U26081 (N_26081,N_22234,N_21099);
xor U26082 (N_26082,N_23378,N_23752);
xnor U26083 (N_26083,N_23645,N_22203);
nand U26084 (N_26084,N_23367,N_22973);
and U26085 (N_26085,N_21333,N_21814);
xnor U26086 (N_26086,N_21088,N_22051);
nand U26087 (N_26087,N_22021,N_21020);
and U26088 (N_26088,N_21720,N_21778);
or U26089 (N_26089,N_23106,N_23149);
nor U26090 (N_26090,N_22684,N_23478);
or U26091 (N_26091,N_23367,N_23038);
nand U26092 (N_26092,N_22906,N_22473);
nand U26093 (N_26093,N_21842,N_23644);
and U26094 (N_26094,N_22033,N_23752);
xor U26095 (N_26095,N_22374,N_22780);
nor U26096 (N_26096,N_23793,N_23227);
nor U26097 (N_26097,N_21919,N_21637);
nand U26098 (N_26098,N_22829,N_21867);
and U26099 (N_26099,N_22481,N_23962);
nand U26100 (N_26100,N_22273,N_21014);
nand U26101 (N_26101,N_23539,N_22752);
and U26102 (N_26102,N_21598,N_23062);
nand U26103 (N_26103,N_23677,N_21513);
nor U26104 (N_26104,N_21465,N_22452);
or U26105 (N_26105,N_22518,N_22280);
nand U26106 (N_26106,N_23306,N_21047);
and U26107 (N_26107,N_21795,N_22545);
nand U26108 (N_26108,N_23009,N_22234);
and U26109 (N_26109,N_21423,N_22090);
and U26110 (N_26110,N_22692,N_23171);
or U26111 (N_26111,N_21072,N_21528);
and U26112 (N_26112,N_21403,N_21390);
nand U26113 (N_26113,N_22870,N_22974);
nand U26114 (N_26114,N_22663,N_23922);
or U26115 (N_26115,N_23896,N_21266);
and U26116 (N_26116,N_21452,N_23999);
nor U26117 (N_26117,N_21220,N_21407);
xnor U26118 (N_26118,N_21334,N_21868);
and U26119 (N_26119,N_22527,N_22765);
nor U26120 (N_26120,N_22600,N_23462);
nand U26121 (N_26121,N_21849,N_22098);
and U26122 (N_26122,N_23036,N_23008);
xnor U26123 (N_26123,N_23782,N_23580);
or U26124 (N_26124,N_22766,N_22180);
nor U26125 (N_26125,N_22106,N_22470);
nor U26126 (N_26126,N_23308,N_23423);
and U26127 (N_26127,N_23262,N_21383);
nor U26128 (N_26128,N_22874,N_21494);
xor U26129 (N_26129,N_23154,N_22088);
nor U26130 (N_26130,N_23736,N_23808);
or U26131 (N_26131,N_22828,N_22696);
and U26132 (N_26132,N_23027,N_22132);
and U26133 (N_26133,N_23477,N_23723);
nor U26134 (N_26134,N_22143,N_22614);
or U26135 (N_26135,N_23252,N_23830);
nor U26136 (N_26136,N_22759,N_22367);
xor U26137 (N_26137,N_23076,N_21179);
or U26138 (N_26138,N_22049,N_23869);
or U26139 (N_26139,N_23303,N_22413);
or U26140 (N_26140,N_21059,N_21863);
nor U26141 (N_26141,N_21606,N_21903);
and U26142 (N_26142,N_22508,N_22156);
nor U26143 (N_26143,N_23224,N_21711);
or U26144 (N_26144,N_23248,N_23025);
nand U26145 (N_26145,N_22987,N_22341);
or U26146 (N_26146,N_23618,N_22926);
or U26147 (N_26147,N_22079,N_21755);
nor U26148 (N_26148,N_23232,N_22547);
nor U26149 (N_26149,N_21697,N_23641);
or U26150 (N_26150,N_22892,N_23024);
and U26151 (N_26151,N_21254,N_23529);
nor U26152 (N_26152,N_21718,N_22652);
or U26153 (N_26153,N_22345,N_21545);
nor U26154 (N_26154,N_21291,N_23177);
nor U26155 (N_26155,N_23453,N_21508);
and U26156 (N_26156,N_22239,N_22900);
and U26157 (N_26157,N_22857,N_22146);
or U26158 (N_26158,N_21022,N_22366);
xnor U26159 (N_26159,N_21874,N_23317);
nor U26160 (N_26160,N_21326,N_22257);
and U26161 (N_26161,N_21152,N_23698);
xnor U26162 (N_26162,N_21793,N_23576);
nor U26163 (N_26163,N_23797,N_23263);
and U26164 (N_26164,N_22330,N_21707);
xor U26165 (N_26165,N_21362,N_23379);
nand U26166 (N_26166,N_22540,N_23842);
nand U26167 (N_26167,N_22688,N_22707);
nand U26168 (N_26168,N_23460,N_21493);
or U26169 (N_26169,N_23786,N_21855);
xnor U26170 (N_26170,N_22318,N_23595);
or U26171 (N_26171,N_21997,N_22972);
and U26172 (N_26172,N_22593,N_22000);
or U26173 (N_26173,N_22048,N_22684);
and U26174 (N_26174,N_22413,N_22460);
or U26175 (N_26175,N_23358,N_21872);
nor U26176 (N_26176,N_23593,N_23207);
nor U26177 (N_26177,N_23289,N_23658);
and U26178 (N_26178,N_23393,N_21772);
nand U26179 (N_26179,N_23128,N_21513);
xnor U26180 (N_26180,N_21014,N_22971);
or U26181 (N_26181,N_23088,N_22545);
nand U26182 (N_26182,N_22073,N_21275);
or U26183 (N_26183,N_23397,N_22067);
or U26184 (N_26184,N_22386,N_22433);
nor U26185 (N_26185,N_21930,N_22641);
nor U26186 (N_26186,N_21337,N_21155);
nand U26187 (N_26187,N_21126,N_22055);
nand U26188 (N_26188,N_22211,N_21973);
nand U26189 (N_26189,N_23555,N_23944);
nand U26190 (N_26190,N_22073,N_22964);
nand U26191 (N_26191,N_21674,N_22405);
nand U26192 (N_26192,N_22789,N_22934);
and U26193 (N_26193,N_23753,N_21540);
nor U26194 (N_26194,N_23562,N_22417);
xor U26195 (N_26195,N_22082,N_21144);
xnor U26196 (N_26196,N_22724,N_22187);
xor U26197 (N_26197,N_23632,N_22858);
nand U26198 (N_26198,N_21931,N_23108);
and U26199 (N_26199,N_22647,N_21256);
and U26200 (N_26200,N_22046,N_22342);
nand U26201 (N_26201,N_21872,N_23954);
xor U26202 (N_26202,N_23081,N_21878);
and U26203 (N_26203,N_21821,N_22802);
xor U26204 (N_26204,N_22925,N_23243);
and U26205 (N_26205,N_21760,N_23411);
xnor U26206 (N_26206,N_22074,N_22658);
or U26207 (N_26207,N_23489,N_21712);
or U26208 (N_26208,N_23641,N_23152);
and U26209 (N_26209,N_22183,N_22541);
nor U26210 (N_26210,N_21177,N_21474);
nand U26211 (N_26211,N_21368,N_22882);
and U26212 (N_26212,N_23893,N_23322);
nand U26213 (N_26213,N_22950,N_22208);
and U26214 (N_26214,N_21086,N_21201);
xor U26215 (N_26215,N_22091,N_23296);
or U26216 (N_26216,N_21779,N_21806);
or U26217 (N_26217,N_23446,N_21212);
xnor U26218 (N_26218,N_23741,N_21427);
nand U26219 (N_26219,N_21832,N_22511);
xor U26220 (N_26220,N_21927,N_23479);
or U26221 (N_26221,N_23932,N_21889);
nor U26222 (N_26222,N_22081,N_21630);
nor U26223 (N_26223,N_21048,N_23548);
and U26224 (N_26224,N_23882,N_21807);
nor U26225 (N_26225,N_21000,N_22481);
xnor U26226 (N_26226,N_22042,N_21045);
nand U26227 (N_26227,N_23314,N_23966);
nor U26228 (N_26228,N_23552,N_21002);
xor U26229 (N_26229,N_22710,N_23333);
nand U26230 (N_26230,N_23352,N_23903);
xnor U26231 (N_26231,N_23743,N_22426);
or U26232 (N_26232,N_22948,N_22896);
xnor U26233 (N_26233,N_21321,N_23230);
or U26234 (N_26234,N_23399,N_23384);
or U26235 (N_26235,N_23178,N_21949);
or U26236 (N_26236,N_22952,N_23928);
and U26237 (N_26237,N_22270,N_22355);
or U26238 (N_26238,N_22172,N_21074);
nor U26239 (N_26239,N_21156,N_23955);
xnor U26240 (N_26240,N_23487,N_21228);
and U26241 (N_26241,N_23704,N_21012);
or U26242 (N_26242,N_23382,N_23174);
nor U26243 (N_26243,N_21953,N_21820);
and U26244 (N_26244,N_21727,N_21739);
xor U26245 (N_26245,N_23717,N_21306);
xor U26246 (N_26246,N_23225,N_22148);
or U26247 (N_26247,N_21851,N_23583);
and U26248 (N_26248,N_23371,N_22241);
nor U26249 (N_26249,N_23367,N_23125);
nand U26250 (N_26250,N_23550,N_21728);
xnor U26251 (N_26251,N_21636,N_22844);
xor U26252 (N_26252,N_21109,N_23478);
and U26253 (N_26253,N_22723,N_21755);
or U26254 (N_26254,N_21946,N_22883);
or U26255 (N_26255,N_23396,N_23423);
nor U26256 (N_26256,N_23919,N_23278);
and U26257 (N_26257,N_23382,N_22230);
xor U26258 (N_26258,N_23135,N_23814);
nor U26259 (N_26259,N_22032,N_21779);
or U26260 (N_26260,N_23767,N_22221);
nor U26261 (N_26261,N_22983,N_22560);
or U26262 (N_26262,N_23773,N_22820);
and U26263 (N_26263,N_22073,N_21951);
nor U26264 (N_26264,N_23663,N_22970);
xor U26265 (N_26265,N_21406,N_22491);
and U26266 (N_26266,N_21971,N_21923);
and U26267 (N_26267,N_22534,N_23037);
or U26268 (N_26268,N_23168,N_21911);
xnor U26269 (N_26269,N_23878,N_23901);
nand U26270 (N_26270,N_22816,N_22691);
nand U26271 (N_26271,N_21700,N_22090);
nor U26272 (N_26272,N_23155,N_21382);
or U26273 (N_26273,N_22492,N_23511);
or U26274 (N_26274,N_23842,N_23014);
or U26275 (N_26275,N_21438,N_22639);
nor U26276 (N_26276,N_22063,N_22383);
xnor U26277 (N_26277,N_22936,N_23256);
nor U26278 (N_26278,N_21178,N_22026);
xor U26279 (N_26279,N_23879,N_22117);
xor U26280 (N_26280,N_21345,N_23532);
and U26281 (N_26281,N_21221,N_21532);
and U26282 (N_26282,N_23718,N_21750);
nand U26283 (N_26283,N_22024,N_22869);
and U26284 (N_26284,N_22539,N_21602);
nand U26285 (N_26285,N_22036,N_23408);
and U26286 (N_26286,N_22041,N_23178);
nor U26287 (N_26287,N_22948,N_23395);
nor U26288 (N_26288,N_23452,N_22683);
or U26289 (N_26289,N_21754,N_21122);
nor U26290 (N_26290,N_21790,N_23033);
xnor U26291 (N_26291,N_22890,N_23066);
or U26292 (N_26292,N_21471,N_21045);
nand U26293 (N_26293,N_21580,N_22163);
and U26294 (N_26294,N_22416,N_23334);
nand U26295 (N_26295,N_23900,N_21364);
or U26296 (N_26296,N_21562,N_21572);
nand U26297 (N_26297,N_23824,N_22897);
and U26298 (N_26298,N_22723,N_21494);
and U26299 (N_26299,N_23480,N_21912);
and U26300 (N_26300,N_22745,N_23236);
and U26301 (N_26301,N_21868,N_21790);
or U26302 (N_26302,N_21259,N_22517);
nor U26303 (N_26303,N_21819,N_23553);
and U26304 (N_26304,N_23419,N_21188);
xor U26305 (N_26305,N_22720,N_23592);
or U26306 (N_26306,N_21048,N_23880);
xor U26307 (N_26307,N_23649,N_23134);
nand U26308 (N_26308,N_21697,N_23949);
nor U26309 (N_26309,N_22082,N_22502);
and U26310 (N_26310,N_21225,N_21647);
and U26311 (N_26311,N_21474,N_22951);
and U26312 (N_26312,N_21110,N_22360);
and U26313 (N_26313,N_21304,N_21005);
and U26314 (N_26314,N_21200,N_22942);
nor U26315 (N_26315,N_22405,N_21038);
and U26316 (N_26316,N_21427,N_23477);
nor U26317 (N_26317,N_22117,N_22305);
or U26318 (N_26318,N_21374,N_21834);
and U26319 (N_26319,N_21454,N_21389);
nand U26320 (N_26320,N_23671,N_21915);
nand U26321 (N_26321,N_21697,N_22915);
or U26322 (N_26322,N_21445,N_22453);
nand U26323 (N_26323,N_22285,N_22844);
nor U26324 (N_26324,N_23506,N_22957);
or U26325 (N_26325,N_22748,N_23596);
or U26326 (N_26326,N_23692,N_22494);
and U26327 (N_26327,N_22682,N_21049);
xor U26328 (N_26328,N_21774,N_23420);
and U26329 (N_26329,N_21957,N_21387);
and U26330 (N_26330,N_23743,N_22500);
nor U26331 (N_26331,N_22995,N_22670);
or U26332 (N_26332,N_23819,N_21022);
nor U26333 (N_26333,N_21794,N_22681);
and U26334 (N_26334,N_22194,N_23293);
xor U26335 (N_26335,N_22394,N_23355);
nand U26336 (N_26336,N_22399,N_21643);
nand U26337 (N_26337,N_21257,N_22386);
xnor U26338 (N_26338,N_23389,N_23500);
nand U26339 (N_26339,N_22333,N_22237);
and U26340 (N_26340,N_21848,N_21863);
and U26341 (N_26341,N_22724,N_23640);
xor U26342 (N_26342,N_22843,N_22301);
xor U26343 (N_26343,N_22302,N_23644);
and U26344 (N_26344,N_21404,N_23357);
nand U26345 (N_26345,N_23558,N_22135);
or U26346 (N_26346,N_22023,N_23128);
and U26347 (N_26347,N_21883,N_21389);
xor U26348 (N_26348,N_22365,N_23991);
or U26349 (N_26349,N_23977,N_21967);
and U26350 (N_26350,N_23358,N_21220);
and U26351 (N_26351,N_22709,N_21970);
xnor U26352 (N_26352,N_22752,N_22764);
xnor U26353 (N_26353,N_23226,N_23645);
or U26354 (N_26354,N_23955,N_22822);
xor U26355 (N_26355,N_22112,N_23840);
or U26356 (N_26356,N_23374,N_21648);
xor U26357 (N_26357,N_22660,N_23365);
or U26358 (N_26358,N_21830,N_23821);
or U26359 (N_26359,N_23937,N_22087);
and U26360 (N_26360,N_23688,N_23201);
nor U26361 (N_26361,N_21709,N_22488);
and U26362 (N_26362,N_22575,N_21010);
nand U26363 (N_26363,N_23721,N_21958);
xor U26364 (N_26364,N_22903,N_22322);
nor U26365 (N_26365,N_23252,N_23761);
nand U26366 (N_26366,N_21553,N_21784);
or U26367 (N_26367,N_21210,N_21527);
nand U26368 (N_26368,N_22061,N_22425);
nand U26369 (N_26369,N_21637,N_22879);
nand U26370 (N_26370,N_22610,N_23892);
xnor U26371 (N_26371,N_23601,N_21468);
or U26372 (N_26372,N_21151,N_21768);
and U26373 (N_26373,N_21341,N_21180);
or U26374 (N_26374,N_23838,N_21806);
and U26375 (N_26375,N_21762,N_22318);
nor U26376 (N_26376,N_21716,N_21428);
xor U26377 (N_26377,N_21262,N_23863);
and U26378 (N_26378,N_22489,N_22897);
nand U26379 (N_26379,N_22905,N_23292);
nand U26380 (N_26380,N_23034,N_23819);
or U26381 (N_26381,N_22849,N_23371);
and U26382 (N_26382,N_21843,N_23538);
nor U26383 (N_26383,N_21097,N_21628);
and U26384 (N_26384,N_22837,N_23560);
or U26385 (N_26385,N_22635,N_23690);
and U26386 (N_26386,N_23923,N_23932);
nor U26387 (N_26387,N_21545,N_22297);
or U26388 (N_26388,N_21779,N_21182);
and U26389 (N_26389,N_22074,N_23948);
or U26390 (N_26390,N_21240,N_22009);
and U26391 (N_26391,N_22282,N_21519);
nand U26392 (N_26392,N_21551,N_22161);
and U26393 (N_26393,N_23778,N_23074);
nor U26394 (N_26394,N_22974,N_22025);
xnor U26395 (N_26395,N_22654,N_22344);
nand U26396 (N_26396,N_21244,N_23896);
nand U26397 (N_26397,N_22493,N_23917);
and U26398 (N_26398,N_23891,N_21307);
nand U26399 (N_26399,N_23627,N_23518);
nand U26400 (N_26400,N_21902,N_22640);
xnor U26401 (N_26401,N_21012,N_21750);
xnor U26402 (N_26402,N_22574,N_22152);
nor U26403 (N_26403,N_21069,N_23685);
or U26404 (N_26404,N_23770,N_22034);
and U26405 (N_26405,N_22575,N_21736);
nor U26406 (N_26406,N_23814,N_22268);
nand U26407 (N_26407,N_23150,N_21510);
nand U26408 (N_26408,N_23028,N_23186);
and U26409 (N_26409,N_23494,N_23056);
xor U26410 (N_26410,N_21689,N_23363);
nand U26411 (N_26411,N_21040,N_21297);
nor U26412 (N_26412,N_21082,N_23947);
or U26413 (N_26413,N_23337,N_22887);
nor U26414 (N_26414,N_23597,N_22819);
xor U26415 (N_26415,N_22894,N_21247);
and U26416 (N_26416,N_21451,N_21112);
nand U26417 (N_26417,N_22785,N_22866);
nand U26418 (N_26418,N_22273,N_23443);
nor U26419 (N_26419,N_21798,N_22261);
or U26420 (N_26420,N_23852,N_21698);
and U26421 (N_26421,N_22059,N_22146);
and U26422 (N_26422,N_22347,N_21271);
or U26423 (N_26423,N_21182,N_22347);
or U26424 (N_26424,N_22713,N_22484);
nor U26425 (N_26425,N_23047,N_23032);
xnor U26426 (N_26426,N_21775,N_22570);
xnor U26427 (N_26427,N_21344,N_22464);
nor U26428 (N_26428,N_23121,N_22816);
nor U26429 (N_26429,N_21318,N_23087);
and U26430 (N_26430,N_23610,N_22172);
and U26431 (N_26431,N_21107,N_21494);
nor U26432 (N_26432,N_23947,N_23388);
nand U26433 (N_26433,N_21287,N_23534);
xor U26434 (N_26434,N_23138,N_21467);
nand U26435 (N_26435,N_22883,N_22689);
nor U26436 (N_26436,N_22162,N_22377);
or U26437 (N_26437,N_23685,N_23127);
or U26438 (N_26438,N_21159,N_21575);
nor U26439 (N_26439,N_21499,N_21293);
xnor U26440 (N_26440,N_22497,N_21874);
nand U26441 (N_26441,N_21123,N_23131);
nor U26442 (N_26442,N_21345,N_22382);
nand U26443 (N_26443,N_21969,N_23808);
and U26444 (N_26444,N_21786,N_22636);
and U26445 (N_26445,N_23585,N_22459);
nor U26446 (N_26446,N_23627,N_22058);
nand U26447 (N_26447,N_21206,N_22840);
nor U26448 (N_26448,N_21994,N_21980);
nor U26449 (N_26449,N_22212,N_21865);
nor U26450 (N_26450,N_22324,N_23095);
nor U26451 (N_26451,N_21874,N_21859);
xnor U26452 (N_26452,N_21281,N_22653);
nor U26453 (N_26453,N_22209,N_23752);
or U26454 (N_26454,N_22872,N_21206);
nand U26455 (N_26455,N_22538,N_22737);
and U26456 (N_26456,N_21437,N_21078);
and U26457 (N_26457,N_23330,N_23119);
and U26458 (N_26458,N_21149,N_23381);
xnor U26459 (N_26459,N_23813,N_22539);
or U26460 (N_26460,N_23666,N_22225);
or U26461 (N_26461,N_21191,N_21604);
or U26462 (N_26462,N_21930,N_22573);
and U26463 (N_26463,N_21346,N_23932);
xnor U26464 (N_26464,N_21231,N_21611);
nor U26465 (N_26465,N_23188,N_22154);
nor U26466 (N_26466,N_21668,N_21100);
and U26467 (N_26467,N_21133,N_23348);
nand U26468 (N_26468,N_22995,N_21733);
xnor U26469 (N_26469,N_21133,N_23457);
nand U26470 (N_26470,N_22146,N_22341);
nand U26471 (N_26471,N_23692,N_22075);
nand U26472 (N_26472,N_23819,N_21164);
nand U26473 (N_26473,N_21661,N_22073);
or U26474 (N_26474,N_21361,N_22915);
xor U26475 (N_26475,N_21926,N_21880);
xnor U26476 (N_26476,N_22055,N_23204);
or U26477 (N_26477,N_22009,N_22970);
xor U26478 (N_26478,N_21939,N_22631);
nand U26479 (N_26479,N_22179,N_21859);
and U26480 (N_26480,N_21795,N_23772);
nor U26481 (N_26481,N_23899,N_23107);
and U26482 (N_26482,N_22881,N_22684);
nor U26483 (N_26483,N_21605,N_23817);
or U26484 (N_26484,N_23055,N_23452);
nand U26485 (N_26485,N_23994,N_21671);
xnor U26486 (N_26486,N_21555,N_21836);
xor U26487 (N_26487,N_21730,N_23327);
nand U26488 (N_26488,N_21432,N_23026);
and U26489 (N_26489,N_23427,N_23824);
and U26490 (N_26490,N_22814,N_21327);
nand U26491 (N_26491,N_23281,N_22942);
and U26492 (N_26492,N_23581,N_22266);
and U26493 (N_26493,N_23692,N_21287);
and U26494 (N_26494,N_21978,N_22696);
nand U26495 (N_26495,N_22967,N_23921);
and U26496 (N_26496,N_21059,N_23896);
nor U26497 (N_26497,N_21782,N_23035);
xor U26498 (N_26498,N_22374,N_23218);
xor U26499 (N_26499,N_23905,N_23855);
or U26500 (N_26500,N_23601,N_21071);
or U26501 (N_26501,N_21107,N_22500);
xnor U26502 (N_26502,N_22054,N_22657);
nand U26503 (N_26503,N_21611,N_23146);
or U26504 (N_26504,N_21363,N_22695);
nor U26505 (N_26505,N_22961,N_22840);
nor U26506 (N_26506,N_23352,N_21926);
nand U26507 (N_26507,N_21942,N_23627);
nor U26508 (N_26508,N_23186,N_23190);
nand U26509 (N_26509,N_23731,N_21674);
and U26510 (N_26510,N_22357,N_21951);
nor U26511 (N_26511,N_21384,N_21004);
nand U26512 (N_26512,N_23588,N_21650);
nand U26513 (N_26513,N_23995,N_23891);
and U26514 (N_26514,N_21822,N_21064);
and U26515 (N_26515,N_21655,N_21214);
or U26516 (N_26516,N_21372,N_22849);
or U26517 (N_26517,N_22666,N_22587);
nand U26518 (N_26518,N_22760,N_21586);
and U26519 (N_26519,N_22568,N_23273);
and U26520 (N_26520,N_23439,N_23787);
or U26521 (N_26521,N_23548,N_21104);
xor U26522 (N_26522,N_23821,N_22175);
xnor U26523 (N_26523,N_22072,N_21319);
or U26524 (N_26524,N_23298,N_21041);
and U26525 (N_26525,N_22996,N_21082);
nand U26526 (N_26526,N_21688,N_21328);
xnor U26527 (N_26527,N_23109,N_22760);
nand U26528 (N_26528,N_23578,N_23520);
and U26529 (N_26529,N_21165,N_23732);
nor U26530 (N_26530,N_21651,N_22533);
nand U26531 (N_26531,N_23869,N_21468);
nor U26532 (N_26532,N_21545,N_23893);
or U26533 (N_26533,N_21128,N_22651);
xor U26534 (N_26534,N_23633,N_22370);
nor U26535 (N_26535,N_22925,N_21369);
nand U26536 (N_26536,N_23001,N_22886);
xor U26537 (N_26537,N_21614,N_21158);
nor U26538 (N_26538,N_22180,N_21449);
or U26539 (N_26539,N_21840,N_21066);
and U26540 (N_26540,N_23499,N_23222);
nor U26541 (N_26541,N_22204,N_23299);
nand U26542 (N_26542,N_21837,N_22157);
and U26543 (N_26543,N_23646,N_23497);
or U26544 (N_26544,N_22621,N_21966);
and U26545 (N_26545,N_22469,N_22447);
or U26546 (N_26546,N_22894,N_21342);
xor U26547 (N_26547,N_21979,N_21250);
xnor U26548 (N_26548,N_22867,N_23431);
xnor U26549 (N_26549,N_22641,N_23110);
or U26550 (N_26550,N_23703,N_21999);
nor U26551 (N_26551,N_22921,N_23095);
xor U26552 (N_26552,N_23632,N_23220);
and U26553 (N_26553,N_21519,N_23971);
and U26554 (N_26554,N_21031,N_21637);
nor U26555 (N_26555,N_21909,N_22597);
nand U26556 (N_26556,N_23908,N_22422);
and U26557 (N_26557,N_22804,N_22494);
and U26558 (N_26558,N_21185,N_21511);
xor U26559 (N_26559,N_23657,N_22534);
xor U26560 (N_26560,N_23396,N_22324);
and U26561 (N_26561,N_21209,N_21091);
xnor U26562 (N_26562,N_21404,N_21288);
or U26563 (N_26563,N_23545,N_22867);
xnor U26564 (N_26564,N_21097,N_23867);
xnor U26565 (N_26565,N_23663,N_21127);
and U26566 (N_26566,N_23274,N_22963);
nand U26567 (N_26567,N_22050,N_21227);
xor U26568 (N_26568,N_23777,N_22528);
nor U26569 (N_26569,N_22683,N_21449);
or U26570 (N_26570,N_21265,N_22716);
nor U26571 (N_26571,N_23033,N_23931);
and U26572 (N_26572,N_22896,N_21497);
or U26573 (N_26573,N_22455,N_22484);
and U26574 (N_26574,N_21370,N_23011);
or U26575 (N_26575,N_22687,N_22989);
nand U26576 (N_26576,N_21485,N_23248);
xor U26577 (N_26577,N_21938,N_21354);
nand U26578 (N_26578,N_22246,N_23113);
nand U26579 (N_26579,N_21791,N_23768);
nand U26580 (N_26580,N_21513,N_23702);
nor U26581 (N_26581,N_23125,N_22192);
and U26582 (N_26582,N_22871,N_23187);
nand U26583 (N_26583,N_23838,N_22166);
xor U26584 (N_26584,N_22658,N_23495);
nand U26585 (N_26585,N_22317,N_22015);
nand U26586 (N_26586,N_21576,N_23800);
xor U26587 (N_26587,N_23281,N_22201);
xnor U26588 (N_26588,N_22575,N_21229);
xnor U26589 (N_26589,N_22398,N_22585);
or U26590 (N_26590,N_23461,N_22632);
and U26591 (N_26591,N_22505,N_22491);
nand U26592 (N_26592,N_21859,N_22851);
and U26593 (N_26593,N_21604,N_22672);
nor U26594 (N_26594,N_21800,N_21955);
and U26595 (N_26595,N_21209,N_21584);
nor U26596 (N_26596,N_23896,N_22338);
nor U26597 (N_26597,N_23459,N_22694);
nor U26598 (N_26598,N_23357,N_23474);
nand U26599 (N_26599,N_23212,N_23037);
and U26600 (N_26600,N_23375,N_22470);
xor U26601 (N_26601,N_22545,N_22973);
nor U26602 (N_26602,N_23330,N_21609);
xor U26603 (N_26603,N_23309,N_22702);
xnor U26604 (N_26604,N_21806,N_22542);
and U26605 (N_26605,N_23260,N_23164);
nand U26606 (N_26606,N_23313,N_23271);
xor U26607 (N_26607,N_22780,N_21595);
xor U26608 (N_26608,N_23491,N_21639);
or U26609 (N_26609,N_23671,N_23923);
xnor U26610 (N_26610,N_22968,N_23415);
or U26611 (N_26611,N_22259,N_22986);
nand U26612 (N_26612,N_23596,N_22821);
and U26613 (N_26613,N_23764,N_21773);
nor U26614 (N_26614,N_21559,N_22608);
and U26615 (N_26615,N_21635,N_23041);
nand U26616 (N_26616,N_21151,N_22847);
nor U26617 (N_26617,N_23972,N_21606);
nor U26618 (N_26618,N_21863,N_23477);
and U26619 (N_26619,N_21791,N_21326);
and U26620 (N_26620,N_22418,N_22333);
xor U26621 (N_26621,N_21507,N_22285);
xnor U26622 (N_26622,N_22962,N_23856);
nor U26623 (N_26623,N_23517,N_23555);
and U26624 (N_26624,N_23507,N_23147);
nand U26625 (N_26625,N_23840,N_21651);
or U26626 (N_26626,N_23756,N_23449);
nor U26627 (N_26627,N_21417,N_22347);
xnor U26628 (N_26628,N_22053,N_23669);
or U26629 (N_26629,N_21030,N_21305);
xnor U26630 (N_26630,N_21983,N_21742);
nand U26631 (N_26631,N_21781,N_21143);
nor U26632 (N_26632,N_23907,N_23075);
and U26633 (N_26633,N_22705,N_21281);
or U26634 (N_26634,N_23857,N_23803);
xor U26635 (N_26635,N_21453,N_22659);
or U26636 (N_26636,N_21633,N_21843);
xnor U26637 (N_26637,N_23464,N_22348);
nand U26638 (N_26638,N_21464,N_21658);
xor U26639 (N_26639,N_21190,N_22230);
or U26640 (N_26640,N_21346,N_21621);
and U26641 (N_26641,N_22635,N_22730);
and U26642 (N_26642,N_21418,N_21264);
or U26643 (N_26643,N_22338,N_21401);
and U26644 (N_26644,N_21325,N_23611);
nor U26645 (N_26645,N_21893,N_23884);
nor U26646 (N_26646,N_22197,N_22730);
and U26647 (N_26647,N_21832,N_21513);
and U26648 (N_26648,N_22270,N_21965);
xor U26649 (N_26649,N_21808,N_23735);
nand U26650 (N_26650,N_21012,N_23437);
nor U26651 (N_26651,N_23710,N_22539);
and U26652 (N_26652,N_23871,N_23227);
nor U26653 (N_26653,N_21944,N_22826);
nand U26654 (N_26654,N_23788,N_22202);
and U26655 (N_26655,N_22372,N_22623);
nor U26656 (N_26656,N_21721,N_22331);
and U26657 (N_26657,N_23558,N_23471);
nand U26658 (N_26658,N_21695,N_22983);
xnor U26659 (N_26659,N_22984,N_22883);
and U26660 (N_26660,N_23879,N_21783);
or U26661 (N_26661,N_23587,N_21596);
xnor U26662 (N_26662,N_23167,N_23389);
or U26663 (N_26663,N_23156,N_22907);
and U26664 (N_26664,N_23261,N_22500);
or U26665 (N_26665,N_22127,N_23852);
xor U26666 (N_26666,N_21707,N_23119);
and U26667 (N_26667,N_22902,N_21482);
xor U26668 (N_26668,N_23403,N_21922);
nand U26669 (N_26669,N_21023,N_21603);
xnor U26670 (N_26670,N_22945,N_22311);
and U26671 (N_26671,N_23592,N_21555);
xor U26672 (N_26672,N_22467,N_21296);
or U26673 (N_26673,N_23611,N_22866);
nand U26674 (N_26674,N_23290,N_23368);
and U26675 (N_26675,N_21426,N_22985);
nand U26676 (N_26676,N_21252,N_22315);
nand U26677 (N_26677,N_22645,N_23540);
nand U26678 (N_26678,N_22666,N_22984);
and U26679 (N_26679,N_21044,N_22028);
nor U26680 (N_26680,N_21158,N_21190);
and U26681 (N_26681,N_21741,N_21235);
nand U26682 (N_26682,N_23752,N_23026);
nand U26683 (N_26683,N_23159,N_23415);
xnor U26684 (N_26684,N_22685,N_21609);
and U26685 (N_26685,N_23859,N_22519);
xnor U26686 (N_26686,N_23197,N_22601);
xor U26687 (N_26687,N_21105,N_22190);
and U26688 (N_26688,N_22071,N_22163);
nor U26689 (N_26689,N_21806,N_23694);
nor U26690 (N_26690,N_22413,N_21028);
or U26691 (N_26691,N_21495,N_23418);
or U26692 (N_26692,N_22438,N_21093);
nor U26693 (N_26693,N_22824,N_21966);
xor U26694 (N_26694,N_21046,N_22260);
nand U26695 (N_26695,N_22612,N_21571);
and U26696 (N_26696,N_23117,N_21393);
or U26697 (N_26697,N_22818,N_21119);
xor U26698 (N_26698,N_21454,N_22292);
xor U26699 (N_26699,N_22425,N_21806);
and U26700 (N_26700,N_22172,N_21704);
or U26701 (N_26701,N_21051,N_23625);
and U26702 (N_26702,N_22002,N_22906);
xnor U26703 (N_26703,N_21202,N_23522);
or U26704 (N_26704,N_22516,N_22826);
nand U26705 (N_26705,N_21884,N_22370);
xnor U26706 (N_26706,N_23033,N_23801);
and U26707 (N_26707,N_22554,N_22346);
or U26708 (N_26708,N_22802,N_23123);
nand U26709 (N_26709,N_23273,N_22875);
nand U26710 (N_26710,N_22299,N_22826);
nand U26711 (N_26711,N_23601,N_22446);
xor U26712 (N_26712,N_22400,N_23746);
nor U26713 (N_26713,N_22233,N_23886);
and U26714 (N_26714,N_22720,N_22337);
or U26715 (N_26715,N_23498,N_22978);
and U26716 (N_26716,N_23099,N_22706);
xor U26717 (N_26717,N_23999,N_22573);
nor U26718 (N_26718,N_22402,N_22927);
and U26719 (N_26719,N_23036,N_22110);
nand U26720 (N_26720,N_23698,N_23690);
xor U26721 (N_26721,N_23947,N_23769);
nor U26722 (N_26722,N_23786,N_22877);
xor U26723 (N_26723,N_23335,N_21526);
nand U26724 (N_26724,N_21081,N_21921);
xnor U26725 (N_26725,N_22821,N_22576);
and U26726 (N_26726,N_23741,N_23848);
xor U26727 (N_26727,N_21890,N_22326);
or U26728 (N_26728,N_23645,N_22234);
or U26729 (N_26729,N_23261,N_23897);
or U26730 (N_26730,N_23321,N_22743);
or U26731 (N_26731,N_23514,N_22511);
xnor U26732 (N_26732,N_21179,N_21595);
or U26733 (N_26733,N_22590,N_22718);
or U26734 (N_26734,N_21225,N_22286);
nand U26735 (N_26735,N_23396,N_21754);
and U26736 (N_26736,N_22748,N_23042);
or U26737 (N_26737,N_23959,N_21907);
xnor U26738 (N_26738,N_22360,N_21299);
and U26739 (N_26739,N_23748,N_21040);
nor U26740 (N_26740,N_22120,N_22291);
nor U26741 (N_26741,N_22924,N_21524);
nor U26742 (N_26742,N_21578,N_23412);
nand U26743 (N_26743,N_22851,N_21865);
xor U26744 (N_26744,N_21291,N_23011);
or U26745 (N_26745,N_23112,N_22034);
and U26746 (N_26746,N_21403,N_21770);
nand U26747 (N_26747,N_22851,N_23476);
nor U26748 (N_26748,N_23344,N_21634);
or U26749 (N_26749,N_22619,N_21496);
xor U26750 (N_26750,N_23217,N_23748);
or U26751 (N_26751,N_23876,N_22255);
or U26752 (N_26752,N_21136,N_22745);
or U26753 (N_26753,N_23288,N_21648);
or U26754 (N_26754,N_23774,N_23469);
nor U26755 (N_26755,N_23228,N_22922);
or U26756 (N_26756,N_21178,N_23371);
nand U26757 (N_26757,N_21206,N_22275);
and U26758 (N_26758,N_23470,N_23264);
xor U26759 (N_26759,N_23052,N_21683);
or U26760 (N_26760,N_23771,N_22149);
nand U26761 (N_26761,N_22607,N_21799);
xnor U26762 (N_26762,N_23065,N_22162);
and U26763 (N_26763,N_21832,N_22549);
nand U26764 (N_26764,N_23433,N_22646);
nand U26765 (N_26765,N_22625,N_21814);
nor U26766 (N_26766,N_23398,N_23597);
nor U26767 (N_26767,N_22911,N_23959);
nand U26768 (N_26768,N_21261,N_23954);
or U26769 (N_26769,N_23050,N_22792);
and U26770 (N_26770,N_23355,N_23112);
nor U26771 (N_26771,N_23705,N_22755);
nand U26772 (N_26772,N_22172,N_22794);
or U26773 (N_26773,N_21852,N_22809);
or U26774 (N_26774,N_22879,N_21389);
xnor U26775 (N_26775,N_22549,N_21633);
nor U26776 (N_26776,N_21605,N_22907);
xor U26777 (N_26777,N_22573,N_22380);
or U26778 (N_26778,N_23545,N_22142);
or U26779 (N_26779,N_22756,N_22585);
and U26780 (N_26780,N_23889,N_22772);
xnor U26781 (N_26781,N_23831,N_21126);
and U26782 (N_26782,N_22857,N_22689);
nor U26783 (N_26783,N_21915,N_22435);
or U26784 (N_26784,N_23122,N_22784);
or U26785 (N_26785,N_22106,N_23385);
xnor U26786 (N_26786,N_21887,N_23043);
or U26787 (N_26787,N_22847,N_23166);
xnor U26788 (N_26788,N_23913,N_23334);
nor U26789 (N_26789,N_22426,N_22862);
or U26790 (N_26790,N_23990,N_23883);
nor U26791 (N_26791,N_21572,N_23351);
and U26792 (N_26792,N_22248,N_23786);
nand U26793 (N_26793,N_22328,N_21021);
xor U26794 (N_26794,N_23666,N_23432);
and U26795 (N_26795,N_22945,N_22804);
nand U26796 (N_26796,N_22574,N_21310);
xnor U26797 (N_26797,N_23332,N_22654);
nand U26798 (N_26798,N_23876,N_22125);
nor U26799 (N_26799,N_21355,N_22255);
or U26800 (N_26800,N_21020,N_23960);
nand U26801 (N_26801,N_23475,N_23930);
nand U26802 (N_26802,N_22985,N_21393);
xnor U26803 (N_26803,N_23441,N_22379);
and U26804 (N_26804,N_22382,N_21261);
nand U26805 (N_26805,N_23077,N_23957);
or U26806 (N_26806,N_22590,N_22659);
xor U26807 (N_26807,N_21149,N_23770);
and U26808 (N_26808,N_21893,N_22232);
nor U26809 (N_26809,N_21198,N_23760);
nand U26810 (N_26810,N_21758,N_23146);
xor U26811 (N_26811,N_22725,N_23223);
nor U26812 (N_26812,N_23554,N_22926);
xnor U26813 (N_26813,N_21187,N_22209);
or U26814 (N_26814,N_21855,N_21350);
or U26815 (N_26815,N_23591,N_22807);
xor U26816 (N_26816,N_21176,N_23053);
xor U26817 (N_26817,N_21902,N_23419);
nand U26818 (N_26818,N_22096,N_23745);
nor U26819 (N_26819,N_23600,N_23574);
xor U26820 (N_26820,N_21853,N_23976);
nand U26821 (N_26821,N_21232,N_21864);
xor U26822 (N_26822,N_23700,N_23928);
nand U26823 (N_26823,N_22548,N_21687);
xnor U26824 (N_26824,N_22678,N_22426);
nand U26825 (N_26825,N_21476,N_23894);
nor U26826 (N_26826,N_23158,N_21610);
nand U26827 (N_26827,N_22311,N_21628);
or U26828 (N_26828,N_21137,N_23429);
xnor U26829 (N_26829,N_22059,N_22122);
or U26830 (N_26830,N_21344,N_23551);
and U26831 (N_26831,N_21089,N_23808);
xor U26832 (N_26832,N_21233,N_22463);
or U26833 (N_26833,N_21898,N_21992);
or U26834 (N_26834,N_22990,N_23572);
nand U26835 (N_26835,N_22983,N_23706);
and U26836 (N_26836,N_23973,N_23144);
nor U26837 (N_26837,N_23808,N_22963);
xnor U26838 (N_26838,N_23666,N_21455);
and U26839 (N_26839,N_21971,N_23300);
and U26840 (N_26840,N_23713,N_21734);
xnor U26841 (N_26841,N_23677,N_21352);
xnor U26842 (N_26842,N_23192,N_23147);
or U26843 (N_26843,N_21269,N_22116);
xor U26844 (N_26844,N_22073,N_21318);
and U26845 (N_26845,N_22674,N_23692);
nand U26846 (N_26846,N_23103,N_21403);
and U26847 (N_26847,N_21977,N_21219);
and U26848 (N_26848,N_23218,N_22160);
nand U26849 (N_26849,N_22079,N_21366);
and U26850 (N_26850,N_22630,N_23315);
nor U26851 (N_26851,N_22244,N_23860);
nor U26852 (N_26852,N_22629,N_21428);
xor U26853 (N_26853,N_23060,N_21470);
and U26854 (N_26854,N_22210,N_21151);
nor U26855 (N_26855,N_21479,N_22820);
nand U26856 (N_26856,N_22182,N_21215);
or U26857 (N_26857,N_21522,N_23704);
and U26858 (N_26858,N_22900,N_21193);
xor U26859 (N_26859,N_23638,N_23621);
nor U26860 (N_26860,N_21739,N_22481);
nand U26861 (N_26861,N_23249,N_23487);
nor U26862 (N_26862,N_21481,N_22960);
and U26863 (N_26863,N_23268,N_23745);
nand U26864 (N_26864,N_21166,N_21002);
or U26865 (N_26865,N_21988,N_23077);
and U26866 (N_26866,N_21395,N_22223);
or U26867 (N_26867,N_21647,N_23344);
xor U26868 (N_26868,N_22276,N_23221);
nor U26869 (N_26869,N_21351,N_22742);
and U26870 (N_26870,N_21729,N_23108);
nor U26871 (N_26871,N_22863,N_22467);
or U26872 (N_26872,N_23692,N_22771);
nor U26873 (N_26873,N_21379,N_21964);
xor U26874 (N_26874,N_22574,N_23961);
xnor U26875 (N_26875,N_23271,N_23113);
nor U26876 (N_26876,N_23113,N_23189);
or U26877 (N_26877,N_22753,N_21779);
and U26878 (N_26878,N_21394,N_22767);
or U26879 (N_26879,N_21017,N_21187);
xnor U26880 (N_26880,N_22817,N_23554);
nor U26881 (N_26881,N_23941,N_23917);
nand U26882 (N_26882,N_21956,N_21288);
nor U26883 (N_26883,N_22530,N_22665);
or U26884 (N_26884,N_23148,N_23245);
nand U26885 (N_26885,N_21937,N_22824);
or U26886 (N_26886,N_23201,N_23068);
or U26887 (N_26887,N_23572,N_21024);
xor U26888 (N_26888,N_23056,N_21408);
nand U26889 (N_26889,N_22597,N_21475);
or U26890 (N_26890,N_23886,N_23553);
xnor U26891 (N_26891,N_23433,N_22098);
or U26892 (N_26892,N_23270,N_21151);
nor U26893 (N_26893,N_22485,N_22203);
xor U26894 (N_26894,N_22216,N_23690);
and U26895 (N_26895,N_23076,N_22117);
or U26896 (N_26896,N_21512,N_22468);
or U26897 (N_26897,N_23102,N_23916);
or U26898 (N_26898,N_22432,N_21499);
nand U26899 (N_26899,N_22950,N_22881);
nand U26900 (N_26900,N_21965,N_22038);
xnor U26901 (N_26901,N_22915,N_21614);
nand U26902 (N_26902,N_22581,N_23170);
nand U26903 (N_26903,N_22819,N_22043);
nand U26904 (N_26904,N_22468,N_22296);
xnor U26905 (N_26905,N_23475,N_21590);
or U26906 (N_26906,N_22427,N_21204);
and U26907 (N_26907,N_23461,N_23055);
xnor U26908 (N_26908,N_23065,N_21664);
nor U26909 (N_26909,N_23791,N_21095);
or U26910 (N_26910,N_22536,N_21853);
nor U26911 (N_26911,N_23321,N_23519);
xnor U26912 (N_26912,N_23392,N_22430);
xor U26913 (N_26913,N_21556,N_21406);
and U26914 (N_26914,N_23660,N_23311);
and U26915 (N_26915,N_23815,N_21004);
xnor U26916 (N_26916,N_22787,N_22052);
nor U26917 (N_26917,N_22894,N_23622);
nand U26918 (N_26918,N_22984,N_21735);
and U26919 (N_26919,N_21462,N_23520);
and U26920 (N_26920,N_22498,N_21244);
nand U26921 (N_26921,N_23598,N_21919);
and U26922 (N_26922,N_21819,N_22739);
or U26923 (N_26923,N_22507,N_22312);
xnor U26924 (N_26924,N_21577,N_23509);
and U26925 (N_26925,N_22890,N_22264);
or U26926 (N_26926,N_23318,N_23481);
xnor U26927 (N_26927,N_21489,N_22656);
nor U26928 (N_26928,N_23946,N_21280);
and U26929 (N_26929,N_21855,N_22036);
and U26930 (N_26930,N_21086,N_22588);
or U26931 (N_26931,N_21887,N_23203);
nor U26932 (N_26932,N_23813,N_22291);
or U26933 (N_26933,N_21999,N_21167);
and U26934 (N_26934,N_22707,N_21054);
xnor U26935 (N_26935,N_21168,N_23555);
or U26936 (N_26936,N_22753,N_23101);
xor U26937 (N_26937,N_22541,N_21175);
and U26938 (N_26938,N_22810,N_23461);
xor U26939 (N_26939,N_21744,N_23200);
nand U26940 (N_26940,N_23193,N_21238);
nor U26941 (N_26941,N_22955,N_22714);
nor U26942 (N_26942,N_23030,N_21627);
and U26943 (N_26943,N_23263,N_22698);
xor U26944 (N_26944,N_21911,N_22032);
nor U26945 (N_26945,N_21178,N_23255);
nand U26946 (N_26946,N_23025,N_22424);
and U26947 (N_26947,N_22267,N_21879);
nand U26948 (N_26948,N_22645,N_22748);
nand U26949 (N_26949,N_22741,N_23573);
and U26950 (N_26950,N_22334,N_21652);
xor U26951 (N_26951,N_21011,N_21668);
and U26952 (N_26952,N_22908,N_22923);
nor U26953 (N_26953,N_22560,N_22699);
or U26954 (N_26954,N_22469,N_21657);
nand U26955 (N_26955,N_22703,N_22853);
xor U26956 (N_26956,N_23770,N_22777);
xnor U26957 (N_26957,N_23430,N_22737);
nor U26958 (N_26958,N_22517,N_23933);
or U26959 (N_26959,N_23125,N_22880);
or U26960 (N_26960,N_21711,N_22096);
and U26961 (N_26961,N_21084,N_23903);
and U26962 (N_26962,N_21664,N_23879);
nand U26963 (N_26963,N_23840,N_21164);
or U26964 (N_26964,N_21765,N_23376);
xor U26965 (N_26965,N_21510,N_23072);
and U26966 (N_26966,N_21474,N_22653);
and U26967 (N_26967,N_23172,N_22868);
nor U26968 (N_26968,N_22200,N_22491);
and U26969 (N_26969,N_23432,N_21965);
nor U26970 (N_26970,N_22691,N_21399);
nand U26971 (N_26971,N_23433,N_23357);
nor U26972 (N_26972,N_21493,N_23234);
or U26973 (N_26973,N_21679,N_22413);
and U26974 (N_26974,N_23030,N_22237);
and U26975 (N_26975,N_21881,N_23999);
nand U26976 (N_26976,N_22514,N_22590);
or U26977 (N_26977,N_21938,N_23939);
xnor U26978 (N_26978,N_23304,N_22944);
or U26979 (N_26979,N_22796,N_22558);
nor U26980 (N_26980,N_22181,N_21852);
or U26981 (N_26981,N_21648,N_23404);
or U26982 (N_26982,N_23260,N_22850);
and U26983 (N_26983,N_21582,N_22740);
xor U26984 (N_26984,N_21149,N_22116);
and U26985 (N_26985,N_23146,N_22611);
nor U26986 (N_26986,N_21013,N_23090);
xor U26987 (N_26987,N_23122,N_23583);
and U26988 (N_26988,N_21708,N_21716);
xor U26989 (N_26989,N_23681,N_23643);
nor U26990 (N_26990,N_23331,N_21691);
nand U26991 (N_26991,N_22003,N_21373);
and U26992 (N_26992,N_21362,N_22237);
and U26993 (N_26993,N_23283,N_23167);
or U26994 (N_26994,N_21812,N_21789);
or U26995 (N_26995,N_23224,N_21180);
xnor U26996 (N_26996,N_23114,N_22418);
and U26997 (N_26997,N_22567,N_23578);
xor U26998 (N_26998,N_21425,N_21476);
nand U26999 (N_26999,N_23053,N_21415);
xor U27000 (N_27000,N_26815,N_24908);
and U27001 (N_27001,N_26402,N_24421);
and U27002 (N_27002,N_26178,N_24382);
and U27003 (N_27003,N_26055,N_26959);
nor U27004 (N_27004,N_26445,N_25466);
and U27005 (N_27005,N_26390,N_25252);
and U27006 (N_27006,N_26406,N_25303);
nor U27007 (N_27007,N_24547,N_24504);
xor U27008 (N_27008,N_26191,N_25016);
nor U27009 (N_27009,N_24842,N_24361);
nand U27010 (N_27010,N_25921,N_24783);
nor U27011 (N_27011,N_25772,N_25004);
or U27012 (N_27012,N_24641,N_24832);
nand U27013 (N_27013,N_25984,N_24067);
nand U27014 (N_27014,N_26833,N_24410);
nor U27015 (N_27015,N_24173,N_26072);
or U27016 (N_27016,N_26995,N_25395);
xor U27017 (N_27017,N_24419,N_25915);
or U27018 (N_27018,N_24223,N_26373);
xnor U27019 (N_27019,N_24843,N_24627);
xor U27020 (N_27020,N_25100,N_25814);
xnor U27021 (N_27021,N_25073,N_24610);
nand U27022 (N_27022,N_24066,N_25233);
nor U27023 (N_27023,N_26693,N_25978);
or U27024 (N_27024,N_26532,N_24405);
xnor U27025 (N_27025,N_24513,N_26614);
and U27026 (N_27026,N_26737,N_26994);
nor U27027 (N_27027,N_26077,N_25549);
nor U27028 (N_27028,N_24986,N_25767);
nand U27029 (N_27029,N_26355,N_26325);
or U27030 (N_27030,N_26853,N_26930);
and U27031 (N_27031,N_24077,N_25131);
nand U27032 (N_27032,N_26269,N_25378);
or U27033 (N_27033,N_26058,N_24852);
nand U27034 (N_27034,N_26050,N_24861);
nor U27035 (N_27035,N_25821,N_24501);
xnor U27036 (N_27036,N_24993,N_26452);
or U27037 (N_27037,N_26159,N_25946);
xor U27038 (N_27038,N_24771,N_25989);
nor U27039 (N_27039,N_26721,N_24640);
and U27040 (N_27040,N_25660,N_25526);
or U27041 (N_27041,N_26429,N_26579);
and U27042 (N_27042,N_24424,N_24830);
and U27043 (N_27043,N_26059,N_25867);
nand U27044 (N_27044,N_26214,N_25026);
and U27045 (N_27045,N_24037,N_25977);
or U27046 (N_27046,N_24375,N_26642);
xor U27047 (N_27047,N_24158,N_25334);
nand U27048 (N_27048,N_26265,N_26589);
nand U27049 (N_27049,N_26510,N_26009);
nor U27050 (N_27050,N_26447,N_25994);
xnor U27051 (N_27051,N_26089,N_24202);
nand U27052 (N_27052,N_24151,N_24990);
xor U27053 (N_27053,N_24427,N_26436);
xnor U27054 (N_27054,N_26256,N_26507);
xnor U27055 (N_27055,N_25329,N_24270);
xor U27056 (N_27056,N_24819,N_24124);
or U27057 (N_27057,N_24761,N_24072);
nand U27058 (N_27058,N_25158,N_26806);
nand U27059 (N_27059,N_25588,N_25700);
nand U27060 (N_27060,N_24668,N_26057);
nand U27061 (N_27061,N_25044,N_26034);
and U27062 (N_27062,N_25823,N_26268);
xnor U27063 (N_27063,N_24715,N_25121);
nor U27064 (N_27064,N_25935,N_25666);
xor U27065 (N_27065,N_24695,N_24679);
or U27066 (N_27066,N_25902,N_26972);
and U27067 (N_27067,N_25434,N_24490);
xnor U27068 (N_27068,N_26914,N_26968);
nand U27069 (N_27069,N_25524,N_25631);
nand U27070 (N_27070,N_24444,N_26011);
and U27071 (N_27071,N_24549,N_26673);
xor U27072 (N_27072,N_26996,N_25920);
and U27073 (N_27073,N_24534,N_26468);
nand U27074 (N_27074,N_26430,N_25725);
nor U27075 (N_27075,N_25277,N_25117);
nand U27076 (N_27076,N_26226,N_26490);
xnor U27077 (N_27077,N_25435,N_24170);
or U27078 (N_27078,N_26871,N_25231);
nor U27079 (N_27079,N_25555,N_26580);
and U27080 (N_27080,N_25265,N_26529);
xnor U27081 (N_27081,N_24972,N_24279);
or U27082 (N_27082,N_24690,N_24566);
xor U27083 (N_27083,N_26215,N_24731);
and U27084 (N_27084,N_25288,N_26915);
xor U27085 (N_27085,N_24409,N_24807);
or U27086 (N_27086,N_26030,N_26841);
nand U27087 (N_27087,N_24229,N_26878);
or U27088 (N_27088,N_24459,N_26453);
or U27089 (N_27089,N_26470,N_24907);
or U27090 (N_27090,N_25143,N_26320);
or U27091 (N_27091,N_26736,N_25890);
nor U27092 (N_27092,N_24743,N_25284);
nand U27093 (N_27093,N_24336,N_25896);
nor U27094 (N_27094,N_24138,N_25177);
or U27095 (N_27095,N_24214,N_24137);
nor U27096 (N_27096,N_25722,N_25628);
or U27097 (N_27097,N_24120,N_25748);
or U27098 (N_27098,N_25719,N_24787);
xor U27099 (N_27099,N_26924,N_26019);
nor U27100 (N_27100,N_25640,N_24484);
nor U27101 (N_27101,N_25908,N_25803);
or U27102 (N_27102,N_26258,N_24928);
and U27103 (N_27103,N_24153,N_26887);
or U27104 (N_27104,N_25112,N_24989);
nand U27105 (N_27105,N_25707,N_24445);
and U27106 (N_27106,N_25626,N_24630);
and U27107 (N_27107,N_25140,N_24727);
nor U27108 (N_27108,N_26640,N_24806);
or U27109 (N_27109,N_24789,N_26442);
nand U27110 (N_27110,N_26259,N_24376);
xor U27111 (N_27111,N_25769,N_25695);
nand U27112 (N_27112,N_24328,N_26353);
nor U27113 (N_27113,N_25097,N_26094);
xnor U27114 (N_27114,N_26318,N_25534);
nor U27115 (N_27115,N_25105,N_26230);
xor U27116 (N_27116,N_26333,N_26829);
or U27117 (N_27117,N_26465,N_25697);
and U27118 (N_27118,N_25339,N_24612);
xor U27119 (N_27119,N_26978,N_25496);
and U27120 (N_27120,N_24091,N_24048);
or U27121 (N_27121,N_25852,N_26377);
xor U27122 (N_27122,N_26300,N_24519);
and U27123 (N_27123,N_24694,N_26856);
or U27124 (N_27124,N_26649,N_25290);
or U27125 (N_27125,N_24291,N_26932);
nor U27126 (N_27126,N_26903,N_24167);
nor U27127 (N_27127,N_24890,N_26337);
or U27128 (N_27128,N_24582,N_26699);
and U27129 (N_27129,N_25881,N_26220);
and U27130 (N_27130,N_24236,N_25703);
nor U27131 (N_27131,N_24043,N_26477);
nand U27132 (N_27132,N_24538,N_26415);
xor U27133 (N_27133,N_24942,N_26905);
xnor U27134 (N_27134,N_25945,N_26124);
and U27135 (N_27135,N_25951,N_24093);
or U27136 (N_27136,N_26204,N_24882);
or U27137 (N_27137,N_24381,N_24929);
nor U27138 (N_27138,N_26123,N_26933);
or U27139 (N_27139,N_25853,N_24316);
or U27140 (N_27140,N_24415,N_25059);
nand U27141 (N_27141,N_25381,N_24536);
nand U27142 (N_27142,N_26264,N_26963);
xor U27143 (N_27143,N_25705,N_25127);
nor U27144 (N_27144,N_26150,N_25924);
nor U27145 (N_27145,N_24065,N_25879);
and U27146 (N_27146,N_26691,N_26462);
nand U27147 (N_27147,N_25980,N_26586);
or U27148 (N_27148,N_24275,N_25027);
nor U27149 (N_27149,N_26745,N_25261);
xnor U27150 (N_27150,N_26083,N_24190);
nand U27151 (N_27151,N_24062,N_26020);
or U27152 (N_27152,N_26970,N_26166);
nand U27153 (N_27153,N_26189,N_25726);
and U27154 (N_27154,N_26664,N_25576);
and U27155 (N_27155,N_26304,N_26350);
nor U27156 (N_27156,N_24286,N_26503);
and U27157 (N_27157,N_24898,N_25355);
xor U27158 (N_27158,N_24313,N_26066);
or U27159 (N_27159,N_25469,N_24924);
nand U27160 (N_27160,N_25540,N_26926);
nor U27161 (N_27161,N_24324,N_24385);
nand U27162 (N_27162,N_24775,N_26308);
and U27163 (N_27163,N_24985,N_24309);
nand U27164 (N_27164,N_26403,N_26454);
nand U27165 (N_27165,N_25262,N_26138);
nand U27166 (N_27166,N_26522,N_25036);
and U27167 (N_27167,N_25562,N_24562);
nand U27168 (N_27168,N_24499,N_25246);
nand U27169 (N_27169,N_26207,N_24212);
or U27170 (N_27170,N_24334,N_25641);
nor U27171 (N_27171,N_26935,N_24474);
or U27172 (N_27172,N_24117,N_24374);
nand U27173 (N_27173,N_25632,N_26735);
xor U27174 (N_27174,N_24317,N_25028);
nor U27175 (N_27175,N_25253,N_26494);
nand U27176 (N_27176,N_24892,N_25436);
xor U27177 (N_27177,N_26061,N_25239);
nor U27178 (N_27178,N_24970,N_26266);
xor U27179 (N_27179,N_24025,N_26224);
xnor U27180 (N_27180,N_26449,N_26272);
nor U27181 (N_27181,N_24577,N_26969);
nor U27182 (N_27182,N_24874,N_25472);
or U27183 (N_27183,N_25001,N_26956);
or U27184 (N_27184,N_25802,N_26511);
or U27185 (N_27185,N_26276,N_25675);
nor U27186 (N_27186,N_26165,N_24941);
xor U27187 (N_27187,N_25900,N_25831);
xnor U27188 (N_27188,N_25053,N_26395);
xor U27189 (N_27189,N_26530,N_24056);
nor U27190 (N_27190,N_25851,N_26385);
xnor U27191 (N_27191,N_25179,N_24156);
and U27192 (N_27192,N_25024,N_25521);
or U27193 (N_27193,N_24607,N_25054);
nor U27194 (N_27194,N_26378,N_25296);
and U27195 (N_27195,N_25522,N_25591);
nor U27196 (N_27196,N_24647,N_25670);
or U27197 (N_27197,N_25464,N_24226);
or U27198 (N_27198,N_26612,N_24732);
and U27199 (N_27199,N_25859,N_24044);
and U27200 (N_27200,N_24526,N_26170);
and U27201 (N_27201,N_24425,N_24502);
and U27202 (N_27202,N_26033,N_25219);
nor U27203 (N_27203,N_25126,N_25471);
nand U27204 (N_27204,N_26407,N_26200);
nand U27205 (N_27205,N_24643,N_24493);
or U27206 (N_27206,N_24981,N_24447);
nor U27207 (N_27207,N_26659,N_26604);
or U27208 (N_27208,N_25518,N_25332);
nor U27209 (N_27209,N_26154,N_24872);
nand U27210 (N_27210,N_24003,N_25553);
or U27211 (N_27211,N_25204,N_25067);
nor U27212 (N_27212,N_26027,N_25954);
or U27213 (N_27213,N_25468,N_26891);
xnor U27214 (N_27214,N_24636,N_24656);
or U27215 (N_27215,N_26720,N_24146);
xor U27216 (N_27216,N_25160,N_24050);
and U27217 (N_27217,N_25556,N_26847);
or U27218 (N_27218,N_25167,N_25183);
xnor U27219 (N_27219,N_24542,N_26032);
and U27220 (N_27220,N_24329,N_26596);
xor U27221 (N_27221,N_24840,N_24758);
nor U27222 (N_27222,N_24207,N_25446);
and U27223 (N_27223,N_26098,N_26424);
nand U27224 (N_27224,N_25706,N_26518);
nor U27225 (N_27225,N_26360,N_25035);
nand U27226 (N_27226,N_24118,N_25130);
xnor U27227 (N_27227,N_25282,N_26791);
xor U27228 (N_27228,N_25586,N_25693);
nand U27229 (N_27229,N_25955,N_24645);
xnor U27230 (N_27230,N_26456,N_25625);
xor U27231 (N_27231,N_24263,N_25872);
nor U27232 (N_27232,N_26158,N_26816);
nand U27233 (N_27233,N_26730,N_24561);
nand U27234 (N_27234,N_26169,N_26792);
xnor U27235 (N_27235,N_24744,N_26684);
nor U27236 (N_27236,N_24491,N_25639);
xnor U27237 (N_27237,N_26760,N_25255);
xor U27238 (N_27238,N_26605,N_25884);
xnor U27239 (N_27239,N_25194,N_25453);
or U27240 (N_27240,N_24274,N_24090);
and U27241 (N_27241,N_26879,N_25101);
or U27242 (N_27242,N_24488,N_25215);
xor U27243 (N_27243,N_26597,N_24088);
nand U27244 (N_27244,N_26814,N_25597);
xor U27245 (N_27245,N_25477,N_24185);
xnor U27246 (N_27246,N_26499,N_26515);
or U27247 (N_27247,N_24299,N_24049);
xnor U27248 (N_27248,N_26203,N_25883);
xnor U27249 (N_27249,N_26989,N_24398);
nand U27250 (N_27250,N_24475,N_25322);
nand U27251 (N_27251,N_25279,N_25025);
nor U27252 (N_27252,N_25806,N_25487);
and U27253 (N_27253,N_26393,N_24133);
xnor U27254 (N_27254,N_24089,N_26912);
nand U27255 (N_27255,N_24883,N_25895);
or U27256 (N_27256,N_26602,N_26495);
and U27257 (N_27257,N_25531,N_26283);
nand U27258 (N_27258,N_25248,N_25444);
and U27259 (N_27259,N_26750,N_24835);
xnor U27260 (N_27260,N_25981,N_24958);
nand U27261 (N_27261,N_26184,N_24633);
xor U27262 (N_27262,N_26650,N_24916);
nand U27263 (N_27263,N_25078,N_25825);
nand U27264 (N_27264,N_24457,N_25629);
xor U27265 (N_27265,N_24805,N_25889);
and U27266 (N_27266,N_24076,N_25386);
or U27267 (N_27267,N_24293,N_26361);
nand U27268 (N_27268,N_26143,N_25120);
xor U27269 (N_27269,N_26942,N_25974);
and U27270 (N_27270,N_25002,N_25805);
nor U27271 (N_27271,N_26267,N_24005);
or U27272 (N_27272,N_24116,N_24403);
nor U27273 (N_27273,N_25321,N_25537);
or U27274 (N_27274,N_24736,N_26014);
and U27275 (N_27275,N_25384,N_26434);
nor U27276 (N_27276,N_24943,N_25571);
xor U27277 (N_27277,N_26139,N_25554);
xnor U27278 (N_27278,N_24967,N_25864);
and U27279 (N_27279,N_24106,N_24784);
nor U27280 (N_27280,N_26254,N_25849);
or U27281 (N_27281,N_26967,N_25478);
nor U27282 (N_27282,N_24754,N_24128);
nand U27283 (N_27283,N_25929,N_24792);
and U27284 (N_27284,N_26389,N_26307);
and U27285 (N_27285,N_24677,N_25756);
nand U27286 (N_27286,N_25958,N_24085);
nand U27287 (N_27287,N_26493,N_25608);
xnor U27288 (N_27288,N_25405,N_26326);
xnor U27289 (N_27289,N_25865,N_26306);
xnor U27290 (N_27290,N_25266,N_26413);
nor U27291 (N_27291,N_25501,N_26433);
xnor U27292 (N_27292,N_24624,N_26686);
nand U27293 (N_27293,N_25732,N_26080);
or U27294 (N_27294,N_24567,N_24438);
or U27295 (N_27295,N_25736,N_25147);
nand U27296 (N_27296,N_26412,N_26130);
and U27297 (N_27297,N_24436,N_26846);
nand U27298 (N_27298,N_26976,N_26576);
nand U27299 (N_27299,N_24543,N_26992);
nand U27300 (N_27300,N_25839,N_24945);
and U27301 (N_27301,N_24682,N_24686);
nand U27302 (N_27302,N_25558,N_25439);
xnor U27303 (N_27303,N_25565,N_25846);
xnor U27304 (N_27304,N_25727,N_26957);
and U27305 (N_27305,N_24494,N_26349);
or U27306 (N_27306,N_26991,N_25717);
nor U27307 (N_27307,N_24255,N_24673);
xnor U27308 (N_27308,N_24234,N_24026);
or U27309 (N_27309,N_25430,N_24082);
or U27310 (N_27310,N_24745,N_25187);
nand U27311 (N_27311,N_24331,N_25835);
xor U27312 (N_27312,N_26253,N_26446);
xnor U27313 (N_27313,N_26091,N_24505);
xor U27314 (N_27314,N_25375,N_25207);
nor U27315 (N_27315,N_25270,N_25647);
and U27316 (N_27316,N_26799,N_25699);
and U27317 (N_27317,N_26983,N_25595);
xnor U27318 (N_27318,N_24795,N_25111);
xor U27319 (N_27319,N_25379,N_24179);
and U27320 (N_27320,N_24858,N_25574);
xnor U27321 (N_27321,N_25794,N_25728);
or U27322 (N_27322,N_25129,N_24777);
and U27323 (N_27323,N_26194,N_25903);
and U27324 (N_27324,N_25635,N_24480);
nand U27325 (N_27325,N_26397,N_25858);
nand U27326 (N_27326,N_25615,N_24407);
and U27327 (N_27327,N_24836,N_26336);
nand U27328 (N_27328,N_24952,N_24800);
or U27329 (N_27329,N_24455,N_26486);
nand U27330 (N_27330,N_26322,N_24834);
and U27331 (N_27331,N_24838,N_25516);
nor U27332 (N_27332,N_26243,N_24804);
and U27333 (N_27333,N_25930,N_26874);
and U27334 (N_27334,N_26862,N_26482);
nor U27335 (N_27335,N_24621,N_25603);
xnor U27336 (N_27336,N_25502,N_24058);
nor U27337 (N_27337,N_26624,N_24318);
xor U27338 (N_27338,N_26504,N_24495);
and U27339 (N_27339,N_24140,N_26718);
or U27340 (N_27340,N_24487,N_25003);
nand U27341 (N_27341,N_24816,N_25015);
and U27342 (N_27342,N_26180,N_26525);
or U27343 (N_27343,N_24984,N_26764);
nor U27344 (N_27344,N_26990,N_26783);
nand U27345 (N_27345,N_24696,N_24098);
xnor U27346 (N_27346,N_26384,N_24905);
xor U27347 (N_27347,N_25861,N_25039);
or U27348 (N_27348,N_25085,N_25891);
nand U27349 (N_27349,N_25776,N_26108);
nor U27350 (N_27350,N_26671,N_24934);
nand U27351 (N_27351,N_26554,N_26723);
or U27352 (N_27352,N_26105,N_25901);
xnor U27353 (N_27353,N_24629,N_24864);
nand U27354 (N_27354,N_24036,N_26010);
nand U27355 (N_27355,N_25730,N_25402);
or U27356 (N_27356,N_24397,N_25820);
xnor U27357 (N_27357,N_25353,N_25933);
and U27358 (N_27358,N_24648,N_25198);
and U27359 (N_27359,N_24352,N_25517);
nor U27360 (N_27360,N_26633,N_26752);
or U27361 (N_27361,N_25503,N_26257);
nor U27362 (N_27362,N_26046,N_26151);
and U27363 (N_27363,N_26068,N_24119);
nand U27364 (N_27364,N_26364,N_25871);
xnor U27365 (N_27365,N_24593,N_26104);
nand U27366 (N_27366,N_26177,N_25245);
nand U27367 (N_27367,N_25673,N_24420);
and U27368 (N_27368,N_26873,N_24471);
xor U27369 (N_27369,N_25461,N_26324);
and U27370 (N_27370,N_26084,N_26206);
and U27371 (N_27371,N_26892,N_26086);
nor U27372 (N_27372,N_24739,N_26354);
xor U27373 (N_27373,N_26164,N_26796);
xnor U27374 (N_27374,N_24897,N_25426);
xnor U27375 (N_27375,N_26509,N_25870);
xor U27376 (N_27376,N_25564,N_24974);
and U27377 (N_27377,N_24276,N_26840);
and U27378 (N_27378,N_25991,N_24553);
nor U27379 (N_27379,N_26909,N_26260);
xor U27380 (N_27380,N_25297,N_26202);
nor U27381 (N_27381,N_24772,N_25512);
xor U27382 (N_27382,N_25287,N_24839);
xor U27383 (N_27383,N_24671,N_24321);
nor U27384 (N_27384,N_26458,N_25021);
nor U27385 (N_27385,N_24107,N_26332);
xnor U27386 (N_27386,N_25237,N_26524);
nor U27387 (N_27387,N_26688,N_25792);
and U27388 (N_27388,N_25046,N_26097);
nand U27389 (N_27389,N_26818,N_24400);
and U27390 (N_27390,N_26753,N_25789);
nand U27391 (N_27391,N_26101,N_25197);
and U27392 (N_27392,N_26843,N_26450);
or U27393 (N_27393,N_24497,N_24540);
nand U27394 (N_27394,N_24155,N_25493);
xnor U27395 (N_27395,N_26656,N_24886);
or U27396 (N_27396,N_25013,N_24717);
xor U27397 (N_27397,N_26645,N_24139);
and U27398 (N_27398,N_26109,N_25498);
nor U27399 (N_27399,N_24295,N_26621);
or U27400 (N_27400,N_26979,N_26535);
nor U27401 (N_27401,N_25696,N_24130);
nor U27402 (N_27402,N_24681,N_25301);
or U27403 (N_27403,N_25927,N_24027);
xor U27404 (N_27404,N_25467,N_26677);
and U27405 (N_27405,N_24971,N_25267);
xnor U27406 (N_27406,N_24416,N_25552);
or U27407 (N_27407,N_26174,N_26961);
and U27408 (N_27408,N_26145,N_25342);
and U27409 (N_27409,N_25932,N_26759);
or U27410 (N_27410,N_25391,N_26323);
xnor U27411 (N_27411,N_25153,N_24238);
and U27412 (N_27412,N_26287,N_25030);
nor U27413 (N_27413,N_26279,N_24844);
nor U27414 (N_27414,N_25637,N_26362);
xnor U27415 (N_27415,N_26794,N_25109);
or U27416 (N_27416,N_24517,N_24466);
and U27417 (N_27417,N_26371,N_26122);
or U27418 (N_27418,N_26769,N_24654);
and U27419 (N_27419,N_24667,N_26551);
xor U27420 (N_27420,N_26618,N_26772);
and U27421 (N_27421,N_25470,N_25985);
xor U27422 (N_27422,N_25777,N_25314);
and U27423 (N_27423,N_24399,N_26830);
nand U27424 (N_27424,N_24964,N_24877);
xor U27425 (N_27425,N_25746,N_26028);
nand U27426 (N_27426,N_25382,N_24033);
and U27427 (N_27427,N_24370,N_24541);
xnor U27428 (N_27428,N_24454,N_26566);
nor U27429 (N_27429,N_25096,N_25917);
nand U27430 (N_27430,N_24362,N_26013);
nand U27431 (N_27431,N_26584,N_25043);
xor U27432 (N_27432,N_25559,N_25302);
and U27433 (N_27433,N_26026,N_24559);
nor U27434 (N_27434,N_26958,N_24194);
nand U27435 (N_27435,N_24569,N_25684);
xor U27436 (N_27436,N_24856,N_25286);
and U27437 (N_27437,N_25715,N_24810);
xor U27438 (N_27438,N_25094,N_25492);
nor U27439 (N_27439,N_24575,N_25420);
and U27440 (N_27440,N_26103,N_24023);
or U27441 (N_27441,N_25336,N_25711);
and U27442 (N_27442,N_24653,N_25357);
nor U27443 (N_27443,N_25863,N_26301);
nor U27444 (N_27444,N_25473,N_24665);
and U27445 (N_27445,N_25782,N_25623);
nand U27446 (N_27446,N_26953,N_24112);
nor U27447 (N_27447,N_24670,N_24253);
or U27448 (N_27448,N_24393,N_25387);
nand U27449 (N_27449,N_24531,N_24652);
or U27450 (N_27450,N_25091,N_26687);
xnor U27451 (N_27451,N_25691,N_25412);
xnor U27452 (N_27452,N_26526,N_25504);
and U27453 (N_27453,N_25940,N_24862);
xor U27454 (N_27454,N_25616,N_26826);
nor U27455 (N_27455,N_26666,N_25235);
or U27456 (N_27456,N_26400,N_25605);
or U27457 (N_27457,N_26100,N_25860);
and U27458 (N_27458,N_25123,N_25643);
or U27459 (N_27459,N_24552,N_24760);
nor U27460 (N_27460,N_25541,N_25681);
nor U27461 (N_27461,N_26727,N_25240);
or U27462 (N_27462,N_25589,N_24738);
and U27463 (N_27463,N_26590,N_26093);
nand U27464 (N_27464,N_26619,N_26156);
and U27465 (N_27465,N_26133,N_24045);
xnor U27466 (N_27466,N_24478,N_26860);
or U27467 (N_27467,N_26778,N_26401);
and U27468 (N_27468,N_26857,N_24750);
xnor U27469 (N_27469,N_24014,N_24606);
and U27470 (N_27470,N_25232,N_24010);
and U27471 (N_27471,N_25442,N_24512);
and U27472 (N_27472,N_26366,N_25486);
and U27473 (N_27473,N_24735,N_26756);
nand U27474 (N_27474,N_26627,N_25850);
xnor U27475 (N_27475,N_24154,N_26635);
or U27476 (N_27476,N_25780,N_24709);
and U27477 (N_27477,N_24599,N_26817);
nand U27478 (N_27478,N_25753,N_26941);
nand U27479 (N_27479,N_25830,N_25328);
xnor U27480 (N_27480,N_24380,N_24973);
or U27481 (N_27481,N_25259,N_24147);
xor U27482 (N_27482,N_25403,N_24343);
xor U27483 (N_27483,N_24017,N_26147);
nand U27484 (N_27484,N_24506,N_24312);
xnor U27485 (N_27485,N_26069,N_25203);
xor U27486 (N_27486,N_24503,N_25743);
nor U27487 (N_27487,N_25022,N_24729);
nand U27488 (N_27488,N_24217,N_26728);
nor U27489 (N_27489,N_25309,N_24662);
and U27490 (N_27490,N_25058,N_24047);
or U27491 (N_27491,N_25809,N_24605);
nand U27492 (N_27492,N_25366,N_26114);
and U27493 (N_27493,N_26466,N_24460);
nand U27494 (N_27494,N_25304,N_25737);
nor U27495 (N_27495,N_24723,N_26461);
and U27496 (N_27496,N_24183,N_25319);
xor U27497 (N_27497,N_24741,N_26487);
nor U27498 (N_27498,N_25271,N_26742);
nor U27499 (N_27499,N_26497,N_25450);
and U27500 (N_27500,N_25546,N_24558);
and U27501 (N_27501,N_25936,N_24189);
xor U27502 (N_27502,N_26303,N_26694);
xnor U27503 (N_27503,N_24991,N_26346);
and U27504 (N_27504,N_26417,N_24000);
nand U27505 (N_27505,N_24518,N_25351);
xor U27506 (N_27506,N_24383,N_24837);
nor U27507 (N_27507,N_26861,N_26911);
nand U27508 (N_27508,N_26965,N_24651);
and U27509 (N_27509,N_24232,N_25414);
nand U27510 (N_27510,N_26228,N_24123);
nand U27511 (N_27511,N_25338,N_25723);
or U27512 (N_27512,N_24351,N_24193);
and U27513 (N_27513,N_24177,N_25771);
nor U27514 (N_27514,N_25424,N_25333);
nor U27515 (N_27515,N_25084,N_26683);
nor U27516 (N_27516,N_26388,N_26929);
xor U27517 (N_27517,N_24759,N_24675);
nor U27518 (N_27518,N_24100,N_25306);
or U27519 (N_27519,N_24191,N_26620);
or U27520 (N_27520,N_26782,N_25071);
or U27521 (N_27521,N_26679,N_25886);
and U27522 (N_27522,N_25390,N_24713);
nand U27523 (N_27523,N_26227,N_26375);
nor U27524 (N_27524,N_25761,N_25652);
and U27525 (N_27525,N_26896,N_26544);
nor U27526 (N_27526,N_25506,N_24615);
and U27527 (N_27527,N_24162,N_26638);
nand U27528 (N_27528,N_26971,N_26644);
nand U27529 (N_27529,N_26917,N_24379);
and U27530 (N_27530,N_24319,N_24585);
and U27531 (N_27531,N_26129,N_24031);
and U27532 (N_27532,N_26351,N_26585);
nor U27533 (N_27533,N_25327,N_25976);
xor U27534 (N_27534,N_25720,N_25077);
and U27535 (N_27535,N_26459,N_24440);
nand U27536 (N_27536,N_24134,N_25755);
and U27537 (N_27537,N_24707,N_25364);
or U27538 (N_27538,N_24465,N_24963);
and U27539 (N_27539,N_24355,N_26327);
nand U27540 (N_27540,N_25817,N_26421);
xnor U27541 (N_27541,N_26328,N_26973);
nand U27542 (N_27542,N_26155,N_25050);
or U27543 (N_27543,N_25686,N_24184);
nand U27544 (N_27544,N_25312,N_26601);
or U27545 (N_27545,N_26670,N_26148);
nand U27546 (N_27546,N_24809,N_26457);
and U27547 (N_27547,N_25729,N_25257);
nor U27548 (N_27548,N_26088,N_24462);
and U27549 (N_27549,N_24638,N_24260);
nor U27550 (N_27550,N_24142,N_25218);
nand U27551 (N_27551,N_25086,N_25797);
nor U27552 (N_27552,N_25051,N_24086);
xnor U27553 (N_27553,N_26600,N_26128);
or U27554 (N_27554,N_25804,N_24642);
and U27555 (N_27555,N_25689,N_26505);
nand U27556 (N_27556,N_24414,N_25760);
xnor U27557 (N_27557,N_25645,N_25837);
xnor U27558 (N_27558,N_26545,N_25186);
nor U27559 (N_27559,N_24280,N_24510);
and U27560 (N_27560,N_24697,N_25581);
or U27561 (N_27561,N_24508,N_25938);
nand U27562 (N_27562,N_25460,N_24979);
xnor U27563 (N_27563,N_25330,N_24594);
and U27564 (N_27564,N_25718,N_26865);
or U27565 (N_27565,N_26125,N_24333);
or U27566 (N_27566,N_26437,N_25567);
xnor U27567 (N_27567,N_25913,N_24372);
and U27568 (N_27568,N_25174,N_26743);
or U27569 (N_27569,N_24479,N_26807);
nand U27570 (N_27570,N_24294,N_25065);
nor U27571 (N_27571,N_25621,N_25798);
nand U27572 (N_27572,N_24557,N_25323);
and U27573 (N_27573,N_25421,N_25742);
xor U27574 (N_27574,N_25841,N_24663);
nand U27575 (N_27575,N_25156,N_26376);
nor U27576 (N_27576,N_25799,N_26591);
xor U27577 (N_27577,N_26501,N_25656);
xnor U27578 (N_27578,N_24525,N_26237);
and U27579 (N_27579,N_26171,N_24431);
and U27580 (N_27580,N_24516,N_24227);
or U27581 (N_27581,N_24261,N_24164);
xor U27582 (N_27582,N_24297,N_25982);
or U27583 (N_27583,N_25500,N_26491);
nor U27584 (N_27584,N_26766,N_25845);
or U27585 (N_27585,N_25205,N_26282);
nor U27586 (N_27586,N_26262,N_26665);
nor U27587 (N_27587,N_25000,N_26435);
nand U27588 (N_27588,N_25161,N_25636);
xor U27589 (N_27589,N_26070,N_25462);
nand U27590 (N_27590,N_25527,N_24721);
nor U27591 (N_27591,N_24204,N_26717);
nand U27592 (N_27592,N_26038,N_26498);
or U27593 (N_27593,N_24925,N_25484);
and U27594 (N_27594,N_24728,N_25409);
xnor U27595 (N_27595,N_26087,N_24244);
and U27596 (N_27596,N_25136,N_26480);
and U27597 (N_27597,N_26460,N_24584);
and U27598 (N_27598,N_25184,N_25214);
or U27599 (N_27599,N_25508,N_25427);
nor U27600 (N_27600,N_24174,N_24007);
nand U27601 (N_27601,N_26374,N_26311);
and U27602 (N_27602,N_25832,N_25494);
nand U27603 (N_27603,N_26071,N_25189);
or U27604 (N_27604,N_26185,N_24104);
or U27605 (N_27605,N_24268,N_24169);
nor U27606 (N_27606,N_24225,N_25714);
and U27607 (N_27607,N_25350,N_25778);
nand U27608 (N_27608,N_25702,N_24032);
and U27609 (N_27609,N_24902,N_26541);
and U27610 (N_27610,N_24870,N_24131);
xnor U27611 (N_27611,N_24939,N_24087);
nand U27612 (N_27612,N_24591,N_24485);
nand U27613 (N_27613,N_26820,N_24685);
or U27614 (N_27614,N_25098,N_25066);
or U27615 (N_27615,N_24604,N_24957);
xnor U27616 (N_27616,N_25244,N_26365);
nand U27617 (N_27617,N_26106,N_26641);
and U27618 (N_27618,N_25888,N_24847);
nor U27619 (N_27619,N_25227,N_25176);
or U27620 (N_27620,N_25230,N_24248);
xor U27621 (N_27621,N_24095,N_25142);
nor U27622 (N_27622,N_26947,N_25211);
nand U27623 (N_27623,N_24136,N_25785);
nor U27624 (N_27624,N_25325,N_24749);
and U27625 (N_27625,N_26703,N_26273);
xor U27626 (N_27626,N_24763,N_24791);
xnor U27627 (N_27627,N_26872,N_26347);
or U27628 (N_27628,N_25770,N_26702);
xor U27629 (N_27629,N_25535,N_24535);
and U27630 (N_27630,N_25163,N_25369);
xor U27631 (N_27631,N_24655,N_25762);
xor U27632 (N_27632,N_26908,N_25868);
nor U27633 (N_27633,N_26255,N_25488);
or U27634 (N_27634,N_26251,N_24669);
and U27635 (N_27635,N_24568,N_26040);
xor U27636 (N_27636,N_24122,N_25548);
nor U27637 (N_27637,N_25489,N_25739);
nand U27638 (N_27638,N_24923,N_24327);
and U27639 (N_27639,N_26527,N_26705);
or U27640 (N_27640,N_26950,N_25115);
xor U27641 (N_27641,N_26539,N_24413);
nor U27642 (N_27642,N_25843,N_24815);
or U27643 (N_27643,N_24166,N_24734);
or U27644 (N_27644,N_25151,N_24278);
nor U27645 (N_27645,N_24978,N_24854);
xor U27646 (N_27646,N_25766,N_25694);
xnor U27647 (N_27647,N_25361,N_25816);
or U27648 (N_27648,N_26825,N_24486);
xor U27649 (N_27649,N_25959,N_26405);
nand U27650 (N_27650,N_24865,N_24285);
xor U27651 (N_27651,N_25281,N_24075);
nor U27652 (N_27652,N_24960,N_25164);
and U27653 (N_27653,N_24780,N_24570);
xnor U27654 (N_27654,N_24586,N_25815);
nand U27655 (N_27655,N_25170,N_25144);
xnor U27656 (N_27656,N_26920,N_24949);
nor U27657 (N_27657,N_24544,N_24115);
xnor U27658 (N_27658,N_25533,N_26653);
nand U27659 (N_27659,N_25665,N_26007);
or U27660 (N_27660,N_24456,N_25064);
nand U27661 (N_27661,N_24693,N_25617);
or U27662 (N_27662,N_25033,N_24521);
and U27663 (N_27663,N_26286,N_25138);
or U27664 (N_27664,N_25926,N_24068);
and U27665 (N_27665,N_26639,N_25679);
nor U27666 (N_27666,N_26758,N_26738);
and U27667 (N_27667,N_26910,N_24850);
and U27668 (N_27668,N_24215,N_25082);
and U27669 (N_27669,N_24720,N_26141);
nor U27670 (N_27670,N_24401,N_24725);
and U27671 (N_27671,N_26570,N_24631);
or U27672 (N_27672,N_24181,N_26002);
nand U27673 (N_27673,N_26572,N_24365);
or U27674 (N_27674,N_24666,N_25885);
or U27675 (N_27675,N_25060,N_26943);
and U27676 (N_27676,N_25916,N_24649);
nand U27677 (N_27677,N_24103,N_25311);
xor U27678 (N_27678,N_26244,N_24110);
or U27679 (N_27679,N_24766,N_25300);
xor U27680 (N_27680,N_25690,N_25988);
or U27681 (N_27681,N_25102,N_26593);
nor U27682 (N_27682,N_24157,N_24245);
nand U27683 (N_27683,N_26611,N_24439);
xor U27684 (N_27684,N_25658,N_24875);
nor U27685 (N_27685,N_24692,N_24698);
xnor U27686 (N_27686,N_25964,N_25912);
and U27687 (N_27687,N_25768,N_25047);
nand U27688 (N_27688,N_24794,N_26075);
xnor U27689 (N_27689,N_25600,N_24676);
nor U27690 (N_27690,N_25661,N_25241);
xor U27691 (N_27691,N_25584,N_24988);
xor U27692 (N_27692,N_26931,N_25220);
xor U27693 (N_27693,N_26060,N_26599);
nor U27694 (N_27694,N_24114,N_24074);
and U27695 (N_27695,N_24081,N_24002);
xor U27696 (N_27696,N_26748,N_24841);
or U27697 (N_27697,N_26977,N_25653);
or U27698 (N_27698,N_26195,N_25348);
and U27699 (N_27699,N_25968,N_25578);
nor U27700 (N_27700,N_26765,N_26289);
nand U27701 (N_27701,N_26280,N_25040);
nand U27702 (N_27702,N_25455,N_25400);
xor U27703 (N_27703,N_26192,N_24144);
xnor U27704 (N_27704,N_25305,N_26701);
and U27705 (N_27705,N_25949,N_26715);
nand U27706 (N_27706,N_25349,N_26848);
xor U27707 (N_27707,N_25834,N_24201);
or U27708 (N_27708,N_25634,N_25188);
nand U27709 (N_27709,N_24386,N_25744);
xnor U27710 (N_27710,N_26054,N_26946);
xnor U27711 (N_27711,N_26363,N_26225);
and U27712 (N_27712,N_26770,N_24823);
or U27713 (N_27713,N_26153,N_25139);
xnor U27714 (N_27714,N_26295,N_25963);
and U27715 (N_27715,N_25135,N_25642);
and U27716 (N_27716,N_25646,N_24867);
and U27717 (N_27717,N_25178,N_26455);
or U27718 (N_27718,N_24477,N_25969);
nor U27719 (N_27719,N_25476,N_25145);
and U27720 (N_27720,N_24339,N_24699);
or U27721 (N_27721,N_26864,N_25423);
and U27722 (N_27722,N_26793,N_25222);
nand U27723 (N_27723,N_25793,N_25856);
nor U27724 (N_27724,N_26934,N_26811);
nor U27725 (N_27725,N_25582,N_26823);
xor U27726 (N_27726,N_25957,N_26073);
xor U27727 (N_27727,N_24171,N_24303);
nor U27728 (N_27728,N_24845,N_24782);
nand U27729 (N_27729,N_25095,N_25709);
or U27730 (N_27730,N_26187,N_26305);
and U27731 (N_27731,N_24442,N_25580);
nor U27732 (N_27732,N_24102,N_25599);
xnor U27733 (N_27733,N_24733,N_26634);
or U27734 (N_27734,N_24786,N_26302);
nor U27735 (N_27735,N_24790,N_26343);
or U27736 (N_27736,N_26126,N_24826);
nor U27737 (N_27737,N_24646,N_25585);
nor U27738 (N_27738,N_24691,N_24396);
or U27739 (N_27739,N_25510,N_26196);
or U27740 (N_27740,N_24152,N_24387);
nand U27741 (N_27741,N_26648,N_25090);
or U27742 (N_27742,N_25909,N_26394);
nor U27743 (N_27743,N_25676,N_24314);
and U27744 (N_27744,N_25614,N_26348);
nor U27745 (N_27745,N_26112,N_25507);
nor U27746 (N_27746,N_25698,N_25377);
or U27747 (N_27747,N_25654,N_26901);
or U27748 (N_27748,N_25326,N_26999);
and U27749 (N_27749,N_26749,N_25848);
xnor U27750 (N_27750,N_26352,N_26063);
or U27751 (N_27751,N_26099,N_26140);
xor U27752 (N_27752,N_26142,N_24539);
xnor U27753 (N_27753,N_26321,N_25898);
xor U27754 (N_27754,N_25292,N_24335);
nor U27755 (N_27755,N_25536,N_26331);
or U27756 (N_27756,N_26676,N_24338);
xnor U27757 (N_27757,N_26132,N_25315);
and U27758 (N_27758,N_26238,N_26242);
and U27759 (N_27759,N_26521,N_24556);
and U27760 (N_27760,N_25528,N_25280);
xor U27761 (N_27761,N_26274,N_26160);
nand U27762 (N_27762,N_26775,N_24041);
nor U27763 (N_27763,N_26583,N_25124);
and U27764 (N_27764,N_25340,N_26987);
or U27765 (N_27765,N_25587,N_24873);
nor U27766 (N_27766,N_26559,N_26469);
or U27767 (N_27767,N_26606,N_24588);
xor U27768 (N_27768,N_25511,N_25800);
and U27769 (N_27769,N_26567,N_24161);
xor U27770 (N_27770,N_25070,N_24701);
or U27771 (N_27771,N_24779,N_26176);
xor U27772 (N_27772,N_24798,N_26278);
xor U27773 (N_27773,N_24483,N_24111);
nor U27774 (N_27774,N_26271,N_26408);
nor U27775 (N_27775,N_26380,N_26223);
xor U27776 (N_27776,N_25371,N_25784);
and U27777 (N_27777,N_26944,N_25181);
nand U27778 (N_27778,N_25998,N_24024);
nand U27779 (N_27779,N_24348,N_26296);
and U27780 (N_27780,N_24936,N_24197);
xor U27781 (N_27781,N_26936,N_26711);
or U27782 (N_27782,N_26779,N_25733);
nor U27783 (N_27783,N_24384,N_24576);
and U27784 (N_27784,N_25657,N_25758);
or U27785 (N_27785,N_26836,N_26432);
and U27786 (N_27786,N_26115,N_26897);
or U27787 (N_27787,N_25914,N_24565);
nand U27788 (N_27788,N_24851,N_26838);
or U27789 (N_27789,N_25458,N_25374);
nor U27790 (N_27790,N_26514,N_24857);
and U27791 (N_27791,N_25055,N_24953);
nand U27792 (N_27792,N_24608,N_24369);
nor U27793 (N_27793,N_26962,N_25074);
nand U27794 (N_27794,N_25020,N_25392);
or U27795 (N_27795,N_26451,N_24453);
xor U27796 (N_27796,N_24757,N_24079);
nand U27797 (N_27797,N_24703,N_25413);
nor U27798 (N_27798,N_25465,N_26418);
nand U27799 (N_27799,N_26921,N_25263);
nor U27800 (N_27800,N_25166,N_25368);
or U27801 (N_27801,N_25389,N_25683);
or U27802 (N_27802,N_25836,N_26516);
or U27803 (N_27803,N_25983,N_26888);
and U27804 (N_27804,N_24982,N_26041);
nand U27805 (N_27805,N_25644,N_25741);
and U27806 (N_27806,N_26233,N_26603);
nor U27807 (N_27807,N_26708,N_24895);
nand U27808 (N_27808,N_24281,N_25272);
nand U27809 (N_27809,N_24938,N_26552);
nand U27810 (N_27810,N_24611,N_25437);
or U27811 (N_27811,N_24449,N_26768);
xor U27812 (N_27812,N_24311,N_24300);
nand U27813 (N_27813,N_24071,N_25372);
and U27814 (N_27814,N_25607,N_26137);
nand U27815 (N_27815,N_26557,N_26235);
nor U27816 (N_27816,N_24004,N_25602);
xor U27817 (N_27817,N_24899,N_25256);
xnor U27818 (N_27818,N_26162,N_25447);
nand U27819 (N_27819,N_26085,N_26236);
nor U27820 (N_27820,N_26609,N_25068);
or U27821 (N_27821,N_26845,N_24209);
nor U27822 (N_27822,N_26808,N_25648);
nand U27823 (N_27823,N_25023,N_24672);
nand U27824 (N_27824,N_26419,N_24868);
or U27825 (N_27825,N_24706,N_24529);
xor U27826 (N_27826,N_25783,N_26954);
xor U27827 (N_27827,N_24678,N_24022);
nand U27828 (N_27828,N_25611,N_25406);
nor U27829 (N_27829,N_26359,N_26519);
or U27830 (N_27830,N_24880,N_25293);
nand U27831 (N_27831,N_26538,N_24951);
nand U27832 (N_27832,N_26485,N_25818);
xor U27833 (N_27833,N_24551,N_24773);
and U27834 (N_27834,N_26188,N_25668);
and U27835 (N_27835,N_25159,N_26428);
nor U27836 (N_27836,N_25480,N_24827);
nand U27837 (N_27837,N_26696,N_24073);
nor U27838 (N_27838,N_26205,N_25229);
and U27839 (N_27839,N_26190,N_25993);
nor U27840 (N_27840,N_24887,N_24940);
or U27841 (N_27841,N_24579,N_26005);
or U27842 (N_27842,N_25243,N_24200);
or U27843 (N_27843,N_26111,N_25076);
xor U27844 (N_27844,N_24277,N_26118);
nand U27845 (N_27845,N_25213,N_25779);
nor U27846 (N_27846,N_26672,N_25970);
or U27847 (N_27847,N_26134,N_26780);
or U27848 (N_27848,N_24931,N_25449);
nand U27849 (N_27849,N_26277,N_25012);
or U27850 (N_27850,N_26313,N_24101);
xnor U27851 (N_27851,N_26918,N_25367);
or U27852 (N_27852,N_25724,N_26062);
xor U27853 (N_27853,N_24482,N_24368);
nor U27854 (N_27854,N_26763,N_24018);
xnor U27855 (N_27855,N_24812,N_25072);
xnor U27856 (N_27856,N_26024,N_24616);
nor U27857 (N_27857,N_25376,N_25356);
or U27858 (N_27858,N_26668,N_24937);
nor U27859 (N_27859,N_24180,N_24496);
and U27860 (N_27860,N_26939,N_24239);
xor U27861 (N_27861,N_26309,N_24659);
xor U27862 (N_27862,N_26001,N_25495);
xor U27863 (N_27863,N_26868,N_24778);
xnor U27864 (N_27864,N_25320,N_26210);
nor U27865 (N_27865,N_24186,N_26212);
nand U27866 (N_27866,N_24289,N_24433);
nand U27867 (N_27867,N_25894,N_25990);
nand U27868 (N_27868,N_26565,N_25010);
or U27869 (N_27869,N_25497,N_25738);
xnor U27870 (N_27870,N_25594,N_25443);
nand U27871 (N_27871,N_26834,N_26179);
xor U27872 (N_27872,N_26439,N_25972);
xor U27873 (N_27873,N_25433,N_25919);
and U27874 (N_27874,N_24927,N_26467);
nor U27875 (N_27875,N_24954,N_24468);
or U27876 (N_27876,N_24785,N_26120);
and U27877 (N_27877,N_26372,N_25757);
nor U27878 (N_27878,N_26065,N_25598);
or U27879 (N_27879,N_26615,N_26299);
and U27880 (N_27880,N_26492,N_25226);
and U27881 (N_27881,N_24282,N_24377);
nor U27882 (N_27882,N_25363,N_25298);
nand U27883 (N_27883,N_26952,N_26975);
or U27884 (N_27884,N_24644,N_25251);
nor U27885 (N_27885,N_26315,N_26960);
nand U27886 (N_27886,N_25677,N_24109);
nand U27887 (N_27887,N_25505,N_26913);
or U27888 (N_27888,N_26734,N_26234);
nor U27889 (N_27889,N_24752,N_26074);
xnor U27890 (N_27890,N_25236,N_26822);
nand U27891 (N_27891,N_24305,N_24175);
nor U27892 (N_27892,N_25208,N_25201);
or U27893 (N_27893,N_24968,N_25146);
and U27894 (N_27894,N_24704,N_25045);
and U27895 (N_27895,N_26344,N_25678);
nand U27896 (N_27896,N_26043,N_24894);
nor U27897 (N_27897,N_26607,N_24797);
or U27898 (N_27898,N_24614,N_24803);
or U27899 (N_27899,N_24587,N_26844);
xnor U27900 (N_27900,N_26193,N_25380);
or U27901 (N_27901,N_25113,N_26367);
and U27902 (N_27902,N_24228,N_25346);
nand U27903 (N_27903,N_26898,N_24719);
and U27904 (N_27904,N_24560,N_25385);
and U27905 (N_27905,N_25459,N_26547);
nand U27906 (N_27906,N_24893,N_25399);
nand U27907 (N_27907,N_26622,N_25721);
or U27908 (N_27908,N_25264,N_26546);
or U27909 (N_27909,N_25995,N_26630);
xnor U27910 (N_27910,N_25876,N_26613);
and U27911 (N_27911,N_24801,N_26483);
nor U27912 (N_27912,N_26250,N_26409);
nor U27913 (N_27913,N_26827,N_26334);
xor U27914 (N_27914,N_25134,N_26680);
nand U27915 (N_27915,N_25141,N_25513);
nor U27916 (N_27916,N_25996,N_25410);
xnor U27917 (N_27917,N_24015,N_25125);
xnor U27918 (N_27918,N_26875,N_24243);
or U27919 (N_27919,N_26785,N_24622);
nor U27920 (N_27920,N_26555,N_25712);
or U27921 (N_27921,N_24829,N_26870);
nand U27922 (N_27922,N_26810,N_26729);
nor U27923 (N_27923,N_24768,N_25150);
nand U27924 (N_27924,N_24035,N_24448);
nor U27925 (N_27925,N_26876,N_24533);
nor U27926 (N_27926,N_26562,N_25283);
xor U27927 (N_27927,N_26199,N_25824);
or U27928 (N_27928,N_24545,N_24564);
or U27929 (N_27929,N_24609,N_24187);
xnor U27930 (N_27930,N_26725,N_25103);
and U27931 (N_27931,N_24901,N_25638);
nor U27932 (N_27932,N_26381,N_26218);
xnor U27933 (N_27933,N_24199,N_26357);
xnor U27934 (N_27934,N_26478,N_25999);
or U27935 (N_27935,N_24350,N_25018);
or U27936 (N_27936,N_26003,N_24241);
and U27937 (N_27937,N_26095,N_26345);
xnor U27938 (N_27938,N_24532,N_26663);
and U27939 (N_27939,N_24213,N_25663);
nor U27940 (N_27940,N_24304,N_25133);
xnor U27941 (N_27941,N_25515,N_24246);
nand U27942 (N_27942,N_26940,N_25137);
xnor U27943 (N_27943,N_25947,N_24983);
or U27944 (N_27944,N_26767,N_25104);
or U27945 (N_27945,N_24249,N_25119);
nor U27946 (N_27946,N_24135,N_26774);
nand U27947 (N_27947,N_26788,N_24113);
nor U27948 (N_27948,N_24206,N_25192);
nand U27949 (N_27949,N_25979,N_25093);
and U27950 (N_27950,N_25795,N_26316);
xnor U27951 (N_27951,N_24814,N_26067);
and U27952 (N_27952,N_24301,N_24863);
nand U27953 (N_27953,N_24467,N_26107);
and U27954 (N_27954,N_24811,N_25200);
xor U27955 (N_27955,N_24571,N_26571);
xnor U27956 (N_27956,N_25922,N_24689);
nand U27957 (N_27957,N_24489,N_26762);
and U27958 (N_27958,N_26790,N_25080);
nand U27959 (N_27959,N_25335,N_25037);
nor U27960 (N_27960,N_24221,N_25971);
and U27961 (N_27961,N_26275,N_26966);
or U27962 (N_27962,N_26484,N_24885);
and U27963 (N_27963,N_24879,N_24220);
xnor U27964 (N_27964,N_25811,N_25953);
or U27965 (N_27965,N_24423,N_25182);
and U27966 (N_27966,N_26015,N_24216);
xnor U27967 (N_27967,N_26714,N_26632);
nor U27968 (N_27968,N_26890,N_26297);
nand U27969 (N_27969,N_26023,N_25731);
and U27970 (N_27970,N_26391,N_24530);
nand U27971 (N_27971,N_24046,N_26369);
or U27972 (N_27972,N_26358,N_25210);
nor U27973 (N_27973,N_25672,N_24443);
xor U27974 (N_27974,N_24718,N_26396);
nor U27975 (N_27975,N_26198,N_26263);
nand U27976 (N_27976,N_25331,N_25075);
and U27977 (N_27977,N_26399,N_24264);
xor U27978 (N_27978,N_25674,N_26157);
nor U27979 (N_27979,N_26899,N_25061);
xnor U27980 (N_27980,N_25118,N_25680);
xor U27981 (N_27981,N_25509,N_24473);
nand U27982 (N_27982,N_26216,N_24019);
xnor U27983 (N_27983,N_24159,N_25411);
or U27984 (N_27984,N_26661,N_25826);
nor U27985 (N_27985,N_24498,N_26884);
and U27986 (N_27986,N_26476,N_26885);
xor U27987 (N_27987,N_25337,N_26732);
nor U27988 (N_27988,N_26813,N_24999);
nor U27989 (N_27989,N_25532,N_24016);
and U27990 (N_27990,N_25948,N_25651);
nor U27991 (N_27991,N_24233,N_25956);
or U27992 (N_27992,N_25196,N_26387);
nand U27993 (N_27993,N_25596,N_26298);
nor U27994 (N_27994,N_24235,N_25155);
and U27995 (N_27995,N_26042,N_24683);
and U27996 (N_27996,N_26082,N_26246);
xor U27997 (N_27997,N_26854,N_24740);
or U27998 (N_27998,N_26837,N_25428);
and U27999 (N_27999,N_25701,N_26802);
nand U28000 (N_28000,N_25960,N_25276);
xor U28001 (N_28001,N_24404,N_25370);
xor U28002 (N_28002,N_26079,N_26855);
xor U28003 (N_28003,N_24432,N_26508);
or U28004 (N_28004,N_24711,N_26747);
and U28005 (N_28005,N_26984,N_26502);
nand U28006 (N_28006,N_25904,N_25781);
and U28007 (N_28007,N_24831,N_24108);
or U28008 (N_28008,N_26773,N_26517);
and U28009 (N_28009,N_26801,N_25454);
nor U28010 (N_28010,N_26037,N_25840);
xor U28011 (N_28011,N_25801,N_24344);
xor U28012 (N_28012,N_24218,N_25416);
xnor U28013 (N_28013,N_26581,N_25031);
nand U28014 (N_28014,N_24619,N_26867);
nand U28015 (N_28015,N_26017,N_26564);
xor U28016 (N_28016,N_24412,N_25844);
nand U28017 (N_28017,N_24054,N_26698);
xor U28018 (N_28018,N_25223,N_24578);
or U28019 (N_28019,N_26444,N_25514);
nand U28020 (N_28020,N_25474,N_25649);
or U28021 (N_28021,N_26726,N_25185);
nand U28022 (N_28022,N_24620,N_24705);
xor U28023 (N_28023,N_24563,N_24203);
nand U28024 (N_28024,N_24262,N_26695);
and U28025 (N_28025,N_24168,N_25195);
nor U28026 (N_28026,N_24959,N_26993);
nand U28027 (N_28027,N_25560,N_25499);
nor U28028 (N_28028,N_24347,N_24708);
nand U28029 (N_28029,N_25734,N_26569);
nand U28030 (N_28030,N_24038,N_24219);
or U28031 (N_28031,N_25692,N_26048);
or U28032 (N_28032,N_26211,N_24751);
nor U28033 (N_28033,N_26598,N_24888);
xor U28034 (N_28034,N_25544,N_25365);
or U28035 (N_28035,N_26078,N_25592);
and U28036 (N_28036,N_26222,N_24781);
nand U28037 (N_28037,N_25819,N_24198);
nand U28038 (N_28038,N_26540,N_24992);
or U28039 (N_28039,N_24097,N_25341);
and U28040 (N_28040,N_25950,N_25790);
nor U28041 (N_28041,N_26675,N_25807);
nand U28042 (N_28042,N_24917,N_24813);
nand U28043 (N_28043,N_24896,N_25260);
xnor U28044 (N_28044,N_26411,N_26281);
xnor U28045 (N_28045,N_26588,N_25216);
nand U28046 (N_28046,N_25659,N_24422);
nand U28047 (N_28047,N_26404,N_25172);
nor U28048 (N_28048,N_26824,N_24946);
nor U28049 (N_28049,N_24126,N_24330);
xnor U28050 (N_28050,N_25937,N_26797);
nor U28051 (N_28051,N_25590,N_24288);
or U28052 (N_28052,N_25907,N_24590);
or U28053 (N_28053,N_25209,N_26370);
nand U28054 (N_28054,N_26631,N_25088);
nand U28055 (N_28055,N_25152,N_26221);
xor U28056 (N_28056,N_25545,N_26651);
nor U28057 (N_28057,N_25561,N_26012);
nor U28058 (N_28058,N_25358,N_24258);
xnor U28059 (N_28059,N_24996,N_26828);
or U28060 (N_28060,N_25899,N_24325);
or U28061 (N_28061,N_24395,N_24013);
nor U28062 (N_28062,N_26803,N_26464);
nor U28063 (N_28063,N_25786,N_26719);
xor U28064 (N_28064,N_26146,N_24378);
and U28065 (N_28065,N_25973,N_24966);
nor U28066 (N_28066,N_24920,N_26662);
xor U28067 (N_28067,N_24891,N_24817);
nor U28068 (N_28068,N_26317,N_24500);
nand U28069 (N_28069,N_24257,N_25313);
nand U28070 (N_28070,N_24764,N_24595);
and U28071 (N_28071,N_26183,N_25622);
xnor U28072 (N_28072,N_25401,N_24769);
and U28073 (N_28073,N_25862,N_25041);
and U28074 (N_28074,N_25965,N_26036);
nand U28075 (N_28075,N_24345,N_24094);
xor U28076 (N_28076,N_25394,N_26949);
xnor U28077 (N_28077,N_24426,N_25568);
nor U28078 (N_28078,N_26981,N_25307);
or U28079 (N_28079,N_24230,N_26869);
nor U28080 (N_28080,N_24617,N_24051);
nand U28081 (N_28081,N_26643,N_26548);
xnor U28082 (N_28082,N_24932,N_24657);
nand U28083 (N_28083,N_24548,N_25132);
nand U28084 (N_28084,N_24296,N_25275);
nand U28085 (N_28085,N_26733,N_24149);
xor U28086 (N_28086,N_24921,N_24320);
xnor U28087 (N_28087,N_24030,N_26617);
nor U28088 (N_28088,N_25258,N_24298);
nor U28089 (N_28089,N_26689,N_25735);
and U28090 (N_28090,N_26379,N_25193);
or U28091 (N_28091,N_25228,N_24354);
nand U28092 (N_28092,N_24520,N_24511);
nor U28093 (N_28093,N_25217,N_25456);
xnor U28094 (N_28094,N_24242,N_24765);
or U28095 (N_28095,N_26948,N_26757);
and U28096 (N_28096,N_25928,N_24323);
xnor U28097 (N_28097,N_26039,N_25048);
and U28098 (N_28098,N_26657,N_24597);
nor U28099 (N_28099,N_24222,N_26092);
nor U28100 (N_28100,N_26900,N_24259);
nor U28101 (N_28101,N_24969,N_26231);
nor U28102 (N_28102,N_24145,N_25092);
nor U28103 (N_28103,N_24042,N_25962);
nand U28104 (N_28104,N_24635,N_24463);
nand U28105 (N_28105,N_24121,N_24254);
nand U28106 (N_28106,N_25206,N_25221);
nor U28107 (N_28107,N_26044,N_24820);
or U28108 (N_28108,N_25463,N_26416);
nand U28109 (N_28109,N_26777,N_25650);
nand U28110 (N_28110,N_25613,N_26923);
nor U28111 (N_28111,N_25485,N_25441);
xor U28112 (N_28112,N_24912,N_26161);
and U28113 (N_28113,N_25250,N_24515);
nand U28114 (N_28114,N_26795,N_24450);
xor U28115 (N_28115,N_24730,N_25751);
nand U28116 (N_28116,N_26831,N_26427);
xnor U28117 (N_28117,N_24172,N_25269);
and U28118 (N_28118,N_25671,N_24524);
and U28119 (N_28119,N_24429,N_26982);
xnor U28120 (N_28120,N_24469,N_26294);
or U28121 (N_28121,N_24132,N_25347);
and U28122 (N_28122,N_26252,N_26582);
xor U28123 (N_28123,N_26731,N_26523);
nand U28124 (N_28124,N_26247,N_24346);
or U28125 (N_28125,N_25986,N_24799);
and U28126 (N_28126,N_24428,N_24746);
or U28127 (N_28127,N_25620,N_26894);
xnor U28128 (N_28128,N_24818,N_26988);
or U28129 (N_28129,N_24029,N_26692);
and U28130 (N_28130,N_26117,N_26163);
or U28131 (N_28131,N_24900,N_25765);
xor U28132 (N_28132,N_24598,N_25827);
nand U28133 (N_28133,N_25038,N_25318);
or U28134 (N_28134,N_26031,N_26463);
or U28135 (N_28135,N_24661,N_26217);
nor U28136 (N_28136,N_24628,N_25682);
nor U28137 (N_28137,N_25490,N_25479);
nand U28138 (N_28138,N_25354,N_26553);
and U28139 (N_28139,N_24451,N_25874);
or U28140 (N_28140,N_26131,N_24250);
nand U28141 (N_28141,N_24006,N_26882);
and U28142 (N_28142,N_26342,N_26902);
and U28143 (N_28143,N_26575,N_25171);
nor U28144 (N_28144,N_25855,N_24251);
and U28145 (N_28145,N_24626,N_24918);
xnor U28146 (N_28146,N_24664,N_26441);
nand U28147 (N_28147,N_24933,N_26512);
nor U28148 (N_28148,N_25373,N_26629);
nor U28149 (N_28149,N_26667,N_25110);
or U28150 (N_28150,N_26472,N_26016);
nor U28151 (N_28151,N_25063,N_25425);
or U28152 (N_28152,N_24915,N_25583);
xnor U28153 (N_28153,N_25934,N_24770);
or U28154 (N_28154,N_26697,N_25154);
xnor U28155 (N_28155,N_25017,N_25716);
or U28156 (N_28156,N_25542,N_26008);
xor U28157 (N_28157,N_24292,N_25396);
xnor U28158 (N_28158,N_25052,N_26239);
nor U28159 (N_28159,N_24418,N_26213);
xor U28160 (N_28160,N_24039,N_26577);
xor U28161 (N_28161,N_25877,N_24390);
nor U28162 (N_28162,N_24084,N_24063);
nor U28163 (N_28163,N_24358,N_25175);
and U28164 (N_28164,N_26974,N_25624);
and U28165 (N_28165,N_25550,N_25008);
and U28166 (N_28166,N_25249,N_25359);
and U28167 (N_28167,N_26076,N_26382);
xor U28168 (N_28168,N_24059,N_25713);
nand U28169 (N_28169,N_26925,N_24522);
nand U28170 (N_28170,N_24240,N_24188);
or U28171 (N_28171,N_24020,N_26740);
nand U28172 (N_28172,N_24163,N_26784);
nand U28173 (N_28173,N_24714,N_25529);
nor U28174 (N_28174,N_24762,N_24881);
nor U28175 (N_28175,N_26563,N_25419);
nand U28176 (N_28176,N_25173,N_26744);
xnor U28177 (N_28177,N_26852,N_26285);
nor U28178 (N_28178,N_26531,N_26489);
xnor U28179 (N_28179,N_24911,N_25708);
nor U28180 (N_28180,N_26883,N_26496);
xnor U28181 (N_28181,N_26249,N_25942);
and U28182 (N_28182,N_24702,N_25397);
xnor U28183 (N_28183,N_25869,N_26471);
and U28184 (N_28184,N_26537,N_26173);
and U28185 (N_28185,N_24446,N_25289);
and U28186 (N_28186,N_25740,N_25882);
or U28187 (N_28187,N_24976,N_26448);
nor U28188 (N_28188,N_25202,N_24528);
nand U28189 (N_28189,N_26819,N_25764);
or U28190 (N_28190,N_25165,N_26674);
or U28191 (N_28191,N_24411,N_24210);
and U28192 (N_28192,N_25062,N_25408);
nor U28193 (N_28193,N_26592,N_24052);
nor U28194 (N_28194,N_25847,N_26398);
xnor U28195 (N_28195,N_24546,N_25149);
xnor U28196 (N_28196,N_25007,N_25422);
and U28197 (N_28197,N_24367,N_26647);
and U28198 (N_28198,N_25388,N_25169);
and U28199 (N_28199,N_24688,N_26004);
nor U28200 (N_28200,N_26628,N_24009);
and U28201 (N_28201,N_25042,N_24574);
nor U28202 (N_28202,N_25575,N_26789);
nand U28203 (N_28203,N_24589,N_25880);
nand U28204 (N_28204,N_24205,N_26021);
nand U28205 (N_28205,N_26053,N_26771);
nand U28206 (N_28206,N_26528,N_24846);
or U28207 (N_28207,N_25752,N_26906);
xnor U28208 (N_28208,N_25285,N_25308);
and U28209 (N_28209,N_24283,N_24148);
nor U28210 (N_28210,N_24034,N_26739);
nand U28211 (N_28211,N_26997,N_25669);
xnor U28212 (N_28212,N_24737,N_24869);
and U28213 (N_28213,N_25543,N_26594);
and U28214 (N_28214,N_24231,N_24833);
or U28215 (N_28215,N_26928,N_25601);
nor U28216 (N_28216,N_24326,N_24083);
or U28217 (N_28217,N_24935,N_24961);
nor U28218 (N_28218,N_25710,N_24596);
xnor U28219 (N_28219,N_25530,N_24859);
nor U28220 (N_28220,N_26805,N_24955);
and U28221 (N_28221,N_25491,N_25087);
nor U28222 (N_28222,N_26284,N_24340);
xnor U28223 (N_28223,N_24315,N_24997);
or U28224 (N_28224,N_24211,N_26414);
nor U28225 (N_28225,N_24322,N_25685);
nor U28226 (N_28226,N_26985,N_25866);
xnor U28227 (N_28227,N_26927,N_24753);
xnor U28228 (N_28228,N_24849,N_25344);
and U28229 (N_28229,N_24700,N_24855);
or U28230 (N_28230,N_26534,N_25069);
nor U28231 (N_28231,N_24848,N_26229);
nand U28232 (N_28232,N_24342,N_24070);
nand U28233 (N_28233,N_26488,N_26209);
or U28234 (N_28234,N_25887,N_25310);
and U28235 (N_28235,N_24995,N_24687);
nand U28236 (N_28236,N_24078,N_25573);
nor U28237 (N_28237,N_25519,N_24922);
nor U28238 (N_28238,N_24271,N_25538);
nand U28239 (N_28239,N_24256,N_26652);
and U28240 (N_28240,N_26741,N_25609);
xor U28241 (N_28241,N_26859,N_26386);
nand U28242 (N_28242,N_26560,N_26724);
xor U28243 (N_28243,N_24099,N_26292);
and U28244 (N_28244,N_25551,N_26029);
nor U28245 (N_28245,N_26842,N_25345);
nand U28246 (N_28246,N_26006,N_26690);
or U28247 (N_28247,N_24371,N_24406);
nor U28248 (N_28248,N_24394,N_24632);
nor U28249 (N_28249,N_26172,N_25057);
nor U28250 (N_28250,N_25106,N_26682);
nor U28251 (N_28251,N_25451,N_26051);
nand U28252 (N_28252,N_24637,N_26025);
or U28253 (N_28253,N_25577,N_26712);
xor U28254 (N_28254,N_26270,N_24176);
nand U28255 (N_28255,N_25606,N_24366);
and U28256 (N_28256,N_26035,N_24755);
nor U28257 (N_28257,N_24061,N_24639);
xor U28258 (N_28258,N_25749,N_25407);
nand U28259 (N_28259,N_25923,N_26658);
and U28260 (N_28260,N_25563,N_24889);
and U28261 (N_28261,N_25254,N_26248);
or U28262 (N_28262,N_26168,N_25049);
xor U28263 (N_28263,N_25525,N_24363);
nand U28264 (N_28264,N_25418,N_24430);
and U28265 (N_28265,N_26938,N_26356);
and U28266 (N_28266,N_24252,N_26685);
and U28267 (N_28267,N_25475,N_26392);
and U28268 (N_28268,N_26481,N_25180);
or U28269 (N_28269,N_25787,N_25191);
nor U28270 (N_28270,N_24208,N_26339);
or U28271 (N_28271,N_24975,N_26136);
and U28272 (N_28272,N_25107,N_25941);
xnor U28273 (N_28273,N_24821,N_25114);
or U28274 (N_28274,N_26000,N_25967);
or U28275 (N_28275,N_25857,N_24267);
or U28276 (N_28276,N_24402,N_26626);
nand U28277 (N_28277,N_24583,N_25316);
nand U28278 (N_28278,N_26706,N_25081);
xor U28279 (N_28279,N_25893,N_25566);
and U28280 (N_28280,N_24127,N_26383);
and U28281 (N_28281,N_25268,N_25557);
and U28282 (N_28282,N_26880,N_26167);
xnor U28283 (N_28283,N_24392,N_24247);
xor U28284 (N_28284,N_26090,N_26616);
nand U28285 (N_28285,N_26558,N_24802);
nor U28286 (N_28286,N_25157,N_24353);
xnor U28287 (N_28287,N_24948,N_25011);
xnor U28288 (N_28288,N_26754,N_26951);
xnor U28289 (N_28289,N_25828,N_24388);
nand U28290 (N_28290,N_26479,N_24272);
or U28291 (N_28291,N_25812,N_24822);
nor U28292 (N_28292,N_24930,N_25966);
nor U28293 (N_28293,N_25238,N_24710);
and U28294 (N_28294,N_26863,N_25892);
nand U28295 (N_28295,N_26440,N_24998);
or U28296 (N_28296,N_24476,N_26625);
or U28297 (N_28297,N_26812,N_24356);
xor U28298 (N_28298,N_24452,N_25009);
nor U28299 (N_28299,N_26186,N_25662);
xnor U28300 (N_28300,N_24634,N_26310);
and U28301 (N_28301,N_26850,N_24359);
nor U28302 (N_28302,N_24064,N_24527);
nand U28303 (N_28303,N_24884,N_25612);
nor U28304 (N_28304,N_24069,N_24572);
and U28305 (N_28305,N_25878,N_24956);
xor U28306 (N_28306,N_26787,N_25910);
nand U28307 (N_28307,N_24310,N_24603);
and U28308 (N_28308,N_26700,N_26722);
nand U28309 (N_28309,N_26410,N_24774);
xnor U28310 (N_28310,N_26047,N_26208);
nor U28311 (N_28311,N_25317,N_24573);
and U28312 (N_28312,N_24021,N_24555);
or U28313 (N_28313,N_26314,N_25754);
nor U28314 (N_28314,N_24793,N_26425);
or U28315 (N_28315,N_24796,N_24550);
or U28316 (N_28316,N_24266,N_25417);
nor U28317 (N_28317,N_25116,N_24011);
xnor U28318 (N_28318,N_24435,N_26549);
or U28319 (N_28319,N_26839,N_25572);
and U28320 (N_28320,N_26710,N_26886);
nor U28321 (N_28321,N_24417,N_24360);
and U28322 (N_28322,N_24125,N_24287);
nand U28323 (N_28323,N_25829,N_26595);
xor U28324 (N_28324,N_25610,N_25343);
or U28325 (N_28325,N_24492,N_26422);
nand U28326 (N_28326,N_26681,N_25992);
nand U28327 (N_28327,N_24592,N_25431);
xnor U28328 (N_28328,N_25019,N_26849);
or U28329 (N_28329,N_25774,N_25593);
nor U28330 (N_28330,N_26574,N_24600);
and U28331 (N_28331,N_25788,N_24364);
nand U28332 (N_28332,N_24674,N_24537);
nand U28333 (N_28333,N_26561,N_25168);
nor U28334 (N_28334,N_24623,N_26809);
and U28335 (N_28335,N_24950,N_25773);
nor U28336 (N_28336,N_24349,N_25796);
nor U28337 (N_28337,N_25579,N_24910);
or U28338 (N_28338,N_24284,N_24903);
or U28339 (N_28339,N_25745,N_26288);
or U28340 (N_28340,N_24825,N_26064);
or U28341 (N_28341,N_25274,N_24012);
or U28342 (N_28342,N_25918,N_24195);
nor U28343 (N_28343,N_24057,N_24105);
and U28344 (N_28344,N_25897,N_24944);
nor U28345 (N_28345,N_24269,N_26102);
and U28346 (N_28346,N_26423,N_24273);
nand U28347 (N_28347,N_26578,N_26556);
nand U28348 (N_28348,N_25199,N_24389);
nor U28349 (N_28349,N_26660,N_26022);
or U28350 (N_28350,N_26420,N_26431);
xor U28351 (N_28351,N_26368,N_24828);
nor U28352 (N_28352,N_24028,N_24129);
nand U28353 (N_28353,N_24055,N_26135);
nor U28354 (N_28354,N_26986,N_26709);
nor U28355 (N_28355,N_26049,N_26955);
xor U28356 (N_28356,N_25089,N_25961);
xor U28357 (N_28357,N_25393,N_26181);
nor U28358 (N_28358,N_24860,N_25630);
and U28359 (N_28359,N_24357,N_24178);
nand U28360 (N_28360,N_26907,N_25822);
and U28361 (N_28361,N_25352,N_24712);
xor U28362 (N_28362,N_25997,N_26197);
nor U28363 (N_28363,N_26786,N_25952);
nand U28364 (N_28364,N_24994,N_25212);
or U28365 (N_28365,N_24507,N_25006);
xnor U28366 (N_28366,N_26866,N_25383);
nand U28367 (N_28367,N_26889,N_25655);
nor U28368 (N_28368,N_24722,N_26500);
and U28369 (N_28369,N_24878,N_24373);
nor U28370 (N_28370,N_26746,N_26240);
or U28371 (N_28371,N_25539,N_26916);
xor U28372 (N_28372,N_25523,N_26335);
xnor U28373 (N_28373,N_24914,N_26056);
nor U28374 (N_28374,N_25034,N_26045);
or U28375 (N_28375,N_25619,N_25032);
xor U28376 (N_28376,N_25520,N_24926);
xnor U28377 (N_28377,N_25448,N_26261);
and U28378 (N_28378,N_25775,N_25360);
nor U28379 (N_28379,N_24514,N_26851);
or U28380 (N_28380,N_26245,N_26655);
or U28381 (N_28381,N_26798,N_25162);
xnor U28382 (N_28382,N_26018,N_24581);
or U28383 (N_28383,N_25842,N_25547);
xor U28384 (N_28384,N_24141,N_26513);
nor U28385 (N_28385,N_25747,N_26341);
nor U28386 (N_28386,N_24237,N_24554);
xnor U28387 (N_28387,N_25833,N_25122);
nor U28388 (N_28388,N_25943,N_26329);
xor U28389 (N_28389,N_26623,N_24776);
or U28390 (N_28390,N_24602,N_25291);
nor U28391 (N_28391,N_24060,N_25791);
and U28392 (N_28392,N_25452,N_25838);
and U28393 (N_28393,N_25763,N_26678);
and U28394 (N_28394,N_24987,N_25906);
and U28395 (N_28395,N_26175,N_25429);
nor U28396 (N_28396,N_24265,N_25911);
or U28397 (N_28397,N_24464,N_26473);
nor U28398 (N_28398,N_26804,N_25604);
nand U28399 (N_28399,N_24332,N_26637);
and U28400 (N_28400,N_24001,N_25569);
nand U28401 (N_28401,N_25128,N_26149);
xor U28402 (N_28402,N_24680,N_26716);
and U28403 (N_28403,N_24391,N_26219);
or U28404 (N_28404,N_25667,N_24182);
and U28405 (N_28405,N_26998,N_25854);
xor U28406 (N_28406,N_24756,N_24906);
or U28407 (N_28407,N_26881,N_25005);
xnor U28408 (N_28408,N_24092,N_24080);
xnor U28409 (N_28409,N_25875,N_24808);
nand U28410 (N_28410,N_25294,N_24307);
or U28411 (N_28411,N_25278,N_24472);
and U28412 (N_28412,N_26232,N_24053);
or U28413 (N_28413,N_25083,N_25570);
or U28414 (N_28414,N_24716,N_24008);
nand U28415 (N_28415,N_25664,N_25190);
or U28416 (N_28416,N_25987,N_24613);
nor U28417 (N_28417,N_26669,N_24726);
or U28418 (N_28418,N_24767,N_24919);
nor U28419 (N_28419,N_26338,N_26152);
xnor U28420 (N_28420,N_26755,N_25704);
nand U28421 (N_28421,N_26426,N_24306);
and U28422 (N_28422,N_24947,N_26761);
xor U28423 (N_28423,N_26835,N_24302);
nor U28424 (N_28424,N_25939,N_24742);
or U28425 (N_28425,N_24308,N_25688);
and U28426 (N_28426,N_26858,N_25440);
and U28427 (N_28427,N_24040,N_26945);
or U28428 (N_28428,N_26781,N_25975);
and U28429 (N_28429,N_25234,N_25627);
nor U28430 (N_28430,N_25056,N_24977);
nand U28431 (N_28431,N_24650,N_26646);
or U28432 (N_28432,N_25944,N_24909);
and U28433 (N_28433,N_26340,N_24461);
xor U28434 (N_28434,N_26573,N_25148);
or U28435 (N_28435,N_25029,N_26241);
or U28436 (N_28436,N_26980,N_25813);
xor U28437 (N_28437,N_24871,N_26751);
nor U28438 (N_28438,N_26704,N_26654);
xnor U28439 (N_28439,N_26319,N_26052);
nand U28440 (N_28440,N_24165,N_26096);
or U28441 (N_28441,N_26144,N_26587);
nand U28442 (N_28442,N_24290,N_24724);
xnor U28443 (N_28443,N_26904,N_24904);
nor U28444 (N_28444,N_25432,N_24962);
xor U28445 (N_28445,N_24160,N_24601);
nand U28446 (N_28446,N_26707,N_25398);
nor U28447 (N_28447,N_25931,N_26113);
nor U28448 (N_28448,N_24192,N_26937);
or U28449 (N_28449,N_25242,N_26293);
and U28450 (N_28450,N_26116,N_24913);
nor U28451 (N_28451,N_25324,N_24684);
or U28452 (N_28452,N_26290,N_26919);
or U28453 (N_28453,N_26964,N_26610);
or U28454 (N_28454,N_24748,N_26821);
xor U28455 (N_28455,N_26438,N_25483);
or U28456 (N_28456,N_24658,N_24458);
nand U28457 (N_28457,N_26330,N_24341);
or U28458 (N_28458,N_26121,N_26893);
and U28459 (N_28459,N_26776,N_24096);
or U28460 (N_28460,N_24876,N_25481);
xnor U28461 (N_28461,N_26081,N_26475);
nand U28462 (N_28462,N_25873,N_24523);
or U28463 (N_28463,N_25108,N_26832);
or U28464 (N_28464,N_26895,N_26636);
xor U28465 (N_28465,N_24866,N_26110);
or U28466 (N_28466,N_26608,N_24143);
xnor U28467 (N_28467,N_25295,N_24150);
xnor U28468 (N_28468,N_25759,N_25438);
nand U28469 (N_28469,N_24660,N_26922);
or U28470 (N_28470,N_25362,N_24965);
and U28471 (N_28471,N_25247,N_24509);
nor U28472 (N_28472,N_25687,N_26506);
nand U28473 (N_28473,N_26182,N_24618);
and U28474 (N_28474,N_24437,N_24824);
or U28475 (N_28475,N_24788,N_25905);
and U28476 (N_28476,N_24434,N_26568);
xor U28477 (N_28477,N_24980,N_25415);
nor U28478 (N_28478,N_26127,N_25079);
nand U28479 (N_28479,N_24224,N_25925);
xnor U28480 (N_28480,N_24747,N_25810);
xnor U28481 (N_28481,N_24580,N_26312);
nor U28482 (N_28482,N_24853,N_25445);
xnor U28483 (N_28483,N_26877,N_26201);
and U28484 (N_28484,N_25299,N_26543);
and U28485 (N_28485,N_24441,N_26542);
xnor U28486 (N_28486,N_25618,N_26713);
nor U28487 (N_28487,N_25633,N_26536);
nor U28488 (N_28488,N_25224,N_25273);
nand U28489 (N_28489,N_26474,N_24337);
or U28490 (N_28490,N_26800,N_25457);
xnor U28491 (N_28491,N_26443,N_25482);
or U28492 (N_28492,N_25225,N_26533);
nand U28493 (N_28493,N_26291,N_24481);
xor U28494 (N_28494,N_25099,N_24625);
nand U28495 (N_28495,N_24470,N_26520);
xnor U28496 (N_28496,N_25750,N_25808);
nand U28497 (N_28497,N_25014,N_25404);
xor U28498 (N_28498,N_26119,N_24196);
or U28499 (N_28499,N_26550,N_24408);
or U28500 (N_28500,N_24146,N_26379);
nor U28501 (N_28501,N_25071,N_24254);
nand U28502 (N_28502,N_24521,N_25127);
xnor U28503 (N_28503,N_25835,N_25690);
or U28504 (N_28504,N_24186,N_24963);
xor U28505 (N_28505,N_26877,N_26866);
nand U28506 (N_28506,N_24965,N_26728);
and U28507 (N_28507,N_25372,N_26401);
and U28508 (N_28508,N_24141,N_24648);
xor U28509 (N_28509,N_24474,N_25284);
nor U28510 (N_28510,N_25213,N_24328);
xor U28511 (N_28511,N_24171,N_26591);
or U28512 (N_28512,N_26443,N_26991);
xor U28513 (N_28513,N_25706,N_25186);
xor U28514 (N_28514,N_26459,N_24922);
and U28515 (N_28515,N_25323,N_26285);
or U28516 (N_28516,N_25915,N_26326);
nand U28517 (N_28517,N_25582,N_25044);
and U28518 (N_28518,N_25428,N_26611);
or U28519 (N_28519,N_24982,N_25629);
and U28520 (N_28520,N_26846,N_24933);
xnor U28521 (N_28521,N_24397,N_26414);
and U28522 (N_28522,N_24837,N_24180);
nor U28523 (N_28523,N_26233,N_25939);
xnor U28524 (N_28524,N_26399,N_24293);
and U28525 (N_28525,N_26345,N_25633);
nor U28526 (N_28526,N_25696,N_26738);
nand U28527 (N_28527,N_25839,N_25971);
xnor U28528 (N_28528,N_25191,N_25620);
nand U28529 (N_28529,N_24558,N_24466);
nand U28530 (N_28530,N_26605,N_24331);
and U28531 (N_28531,N_24806,N_26875);
nor U28532 (N_28532,N_24656,N_25976);
xnor U28533 (N_28533,N_25074,N_25786);
nand U28534 (N_28534,N_24079,N_26300);
and U28535 (N_28535,N_24128,N_26102);
or U28536 (N_28536,N_25005,N_24594);
nand U28537 (N_28537,N_24018,N_25802);
nor U28538 (N_28538,N_25333,N_26282);
and U28539 (N_28539,N_24006,N_25282);
xor U28540 (N_28540,N_24278,N_25644);
nor U28541 (N_28541,N_24979,N_25016);
and U28542 (N_28542,N_26780,N_24714);
nand U28543 (N_28543,N_24129,N_26895);
xor U28544 (N_28544,N_25232,N_26548);
xnor U28545 (N_28545,N_25166,N_26323);
nand U28546 (N_28546,N_24106,N_25214);
and U28547 (N_28547,N_25302,N_26436);
nand U28548 (N_28548,N_26518,N_24717);
and U28549 (N_28549,N_26964,N_24988);
nor U28550 (N_28550,N_24880,N_25348);
xor U28551 (N_28551,N_26931,N_26244);
xor U28552 (N_28552,N_24869,N_26434);
or U28553 (N_28553,N_26391,N_24646);
nor U28554 (N_28554,N_26120,N_24235);
and U28555 (N_28555,N_25724,N_25433);
and U28556 (N_28556,N_26640,N_24235);
xor U28557 (N_28557,N_25507,N_25893);
nand U28558 (N_28558,N_24804,N_25618);
xnor U28559 (N_28559,N_25712,N_26650);
and U28560 (N_28560,N_26360,N_25335);
xnor U28561 (N_28561,N_24447,N_26454);
xnor U28562 (N_28562,N_25178,N_26162);
xnor U28563 (N_28563,N_26707,N_25563);
nand U28564 (N_28564,N_24948,N_25241);
xnor U28565 (N_28565,N_25860,N_26333);
or U28566 (N_28566,N_24627,N_25943);
nor U28567 (N_28567,N_26646,N_26180);
nand U28568 (N_28568,N_24174,N_25308);
or U28569 (N_28569,N_25209,N_25814);
nor U28570 (N_28570,N_25102,N_26840);
xnor U28571 (N_28571,N_24751,N_26398);
or U28572 (N_28572,N_24871,N_25378);
xor U28573 (N_28573,N_26594,N_24220);
nor U28574 (N_28574,N_25245,N_25201);
or U28575 (N_28575,N_26390,N_26606);
nor U28576 (N_28576,N_26423,N_24759);
and U28577 (N_28577,N_25912,N_24402);
or U28578 (N_28578,N_24861,N_25002);
and U28579 (N_28579,N_24097,N_24539);
and U28580 (N_28580,N_24996,N_26756);
and U28581 (N_28581,N_25628,N_26638);
and U28582 (N_28582,N_25987,N_26155);
nand U28583 (N_28583,N_24998,N_25590);
nand U28584 (N_28584,N_24289,N_26416);
xor U28585 (N_28585,N_26319,N_25797);
xnor U28586 (N_28586,N_25860,N_25152);
or U28587 (N_28587,N_25545,N_25286);
and U28588 (N_28588,N_24280,N_25133);
nand U28589 (N_28589,N_26868,N_25777);
and U28590 (N_28590,N_24949,N_24035);
nor U28591 (N_28591,N_26650,N_26505);
or U28592 (N_28592,N_24727,N_25944);
xnor U28593 (N_28593,N_25414,N_24436);
nor U28594 (N_28594,N_25410,N_25710);
or U28595 (N_28595,N_26759,N_26184);
or U28596 (N_28596,N_24384,N_24463);
nor U28597 (N_28597,N_25237,N_25098);
nor U28598 (N_28598,N_24138,N_24237);
or U28599 (N_28599,N_25862,N_25045);
or U28600 (N_28600,N_25843,N_25935);
nor U28601 (N_28601,N_25607,N_26523);
or U28602 (N_28602,N_25976,N_24910);
nor U28603 (N_28603,N_24384,N_26821);
and U28604 (N_28604,N_26753,N_25519);
nor U28605 (N_28605,N_25740,N_26828);
nand U28606 (N_28606,N_24782,N_24398);
or U28607 (N_28607,N_26558,N_24995);
and U28608 (N_28608,N_24638,N_26061);
nand U28609 (N_28609,N_24980,N_25921);
nor U28610 (N_28610,N_26981,N_25978);
and U28611 (N_28611,N_26237,N_24846);
nand U28612 (N_28612,N_24273,N_25333);
or U28613 (N_28613,N_24617,N_26066);
or U28614 (N_28614,N_25971,N_26843);
nand U28615 (N_28615,N_26083,N_26358);
nand U28616 (N_28616,N_24874,N_24226);
nand U28617 (N_28617,N_24804,N_26364);
nor U28618 (N_28618,N_25411,N_24214);
nor U28619 (N_28619,N_24683,N_24590);
nand U28620 (N_28620,N_24950,N_26179);
and U28621 (N_28621,N_24117,N_26376);
and U28622 (N_28622,N_25578,N_26764);
nand U28623 (N_28623,N_26688,N_26894);
and U28624 (N_28624,N_24651,N_24442);
nand U28625 (N_28625,N_25875,N_25207);
nand U28626 (N_28626,N_25394,N_24511);
xnor U28627 (N_28627,N_26794,N_25583);
nor U28628 (N_28628,N_26025,N_26093);
and U28629 (N_28629,N_24650,N_25742);
or U28630 (N_28630,N_26707,N_26404);
and U28631 (N_28631,N_25398,N_25597);
nand U28632 (N_28632,N_26993,N_25411);
nand U28633 (N_28633,N_26709,N_25671);
and U28634 (N_28634,N_25072,N_25093);
nor U28635 (N_28635,N_25449,N_25695);
or U28636 (N_28636,N_24604,N_25424);
or U28637 (N_28637,N_26008,N_25239);
xor U28638 (N_28638,N_24752,N_24259);
nor U28639 (N_28639,N_26027,N_25761);
and U28640 (N_28640,N_24584,N_24948);
or U28641 (N_28641,N_24617,N_25733);
nand U28642 (N_28642,N_25153,N_24126);
and U28643 (N_28643,N_24475,N_25090);
xnor U28644 (N_28644,N_26485,N_26135);
or U28645 (N_28645,N_24366,N_26391);
nor U28646 (N_28646,N_26921,N_26186);
and U28647 (N_28647,N_26439,N_26502);
nor U28648 (N_28648,N_24539,N_25620);
xor U28649 (N_28649,N_26530,N_25978);
and U28650 (N_28650,N_25201,N_24677);
nand U28651 (N_28651,N_26626,N_24356);
and U28652 (N_28652,N_26629,N_24326);
xnor U28653 (N_28653,N_25378,N_25408);
and U28654 (N_28654,N_26794,N_26705);
and U28655 (N_28655,N_26103,N_24853);
nand U28656 (N_28656,N_25919,N_26664);
or U28657 (N_28657,N_25257,N_26033);
or U28658 (N_28658,N_25485,N_25785);
nand U28659 (N_28659,N_24101,N_25008);
nor U28660 (N_28660,N_24933,N_24448);
nand U28661 (N_28661,N_26910,N_24234);
nand U28662 (N_28662,N_25344,N_25125);
and U28663 (N_28663,N_24676,N_24915);
nand U28664 (N_28664,N_25674,N_25585);
nand U28665 (N_28665,N_24742,N_24441);
nand U28666 (N_28666,N_24729,N_25100);
nand U28667 (N_28667,N_24148,N_24102);
or U28668 (N_28668,N_26484,N_24343);
nor U28669 (N_28669,N_24177,N_26784);
or U28670 (N_28670,N_24146,N_24302);
or U28671 (N_28671,N_26009,N_24111);
xnor U28672 (N_28672,N_26030,N_25241);
nor U28673 (N_28673,N_26444,N_26139);
and U28674 (N_28674,N_26148,N_25515);
nor U28675 (N_28675,N_25317,N_26411);
and U28676 (N_28676,N_26696,N_24621);
xnor U28677 (N_28677,N_26545,N_26698);
and U28678 (N_28678,N_26488,N_26337);
and U28679 (N_28679,N_25557,N_26478);
nor U28680 (N_28680,N_25904,N_26016);
nand U28681 (N_28681,N_25645,N_25931);
and U28682 (N_28682,N_26139,N_24373);
and U28683 (N_28683,N_26275,N_25264);
nand U28684 (N_28684,N_24092,N_25265);
and U28685 (N_28685,N_26976,N_24088);
nor U28686 (N_28686,N_24159,N_25928);
nand U28687 (N_28687,N_25308,N_24564);
nor U28688 (N_28688,N_24394,N_26427);
xor U28689 (N_28689,N_25364,N_24585);
nor U28690 (N_28690,N_25139,N_26658);
and U28691 (N_28691,N_26809,N_26640);
nor U28692 (N_28692,N_26391,N_24527);
and U28693 (N_28693,N_25087,N_25723);
and U28694 (N_28694,N_24057,N_26058);
nor U28695 (N_28695,N_24464,N_25759);
nand U28696 (N_28696,N_25529,N_24488);
and U28697 (N_28697,N_24200,N_25464);
or U28698 (N_28698,N_26270,N_26468);
and U28699 (N_28699,N_26646,N_25498);
xnor U28700 (N_28700,N_25521,N_26371);
nand U28701 (N_28701,N_24029,N_24898);
and U28702 (N_28702,N_24150,N_25649);
and U28703 (N_28703,N_26724,N_26763);
and U28704 (N_28704,N_25352,N_26376);
or U28705 (N_28705,N_26369,N_25024);
xor U28706 (N_28706,N_26156,N_26399);
and U28707 (N_28707,N_24698,N_24037);
or U28708 (N_28708,N_24543,N_25102);
xnor U28709 (N_28709,N_24347,N_26351);
and U28710 (N_28710,N_25509,N_25752);
xor U28711 (N_28711,N_24419,N_26032);
or U28712 (N_28712,N_25221,N_24159);
or U28713 (N_28713,N_24031,N_25662);
nor U28714 (N_28714,N_26058,N_26556);
and U28715 (N_28715,N_26339,N_24552);
nand U28716 (N_28716,N_25422,N_24561);
nand U28717 (N_28717,N_24585,N_24548);
xor U28718 (N_28718,N_26771,N_26587);
nor U28719 (N_28719,N_26387,N_24722);
and U28720 (N_28720,N_26830,N_26129);
or U28721 (N_28721,N_24887,N_25304);
nor U28722 (N_28722,N_26365,N_24880);
nor U28723 (N_28723,N_25905,N_24653);
nand U28724 (N_28724,N_24839,N_26585);
nand U28725 (N_28725,N_26133,N_25315);
nand U28726 (N_28726,N_25342,N_26528);
or U28727 (N_28727,N_26010,N_26317);
and U28728 (N_28728,N_26406,N_26869);
and U28729 (N_28729,N_24388,N_24659);
or U28730 (N_28730,N_26767,N_25066);
and U28731 (N_28731,N_24020,N_24961);
xnor U28732 (N_28732,N_24114,N_24041);
nor U28733 (N_28733,N_25167,N_24232);
nand U28734 (N_28734,N_26031,N_25759);
xnor U28735 (N_28735,N_26024,N_25595);
nand U28736 (N_28736,N_24740,N_25084);
and U28737 (N_28737,N_26208,N_25883);
xnor U28738 (N_28738,N_26594,N_24654);
or U28739 (N_28739,N_26016,N_26715);
xor U28740 (N_28740,N_24344,N_25602);
and U28741 (N_28741,N_25986,N_25466);
nor U28742 (N_28742,N_25346,N_25296);
nand U28743 (N_28743,N_24591,N_24534);
xor U28744 (N_28744,N_24203,N_25405);
and U28745 (N_28745,N_24931,N_25674);
xnor U28746 (N_28746,N_24629,N_25117);
or U28747 (N_28747,N_24806,N_24239);
or U28748 (N_28748,N_26084,N_26940);
nand U28749 (N_28749,N_26895,N_24699);
nand U28750 (N_28750,N_25050,N_25939);
nand U28751 (N_28751,N_25999,N_25396);
xnor U28752 (N_28752,N_25141,N_26749);
nand U28753 (N_28753,N_26818,N_26046);
xor U28754 (N_28754,N_26561,N_26982);
xnor U28755 (N_28755,N_25758,N_25878);
nor U28756 (N_28756,N_25715,N_25287);
xor U28757 (N_28757,N_25219,N_25189);
nand U28758 (N_28758,N_25039,N_26061);
and U28759 (N_28759,N_26139,N_26114);
nand U28760 (N_28760,N_26361,N_26493);
and U28761 (N_28761,N_24711,N_24063);
xor U28762 (N_28762,N_24184,N_26695);
nor U28763 (N_28763,N_24923,N_24410);
nor U28764 (N_28764,N_26493,N_25516);
or U28765 (N_28765,N_24260,N_26837);
nor U28766 (N_28766,N_26116,N_26041);
xnor U28767 (N_28767,N_24502,N_24018);
xor U28768 (N_28768,N_25693,N_25041);
nand U28769 (N_28769,N_25899,N_26404);
or U28770 (N_28770,N_24939,N_25388);
nand U28771 (N_28771,N_25228,N_25456);
or U28772 (N_28772,N_25223,N_24879);
xnor U28773 (N_28773,N_24355,N_25737);
nand U28774 (N_28774,N_25843,N_24511);
and U28775 (N_28775,N_24561,N_26000);
xor U28776 (N_28776,N_25357,N_24762);
nand U28777 (N_28777,N_25328,N_24309);
and U28778 (N_28778,N_26824,N_25098);
xor U28779 (N_28779,N_26400,N_25589);
or U28780 (N_28780,N_25011,N_26914);
xor U28781 (N_28781,N_26003,N_24100);
nor U28782 (N_28782,N_24920,N_26545);
or U28783 (N_28783,N_24305,N_26109);
nor U28784 (N_28784,N_25235,N_26965);
xor U28785 (N_28785,N_25376,N_24696);
xor U28786 (N_28786,N_26488,N_24940);
xnor U28787 (N_28787,N_25022,N_24493);
and U28788 (N_28788,N_25369,N_25433);
and U28789 (N_28789,N_24566,N_26627);
nor U28790 (N_28790,N_24649,N_26500);
nand U28791 (N_28791,N_26445,N_25321);
nor U28792 (N_28792,N_25823,N_24568);
nand U28793 (N_28793,N_26987,N_25691);
and U28794 (N_28794,N_25851,N_24128);
nor U28795 (N_28795,N_24611,N_26370);
or U28796 (N_28796,N_26241,N_26239);
or U28797 (N_28797,N_26227,N_25478);
and U28798 (N_28798,N_24835,N_26238);
and U28799 (N_28799,N_25251,N_26508);
and U28800 (N_28800,N_26782,N_25977);
and U28801 (N_28801,N_26263,N_26919);
and U28802 (N_28802,N_24759,N_26227);
nor U28803 (N_28803,N_24195,N_26598);
nor U28804 (N_28804,N_24278,N_26553);
nand U28805 (N_28805,N_24958,N_24444);
or U28806 (N_28806,N_24283,N_25398);
nand U28807 (N_28807,N_24982,N_24838);
xor U28808 (N_28808,N_25018,N_25403);
or U28809 (N_28809,N_26879,N_26195);
xor U28810 (N_28810,N_26900,N_26477);
nand U28811 (N_28811,N_25248,N_25421);
and U28812 (N_28812,N_25389,N_24668);
xor U28813 (N_28813,N_26459,N_25912);
or U28814 (N_28814,N_26914,N_24462);
or U28815 (N_28815,N_26476,N_26061);
and U28816 (N_28816,N_26085,N_25133);
or U28817 (N_28817,N_24474,N_25835);
or U28818 (N_28818,N_25280,N_24393);
nor U28819 (N_28819,N_24214,N_25445);
and U28820 (N_28820,N_24700,N_25637);
and U28821 (N_28821,N_25891,N_24835);
nand U28822 (N_28822,N_26123,N_26959);
xnor U28823 (N_28823,N_24077,N_24151);
or U28824 (N_28824,N_26081,N_26084);
xnor U28825 (N_28825,N_24168,N_24159);
or U28826 (N_28826,N_25111,N_26793);
xor U28827 (N_28827,N_24875,N_25315);
or U28828 (N_28828,N_26910,N_26744);
or U28829 (N_28829,N_24719,N_26685);
nor U28830 (N_28830,N_26580,N_24972);
or U28831 (N_28831,N_25610,N_25547);
nand U28832 (N_28832,N_24793,N_26898);
nand U28833 (N_28833,N_25525,N_24850);
xor U28834 (N_28834,N_25206,N_26162);
xor U28835 (N_28835,N_26249,N_25157);
nand U28836 (N_28836,N_26248,N_26882);
or U28837 (N_28837,N_24291,N_26984);
nand U28838 (N_28838,N_24586,N_24849);
xnor U28839 (N_28839,N_24718,N_25140);
nand U28840 (N_28840,N_26416,N_24395);
nand U28841 (N_28841,N_24989,N_25414);
nor U28842 (N_28842,N_26267,N_25858);
xor U28843 (N_28843,N_24393,N_24823);
nand U28844 (N_28844,N_25097,N_24291);
or U28845 (N_28845,N_26122,N_25505);
nand U28846 (N_28846,N_25974,N_26193);
xnor U28847 (N_28847,N_26610,N_26936);
nor U28848 (N_28848,N_24690,N_26398);
or U28849 (N_28849,N_26018,N_26084);
nand U28850 (N_28850,N_25194,N_25821);
or U28851 (N_28851,N_26667,N_24692);
or U28852 (N_28852,N_26277,N_25557);
xnor U28853 (N_28853,N_25485,N_26021);
and U28854 (N_28854,N_24999,N_24945);
xor U28855 (N_28855,N_26714,N_25164);
nand U28856 (N_28856,N_24129,N_25880);
and U28857 (N_28857,N_25295,N_25620);
nor U28858 (N_28858,N_25993,N_26286);
xnor U28859 (N_28859,N_25932,N_24705);
nor U28860 (N_28860,N_26230,N_25317);
nand U28861 (N_28861,N_25014,N_26821);
or U28862 (N_28862,N_25645,N_24922);
nor U28863 (N_28863,N_25948,N_26897);
and U28864 (N_28864,N_24708,N_24934);
nand U28865 (N_28865,N_26390,N_25604);
and U28866 (N_28866,N_26112,N_26013);
nand U28867 (N_28867,N_24121,N_25790);
or U28868 (N_28868,N_25261,N_24693);
xor U28869 (N_28869,N_24988,N_25693);
or U28870 (N_28870,N_24534,N_25339);
or U28871 (N_28871,N_24793,N_24089);
xor U28872 (N_28872,N_25790,N_24377);
nand U28873 (N_28873,N_24916,N_24725);
and U28874 (N_28874,N_26898,N_25668);
and U28875 (N_28875,N_25338,N_26316);
or U28876 (N_28876,N_24987,N_26378);
xor U28877 (N_28877,N_25917,N_25143);
or U28878 (N_28878,N_25261,N_24288);
or U28879 (N_28879,N_26494,N_24446);
or U28880 (N_28880,N_26205,N_24812);
and U28881 (N_28881,N_26163,N_26356);
nand U28882 (N_28882,N_24873,N_24234);
or U28883 (N_28883,N_25536,N_26281);
nor U28884 (N_28884,N_25151,N_26922);
xnor U28885 (N_28885,N_26100,N_26140);
and U28886 (N_28886,N_25627,N_24151);
and U28887 (N_28887,N_25282,N_24597);
nand U28888 (N_28888,N_24386,N_24195);
nor U28889 (N_28889,N_26544,N_24871);
xnor U28890 (N_28890,N_26540,N_24056);
xor U28891 (N_28891,N_26472,N_25571);
and U28892 (N_28892,N_26943,N_25482);
nand U28893 (N_28893,N_26188,N_25363);
or U28894 (N_28894,N_25027,N_24183);
and U28895 (N_28895,N_24855,N_26890);
or U28896 (N_28896,N_26283,N_25913);
xnor U28897 (N_28897,N_24648,N_24798);
or U28898 (N_28898,N_26520,N_25501);
and U28899 (N_28899,N_24802,N_25297);
nor U28900 (N_28900,N_26018,N_24911);
nand U28901 (N_28901,N_26718,N_26796);
nor U28902 (N_28902,N_25365,N_24407);
xor U28903 (N_28903,N_24248,N_25955);
xnor U28904 (N_28904,N_24915,N_24921);
nor U28905 (N_28905,N_24140,N_26937);
xor U28906 (N_28906,N_24133,N_26909);
xnor U28907 (N_28907,N_26570,N_26402);
nand U28908 (N_28908,N_24021,N_24747);
or U28909 (N_28909,N_25342,N_24325);
xor U28910 (N_28910,N_26530,N_26261);
and U28911 (N_28911,N_25587,N_26877);
or U28912 (N_28912,N_24964,N_24042);
and U28913 (N_28913,N_25015,N_24922);
or U28914 (N_28914,N_24809,N_24485);
or U28915 (N_28915,N_24568,N_24865);
nand U28916 (N_28916,N_25309,N_24427);
or U28917 (N_28917,N_24656,N_26232);
nand U28918 (N_28918,N_25286,N_25935);
nor U28919 (N_28919,N_26722,N_25180);
xor U28920 (N_28920,N_26977,N_24513);
or U28921 (N_28921,N_26159,N_24099);
nor U28922 (N_28922,N_24449,N_26570);
xnor U28923 (N_28923,N_25083,N_24366);
and U28924 (N_28924,N_25101,N_25728);
or U28925 (N_28925,N_26085,N_26423);
and U28926 (N_28926,N_24317,N_25525);
nand U28927 (N_28927,N_24825,N_26747);
and U28928 (N_28928,N_25886,N_26322);
nand U28929 (N_28929,N_24482,N_26537);
or U28930 (N_28930,N_25520,N_25367);
nor U28931 (N_28931,N_24779,N_26635);
nor U28932 (N_28932,N_24313,N_24391);
nand U28933 (N_28933,N_26928,N_26884);
nand U28934 (N_28934,N_26073,N_24570);
nand U28935 (N_28935,N_25373,N_25150);
xor U28936 (N_28936,N_24321,N_24894);
nand U28937 (N_28937,N_26235,N_26110);
xor U28938 (N_28938,N_26216,N_24049);
nor U28939 (N_28939,N_26100,N_25000);
or U28940 (N_28940,N_26488,N_26757);
or U28941 (N_28941,N_25206,N_24706);
nor U28942 (N_28942,N_25005,N_25665);
nor U28943 (N_28943,N_25313,N_24694);
nand U28944 (N_28944,N_26734,N_26230);
nand U28945 (N_28945,N_24481,N_24894);
xnor U28946 (N_28946,N_25206,N_25118);
or U28947 (N_28947,N_24112,N_25706);
nand U28948 (N_28948,N_26567,N_24460);
xnor U28949 (N_28949,N_26695,N_26200);
and U28950 (N_28950,N_24705,N_24591);
nand U28951 (N_28951,N_25771,N_26929);
xnor U28952 (N_28952,N_25109,N_25102);
nor U28953 (N_28953,N_25756,N_24540);
xnor U28954 (N_28954,N_24242,N_25985);
xor U28955 (N_28955,N_25157,N_26986);
nand U28956 (N_28956,N_24314,N_26948);
nor U28957 (N_28957,N_25435,N_26037);
and U28958 (N_28958,N_24912,N_26876);
nor U28959 (N_28959,N_25238,N_26111);
nand U28960 (N_28960,N_25150,N_25313);
nor U28961 (N_28961,N_25612,N_26632);
nand U28962 (N_28962,N_26395,N_26367);
xor U28963 (N_28963,N_24859,N_25487);
xnor U28964 (N_28964,N_25851,N_25518);
nor U28965 (N_28965,N_24421,N_24002);
nor U28966 (N_28966,N_26453,N_26721);
and U28967 (N_28967,N_25055,N_25753);
nor U28968 (N_28968,N_25900,N_24067);
nor U28969 (N_28969,N_26937,N_26659);
nand U28970 (N_28970,N_25843,N_26613);
or U28971 (N_28971,N_25623,N_25343);
xor U28972 (N_28972,N_24582,N_24190);
and U28973 (N_28973,N_24249,N_24818);
and U28974 (N_28974,N_25172,N_24649);
or U28975 (N_28975,N_24981,N_24985);
nor U28976 (N_28976,N_25417,N_26941);
nand U28977 (N_28977,N_25438,N_25199);
or U28978 (N_28978,N_24837,N_24594);
nor U28979 (N_28979,N_24806,N_25944);
and U28980 (N_28980,N_24321,N_25953);
nand U28981 (N_28981,N_24241,N_24041);
nor U28982 (N_28982,N_24674,N_24910);
xor U28983 (N_28983,N_26581,N_25667);
or U28984 (N_28984,N_24482,N_24530);
xnor U28985 (N_28985,N_24154,N_25819);
or U28986 (N_28986,N_25349,N_26786);
and U28987 (N_28987,N_25678,N_26312);
xor U28988 (N_28988,N_25094,N_26693);
nor U28989 (N_28989,N_25753,N_26029);
nor U28990 (N_28990,N_24353,N_26659);
nor U28991 (N_28991,N_25943,N_25350);
nand U28992 (N_28992,N_26135,N_26844);
and U28993 (N_28993,N_24778,N_26482);
and U28994 (N_28994,N_25194,N_24733);
xor U28995 (N_28995,N_26533,N_26682);
or U28996 (N_28996,N_26112,N_25091);
nor U28997 (N_28997,N_24158,N_26143);
xor U28998 (N_28998,N_25357,N_25976);
and U28999 (N_28999,N_24718,N_25450);
and U29000 (N_29000,N_24649,N_26687);
and U29001 (N_29001,N_25674,N_26380);
xor U29002 (N_29002,N_24849,N_25526);
and U29003 (N_29003,N_26092,N_26005);
nor U29004 (N_29004,N_26008,N_24413);
and U29005 (N_29005,N_25183,N_24291);
and U29006 (N_29006,N_26668,N_24501);
or U29007 (N_29007,N_24504,N_24935);
and U29008 (N_29008,N_25381,N_25681);
nand U29009 (N_29009,N_24195,N_24674);
nand U29010 (N_29010,N_26139,N_25956);
nand U29011 (N_29011,N_26128,N_24617);
and U29012 (N_29012,N_25203,N_26043);
nor U29013 (N_29013,N_24271,N_26643);
nor U29014 (N_29014,N_26010,N_24141);
and U29015 (N_29015,N_26157,N_26197);
and U29016 (N_29016,N_24906,N_26033);
and U29017 (N_29017,N_24719,N_25033);
xor U29018 (N_29018,N_25204,N_24116);
nor U29019 (N_29019,N_25675,N_26326);
xor U29020 (N_29020,N_25763,N_24045);
or U29021 (N_29021,N_24006,N_24280);
nand U29022 (N_29022,N_26931,N_26182);
nand U29023 (N_29023,N_25340,N_24027);
or U29024 (N_29024,N_26933,N_26857);
nand U29025 (N_29025,N_25605,N_24151);
nor U29026 (N_29026,N_25638,N_26792);
xnor U29027 (N_29027,N_25902,N_25916);
nand U29028 (N_29028,N_25390,N_24622);
nand U29029 (N_29029,N_24369,N_25099);
xnor U29030 (N_29030,N_26691,N_24214);
nand U29031 (N_29031,N_25312,N_24727);
nand U29032 (N_29032,N_25197,N_24045);
or U29033 (N_29033,N_24705,N_25108);
or U29034 (N_29034,N_25447,N_25150);
nand U29035 (N_29035,N_24941,N_24503);
nor U29036 (N_29036,N_24039,N_25395);
or U29037 (N_29037,N_25806,N_24667);
nand U29038 (N_29038,N_24358,N_24530);
nor U29039 (N_29039,N_26170,N_26891);
or U29040 (N_29040,N_24357,N_26744);
nand U29041 (N_29041,N_24665,N_26210);
nor U29042 (N_29042,N_24470,N_26930);
nor U29043 (N_29043,N_24002,N_25955);
or U29044 (N_29044,N_25107,N_25813);
and U29045 (N_29045,N_26765,N_24897);
xnor U29046 (N_29046,N_25407,N_26355);
and U29047 (N_29047,N_25779,N_24757);
and U29048 (N_29048,N_25565,N_24110);
and U29049 (N_29049,N_24989,N_25038);
xor U29050 (N_29050,N_26931,N_25835);
xor U29051 (N_29051,N_24572,N_26789);
nor U29052 (N_29052,N_24503,N_26769);
and U29053 (N_29053,N_24737,N_26632);
nand U29054 (N_29054,N_24376,N_26404);
or U29055 (N_29055,N_26309,N_24070);
nand U29056 (N_29056,N_26316,N_24691);
and U29057 (N_29057,N_26300,N_25424);
nand U29058 (N_29058,N_24903,N_25205);
or U29059 (N_29059,N_26939,N_25121);
xor U29060 (N_29060,N_25034,N_25723);
nand U29061 (N_29061,N_24651,N_24423);
xnor U29062 (N_29062,N_24104,N_25067);
and U29063 (N_29063,N_24716,N_24954);
nand U29064 (N_29064,N_24074,N_24300);
and U29065 (N_29065,N_24297,N_24425);
nand U29066 (N_29066,N_24126,N_24846);
nand U29067 (N_29067,N_26329,N_25406);
or U29068 (N_29068,N_25021,N_25642);
and U29069 (N_29069,N_25428,N_26684);
and U29070 (N_29070,N_24765,N_24613);
or U29071 (N_29071,N_26931,N_25290);
nor U29072 (N_29072,N_26101,N_26035);
or U29073 (N_29073,N_24675,N_25219);
nor U29074 (N_29074,N_24969,N_25710);
and U29075 (N_29075,N_24684,N_26295);
and U29076 (N_29076,N_25324,N_26976);
nor U29077 (N_29077,N_25357,N_24224);
nand U29078 (N_29078,N_24294,N_26249);
nand U29079 (N_29079,N_24195,N_25181);
or U29080 (N_29080,N_24076,N_24858);
xnor U29081 (N_29081,N_24433,N_26059);
and U29082 (N_29082,N_25715,N_24087);
nand U29083 (N_29083,N_26787,N_25783);
or U29084 (N_29084,N_25227,N_24783);
and U29085 (N_29085,N_26368,N_25244);
xor U29086 (N_29086,N_24811,N_26698);
nor U29087 (N_29087,N_25252,N_24770);
xor U29088 (N_29088,N_26756,N_24192);
xnor U29089 (N_29089,N_26466,N_26612);
and U29090 (N_29090,N_24289,N_25923);
or U29091 (N_29091,N_25779,N_24059);
nand U29092 (N_29092,N_26531,N_24240);
xor U29093 (N_29093,N_24534,N_26012);
nor U29094 (N_29094,N_24833,N_25885);
and U29095 (N_29095,N_24180,N_24652);
nand U29096 (N_29096,N_24696,N_25356);
or U29097 (N_29097,N_26980,N_26957);
xnor U29098 (N_29098,N_26684,N_24021);
and U29099 (N_29099,N_24981,N_24161);
or U29100 (N_29100,N_26101,N_25373);
nor U29101 (N_29101,N_24561,N_25216);
xor U29102 (N_29102,N_25097,N_24569);
or U29103 (N_29103,N_26895,N_26272);
and U29104 (N_29104,N_24415,N_24682);
xnor U29105 (N_29105,N_24233,N_25636);
or U29106 (N_29106,N_24589,N_25149);
or U29107 (N_29107,N_26322,N_25703);
and U29108 (N_29108,N_25633,N_26791);
xnor U29109 (N_29109,N_26764,N_25194);
and U29110 (N_29110,N_24175,N_24404);
nor U29111 (N_29111,N_26639,N_25872);
or U29112 (N_29112,N_26054,N_26346);
nor U29113 (N_29113,N_24252,N_25004);
xor U29114 (N_29114,N_24158,N_24560);
or U29115 (N_29115,N_24772,N_26782);
and U29116 (N_29116,N_24979,N_25228);
nand U29117 (N_29117,N_24704,N_26568);
xnor U29118 (N_29118,N_26160,N_24371);
nand U29119 (N_29119,N_26560,N_24398);
xor U29120 (N_29120,N_25027,N_26640);
nor U29121 (N_29121,N_25354,N_26053);
nand U29122 (N_29122,N_24256,N_24384);
and U29123 (N_29123,N_24857,N_24315);
xnor U29124 (N_29124,N_26344,N_25404);
and U29125 (N_29125,N_24813,N_26494);
nand U29126 (N_29126,N_24091,N_26814);
or U29127 (N_29127,N_25638,N_26772);
nand U29128 (N_29128,N_26278,N_24337);
nand U29129 (N_29129,N_26201,N_24816);
or U29130 (N_29130,N_25842,N_25827);
nor U29131 (N_29131,N_26422,N_24003);
nand U29132 (N_29132,N_24298,N_25969);
xor U29133 (N_29133,N_25125,N_25919);
nand U29134 (N_29134,N_25226,N_24489);
nor U29135 (N_29135,N_26134,N_26849);
xnor U29136 (N_29136,N_25252,N_24494);
or U29137 (N_29137,N_24925,N_25215);
or U29138 (N_29138,N_26220,N_26710);
xnor U29139 (N_29139,N_24695,N_24659);
nand U29140 (N_29140,N_26418,N_25463);
or U29141 (N_29141,N_25563,N_24848);
xnor U29142 (N_29142,N_24296,N_24986);
nand U29143 (N_29143,N_25965,N_25813);
and U29144 (N_29144,N_25564,N_26022);
or U29145 (N_29145,N_25488,N_26245);
and U29146 (N_29146,N_24058,N_24204);
nand U29147 (N_29147,N_26388,N_24327);
nand U29148 (N_29148,N_25829,N_24510);
nand U29149 (N_29149,N_24126,N_26523);
xnor U29150 (N_29150,N_24051,N_26423);
nor U29151 (N_29151,N_26097,N_26314);
and U29152 (N_29152,N_24198,N_24269);
nor U29153 (N_29153,N_24946,N_26835);
xor U29154 (N_29154,N_24590,N_26238);
xnor U29155 (N_29155,N_25317,N_26947);
or U29156 (N_29156,N_26503,N_25628);
and U29157 (N_29157,N_26373,N_26591);
nand U29158 (N_29158,N_26307,N_26445);
or U29159 (N_29159,N_25791,N_26168);
nand U29160 (N_29160,N_24720,N_25807);
and U29161 (N_29161,N_26806,N_25071);
nor U29162 (N_29162,N_25423,N_25864);
nand U29163 (N_29163,N_26937,N_26664);
and U29164 (N_29164,N_24948,N_25262);
nor U29165 (N_29165,N_24540,N_26464);
or U29166 (N_29166,N_25517,N_25415);
xnor U29167 (N_29167,N_25537,N_25249);
and U29168 (N_29168,N_24990,N_26029);
or U29169 (N_29169,N_25221,N_24096);
xor U29170 (N_29170,N_26364,N_25132);
xnor U29171 (N_29171,N_25109,N_24108);
nand U29172 (N_29172,N_25658,N_26220);
nor U29173 (N_29173,N_26095,N_26598);
nand U29174 (N_29174,N_24914,N_26973);
nor U29175 (N_29175,N_26410,N_25914);
nor U29176 (N_29176,N_24829,N_24956);
or U29177 (N_29177,N_26907,N_25105);
and U29178 (N_29178,N_26082,N_25130);
or U29179 (N_29179,N_24759,N_24183);
or U29180 (N_29180,N_26100,N_25375);
nor U29181 (N_29181,N_25680,N_25812);
nand U29182 (N_29182,N_24538,N_24888);
nor U29183 (N_29183,N_26333,N_25062);
xor U29184 (N_29184,N_26657,N_24330);
and U29185 (N_29185,N_26361,N_25497);
nor U29186 (N_29186,N_25329,N_24726);
and U29187 (N_29187,N_26072,N_24712);
and U29188 (N_29188,N_25494,N_26043);
nor U29189 (N_29189,N_26540,N_26788);
xor U29190 (N_29190,N_25340,N_24314);
nand U29191 (N_29191,N_24164,N_25552);
xor U29192 (N_29192,N_26623,N_24788);
nand U29193 (N_29193,N_25186,N_25564);
xor U29194 (N_29194,N_24384,N_26680);
nor U29195 (N_29195,N_25538,N_26310);
and U29196 (N_29196,N_24775,N_24593);
xor U29197 (N_29197,N_24442,N_25748);
or U29198 (N_29198,N_24167,N_25122);
xor U29199 (N_29199,N_24397,N_26821);
nor U29200 (N_29200,N_24770,N_26482);
and U29201 (N_29201,N_25398,N_26050);
and U29202 (N_29202,N_24725,N_26726);
or U29203 (N_29203,N_26754,N_26684);
and U29204 (N_29204,N_24796,N_25432);
nand U29205 (N_29205,N_25953,N_24686);
nor U29206 (N_29206,N_25020,N_26205);
xor U29207 (N_29207,N_24459,N_26059);
or U29208 (N_29208,N_26627,N_24788);
xor U29209 (N_29209,N_26045,N_26486);
nand U29210 (N_29210,N_25549,N_26711);
xnor U29211 (N_29211,N_25325,N_24927);
xnor U29212 (N_29212,N_26825,N_25728);
or U29213 (N_29213,N_26605,N_24085);
or U29214 (N_29214,N_24787,N_26940);
nand U29215 (N_29215,N_26040,N_26229);
xnor U29216 (N_29216,N_25436,N_25035);
and U29217 (N_29217,N_26190,N_26689);
nand U29218 (N_29218,N_24352,N_24381);
or U29219 (N_29219,N_26832,N_25919);
xnor U29220 (N_29220,N_26816,N_25713);
nand U29221 (N_29221,N_25344,N_26175);
and U29222 (N_29222,N_26968,N_25602);
or U29223 (N_29223,N_24545,N_26612);
nor U29224 (N_29224,N_25066,N_26745);
nand U29225 (N_29225,N_25129,N_24906);
and U29226 (N_29226,N_26063,N_26764);
and U29227 (N_29227,N_26820,N_26399);
or U29228 (N_29228,N_25777,N_25527);
or U29229 (N_29229,N_26750,N_25531);
or U29230 (N_29230,N_24541,N_24912);
or U29231 (N_29231,N_25671,N_25135);
nand U29232 (N_29232,N_26321,N_25149);
nand U29233 (N_29233,N_24517,N_25646);
xnor U29234 (N_29234,N_25441,N_24527);
nor U29235 (N_29235,N_26074,N_26739);
xnor U29236 (N_29236,N_25585,N_24297);
nor U29237 (N_29237,N_25113,N_26288);
xor U29238 (N_29238,N_25982,N_24089);
nand U29239 (N_29239,N_26546,N_25137);
and U29240 (N_29240,N_24269,N_24671);
xnor U29241 (N_29241,N_26509,N_25471);
or U29242 (N_29242,N_24628,N_25686);
nor U29243 (N_29243,N_26673,N_26385);
and U29244 (N_29244,N_26860,N_25171);
nand U29245 (N_29245,N_26728,N_24934);
nand U29246 (N_29246,N_26729,N_24413);
nor U29247 (N_29247,N_24341,N_24951);
and U29248 (N_29248,N_25651,N_26681);
nand U29249 (N_29249,N_25360,N_24287);
or U29250 (N_29250,N_25910,N_26920);
or U29251 (N_29251,N_24387,N_26612);
or U29252 (N_29252,N_25322,N_24539);
nand U29253 (N_29253,N_24453,N_24297);
or U29254 (N_29254,N_24787,N_24972);
xnor U29255 (N_29255,N_24682,N_26489);
nand U29256 (N_29256,N_26006,N_25557);
and U29257 (N_29257,N_26708,N_24626);
xor U29258 (N_29258,N_24631,N_24220);
nor U29259 (N_29259,N_26401,N_26922);
nor U29260 (N_29260,N_25096,N_24943);
nand U29261 (N_29261,N_26870,N_25905);
or U29262 (N_29262,N_26629,N_24351);
xnor U29263 (N_29263,N_25266,N_24324);
and U29264 (N_29264,N_26098,N_24561);
or U29265 (N_29265,N_24609,N_26407);
nand U29266 (N_29266,N_24801,N_26295);
xor U29267 (N_29267,N_24853,N_26228);
xnor U29268 (N_29268,N_25805,N_24910);
nand U29269 (N_29269,N_26103,N_26766);
or U29270 (N_29270,N_24665,N_26160);
xnor U29271 (N_29271,N_25890,N_25073);
xnor U29272 (N_29272,N_24364,N_25469);
nand U29273 (N_29273,N_26868,N_25415);
nand U29274 (N_29274,N_25630,N_25343);
or U29275 (N_29275,N_25539,N_26503);
nand U29276 (N_29276,N_25448,N_24173);
xnor U29277 (N_29277,N_24127,N_26078);
and U29278 (N_29278,N_25260,N_24505);
or U29279 (N_29279,N_26889,N_25309);
and U29280 (N_29280,N_24883,N_26632);
or U29281 (N_29281,N_25447,N_24609);
and U29282 (N_29282,N_24406,N_24664);
and U29283 (N_29283,N_25023,N_25631);
or U29284 (N_29284,N_26471,N_25849);
and U29285 (N_29285,N_25316,N_26557);
xor U29286 (N_29286,N_26897,N_24531);
or U29287 (N_29287,N_26695,N_26321);
xor U29288 (N_29288,N_25446,N_24391);
xor U29289 (N_29289,N_24763,N_24435);
or U29290 (N_29290,N_26958,N_25890);
or U29291 (N_29291,N_25270,N_25567);
xor U29292 (N_29292,N_25737,N_25493);
nor U29293 (N_29293,N_26479,N_25953);
xnor U29294 (N_29294,N_26767,N_25122);
xnor U29295 (N_29295,N_25750,N_25767);
xnor U29296 (N_29296,N_25198,N_24383);
nor U29297 (N_29297,N_25731,N_25566);
or U29298 (N_29298,N_24950,N_26404);
nor U29299 (N_29299,N_25511,N_26397);
nor U29300 (N_29300,N_26510,N_26718);
nand U29301 (N_29301,N_26142,N_26045);
and U29302 (N_29302,N_24132,N_24929);
or U29303 (N_29303,N_24461,N_24545);
and U29304 (N_29304,N_24156,N_26717);
nand U29305 (N_29305,N_25289,N_25914);
nand U29306 (N_29306,N_25053,N_26718);
xor U29307 (N_29307,N_25844,N_25256);
nand U29308 (N_29308,N_24635,N_24253);
or U29309 (N_29309,N_24689,N_24976);
or U29310 (N_29310,N_24732,N_26155);
nand U29311 (N_29311,N_26198,N_24798);
nand U29312 (N_29312,N_26840,N_24500);
nand U29313 (N_29313,N_26634,N_25537);
xnor U29314 (N_29314,N_26628,N_24709);
xnor U29315 (N_29315,N_25870,N_24538);
and U29316 (N_29316,N_25499,N_26269);
and U29317 (N_29317,N_26585,N_26434);
or U29318 (N_29318,N_25023,N_25185);
and U29319 (N_29319,N_24418,N_24325);
or U29320 (N_29320,N_24618,N_24600);
nor U29321 (N_29321,N_25702,N_24256);
xor U29322 (N_29322,N_24353,N_26025);
nor U29323 (N_29323,N_24669,N_25842);
nor U29324 (N_29324,N_26578,N_24312);
nor U29325 (N_29325,N_25893,N_25038);
xnor U29326 (N_29326,N_26229,N_25404);
and U29327 (N_29327,N_25271,N_25560);
xnor U29328 (N_29328,N_26490,N_25046);
nand U29329 (N_29329,N_25514,N_26586);
and U29330 (N_29330,N_24700,N_24677);
nand U29331 (N_29331,N_24062,N_26505);
nand U29332 (N_29332,N_25660,N_25248);
nand U29333 (N_29333,N_25477,N_25088);
nor U29334 (N_29334,N_26481,N_25936);
or U29335 (N_29335,N_26032,N_24700);
nand U29336 (N_29336,N_25386,N_26444);
nand U29337 (N_29337,N_26419,N_24132);
nand U29338 (N_29338,N_25651,N_25310);
nand U29339 (N_29339,N_24785,N_25824);
xor U29340 (N_29340,N_24935,N_25355);
nor U29341 (N_29341,N_25779,N_26013);
nor U29342 (N_29342,N_24365,N_25779);
xor U29343 (N_29343,N_24212,N_24256);
or U29344 (N_29344,N_24418,N_24328);
or U29345 (N_29345,N_24379,N_24332);
nand U29346 (N_29346,N_24570,N_25481);
or U29347 (N_29347,N_25694,N_26653);
xnor U29348 (N_29348,N_24195,N_26478);
nand U29349 (N_29349,N_26117,N_24756);
and U29350 (N_29350,N_26591,N_24223);
and U29351 (N_29351,N_24699,N_25996);
xnor U29352 (N_29352,N_26021,N_26195);
nand U29353 (N_29353,N_24034,N_26013);
xor U29354 (N_29354,N_26573,N_25154);
and U29355 (N_29355,N_25448,N_25340);
nor U29356 (N_29356,N_26547,N_24450);
xnor U29357 (N_29357,N_24685,N_26783);
nand U29358 (N_29358,N_25681,N_26432);
nand U29359 (N_29359,N_25754,N_24489);
xnor U29360 (N_29360,N_24302,N_26460);
or U29361 (N_29361,N_24691,N_25377);
or U29362 (N_29362,N_24968,N_25360);
nor U29363 (N_29363,N_25754,N_24465);
or U29364 (N_29364,N_24060,N_26697);
nor U29365 (N_29365,N_25709,N_25021);
or U29366 (N_29366,N_25918,N_26231);
nand U29367 (N_29367,N_25933,N_26574);
or U29368 (N_29368,N_24911,N_26547);
and U29369 (N_29369,N_26449,N_25828);
nand U29370 (N_29370,N_26816,N_26169);
xnor U29371 (N_29371,N_25183,N_26041);
nand U29372 (N_29372,N_24802,N_26953);
and U29373 (N_29373,N_25045,N_25057);
nor U29374 (N_29374,N_26100,N_25820);
or U29375 (N_29375,N_24555,N_26794);
xnor U29376 (N_29376,N_26916,N_26040);
and U29377 (N_29377,N_25144,N_26663);
or U29378 (N_29378,N_24287,N_24732);
nor U29379 (N_29379,N_25562,N_25365);
or U29380 (N_29380,N_26813,N_24639);
nand U29381 (N_29381,N_26436,N_26149);
and U29382 (N_29382,N_24958,N_26908);
nand U29383 (N_29383,N_24390,N_26132);
and U29384 (N_29384,N_26495,N_26990);
or U29385 (N_29385,N_24592,N_25722);
xnor U29386 (N_29386,N_25868,N_24025);
nor U29387 (N_29387,N_25354,N_25630);
or U29388 (N_29388,N_25541,N_24784);
xor U29389 (N_29389,N_24698,N_25866);
xor U29390 (N_29390,N_25861,N_24754);
or U29391 (N_29391,N_25288,N_25735);
and U29392 (N_29392,N_26186,N_25031);
and U29393 (N_29393,N_24723,N_26989);
xor U29394 (N_29394,N_24044,N_25846);
and U29395 (N_29395,N_25908,N_25809);
or U29396 (N_29396,N_26377,N_24369);
xnor U29397 (N_29397,N_24424,N_24134);
or U29398 (N_29398,N_26842,N_26348);
and U29399 (N_29399,N_24130,N_25766);
nor U29400 (N_29400,N_24086,N_24701);
xor U29401 (N_29401,N_26947,N_24361);
xnor U29402 (N_29402,N_24085,N_24158);
and U29403 (N_29403,N_24198,N_26470);
or U29404 (N_29404,N_26256,N_24294);
and U29405 (N_29405,N_24764,N_26643);
and U29406 (N_29406,N_25832,N_24690);
and U29407 (N_29407,N_26453,N_25048);
and U29408 (N_29408,N_24528,N_24649);
and U29409 (N_29409,N_24354,N_26915);
or U29410 (N_29410,N_25104,N_26968);
nand U29411 (N_29411,N_24944,N_24069);
xor U29412 (N_29412,N_26912,N_24646);
and U29413 (N_29413,N_25839,N_25411);
and U29414 (N_29414,N_24629,N_24042);
or U29415 (N_29415,N_25595,N_24825);
nand U29416 (N_29416,N_25059,N_24458);
or U29417 (N_29417,N_26797,N_24596);
or U29418 (N_29418,N_25815,N_25821);
nand U29419 (N_29419,N_24150,N_24779);
xor U29420 (N_29420,N_24518,N_24106);
xor U29421 (N_29421,N_24323,N_25318);
xor U29422 (N_29422,N_26875,N_24218);
xor U29423 (N_29423,N_24013,N_24342);
xor U29424 (N_29424,N_26315,N_24147);
xnor U29425 (N_29425,N_24582,N_24063);
or U29426 (N_29426,N_26254,N_25301);
nor U29427 (N_29427,N_25078,N_24224);
nor U29428 (N_29428,N_26743,N_24372);
nor U29429 (N_29429,N_24970,N_24802);
or U29430 (N_29430,N_24120,N_26364);
and U29431 (N_29431,N_24601,N_24723);
nor U29432 (N_29432,N_25958,N_26587);
nand U29433 (N_29433,N_26884,N_26064);
xnor U29434 (N_29434,N_24632,N_26672);
nor U29435 (N_29435,N_26603,N_24728);
xor U29436 (N_29436,N_26543,N_26386);
xor U29437 (N_29437,N_26577,N_26072);
or U29438 (N_29438,N_24706,N_24476);
nor U29439 (N_29439,N_24544,N_25058);
nor U29440 (N_29440,N_26794,N_24554);
and U29441 (N_29441,N_26107,N_26275);
and U29442 (N_29442,N_25322,N_25384);
and U29443 (N_29443,N_26163,N_25853);
and U29444 (N_29444,N_26538,N_24849);
nor U29445 (N_29445,N_24786,N_25050);
nand U29446 (N_29446,N_25686,N_25696);
nor U29447 (N_29447,N_24005,N_25940);
xor U29448 (N_29448,N_25489,N_26087);
xor U29449 (N_29449,N_24419,N_26743);
nand U29450 (N_29450,N_26692,N_24752);
or U29451 (N_29451,N_25654,N_24587);
xnor U29452 (N_29452,N_25381,N_24029);
nor U29453 (N_29453,N_24976,N_26078);
xnor U29454 (N_29454,N_25998,N_25322);
nand U29455 (N_29455,N_26583,N_24514);
nand U29456 (N_29456,N_24883,N_24406);
xnor U29457 (N_29457,N_25527,N_26687);
xor U29458 (N_29458,N_25564,N_25242);
and U29459 (N_29459,N_24172,N_26317);
nor U29460 (N_29460,N_24095,N_26739);
nor U29461 (N_29461,N_24605,N_24398);
or U29462 (N_29462,N_24863,N_24374);
and U29463 (N_29463,N_25777,N_24441);
or U29464 (N_29464,N_25992,N_26852);
nand U29465 (N_29465,N_25193,N_25554);
nor U29466 (N_29466,N_26205,N_26640);
nand U29467 (N_29467,N_26120,N_25906);
xnor U29468 (N_29468,N_24688,N_25189);
xnor U29469 (N_29469,N_24406,N_26930);
or U29470 (N_29470,N_26590,N_26699);
nor U29471 (N_29471,N_24582,N_25205);
nor U29472 (N_29472,N_25883,N_24694);
xor U29473 (N_29473,N_24479,N_24731);
xnor U29474 (N_29474,N_25190,N_26638);
xnor U29475 (N_29475,N_25745,N_24336);
or U29476 (N_29476,N_25014,N_24808);
xnor U29477 (N_29477,N_24506,N_25036);
nor U29478 (N_29478,N_25220,N_25170);
nand U29479 (N_29479,N_26040,N_26746);
or U29480 (N_29480,N_25045,N_24010);
nor U29481 (N_29481,N_26803,N_24842);
and U29482 (N_29482,N_25151,N_25236);
nor U29483 (N_29483,N_25931,N_26870);
and U29484 (N_29484,N_24345,N_25698);
and U29485 (N_29485,N_26804,N_26334);
or U29486 (N_29486,N_26719,N_24914);
and U29487 (N_29487,N_25560,N_26722);
and U29488 (N_29488,N_25316,N_26576);
nand U29489 (N_29489,N_25921,N_25636);
nor U29490 (N_29490,N_26617,N_26930);
and U29491 (N_29491,N_25244,N_24985);
nand U29492 (N_29492,N_24877,N_25883);
nand U29493 (N_29493,N_25411,N_25744);
or U29494 (N_29494,N_25476,N_26913);
nor U29495 (N_29495,N_25905,N_26242);
and U29496 (N_29496,N_26245,N_26301);
xnor U29497 (N_29497,N_26784,N_26924);
nand U29498 (N_29498,N_25634,N_25195);
nand U29499 (N_29499,N_26911,N_25048);
and U29500 (N_29500,N_24443,N_25033);
and U29501 (N_29501,N_26076,N_25148);
nor U29502 (N_29502,N_24778,N_25281);
or U29503 (N_29503,N_24656,N_26797);
nor U29504 (N_29504,N_24891,N_26187);
or U29505 (N_29505,N_24128,N_25506);
nor U29506 (N_29506,N_24186,N_24980);
nor U29507 (N_29507,N_26656,N_25573);
and U29508 (N_29508,N_24746,N_26404);
or U29509 (N_29509,N_26700,N_26272);
or U29510 (N_29510,N_24520,N_24922);
and U29511 (N_29511,N_24863,N_25856);
nor U29512 (N_29512,N_26620,N_25094);
nand U29513 (N_29513,N_25765,N_26504);
nor U29514 (N_29514,N_26596,N_25485);
xor U29515 (N_29515,N_24413,N_26352);
nand U29516 (N_29516,N_24139,N_25954);
and U29517 (N_29517,N_24533,N_26157);
nor U29518 (N_29518,N_26357,N_26582);
xnor U29519 (N_29519,N_25467,N_24577);
nor U29520 (N_29520,N_25811,N_26902);
nor U29521 (N_29521,N_25567,N_26699);
xor U29522 (N_29522,N_26516,N_26250);
xnor U29523 (N_29523,N_26872,N_26565);
or U29524 (N_29524,N_25569,N_25716);
or U29525 (N_29525,N_25264,N_25547);
nor U29526 (N_29526,N_25266,N_26000);
or U29527 (N_29527,N_25874,N_24900);
nor U29528 (N_29528,N_25731,N_26192);
nand U29529 (N_29529,N_25433,N_26416);
and U29530 (N_29530,N_24821,N_25948);
or U29531 (N_29531,N_26135,N_25804);
and U29532 (N_29532,N_25452,N_25096);
xnor U29533 (N_29533,N_24686,N_26937);
nand U29534 (N_29534,N_26643,N_25115);
nor U29535 (N_29535,N_26086,N_26820);
nor U29536 (N_29536,N_26753,N_24659);
and U29537 (N_29537,N_24427,N_25847);
nor U29538 (N_29538,N_26281,N_24188);
nand U29539 (N_29539,N_26279,N_26179);
nor U29540 (N_29540,N_26176,N_26516);
or U29541 (N_29541,N_26815,N_24157);
xor U29542 (N_29542,N_25334,N_24726);
nand U29543 (N_29543,N_25717,N_26300);
xnor U29544 (N_29544,N_25830,N_26265);
and U29545 (N_29545,N_24964,N_24139);
nand U29546 (N_29546,N_25488,N_25862);
and U29547 (N_29547,N_26964,N_26415);
nand U29548 (N_29548,N_26072,N_26190);
nand U29549 (N_29549,N_25992,N_26272);
xnor U29550 (N_29550,N_24137,N_25963);
and U29551 (N_29551,N_26426,N_26741);
nand U29552 (N_29552,N_24568,N_25476);
and U29553 (N_29553,N_24218,N_26634);
nor U29554 (N_29554,N_26255,N_24347);
and U29555 (N_29555,N_25952,N_26411);
nand U29556 (N_29556,N_25552,N_24079);
xor U29557 (N_29557,N_26609,N_24182);
nor U29558 (N_29558,N_24123,N_24773);
nor U29559 (N_29559,N_25549,N_26158);
nor U29560 (N_29560,N_24011,N_26434);
or U29561 (N_29561,N_26923,N_26979);
xnor U29562 (N_29562,N_24422,N_25510);
or U29563 (N_29563,N_25861,N_25783);
nand U29564 (N_29564,N_24690,N_25293);
and U29565 (N_29565,N_25718,N_26573);
nand U29566 (N_29566,N_24540,N_25699);
nand U29567 (N_29567,N_26528,N_25409);
and U29568 (N_29568,N_26206,N_24315);
xnor U29569 (N_29569,N_26848,N_26505);
nor U29570 (N_29570,N_24913,N_24467);
and U29571 (N_29571,N_24775,N_24659);
and U29572 (N_29572,N_24770,N_26496);
xor U29573 (N_29573,N_26064,N_26737);
xor U29574 (N_29574,N_24283,N_25498);
nand U29575 (N_29575,N_25841,N_26423);
nor U29576 (N_29576,N_24169,N_25790);
nor U29577 (N_29577,N_24373,N_26529);
xor U29578 (N_29578,N_25840,N_24307);
xor U29579 (N_29579,N_26106,N_24531);
and U29580 (N_29580,N_26706,N_26159);
xor U29581 (N_29581,N_26552,N_25973);
nor U29582 (N_29582,N_26489,N_24681);
or U29583 (N_29583,N_24030,N_25830);
or U29584 (N_29584,N_26029,N_25700);
nor U29585 (N_29585,N_24662,N_24669);
and U29586 (N_29586,N_25208,N_26746);
and U29587 (N_29587,N_26047,N_25710);
or U29588 (N_29588,N_24021,N_26973);
nor U29589 (N_29589,N_24322,N_25015);
nor U29590 (N_29590,N_24107,N_24855);
or U29591 (N_29591,N_25634,N_26183);
and U29592 (N_29592,N_25544,N_25844);
nor U29593 (N_29593,N_25298,N_24568);
nor U29594 (N_29594,N_26150,N_25352);
xor U29595 (N_29595,N_26734,N_26501);
nor U29596 (N_29596,N_24979,N_24919);
and U29597 (N_29597,N_25532,N_26604);
and U29598 (N_29598,N_24627,N_25302);
nand U29599 (N_29599,N_25370,N_24861);
or U29600 (N_29600,N_26882,N_24089);
or U29601 (N_29601,N_24791,N_24895);
or U29602 (N_29602,N_24281,N_24112);
nand U29603 (N_29603,N_25288,N_25404);
nor U29604 (N_29604,N_26121,N_24051);
nand U29605 (N_29605,N_25630,N_26057);
nand U29606 (N_29606,N_26099,N_24109);
xor U29607 (N_29607,N_24296,N_25182);
or U29608 (N_29608,N_25841,N_24414);
or U29609 (N_29609,N_24801,N_26252);
nor U29610 (N_29610,N_26784,N_24487);
nor U29611 (N_29611,N_25034,N_24121);
nand U29612 (N_29612,N_25408,N_26085);
nor U29613 (N_29613,N_26946,N_24897);
nand U29614 (N_29614,N_26730,N_24208);
nand U29615 (N_29615,N_26583,N_25739);
nand U29616 (N_29616,N_26397,N_26873);
nor U29617 (N_29617,N_24764,N_25394);
nand U29618 (N_29618,N_26065,N_24290);
nor U29619 (N_29619,N_25851,N_25981);
and U29620 (N_29620,N_25860,N_26746);
and U29621 (N_29621,N_26093,N_24017);
xor U29622 (N_29622,N_26828,N_24502);
nor U29623 (N_29623,N_25780,N_24833);
xor U29624 (N_29624,N_25369,N_24240);
xor U29625 (N_29625,N_25660,N_25000);
xor U29626 (N_29626,N_26840,N_24245);
xor U29627 (N_29627,N_26240,N_25810);
xor U29628 (N_29628,N_24030,N_25225);
xnor U29629 (N_29629,N_24573,N_25929);
nand U29630 (N_29630,N_26382,N_25300);
or U29631 (N_29631,N_26045,N_26575);
nor U29632 (N_29632,N_25345,N_26246);
nor U29633 (N_29633,N_24244,N_26800);
xor U29634 (N_29634,N_25789,N_26030);
nand U29635 (N_29635,N_24350,N_25487);
or U29636 (N_29636,N_24516,N_24314);
nand U29637 (N_29637,N_26704,N_24531);
nand U29638 (N_29638,N_25487,N_26891);
and U29639 (N_29639,N_26455,N_26933);
xor U29640 (N_29640,N_26603,N_25653);
nand U29641 (N_29641,N_26536,N_26616);
xnor U29642 (N_29642,N_24996,N_26999);
nand U29643 (N_29643,N_24421,N_24003);
nor U29644 (N_29644,N_24136,N_26357);
and U29645 (N_29645,N_26096,N_25799);
and U29646 (N_29646,N_26623,N_26179);
or U29647 (N_29647,N_26012,N_24046);
nand U29648 (N_29648,N_25588,N_26099);
and U29649 (N_29649,N_26207,N_24422);
or U29650 (N_29650,N_25050,N_26544);
nor U29651 (N_29651,N_24766,N_25705);
and U29652 (N_29652,N_26393,N_25192);
and U29653 (N_29653,N_25095,N_24724);
and U29654 (N_29654,N_25250,N_24684);
xnor U29655 (N_29655,N_26366,N_24084);
xor U29656 (N_29656,N_26965,N_25352);
and U29657 (N_29657,N_24129,N_25976);
nand U29658 (N_29658,N_26212,N_26433);
and U29659 (N_29659,N_26330,N_26437);
and U29660 (N_29660,N_26461,N_25519);
and U29661 (N_29661,N_24200,N_24394);
nor U29662 (N_29662,N_24191,N_26966);
nor U29663 (N_29663,N_25504,N_26701);
nor U29664 (N_29664,N_24499,N_24800);
and U29665 (N_29665,N_26307,N_24093);
nor U29666 (N_29666,N_26969,N_26694);
or U29667 (N_29667,N_26198,N_25646);
nand U29668 (N_29668,N_26891,N_25136);
nor U29669 (N_29669,N_26735,N_25906);
nor U29670 (N_29670,N_25493,N_26754);
xnor U29671 (N_29671,N_25408,N_24639);
and U29672 (N_29672,N_24302,N_26463);
nand U29673 (N_29673,N_26868,N_24123);
nand U29674 (N_29674,N_25991,N_26039);
xnor U29675 (N_29675,N_25916,N_26892);
nor U29676 (N_29676,N_24177,N_24514);
or U29677 (N_29677,N_26053,N_25751);
and U29678 (N_29678,N_24995,N_26471);
and U29679 (N_29679,N_24257,N_26167);
nor U29680 (N_29680,N_26122,N_25432);
nor U29681 (N_29681,N_26890,N_25164);
or U29682 (N_29682,N_24302,N_25047);
xnor U29683 (N_29683,N_24464,N_26771);
nand U29684 (N_29684,N_26240,N_26057);
and U29685 (N_29685,N_26039,N_25286);
nor U29686 (N_29686,N_24380,N_24193);
nor U29687 (N_29687,N_24886,N_25308);
or U29688 (N_29688,N_26213,N_24820);
nand U29689 (N_29689,N_25250,N_25069);
xnor U29690 (N_29690,N_25527,N_26909);
nand U29691 (N_29691,N_26731,N_24663);
nand U29692 (N_29692,N_24516,N_25497);
xnor U29693 (N_29693,N_25882,N_25136);
nor U29694 (N_29694,N_25971,N_25435);
or U29695 (N_29695,N_25327,N_25061);
and U29696 (N_29696,N_26685,N_24916);
xor U29697 (N_29697,N_25238,N_25783);
and U29698 (N_29698,N_26335,N_25805);
and U29699 (N_29699,N_24519,N_24359);
nand U29700 (N_29700,N_25217,N_26194);
and U29701 (N_29701,N_24905,N_26605);
and U29702 (N_29702,N_26663,N_25452);
nand U29703 (N_29703,N_25764,N_26077);
xor U29704 (N_29704,N_25239,N_25533);
or U29705 (N_29705,N_25904,N_24644);
and U29706 (N_29706,N_26408,N_26195);
nand U29707 (N_29707,N_24446,N_26152);
nand U29708 (N_29708,N_24401,N_26094);
and U29709 (N_29709,N_26029,N_25567);
or U29710 (N_29710,N_25898,N_25645);
and U29711 (N_29711,N_24306,N_26794);
nand U29712 (N_29712,N_25897,N_25016);
nand U29713 (N_29713,N_24090,N_24947);
or U29714 (N_29714,N_26811,N_26498);
and U29715 (N_29715,N_25408,N_25061);
and U29716 (N_29716,N_25553,N_24313);
nand U29717 (N_29717,N_24917,N_24037);
xnor U29718 (N_29718,N_24106,N_26317);
xnor U29719 (N_29719,N_24199,N_25464);
nor U29720 (N_29720,N_25744,N_24301);
nand U29721 (N_29721,N_25590,N_24545);
and U29722 (N_29722,N_24615,N_24321);
nor U29723 (N_29723,N_24476,N_24935);
xnor U29724 (N_29724,N_26274,N_26507);
nor U29725 (N_29725,N_24782,N_25153);
nor U29726 (N_29726,N_24435,N_26499);
or U29727 (N_29727,N_24837,N_26930);
nand U29728 (N_29728,N_25768,N_26379);
and U29729 (N_29729,N_26067,N_24736);
nor U29730 (N_29730,N_25246,N_24615);
xnor U29731 (N_29731,N_24590,N_25802);
nand U29732 (N_29732,N_24206,N_26144);
or U29733 (N_29733,N_26834,N_24521);
nor U29734 (N_29734,N_24666,N_24778);
or U29735 (N_29735,N_24735,N_24949);
or U29736 (N_29736,N_24956,N_24163);
nand U29737 (N_29737,N_24581,N_24298);
nor U29738 (N_29738,N_24355,N_26382);
nand U29739 (N_29739,N_25551,N_24777);
nand U29740 (N_29740,N_25539,N_24575);
and U29741 (N_29741,N_24661,N_26253);
nand U29742 (N_29742,N_25978,N_24875);
or U29743 (N_29743,N_26922,N_26056);
xor U29744 (N_29744,N_25646,N_25388);
nor U29745 (N_29745,N_25945,N_24200);
xor U29746 (N_29746,N_26889,N_26946);
xnor U29747 (N_29747,N_26129,N_25304);
and U29748 (N_29748,N_25441,N_26594);
and U29749 (N_29749,N_25720,N_24655);
or U29750 (N_29750,N_26154,N_26650);
nor U29751 (N_29751,N_24636,N_25661);
nand U29752 (N_29752,N_24900,N_25245);
nor U29753 (N_29753,N_26561,N_24478);
xor U29754 (N_29754,N_25388,N_25015);
nand U29755 (N_29755,N_26103,N_26759);
nand U29756 (N_29756,N_24675,N_25058);
xor U29757 (N_29757,N_24912,N_26043);
nor U29758 (N_29758,N_24733,N_25618);
and U29759 (N_29759,N_25303,N_26187);
and U29760 (N_29760,N_26100,N_26848);
xor U29761 (N_29761,N_25317,N_26196);
nand U29762 (N_29762,N_25778,N_26174);
xnor U29763 (N_29763,N_25935,N_25893);
or U29764 (N_29764,N_24683,N_26083);
nor U29765 (N_29765,N_24438,N_26603);
and U29766 (N_29766,N_25356,N_24613);
nand U29767 (N_29767,N_24444,N_25569);
nand U29768 (N_29768,N_26417,N_26161);
xnor U29769 (N_29769,N_26545,N_25369);
nand U29770 (N_29770,N_25475,N_24574);
nand U29771 (N_29771,N_25550,N_24820);
and U29772 (N_29772,N_24875,N_26908);
xnor U29773 (N_29773,N_24398,N_26696);
nor U29774 (N_29774,N_25293,N_25018);
or U29775 (N_29775,N_26302,N_24808);
xor U29776 (N_29776,N_26401,N_24506);
and U29777 (N_29777,N_25538,N_24676);
nor U29778 (N_29778,N_26592,N_25552);
and U29779 (N_29779,N_24179,N_26301);
xor U29780 (N_29780,N_25648,N_25315);
xor U29781 (N_29781,N_25935,N_25837);
nor U29782 (N_29782,N_24204,N_25179);
xor U29783 (N_29783,N_24856,N_25809);
nor U29784 (N_29784,N_25836,N_25152);
nor U29785 (N_29785,N_24253,N_26417);
xnor U29786 (N_29786,N_26408,N_26128);
nand U29787 (N_29787,N_26002,N_25230);
or U29788 (N_29788,N_25366,N_24869);
or U29789 (N_29789,N_24750,N_25871);
nand U29790 (N_29790,N_25201,N_24676);
nor U29791 (N_29791,N_25581,N_26548);
nor U29792 (N_29792,N_25933,N_24623);
or U29793 (N_29793,N_25787,N_25979);
nand U29794 (N_29794,N_24563,N_24778);
and U29795 (N_29795,N_24794,N_24195);
xor U29796 (N_29796,N_26565,N_25186);
or U29797 (N_29797,N_26071,N_25923);
xnor U29798 (N_29798,N_25394,N_26696);
xnor U29799 (N_29799,N_24041,N_26945);
nand U29800 (N_29800,N_24671,N_24499);
or U29801 (N_29801,N_26493,N_25682);
and U29802 (N_29802,N_24504,N_26565);
and U29803 (N_29803,N_26733,N_25057);
xor U29804 (N_29804,N_25316,N_25629);
nor U29805 (N_29805,N_26612,N_24668);
or U29806 (N_29806,N_26566,N_24990);
or U29807 (N_29807,N_26574,N_26674);
nor U29808 (N_29808,N_24691,N_24024);
and U29809 (N_29809,N_24547,N_24577);
and U29810 (N_29810,N_25112,N_26680);
and U29811 (N_29811,N_26944,N_25190);
and U29812 (N_29812,N_26387,N_25058);
or U29813 (N_29813,N_26443,N_24574);
nor U29814 (N_29814,N_24839,N_25913);
nand U29815 (N_29815,N_26530,N_26385);
nor U29816 (N_29816,N_24142,N_26441);
nand U29817 (N_29817,N_24340,N_26792);
xnor U29818 (N_29818,N_24557,N_25789);
or U29819 (N_29819,N_26830,N_26382);
and U29820 (N_29820,N_24292,N_24761);
and U29821 (N_29821,N_25473,N_24511);
xnor U29822 (N_29822,N_26346,N_26235);
and U29823 (N_29823,N_24427,N_24214);
nor U29824 (N_29824,N_25477,N_24593);
or U29825 (N_29825,N_26130,N_24000);
nor U29826 (N_29826,N_24142,N_24036);
xor U29827 (N_29827,N_25033,N_24203);
and U29828 (N_29828,N_25366,N_24935);
nand U29829 (N_29829,N_25118,N_24514);
or U29830 (N_29830,N_26276,N_26746);
nand U29831 (N_29831,N_25786,N_25563);
or U29832 (N_29832,N_25505,N_26609);
or U29833 (N_29833,N_26376,N_25933);
or U29834 (N_29834,N_24187,N_26436);
xnor U29835 (N_29835,N_24659,N_26517);
xor U29836 (N_29836,N_25391,N_25864);
nand U29837 (N_29837,N_26186,N_25545);
nor U29838 (N_29838,N_26674,N_25629);
nor U29839 (N_29839,N_24104,N_26449);
xnor U29840 (N_29840,N_26786,N_26067);
nand U29841 (N_29841,N_25897,N_25719);
or U29842 (N_29842,N_26315,N_24307);
and U29843 (N_29843,N_26271,N_24777);
xnor U29844 (N_29844,N_26555,N_26174);
or U29845 (N_29845,N_25548,N_25602);
xnor U29846 (N_29846,N_26170,N_25830);
nor U29847 (N_29847,N_24835,N_25336);
xor U29848 (N_29848,N_24129,N_25349);
xor U29849 (N_29849,N_25699,N_26051);
nor U29850 (N_29850,N_25032,N_24577);
xnor U29851 (N_29851,N_25017,N_25574);
or U29852 (N_29852,N_26130,N_24149);
xnor U29853 (N_29853,N_24343,N_24193);
nand U29854 (N_29854,N_25153,N_24635);
xor U29855 (N_29855,N_26430,N_25746);
and U29856 (N_29856,N_25790,N_24331);
nor U29857 (N_29857,N_24186,N_24552);
xor U29858 (N_29858,N_24871,N_25790);
and U29859 (N_29859,N_25260,N_26523);
or U29860 (N_29860,N_26314,N_26401);
nor U29861 (N_29861,N_26676,N_25303);
or U29862 (N_29862,N_25796,N_25226);
or U29863 (N_29863,N_25728,N_24590);
and U29864 (N_29864,N_26862,N_25373);
and U29865 (N_29865,N_24022,N_25925);
nor U29866 (N_29866,N_26820,N_26438);
or U29867 (N_29867,N_26747,N_25757);
or U29868 (N_29868,N_25039,N_24731);
xnor U29869 (N_29869,N_26161,N_26575);
nand U29870 (N_29870,N_24677,N_25254);
and U29871 (N_29871,N_25897,N_25566);
xor U29872 (N_29872,N_24638,N_25200);
xor U29873 (N_29873,N_26375,N_24636);
xnor U29874 (N_29874,N_26635,N_25585);
nor U29875 (N_29875,N_25304,N_25632);
and U29876 (N_29876,N_24299,N_26557);
nor U29877 (N_29877,N_26884,N_26198);
and U29878 (N_29878,N_25747,N_24642);
nand U29879 (N_29879,N_25417,N_24958);
nor U29880 (N_29880,N_26777,N_25384);
nor U29881 (N_29881,N_25633,N_26370);
or U29882 (N_29882,N_24505,N_24150);
xor U29883 (N_29883,N_26286,N_25481);
nor U29884 (N_29884,N_24671,N_26209);
or U29885 (N_29885,N_26476,N_26537);
xnor U29886 (N_29886,N_26435,N_24488);
nand U29887 (N_29887,N_24498,N_26932);
and U29888 (N_29888,N_25362,N_26126);
or U29889 (N_29889,N_26535,N_24290);
nor U29890 (N_29890,N_25269,N_26372);
nor U29891 (N_29891,N_25438,N_25034);
or U29892 (N_29892,N_24730,N_24976);
nor U29893 (N_29893,N_25775,N_24541);
xnor U29894 (N_29894,N_24918,N_26629);
or U29895 (N_29895,N_25410,N_25250);
xnor U29896 (N_29896,N_24320,N_24843);
nor U29897 (N_29897,N_25870,N_24390);
nor U29898 (N_29898,N_26977,N_26754);
and U29899 (N_29899,N_24682,N_24236);
or U29900 (N_29900,N_25357,N_24250);
or U29901 (N_29901,N_25809,N_26734);
nand U29902 (N_29902,N_24773,N_24825);
nor U29903 (N_29903,N_24349,N_24153);
or U29904 (N_29904,N_24594,N_24771);
and U29905 (N_29905,N_25504,N_24850);
or U29906 (N_29906,N_26775,N_25710);
nor U29907 (N_29907,N_24607,N_25376);
or U29908 (N_29908,N_25863,N_25892);
nor U29909 (N_29909,N_26037,N_24252);
nand U29910 (N_29910,N_26050,N_26854);
xor U29911 (N_29911,N_24978,N_26682);
nor U29912 (N_29912,N_25862,N_24304);
or U29913 (N_29913,N_24323,N_25223);
xor U29914 (N_29914,N_24543,N_26759);
nand U29915 (N_29915,N_25053,N_25002);
and U29916 (N_29916,N_24598,N_25707);
or U29917 (N_29917,N_24336,N_24723);
and U29918 (N_29918,N_25750,N_25593);
xnor U29919 (N_29919,N_24036,N_25691);
or U29920 (N_29920,N_26148,N_25271);
and U29921 (N_29921,N_25121,N_24752);
nor U29922 (N_29922,N_26022,N_24910);
xor U29923 (N_29923,N_24304,N_24778);
and U29924 (N_29924,N_25012,N_24954);
nand U29925 (N_29925,N_25437,N_24332);
xor U29926 (N_29926,N_25858,N_26055);
nor U29927 (N_29927,N_25814,N_25089);
or U29928 (N_29928,N_25102,N_24317);
or U29929 (N_29929,N_24049,N_26028);
nand U29930 (N_29930,N_26062,N_25811);
xor U29931 (N_29931,N_26372,N_24025);
and U29932 (N_29932,N_25692,N_25110);
and U29933 (N_29933,N_26366,N_24272);
xor U29934 (N_29934,N_26112,N_24504);
nand U29935 (N_29935,N_25973,N_24587);
xor U29936 (N_29936,N_24501,N_25845);
xor U29937 (N_29937,N_26964,N_24499);
nand U29938 (N_29938,N_26255,N_25797);
nand U29939 (N_29939,N_25641,N_24652);
xnor U29940 (N_29940,N_24313,N_24301);
nor U29941 (N_29941,N_25742,N_26857);
nor U29942 (N_29942,N_25719,N_24758);
xor U29943 (N_29943,N_25887,N_24200);
or U29944 (N_29944,N_26233,N_26268);
and U29945 (N_29945,N_26620,N_26871);
nor U29946 (N_29946,N_25877,N_24044);
and U29947 (N_29947,N_24099,N_24891);
or U29948 (N_29948,N_26053,N_24323);
or U29949 (N_29949,N_26834,N_25123);
nor U29950 (N_29950,N_25445,N_26322);
xnor U29951 (N_29951,N_25008,N_24068);
or U29952 (N_29952,N_24959,N_24400);
or U29953 (N_29953,N_24661,N_25778);
xnor U29954 (N_29954,N_24575,N_24332);
xor U29955 (N_29955,N_24390,N_25152);
or U29956 (N_29956,N_26097,N_26224);
nand U29957 (N_29957,N_25901,N_24357);
or U29958 (N_29958,N_24432,N_24780);
nor U29959 (N_29959,N_26453,N_25846);
or U29960 (N_29960,N_24539,N_24743);
or U29961 (N_29961,N_24320,N_25379);
or U29962 (N_29962,N_26668,N_24827);
and U29963 (N_29963,N_24891,N_24724);
and U29964 (N_29964,N_25689,N_25839);
xor U29965 (N_29965,N_24708,N_25155);
xnor U29966 (N_29966,N_25618,N_26012);
or U29967 (N_29967,N_25961,N_25535);
or U29968 (N_29968,N_24445,N_24682);
or U29969 (N_29969,N_26352,N_25724);
nor U29970 (N_29970,N_26864,N_25385);
xnor U29971 (N_29971,N_26055,N_24723);
xnor U29972 (N_29972,N_25658,N_25970);
nand U29973 (N_29973,N_26422,N_24252);
nor U29974 (N_29974,N_25189,N_26275);
nand U29975 (N_29975,N_26429,N_26361);
and U29976 (N_29976,N_24264,N_24644);
or U29977 (N_29977,N_26406,N_24507);
xor U29978 (N_29978,N_24247,N_24386);
nand U29979 (N_29979,N_26412,N_26071);
nand U29980 (N_29980,N_25122,N_25982);
or U29981 (N_29981,N_24120,N_26225);
xor U29982 (N_29982,N_25130,N_24392);
and U29983 (N_29983,N_25303,N_24065);
xnor U29984 (N_29984,N_25236,N_25699);
nor U29985 (N_29985,N_25942,N_26447);
or U29986 (N_29986,N_25343,N_26299);
nor U29987 (N_29987,N_25795,N_24682);
nor U29988 (N_29988,N_25385,N_26367);
and U29989 (N_29989,N_26274,N_26578);
nor U29990 (N_29990,N_25405,N_25044);
xor U29991 (N_29991,N_24474,N_26841);
nor U29992 (N_29992,N_25692,N_26582);
and U29993 (N_29993,N_25752,N_26404);
or U29994 (N_29994,N_26330,N_25497);
and U29995 (N_29995,N_25332,N_24288);
nor U29996 (N_29996,N_26331,N_25427);
nor U29997 (N_29997,N_24240,N_25944);
or U29998 (N_29998,N_24935,N_25401);
xor U29999 (N_29999,N_24568,N_24610);
xnor UO_0 (O_0,N_29955,N_29271);
nand UO_1 (O_1,N_29056,N_27261);
or UO_2 (O_2,N_28996,N_27389);
and UO_3 (O_3,N_28631,N_28223);
nand UO_4 (O_4,N_29917,N_29313);
xor UO_5 (O_5,N_28615,N_28436);
and UO_6 (O_6,N_28699,N_29558);
and UO_7 (O_7,N_29352,N_28005);
or UO_8 (O_8,N_29262,N_27100);
or UO_9 (O_9,N_27891,N_28767);
or UO_10 (O_10,N_28067,N_28637);
and UO_11 (O_11,N_29025,N_29930);
and UO_12 (O_12,N_28925,N_28167);
xor UO_13 (O_13,N_27072,N_28449);
nand UO_14 (O_14,N_28183,N_29153);
nand UO_15 (O_15,N_29308,N_28232);
nor UO_16 (O_16,N_28219,N_29230);
and UO_17 (O_17,N_29004,N_29291);
xor UO_18 (O_18,N_29422,N_28203);
or UO_19 (O_19,N_27413,N_29003);
nor UO_20 (O_20,N_28195,N_27673);
and UO_21 (O_21,N_29761,N_29042);
and UO_22 (O_22,N_29831,N_27635);
xnor UO_23 (O_23,N_27031,N_28603);
or UO_24 (O_24,N_29502,N_27664);
nand UO_25 (O_25,N_29724,N_29898);
nand UO_26 (O_26,N_29924,N_27535);
xnor UO_27 (O_27,N_29106,N_28485);
xnor UO_28 (O_28,N_28052,N_27213);
or UO_29 (O_29,N_28759,N_27161);
nor UO_30 (O_30,N_27479,N_28434);
xnor UO_31 (O_31,N_27536,N_28374);
nand UO_32 (O_32,N_29981,N_29903);
or UO_33 (O_33,N_29904,N_28487);
nand UO_34 (O_34,N_27960,N_29604);
nor UO_35 (O_35,N_27944,N_28537);
nand UO_36 (O_36,N_29733,N_28983);
nand UO_37 (O_37,N_27822,N_27600);
xor UO_38 (O_38,N_28505,N_29293);
and UO_39 (O_39,N_27777,N_29988);
and UO_40 (O_40,N_27178,N_29492);
and UO_41 (O_41,N_27328,N_29404);
and UO_42 (O_42,N_28033,N_27611);
or UO_43 (O_43,N_29397,N_29549);
nand UO_44 (O_44,N_28519,N_27314);
nor UO_45 (O_45,N_27561,N_28225);
xnor UO_46 (O_46,N_28278,N_27268);
or UO_47 (O_47,N_29169,N_27110);
xor UO_48 (O_48,N_29157,N_27106);
nor UO_49 (O_49,N_29662,N_28504);
and UO_50 (O_50,N_29695,N_29031);
nor UO_51 (O_51,N_27377,N_29769);
xnor UO_52 (O_52,N_29253,N_27878);
and UO_53 (O_53,N_29447,N_28113);
xnor UO_54 (O_54,N_29163,N_28105);
nor UO_55 (O_55,N_28212,N_27453);
nor UO_56 (O_56,N_28660,N_28517);
xnor UO_57 (O_57,N_27608,N_27010);
xor UO_58 (O_58,N_29252,N_29837);
nand UO_59 (O_59,N_29997,N_29569);
nand UO_60 (O_60,N_28139,N_28150);
nor UO_61 (O_61,N_27175,N_29865);
nand UO_62 (O_62,N_27484,N_27671);
nor UO_63 (O_63,N_28679,N_29869);
nor UO_64 (O_64,N_28456,N_29848);
nor UO_65 (O_65,N_29358,N_28815);
xor UO_66 (O_66,N_28286,N_29192);
nand UO_67 (O_67,N_28502,N_27696);
and UO_68 (O_68,N_27816,N_28410);
or UO_69 (O_69,N_27419,N_28110);
and UO_70 (O_70,N_27787,N_28227);
xnor UO_71 (O_71,N_29793,N_27636);
nor UO_72 (O_72,N_29998,N_28606);
or UO_73 (O_73,N_27245,N_28403);
nand UO_74 (O_74,N_27667,N_27494);
and UO_75 (O_75,N_29684,N_29914);
xor UO_76 (O_76,N_29611,N_29841);
and UO_77 (O_77,N_27588,N_29249);
nor UO_78 (O_78,N_27622,N_29757);
and UO_79 (O_79,N_28642,N_27058);
nor UO_80 (O_80,N_28211,N_28848);
nor UO_81 (O_81,N_29780,N_28459);
xor UO_82 (O_82,N_29199,N_28307);
xor UO_83 (O_83,N_27024,N_27590);
nand UO_84 (O_84,N_28712,N_28906);
and UO_85 (O_85,N_29941,N_28088);
or UO_86 (O_86,N_29952,N_27862);
xor UO_87 (O_87,N_29797,N_29136);
and UO_88 (O_88,N_27784,N_29779);
xor UO_89 (O_89,N_28064,N_27294);
nor UO_90 (O_90,N_28316,N_27235);
xor UO_91 (O_91,N_27525,N_27919);
or UO_92 (O_92,N_29918,N_27420);
nor UO_93 (O_93,N_28412,N_29643);
nor UO_94 (O_94,N_29024,N_29411);
and UO_95 (O_95,N_29150,N_28473);
or UO_96 (O_96,N_28454,N_28457);
xnor UO_97 (O_97,N_27633,N_27527);
and UO_98 (O_98,N_27128,N_28509);
xnor UO_99 (O_99,N_28363,N_28920);
nand UO_100 (O_100,N_28216,N_27382);
or UO_101 (O_101,N_29123,N_28243);
nor UO_102 (O_102,N_27360,N_27693);
xor UO_103 (O_103,N_28790,N_28241);
nor UO_104 (O_104,N_29139,N_27158);
xor UO_105 (O_105,N_28035,N_28400);
xnor UO_106 (O_106,N_28069,N_27032);
or UO_107 (O_107,N_27613,N_27039);
xor UO_108 (O_108,N_28799,N_29138);
nand UO_109 (O_109,N_29834,N_28168);
xnor UO_110 (O_110,N_27904,N_29812);
or UO_111 (O_111,N_28065,N_28002);
xor UO_112 (O_112,N_27978,N_29204);
or UO_113 (O_113,N_28582,N_27576);
xor UO_114 (O_114,N_27977,N_28467);
and UO_115 (O_115,N_28599,N_28813);
nor UO_116 (O_116,N_29129,N_29525);
xor UO_117 (O_117,N_27095,N_28725);
nor UO_118 (O_118,N_29175,N_29939);
and UO_119 (O_119,N_28226,N_27103);
nand UO_120 (O_120,N_28377,N_27899);
nand UO_121 (O_121,N_28433,N_27012);
and UO_122 (O_122,N_27201,N_28944);
nand UO_123 (O_123,N_27283,N_29882);
and UO_124 (O_124,N_28010,N_28146);
xor UO_125 (O_125,N_29122,N_27749);
nand UO_126 (O_126,N_27312,N_27874);
nor UO_127 (O_127,N_27866,N_29061);
or UO_128 (O_128,N_28273,N_27873);
xnor UO_129 (O_129,N_29664,N_27928);
and UO_130 (O_130,N_28826,N_29995);
xnor UO_131 (O_131,N_29279,N_29171);
nor UO_132 (O_132,N_29266,N_27317);
and UO_133 (O_133,N_28758,N_27371);
xor UO_134 (O_134,N_29176,N_27473);
xnor UO_135 (O_135,N_29702,N_27192);
and UO_136 (O_136,N_28391,N_27188);
and UO_137 (O_137,N_28722,N_29333);
nor UO_138 (O_138,N_28570,N_29720);
and UO_139 (O_139,N_29661,N_29760);
and UO_140 (O_140,N_27686,N_28738);
nor UO_141 (O_141,N_28998,N_29573);
nor UO_142 (O_142,N_27991,N_27480);
and UO_143 (O_143,N_27586,N_28928);
or UO_144 (O_144,N_29181,N_29329);
nand UO_145 (O_145,N_28420,N_28240);
nor UO_146 (O_146,N_29351,N_28149);
and UO_147 (O_147,N_27859,N_27096);
and UO_148 (O_148,N_29993,N_29620);
and UO_149 (O_149,N_28109,N_29172);
or UO_150 (O_150,N_29883,N_28828);
and UO_151 (O_151,N_29096,N_28927);
nor UO_152 (O_152,N_29739,N_27470);
xnor UO_153 (O_153,N_27153,N_28032);
or UO_154 (O_154,N_27451,N_27515);
nor UO_155 (O_155,N_27378,N_28288);
or UO_156 (O_156,N_29730,N_28342);
nor UO_157 (O_157,N_29033,N_28174);
nor UO_158 (O_158,N_28484,N_28869);
or UO_159 (O_159,N_28413,N_28562);
nor UO_160 (O_160,N_27387,N_29946);
nor UO_161 (O_161,N_28770,N_27794);
or UO_162 (O_162,N_27144,N_27523);
xnor UO_163 (O_163,N_27560,N_29101);
and UO_164 (O_164,N_27246,N_28074);
or UO_165 (O_165,N_28737,N_29005);
nand UO_166 (O_166,N_28127,N_29305);
xnor UO_167 (O_167,N_27281,N_28675);
and UO_168 (O_168,N_28215,N_29294);
nand UO_169 (O_169,N_27951,N_27884);
nand UO_170 (O_170,N_27895,N_28780);
nor UO_171 (O_171,N_27680,N_28971);
or UO_172 (O_172,N_29234,N_27547);
and UO_173 (O_173,N_27155,N_27579);
xnor UO_174 (O_174,N_27423,N_27203);
nor UO_175 (O_175,N_28846,N_28244);
nand UO_176 (O_176,N_29211,N_28483);
and UO_177 (O_177,N_28355,N_29973);
or UO_178 (O_178,N_29556,N_27701);
xor UO_179 (O_179,N_27087,N_27882);
nor UO_180 (O_180,N_27141,N_27214);
and UO_181 (O_181,N_27455,N_27077);
or UO_182 (O_182,N_28945,N_29484);
and UO_183 (O_183,N_29531,N_28480);
or UO_184 (O_184,N_28914,N_27861);
nand UO_185 (O_185,N_27939,N_28026);
or UO_186 (O_186,N_29615,N_29270);
nand UO_187 (O_187,N_27388,N_27887);
or UO_188 (O_188,N_29445,N_27638);
nor UO_189 (O_189,N_28023,N_28047);
or UO_190 (O_190,N_28321,N_28408);
or UO_191 (O_191,N_29663,N_29921);
or UO_192 (O_192,N_29544,N_28789);
or UO_193 (O_193,N_27856,N_28867);
xnor UO_194 (O_194,N_27783,N_28531);
or UO_195 (O_195,N_27107,N_29207);
nor UO_196 (O_196,N_28339,N_28809);
xnor UO_197 (O_197,N_28380,N_27810);
and UO_198 (O_198,N_28124,N_27612);
nand UO_199 (O_199,N_28702,N_29110);
and UO_200 (O_200,N_28112,N_28888);
or UO_201 (O_201,N_27775,N_27168);
and UO_202 (O_202,N_27081,N_29514);
and UO_203 (O_203,N_27826,N_28585);
or UO_204 (O_204,N_29160,N_28879);
and UO_205 (O_205,N_29020,N_27559);
nand UO_206 (O_206,N_28808,N_27132);
nand UO_207 (O_207,N_27599,N_28267);
nor UO_208 (O_208,N_27662,N_29501);
nor UO_209 (O_209,N_27068,N_28624);
nor UO_210 (O_210,N_28042,N_28806);
nand UO_211 (O_211,N_28651,N_28486);
and UO_212 (O_212,N_28025,N_27057);
nand UO_213 (O_213,N_29519,N_28892);
and UO_214 (O_214,N_27832,N_27018);
or UO_215 (O_215,N_27989,N_29623);
or UO_216 (O_216,N_29855,N_29185);
nand UO_217 (O_217,N_29506,N_28668);
nand UO_218 (O_218,N_27804,N_29594);
nand UO_219 (O_219,N_29335,N_28249);
xor UO_220 (O_220,N_28787,N_27257);
nor UO_221 (O_221,N_28401,N_29390);
or UO_222 (O_222,N_28089,N_29711);
nor UO_223 (O_223,N_28349,N_29037);
or UO_224 (O_224,N_27914,N_27477);
nand UO_225 (O_225,N_27459,N_28008);
and UO_226 (O_226,N_29121,N_28994);
nor UO_227 (O_227,N_28807,N_29016);
nand UO_228 (O_228,N_27184,N_27946);
and UO_229 (O_229,N_29665,N_29434);
and UO_230 (O_230,N_29375,N_29449);
nand UO_231 (O_231,N_27011,N_29919);
xor UO_232 (O_232,N_27123,N_29732);
nor UO_233 (O_233,N_29217,N_29376);
or UO_234 (O_234,N_29959,N_28359);
xor UO_235 (O_235,N_28620,N_29692);
and UO_236 (O_236,N_27618,N_29710);
xor UO_237 (O_237,N_27949,N_27952);
xor UO_238 (O_238,N_28987,N_27071);
and UO_239 (O_239,N_28070,N_28716);
and UO_240 (O_240,N_27481,N_29605);
and UO_241 (O_241,N_27570,N_27157);
or UO_242 (O_242,N_27631,N_28075);
nand UO_243 (O_243,N_28426,N_29480);
nand UO_244 (O_244,N_28810,N_28082);
nand UO_245 (O_245,N_28394,N_27052);
nor UO_246 (O_246,N_29010,N_27177);
nand UO_247 (O_247,N_28742,N_27567);
nor UO_248 (O_248,N_29022,N_28794);
and UO_249 (O_249,N_28686,N_27198);
xnor UO_250 (O_250,N_28491,N_28283);
and UO_251 (O_251,N_28255,N_28850);
or UO_252 (O_252,N_27835,N_27705);
and UO_253 (O_253,N_29499,N_27778);
xor UO_254 (O_254,N_27362,N_29627);
nor UO_255 (O_255,N_29740,N_29628);
and UO_256 (O_256,N_28136,N_27913);
or UO_257 (O_257,N_28908,N_29088);
or UO_258 (O_258,N_28282,N_29255);
xor UO_259 (O_259,N_27838,N_28918);
and UO_260 (O_260,N_29269,N_27185);
and UO_261 (O_261,N_28445,N_27359);
and UO_262 (O_262,N_28719,N_27137);
nand UO_263 (O_263,N_28823,N_28543);
xor UO_264 (O_264,N_27485,N_29507);
nand UO_265 (O_265,N_29448,N_27996);
nand UO_266 (O_266,N_29331,N_28859);
xor UO_267 (O_267,N_29045,N_28550);
xnor UO_268 (O_268,N_29453,N_29147);
nand UO_269 (O_269,N_27027,N_28793);
nor UO_270 (O_270,N_29585,N_28833);
or UO_271 (O_271,N_27392,N_28322);
nand UO_272 (O_272,N_28508,N_29555);
or UO_273 (O_273,N_29144,N_27722);
xor UO_274 (O_274,N_28302,N_27806);
or UO_275 (O_275,N_29301,N_28559);
or UO_276 (O_276,N_29667,N_28577);
xor UO_277 (O_277,N_28123,N_28043);
or UO_278 (O_278,N_28118,N_28430);
and UO_279 (O_279,N_27326,N_27520);
xor UO_280 (O_280,N_27207,N_29971);
and UO_281 (O_281,N_28720,N_27179);
xor UO_282 (O_282,N_27465,N_29897);
xor UO_283 (O_283,N_29547,N_29191);
or UO_284 (O_284,N_29465,N_29057);
nor UO_285 (O_285,N_29328,N_28335);
xnor UO_286 (O_286,N_27801,N_28027);
nand UO_287 (O_287,N_27251,N_28341);
nor UO_288 (O_288,N_27467,N_29155);
or UO_289 (O_289,N_27578,N_29963);
xor UO_290 (O_290,N_29112,N_29906);
nor UO_291 (O_291,N_29395,N_28234);
nand UO_292 (O_292,N_28134,N_27898);
or UO_293 (O_293,N_27981,N_27379);
and UO_294 (O_294,N_28894,N_29134);
nand UO_295 (O_295,N_28334,N_27511);
nand UO_296 (O_296,N_27365,N_27677);
or UO_297 (O_297,N_29215,N_27720);
and UO_298 (O_298,N_29391,N_27444);
nor UO_299 (O_299,N_27774,N_27212);
nor UO_300 (O_300,N_27566,N_27751);
and UO_301 (O_301,N_29942,N_27974);
nand UO_302 (O_302,N_29912,N_28788);
xnor UO_303 (O_303,N_28930,N_28298);
nand UO_304 (O_304,N_27117,N_27236);
xor UO_305 (O_305,N_28545,N_29379);
nor UO_306 (O_306,N_29315,N_28511);
nand UO_307 (O_307,N_29454,N_27607);
or UO_308 (O_308,N_28164,N_28315);
nand UO_309 (O_309,N_28761,N_29802);
nand UO_310 (O_310,N_28049,N_29392);
or UO_311 (O_311,N_29572,N_29950);
and UO_312 (O_312,N_29637,N_29413);
nand UO_313 (O_313,N_27145,N_29074);
and UO_314 (O_314,N_27475,N_29978);
nand UO_315 (O_315,N_27313,N_27393);
and UO_316 (O_316,N_28617,N_29595);
nor UO_317 (O_317,N_28407,N_29443);
xnor UO_318 (O_318,N_27616,N_28801);
xnor UO_319 (O_319,N_28352,N_27329);
and UO_320 (O_320,N_27112,N_28804);
and UO_321 (O_321,N_27228,N_29178);
or UO_322 (O_322,N_27311,N_28985);
nor UO_323 (O_323,N_29670,N_29124);
nand UO_324 (O_324,N_27512,N_28956);
nor UO_325 (O_325,N_29895,N_29164);
nor UO_326 (O_326,N_28547,N_27008);
xnor UO_327 (O_327,N_29938,N_29093);
nand UO_328 (O_328,N_29884,N_28776);
and UO_329 (O_329,N_27718,N_27152);
nand UO_330 (O_330,N_29070,N_28347);
xnor UO_331 (O_331,N_29052,N_27262);
nor UO_332 (O_332,N_29188,N_29618);
xor UO_333 (O_333,N_27640,N_28728);
xnor UO_334 (O_334,N_28865,N_29489);
xnor UO_335 (O_335,N_27334,N_28265);
xnor UO_336 (O_336,N_29205,N_29463);
and UO_337 (O_337,N_27487,N_28197);
or UO_338 (O_338,N_27966,N_27972);
xnor UO_339 (O_339,N_29055,N_28544);
or UO_340 (O_340,N_29084,N_28614);
xor UO_341 (O_341,N_29767,N_28692);
or UO_342 (O_342,N_27015,N_29421);
and UO_343 (O_343,N_27042,N_27865);
xor UO_344 (O_344,N_28522,N_29994);
and UO_345 (O_345,N_29246,N_29048);
or UO_346 (O_346,N_29140,N_28836);
nor UO_347 (O_347,N_27468,N_29356);
xor UO_348 (O_348,N_27504,N_29584);
nand UO_349 (O_349,N_27217,N_29888);
xor UO_350 (O_350,N_27344,N_29681);
or UO_351 (O_351,N_28510,N_28791);
nor UO_352 (O_352,N_29726,N_27463);
or UO_353 (O_353,N_28604,N_27164);
or UO_354 (O_354,N_29259,N_27256);
nand UO_355 (O_355,N_29113,N_27428);
xor UO_356 (O_356,N_29565,N_27736);
and UO_357 (O_357,N_27795,N_27061);
and UO_358 (O_358,N_28648,N_27374);
xor UO_359 (O_359,N_27290,N_29872);
nor UO_360 (O_360,N_29817,N_28180);
nor UO_361 (O_361,N_27211,N_27224);
nand UO_362 (O_362,N_28022,N_27458);
and UO_363 (O_363,N_29648,N_29986);
or UO_364 (O_364,N_29274,N_28329);
and UO_365 (O_365,N_28703,N_28520);
or UO_366 (O_366,N_28091,N_29861);
and UO_367 (O_367,N_28609,N_28220);
xor UO_368 (O_368,N_29516,N_28166);
and UO_369 (O_369,N_27337,N_29455);
or UO_370 (O_370,N_28007,N_29715);
nand UO_371 (O_371,N_28000,N_29947);
or UO_372 (O_372,N_29829,N_29469);
xnor UO_373 (O_373,N_27843,N_28084);
and UO_374 (O_374,N_29653,N_27133);
and UO_375 (O_375,N_29660,N_27513);
xor UO_376 (O_376,N_29989,N_28441);
nand UO_377 (O_377,N_27037,N_28418);
nand UO_378 (O_378,N_29340,N_28698);
and UO_379 (O_379,N_28272,N_27051);
or UO_380 (O_380,N_29583,N_29082);
nand UO_381 (O_381,N_28652,N_29878);
xor UO_382 (O_382,N_27354,N_27752);
and UO_383 (O_383,N_28125,N_27764);
and UO_384 (O_384,N_28100,N_28452);
or UO_385 (O_385,N_28235,N_27358);
xor UO_386 (O_386,N_29467,N_29568);
or UO_387 (O_387,N_27048,N_29626);
nor UO_388 (O_388,N_28602,N_28764);
nand UO_389 (O_389,N_27927,N_28530);
nor UO_390 (O_390,N_29401,N_28156);
nand UO_391 (O_391,N_28160,N_29880);
or UO_392 (O_392,N_28524,N_27282);
nor UO_393 (O_393,N_28422,N_29578);
xnor UO_394 (O_394,N_28934,N_28571);
nand UO_395 (O_395,N_29579,N_28576);
nand UO_396 (O_396,N_27768,N_28636);
xor UO_397 (O_397,N_28816,N_29886);
nor UO_398 (O_398,N_27398,N_27406);
nor UO_399 (O_399,N_28919,N_29874);
and UO_400 (O_400,N_29423,N_27624);
nand UO_401 (O_401,N_27316,N_28428);
xor UO_402 (O_402,N_29592,N_29366);
or UO_403 (O_403,N_28729,N_29580);
nor UO_404 (O_404,N_27293,N_27482);
xnor UO_405 (O_405,N_29384,N_29983);
xnor UO_406 (O_406,N_27648,N_27028);
nor UO_407 (O_407,N_29546,N_27279);
or UO_408 (O_408,N_29617,N_27528);
xnor UO_409 (O_409,N_29195,N_27324);
nor UO_410 (O_410,N_28475,N_29777);
xnor UO_411 (O_411,N_27020,N_29382);
or UO_412 (O_412,N_27756,N_28356);
and UO_413 (O_413,N_29148,N_27265);
nand UO_414 (O_414,N_27429,N_27524);
or UO_415 (O_415,N_29790,N_27017);
nor UO_416 (O_416,N_28402,N_28293);
xnor UO_417 (O_417,N_29430,N_29035);
or UO_418 (O_418,N_28901,N_27791);
xor UO_419 (O_419,N_29735,N_27872);
nor UO_420 (O_420,N_27833,N_29203);
xor UO_421 (O_421,N_27734,N_27260);
xor UO_422 (O_422,N_29638,N_27564);
nand UO_423 (O_423,N_28965,N_27780);
nand UO_424 (O_424,N_27690,N_27993);
or UO_425 (O_425,N_28192,N_28959);
and UO_426 (O_426,N_28176,N_27171);
or UO_427 (O_427,N_27227,N_27990);
or UO_428 (O_428,N_27304,N_27506);
nor UO_429 (O_429,N_27248,N_27765);
nand UO_430 (O_430,N_29137,N_27836);
xnor UO_431 (O_431,N_29808,N_27291);
nor UO_432 (O_432,N_29945,N_29844);
nand UO_433 (O_433,N_28479,N_27584);
or UO_434 (O_434,N_28396,N_28515);
nand UO_435 (O_435,N_29241,N_29932);
or UO_436 (O_436,N_27376,N_27094);
nor UO_437 (O_437,N_28546,N_28344);
or UO_438 (O_438,N_27197,N_29539);
xnor UO_439 (O_439,N_29302,N_27741);
nor UO_440 (O_440,N_28845,N_29370);
xor UO_441 (O_441,N_27811,N_29717);
nor UO_442 (O_442,N_28498,N_28924);
nand UO_443 (O_443,N_28465,N_27418);
and UO_444 (O_444,N_29508,N_27967);
or UO_445 (O_445,N_27649,N_28549);
nand UO_446 (O_446,N_27000,N_29407);
xor UO_447 (O_447,N_27926,N_28558);
and UO_448 (O_448,N_27670,N_29826);
xnor UO_449 (O_449,N_27743,N_29159);
nor UO_450 (O_450,N_27434,N_29001);
xnor UO_451 (O_451,N_29077,N_28437);
nor UO_452 (O_452,N_29689,N_27647);
nand UO_453 (O_453,N_29091,N_29372);
nor UO_454 (O_454,N_28337,N_27395);
or UO_455 (O_455,N_28497,N_28063);
and UO_456 (O_456,N_27685,N_28157);
nand UO_457 (O_457,N_28458,N_29131);
nor UO_458 (O_458,N_29051,N_28425);
xnor UO_459 (O_459,N_29126,N_29535);
nand UO_460 (O_460,N_27270,N_28263);
nand UO_461 (O_461,N_29151,N_29498);
nand UO_462 (O_462,N_29712,N_27642);
xor UO_463 (O_463,N_29833,N_29840);
or UO_464 (O_464,N_28464,N_27263);
xnor UO_465 (O_465,N_28542,N_29424);
or UO_466 (O_466,N_27180,N_27476);
nand UO_467 (O_467,N_28299,N_28727);
nand UO_468 (O_468,N_27274,N_29783);
and UO_469 (O_469,N_27383,N_28557);
or UO_470 (O_470,N_28138,N_29312);
nand UO_471 (O_471,N_27735,N_29278);
xor UO_472 (O_472,N_28656,N_27066);
nand UO_473 (O_473,N_27125,N_29450);
and UO_474 (O_474,N_29723,N_28536);
and UO_475 (O_475,N_29251,N_29075);
and UO_476 (O_476,N_29054,N_28739);
nand UO_477 (O_477,N_29889,N_28085);
xor UO_478 (O_478,N_29478,N_27970);
xnor UO_479 (O_479,N_28704,N_27727);
xnor UO_480 (O_480,N_27830,N_29161);
nand UO_481 (O_481,N_28916,N_29901);
or UO_482 (O_482,N_28644,N_28367);
xor UO_483 (O_483,N_27505,N_27014);
xor UO_484 (O_484,N_27658,N_29190);
and UO_485 (O_485,N_29283,N_27805);
and UO_486 (O_486,N_28817,N_27712);
xnor UO_487 (O_487,N_29257,N_28943);
and UO_488 (O_488,N_29713,N_27210);
nand UO_489 (O_489,N_27786,N_28782);
nor UO_490 (O_490,N_28990,N_29613);
nand UO_491 (O_491,N_29418,N_29642);
and UO_492 (O_492,N_29629,N_27592);
xor UO_493 (O_493,N_27206,N_28169);
nand UO_494 (O_494,N_28805,N_28490);
and UO_495 (O_495,N_27421,N_28744);
and UO_496 (O_496,N_29859,N_27143);
nand UO_497 (O_497,N_28619,N_27645);
or UO_498 (O_498,N_29676,N_29023);
and UO_499 (O_499,N_28097,N_28364);
nor UO_500 (O_500,N_29267,N_28685);
nor UO_501 (O_501,N_27307,N_27483);
nor UO_502 (O_502,N_27955,N_29916);
or UO_503 (O_503,N_28590,N_29388);
xnor UO_504 (O_504,N_28763,N_27726);
nand UO_505 (O_505,N_29344,N_28607);
nor UO_506 (O_506,N_27089,N_29095);
nand UO_507 (O_507,N_27797,N_29591);
xor UO_508 (O_508,N_29510,N_28680);
and UO_509 (O_509,N_29482,N_29245);
nand UO_510 (O_510,N_29589,N_27150);
xor UO_511 (O_511,N_28297,N_29563);
nor UO_512 (O_512,N_28783,N_28379);
xnor UO_513 (O_513,N_29201,N_29458);
and UO_514 (O_514,N_29087,N_27043);
and UO_515 (O_515,N_29426,N_28989);
nand UO_516 (O_516,N_28256,N_28527);
or UO_517 (O_517,N_29038,N_28252);
and UO_518 (O_518,N_29784,N_27375);
xnor UO_519 (O_519,N_27992,N_28133);
and UO_520 (O_520,N_27204,N_29438);
nor UO_521 (O_521,N_27055,N_28866);
nor UO_522 (O_522,N_29899,N_29871);
or UO_523 (O_523,N_27557,N_29527);
and UO_524 (O_524,N_29644,N_28264);
or UO_525 (O_525,N_28046,N_28909);
nor UO_526 (O_526,N_27848,N_29678);
or UO_527 (O_527,N_28820,N_28891);
or UO_528 (O_528,N_29470,N_27845);
or UO_529 (O_529,N_27875,N_27102);
and UO_530 (O_530,N_28872,N_29513);
or UO_531 (O_531,N_27396,N_27773);
and UO_532 (O_532,N_27994,N_28248);
nand UO_533 (O_533,N_27907,N_27500);
xor UO_534 (O_534,N_29835,N_28311);
and UO_535 (O_535,N_27169,N_29260);
xor UO_536 (O_536,N_29847,N_28336);
or UO_537 (O_537,N_27782,N_28414);
nor UO_538 (O_538,N_29647,N_27044);
xor UO_539 (O_539,N_27819,N_27076);
and UO_540 (O_540,N_27433,N_29951);
nand UO_541 (O_541,N_27562,N_27985);
nor UO_542 (O_542,N_28201,N_28466);
nand UO_543 (O_543,N_27183,N_29338);
nand UO_544 (O_544,N_27182,N_27047);
nor UO_545 (O_545,N_27229,N_28640);
or UO_546 (O_546,N_28371,N_29365);
nor UO_547 (O_547,N_28245,N_27437);
nand UO_548 (O_548,N_28958,N_28472);
xnor UO_549 (O_549,N_28194,N_27738);
or UO_550 (O_550,N_29851,N_27219);
nor UO_551 (O_551,N_27920,N_28081);
xor UO_552 (O_552,N_27641,N_29452);
or UO_553 (O_553,N_28303,N_29738);
or UO_554 (O_554,N_27620,N_28541);
or UO_555 (O_555,N_27046,N_27099);
nor UO_556 (O_556,N_28102,N_28093);
or UO_557 (O_557,N_29956,N_27486);
nor UO_558 (O_558,N_28224,N_29049);
or UO_559 (O_559,N_27663,N_28221);
xor UO_560 (O_560,N_28271,N_27343);
xnor UO_561 (O_561,N_28688,N_28654);
nand UO_562 (O_562,N_27109,N_27216);
or UO_563 (O_563,N_29170,N_29477);
or UO_564 (O_564,N_27321,N_27439);
nor UO_565 (O_565,N_28460,N_29795);
or UO_566 (O_566,N_27063,N_28295);
and UO_567 (O_567,N_29102,N_29474);
nor UO_568 (O_568,N_28724,N_27114);
nor UO_569 (O_569,N_27879,N_29813);
and UO_570 (O_570,N_28447,N_28242);
nor UO_571 (O_571,N_28760,N_27386);
xor UO_572 (O_572,N_27340,N_29494);
or UO_573 (O_573,N_27921,N_28314);
xnor UO_574 (O_574,N_27998,N_28964);
nand UO_575 (O_575,N_28128,N_27253);
nand UO_576 (O_576,N_28878,N_29806);
xor UO_577 (O_577,N_29616,N_28960);
and UO_578 (O_578,N_29142,N_27747);
nor UO_579 (O_579,N_28895,N_28055);
nor UO_580 (O_580,N_28825,N_27069);
xor UO_581 (O_581,N_29398,N_29177);
nor UO_582 (O_582,N_29187,N_28442);
nand UO_583 (O_583,N_28382,N_27490);
nor UO_584 (O_584,N_27163,N_29183);
xor UO_585 (O_585,N_29496,N_29184);
and UO_586 (O_586,N_29749,N_28535);
nand UO_587 (O_587,N_29809,N_28625);
and UO_588 (O_588,N_27753,N_27853);
xor UO_589 (O_589,N_29666,N_28967);
nand UO_590 (O_590,N_27021,N_28006);
xnor UO_591 (O_591,N_27165,N_29736);
and UO_592 (O_592,N_29853,N_28198);
nand UO_593 (O_593,N_28236,N_27456);
xor UO_594 (O_594,N_29577,N_28208);
xor UO_595 (O_595,N_27462,N_29818);
and UO_596 (O_596,N_27697,N_28068);
nor UO_597 (O_597,N_27573,N_27200);
nand UO_598 (O_598,N_28753,N_28348);
xor UO_599 (O_599,N_28976,N_27399);
xor UO_600 (O_600,N_29640,N_27067);
nand UO_601 (O_601,N_29511,N_27759);
xor UO_602 (O_602,N_27660,N_28896);
xor UO_603 (O_603,N_29242,N_29414);
nand UO_604 (O_604,N_28948,N_28300);
xnor UO_605 (O_605,N_28350,N_29860);
or UO_606 (O_606,N_29575,N_28090);
nand UO_607 (O_607,N_29553,N_29683);
and UO_608 (O_608,N_28565,N_27661);
xor UO_609 (O_609,N_29306,N_29325);
xor UO_610 (O_610,N_27918,N_29805);
xnor UO_611 (O_611,N_28031,N_29687);
or UO_612 (O_612,N_29263,N_29236);
or UO_613 (O_613,N_28732,N_28182);
nand UO_614 (O_614,N_29268,N_28605);
and UO_615 (O_615,N_28681,N_28641);
xor UO_616 (O_616,N_27617,N_29107);
and UO_617 (O_617,N_27781,N_28669);
or UO_618 (O_618,N_29248,N_28772);
xor UO_619 (O_619,N_28755,N_29927);
or UO_620 (O_620,N_29574,N_29179);
or UO_621 (O_621,N_29303,N_27917);
nor UO_622 (O_622,N_29693,N_27121);
nor UO_623 (O_623,N_28373,N_28210);
and UO_624 (O_624,N_28822,N_28238);
xor UO_625 (O_625,N_28684,N_27594);
xor UO_626 (O_626,N_28059,N_27770);
or UO_627 (O_627,N_29650,N_28616);
or UO_628 (O_628,N_29744,N_27308);
and UO_629 (O_629,N_28276,N_29741);
and UO_630 (O_630,N_29440,N_28114);
xnor UO_631 (O_631,N_28829,N_27159);
and UO_632 (O_632,N_29542,N_28148);
and UO_633 (O_633,N_27615,N_27892);
nand UO_634 (O_634,N_29999,N_27880);
nor UO_635 (O_635,N_29487,N_29517);
xnor UO_636 (O_636,N_29186,N_29567);
xnor UO_637 (O_637,N_29468,N_27442);
xnor UO_638 (O_638,N_27241,N_28942);
and UO_639 (O_639,N_29529,N_27812);
nor UO_640 (O_640,N_27834,N_28370);
and UO_641 (O_641,N_28421,N_27644);
nor UO_642 (O_642,N_27466,N_28092);
nor UO_643 (O_643,N_28649,N_28158);
and UO_644 (O_644,N_27302,N_28254);
and UO_645 (O_645,N_27754,N_29731);
nand UO_646 (O_646,N_27850,N_28752);
nor UO_647 (O_647,N_29111,N_27923);
nor UO_648 (O_648,N_27060,N_27569);
nand UO_649 (O_649,N_28269,N_27336);
and UO_650 (O_650,N_28062,N_27837);
nor UO_651 (O_651,N_27361,N_28591);
or UO_652 (O_652,N_29034,N_29261);
xnor UO_653 (O_653,N_27903,N_27863);
nand UO_654 (O_654,N_27911,N_29094);
and UO_655 (O_655,N_28213,N_28378);
xnor UO_656 (O_656,N_29699,N_28087);
xnor UO_657 (O_657,N_27139,N_27319);
and UO_658 (O_658,N_29310,N_28345);
and UO_659 (O_659,N_29357,N_28121);
and UO_660 (O_660,N_27860,N_29518);
nor UO_661 (O_661,N_28262,N_27971);
xnor UO_662 (O_662,N_28961,N_28953);
xor UO_663 (O_663,N_29718,N_29288);
and UO_664 (O_664,N_29936,N_29933);
and UO_665 (O_665,N_27170,N_28496);
and UO_666 (O_666,N_28905,N_28634);
nand UO_667 (O_667,N_29119,N_27495);
or UO_668 (O_668,N_28333,N_28104);
and UO_669 (O_669,N_29222,N_27698);
or UO_670 (O_670,N_28997,N_28332);
xor UO_671 (O_671,N_28187,N_27529);
or UO_672 (O_672,N_29982,N_29300);
nor UO_673 (O_673,N_29040,N_27630);
nor UO_674 (O_674,N_27005,N_29621);
nor UO_675 (O_675,N_29686,N_29080);
or UO_676 (O_676,N_27571,N_27601);
nor UO_677 (O_677,N_28765,N_29433);
or UO_678 (O_678,N_29218,N_28390);
xnor UO_679 (O_679,N_28493,N_27945);
or UO_680 (O_680,N_28366,N_28455);
xor UO_681 (O_681,N_27394,N_28743);
nand UO_682 (O_682,N_29928,N_29265);
nor UO_683 (O_683,N_28781,N_28650);
and UO_684 (O_684,N_27176,N_27936);
nand UO_685 (O_685,N_29854,N_27807);
nor UO_686 (O_686,N_29537,N_28750);
xnor UO_687 (O_687,N_28018,N_27924);
xor UO_688 (O_688,N_29223,N_27957);
nand UO_689 (O_689,N_29512,N_27287);
nand UO_690 (O_690,N_27405,N_27381);
xor UO_691 (O_691,N_28024,N_29221);
xnor UO_692 (O_692,N_29788,N_27167);
and UO_693 (O_693,N_29852,N_27637);
or UO_694 (O_694,N_29298,N_28981);
nand UO_695 (O_695,N_28417,N_27912);
and UO_696 (O_696,N_27530,N_29624);
xor UO_697 (O_697,N_28096,N_27040);
nand UO_698 (O_698,N_27083,N_28529);
nor UO_699 (O_699,N_29457,N_28970);
or UO_700 (O_700,N_28844,N_28933);
nor UO_701 (O_701,N_29654,N_29564);
and UO_702 (O_702,N_27745,N_29432);
xnor UO_703 (O_703,N_29771,N_27003);
or UO_704 (O_704,N_27675,N_27545);
nand UO_705 (O_705,N_28999,N_27342);
nand UO_706 (O_706,N_27956,N_28162);
or UO_707 (O_707,N_27034,N_28036);
or UO_708 (O_708,N_28575,N_29839);
and UO_709 (O_709,N_28111,N_29322);
or UO_710 (O_710,N_27950,N_27984);
or UO_711 (O_711,N_28330,N_28811);
nand UO_712 (O_712,N_27284,N_27813);
xor UO_713 (O_713,N_29237,N_27916);
nand UO_714 (O_714,N_29875,N_28855);
nand UO_715 (O_715,N_27215,N_27708);
nor UO_716 (O_716,N_27412,N_27713);
nor UO_717 (O_717,N_27702,N_29582);
xor UO_718 (O_718,N_28768,N_29870);
xnor UO_719 (O_719,N_28709,N_28682);
or UO_720 (O_720,N_29258,N_29566);
and UO_721 (O_721,N_29063,N_27491);
and UO_722 (O_722,N_28757,N_29929);
or UO_723 (O_723,N_28834,N_28986);
or UO_724 (O_724,N_29934,N_28568);
xor UO_725 (O_725,N_28980,N_28773);
or UO_726 (O_726,N_28982,N_27135);
and UO_727 (O_727,N_27492,N_28086);
nor UO_728 (O_728,N_29360,N_29311);
nor UO_729 (O_729,N_29593,N_28048);
and UO_730 (O_730,N_27223,N_29041);
and UO_731 (O_731,N_29677,N_27650);
nor UO_732 (O_732,N_28041,N_27232);
and UO_733 (O_733,N_28482,N_27531);
and UO_734 (O_734,N_28697,N_29534);
xnor UO_735 (O_735,N_29727,N_27857);
or UO_736 (O_736,N_29596,N_27323);
and UO_737 (O_737,N_29287,N_29479);
nor UO_738 (O_738,N_27277,N_28494);
and UO_739 (O_739,N_29943,N_29515);
and UO_740 (O_740,N_27968,N_27348);
nor UO_741 (O_741,N_29915,N_28435);
and UO_742 (O_742,N_29476,N_29543);
nand UO_743 (O_743,N_27674,N_27300);
or UO_744 (O_744,N_29863,N_29940);
nor UO_745 (O_745,N_27154,N_29864);
or UO_746 (O_746,N_28443,N_28229);
xor UO_747 (O_747,N_27240,N_27683);
nand UO_748 (O_748,N_29816,N_29907);
xnor UO_749 (O_749,N_27113,N_29373);
or UO_750 (O_750,N_29345,N_27606);
or UO_751 (O_751,N_28701,N_27869);
nor UO_752 (O_752,N_29752,N_28777);
and UO_753 (O_753,N_28935,N_29530);
or UO_754 (O_754,N_28185,N_29659);
xnor UO_755 (O_755,N_27716,N_28882);
nand UO_756 (O_756,N_28319,N_28883);
or UO_757 (O_757,N_29656,N_29785);
and UO_758 (O_758,N_28015,N_27289);
nand UO_759 (O_759,N_29775,N_29158);
xnor UO_760 (O_760,N_27544,N_27191);
or UO_761 (O_761,N_27983,N_27286);
nand UO_762 (O_762,N_29991,N_29026);
xor UO_763 (O_763,N_27390,N_29320);
nor UO_764 (O_764,N_27551,N_27733);
and UO_765 (O_765,N_29068,N_27572);
nand UO_766 (O_766,N_29118,N_27309);
xnor UO_767 (O_767,N_29896,N_28646);
or UO_768 (O_768,N_28858,N_28147);
nor UO_769 (O_769,N_29984,N_27541);
and UO_770 (O_770,N_28735,N_27496);
nor UO_771 (O_771,N_29402,N_29032);
nor UO_772 (O_772,N_28285,N_27339);
nand UO_773 (O_773,N_29009,N_29167);
nand UO_774 (O_774,N_27533,N_29180);
nand UO_775 (O_775,N_29441,N_28320);
or UO_776 (O_776,N_27105,N_27706);
and UO_777 (O_777,N_28747,N_28397);
and UO_778 (O_778,N_27075,N_27285);
and UO_779 (O_779,N_29359,N_28386);
or UO_780 (O_780,N_27846,N_28832);
and UO_781 (O_781,N_27231,N_27411);
and UO_782 (O_782,N_28792,N_28039);
and UO_783 (O_783,N_29762,N_28706);
nand UO_784 (O_784,N_29704,N_27803);
and UO_785 (O_785,N_28911,N_28440);
xnor UO_786 (O_786,N_28078,N_27130);
xor UO_787 (O_787,N_29587,N_28423);
nand UO_788 (O_788,N_27715,N_29227);
nor UO_789 (O_789,N_28186,N_27267);
nor UO_790 (O_790,N_27627,N_29866);
nor UO_791 (O_791,N_29690,N_29714);
nand UO_792 (O_792,N_28630,N_27244);
and UO_793 (O_793,N_27269,N_29913);
nor UO_794 (O_794,N_28406,N_29570);
and UO_795 (O_795,N_29935,N_29109);
nand UO_796 (O_796,N_29060,N_28431);
xnor UO_797 (O_797,N_27961,N_27888);
nor UO_798 (O_798,N_27554,N_28044);
or UO_799 (O_799,N_28864,N_29557);
and UO_800 (O_800,N_29766,N_29965);
nand UO_801 (O_801,N_28854,N_27980);
nor UO_802 (O_802,N_28708,N_27138);
nand UO_803 (O_803,N_27796,N_28247);
and UO_804 (O_804,N_28946,N_28132);
and UO_805 (O_805,N_28222,N_28596);
nor UO_806 (O_806,N_28874,N_29304);
or UO_807 (O_807,N_27851,N_29436);
nand UO_808 (O_808,N_27687,N_28618);
and UO_809 (O_809,N_28532,N_29027);
xnor UO_810 (O_810,N_29614,N_28281);
or UO_811 (O_811,N_29321,N_27050);
or UO_812 (O_812,N_27986,N_29923);
nand UO_813 (O_813,N_28060,N_29299);
nor UO_814 (O_814,N_29324,N_29473);
or UO_815 (O_815,N_29347,N_28172);
nor UO_816 (O_816,N_27934,N_27883);
nand UO_817 (O_817,N_28707,N_27409);
xor UO_818 (O_818,N_27199,N_27449);
nand UO_819 (O_819,N_29330,N_27147);
nand UO_820 (O_820,N_29786,N_29256);
or UO_821 (O_821,N_27410,N_29165);
nor UO_822 (O_822,N_29314,N_27435);
or UO_823 (O_823,N_29319,N_29728);
nand UO_824 (O_824,N_28843,N_27632);
and UO_825 (O_825,N_27186,N_27258);
or UO_826 (O_826,N_27151,N_29856);
xor UO_827 (O_827,N_28346,N_28672);
nand UO_828 (O_828,N_28573,N_27445);
nor UO_829 (O_829,N_27943,N_29381);
nor UO_830 (O_830,N_28137,N_28338);
xor UO_831 (O_831,N_29755,N_29560);
xnor UO_832 (O_832,N_28931,N_27785);
or UO_833 (O_833,N_28108,N_27427);
or UO_834 (O_834,N_28003,N_28628);
nor UO_835 (O_835,N_27416,N_28907);
nand UO_836 (O_836,N_27436,N_28786);
or UO_837 (O_837,N_27808,N_28304);
nor UO_838 (O_838,N_28915,N_29342);
xnor UO_839 (O_839,N_28674,N_28551);
or UO_840 (O_840,N_27694,N_29078);
nand UO_841 (O_841,N_29729,N_28004);
nand UO_842 (O_842,N_29343,N_29162);
xnor UO_843 (O_843,N_29355,N_28292);
nor UO_844 (O_844,N_28388,N_27672);
nand UO_845 (O_845,N_28462,N_27367);
and UO_846 (O_846,N_29701,N_29622);
nand UO_847 (O_847,N_29842,N_27937);
nand UO_848 (O_848,N_28947,N_27695);
xnor UO_849 (O_849,N_28839,N_29830);
and UO_850 (O_850,N_28163,N_28419);
or UO_851 (O_851,N_27522,N_29719);
or UO_852 (O_852,N_27868,N_27652);
and UO_853 (O_853,N_28372,N_29576);
xnor UO_854 (O_854,N_27054,N_29368);
and UO_855 (O_855,N_27876,N_27821);
or UO_856 (O_856,N_29198,N_27729);
xnor UO_857 (O_857,N_27656,N_28237);
nand UO_858 (O_858,N_29706,N_28470);
and UO_859 (O_859,N_29590,N_29911);
xor UO_860 (O_860,N_28731,N_27827);
xnor UO_861 (O_861,N_28119,N_29387);
or UO_862 (O_862,N_27009,N_28870);
nor UO_863 (O_863,N_27582,N_27609);
nand UO_864 (O_864,N_27779,N_28635);
xor UO_865 (O_865,N_28610,N_28949);
xor UO_866 (O_866,N_29386,N_29533);
nand UO_867 (O_867,N_29532,N_27555);
nor UO_868 (O_868,N_27218,N_27438);
nand UO_869 (O_869,N_27610,N_28309);
and UO_870 (O_870,N_27338,N_27975);
nor UO_871 (O_871,N_29619,N_29115);
nand UO_872 (O_872,N_28409,N_27750);
nand UO_873 (O_873,N_27038,N_28754);
and UO_874 (O_874,N_28523,N_29332);
and UO_875 (O_875,N_29781,N_27401);
or UO_876 (O_876,N_29505,N_28488);
xnor UO_877 (O_877,N_27651,N_27297);
nand UO_878 (O_878,N_28751,N_27840);
and UO_879 (O_879,N_28019,N_27999);
and UO_880 (O_880,N_27707,N_29554);
or UO_881 (O_881,N_29296,N_28655);
or UO_882 (O_882,N_27356,N_29285);
nor UO_883 (O_883,N_28748,N_29280);
nor UO_884 (O_884,N_28734,N_27864);
nor UO_885 (O_885,N_27540,N_28884);
or UO_886 (O_886,N_27885,N_27682);
nand UO_887 (O_887,N_29197,N_29208);
or UO_888 (O_888,N_28429,N_29979);
xor UO_889 (O_889,N_29523,N_28270);
nand UO_890 (O_890,N_27173,N_27202);
nor UO_891 (O_891,N_29691,N_28251);
xnor UO_892 (O_892,N_28877,N_27725);
nor UO_893 (O_893,N_29571,N_27519);
nor UO_894 (O_894,N_28057,N_27849);
and UO_895 (O_895,N_29168,N_27521);
xnor UO_896 (O_896,N_28274,N_29132);
xor UO_897 (O_897,N_28841,N_28926);
xor UO_898 (O_898,N_29350,N_27305);
and UO_899 (O_899,N_28762,N_27346);
or UO_900 (O_900,N_29980,N_27510);
nand UO_901 (O_901,N_29276,N_27509);
or UO_902 (O_902,N_27448,N_28972);
nor UO_903 (O_903,N_29028,N_27295);
xor UO_904 (O_904,N_29894,N_27194);
nor UO_905 (O_905,N_28670,N_27621);
nand UO_906 (O_906,N_27250,N_28730);
xnor UO_907 (O_907,N_29064,N_29233);
or UO_908 (O_908,N_28438,N_28871);
xor UO_909 (O_909,N_27798,N_28671);
and UO_910 (O_910,N_29700,N_29763);
or UO_911 (O_911,N_28941,N_29002);
or UO_912 (O_912,N_29410,N_27553);
nand UO_913 (O_913,N_29214,N_29598);
nand UO_914 (O_914,N_29810,N_29658);
xnor UO_915 (O_915,N_29206,N_29977);
nor UO_916 (O_916,N_28555,N_27908);
xor UO_917 (O_917,N_27737,N_27292);
nand UO_918 (O_918,N_27148,N_27301);
nand UO_919 (O_919,N_27472,N_29964);
nand UO_920 (O_920,N_27858,N_27140);
nand UO_921 (O_921,N_27855,N_28538);
and UO_922 (O_922,N_29603,N_27575);
or UO_923 (O_923,N_28957,N_28012);
nand UO_924 (O_924,N_27035,N_29734);
xnor UO_925 (O_925,N_27432,N_28145);
nor UO_926 (O_926,N_29475,N_27623);
nor UO_927 (O_927,N_29046,N_28814);
nand UO_928 (O_928,N_28323,N_27469);
nand UO_929 (O_929,N_27368,N_28468);
nand UO_930 (O_930,N_27266,N_27678);
nand UO_931 (O_931,N_27026,N_29275);
xor UO_932 (O_932,N_28900,N_28107);
nand UO_933 (O_933,N_27181,N_27298);
nand UO_934 (O_934,N_28313,N_29825);
and UO_935 (O_935,N_28054,N_29600);
nand UO_936 (O_936,N_28910,N_29522);
or UO_937 (O_937,N_27585,N_28280);
nand UO_938 (O_938,N_29431,N_29944);
xnor UO_939 (O_939,N_28638,N_28340);
nor UO_940 (O_940,N_29065,N_27922);
xor UO_941 (O_941,N_29243,N_29405);
xnor UO_942 (O_942,N_29146,N_29014);
xor UO_943 (O_943,N_29748,N_29996);
and UO_944 (O_944,N_28673,N_28343);
nor UO_945 (O_945,N_28653,N_28665);
nor UO_946 (O_946,N_27772,N_27893);
and UO_947 (O_947,N_28103,N_29250);
nand UO_948 (O_948,N_29318,N_29873);
nand UO_949 (O_949,N_28993,N_29389);
nor UO_950 (O_950,N_29353,N_29166);
nor UO_951 (O_951,N_28969,N_28795);
or UO_952 (O_952,N_28284,N_29429);
nand UO_953 (O_953,N_29646,N_28539);
xnor UO_954 (O_954,N_28819,N_29838);
nor UO_955 (O_955,N_28885,N_28663);
nand UO_956 (O_956,N_29609,N_29108);
xnor UO_957 (O_957,N_29669,N_27619);
xor UO_958 (O_958,N_27078,N_29694);
xnor UO_959 (O_959,N_27127,N_27769);
nor UO_960 (O_960,N_27414,N_27982);
nand UO_961 (O_961,N_27901,N_28554);
and UO_962 (O_962,N_28838,N_29133);
or UO_963 (O_963,N_29297,N_28050);
nand UO_964 (O_964,N_28116,N_28305);
or UO_965 (O_965,N_29062,N_28584);
nor UO_966 (O_966,N_27767,N_29385);
xor UO_967 (O_967,N_27995,N_27347);
or UO_968 (O_968,N_28395,N_27755);
or UO_969 (O_969,N_27842,N_29145);
nor UO_970 (O_970,N_28857,N_29796);
and UO_971 (O_971,N_29341,N_29067);
or UO_972 (O_972,N_29015,N_27565);
or UO_973 (O_973,N_29105,N_29636);
nor UO_974 (O_974,N_28361,N_29641);
and UO_975 (O_975,N_27959,N_29406);
and UO_976 (O_976,N_29987,N_28011);
nand UO_977 (O_977,N_27684,N_29209);
and UO_978 (O_978,N_27108,N_27538);
nand UO_979 (O_979,N_27593,N_28478);
xor UO_980 (O_980,N_28030,N_28534);
xnor UO_981 (O_981,N_27867,N_28643);
and UO_982 (O_982,N_29377,N_27829);
or UO_983 (O_983,N_27910,N_29213);
nand UO_984 (O_984,N_29226,N_28597);
xnor UO_985 (O_985,N_29290,N_29059);
and UO_986 (O_986,N_27628,N_28561);
nand UO_987 (O_987,N_28847,N_27254);
xor UO_988 (O_988,N_29750,N_28489);
or UO_989 (O_989,N_29612,N_27208);
or UO_990 (O_990,N_29120,N_27665);
and UO_991 (O_991,N_29867,N_29210);
nand UO_992 (O_992,N_29408,N_27776);
nor UO_993 (O_993,N_27424,N_27497);
xnor UO_994 (O_994,N_28831,N_27440);
or UO_995 (O_995,N_28661,N_28917);
or UO_996 (O_996,N_28261,N_27932);
or UO_997 (O_997,N_28277,N_29900);
nor UO_998 (O_998,N_28563,N_27325);
xnor UO_999 (O_999,N_28733,N_28612);
nand UO_1000 (O_1000,N_29931,N_28029);
xor UO_1001 (O_1001,N_27303,N_28862);
xor UO_1002 (O_1002,N_28569,N_28206);
xnor UO_1003 (O_1003,N_27761,N_29053);
xor UO_1004 (O_1004,N_29703,N_29295);
nor UO_1005 (O_1005,N_29922,N_27877);
nor UO_1006 (O_1006,N_27723,N_27460);
nor UO_1007 (O_1007,N_29823,N_27234);
nand UO_1008 (O_1008,N_28231,N_27264);
nand UO_1009 (O_1009,N_29451,N_27242);
or UO_1010 (O_1010,N_29881,N_28830);
or UO_1011 (O_1011,N_29791,N_28842);
nor UO_1012 (O_1012,N_29960,N_28141);
nor UO_1013 (O_1013,N_28385,N_28902);
nor UO_1014 (O_1014,N_28196,N_28835);
nand UO_1015 (O_1015,N_28159,N_29403);
or UO_1016 (O_1016,N_27517,N_27938);
xnor UO_1017 (O_1017,N_29420,N_29581);
nor UO_1018 (O_1018,N_27703,N_27711);
xnor UO_1019 (O_1019,N_29072,N_27430);
xor UO_1020 (O_1020,N_29127,N_27719);
or UO_1021 (O_1021,N_29007,N_28291);
xor UO_1022 (O_1022,N_29602,N_27692);
xor UO_1023 (O_1023,N_27550,N_28246);
nor UO_1024 (O_1024,N_29649,N_29363);
xor UO_1025 (O_1025,N_29559,N_27969);
nand UO_1026 (O_1026,N_29277,N_27275);
and UO_1027 (O_1027,N_28721,N_29425);
nor UO_1028 (O_1028,N_27259,N_28984);
nand UO_1029 (O_1029,N_29130,N_27471);
nor UO_1030 (O_1030,N_28177,N_29066);
and UO_1031 (O_1031,N_28020,N_27457);
xnor UO_1032 (O_1032,N_27116,N_29419);
nand UO_1033 (O_1033,N_27272,N_28130);
xnor UO_1034 (O_1034,N_27142,N_28932);
nand UO_1035 (O_1035,N_29239,N_27091);
xor UO_1036 (O_1036,N_29685,N_27350);
and UO_1037 (O_1037,N_27709,N_28383);
or UO_1038 (O_1038,N_27841,N_29705);
nand UO_1039 (O_1039,N_28171,N_27915);
and UO_1040 (O_1040,N_28873,N_28126);
xor UO_1041 (O_1041,N_28463,N_28921);
or UO_1042 (O_1042,N_28135,N_28647);
xor UO_1043 (O_1043,N_27049,N_27403);
nor UO_1044 (O_1044,N_29083,N_29317);
and UO_1045 (O_1045,N_27493,N_28645);
and UO_1046 (O_1046,N_28802,N_27345);
and UO_1047 (O_1047,N_29461,N_29481);
nand UO_1048 (O_1048,N_29346,N_29820);
nand UO_1049 (O_1049,N_29036,N_29639);
nand UO_1050 (O_1050,N_29493,N_27407);
nor UO_1051 (O_1051,N_27526,N_28800);
nand UO_1052 (O_1052,N_27549,N_27056);
and UO_1053 (O_1053,N_27196,N_27534);
nor UO_1054 (O_1054,N_27441,N_29891);
nand UO_1055 (O_1055,N_29235,N_27001);
nand UO_1056 (O_1056,N_29902,N_27230);
nor UO_1057 (O_1057,N_29019,N_27209);
and UO_1058 (O_1058,N_28950,N_27963);
or UO_1059 (O_1059,N_28106,N_27931);
nand UO_1060 (O_1060,N_27691,N_28193);
or UO_1061 (O_1061,N_27595,N_27417);
xnor UO_1062 (O_1062,N_28188,N_29743);
nor UO_1063 (O_1063,N_29789,N_29774);
and UO_1064 (O_1064,N_28144,N_27415);
or UO_1065 (O_1065,N_27172,N_27947);
nor UO_1066 (O_1066,N_29746,N_27327);
nand UO_1067 (O_1067,N_29990,N_28592);
xor UO_1068 (O_1068,N_28506,N_27581);
nand UO_1069 (O_1069,N_28161,N_29803);
or UO_1070 (O_1070,N_28952,N_28325);
or UO_1071 (O_1071,N_27792,N_29104);
and UO_1072 (O_1072,N_28200,N_28937);
or UO_1073 (O_1073,N_28207,N_29937);
nor UO_1074 (O_1074,N_29017,N_28173);
nor UO_1075 (O_1075,N_29076,N_28317);
or UO_1076 (O_1076,N_27013,N_29697);
nand UO_1077 (O_1077,N_28903,N_28938);
nand UO_1078 (O_1078,N_29089,N_29435);
and UO_1079 (O_1079,N_29759,N_28564);
and UO_1080 (O_1080,N_28627,N_27669);
xnor UO_1081 (O_1081,N_29607,N_27508);
nor UO_1082 (O_1082,N_29272,N_27239);
and UO_1083 (O_1083,N_29500,N_28120);
xor UO_1084 (O_1084,N_28991,N_28746);
or UO_1085 (O_1085,N_28205,N_28658);
or UO_1086 (O_1086,N_27625,N_27370);
xnor UO_1087 (O_1087,N_29975,N_28977);
xnor UO_1088 (O_1088,N_29821,N_28250);
and UO_1089 (O_1089,N_27384,N_27079);
or UO_1090 (O_1090,N_28713,N_29819);
and UO_1091 (O_1091,N_27400,N_28028);
xnor UO_1092 (O_1092,N_27598,N_27580);
and UO_1093 (O_1093,N_27614,N_27062);
xor UO_1094 (O_1094,N_29526,N_29772);
nand UO_1095 (O_1095,N_29680,N_29674);
xor UO_1096 (O_1096,N_29538,N_29364);
and UO_1097 (O_1097,N_28723,N_27704);
and UO_1098 (O_1098,N_27243,N_29339);
nand UO_1099 (O_1099,N_29846,N_27097);
or UO_1100 (O_1100,N_29081,N_29972);
xnor UO_1101 (O_1101,N_27940,N_29961);
nor UO_1102 (O_1102,N_28821,N_27007);
nand UO_1103 (O_1103,N_27187,N_29910);
and UO_1104 (O_1104,N_28889,N_27247);
nand UO_1105 (O_1105,N_29497,N_29630);
nor UO_1106 (O_1106,N_27689,N_28415);
xnor UO_1107 (O_1107,N_27499,N_28852);
nand UO_1108 (O_1108,N_28621,N_29444);
or UO_1109 (O_1109,N_28275,N_27002);
or UO_1110 (O_1110,N_29491,N_28037);
nor UO_1111 (O_1111,N_27514,N_28856);
or UO_1112 (O_1112,N_27220,N_27464);
and UO_1113 (O_1113,N_29608,N_29671);
nor UO_1114 (O_1114,N_27583,N_28389);
xor UO_1115 (O_1115,N_28553,N_27425);
nor UO_1116 (O_1116,N_28579,N_27854);
and UO_1117 (O_1117,N_29462,N_28955);
nor UO_1118 (O_1118,N_29962,N_28444);
xor UO_1119 (O_1119,N_29958,N_27894);
xor UO_1120 (O_1120,N_28897,N_29634);
nand UO_1121 (O_1121,N_28516,N_29254);
nor UO_1122 (O_1122,N_27793,N_27070);
xor UO_1123 (O_1123,N_28778,N_28368);
and UO_1124 (O_1124,N_28583,N_29152);
nand UO_1125 (O_1125,N_27352,N_27131);
nor UO_1126 (O_1126,N_28886,N_29374);
or UO_1127 (O_1127,N_29801,N_29446);
nor UO_1128 (O_1128,N_28365,N_29551);
and UO_1129 (O_1129,N_28204,N_28700);
or UO_1130 (O_1130,N_29588,N_28893);
xnor UO_1131 (O_1131,N_29655,N_27518);
xnor UO_1132 (O_1132,N_29758,N_27461);
xnor UO_1133 (O_1133,N_27679,N_28528);
and UO_1134 (O_1134,N_28608,N_29843);
xnor UO_1135 (O_1135,N_28678,N_27731);
or UO_1136 (O_1136,N_28705,N_27082);
or UO_1137 (O_1137,N_27766,N_28165);
xnor UO_1138 (O_1138,N_29173,N_27115);
and UO_1139 (O_1139,N_28860,N_28101);
and UO_1140 (O_1140,N_29231,N_29631);
or UO_1141 (O_1141,N_28471,N_27935);
and UO_1142 (O_1142,N_28951,N_28098);
nand UO_1143 (O_1143,N_27341,N_27507);
and UO_1144 (O_1144,N_28899,N_29399);
and UO_1145 (O_1145,N_27104,N_28868);
or UO_1146 (O_1146,N_29682,N_27714);
nor UO_1147 (O_1147,N_28117,N_27088);
nor UO_1148 (O_1148,N_27552,N_29327);
nand UO_1149 (O_1149,N_28974,N_28260);
and UO_1150 (O_1150,N_27831,N_28217);
or UO_1151 (O_1151,N_29117,N_27676);
xnor UO_1152 (O_1152,N_27596,N_27800);
and UO_1153 (O_1153,N_28376,N_27238);
nand UO_1154 (O_1154,N_27643,N_27162);
nand UO_1155 (O_1155,N_27160,N_29550);
and UO_1156 (O_1156,N_29006,N_28587);
or UO_1157 (O_1157,N_27721,N_28693);
or UO_1158 (O_1158,N_29754,N_28289);
xor UO_1159 (O_1159,N_28051,N_29747);
xnor UO_1160 (O_1160,N_28567,N_27447);
nor UO_1161 (O_1161,N_28427,N_27357);
xor UO_1162 (O_1162,N_27205,N_29792);
xnor UO_1163 (O_1163,N_29668,N_29114);
or UO_1164 (O_1164,N_27646,N_27030);
nand UO_1165 (O_1165,N_28756,N_28639);
or UO_1166 (O_1166,N_27431,N_29100);
nand UO_1167 (O_1167,N_28501,N_28863);
or UO_1168 (O_1168,N_28140,N_29361);
nand UO_1169 (O_1169,N_27353,N_27333);
and UO_1170 (O_1170,N_27543,N_29586);
or UO_1171 (O_1171,N_29212,N_27954);
nand UO_1172 (O_1172,N_29974,N_29099);
nor UO_1173 (O_1173,N_28687,N_28094);
nor UO_1174 (O_1174,N_29486,N_27668);
nand UO_1175 (O_1175,N_27700,N_29985);
nor UO_1176 (O_1176,N_28975,N_29597);
or UO_1177 (O_1177,N_27948,N_28922);
xnor UO_1178 (O_1178,N_28357,N_28696);
xnor UO_1179 (O_1179,N_27059,N_27288);
or UO_1180 (O_1180,N_27577,N_29018);
nand UO_1181 (O_1181,N_29601,N_28184);
nor UO_1182 (O_1182,N_29380,N_27654);
and UO_1183 (O_1183,N_27189,N_29442);
nand UO_1184 (O_1184,N_29756,N_28861);
xor UO_1185 (O_1185,N_29073,N_29264);
nand UO_1186 (O_1186,N_29814,N_27397);
nand UO_1187 (O_1187,N_28461,N_28129);
nand UO_1188 (O_1188,N_27503,N_28540);
nor UO_1189 (O_1189,N_28155,N_29708);
or UO_1190 (O_1190,N_27758,N_28021);
nand UO_1191 (O_1191,N_28689,N_28001);
xor UO_1192 (O_1192,N_29966,N_28477);
nand UO_1193 (O_1193,N_29673,N_28257);
nand UO_1194 (O_1194,N_28279,N_28294);
or UO_1195 (O_1195,N_28034,N_27742);
and UO_1196 (O_1196,N_28079,N_28533);
xor UO_1197 (O_1197,N_28598,N_28404);
or UO_1198 (O_1198,N_27930,N_27591);
nor UO_1199 (O_1199,N_29969,N_29471);
xnor UO_1200 (O_1200,N_28077,N_27349);
or UO_1201 (O_1201,N_27556,N_27149);
xnor UO_1202 (O_1202,N_27364,N_27299);
or UO_1203 (O_1203,N_27653,N_29354);
or UO_1204 (O_1204,N_27870,N_27408);
or UO_1205 (O_1205,N_28593,N_29606);
or UO_1206 (O_1206,N_27252,N_28306);
and UO_1207 (O_1207,N_29887,N_29394);
nand UO_1208 (O_1208,N_27563,N_27053);
or UO_1209 (O_1209,N_29273,N_27193);
or UO_1210 (O_1210,N_27976,N_27710);
or UO_1211 (O_1211,N_27016,N_29845);
nor UO_1212 (O_1212,N_29976,N_29716);
and UO_1213 (O_1213,N_27373,N_28978);
nand UO_1214 (O_1214,N_27659,N_28066);
xor UO_1215 (O_1215,N_29459,N_29085);
or UO_1216 (O_1216,N_28453,N_28968);
xor UO_1217 (O_1217,N_28381,N_27136);
xnor UO_1218 (O_1218,N_27004,N_28560);
xor UO_1219 (O_1219,N_27933,N_29967);
xor UO_1220 (O_1220,N_27906,N_29800);
and UO_1221 (O_1221,N_29000,N_27306);
and UO_1222 (O_1222,N_27129,N_28629);
and UO_1223 (O_1223,N_28875,N_28939);
nor UO_1224 (O_1224,N_29828,N_27029);
and UO_1225 (O_1225,N_27757,N_27385);
xor UO_1226 (O_1226,N_29141,N_29815);
nand UO_1227 (O_1227,N_29776,N_28623);
nand UO_1228 (O_1228,N_29610,N_28446);
or UO_1229 (O_1229,N_29369,N_29058);
and UO_1230 (O_1230,N_28574,N_27320);
xor UO_1231 (O_1231,N_29773,N_28290);
xnor UO_1232 (O_1232,N_29143,N_27717);
nor UO_1233 (O_1233,N_27639,N_28416);
xnor UO_1234 (O_1234,N_29008,N_27558);
xor UO_1235 (O_1235,N_29545,N_28881);
or UO_1236 (O_1236,N_28512,N_29286);
nand UO_1237 (O_1237,N_28095,N_28405);
nand UO_1238 (O_1238,N_27847,N_28178);
or UO_1239 (O_1239,N_27802,N_28218);
or UO_1240 (O_1240,N_27351,N_28711);
xor UO_1241 (O_1241,N_28014,N_29908);
xor UO_1242 (O_1242,N_27085,N_28253);
and UO_1243 (O_1243,N_29367,N_29737);
or UO_1244 (O_1244,N_27222,N_29292);
nor UO_1245 (O_1245,N_28481,N_27548);
nand UO_1246 (O_1246,N_29909,N_27280);
nand UO_1247 (O_1247,N_29483,N_27330);
xor UO_1248 (O_1248,N_27587,N_27997);
and UO_1249 (O_1249,N_28214,N_28518);
nand UO_1250 (O_1250,N_28360,N_29877);
and UO_1251 (O_1251,N_27820,N_29521);
nor UO_1252 (O_1252,N_28038,N_28962);
xor UO_1253 (O_1253,N_27111,N_28572);
and UO_1254 (O_1254,N_29030,N_29464);
or UO_1255 (O_1255,N_29039,N_28362);
and UO_1256 (O_1256,N_29970,N_28779);
nor UO_1257 (O_1257,N_29675,N_27881);
or UO_1258 (O_1258,N_28659,N_27788);
xnor UO_1259 (O_1259,N_28566,N_29520);
nand UO_1260 (O_1260,N_28239,N_27119);
xnor UO_1261 (O_1261,N_28657,N_29798);
or UO_1262 (O_1262,N_27249,N_27539);
or UO_1263 (O_1263,N_27728,N_29721);
or UO_1264 (O_1264,N_27871,N_27799);
and UO_1265 (O_1265,N_29832,N_28228);
nor UO_1266 (O_1266,N_27422,N_28312);
nor UO_1267 (O_1267,N_29383,N_29885);
or UO_1268 (O_1268,N_29536,N_27271);
or UO_1269 (O_1269,N_27478,N_28581);
nand UO_1270 (O_1270,N_29284,N_29282);
and UO_1271 (O_1271,N_27958,N_28771);
xor UO_1272 (O_1272,N_28268,N_28718);
and UO_1273 (O_1273,N_29787,N_27174);
nor UO_1274 (O_1274,N_28310,N_29540);
nor UO_1275 (O_1275,N_27987,N_29778);
nand UO_1276 (O_1276,N_28469,N_29224);
xor UO_1277 (O_1277,N_29098,N_27443);
or UO_1278 (O_1278,N_28451,N_29193);
xor UO_1279 (O_1279,N_29348,N_28318);
nor UO_1280 (O_1280,N_28851,N_27902);
and UO_1281 (O_1281,N_29182,N_27886);
nand UO_1282 (O_1282,N_28507,N_29707);
xor UO_1283 (O_1283,N_28514,N_27064);
xor UO_1284 (O_1284,N_29196,N_27815);
nand UO_1285 (O_1285,N_27093,N_28083);
or UO_1286 (O_1286,N_29011,N_27666);
xor UO_1287 (O_1287,N_29485,N_29326);
xnor UO_1288 (O_1288,N_29416,N_28717);
nand UO_1289 (O_1289,N_27315,N_29156);
nor UO_1290 (O_1290,N_28076,N_27426);
and UO_1291 (O_1291,N_27036,N_28152);
or UO_1292 (O_1292,N_28827,N_29232);
nand UO_1293 (O_1293,N_27454,N_29071);
and UO_1294 (O_1294,N_28393,N_27516);
nor UO_1295 (O_1295,N_29281,N_27092);
nand UO_1296 (O_1296,N_28662,N_27744);
and UO_1297 (O_1297,N_29220,N_29069);
and UO_1298 (O_1298,N_28611,N_29561);
xor UO_1299 (O_1299,N_29552,N_28513);
or UO_1300 (O_1300,N_27331,N_28766);
or UO_1301 (O_1301,N_27568,N_29247);
and UO_1302 (O_1302,N_29599,N_28301);
and UO_1303 (O_1303,N_27025,N_27979);
xnor UO_1304 (O_1304,N_27929,N_28769);
xnor UO_1305 (O_1305,N_28009,N_28190);
and UO_1306 (O_1306,N_27074,N_27195);
xnor UO_1307 (O_1307,N_27090,N_28189);
nor UO_1308 (O_1308,N_29396,N_27474);
xnor UO_1309 (O_1309,N_28979,N_28588);
xnor UO_1310 (O_1310,N_29524,N_27626);
nor UO_1311 (O_1311,N_27080,N_29427);
and UO_1312 (O_1312,N_27118,N_29050);
nor UO_1313 (O_1313,N_28258,N_28966);
nor UO_1314 (O_1314,N_28890,N_27073);
nand UO_1315 (O_1315,N_28324,N_28812);
and UO_1316 (O_1316,N_27086,N_28017);
and UO_1317 (O_1317,N_29289,N_28694);
nor UO_1318 (O_1318,N_28633,N_28691);
xor UO_1319 (O_1319,N_29799,N_27953);
and UO_1320 (O_1320,N_29128,N_28887);
nand UO_1321 (O_1321,N_27023,N_27763);
or UO_1322 (O_1322,N_27739,N_27488);
or UO_1323 (O_1323,N_27905,N_28115);
nand UO_1324 (O_1324,N_28940,N_28578);
nor UO_1325 (O_1325,N_29632,N_29696);
and UO_1326 (O_1326,N_28191,N_28179);
nand UO_1327 (O_1327,N_27732,N_28594);
nor UO_1328 (O_1328,N_28358,N_29633);
nor UO_1329 (O_1329,N_27134,N_28923);
and UO_1330 (O_1330,N_28351,N_27790);
or UO_1331 (O_1331,N_29316,N_28384);
or UO_1332 (O_1332,N_28392,N_29400);
nor UO_1333 (O_1333,N_28492,N_29244);
and UO_1334 (O_1334,N_27688,N_27925);
and UO_1335 (O_1335,N_28840,N_28853);
nand UO_1336 (O_1336,N_27126,N_28626);
nand UO_1337 (O_1337,N_28399,N_29021);
nor UO_1338 (O_1338,N_27450,N_27574);
or UO_1339 (O_1339,N_29090,N_28589);
nor UO_1340 (O_1340,N_29336,N_27166);
and UO_1341 (O_1341,N_27273,N_28904);
nand UO_1342 (O_1342,N_27973,N_28774);
or UO_1343 (O_1343,N_27988,N_29509);
and UO_1344 (O_1344,N_27942,N_29635);
nor UO_1345 (O_1345,N_29765,N_29745);
nor UO_1346 (O_1346,N_28736,N_27380);
xnor UO_1347 (O_1347,N_29698,N_28595);
and UO_1348 (O_1348,N_27889,N_27502);
nand UO_1349 (O_1349,N_29625,N_28992);
xor UO_1350 (O_1350,N_28369,N_29047);
nand UO_1351 (O_1351,N_27657,N_28142);
xor UO_1352 (O_1352,N_28548,N_27335);
and UO_1353 (O_1353,N_29742,N_28954);
xor UO_1354 (O_1354,N_29822,N_27322);
and UO_1355 (O_1355,N_29472,N_29657);
and UO_1356 (O_1356,N_29709,N_29309);
nand UO_1357 (O_1357,N_27296,N_29228);
and UO_1358 (O_1358,N_29116,N_28331);
nand UO_1359 (O_1359,N_29849,N_28929);
nand UO_1360 (O_1360,N_27771,N_27084);
xnor UO_1361 (O_1361,N_29456,N_27233);
nand UO_1362 (O_1362,N_29135,N_29807);
nand UO_1363 (O_1363,N_29219,N_28525);
or UO_1364 (O_1364,N_29092,N_29770);
xnor UO_1365 (O_1365,N_28824,N_28439);
or UO_1366 (O_1366,N_29722,N_27101);
and UO_1367 (O_1367,N_28715,N_27746);
or UO_1368 (O_1368,N_27369,N_28154);
nor UO_1369 (O_1369,N_28898,N_28353);
or UO_1370 (O_1370,N_28202,N_27760);
or UO_1371 (O_1371,N_29827,N_29409);
xnor UO_1372 (O_1372,N_29651,N_28556);
xnor UO_1373 (O_1373,N_29200,N_28749);
and UO_1374 (O_1374,N_28622,N_28818);
xnor UO_1375 (O_1375,N_28784,N_27363);
and UO_1376 (O_1376,N_29460,N_28080);
nor UO_1377 (O_1377,N_29154,N_28526);
xnor UO_1378 (O_1378,N_29216,N_27226);
xor UO_1379 (O_1379,N_28503,N_28151);
nor UO_1380 (O_1380,N_28666,N_28058);
xnor UO_1381 (O_1381,N_27844,N_29371);
xnor UO_1382 (O_1382,N_29953,N_28072);
xor UO_1383 (O_1383,N_28071,N_27402);
nor UO_1384 (O_1384,N_28667,N_28045);
and UO_1385 (O_1385,N_29948,N_29439);
xor UO_1386 (O_1386,N_29149,N_28448);
nand UO_1387 (O_1387,N_28424,N_29925);
and UO_1388 (O_1388,N_27355,N_28745);
nand UO_1389 (O_1389,N_27190,N_28988);
and UO_1390 (O_1390,N_27629,N_29688);
nor UO_1391 (O_1391,N_27033,N_28099);
nand UO_1392 (O_1392,N_29811,N_28209);
nand UO_1393 (O_1393,N_29225,N_27391);
nand UO_1394 (O_1394,N_29194,N_27446);
xnor UO_1395 (O_1395,N_29890,N_29672);
or UO_1396 (O_1396,N_28963,N_28266);
and UO_1397 (O_1397,N_27589,N_29862);
xor UO_1398 (O_1398,N_27372,N_29378);
nand UO_1399 (O_1399,N_29879,N_28552);
xnor UO_1400 (O_1400,N_27818,N_29238);
nor UO_1401 (O_1401,N_28995,N_27278);
nand UO_1402 (O_1402,N_28053,N_28601);
and UO_1403 (O_1403,N_28056,N_28613);
or UO_1404 (O_1404,N_27065,N_28880);
nor UO_1405 (O_1405,N_27366,N_28876);
nor UO_1406 (O_1406,N_28287,N_27255);
and UO_1407 (O_1407,N_29850,N_29013);
nor UO_1408 (O_1408,N_28676,N_29086);
nand UO_1409 (O_1409,N_29541,N_28632);
xor UO_1410 (O_1410,N_29876,N_27124);
nand UO_1411 (O_1411,N_27019,N_28259);
or UO_1412 (O_1412,N_27900,N_27655);
xor UO_1413 (O_1413,N_29892,N_29824);
or UO_1414 (O_1414,N_29202,N_29044);
xor UO_1415 (O_1415,N_29905,N_27817);
nand UO_1416 (O_1416,N_27501,N_28726);
and UO_1417 (O_1417,N_27537,N_29920);
nand UO_1418 (O_1418,N_28936,N_27809);
nand UO_1419 (O_1419,N_28432,N_28476);
xor UO_1420 (O_1420,N_29968,N_27022);
or UO_1421 (O_1421,N_29751,N_27546);
xor UO_1422 (O_1422,N_29415,N_28061);
or UO_1423 (O_1423,N_28803,N_28131);
nand UO_1424 (O_1424,N_27318,N_27724);
xor UO_1425 (O_1425,N_27602,N_28398);
nor UO_1426 (O_1426,N_29097,N_29490);
xor UO_1427 (O_1427,N_28664,N_28375);
nor UO_1428 (O_1428,N_29782,N_27452);
nor UO_1429 (O_1429,N_27762,N_28837);
nor UO_1430 (O_1430,N_29528,N_29548);
and UO_1431 (O_1431,N_27839,N_29858);
nor UO_1432 (O_1432,N_29804,N_28849);
and UO_1433 (O_1433,N_29417,N_28016);
and UO_1434 (O_1434,N_29504,N_28308);
and UO_1435 (O_1435,N_29012,N_28695);
nand UO_1436 (O_1436,N_29229,N_29240);
nor UO_1437 (O_1437,N_29334,N_28327);
xor UO_1438 (O_1438,N_29362,N_29893);
and UO_1439 (O_1439,N_27498,N_27897);
and UO_1440 (O_1440,N_27740,N_28181);
nand UO_1441 (O_1441,N_28387,N_27965);
and UO_1442 (O_1442,N_28230,N_27603);
nand UO_1443 (O_1443,N_29768,N_27237);
nor UO_1444 (O_1444,N_27310,N_28175);
nor UO_1445 (O_1445,N_29645,N_29337);
and UO_1446 (O_1446,N_27532,N_29652);
and UO_1447 (O_1447,N_29949,N_28714);
and UO_1448 (O_1448,N_27890,N_27824);
nand UO_1449 (O_1449,N_29079,N_29794);
or UO_1450 (O_1450,N_28122,N_27098);
and UO_1451 (O_1451,N_27634,N_29868);
xor UO_1452 (O_1452,N_27896,N_29323);
xnor UO_1453 (O_1453,N_27605,N_29437);
xnor UO_1454 (O_1454,N_27789,N_28741);
xor UO_1455 (O_1455,N_27045,N_28580);
or UO_1456 (O_1456,N_28683,N_28326);
and UO_1457 (O_1457,N_29764,N_27730);
or UO_1458 (O_1458,N_27122,N_27814);
xnor UO_1459 (O_1459,N_27597,N_28600);
and UO_1460 (O_1460,N_29103,N_27699);
xor UO_1461 (O_1461,N_28450,N_29428);
or UO_1462 (O_1462,N_28690,N_28153);
or UO_1463 (O_1463,N_28143,N_29753);
nor UO_1464 (O_1464,N_27604,N_29307);
nor UO_1465 (O_1465,N_29349,N_29189);
xor UO_1466 (O_1466,N_27156,N_28973);
xor UO_1467 (O_1467,N_27542,N_29562);
xor UO_1468 (O_1468,N_28775,N_29488);
nand UO_1469 (O_1469,N_29503,N_27828);
nor UO_1470 (O_1470,N_29495,N_28170);
or UO_1471 (O_1471,N_29412,N_27748);
or UO_1472 (O_1472,N_27276,N_28040);
or UO_1473 (O_1473,N_27404,N_27962);
nor UO_1474 (O_1474,N_27146,N_27681);
nand UO_1475 (O_1475,N_28233,N_28474);
or UO_1476 (O_1476,N_27120,N_27852);
or UO_1477 (O_1477,N_27825,N_28521);
nand UO_1478 (O_1478,N_29125,N_29954);
or UO_1479 (O_1479,N_28073,N_28499);
or UO_1480 (O_1480,N_27332,N_28785);
xor UO_1481 (O_1481,N_28296,N_28500);
xor UO_1482 (O_1482,N_29029,N_28199);
and UO_1483 (O_1483,N_29992,N_27489);
and UO_1484 (O_1484,N_28913,N_29957);
and UO_1485 (O_1485,N_28328,N_29466);
xnor UO_1486 (O_1486,N_29679,N_27941);
nand UO_1487 (O_1487,N_29043,N_27964);
xor UO_1488 (O_1488,N_29393,N_29174);
nand UO_1489 (O_1489,N_27225,N_28013);
nand UO_1490 (O_1490,N_28677,N_29926);
xnor UO_1491 (O_1491,N_27221,N_28586);
or UO_1492 (O_1492,N_27006,N_29725);
nand UO_1493 (O_1493,N_28796,N_27041);
nor UO_1494 (O_1494,N_27909,N_28354);
or UO_1495 (O_1495,N_28797,N_28912);
or UO_1496 (O_1496,N_28798,N_27823);
nor UO_1497 (O_1497,N_28740,N_28710);
nand UO_1498 (O_1498,N_29836,N_29857);
nor UO_1499 (O_1499,N_28411,N_28495);
nand UO_1500 (O_1500,N_27755,N_28125);
xor UO_1501 (O_1501,N_27718,N_27894);
or UO_1502 (O_1502,N_27658,N_29466);
or UO_1503 (O_1503,N_29359,N_28016);
nor UO_1504 (O_1504,N_29243,N_28340);
or UO_1505 (O_1505,N_27316,N_29031);
and UO_1506 (O_1506,N_28505,N_28603);
nor UO_1507 (O_1507,N_27748,N_27833);
or UO_1508 (O_1508,N_27068,N_27438);
nor UO_1509 (O_1509,N_28385,N_29324);
nand UO_1510 (O_1510,N_28892,N_28863);
or UO_1511 (O_1511,N_27398,N_29298);
nand UO_1512 (O_1512,N_27315,N_29258);
nand UO_1513 (O_1513,N_27307,N_28551);
xnor UO_1514 (O_1514,N_28804,N_29355);
nor UO_1515 (O_1515,N_29279,N_28161);
nand UO_1516 (O_1516,N_28376,N_28570);
and UO_1517 (O_1517,N_29541,N_29407);
and UO_1518 (O_1518,N_28413,N_29705);
or UO_1519 (O_1519,N_27653,N_27310);
nor UO_1520 (O_1520,N_28298,N_28469);
nand UO_1521 (O_1521,N_29579,N_27790);
and UO_1522 (O_1522,N_28174,N_27520);
and UO_1523 (O_1523,N_29445,N_29677);
and UO_1524 (O_1524,N_27437,N_28119);
nor UO_1525 (O_1525,N_29135,N_28404);
xor UO_1526 (O_1526,N_28177,N_28611);
nand UO_1527 (O_1527,N_27452,N_29927);
nor UO_1528 (O_1528,N_28390,N_27992);
or UO_1529 (O_1529,N_29065,N_27564);
xnor UO_1530 (O_1530,N_29770,N_28628);
xnor UO_1531 (O_1531,N_29809,N_29227);
nand UO_1532 (O_1532,N_27248,N_27048);
nor UO_1533 (O_1533,N_29886,N_27925);
or UO_1534 (O_1534,N_27961,N_29255);
nor UO_1535 (O_1535,N_28008,N_28636);
nand UO_1536 (O_1536,N_27707,N_27681);
or UO_1537 (O_1537,N_27103,N_29834);
xor UO_1538 (O_1538,N_28453,N_28962);
or UO_1539 (O_1539,N_27787,N_29716);
or UO_1540 (O_1540,N_27832,N_28670);
and UO_1541 (O_1541,N_27166,N_28133);
and UO_1542 (O_1542,N_27616,N_28775);
xor UO_1543 (O_1543,N_29890,N_28612);
and UO_1544 (O_1544,N_29399,N_27296);
and UO_1545 (O_1545,N_27501,N_29872);
and UO_1546 (O_1546,N_29199,N_28456);
and UO_1547 (O_1547,N_28499,N_29872);
or UO_1548 (O_1548,N_27414,N_27736);
nor UO_1549 (O_1549,N_29342,N_28930);
xor UO_1550 (O_1550,N_29264,N_27036);
nand UO_1551 (O_1551,N_29569,N_27597);
and UO_1552 (O_1552,N_29400,N_29203);
xnor UO_1553 (O_1553,N_28197,N_29678);
or UO_1554 (O_1554,N_27789,N_29813);
nand UO_1555 (O_1555,N_27458,N_27546);
nand UO_1556 (O_1556,N_27119,N_28599);
xor UO_1557 (O_1557,N_28769,N_29881);
and UO_1558 (O_1558,N_29002,N_28302);
xor UO_1559 (O_1559,N_28731,N_29886);
nor UO_1560 (O_1560,N_28284,N_28918);
or UO_1561 (O_1561,N_27486,N_27363);
nor UO_1562 (O_1562,N_29719,N_27517);
and UO_1563 (O_1563,N_27584,N_28105);
and UO_1564 (O_1564,N_29443,N_28622);
nand UO_1565 (O_1565,N_28911,N_29885);
or UO_1566 (O_1566,N_29670,N_29507);
xnor UO_1567 (O_1567,N_28524,N_28958);
or UO_1568 (O_1568,N_27645,N_27841);
or UO_1569 (O_1569,N_29587,N_28531);
nor UO_1570 (O_1570,N_28694,N_29308);
or UO_1571 (O_1571,N_27443,N_27915);
or UO_1572 (O_1572,N_28236,N_27728);
nor UO_1573 (O_1573,N_28414,N_29204);
xnor UO_1574 (O_1574,N_29168,N_29389);
and UO_1575 (O_1575,N_28140,N_27702);
xnor UO_1576 (O_1576,N_27203,N_27126);
nor UO_1577 (O_1577,N_27373,N_29727);
or UO_1578 (O_1578,N_28141,N_27236);
xor UO_1579 (O_1579,N_28124,N_28713);
xnor UO_1580 (O_1580,N_27515,N_29621);
or UO_1581 (O_1581,N_28460,N_28276);
xnor UO_1582 (O_1582,N_28133,N_27169);
or UO_1583 (O_1583,N_29836,N_29742);
nor UO_1584 (O_1584,N_28654,N_28515);
xor UO_1585 (O_1585,N_27388,N_29257);
or UO_1586 (O_1586,N_29843,N_28339);
xor UO_1587 (O_1587,N_28019,N_27769);
and UO_1588 (O_1588,N_29425,N_29917);
xnor UO_1589 (O_1589,N_29537,N_28927);
and UO_1590 (O_1590,N_29488,N_28619);
and UO_1591 (O_1591,N_27127,N_28037);
nor UO_1592 (O_1592,N_27269,N_27167);
or UO_1593 (O_1593,N_28429,N_29420);
nor UO_1594 (O_1594,N_27106,N_27942);
nor UO_1595 (O_1595,N_29168,N_27797);
xor UO_1596 (O_1596,N_29568,N_27380);
or UO_1597 (O_1597,N_28948,N_29038);
nor UO_1598 (O_1598,N_27572,N_29457);
and UO_1599 (O_1599,N_28132,N_27497);
nand UO_1600 (O_1600,N_28208,N_29312);
nand UO_1601 (O_1601,N_27648,N_29439);
xor UO_1602 (O_1602,N_27718,N_27934);
nand UO_1603 (O_1603,N_29254,N_27743);
or UO_1604 (O_1604,N_28964,N_27878);
or UO_1605 (O_1605,N_28601,N_28450);
xor UO_1606 (O_1606,N_28873,N_27012);
nand UO_1607 (O_1607,N_27669,N_28647);
or UO_1608 (O_1608,N_27246,N_29075);
or UO_1609 (O_1609,N_28748,N_29363);
nand UO_1610 (O_1610,N_27620,N_28184);
and UO_1611 (O_1611,N_28819,N_27687);
and UO_1612 (O_1612,N_29240,N_27122);
nor UO_1613 (O_1613,N_27469,N_27150);
or UO_1614 (O_1614,N_29979,N_28297);
nor UO_1615 (O_1615,N_28696,N_27354);
nor UO_1616 (O_1616,N_28534,N_27799);
nor UO_1617 (O_1617,N_29300,N_28070);
or UO_1618 (O_1618,N_27533,N_29435);
nand UO_1619 (O_1619,N_27531,N_29106);
xor UO_1620 (O_1620,N_27769,N_27093);
and UO_1621 (O_1621,N_27859,N_29874);
and UO_1622 (O_1622,N_27193,N_28606);
nor UO_1623 (O_1623,N_29116,N_29525);
nor UO_1624 (O_1624,N_29044,N_27303);
or UO_1625 (O_1625,N_29160,N_27737);
nand UO_1626 (O_1626,N_29484,N_27932);
or UO_1627 (O_1627,N_29586,N_28421);
nor UO_1628 (O_1628,N_29317,N_28552);
or UO_1629 (O_1629,N_27134,N_29782);
nor UO_1630 (O_1630,N_28105,N_28071);
xor UO_1631 (O_1631,N_27157,N_27161);
nand UO_1632 (O_1632,N_27414,N_29829);
xor UO_1633 (O_1633,N_27855,N_28413);
nand UO_1634 (O_1634,N_27632,N_27945);
nand UO_1635 (O_1635,N_28644,N_27783);
or UO_1636 (O_1636,N_29212,N_28794);
nand UO_1637 (O_1637,N_29949,N_28116);
nor UO_1638 (O_1638,N_27740,N_28769);
or UO_1639 (O_1639,N_29721,N_28017);
and UO_1640 (O_1640,N_27130,N_28536);
nor UO_1641 (O_1641,N_27335,N_28898);
and UO_1642 (O_1642,N_29263,N_27876);
nand UO_1643 (O_1643,N_27091,N_27370);
and UO_1644 (O_1644,N_28814,N_27760);
nand UO_1645 (O_1645,N_29608,N_29778);
or UO_1646 (O_1646,N_29022,N_27222);
nor UO_1647 (O_1647,N_29076,N_29014);
xor UO_1648 (O_1648,N_29780,N_28377);
nand UO_1649 (O_1649,N_28547,N_27106);
nor UO_1650 (O_1650,N_29542,N_27231);
nor UO_1651 (O_1651,N_28207,N_28987);
or UO_1652 (O_1652,N_27164,N_29547);
nor UO_1653 (O_1653,N_29840,N_28342);
xor UO_1654 (O_1654,N_28190,N_27989);
xnor UO_1655 (O_1655,N_29948,N_28035);
nor UO_1656 (O_1656,N_29794,N_28407);
and UO_1657 (O_1657,N_27133,N_27927);
xnor UO_1658 (O_1658,N_28166,N_28680);
nor UO_1659 (O_1659,N_27685,N_29858);
xnor UO_1660 (O_1660,N_29367,N_27075);
or UO_1661 (O_1661,N_28076,N_29841);
xnor UO_1662 (O_1662,N_29722,N_29916);
or UO_1663 (O_1663,N_27793,N_27876);
nand UO_1664 (O_1664,N_27345,N_28496);
or UO_1665 (O_1665,N_29888,N_28079);
or UO_1666 (O_1666,N_29025,N_27320);
nor UO_1667 (O_1667,N_27467,N_27072);
nand UO_1668 (O_1668,N_28408,N_29335);
nor UO_1669 (O_1669,N_29406,N_28645);
and UO_1670 (O_1670,N_28794,N_27146);
nand UO_1671 (O_1671,N_27490,N_28586);
xor UO_1672 (O_1672,N_29911,N_28734);
and UO_1673 (O_1673,N_29520,N_27990);
or UO_1674 (O_1674,N_29095,N_29120);
xor UO_1675 (O_1675,N_27579,N_28315);
nor UO_1676 (O_1676,N_29570,N_29404);
and UO_1677 (O_1677,N_27736,N_28331);
nand UO_1678 (O_1678,N_29645,N_28920);
or UO_1679 (O_1679,N_29993,N_28841);
nand UO_1680 (O_1680,N_28339,N_29577);
nor UO_1681 (O_1681,N_28165,N_29170);
nand UO_1682 (O_1682,N_29165,N_28500);
and UO_1683 (O_1683,N_29955,N_28637);
and UO_1684 (O_1684,N_29323,N_29495);
nand UO_1685 (O_1685,N_27245,N_28661);
nor UO_1686 (O_1686,N_27070,N_27620);
nand UO_1687 (O_1687,N_27046,N_29062);
and UO_1688 (O_1688,N_27178,N_27055);
and UO_1689 (O_1689,N_29869,N_28248);
or UO_1690 (O_1690,N_29889,N_29869);
nand UO_1691 (O_1691,N_29996,N_28659);
nand UO_1692 (O_1692,N_28757,N_27522);
nor UO_1693 (O_1693,N_28146,N_28233);
nand UO_1694 (O_1694,N_29745,N_27414);
xnor UO_1695 (O_1695,N_29930,N_29702);
nand UO_1696 (O_1696,N_29887,N_29278);
xnor UO_1697 (O_1697,N_28346,N_29440);
nand UO_1698 (O_1698,N_28463,N_27976);
nand UO_1699 (O_1699,N_27509,N_28133);
nand UO_1700 (O_1700,N_29230,N_27082);
nor UO_1701 (O_1701,N_29332,N_29698);
or UO_1702 (O_1702,N_28645,N_29504);
or UO_1703 (O_1703,N_28632,N_27792);
xnor UO_1704 (O_1704,N_29473,N_29371);
nor UO_1705 (O_1705,N_29242,N_27604);
nand UO_1706 (O_1706,N_28002,N_27601);
nand UO_1707 (O_1707,N_29307,N_29454);
or UO_1708 (O_1708,N_27955,N_28129);
and UO_1709 (O_1709,N_27647,N_29200);
or UO_1710 (O_1710,N_28562,N_27656);
nand UO_1711 (O_1711,N_28451,N_28121);
nand UO_1712 (O_1712,N_29349,N_29413);
nor UO_1713 (O_1713,N_27264,N_27551);
xor UO_1714 (O_1714,N_29539,N_27007);
xor UO_1715 (O_1715,N_28315,N_28960);
xnor UO_1716 (O_1716,N_27624,N_29367);
nor UO_1717 (O_1717,N_28019,N_28486);
or UO_1718 (O_1718,N_29677,N_28942);
or UO_1719 (O_1719,N_28630,N_27975);
nor UO_1720 (O_1720,N_27924,N_28892);
nand UO_1721 (O_1721,N_29125,N_27295);
and UO_1722 (O_1722,N_29561,N_28535);
nor UO_1723 (O_1723,N_29847,N_27196);
xor UO_1724 (O_1724,N_29323,N_29215);
or UO_1725 (O_1725,N_29939,N_29150);
or UO_1726 (O_1726,N_29828,N_27866);
nor UO_1727 (O_1727,N_27240,N_27430);
or UO_1728 (O_1728,N_28250,N_27835);
and UO_1729 (O_1729,N_27779,N_27866);
nor UO_1730 (O_1730,N_29158,N_28456);
nand UO_1731 (O_1731,N_27554,N_27877);
xnor UO_1732 (O_1732,N_27937,N_28765);
or UO_1733 (O_1733,N_28729,N_27412);
or UO_1734 (O_1734,N_28731,N_28886);
and UO_1735 (O_1735,N_29136,N_28559);
nand UO_1736 (O_1736,N_29230,N_29901);
nor UO_1737 (O_1737,N_29520,N_28626);
nor UO_1738 (O_1738,N_27353,N_29423);
nand UO_1739 (O_1739,N_29615,N_27879);
and UO_1740 (O_1740,N_28505,N_27146);
xor UO_1741 (O_1741,N_28585,N_29194);
or UO_1742 (O_1742,N_29675,N_28118);
nor UO_1743 (O_1743,N_28747,N_27416);
nor UO_1744 (O_1744,N_29226,N_28818);
xor UO_1745 (O_1745,N_28897,N_27375);
or UO_1746 (O_1746,N_27933,N_27690);
xor UO_1747 (O_1747,N_28341,N_29966);
xor UO_1748 (O_1748,N_27399,N_28710);
nor UO_1749 (O_1749,N_28673,N_28435);
or UO_1750 (O_1750,N_28412,N_28597);
nand UO_1751 (O_1751,N_29607,N_27973);
xor UO_1752 (O_1752,N_29966,N_28270);
nor UO_1753 (O_1753,N_28868,N_29528);
or UO_1754 (O_1754,N_28002,N_29627);
and UO_1755 (O_1755,N_27238,N_28340);
and UO_1756 (O_1756,N_27155,N_27616);
nor UO_1757 (O_1757,N_27357,N_29601);
xor UO_1758 (O_1758,N_29019,N_29810);
xor UO_1759 (O_1759,N_29499,N_29946);
nand UO_1760 (O_1760,N_29586,N_27214);
or UO_1761 (O_1761,N_27804,N_29781);
or UO_1762 (O_1762,N_27581,N_27492);
nor UO_1763 (O_1763,N_27466,N_27230);
nand UO_1764 (O_1764,N_29680,N_29243);
nand UO_1765 (O_1765,N_28550,N_27304);
nand UO_1766 (O_1766,N_29904,N_29715);
xnor UO_1767 (O_1767,N_28398,N_27279);
nand UO_1768 (O_1768,N_27203,N_28243);
nor UO_1769 (O_1769,N_29056,N_27223);
xor UO_1770 (O_1770,N_28070,N_29144);
or UO_1771 (O_1771,N_27050,N_29598);
nand UO_1772 (O_1772,N_27742,N_28293);
or UO_1773 (O_1773,N_28097,N_29057);
or UO_1774 (O_1774,N_27492,N_27229);
nand UO_1775 (O_1775,N_29128,N_27431);
nor UO_1776 (O_1776,N_27426,N_28370);
xnor UO_1777 (O_1777,N_29258,N_28821);
and UO_1778 (O_1778,N_29295,N_27253);
or UO_1779 (O_1779,N_28562,N_29844);
xnor UO_1780 (O_1780,N_27399,N_27710);
or UO_1781 (O_1781,N_27933,N_28344);
and UO_1782 (O_1782,N_28848,N_28875);
and UO_1783 (O_1783,N_28215,N_29504);
xor UO_1784 (O_1784,N_28295,N_29635);
xnor UO_1785 (O_1785,N_27952,N_29871);
or UO_1786 (O_1786,N_28814,N_27673);
nand UO_1787 (O_1787,N_29163,N_29421);
and UO_1788 (O_1788,N_29469,N_28487);
and UO_1789 (O_1789,N_29160,N_27060);
nor UO_1790 (O_1790,N_29617,N_29525);
xor UO_1791 (O_1791,N_28066,N_29136);
xor UO_1792 (O_1792,N_27483,N_29141);
nand UO_1793 (O_1793,N_28867,N_28309);
nand UO_1794 (O_1794,N_28885,N_29489);
nor UO_1795 (O_1795,N_27991,N_29943);
nor UO_1796 (O_1796,N_29411,N_27921);
and UO_1797 (O_1797,N_27503,N_27462);
nor UO_1798 (O_1798,N_27446,N_29321);
nand UO_1799 (O_1799,N_28104,N_28555);
xor UO_1800 (O_1800,N_27974,N_29351);
and UO_1801 (O_1801,N_28165,N_28376);
nor UO_1802 (O_1802,N_29383,N_29753);
nor UO_1803 (O_1803,N_27945,N_27815);
nand UO_1804 (O_1804,N_29657,N_28620);
and UO_1805 (O_1805,N_29367,N_29989);
nor UO_1806 (O_1806,N_27837,N_28557);
or UO_1807 (O_1807,N_28274,N_27848);
xnor UO_1808 (O_1808,N_29371,N_27160);
xor UO_1809 (O_1809,N_27432,N_28521);
nor UO_1810 (O_1810,N_28215,N_27516);
and UO_1811 (O_1811,N_29360,N_27485);
or UO_1812 (O_1812,N_27051,N_28872);
xor UO_1813 (O_1813,N_28703,N_29675);
xor UO_1814 (O_1814,N_28598,N_29743);
nand UO_1815 (O_1815,N_28033,N_29538);
or UO_1816 (O_1816,N_27107,N_27620);
nand UO_1817 (O_1817,N_27283,N_28093);
and UO_1818 (O_1818,N_27482,N_27235);
or UO_1819 (O_1819,N_29334,N_28187);
and UO_1820 (O_1820,N_28322,N_28900);
and UO_1821 (O_1821,N_28911,N_29785);
or UO_1822 (O_1822,N_29478,N_28772);
or UO_1823 (O_1823,N_28531,N_27788);
nand UO_1824 (O_1824,N_27353,N_27472);
or UO_1825 (O_1825,N_27539,N_28507);
nand UO_1826 (O_1826,N_28406,N_28739);
nand UO_1827 (O_1827,N_28681,N_28883);
nand UO_1828 (O_1828,N_29756,N_29556);
nor UO_1829 (O_1829,N_27940,N_29723);
nand UO_1830 (O_1830,N_27333,N_27943);
nand UO_1831 (O_1831,N_28416,N_29747);
nor UO_1832 (O_1832,N_27226,N_28135);
nand UO_1833 (O_1833,N_29990,N_28606);
or UO_1834 (O_1834,N_28686,N_27756);
or UO_1835 (O_1835,N_27663,N_28900);
and UO_1836 (O_1836,N_27581,N_27568);
or UO_1837 (O_1837,N_29618,N_27740);
xor UO_1838 (O_1838,N_29275,N_29015);
or UO_1839 (O_1839,N_27924,N_29983);
nor UO_1840 (O_1840,N_27531,N_28586);
nor UO_1841 (O_1841,N_28700,N_29873);
nand UO_1842 (O_1842,N_28853,N_27482);
or UO_1843 (O_1843,N_27881,N_27363);
and UO_1844 (O_1844,N_28020,N_29512);
xor UO_1845 (O_1845,N_28276,N_29973);
xor UO_1846 (O_1846,N_27562,N_27962);
nor UO_1847 (O_1847,N_29625,N_28549);
and UO_1848 (O_1848,N_28950,N_28402);
nor UO_1849 (O_1849,N_29544,N_28001);
and UO_1850 (O_1850,N_29696,N_28824);
xnor UO_1851 (O_1851,N_27263,N_28973);
and UO_1852 (O_1852,N_27845,N_29576);
nor UO_1853 (O_1853,N_28316,N_27903);
nor UO_1854 (O_1854,N_27771,N_27991);
xor UO_1855 (O_1855,N_29829,N_28136);
and UO_1856 (O_1856,N_29510,N_28494);
xor UO_1857 (O_1857,N_29897,N_27792);
and UO_1858 (O_1858,N_29450,N_29330);
and UO_1859 (O_1859,N_27328,N_28631);
or UO_1860 (O_1860,N_29267,N_28225);
xor UO_1861 (O_1861,N_27865,N_29333);
or UO_1862 (O_1862,N_28232,N_28116);
xnor UO_1863 (O_1863,N_27485,N_27229);
xnor UO_1864 (O_1864,N_28208,N_29256);
and UO_1865 (O_1865,N_28985,N_27048);
nand UO_1866 (O_1866,N_28236,N_29632);
xor UO_1867 (O_1867,N_27499,N_29125);
or UO_1868 (O_1868,N_27480,N_28727);
or UO_1869 (O_1869,N_29811,N_29791);
nor UO_1870 (O_1870,N_27958,N_27691);
nand UO_1871 (O_1871,N_27436,N_27931);
and UO_1872 (O_1872,N_27971,N_28516);
xnor UO_1873 (O_1873,N_27259,N_28932);
nand UO_1874 (O_1874,N_27325,N_28362);
nand UO_1875 (O_1875,N_29762,N_28073);
or UO_1876 (O_1876,N_27679,N_27247);
xor UO_1877 (O_1877,N_29798,N_29524);
nor UO_1878 (O_1878,N_29779,N_29941);
and UO_1879 (O_1879,N_28402,N_28646);
or UO_1880 (O_1880,N_27302,N_27931);
nor UO_1881 (O_1881,N_29776,N_28655);
xnor UO_1882 (O_1882,N_29275,N_29162);
xnor UO_1883 (O_1883,N_29354,N_29217);
nor UO_1884 (O_1884,N_28806,N_29119);
nand UO_1885 (O_1885,N_28823,N_27533);
nor UO_1886 (O_1886,N_29155,N_29816);
or UO_1887 (O_1887,N_27215,N_28644);
nor UO_1888 (O_1888,N_29258,N_28985);
nand UO_1889 (O_1889,N_28475,N_28700);
and UO_1890 (O_1890,N_27344,N_29373);
nor UO_1891 (O_1891,N_28050,N_27432);
xor UO_1892 (O_1892,N_28675,N_28881);
and UO_1893 (O_1893,N_29387,N_29843);
or UO_1894 (O_1894,N_29081,N_28442);
xor UO_1895 (O_1895,N_29002,N_27241);
and UO_1896 (O_1896,N_27730,N_27014);
and UO_1897 (O_1897,N_28868,N_27237);
nor UO_1898 (O_1898,N_29424,N_27672);
or UO_1899 (O_1899,N_28188,N_27510);
or UO_1900 (O_1900,N_29105,N_28819);
nor UO_1901 (O_1901,N_29697,N_27694);
and UO_1902 (O_1902,N_27888,N_28973);
nand UO_1903 (O_1903,N_28574,N_28081);
or UO_1904 (O_1904,N_27812,N_29910);
and UO_1905 (O_1905,N_29860,N_27000);
and UO_1906 (O_1906,N_29875,N_29205);
xnor UO_1907 (O_1907,N_29095,N_27424);
nor UO_1908 (O_1908,N_29964,N_29456);
xor UO_1909 (O_1909,N_28519,N_28487);
nor UO_1910 (O_1910,N_28689,N_28162);
nand UO_1911 (O_1911,N_27906,N_29463);
and UO_1912 (O_1912,N_27651,N_29627);
nand UO_1913 (O_1913,N_28924,N_28741);
or UO_1914 (O_1914,N_27060,N_28242);
and UO_1915 (O_1915,N_28766,N_28519);
and UO_1916 (O_1916,N_27739,N_28734);
or UO_1917 (O_1917,N_27853,N_28870);
or UO_1918 (O_1918,N_28078,N_27887);
or UO_1919 (O_1919,N_28201,N_28622);
nor UO_1920 (O_1920,N_29906,N_29755);
nor UO_1921 (O_1921,N_29921,N_28261);
xor UO_1922 (O_1922,N_29097,N_27067);
xnor UO_1923 (O_1923,N_29672,N_28817);
and UO_1924 (O_1924,N_27843,N_28531);
nor UO_1925 (O_1925,N_27635,N_27938);
or UO_1926 (O_1926,N_29912,N_29794);
nor UO_1927 (O_1927,N_29552,N_28093);
xnor UO_1928 (O_1928,N_28612,N_27646);
or UO_1929 (O_1929,N_27145,N_28965);
or UO_1930 (O_1930,N_28679,N_27625);
and UO_1931 (O_1931,N_29689,N_27265);
or UO_1932 (O_1932,N_28811,N_27204);
or UO_1933 (O_1933,N_28461,N_27022);
and UO_1934 (O_1934,N_28692,N_29093);
xnor UO_1935 (O_1935,N_29510,N_27858);
nor UO_1936 (O_1936,N_28897,N_29167);
nand UO_1937 (O_1937,N_27800,N_28968);
or UO_1938 (O_1938,N_29314,N_29879);
nor UO_1939 (O_1939,N_27089,N_29637);
and UO_1940 (O_1940,N_29017,N_28644);
xnor UO_1941 (O_1941,N_29825,N_27567);
and UO_1942 (O_1942,N_27120,N_27373);
and UO_1943 (O_1943,N_29687,N_28951);
xnor UO_1944 (O_1944,N_27696,N_29125);
nand UO_1945 (O_1945,N_27293,N_29910);
or UO_1946 (O_1946,N_28565,N_28525);
nand UO_1947 (O_1947,N_28734,N_27490);
nand UO_1948 (O_1948,N_27226,N_27188);
nand UO_1949 (O_1949,N_29700,N_29729);
nor UO_1950 (O_1950,N_28743,N_28711);
and UO_1951 (O_1951,N_29789,N_27399);
and UO_1952 (O_1952,N_27834,N_28182);
xnor UO_1953 (O_1953,N_29895,N_27239);
or UO_1954 (O_1954,N_29276,N_29638);
xnor UO_1955 (O_1955,N_27722,N_27667);
nand UO_1956 (O_1956,N_27841,N_27876);
and UO_1957 (O_1957,N_27386,N_29435);
xor UO_1958 (O_1958,N_27250,N_27884);
and UO_1959 (O_1959,N_27635,N_28720);
and UO_1960 (O_1960,N_27311,N_28191);
nand UO_1961 (O_1961,N_29830,N_27651);
xnor UO_1962 (O_1962,N_27977,N_27860);
nor UO_1963 (O_1963,N_28560,N_27289);
nor UO_1964 (O_1964,N_28366,N_27961);
and UO_1965 (O_1965,N_27277,N_29669);
and UO_1966 (O_1966,N_27511,N_29873);
nor UO_1967 (O_1967,N_27505,N_27540);
nor UO_1968 (O_1968,N_29752,N_27905);
or UO_1969 (O_1969,N_28059,N_28243);
and UO_1970 (O_1970,N_28980,N_27904);
xnor UO_1971 (O_1971,N_27404,N_27291);
nand UO_1972 (O_1972,N_29879,N_29639);
nand UO_1973 (O_1973,N_27656,N_28457);
or UO_1974 (O_1974,N_28297,N_28356);
xor UO_1975 (O_1975,N_28158,N_28865);
xor UO_1976 (O_1976,N_29320,N_27045);
or UO_1977 (O_1977,N_27129,N_28151);
and UO_1978 (O_1978,N_29723,N_28782);
nor UO_1979 (O_1979,N_29558,N_28024);
and UO_1980 (O_1980,N_29578,N_27396);
xor UO_1981 (O_1981,N_29057,N_27849);
nor UO_1982 (O_1982,N_28483,N_27103);
xor UO_1983 (O_1983,N_28051,N_28426);
and UO_1984 (O_1984,N_29107,N_28680);
nand UO_1985 (O_1985,N_28350,N_28742);
nand UO_1986 (O_1986,N_27930,N_27683);
xor UO_1987 (O_1987,N_29333,N_28747);
nor UO_1988 (O_1988,N_27179,N_28223);
nand UO_1989 (O_1989,N_27294,N_27678);
nand UO_1990 (O_1990,N_28885,N_28963);
or UO_1991 (O_1991,N_27711,N_28004);
or UO_1992 (O_1992,N_29774,N_27617);
or UO_1993 (O_1993,N_28087,N_29728);
nand UO_1994 (O_1994,N_27242,N_29183);
and UO_1995 (O_1995,N_28444,N_27780);
or UO_1996 (O_1996,N_27826,N_28194);
and UO_1997 (O_1997,N_28972,N_27418);
nor UO_1998 (O_1998,N_28283,N_28550);
or UO_1999 (O_1999,N_28347,N_28135);
and UO_2000 (O_2000,N_29331,N_27272);
or UO_2001 (O_2001,N_27062,N_28343);
xor UO_2002 (O_2002,N_27936,N_29093);
or UO_2003 (O_2003,N_27802,N_29145);
xor UO_2004 (O_2004,N_28578,N_29682);
and UO_2005 (O_2005,N_29568,N_28990);
and UO_2006 (O_2006,N_29434,N_28866);
xor UO_2007 (O_2007,N_28058,N_27908);
or UO_2008 (O_2008,N_28789,N_29671);
nor UO_2009 (O_2009,N_29239,N_27957);
nor UO_2010 (O_2010,N_27257,N_27796);
nand UO_2011 (O_2011,N_27088,N_29298);
or UO_2012 (O_2012,N_27590,N_28624);
and UO_2013 (O_2013,N_29169,N_28534);
xnor UO_2014 (O_2014,N_29235,N_28486);
xor UO_2015 (O_2015,N_29210,N_28605);
or UO_2016 (O_2016,N_27936,N_29983);
xnor UO_2017 (O_2017,N_28234,N_29665);
nand UO_2018 (O_2018,N_28265,N_29531);
and UO_2019 (O_2019,N_29614,N_28318);
and UO_2020 (O_2020,N_27518,N_29995);
and UO_2021 (O_2021,N_27217,N_28797);
nor UO_2022 (O_2022,N_27960,N_28341);
or UO_2023 (O_2023,N_29532,N_28840);
or UO_2024 (O_2024,N_27719,N_27357);
nand UO_2025 (O_2025,N_28858,N_28799);
nor UO_2026 (O_2026,N_28416,N_29880);
and UO_2027 (O_2027,N_28530,N_29236);
nor UO_2028 (O_2028,N_27068,N_28094);
nand UO_2029 (O_2029,N_27856,N_27694);
or UO_2030 (O_2030,N_27702,N_27984);
nand UO_2031 (O_2031,N_28749,N_29052);
nand UO_2032 (O_2032,N_28584,N_29802);
nand UO_2033 (O_2033,N_27504,N_29311);
and UO_2034 (O_2034,N_27209,N_27390);
xnor UO_2035 (O_2035,N_28481,N_27330);
xor UO_2036 (O_2036,N_28045,N_27160);
xnor UO_2037 (O_2037,N_28455,N_29704);
nor UO_2038 (O_2038,N_27515,N_28154);
xor UO_2039 (O_2039,N_27227,N_27985);
or UO_2040 (O_2040,N_28228,N_29558);
nor UO_2041 (O_2041,N_28941,N_29911);
nor UO_2042 (O_2042,N_28464,N_29871);
xnor UO_2043 (O_2043,N_27161,N_29414);
and UO_2044 (O_2044,N_28889,N_28101);
and UO_2045 (O_2045,N_27610,N_29297);
nor UO_2046 (O_2046,N_27923,N_28413);
nor UO_2047 (O_2047,N_29616,N_27374);
or UO_2048 (O_2048,N_29613,N_27455);
or UO_2049 (O_2049,N_27917,N_29571);
nand UO_2050 (O_2050,N_28408,N_29225);
xor UO_2051 (O_2051,N_28654,N_29475);
nor UO_2052 (O_2052,N_29618,N_27721);
nand UO_2053 (O_2053,N_29973,N_27547);
nand UO_2054 (O_2054,N_28477,N_28886);
nor UO_2055 (O_2055,N_27050,N_28169);
nor UO_2056 (O_2056,N_29749,N_29255);
or UO_2057 (O_2057,N_27494,N_29013);
nand UO_2058 (O_2058,N_28089,N_27070);
xor UO_2059 (O_2059,N_29851,N_28712);
nand UO_2060 (O_2060,N_29259,N_29419);
or UO_2061 (O_2061,N_29734,N_28042);
nor UO_2062 (O_2062,N_29271,N_27093);
nor UO_2063 (O_2063,N_28141,N_29447);
and UO_2064 (O_2064,N_27763,N_28218);
or UO_2065 (O_2065,N_27130,N_29117);
and UO_2066 (O_2066,N_29790,N_28824);
nor UO_2067 (O_2067,N_27353,N_29491);
xor UO_2068 (O_2068,N_27960,N_28140);
nand UO_2069 (O_2069,N_29117,N_29647);
or UO_2070 (O_2070,N_29756,N_29776);
nor UO_2071 (O_2071,N_27952,N_28465);
nor UO_2072 (O_2072,N_29806,N_27936);
and UO_2073 (O_2073,N_29837,N_29030);
nand UO_2074 (O_2074,N_28230,N_27826);
or UO_2075 (O_2075,N_28967,N_27971);
nand UO_2076 (O_2076,N_28791,N_28276);
and UO_2077 (O_2077,N_29316,N_29745);
and UO_2078 (O_2078,N_28918,N_27095);
or UO_2079 (O_2079,N_28633,N_28018);
nor UO_2080 (O_2080,N_29925,N_27854);
xnor UO_2081 (O_2081,N_28485,N_28227);
nand UO_2082 (O_2082,N_28699,N_29443);
or UO_2083 (O_2083,N_27481,N_28703);
nand UO_2084 (O_2084,N_28417,N_27984);
and UO_2085 (O_2085,N_29315,N_29328);
xor UO_2086 (O_2086,N_29667,N_29256);
xnor UO_2087 (O_2087,N_27779,N_29026);
nand UO_2088 (O_2088,N_29401,N_28675);
nand UO_2089 (O_2089,N_28820,N_29918);
or UO_2090 (O_2090,N_27768,N_29782);
or UO_2091 (O_2091,N_29869,N_27259);
nor UO_2092 (O_2092,N_27483,N_28217);
xor UO_2093 (O_2093,N_27821,N_28816);
nor UO_2094 (O_2094,N_28272,N_28668);
nand UO_2095 (O_2095,N_27199,N_28353);
nor UO_2096 (O_2096,N_28347,N_29543);
and UO_2097 (O_2097,N_29092,N_29799);
xnor UO_2098 (O_2098,N_28684,N_29805);
or UO_2099 (O_2099,N_27822,N_28712);
and UO_2100 (O_2100,N_28359,N_28940);
nand UO_2101 (O_2101,N_28909,N_27521);
nand UO_2102 (O_2102,N_27522,N_28314);
or UO_2103 (O_2103,N_28706,N_27100);
or UO_2104 (O_2104,N_28058,N_28755);
and UO_2105 (O_2105,N_27778,N_28575);
nand UO_2106 (O_2106,N_27760,N_27963);
and UO_2107 (O_2107,N_29605,N_28863);
nor UO_2108 (O_2108,N_28560,N_27270);
nand UO_2109 (O_2109,N_27812,N_28615);
and UO_2110 (O_2110,N_27330,N_27486);
xnor UO_2111 (O_2111,N_28625,N_28459);
nor UO_2112 (O_2112,N_28133,N_28158);
or UO_2113 (O_2113,N_28626,N_29361);
and UO_2114 (O_2114,N_28482,N_29839);
xor UO_2115 (O_2115,N_28944,N_28470);
nor UO_2116 (O_2116,N_27118,N_27571);
or UO_2117 (O_2117,N_28948,N_27655);
nand UO_2118 (O_2118,N_27897,N_27481);
xnor UO_2119 (O_2119,N_28239,N_28134);
xnor UO_2120 (O_2120,N_28486,N_29503);
and UO_2121 (O_2121,N_27093,N_27356);
xor UO_2122 (O_2122,N_28496,N_28767);
or UO_2123 (O_2123,N_27211,N_29104);
and UO_2124 (O_2124,N_28782,N_29882);
nand UO_2125 (O_2125,N_27289,N_27573);
nand UO_2126 (O_2126,N_27062,N_28077);
xnor UO_2127 (O_2127,N_27143,N_29718);
xor UO_2128 (O_2128,N_28627,N_29244);
xnor UO_2129 (O_2129,N_28057,N_28737);
nand UO_2130 (O_2130,N_27531,N_28216);
nor UO_2131 (O_2131,N_28398,N_29745);
nor UO_2132 (O_2132,N_29840,N_27411);
and UO_2133 (O_2133,N_27040,N_27525);
or UO_2134 (O_2134,N_28083,N_29913);
nor UO_2135 (O_2135,N_27837,N_28989);
nor UO_2136 (O_2136,N_29307,N_29659);
xor UO_2137 (O_2137,N_28203,N_29435);
nand UO_2138 (O_2138,N_29183,N_29656);
nand UO_2139 (O_2139,N_29924,N_28758);
and UO_2140 (O_2140,N_28171,N_27434);
nand UO_2141 (O_2141,N_28965,N_27311);
nor UO_2142 (O_2142,N_29344,N_29591);
nor UO_2143 (O_2143,N_29702,N_27069);
or UO_2144 (O_2144,N_27635,N_28628);
and UO_2145 (O_2145,N_29395,N_29364);
xor UO_2146 (O_2146,N_27203,N_29738);
or UO_2147 (O_2147,N_29284,N_27084);
or UO_2148 (O_2148,N_28766,N_28177);
nand UO_2149 (O_2149,N_27447,N_27057);
xor UO_2150 (O_2150,N_29427,N_28779);
nor UO_2151 (O_2151,N_28778,N_27699);
nor UO_2152 (O_2152,N_28992,N_29908);
and UO_2153 (O_2153,N_29283,N_29802);
nor UO_2154 (O_2154,N_29854,N_29245);
and UO_2155 (O_2155,N_28956,N_27470);
xor UO_2156 (O_2156,N_29153,N_27058);
and UO_2157 (O_2157,N_28255,N_29076);
and UO_2158 (O_2158,N_29077,N_27253);
xor UO_2159 (O_2159,N_27829,N_29241);
and UO_2160 (O_2160,N_28911,N_27042);
nand UO_2161 (O_2161,N_28003,N_29920);
nand UO_2162 (O_2162,N_27123,N_28946);
and UO_2163 (O_2163,N_28129,N_28480);
or UO_2164 (O_2164,N_28409,N_29827);
xor UO_2165 (O_2165,N_27746,N_29550);
or UO_2166 (O_2166,N_29891,N_28905);
nor UO_2167 (O_2167,N_29713,N_29735);
nand UO_2168 (O_2168,N_28175,N_27092);
xnor UO_2169 (O_2169,N_27849,N_27810);
nand UO_2170 (O_2170,N_27044,N_29016);
or UO_2171 (O_2171,N_27322,N_29687);
and UO_2172 (O_2172,N_28988,N_29627);
xnor UO_2173 (O_2173,N_28065,N_29749);
nand UO_2174 (O_2174,N_28832,N_29876);
xnor UO_2175 (O_2175,N_27560,N_27313);
nand UO_2176 (O_2176,N_28895,N_28593);
or UO_2177 (O_2177,N_27461,N_29971);
nor UO_2178 (O_2178,N_28243,N_27574);
xnor UO_2179 (O_2179,N_27631,N_27874);
nand UO_2180 (O_2180,N_27933,N_29902);
nand UO_2181 (O_2181,N_29555,N_29081);
and UO_2182 (O_2182,N_29787,N_28894);
and UO_2183 (O_2183,N_27063,N_28813);
or UO_2184 (O_2184,N_27393,N_28002);
nand UO_2185 (O_2185,N_27477,N_27671);
and UO_2186 (O_2186,N_29749,N_28754);
nand UO_2187 (O_2187,N_28203,N_29781);
or UO_2188 (O_2188,N_28862,N_29471);
xnor UO_2189 (O_2189,N_28716,N_28841);
nand UO_2190 (O_2190,N_28635,N_29767);
and UO_2191 (O_2191,N_29147,N_29585);
xor UO_2192 (O_2192,N_28669,N_28747);
xor UO_2193 (O_2193,N_29781,N_27436);
and UO_2194 (O_2194,N_29569,N_28022);
nor UO_2195 (O_2195,N_27297,N_27187);
nor UO_2196 (O_2196,N_27829,N_29676);
and UO_2197 (O_2197,N_28078,N_29715);
or UO_2198 (O_2198,N_27009,N_28987);
nor UO_2199 (O_2199,N_28820,N_27174);
or UO_2200 (O_2200,N_29173,N_27821);
nand UO_2201 (O_2201,N_29359,N_28620);
nand UO_2202 (O_2202,N_28421,N_27974);
or UO_2203 (O_2203,N_29872,N_28827);
or UO_2204 (O_2204,N_28222,N_29334);
nor UO_2205 (O_2205,N_28233,N_29969);
or UO_2206 (O_2206,N_27539,N_27147);
nor UO_2207 (O_2207,N_28585,N_28935);
nor UO_2208 (O_2208,N_29145,N_29984);
nand UO_2209 (O_2209,N_28665,N_29760);
nand UO_2210 (O_2210,N_29738,N_27933);
xnor UO_2211 (O_2211,N_28316,N_29804);
or UO_2212 (O_2212,N_27281,N_29743);
or UO_2213 (O_2213,N_29187,N_28057);
xor UO_2214 (O_2214,N_27189,N_28498);
xnor UO_2215 (O_2215,N_28141,N_27193);
nor UO_2216 (O_2216,N_29002,N_29028);
or UO_2217 (O_2217,N_28868,N_28865);
and UO_2218 (O_2218,N_29845,N_27690);
nor UO_2219 (O_2219,N_27558,N_28577);
nand UO_2220 (O_2220,N_28388,N_29677);
nand UO_2221 (O_2221,N_28936,N_27711);
xnor UO_2222 (O_2222,N_27149,N_29505);
nor UO_2223 (O_2223,N_27182,N_28094);
nand UO_2224 (O_2224,N_29946,N_29298);
or UO_2225 (O_2225,N_29803,N_28368);
or UO_2226 (O_2226,N_29041,N_29997);
xor UO_2227 (O_2227,N_29083,N_29708);
or UO_2228 (O_2228,N_27390,N_28851);
nor UO_2229 (O_2229,N_27955,N_27008);
and UO_2230 (O_2230,N_28638,N_29321);
nand UO_2231 (O_2231,N_28344,N_29148);
xnor UO_2232 (O_2232,N_27553,N_28214);
xnor UO_2233 (O_2233,N_29004,N_27998);
or UO_2234 (O_2234,N_29524,N_28033);
or UO_2235 (O_2235,N_28258,N_27985);
nor UO_2236 (O_2236,N_27399,N_28218);
nand UO_2237 (O_2237,N_27584,N_28751);
nand UO_2238 (O_2238,N_28584,N_27838);
nor UO_2239 (O_2239,N_28322,N_28524);
xor UO_2240 (O_2240,N_29310,N_29100);
xor UO_2241 (O_2241,N_27166,N_28707);
and UO_2242 (O_2242,N_28848,N_28425);
or UO_2243 (O_2243,N_29691,N_29220);
or UO_2244 (O_2244,N_28786,N_27174);
xor UO_2245 (O_2245,N_28999,N_27550);
and UO_2246 (O_2246,N_27067,N_28243);
and UO_2247 (O_2247,N_28759,N_28636);
nand UO_2248 (O_2248,N_27442,N_29890);
nor UO_2249 (O_2249,N_28490,N_27254);
nor UO_2250 (O_2250,N_27247,N_27578);
nand UO_2251 (O_2251,N_29131,N_27263);
xor UO_2252 (O_2252,N_28773,N_27101);
and UO_2253 (O_2253,N_27561,N_28507);
xnor UO_2254 (O_2254,N_27250,N_28444);
xor UO_2255 (O_2255,N_28388,N_28371);
nor UO_2256 (O_2256,N_27051,N_27287);
nor UO_2257 (O_2257,N_27045,N_29039);
nor UO_2258 (O_2258,N_27144,N_29723);
nor UO_2259 (O_2259,N_28258,N_27978);
or UO_2260 (O_2260,N_29310,N_28344);
nand UO_2261 (O_2261,N_28009,N_28650);
nor UO_2262 (O_2262,N_28824,N_28781);
nand UO_2263 (O_2263,N_29852,N_27874);
or UO_2264 (O_2264,N_29197,N_27686);
nand UO_2265 (O_2265,N_29234,N_28729);
xnor UO_2266 (O_2266,N_28152,N_28166);
nor UO_2267 (O_2267,N_28674,N_29929);
nand UO_2268 (O_2268,N_27168,N_27584);
xnor UO_2269 (O_2269,N_29594,N_27786);
nand UO_2270 (O_2270,N_28293,N_27447);
and UO_2271 (O_2271,N_29139,N_28030);
nor UO_2272 (O_2272,N_28744,N_28862);
nor UO_2273 (O_2273,N_28167,N_29368);
nor UO_2274 (O_2274,N_28755,N_29426);
nand UO_2275 (O_2275,N_27344,N_28161);
nor UO_2276 (O_2276,N_27662,N_28064);
xnor UO_2277 (O_2277,N_29916,N_27041);
and UO_2278 (O_2278,N_27028,N_27865);
and UO_2279 (O_2279,N_27839,N_27868);
nor UO_2280 (O_2280,N_27838,N_29388);
nor UO_2281 (O_2281,N_28497,N_27194);
or UO_2282 (O_2282,N_27498,N_29872);
or UO_2283 (O_2283,N_27863,N_29369);
xnor UO_2284 (O_2284,N_27401,N_27148);
and UO_2285 (O_2285,N_27676,N_28590);
xnor UO_2286 (O_2286,N_28649,N_28364);
and UO_2287 (O_2287,N_29916,N_27931);
or UO_2288 (O_2288,N_28421,N_28875);
or UO_2289 (O_2289,N_27640,N_28557);
or UO_2290 (O_2290,N_29472,N_28354);
nor UO_2291 (O_2291,N_28615,N_28887);
or UO_2292 (O_2292,N_29953,N_27584);
nor UO_2293 (O_2293,N_28189,N_27218);
nand UO_2294 (O_2294,N_29724,N_27587);
nand UO_2295 (O_2295,N_29691,N_27163);
nand UO_2296 (O_2296,N_27597,N_28405);
xnor UO_2297 (O_2297,N_28568,N_28840);
nand UO_2298 (O_2298,N_29461,N_28303);
xnor UO_2299 (O_2299,N_27636,N_28749);
and UO_2300 (O_2300,N_28243,N_28657);
or UO_2301 (O_2301,N_27204,N_27181);
nor UO_2302 (O_2302,N_27235,N_27232);
nor UO_2303 (O_2303,N_29007,N_27328);
and UO_2304 (O_2304,N_28666,N_28676);
or UO_2305 (O_2305,N_29102,N_29221);
and UO_2306 (O_2306,N_28400,N_27288);
or UO_2307 (O_2307,N_27304,N_27432);
xnor UO_2308 (O_2308,N_27280,N_27269);
nor UO_2309 (O_2309,N_28211,N_28094);
nor UO_2310 (O_2310,N_27158,N_29801);
or UO_2311 (O_2311,N_28714,N_29362);
nor UO_2312 (O_2312,N_27972,N_28504);
nor UO_2313 (O_2313,N_28987,N_27731);
or UO_2314 (O_2314,N_28216,N_28700);
nor UO_2315 (O_2315,N_29407,N_27411);
nor UO_2316 (O_2316,N_29669,N_28106);
nor UO_2317 (O_2317,N_27385,N_29629);
xnor UO_2318 (O_2318,N_28047,N_27986);
or UO_2319 (O_2319,N_27910,N_27604);
nor UO_2320 (O_2320,N_28554,N_29559);
or UO_2321 (O_2321,N_28063,N_28502);
and UO_2322 (O_2322,N_27032,N_28953);
nand UO_2323 (O_2323,N_28793,N_29099);
xor UO_2324 (O_2324,N_27532,N_29501);
nor UO_2325 (O_2325,N_28136,N_27637);
nand UO_2326 (O_2326,N_29088,N_28765);
nand UO_2327 (O_2327,N_27278,N_29657);
nor UO_2328 (O_2328,N_27787,N_27149);
or UO_2329 (O_2329,N_29869,N_29881);
nand UO_2330 (O_2330,N_27680,N_28316);
nand UO_2331 (O_2331,N_27997,N_28480);
xnor UO_2332 (O_2332,N_27163,N_28231);
nand UO_2333 (O_2333,N_27996,N_28425);
or UO_2334 (O_2334,N_29331,N_28839);
nor UO_2335 (O_2335,N_28891,N_28086);
and UO_2336 (O_2336,N_28915,N_29060);
or UO_2337 (O_2337,N_27813,N_29929);
nand UO_2338 (O_2338,N_28320,N_28099);
and UO_2339 (O_2339,N_27325,N_28417);
xnor UO_2340 (O_2340,N_29132,N_29999);
and UO_2341 (O_2341,N_28694,N_28567);
and UO_2342 (O_2342,N_27966,N_28691);
and UO_2343 (O_2343,N_27109,N_29842);
and UO_2344 (O_2344,N_28975,N_28101);
nor UO_2345 (O_2345,N_28327,N_27819);
nor UO_2346 (O_2346,N_28356,N_28491);
nand UO_2347 (O_2347,N_27111,N_29785);
and UO_2348 (O_2348,N_29022,N_29480);
and UO_2349 (O_2349,N_27080,N_27561);
xor UO_2350 (O_2350,N_28438,N_29340);
nor UO_2351 (O_2351,N_28025,N_29129);
and UO_2352 (O_2352,N_27381,N_29969);
xnor UO_2353 (O_2353,N_27751,N_27367);
nor UO_2354 (O_2354,N_28266,N_29688);
or UO_2355 (O_2355,N_28048,N_28925);
xor UO_2356 (O_2356,N_28553,N_29128);
and UO_2357 (O_2357,N_27878,N_28755);
or UO_2358 (O_2358,N_29767,N_28931);
nor UO_2359 (O_2359,N_27801,N_27041);
xor UO_2360 (O_2360,N_28136,N_27793);
xnor UO_2361 (O_2361,N_27389,N_27234);
xor UO_2362 (O_2362,N_29968,N_28892);
nand UO_2363 (O_2363,N_27788,N_27839);
and UO_2364 (O_2364,N_27373,N_29522);
xor UO_2365 (O_2365,N_29895,N_27133);
nand UO_2366 (O_2366,N_27178,N_27905);
xor UO_2367 (O_2367,N_28345,N_27209);
and UO_2368 (O_2368,N_28621,N_28077);
and UO_2369 (O_2369,N_27495,N_28332);
xor UO_2370 (O_2370,N_29099,N_29902);
nor UO_2371 (O_2371,N_29706,N_29191);
nor UO_2372 (O_2372,N_27199,N_29185);
xnor UO_2373 (O_2373,N_28339,N_28447);
xnor UO_2374 (O_2374,N_27824,N_27647);
and UO_2375 (O_2375,N_28629,N_27789);
nand UO_2376 (O_2376,N_28529,N_28823);
and UO_2377 (O_2377,N_29574,N_28227);
and UO_2378 (O_2378,N_28232,N_29759);
nand UO_2379 (O_2379,N_29252,N_27123);
xor UO_2380 (O_2380,N_28685,N_28168);
or UO_2381 (O_2381,N_27071,N_29119);
or UO_2382 (O_2382,N_29158,N_28138);
nor UO_2383 (O_2383,N_28430,N_27899);
nor UO_2384 (O_2384,N_27097,N_29650);
and UO_2385 (O_2385,N_28030,N_27705);
nand UO_2386 (O_2386,N_29323,N_27710);
or UO_2387 (O_2387,N_27210,N_28939);
nand UO_2388 (O_2388,N_28386,N_29788);
nand UO_2389 (O_2389,N_28555,N_27081);
xnor UO_2390 (O_2390,N_28919,N_27731);
and UO_2391 (O_2391,N_29576,N_27980);
nand UO_2392 (O_2392,N_29967,N_27135);
nand UO_2393 (O_2393,N_27866,N_27484);
and UO_2394 (O_2394,N_28039,N_27401);
or UO_2395 (O_2395,N_27294,N_27004);
nor UO_2396 (O_2396,N_28796,N_27597);
nor UO_2397 (O_2397,N_29359,N_28926);
xnor UO_2398 (O_2398,N_29196,N_27233);
xor UO_2399 (O_2399,N_28999,N_28214);
xnor UO_2400 (O_2400,N_29137,N_29752);
nor UO_2401 (O_2401,N_27783,N_28726);
nand UO_2402 (O_2402,N_28626,N_29340);
nor UO_2403 (O_2403,N_27404,N_29426);
xnor UO_2404 (O_2404,N_29310,N_28522);
nand UO_2405 (O_2405,N_28913,N_29188);
xnor UO_2406 (O_2406,N_27068,N_29688);
nor UO_2407 (O_2407,N_29081,N_29931);
or UO_2408 (O_2408,N_28763,N_29344);
or UO_2409 (O_2409,N_27739,N_28206);
nor UO_2410 (O_2410,N_28483,N_27441);
nand UO_2411 (O_2411,N_28380,N_27459);
nand UO_2412 (O_2412,N_27342,N_27232);
nor UO_2413 (O_2413,N_28218,N_28638);
nor UO_2414 (O_2414,N_28365,N_28090);
xor UO_2415 (O_2415,N_27205,N_29547);
nor UO_2416 (O_2416,N_29282,N_27226);
xor UO_2417 (O_2417,N_28797,N_28897);
xor UO_2418 (O_2418,N_28888,N_27026);
nand UO_2419 (O_2419,N_27818,N_29755);
nor UO_2420 (O_2420,N_27626,N_28942);
or UO_2421 (O_2421,N_28835,N_28269);
or UO_2422 (O_2422,N_29675,N_27071);
and UO_2423 (O_2423,N_28965,N_28578);
or UO_2424 (O_2424,N_27095,N_27313);
xor UO_2425 (O_2425,N_27898,N_28165);
xor UO_2426 (O_2426,N_28313,N_28644);
xor UO_2427 (O_2427,N_27410,N_28630);
nor UO_2428 (O_2428,N_28747,N_29590);
or UO_2429 (O_2429,N_27710,N_28045);
or UO_2430 (O_2430,N_28657,N_27223);
xnor UO_2431 (O_2431,N_28092,N_27859);
or UO_2432 (O_2432,N_29336,N_28334);
or UO_2433 (O_2433,N_29600,N_29068);
xor UO_2434 (O_2434,N_29615,N_28005);
xor UO_2435 (O_2435,N_28539,N_29194);
nor UO_2436 (O_2436,N_28381,N_27410);
and UO_2437 (O_2437,N_27328,N_27098);
nor UO_2438 (O_2438,N_27101,N_28796);
nand UO_2439 (O_2439,N_27312,N_29767);
xor UO_2440 (O_2440,N_27617,N_27466);
and UO_2441 (O_2441,N_27778,N_27591);
nor UO_2442 (O_2442,N_27409,N_28549);
nor UO_2443 (O_2443,N_27849,N_27180);
and UO_2444 (O_2444,N_27754,N_27145);
nand UO_2445 (O_2445,N_28284,N_29219);
or UO_2446 (O_2446,N_27279,N_28505);
or UO_2447 (O_2447,N_27657,N_29380);
nor UO_2448 (O_2448,N_29071,N_28889);
and UO_2449 (O_2449,N_28938,N_28099);
or UO_2450 (O_2450,N_28452,N_27081);
or UO_2451 (O_2451,N_29280,N_29986);
or UO_2452 (O_2452,N_28283,N_29223);
nor UO_2453 (O_2453,N_28788,N_28569);
and UO_2454 (O_2454,N_28424,N_28219);
xor UO_2455 (O_2455,N_27803,N_27008);
and UO_2456 (O_2456,N_29017,N_27318);
xor UO_2457 (O_2457,N_27189,N_29269);
or UO_2458 (O_2458,N_27094,N_29434);
nand UO_2459 (O_2459,N_27062,N_27182);
or UO_2460 (O_2460,N_27620,N_28851);
and UO_2461 (O_2461,N_28379,N_29087);
nor UO_2462 (O_2462,N_29931,N_29254);
nor UO_2463 (O_2463,N_28166,N_28027);
xor UO_2464 (O_2464,N_29948,N_29052);
and UO_2465 (O_2465,N_29713,N_27460);
and UO_2466 (O_2466,N_29327,N_27932);
xor UO_2467 (O_2467,N_27928,N_28073);
nand UO_2468 (O_2468,N_29093,N_29939);
xnor UO_2469 (O_2469,N_28625,N_28346);
or UO_2470 (O_2470,N_29968,N_29024);
nor UO_2471 (O_2471,N_27076,N_28344);
and UO_2472 (O_2472,N_27308,N_28473);
nor UO_2473 (O_2473,N_27216,N_27983);
or UO_2474 (O_2474,N_29369,N_27385);
xor UO_2475 (O_2475,N_27310,N_27123);
nor UO_2476 (O_2476,N_29103,N_28561);
xnor UO_2477 (O_2477,N_28772,N_28988);
xor UO_2478 (O_2478,N_27969,N_29885);
nor UO_2479 (O_2479,N_28014,N_27190);
nor UO_2480 (O_2480,N_29580,N_28333);
nor UO_2481 (O_2481,N_27764,N_29714);
and UO_2482 (O_2482,N_27390,N_29562);
nor UO_2483 (O_2483,N_28652,N_27080);
or UO_2484 (O_2484,N_29835,N_29135);
nor UO_2485 (O_2485,N_29131,N_28361);
nor UO_2486 (O_2486,N_27718,N_27090);
nor UO_2487 (O_2487,N_28520,N_27028);
nand UO_2488 (O_2488,N_29109,N_27446);
nor UO_2489 (O_2489,N_28932,N_29931);
xor UO_2490 (O_2490,N_29893,N_28139);
nand UO_2491 (O_2491,N_28937,N_29593);
and UO_2492 (O_2492,N_27581,N_28815);
or UO_2493 (O_2493,N_27577,N_28773);
xor UO_2494 (O_2494,N_28825,N_27128);
and UO_2495 (O_2495,N_29403,N_28027);
or UO_2496 (O_2496,N_28950,N_28899);
xnor UO_2497 (O_2497,N_28225,N_27916);
nor UO_2498 (O_2498,N_29909,N_28132);
or UO_2499 (O_2499,N_28905,N_28214);
xor UO_2500 (O_2500,N_27115,N_29875);
nor UO_2501 (O_2501,N_28486,N_28541);
xor UO_2502 (O_2502,N_28781,N_27973);
nor UO_2503 (O_2503,N_29711,N_29071);
nand UO_2504 (O_2504,N_27447,N_27140);
nor UO_2505 (O_2505,N_27543,N_28416);
and UO_2506 (O_2506,N_27639,N_28145);
or UO_2507 (O_2507,N_28063,N_27747);
nand UO_2508 (O_2508,N_29727,N_28325);
xnor UO_2509 (O_2509,N_27518,N_27250);
xnor UO_2510 (O_2510,N_28535,N_28632);
nand UO_2511 (O_2511,N_28838,N_28327);
nand UO_2512 (O_2512,N_28429,N_29041);
nor UO_2513 (O_2513,N_29359,N_27178);
xor UO_2514 (O_2514,N_27578,N_27963);
nor UO_2515 (O_2515,N_27501,N_27328);
and UO_2516 (O_2516,N_28576,N_27715);
xnor UO_2517 (O_2517,N_27346,N_27588);
or UO_2518 (O_2518,N_27281,N_27259);
and UO_2519 (O_2519,N_29991,N_27192);
and UO_2520 (O_2520,N_29548,N_28869);
or UO_2521 (O_2521,N_29035,N_29654);
nor UO_2522 (O_2522,N_28183,N_28466);
and UO_2523 (O_2523,N_29024,N_27329);
or UO_2524 (O_2524,N_29192,N_27338);
or UO_2525 (O_2525,N_27849,N_28741);
xor UO_2526 (O_2526,N_29344,N_27820);
and UO_2527 (O_2527,N_29409,N_27889);
or UO_2528 (O_2528,N_28585,N_27803);
or UO_2529 (O_2529,N_28072,N_29951);
or UO_2530 (O_2530,N_27648,N_28407);
or UO_2531 (O_2531,N_29929,N_27101);
nor UO_2532 (O_2532,N_29899,N_29208);
or UO_2533 (O_2533,N_27557,N_27263);
nand UO_2534 (O_2534,N_27942,N_28768);
or UO_2535 (O_2535,N_27961,N_27471);
and UO_2536 (O_2536,N_28869,N_28165);
or UO_2537 (O_2537,N_29146,N_28141);
nand UO_2538 (O_2538,N_27376,N_28076);
nand UO_2539 (O_2539,N_28877,N_27803);
xor UO_2540 (O_2540,N_27924,N_28554);
or UO_2541 (O_2541,N_27651,N_27849);
nor UO_2542 (O_2542,N_28594,N_27353);
or UO_2543 (O_2543,N_27383,N_29732);
nor UO_2544 (O_2544,N_29619,N_29211);
nor UO_2545 (O_2545,N_28922,N_28775);
nor UO_2546 (O_2546,N_29698,N_29310);
or UO_2547 (O_2547,N_27795,N_27583);
or UO_2548 (O_2548,N_29159,N_28777);
and UO_2549 (O_2549,N_27814,N_28737);
and UO_2550 (O_2550,N_28022,N_29130);
nor UO_2551 (O_2551,N_27465,N_28158);
xor UO_2552 (O_2552,N_28606,N_27200);
nand UO_2553 (O_2553,N_29978,N_29049);
nor UO_2554 (O_2554,N_27740,N_29465);
nand UO_2555 (O_2555,N_28161,N_29420);
xor UO_2556 (O_2556,N_29441,N_28635);
nor UO_2557 (O_2557,N_28744,N_29964);
nor UO_2558 (O_2558,N_29293,N_27058);
nor UO_2559 (O_2559,N_28606,N_27992);
nand UO_2560 (O_2560,N_27856,N_29786);
nand UO_2561 (O_2561,N_28312,N_27217);
nand UO_2562 (O_2562,N_28124,N_29156);
xor UO_2563 (O_2563,N_29251,N_29206);
and UO_2564 (O_2564,N_29679,N_29139);
nand UO_2565 (O_2565,N_27480,N_29088);
nor UO_2566 (O_2566,N_28482,N_29265);
and UO_2567 (O_2567,N_29600,N_28489);
xnor UO_2568 (O_2568,N_28271,N_27009);
or UO_2569 (O_2569,N_27813,N_28399);
or UO_2570 (O_2570,N_28205,N_27563);
nor UO_2571 (O_2571,N_27718,N_27007);
nor UO_2572 (O_2572,N_29890,N_28150);
xnor UO_2573 (O_2573,N_27576,N_29736);
or UO_2574 (O_2574,N_28247,N_27542);
nor UO_2575 (O_2575,N_28414,N_27784);
xor UO_2576 (O_2576,N_28848,N_27075);
nor UO_2577 (O_2577,N_29804,N_27132);
nand UO_2578 (O_2578,N_27984,N_27871);
or UO_2579 (O_2579,N_27202,N_27776);
or UO_2580 (O_2580,N_27952,N_28651);
and UO_2581 (O_2581,N_27054,N_29036);
nand UO_2582 (O_2582,N_29879,N_28822);
nor UO_2583 (O_2583,N_27677,N_29457);
nand UO_2584 (O_2584,N_29752,N_28151);
or UO_2585 (O_2585,N_27079,N_29444);
or UO_2586 (O_2586,N_28096,N_29489);
xnor UO_2587 (O_2587,N_27735,N_29189);
nand UO_2588 (O_2588,N_29526,N_28908);
or UO_2589 (O_2589,N_28567,N_29732);
xor UO_2590 (O_2590,N_27214,N_27553);
or UO_2591 (O_2591,N_29232,N_27936);
nand UO_2592 (O_2592,N_29522,N_29314);
xnor UO_2593 (O_2593,N_29188,N_28055);
nand UO_2594 (O_2594,N_29741,N_27440);
xor UO_2595 (O_2595,N_28117,N_27868);
or UO_2596 (O_2596,N_29287,N_29586);
or UO_2597 (O_2597,N_27404,N_28036);
nor UO_2598 (O_2598,N_28870,N_29566);
and UO_2599 (O_2599,N_27116,N_27345);
and UO_2600 (O_2600,N_29575,N_28059);
and UO_2601 (O_2601,N_28012,N_28669);
nor UO_2602 (O_2602,N_28197,N_27450);
and UO_2603 (O_2603,N_29707,N_28592);
or UO_2604 (O_2604,N_27723,N_28818);
nor UO_2605 (O_2605,N_28045,N_28851);
and UO_2606 (O_2606,N_28207,N_29730);
nor UO_2607 (O_2607,N_28961,N_29354);
and UO_2608 (O_2608,N_28494,N_29281);
xnor UO_2609 (O_2609,N_27692,N_29435);
xnor UO_2610 (O_2610,N_29179,N_28042);
nand UO_2611 (O_2611,N_29614,N_27505);
or UO_2612 (O_2612,N_27524,N_29978);
xor UO_2613 (O_2613,N_29658,N_29362);
and UO_2614 (O_2614,N_27713,N_29586);
nor UO_2615 (O_2615,N_29748,N_27365);
xor UO_2616 (O_2616,N_28626,N_27420);
nor UO_2617 (O_2617,N_28487,N_27574);
xor UO_2618 (O_2618,N_29979,N_29753);
nand UO_2619 (O_2619,N_29087,N_29546);
and UO_2620 (O_2620,N_27036,N_27975);
xnor UO_2621 (O_2621,N_28149,N_27106);
nor UO_2622 (O_2622,N_28554,N_29662);
and UO_2623 (O_2623,N_29431,N_28176);
or UO_2624 (O_2624,N_28139,N_28871);
and UO_2625 (O_2625,N_27116,N_29718);
nand UO_2626 (O_2626,N_29862,N_29371);
or UO_2627 (O_2627,N_27817,N_29724);
xnor UO_2628 (O_2628,N_29949,N_27218);
xnor UO_2629 (O_2629,N_28777,N_28646);
or UO_2630 (O_2630,N_29451,N_28224);
nand UO_2631 (O_2631,N_27653,N_29532);
and UO_2632 (O_2632,N_27878,N_29529);
nor UO_2633 (O_2633,N_29094,N_29129);
and UO_2634 (O_2634,N_27524,N_27367);
xor UO_2635 (O_2635,N_27493,N_28598);
xnor UO_2636 (O_2636,N_28459,N_28982);
and UO_2637 (O_2637,N_28340,N_29429);
nor UO_2638 (O_2638,N_29545,N_28703);
xnor UO_2639 (O_2639,N_28110,N_28897);
nor UO_2640 (O_2640,N_28045,N_28282);
or UO_2641 (O_2641,N_29323,N_29735);
nor UO_2642 (O_2642,N_29108,N_29605);
and UO_2643 (O_2643,N_29014,N_29987);
and UO_2644 (O_2644,N_28863,N_29839);
xor UO_2645 (O_2645,N_27529,N_28415);
xnor UO_2646 (O_2646,N_28736,N_27653);
nand UO_2647 (O_2647,N_28534,N_28863);
and UO_2648 (O_2648,N_29013,N_29098);
or UO_2649 (O_2649,N_27223,N_29063);
nand UO_2650 (O_2650,N_27270,N_28708);
or UO_2651 (O_2651,N_27697,N_27150);
nand UO_2652 (O_2652,N_29757,N_27586);
nand UO_2653 (O_2653,N_29161,N_28611);
xnor UO_2654 (O_2654,N_28953,N_27297);
and UO_2655 (O_2655,N_29662,N_28704);
nor UO_2656 (O_2656,N_28354,N_28039);
and UO_2657 (O_2657,N_27087,N_29724);
nor UO_2658 (O_2658,N_29078,N_27852);
or UO_2659 (O_2659,N_29506,N_28399);
nor UO_2660 (O_2660,N_28523,N_28735);
xor UO_2661 (O_2661,N_29845,N_28948);
and UO_2662 (O_2662,N_27655,N_29489);
nand UO_2663 (O_2663,N_29972,N_29356);
nor UO_2664 (O_2664,N_27334,N_27586);
or UO_2665 (O_2665,N_27350,N_28014);
or UO_2666 (O_2666,N_27033,N_29640);
xor UO_2667 (O_2667,N_28259,N_27049);
nand UO_2668 (O_2668,N_29073,N_29060);
nor UO_2669 (O_2669,N_29163,N_29833);
xnor UO_2670 (O_2670,N_29416,N_29509);
and UO_2671 (O_2671,N_29925,N_29965);
or UO_2672 (O_2672,N_29244,N_29824);
or UO_2673 (O_2673,N_28927,N_28255);
or UO_2674 (O_2674,N_27692,N_28804);
nand UO_2675 (O_2675,N_29297,N_28213);
nand UO_2676 (O_2676,N_28792,N_28883);
nor UO_2677 (O_2677,N_29436,N_28236);
nor UO_2678 (O_2678,N_27864,N_28647);
or UO_2679 (O_2679,N_29021,N_27818);
or UO_2680 (O_2680,N_27413,N_29394);
and UO_2681 (O_2681,N_27107,N_27427);
nor UO_2682 (O_2682,N_28515,N_27596);
nor UO_2683 (O_2683,N_27847,N_27355);
and UO_2684 (O_2684,N_27604,N_27289);
nand UO_2685 (O_2685,N_28316,N_28897);
or UO_2686 (O_2686,N_28755,N_28334);
nand UO_2687 (O_2687,N_29531,N_29586);
nor UO_2688 (O_2688,N_28097,N_29887);
and UO_2689 (O_2689,N_28917,N_27467);
nand UO_2690 (O_2690,N_29259,N_28915);
or UO_2691 (O_2691,N_28493,N_29053);
or UO_2692 (O_2692,N_28814,N_28862);
and UO_2693 (O_2693,N_28011,N_28741);
nor UO_2694 (O_2694,N_27313,N_29954);
and UO_2695 (O_2695,N_27190,N_27443);
nand UO_2696 (O_2696,N_29639,N_28220);
xnor UO_2697 (O_2697,N_27935,N_28229);
nand UO_2698 (O_2698,N_28090,N_29952);
nor UO_2699 (O_2699,N_29958,N_28401);
xor UO_2700 (O_2700,N_29570,N_28487);
and UO_2701 (O_2701,N_27517,N_27981);
nand UO_2702 (O_2702,N_29425,N_29388);
nor UO_2703 (O_2703,N_29595,N_28306);
xnor UO_2704 (O_2704,N_28387,N_29918);
nand UO_2705 (O_2705,N_27223,N_29958);
or UO_2706 (O_2706,N_27928,N_27613);
nor UO_2707 (O_2707,N_27568,N_29100);
and UO_2708 (O_2708,N_27253,N_27654);
or UO_2709 (O_2709,N_29643,N_27425);
and UO_2710 (O_2710,N_27608,N_28213);
and UO_2711 (O_2711,N_28759,N_29368);
nor UO_2712 (O_2712,N_28937,N_28239);
nand UO_2713 (O_2713,N_27831,N_27811);
nor UO_2714 (O_2714,N_29865,N_29489);
nor UO_2715 (O_2715,N_29957,N_27744);
or UO_2716 (O_2716,N_29456,N_29207);
nand UO_2717 (O_2717,N_27046,N_28938);
nand UO_2718 (O_2718,N_29970,N_28171);
and UO_2719 (O_2719,N_27091,N_28250);
xnor UO_2720 (O_2720,N_27033,N_28792);
and UO_2721 (O_2721,N_29106,N_29704);
xor UO_2722 (O_2722,N_28447,N_27447);
nor UO_2723 (O_2723,N_29106,N_28139);
nor UO_2724 (O_2724,N_29130,N_27049);
nand UO_2725 (O_2725,N_27409,N_27902);
and UO_2726 (O_2726,N_27317,N_29388);
or UO_2727 (O_2727,N_27127,N_28877);
and UO_2728 (O_2728,N_28299,N_28233);
and UO_2729 (O_2729,N_29663,N_28983);
nor UO_2730 (O_2730,N_28783,N_27103);
nand UO_2731 (O_2731,N_27473,N_28956);
nand UO_2732 (O_2732,N_27974,N_29986);
nand UO_2733 (O_2733,N_27968,N_27907);
or UO_2734 (O_2734,N_27825,N_28584);
or UO_2735 (O_2735,N_27084,N_27389);
nand UO_2736 (O_2736,N_27723,N_27233);
or UO_2737 (O_2737,N_29312,N_29107);
xor UO_2738 (O_2738,N_27546,N_29392);
or UO_2739 (O_2739,N_28264,N_29601);
nor UO_2740 (O_2740,N_27905,N_27646);
nand UO_2741 (O_2741,N_28613,N_28887);
nor UO_2742 (O_2742,N_28731,N_29761);
nand UO_2743 (O_2743,N_27014,N_29984);
nor UO_2744 (O_2744,N_28355,N_29810);
xnor UO_2745 (O_2745,N_28348,N_28141);
xor UO_2746 (O_2746,N_27668,N_28343);
nand UO_2747 (O_2747,N_29770,N_27722);
nor UO_2748 (O_2748,N_28126,N_28946);
nand UO_2749 (O_2749,N_27599,N_27736);
nand UO_2750 (O_2750,N_29593,N_28409);
or UO_2751 (O_2751,N_27673,N_27111);
xor UO_2752 (O_2752,N_29077,N_29054);
and UO_2753 (O_2753,N_27808,N_29665);
nor UO_2754 (O_2754,N_28496,N_28356);
nor UO_2755 (O_2755,N_28915,N_28432);
and UO_2756 (O_2756,N_27778,N_28939);
and UO_2757 (O_2757,N_28044,N_29417);
xnor UO_2758 (O_2758,N_28941,N_28120);
and UO_2759 (O_2759,N_27936,N_27265);
and UO_2760 (O_2760,N_29924,N_27630);
nor UO_2761 (O_2761,N_27888,N_27905);
and UO_2762 (O_2762,N_28263,N_29197);
nand UO_2763 (O_2763,N_29825,N_29650);
or UO_2764 (O_2764,N_28213,N_27662);
and UO_2765 (O_2765,N_27073,N_27959);
nor UO_2766 (O_2766,N_28471,N_27424);
and UO_2767 (O_2767,N_28364,N_27963);
xnor UO_2768 (O_2768,N_28031,N_28162);
and UO_2769 (O_2769,N_28830,N_29498);
or UO_2770 (O_2770,N_27331,N_28100);
nor UO_2771 (O_2771,N_28296,N_28115);
xor UO_2772 (O_2772,N_29288,N_28580);
xnor UO_2773 (O_2773,N_28882,N_28838);
nor UO_2774 (O_2774,N_27491,N_29549);
and UO_2775 (O_2775,N_29980,N_27589);
xor UO_2776 (O_2776,N_29114,N_28731);
nor UO_2777 (O_2777,N_27220,N_28288);
and UO_2778 (O_2778,N_27871,N_29594);
nor UO_2779 (O_2779,N_29310,N_29472);
nand UO_2780 (O_2780,N_27505,N_29003);
nor UO_2781 (O_2781,N_28662,N_28059);
nand UO_2782 (O_2782,N_27280,N_28990);
nand UO_2783 (O_2783,N_29398,N_29625);
or UO_2784 (O_2784,N_29059,N_27695);
nand UO_2785 (O_2785,N_29334,N_27012);
xnor UO_2786 (O_2786,N_27315,N_27216);
and UO_2787 (O_2787,N_28698,N_27816);
nand UO_2788 (O_2788,N_27864,N_27965);
nand UO_2789 (O_2789,N_29596,N_29786);
and UO_2790 (O_2790,N_27709,N_27994);
nand UO_2791 (O_2791,N_29351,N_29290);
nor UO_2792 (O_2792,N_27802,N_28470);
and UO_2793 (O_2793,N_27069,N_29776);
nor UO_2794 (O_2794,N_28313,N_29420);
nand UO_2795 (O_2795,N_28220,N_29070);
or UO_2796 (O_2796,N_27789,N_28685);
and UO_2797 (O_2797,N_28808,N_29560);
nand UO_2798 (O_2798,N_27880,N_28149);
xor UO_2799 (O_2799,N_27658,N_29594);
or UO_2800 (O_2800,N_28010,N_27748);
nor UO_2801 (O_2801,N_29967,N_28701);
and UO_2802 (O_2802,N_28110,N_29409);
nand UO_2803 (O_2803,N_28406,N_29042);
nand UO_2804 (O_2804,N_27654,N_28786);
nand UO_2805 (O_2805,N_27515,N_27465);
nand UO_2806 (O_2806,N_27877,N_28045);
or UO_2807 (O_2807,N_28316,N_29361);
and UO_2808 (O_2808,N_27346,N_27697);
nor UO_2809 (O_2809,N_27435,N_28379);
xor UO_2810 (O_2810,N_27314,N_28341);
nand UO_2811 (O_2811,N_29328,N_27536);
nand UO_2812 (O_2812,N_28287,N_27257);
and UO_2813 (O_2813,N_28251,N_29776);
nand UO_2814 (O_2814,N_28757,N_29684);
and UO_2815 (O_2815,N_28726,N_28376);
nand UO_2816 (O_2816,N_27067,N_29906);
or UO_2817 (O_2817,N_29403,N_28151);
nand UO_2818 (O_2818,N_27105,N_27757);
or UO_2819 (O_2819,N_28025,N_27938);
or UO_2820 (O_2820,N_28654,N_28476);
and UO_2821 (O_2821,N_29247,N_29157);
nand UO_2822 (O_2822,N_29566,N_29964);
or UO_2823 (O_2823,N_27065,N_28489);
or UO_2824 (O_2824,N_28040,N_28808);
xnor UO_2825 (O_2825,N_29049,N_29931);
nor UO_2826 (O_2826,N_27359,N_29186);
xnor UO_2827 (O_2827,N_28233,N_27571);
nand UO_2828 (O_2828,N_29035,N_29398);
nand UO_2829 (O_2829,N_27192,N_27218);
and UO_2830 (O_2830,N_27569,N_28370);
or UO_2831 (O_2831,N_28625,N_29134);
or UO_2832 (O_2832,N_27130,N_27537);
nand UO_2833 (O_2833,N_27367,N_29121);
and UO_2834 (O_2834,N_29883,N_28904);
nor UO_2835 (O_2835,N_27875,N_29462);
or UO_2836 (O_2836,N_29857,N_27518);
and UO_2837 (O_2837,N_27156,N_28942);
or UO_2838 (O_2838,N_27561,N_28043);
and UO_2839 (O_2839,N_29805,N_28673);
xor UO_2840 (O_2840,N_28111,N_29502);
nand UO_2841 (O_2841,N_27106,N_28558);
xnor UO_2842 (O_2842,N_27972,N_29219);
nand UO_2843 (O_2843,N_28502,N_28772);
and UO_2844 (O_2844,N_28989,N_28197);
and UO_2845 (O_2845,N_29175,N_28582);
and UO_2846 (O_2846,N_29805,N_29651);
or UO_2847 (O_2847,N_29928,N_27382);
or UO_2848 (O_2848,N_28776,N_27938);
nor UO_2849 (O_2849,N_28404,N_28549);
nor UO_2850 (O_2850,N_29271,N_27057);
nor UO_2851 (O_2851,N_28750,N_29022);
or UO_2852 (O_2852,N_29708,N_29909);
nand UO_2853 (O_2853,N_29060,N_28359);
nor UO_2854 (O_2854,N_28860,N_29067);
or UO_2855 (O_2855,N_27917,N_27891);
and UO_2856 (O_2856,N_27853,N_29598);
nor UO_2857 (O_2857,N_27244,N_27793);
nor UO_2858 (O_2858,N_29271,N_27834);
and UO_2859 (O_2859,N_28760,N_28272);
and UO_2860 (O_2860,N_29673,N_27174);
or UO_2861 (O_2861,N_27406,N_29534);
nor UO_2862 (O_2862,N_29948,N_28590);
nor UO_2863 (O_2863,N_27097,N_29058);
xnor UO_2864 (O_2864,N_27159,N_27947);
and UO_2865 (O_2865,N_28767,N_29493);
and UO_2866 (O_2866,N_28798,N_28745);
nand UO_2867 (O_2867,N_28252,N_28680);
or UO_2868 (O_2868,N_28835,N_27753);
xor UO_2869 (O_2869,N_27200,N_28030);
or UO_2870 (O_2870,N_28850,N_27832);
or UO_2871 (O_2871,N_29930,N_27234);
or UO_2872 (O_2872,N_27375,N_27022);
or UO_2873 (O_2873,N_29082,N_29067);
xnor UO_2874 (O_2874,N_28534,N_27203);
xnor UO_2875 (O_2875,N_27068,N_27350);
or UO_2876 (O_2876,N_28108,N_28417);
xnor UO_2877 (O_2877,N_29492,N_28015);
and UO_2878 (O_2878,N_29969,N_29821);
and UO_2879 (O_2879,N_29646,N_29891);
nor UO_2880 (O_2880,N_28897,N_27282);
nand UO_2881 (O_2881,N_27625,N_27483);
xor UO_2882 (O_2882,N_29782,N_29172);
nand UO_2883 (O_2883,N_29335,N_27538);
nand UO_2884 (O_2884,N_28198,N_27946);
nor UO_2885 (O_2885,N_29711,N_28288);
nand UO_2886 (O_2886,N_28663,N_29449);
or UO_2887 (O_2887,N_28580,N_29610);
xor UO_2888 (O_2888,N_28172,N_29467);
nor UO_2889 (O_2889,N_28721,N_29562);
xnor UO_2890 (O_2890,N_29784,N_29841);
or UO_2891 (O_2891,N_27709,N_29380);
or UO_2892 (O_2892,N_29313,N_28797);
nand UO_2893 (O_2893,N_27228,N_29292);
and UO_2894 (O_2894,N_28150,N_27597);
and UO_2895 (O_2895,N_29562,N_29833);
nand UO_2896 (O_2896,N_28673,N_27177);
nand UO_2897 (O_2897,N_28384,N_28178);
or UO_2898 (O_2898,N_27119,N_27890);
nand UO_2899 (O_2899,N_29850,N_27218);
and UO_2900 (O_2900,N_29899,N_28094);
or UO_2901 (O_2901,N_28993,N_29558);
nand UO_2902 (O_2902,N_28708,N_27387);
xor UO_2903 (O_2903,N_27645,N_27387);
and UO_2904 (O_2904,N_27040,N_28257);
and UO_2905 (O_2905,N_28877,N_27040);
nor UO_2906 (O_2906,N_27960,N_29598);
xor UO_2907 (O_2907,N_29219,N_29218);
nor UO_2908 (O_2908,N_27079,N_27165);
or UO_2909 (O_2909,N_29157,N_29621);
nor UO_2910 (O_2910,N_29267,N_29406);
nor UO_2911 (O_2911,N_27703,N_28240);
nor UO_2912 (O_2912,N_28044,N_29199);
nand UO_2913 (O_2913,N_27576,N_27283);
nand UO_2914 (O_2914,N_27513,N_29537);
and UO_2915 (O_2915,N_28772,N_29397);
nor UO_2916 (O_2916,N_27000,N_28162);
and UO_2917 (O_2917,N_27107,N_28989);
nand UO_2918 (O_2918,N_29903,N_28008);
nor UO_2919 (O_2919,N_27740,N_27386);
nor UO_2920 (O_2920,N_29117,N_29568);
nand UO_2921 (O_2921,N_28199,N_29184);
and UO_2922 (O_2922,N_29233,N_29004);
nand UO_2923 (O_2923,N_28765,N_28617);
xor UO_2924 (O_2924,N_29648,N_28835);
nand UO_2925 (O_2925,N_29300,N_29896);
nand UO_2926 (O_2926,N_28725,N_29342);
nand UO_2927 (O_2927,N_29038,N_28074);
xnor UO_2928 (O_2928,N_27409,N_29951);
and UO_2929 (O_2929,N_28419,N_29459);
and UO_2930 (O_2930,N_28228,N_28983);
or UO_2931 (O_2931,N_27463,N_27704);
or UO_2932 (O_2932,N_29567,N_27914);
and UO_2933 (O_2933,N_27148,N_29247);
and UO_2934 (O_2934,N_29133,N_29286);
or UO_2935 (O_2935,N_28945,N_27134);
or UO_2936 (O_2936,N_28944,N_28584);
xor UO_2937 (O_2937,N_28500,N_27261);
and UO_2938 (O_2938,N_27250,N_29829);
xor UO_2939 (O_2939,N_27389,N_29659);
and UO_2940 (O_2940,N_29794,N_27121);
xor UO_2941 (O_2941,N_28171,N_27435);
xor UO_2942 (O_2942,N_27155,N_29897);
xor UO_2943 (O_2943,N_29123,N_27117);
xnor UO_2944 (O_2944,N_27345,N_27275);
or UO_2945 (O_2945,N_28310,N_28666);
or UO_2946 (O_2946,N_28829,N_28741);
nand UO_2947 (O_2947,N_29301,N_27487);
xor UO_2948 (O_2948,N_28844,N_29550);
nand UO_2949 (O_2949,N_29102,N_27377);
xor UO_2950 (O_2950,N_28682,N_29765);
nor UO_2951 (O_2951,N_29387,N_27906);
or UO_2952 (O_2952,N_28249,N_27483);
or UO_2953 (O_2953,N_28161,N_27164);
nor UO_2954 (O_2954,N_29094,N_28478);
nand UO_2955 (O_2955,N_28574,N_28759);
and UO_2956 (O_2956,N_27371,N_28490);
xnor UO_2957 (O_2957,N_28284,N_28780);
nor UO_2958 (O_2958,N_28493,N_29525);
xnor UO_2959 (O_2959,N_27657,N_29506);
or UO_2960 (O_2960,N_29399,N_29935);
xnor UO_2961 (O_2961,N_29687,N_29092);
and UO_2962 (O_2962,N_27942,N_29902);
or UO_2963 (O_2963,N_27054,N_28911);
and UO_2964 (O_2964,N_29097,N_28772);
xor UO_2965 (O_2965,N_27256,N_27682);
or UO_2966 (O_2966,N_27421,N_29272);
nand UO_2967 (O_2967,N_27557,N_28719);
and UO_2968 (O_2968,N_28066,N_27188);
nand UO_2969 (O_2969,N_29010,N_28023);
or UO_2970 (O_2970,N_29852,N_28307);
xnor UO_2971 (O_2971,N_27255,N_28372);
xor UO_2972 (O_2972,N_27882,N_29629);
nor UO_2973 (O_2973,N_27120,N_27251);
nand UO_2974 (O_2974,N_27885,N_28349);
or UO_2975 (O_2975,N_27988,N_27790);
nor UO_2976 (O_2976,N_28442,N_29349);
or UO_2977 (O_2977,N_29683,N_27743);
or UO_2978 (O_2978,N_28021,N_27857);
and UO_2979 (O_2979,N_27515,N_27496);
nor UO_2980 (O_2980,N_29977,N_27942);
xor UO_2981 (O_2981,N_28748,N_27815);
and UO_2982 (O_2982,N_28638,N_27770);
nor UO_2983 (O_2983,N_28473,N_28018);
nor UO_2984 (O_2984,N_28207,N_28770);
nor UO_2985 (O_2985,N_28692,N_29172);
nor UO_2986 (O_2986,N_29004,N_29447);
nand UO_2987 (O_2987,N_27132,N_29272);
nor UO_2988 (O_2988,N_28634,N_29272);
and UO_2989 (O_2989,N_27591,N_29612);
xnor UO_2990 (O_2990,N_28156,N_28888);
or UO_2991 (O_2991,N_28164,N_29763);
nand UO_2992 (O_2992,N_29195,N_27529);
nand UO_2993 (O_2993,N_28362,N_27002);
nand UO_2994 (O_2994,N_29329,N_27506);
xor UO_2995 (O_2995,N_29544,N_28171);
and UO_2996 (O_2996,N_29949,N_28507);
and UO_2997 (O_2997,N_29787,N_29713);
nor UO_2998 (O_2998,N_28286,N_29822);
nand UO_2999 (O_2999,N_29170,N_27035);
or UO_3000 (O_3000,N_29385,N_28349);
nand UO_3001 (O_3001,N_28595,N_29517);
xnor UO_3002 (O_3002,N_29938,N_29440);
or UO_3003 (O_3003,N_28935,N_27706);
xnor UO_3004 (O_3004,N_27170,N_28853);
nor UO_3005 (O_3005,N_27226,N_28418);
and UO_3006 (O_3006,N_28386,N_29588);
nand UO_3007 (O_3007,N_27097,N_29008);
nor UO_3008 (O_3008,N_28538,N_29340);
nand UO_3009 (O_3009,N_27188,N_29213);
xnor UO_3010 (O_3010,N_27327,N_28577);
xor UO_3011 (O_3011,N_27919,N_29996);
xor UO_3012 (O_3012,N_27007,N_28546);
or UO_3013 (O_3013,N_28782,N_29179);
xnor UO_3014 (O_3014,N_28254,N_27996);
nand UO_3015 (O_3015,N_27136,N_29261);
xnor UO_3016 (O_3016,N_27694,N_29618);
xor UO_3017 (O_3017,N_28075,N_29764);
xnor UO_3018 (O_3018,N_29230,N_28452);
or UO_3019 (O_3019,N_28984,N_28496);
nand UO_3020 (O_3020,N_27130,N_29021);
nand UO_3021 (O_3021,N_29574,N_27971);
xnor UO_3022 (O_3022,N_28197,N_28613);
nand UO_3023 (O_3023,N_29090,N_29007);
nor UO_3024 (O_3024,N_28590,N_28784);
and UO_3025 (O_3025,N_28087,N_27120);
nand UO_3026 (O_3026,N_29559,N_28615);
or UO_3027 (O_3027,N_29865,N_29627);
nand UO_3028 (O_3028,N_29650,N_28906);
nor UO_3029 (O_3029,N_27975,N_29405);
nand UO_3030 (O_3030,N_29218,N_29901);
and UO_3031 (O_3031,N_29014,N_28202);
xnor UO_3032 (O_3032,N_27316,N_27249);
and UO_3033 (O_3033,N_28921,N_27915);
nand UO_3034 (O_3034,N_29706,N_27460);
nor UO_3035 (O_3035,N_29518,N_29730);
and UO_3036 (O_3036,N_28113,N_28152);
xor UO_3037 (O_3037,N_27726,N_28827);
and UO_3038 (O_3038,N_29920,N_27559);
and UO_3039 (O_3039,N_29789,N_27647);
or UO_3040 (O_3040,N_27909,N_27764);
and UO_3041 (O_3041,N_29387,N_29227);
and UO_3042 (O_3042,N_27761,N_28619);
xnor UO_3043 (O_3043,N_27867,N_27396);
nor UO_3044 (O_3044,N_27485,N_27008);
xor UO_3045 (O_3045,N_29158,N_27716);
nand UO_3046 (O_3046,N_29632,N_29227);
nor UO_3047 (O_3047,N_27043,N_28590);
nand UO_3048 (O_3048,N_29346,N_28514);
nor UO_3049 (O_3049,N_29633,N_29547);
xnor UO_3050 (O_3050,N_28905,N_28290);
or UO_3051 (O_3051,N_29707,N_29849);
and UO_3052 (O_3052,N_28356,N_29618);
xnor UO_3053 (O_3053,N_27430,N_29668);
nand UO_3054 (O_3054,N_28784,N_27351);
xor UO_3055 (O_3055,N_27385,N_28530);
or UO_3056 (O_3056,N_28524,N_27223);
nand UO_3057 (O_3057,N_29556,N_28661);
or UO_3058 (O_3058,N_28066,N_29225);
nor UO_3059 (O_3059,N_27276,N_29467);
and UO_3060 (O_3060,N_29430,N_27434);
and UO_3061 (O_3061,N_28219,N_28738);
nor UO_3062 (O_3062,N_29302,N_29101);
or UO_3063 (O_3063,N_29614,N_27386);
and UO_3064 (O_3064,N_28536,N_29584);
xor UO_3065 (O_3065,N_28538,N_27517);
nor UO_3066 (O_3066,N_28883,N_28444);
xor UO_3067 (O_3067,N_28810,N_27012);
nor UO_3068 (O_3068,N_29584,N_29425);
and UO_3069 (O_3069,N_29169,N_27815);
nand UO_3070 (O_3070,N_29029,N_27754);
xnor UO_3071 (O_3071,N_29144,N_27535);
or UO_3072 (O_3072,N_28921,N_27949);
and UO_3073 (O_3073,N_28049,N_27870);
and UO_3074 (O_3074,N_29689,N_27833);
or UO_3075 (O_3075,N_28492,N_28052);
and UO_3076 (O_3076,N_29489,N_29858);
nand UO_3077 (O_3077,N_27628,N_27005);
nand UO_3078 (O_3078,N_29890,N_27379);
or UO_3079 (O_3079,N_28164,N_29276);
and UO_3080 (O_3080,N_28367,N_27199);
or UO_3081 (O_3081,N_27436,N_29873);
xor UO_3082 (O_3082,N_28159,N_27692);
or UO_3083 (O_3083,N_27826,N_27132);
and UO_3084 (O_3084,N_28835,N_27291);
nor UO_3085 (O_3085,N_28490,N_27946);
or UO_3086 (O_3086,N_27499,N_28669);
xor UO_3087 (O_3087,N_28569,N_29057);
nor UO_3088 (O_3088,N_27769,N_29475);
xor UO_3089 (O_3089,N_27503,N_27529);
or UO_3090 (O_3090,N_28822,N_27454);
xnor UO_3091 (O_3091,N_29079,N_28308);
nor UO_3092 (O_3092,N_27117,N_29129);
and UO_3093 (O_3093,N_29930,N_27607);
nor UO_3094 (O_3094,N_27165,N_28165);
nor UO_3095 (O_3095,N_29918,N_28428);
xnor UO_3096 (O_3096,N_28913,N_27492);
and UO_3097 (O_3097,N_29756,N_29353);
xnor UO_3098 (O_3098,N_28031,N_27239);
nor UO_3099 (O_3099,N_27561,N_29577);
or UO_3100 (O_3100,N_29778,N_29056);
xor UO_3101 (O_3101,N_27356,N_28343);
nand UO_3102 (O_3102,N_29702,N_29921);
nand UO_3103 (O_3103,N_29694,N_29692);
nor UO_3104 (O_3104,N_28232,N_29359);
xnor UO_3105 (O_3105,N_28751,N_28019);
nor UO_3106 (O_3106,N_28567,N_29541);
and UO_3107 (O_3107,N_27441,N_28095);
and UO_3108 (O_3108,N_28211,N_28778);
and UO_3109 (O_3109,N_28661,N_29033);
and UO_3110 (O_3110,N_29494,N_28133);
nand UO_3111 (O_3111,N_28306,N_29391);
nand UO_3112 (O_3112,N_28607,N_29019);
and UO_3113 (O_3113,N_27563,N_28265);
or UO_3114 (O_3114,N_28867,N_29601);
nor UO_3115 (O_3115,N_27784,N_28667);
nor UO_3116 (O_3116,N_29222,N_27994);
xor UO_3117 (O_3117,N_28116,N_27466);
and UO_3118 (O_3118,N_27142,N_27776);
nand UO_3119 (O_3119,N_29213,N_28769);
and UO_3120 (O_3120,N_27964,N_28019);
or UO_3121 (O_3121,N_28264,N_29093);
and UO_3122 (O_3122,N_28675,N_27533);
nand UO_3123 (O_3123,N_27919,N_28318);
xnor UO_3124 (O_3124,N_29867,N_29729);
nor UO_3125 (O_3125,N_28257,N_29111);
xnor UO_3126 (O_3126,N_28356,N_27451);
nand UO_3127 (O_3127,N_29132,N_28086);
or UO_3128 (O_3128,N_29535,N_28766);
xnor UO_3129 (O_3129,N_29431,N_29948);
xor UO_3130 (O_3130,N_27569,N_29533);
nand UO_3131 (O_3131,N_28869,N_27500);
or UO_3132 (O_3132,N_28304,N_28307);
nand UO_3133 (O_3133,N_29718,N_28933);
or UO_3134 (O_3134,N_28632,N_27507);
nand UO_3135 (O_3135,N_27889,N_28331);
nand UO_3136 (O_3136,N_27660,N_29094);
nor UO_3137 (O_3137,N_29019,N_29671);
nand UO_3138 (O_3138,N_27393,N_28438);
nand UO_3139 (O_3139,N_27299,N_29450);
nor UO_3140 (O_3140,N_29476,N_28722);
and UO_3141 (O_3141,N_29932,N_29681);
xnor UO_3142 (O_3142,N_27797,N_27530);
xor UO_3143 (O_3143,N_27690,N_29769);
nand UO_3144 (O_3144,N_29077,N_29395);
xor UO_3145 (O_3145,N_27320,N_27614);
nor UO_3146 (O_3146,N_27200,N_27380);
or UO_3147 (O_3147,N_27789,N_29905);
or UO_3148 (O_3148,N_27265,N_29734);
and UO_3149 (O_3149,N_29047,N_28832);
nand UO_3150 (O_3150,N_28424,N_28189);
nor UO_3151 (O_3151,N_28173,N_28380);
nor UO_3152 (O_3152,N_28486,N_29497);
xor UO_3153 (O_3153,N_28213,N_27261);
or UO_3154 (O_3154,N_29111,N_27215);
xnor UO_3155 (O_3155,N_28307,N_27355);
or UO_3156 (O_3156,N_28222,N_28287);
xor UO_3157 (O_3157,N_27140,N_27625);
nand UO_3158 (O_3158,N_28402,N_29591);
xnor UO_3159 (O_3159,N_29262,N_27331);
or UO_3160 (O_3160,N_27335,N_28924);
and UO_3161 (O_3161,N_29909,N_29058);
nand UO_3162 (O_3162,N_27956,N_28581);
nand UO_3163 (O_3163,N_29082,N_27036);
xor UO_3164 (O_3164,N_29385,N_27392);
or UO_3165 (O_3165,N_27231,N_29563);
and UO_3166 (O_3166,N_29071,N_27545);
xor UO_3167 (O_3167,N_29246,N_27379);
nor UO_3168 (O_3168,N_28658,N_27266);
xor UO_3169 (O_3169,N_27515,N_28613);
xnor UO_3170 (O_3170,N_29423,N_29919);
xor UO_3171 (O_3171,N_29821,N_27970);
xor UO_3172 (O_3172,N_28953,N_27781);
and UO_3173 (O_3173,N_28819,N_27227);
nor UO_3174 (O_3174,N_29998,N_29256);
xnor UO_3175 (O_3175,N_29671,N_28546);
and UO_3176 (O_3176,N_29873,N_29520);
nor UO_3177 (O_3177,N_27895,N_28788);
and UO_3178 (O_3178,N_28811,N_27612);
nor UO_3179 (O_3179,N_29144,N_29635);
and UO_3180 (O_3180,N_29337,N_28936);
xnor UO_3181 (O_3181,N_27012,N_28684);
and UO_3182 (O_3182,N_27278,N_28870);
or UO_3183 (O_3183,N_27711,N_28109);
nand UO_3184 (O_3184,N_27180,N_29964);
or UO_3185 (O_3185,N_28919,N_29272);
xor UO_3186 (O_3186,N_28607,N_27973);
nor UO_3187 (O_3187,N_29951,N_29475);
and UO_3188 (O_3188,N_28142,N_29059);
nand UO_3189 (O_3189,N_29330,N_28251);
or UO_3190 (O_3190,N_28579,N_28761);
or UO_3191 (O_3191,N_27094,N_28607);
nand UO_3192 (O_3192,N_29241,N_27879);
and UO_3193 (O_3193,N_27207,N_27842);
or UO_3194 (O_3194,N_27725,N_28335);
and UO_3195 (O_3195,N_29564,N_28079);
nand UO_3196 (O_3196,N_27720,N_29743);
nor UO_3197 (O_3197,N_28697,N_29489);
nand UO_3198 (O_3198,N_28562,N_28941);
nor UO_3199 (O_3199,N_28244,N_27443);
or UO_3200 (O_3200,N_27823,N_27973);
or UO_3201 (O_3201,N_28709,N_27720);
nand UO_3202 (O_3202,N_28830,N_27888);
nor UO_3203 (O_3203,N_28185,N_29468);
or UO_3204 (O_3204,N_29049,N_29915);
or UO_3205 (O_3205,N_28827,N_28198);
or UO_3206 (O_3206,N_29074,N_28350);
and UO_3207 (O_3207,N_29198,N_28120);
and UO_3208 (O_3208,N_29925,N_29185);
nand UO_3209 (O_3209,N_28387,N_29260);
and UO_3210 (O_3210,N_28798,N_29283);
nand UO_3211 (O_3211,N_29180,N_27112);
xnor UO_3212 (O_3212,N_29318,N_28793);
nor UO_3213 (O_3213,N_28884,N_27577);
and UO_3214 (O_3214,N_28013,N_27893);
and UO_3215 (O_3215,N_28874,N_27553);
and UO_3216 (O_3216,N_29282,N_27987);
and UO_3217 (O_3217,N_28665,N_29395);
nand UO_3218 (O_3218,N_28939,N_27018);
and UO_3219 (O_3219,N_29056,N_29063);
nor UO_3220 (O_3220,N_29802,N_29208);
xor UO_3221 (O_3221,N_29397,N_29139);
or UO_3222 (O_3222,N_27651,N_27205);
nor UO_3223 (O_3223,N_29167,N_27960);
nor UO_3224 (O_3224,N_28972,N_29941);
nor UO_3225 (O_3225,N_27504,N_28368);
and UO_3226 (O_3226,N_28560,N_27253);
nand UO_3227 (O_3227,N_29041,N_28025);
nand UO_3228 (O_3228,N_28679,N_29488);
or UO_3229 (O_3229,N_27496,N_27285);
and UO_3230 (O_3230,N_27770,N_28358);
and UO_3231 (O_3231,N_29929,N_27042);
and UO_3232 (O_3232,N_28820,N_29178);
and UO_3233 (O_3233,N_27843,N_29884);
nor UO_3234 (O_3234,N_29977,N_27785);
xnor UO_3235 (O_3235,N_28572,N_28849);
nor UO_3236 (O_3236,N_29898,N_29920);
and UO_3237 (O_3237,N_27530,N_27925);
nor UO_3238 (O_3238,N_27297,N_27753);
xor UO_3239 (O_3239,N_27520,N_29640);
nor UO_3240 (O_3240,N_29011,N_27637);
or UO_3241 (O_3241,N_27194,N_27401);
and UO_3242 (O_3242,N_27721,N_28113);
xnor UO_3243 (O_3243,N_27980,N_28636);
nor UO_3244 (O_3244,N_28545,N_29440);
nor UO_3245 (O_3245,N_28077,N_27274);
and UO_3246 (O_3246,N_29091,N_28112);
or UO_3247 (O_3247,N_27873,N_27728);
nand UO_3248 (O_3248,N_27337,N_28836);
nand UO_3249 (O_3249,N_29887,N_27268);
and UO_3250 (O_3250,N_28513,N_27341);
or UO_3251 (O_3251,N_29019,N_28252);
nand UO_3252 (O_3252,N_28567,N_29477);
xnor UO_3253 (O_3253,N_27245,N_28580);
and UO_3254 (O_3254,N_28681,N_28803);
and UO_3255 (O_3255,N_29661,N_29750);
xor UO_3256 (O_3256,N_29547,N_29804);
and UO_3257 (O_3257,N_28576,N_29145);
and UO_3258 (O_3258,N_29330,N_29561);
nand UO_3259 (O_3259,N_28185,N_28508);
and UO_3260 (O_3260,N_28966,N_28777);
nor UO_3261 (O_3261,N_27707,N_27513);
and UO_3262 (O_3262,N_27631,N_27871);
or UO_3263 (O_3263,N_29826,N_29179);
nand UO_3264 (O_3264,N_27706,N_27966);
nand UO_3265 (O_3265,N_29028,N_29316);
or UO_3266 (O_3266,N_28399,N_28566);
nand UO_3267 (O_3267,N_27640,N_28835);
nand UO_3268 (O_3268,N_27174,N_27346);
xor UO_3269 (O_3269,N_27016,N_27246);
or UO_3270 (O_3270,N_28008,N_29251);
or UO_3271 (O_3271,N_29899,N_28172);
and UO_3272 (O_3272,N_28154,N_28064);
nand UO_3273 (O_3273,N_29783,N_28577);
or UO_3274 (O_3274,N_28398,N_27911);
or UO_3275 (O_3275,N_28590,N_29704);
nor UO_3276 (O_3276,N_28028,N_28643);
nor UO_3277 (O_3277,N_27708,N_28171);
nand UO_3278 (O_3278,N_29909,N_27119);
nor UO_3279 (O_3279,N_29364,N_28565);
nand UO_3280 (O_3280,N_29895,N_29321);
nand UO_3281 (O_3281,N_27915,N_29388);
or UO_3282 (O_3282,N_27929,N_27949);
nor UO_3283 (O_3283,N_29270,N_28080);
or UO_3284 (O_3284,N_27671,N_28878);
and UO_3285 (O_3285,N_27163,N_29941);
nand UO_3286 (O_3286,N_28905,N_28255);
nand UO_3287 (O_3287,N_29843,N_27026);
nor UO_3288 (O_3288,N_28010,N_27985);
and UO_3289 (O_3289,N_28107,N_27815);
xor UO_3290 (O_3290,N_27823,N_29134);
and UO_3291 (O_3291,N_28372,N_29380);
nand UO_3292 (O_3292,N_28947,N_28683);
and UO_3293 (O_3293,N_29760,N_29199);
nor UO_3294 (O_3294,N_29861,N_29199);
nor UO_3295 (O_3295,N_29991,N_29957);
and UO_3296 (O_3296,N_27633,N_27261);
nor UO_3297 (O_3297,N_29801,N_27224);
and UO_3298 (O_3298,N_28809,N_27354);
or UO_3299 (O_3299,N_29536,N_29486);
or UO_3300 (O_3300,N_28541,N_27484);
and UO_3301 (O_3301,N_29984,N_28878);
nor UO_3302 (O_3302,N_28526,N_29620);
and UO_3303 (O_3303,N_28062,N_27619);
nand UO_3304 (O_3304,N_29042,N_28227);
or UO_3305 (O_3305,N_27412,N_27815);
or UO_3306 (O_3306,N_29428,N_29382);
xnor UO_3307 (O_3307,N_27479,N_29882);
xor UO_3308 (O_3308,N_28062,N_27926);
nand UO_3309 (O_3309,N_27566,N_28469);
or UO_3310 (O_3310,N_28947,N_28287);
xor UO_3311 (O_3311,N_27383,N_29424);
xor UO_3312 (O_3312,N_28803,N_28144);
nand UO_3313 (O_3313,N_27773,N_29252);
nor UO_3314 (O_3314,N_29093,N_29165);
or UO_3315 (O_3315,N_29386,N_27899);
nor UO_3316 (O_3316,N_28162,N_27493);
and UO_3317 (O_3317,N_29268,N_27275);
or UO_3318 (O_3318,N_27004,N_27269);
nor UO_3319 (O_3319,N_27779,N_28933);
and UO_3320 (O_3320,N_28801,N_29781);
and UO_3321 (O_3321,N_29929,N_27287);
and UO_3322 (O_3322,N_28051,N_29361);
or UO_3323 (O_3323,N_29651,N_27900);
nand UO_3324 (O_3324,N_29421,N_28055);
xor UO_3325 (O_3325,N_27992,N_28842);
nand UO_3326 (O_3326,N_27841,N_27025);
nand UO_3327 (O_3327,N_28729,N_27286);
xnor UO_3328 (O_3328,N_29788,N_27158);
nand UO_3329 (O_3329,N_29647,N_27436);
nand UO_3330 (O_3330,N_27010,N_28456);
or UO_3331 (O_3331,N_29059,N_28468);
or UO_3332 (O_3332,N_29896,N_28954);
and UO_3333 (O_3333,N_29086,N_27401);
nand UO_3334 (O_3334,N_27910,N_29794);
or UO_3335 (O_3335,N_28280,N_29806);
and UO_3336 (O_3336,N_28619,N_27859);
nand UO_3337 (O_3337,N_29231,N_28170);
xor UO_3338 (O_3338,N_27003,N_29372);
nor UO_3339 (O_3339,N_29538,N_29022);
and UO_3340 (O_3340,N_27254,N_28451);
nor UO_3341 (O_3341,N_29750,N_27499);
xor UO_3342 (O_3342,N_28993,N_29573);
xor UO_3343 (O_3343,N_29907,N_28289);
nor UO_3344 (O_3344,N_28653,N_28504);
or UO_3345 (O_3345,N_28035,N_29203);
nand UO_3346 (O_3346,N_27965,N_27722);
and UO_3347 (O_3347,N_29453,N_28529);
or UO_3348 (O_3348,N_28127,N_27529);
xor UO_3349 (O_3349,N_29999,N_28983);
or UO_3350 (O_3350,N_27741,N_28152);
or UO_3351 (O_3351,N_28138,N_27687);
nor UO_3352 (O_3352,N_29117,N_27480);
nand UO_3353 (O_3353,N_28075,N_27476);
xnor UO_3354 (O_3354,N_29291,N_28482);
xor UO_3355 (O_3355,N_27265,N_28928);
and UO_3356 (O_3356,N_29371,N_27855);
and UO_3357 (O_3357,N_28224,N_29381);
nor UO_3358 (O_3358,N_29971,N_27225);
xor UO_3359 (O_3359,N_27108,N_28472);
or UO_3360 (O_3360,N_27571,N_29208);
nand UO_3361 (O_3361,N_29236,N_27023);
xor UO_3362 (O_3362,N_27445,N_29753);
and UO_3363 (O_3363,N_27804,N_29138);
nor UO_3364 (O_3364,N_27744,N_27789);
and UO_3365 (O_3365,N_28274,N_29535);
and UO_3366 (O_3366,N_27814,N_29581);
nand UO_3367 (O_3367,N_27811,N_27724);
xor UO_3368 (O_3368,N_29670,N_27770);
xnor UO_3369 (O_3369,N_27179,N_29098);
and UO_3370 (O_3370,N_27843,N_28877);
or UO_3371 (O_3371,N_29999,N_29600);
or UO_3372 (O_3372,N_27883,N_27871);
or UO_3373 (O_3373,N_29486,N_28495);
xnor UO_3374 (O_3374,N_29586,N_27660);
and UO_3375 (O_3375,N_27746,N_27591);
xnor UO_3376 (O_3376,N_28605,N_28337);
and UO_3377 (O_3377,N_27934,N_28564);
nor UO_3378 (O_3378,N_29514,N_29288);
or UO_3379 (O_3379,N_29932,N_28824);
nor UO_3380 (O_3380,N_29224,N_29629);
nand UO_3381 (O_3381,N_28997,N_29658);
nand UO_3382 (O_3382,N_27981,N_29075);
or UO_3383 (O_3383,N_29410,N_27390);
nor UO_3384 (O_3384,N_27942,N_27774);
and UO_3385 (O_3385,N_29930,N_28357);
xor UO_3386 (O_3386,N_28554,N_27741);
or UO_3387 (O_3387,N_29027,N_29556);
and UO_3388 (O_3388,N_27633,N_27532);
and UO_3389 (O_3389,N_27176,N_28656);
or UO_3390 (O_3390,N_29465,N_28939);
nor UO_3391 (O_3391,N_29311,N_27017);
xor UO_3392 (O_3392,N_28601,N_29792);
xor UO_3393 (O_3393,N_28501,N_28753);
or UO_3394 (O_3394,N_28360,N_28430);
and UO_3395 (O_3395,N_29763,N_28486);
nor UO_3396 (O_3396,N_28011,N_27296);
and UO_3397 (O_3397,N_27757,N_27846);
xor UO_3398 (O_3398,N_27395,N_28259);
nand UO_3399 (O_3399,N_29563,N_28558);
or UO_3400 (O_3400,N_29639,N_27155);
nor UO_3401 (O_3401,N_28034,N_27073);
nand UO_3402 (O_3402,N_29750,N_29397);
and UO_3403 (O_3403,N_27397,N_29375);
nor UO_3404 (O_3404,N_28037,N_28065);
and UO_3405 (O_3405,N_29858,N_29957);
xnor UO_3406 (O_3406,N_28544,N_27173);
nor UO_3407 (O_3407,N_29682,N_28099);
nor UO_3408 (O_3408,N_27789,N_28415);
or UO_3409 (O_3409,N_27902,N_29925);
nand UO_3410 (O_3410,N_28172,N_29811);
and UO_3411 (O_3411,N_27915,N_29859);
nand UO_3412 (O_3412,N_27049,N_27572);
nor UO_3413 (O_3413,N_27509,N_29104);
xor UO_3414 (O_3414,N_29195,N_28333);
nand UO_3415 (O_3415,N_28989,N_27732);
nor UO_3416 (O_3416,N_29053,N_27633);
xnor UO_3417 (O_3417,N_27074,N_28699);
nand UO_3418 (O_3418,N_28564,N_29263);
or UO_3419 (O_3419,N_27541,N_28649);
nand UO_3420 (O_3420,N_27598,N_28824);
or UO_3421 (O_3421,N_29999,N_29013);
or UO_3422 (O_3422,N_29064,N_27586);
or UO_3423 (O_3423,N_28503,N_28245);
and UO_3424 (O_3424,N_28205,N_27894);
and UO_3425 (O_3425,N_28616,N_29522);
or UO_3426 (O_3426,N_29821,N_28290);
or UO_3427 (O_3427,N_29358,N_28154);
nor UO_3428 (O_3428,N_28631,N_27103);
xor UO_3429 (O_3429,N_28034,N_29642);
nor UO_3430 (O_3430,N_27106,N_28137);
nand UO_3431 (O_3431,N_29403,N_28842);
or UO_3432 (O_3432,N_27896,N_29852);
and UO_3433 (O_3433,N_27180,N_28324);
or UO_3434 (O_3434,N_27450,N_29265);
nand UO_3435 (O_3435,N_28888,N_29764);
nand UO_3436 (O_3436,N_29204,N_29788);
and UO_3437 (O_3437,N_29290,N_28693);
nor UO_3438 (O_3438,N_27148,N_28305);
or UO_3439 (O_3439,N_28619,N_29567);
and UO_3440 (O_3440,N_29532,N_28110);
nor UO_3441 (O_3441,N_28587,N_28254);
or UO_3442 (O_3442,N_27750,N_27153);
nand UO_3443 (O_3443,N_27484,N_29636);
or UO_3444 (O_3444,N_29681,N_29501);
and UO_3445 (O_3445,N_29533,N_29402);
or UO_3446 (O_3446,N_29532,N_28612);
nand UO_3447 (O_3447,N_29747,N_27601);
or UO_3448 (O_3448,N_28914,N_28592);
and UO_3449 (O_3449,N_27173,N_29336);
nand UO_3450 (O_3450,N_29107,N_28481);
xor UO_3451 (O_3451,N_27906,N_28729);
xor UO_3452 (O_3452,N_27054,N_27754);
xor UO_3453 (O_3453,N_29579,N_28879);
xnor UO_3454 (O_3454,N_28568,N_29232);
nand UO_3455 (O_3455,N_27023,N_28531);
or UO_3456 (O_3456,N_29668,N_28239);
and UO_3457 (O_3457,N_28496,N_28339);
nor UO_3458 (O_3458,N_29948,N_29553);
xor UO_3459 (O_3459,N_29595,N_29811);
or UO_3460 (O_3460,N_28012,N_29839);
and UO_3461 (O_3461,N_27309,N_29337);
xnor UO_3462 (O_3462,N_29866,N_28919);
and UO_3463 (O_3463,N_27960,N_27478);
or UO_3464 (O_3464,N_29039,N_29767);
xnor UO_3465 (O_3465,N_29847,N_29108);
or UO_3466 (O_3466,N_27462,N_29185);
xnor UO_3467 (O_3467,N_28923,N_28952);
and UO_3468 (O_3468,N_27156,N_28570);
and UO_3469 (O_3469,N_29579,N_28203);
xnor UO_3470 (O_3470,N_28558,N_27322);
nor UO_3471 (O_3471,N_28960,N_27851);
nand UO_3472 (O_3472,N_27934,N_29265);
nand UO_3473 (O_3473,N_27221,N_27265);
nor UO_3474 (O_3474,N_27445,N_27003);
nand UO_3475 (O_3475,N_29985,N_27849);
or UO_3476 (O_3476,N_29937,N_28140);
xnor UO_3477 (O_3477,N_27560,N_29558);
or UO_3478 (O_3478,N_27272,N_28525);
nand UO_3479 (O_3479,N_28533,N_27086);
and UO_3480 (O_3480,N_29483,N_27051);
xnor UO_3481 (O_3481,N_29609,N_27555);
nand UO_3482 (O_3482,N_28798,N_29291);
nor UO_3483 (O_3483,N_29154,N_27853);
and UO_3484 (O_3484,N_28632,N_28148);
and UO_3485 (O_3485,N_28784,N_27339);
or UO_3486 (O_3486,N_27336,N_28640);
or UO_3487 (O_3487,N_28427,N_28148);
or UO_3488 (O_3488,N_27623,N_27106);
nor UO_3489 (O_3489,N_29408,N_29161);
nor UO_3490 (O_3490,N_29679,N_27400);
or UO_3491 (O_3491,N_28134,N_29229);
xnor UO_3492 (O_3492,N_28822,N_29145);
or UO_3493 (O_3493,N_27692,N_27166);
or UO_3494 (O_3494,N_29509,N_28721);
nand UO_3495 (O_3495,N_28526,N_27546);
nor UO_3496 (O_3496,N_29381,N_27555);
and UO_3497 (O_3497,N_29030,N_29117);
xor UO_3498 (O_3498,N_27150,N_28695);
nand UO_3499 (O_3499,N_28374,N_28404);
endmodule