module basic_500_3000_500_40_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_202,In_370);
and U1 (N_1,In_27,In_372);
xnor U2 (N_2,In_339,In_115);
or U3 (N_3,In_389,In_469);
and U4 (N_4,In_496,In_277);
xor U5 (N_5,In_95,In_465);
nor U6 (N_6,In_461,In_101);
nand U7 (N_7,In_369,In_429);
or U8 (N_8,In_266,In_458);
xor U9 (N_9,In_35,In_274);
nand U10 (N_10,In_248,In_445);
xnor U11 (N_11,In_474,In_414);
and U12 (N_12,In_334,In_156);
or U13 (N_13,In_417,In_144);
nand U14 (N_14,In_270,In_160);
or U15 (N_15,In_359,In_100);
nand U16 (N_16,In_399,In_82);
or U17 (N_17,In_121,In_470);
and U18 (N_18,In_222,In_163);
and U19 (N_19,In_87,In_211);
or U20 (N_20,In_335,In_418);
nor U21 (N_21,In_21,In_215);
nor U22 (N_22,In_209,In_84);
or U23 (N_23,In_410,In_191);
or U24 (N_24,In_340,In_436);
nor U25 (N_25,In_499,In_392);
xnor U26 (N_26,In_12,In_301);
nand U27 (N_27,In_310,In_174);
xor U28 (N_28,In_381,In_261);
xnor U29 (N_29,In_18,In_498);
nand U30 (N_30,In_492,In_201);
and U31 (N_31,In_5,In_104);
or U32 (N_32,In_348,In_432);
nor U33 (N_33,In_276,In_294);
or U34 (N_34,In_168,In_46);
nand U35 (N_35,In_403,In_364);
xnor U36 (N_36,In_398,In_446);
nor U37 (N_37,In_391,In_443);
and U38 (N_38,In_118,In_90);
nand U39 (N_39,In_473,In_363);
nand U40 (N_40,In_152,In_108);
or U41 (N_41,In_493,In_377);
or U42 (N_42,In_253,In_353);
and U43 (N_43,In_302,In_350);
or U44 (N_44,In_228,In_243);
or U45 (N_45,In_70,In_162);
and U46 (N_46,In_425,In_47);
and U47 (N_47,In_400,In_89);
nand U48 (N_48,In_49,In_34);
or U49 (N_49,In_52,In_305);
nor U50 (N_50,In_472,In_42);
xnor U51 (N_51,In_246,In_44);
nor U52 (N_52,In_64,In_497);
nand U53 (N_53,In_267,In_56);
and U54 (N_54,In_286,In_236);
nor U55 (N_55,In_379,In_145);
nand U56 (N_56,In_483,In_207);
or U57 (N_57,In_91,In_176);
nand U58 (N_58,In_155,In_10);
xnor U59 (N_59,In_140,In_488);
and U60 (N_60,In_284,In_40);
or U61 (N_61,In_264,In_378);
or U62 (N_62,In_451,In_412);
xor U63 (N_63,In_252,In_29);
nor U64 (N_64,In_448,In_3);
nor U65 (N_65,In_426,In_67);
nand U66 (N_66,In_452,In_439);
or U67 (N_67,In_33,In_116);
or U68 (N_68,In_62,In_143);
and U69 (N_69,In_440,In_419);
nor U70 (N_70,In_380,In_125);
nor U71 (N_71,In_298,In_26);
xnor U72 (N_72,In_72,In_349);
and U73 (N_73,In_186,In_324);
or U74 (N_74,In_226,In_281);
and U75 (N_75,In_291,In_300);
xor U76 (N_76,N_42,In_20);
and U77 (N_77,In_329,N_25);
and U78 (N_78,In_0,In_217);
or U79 (N_79,N_52,In_311);
nand U80 (N_80,N_66,N_7);
or U81 (N_81,In_208,In_427);
xor U82 (N_82,In_124,In_135);
nand U83 (N_83,In_476,In_14);
xor U84 (N_84,In_88,In_106);
nor U85 (N_85,In_455,In_221);
nand U86 (N_86,In_107,In_203);
xor U87 (N_87,In_130,In_257);
or U88 (N_88,In_289,In_131);
nor U89 (N_89,In_312,In_109);
nand U90 (N_90,In_317,N_19);
or U91 (N_91,In_195,In_51);
xnor U92 (N_92,In_299,In_457);
or U93 (N_93,In_213,In_210);
and U94 (N_94,In_7,In_367);
and U95 (N_95,In_31,In_63);
or U96 (N_96,In_481,In_288);
or U97 (N_97,In_325,In_200);
nor U98 (N_98,N_46,In_424);
or U99 (N_99,N_68,In_245);
nand U100 (N_100,N_49,In_69);
or U101 (N_101,In_187,N_12);
nor U102 (N_102,In_113,In_61);
nand U103 (N_103,In_164,In_279);
or U104 (N_104,In_8,N_35);
or U105 (N_105,N_6,In_268);
xnor U106 (N_106,In_395,In_59);
nand U107 (N_107,N_26,In_292);
and U108 (N_108,In_447,In_468);
nor U109 (N_109,In_81,In_66);
nand U110 (N_110,In_78,N_65);
xnor U111 (N_111,In_178,In_133);
nand U112 (N_112,In_205,In_278);
and U113 (N_113,In_409,In_411);
and U114 (N_114,In_229,In_28);
nor U115 (N_115,In_464,In_265);
and U116 (N_116,In_102,In_128);
xnor U117 (N_117,In_450,In_68);
xor U118 (N_118,In_453,In_295);
nand U119 (N_119,In_111,In_73);
nor U120 (N_120,In_368,In_323);
nor U121 (N_121,In_489,In_25);
nand U122 (N_122,In_117,N_38);
xor U123 (N_123,In_313,In_309);
nand U124 (N_124,In_356,In_183);
xor U125 (N_125,In_165,N_69);
and U126 (N_126,In_149,In_132);
nor U127 (N_127,In_347,N_48);
xor U128 (N_128,In_166,In_159);
nor U129 (N_129,In_39,In_394);
xor U130 (N_130,In_431,N_53);
xor U131 (N_131,N_58,In_249);
xor U132 (N_132,N_31,In_19);
or U133 (N_133,In_13,In_303);
xor U134 (N_134,In_38,In_173);
or U135 (N_135,In_184,In_172);
nand U136 (N_136,In_224,In_79);
nor U137 (N_137,N_3,N_62);
and U138 (N_138,N_30,In_491);
or U139 (N_139,In_196,In_180);
nor U140 (N_140,In_94,In_415);
nand U141 (N_141,In_110,N_9);
and U142 (N_142,N_36,In_442);
nor U143 (N_143,In_371,In_479);
nor U144 (N_144,In_385,N_16);
xnor U145 (N_145,In_6,In_139);
xor U146 (N_146,In_74,In_471);
xnor U147 (N_147,In_456,N_73);
or U148 (N_148,In_346,In_420);
and U149 (N_149,N_72,N_47);
nand U150 (N_150,In_216,N_43);
nand U151 (N_151,In_232,N_78);
xor U152 (N_152,In_179,In_151);
nand U153 (N_153,N_85,In_322);
nor U154 (N_154,N_100,In_50);
nand U155 (N_155,N_82,In_360);
nand U156 (N_156,In_223,In_53);
nor U157 (N_157,In_123,In_404);
xnor U158 (N_158,In_197,In_251);
or U159 (N_159,In_321,In_307);
nor U160 (N_160,In_421,In_485);
nand U161 (N_161,In_230,In_283);
or U162 (N_162,In_331,In_241);
and U163 (N_163,In_199,In_161);
and U164 (N_164,N_121,In_390);
nor U165 (N_165,In_328,N_137);
nand U166 (N_166,In_147,In_57);
xnor U167 (N_167,N_135,N_113);
and U168 (N_168,N_1,N_102);
or U169 (N_169,N_98,N_119);
or U170 (N_170,N_86,In_99);
and U171 (N_171,N_27,In_343);
or U172 (N_172,In_422,In_83);
xnor U173 (N_173,In_254,In_37);
or U174 (N_174,N_34,In_76);
and U175 (N_175,In_352,N_13);
and U176 (N_176,N_142,N_64);
or U177 (N_177,In_170,In_351);
nor U178 (N_178,In_218,In_304);
nor U179 (N_179,N_110,In_233);
nor U180 (N_180,In_438,N_77);
and U181 (N_181,N_15,N_109);
nand U182 (N_182,In_129,In_240);
nor U183 (N_183,N_33,In_397);
and U184 (N_184,In_280,N_44);
nor U185 (N_185,In_262,N_14);
or U186 (N_186,N_0,In_142);
and U187 (N_187,N_148,In_361);
nor U188 (N_188,N_94,N_5);
and U189 (N_189,N_120,N_74);
nand U190 (N_190,In_290,In_9);
or U191 (N_191,N_126,In_354);
and U192 (N_192,In_285,In_484);
xnor U193 (N_193,N_136,In_169);
xor U194 (N_194,In_220,In_401);
nor U195 (N_195,In_234,In_258);
and U196 (N_196,In_387,In_96);
nand U197 (N_197,N_45,In_462);
and U198 (N_198,N_141,In_408);
nor U199 (N_199,In_15,N_4);
nand U200 (N_200,In_239,N_138);
and U201 (N_201,In_242,N_21);
and U202 (N_202,In_194,N_101);
xor U203 (N_203,N_54,In_153);
nand U204 (N_204,N_76,N_143);
nor U205 (N_205,N_106,In_382);
or U206 (N_206,In_341,In_388);
xnor U207 (N_207,In_105,In_30);
xor U208 (N_208,N_112,In_126);
or U209 (N_209,N_129,In_237);
nor U210 (N_210,In_407,N_67);
or U211 (N_211,In_65,In_428);
nor U212 (N_212,In_345,In_374);
nand U213 (N_213,In_293,In_58);
and U214 (N_214,In_263,N_130);
or U215 (N_215,In_17,In_366);
xnor U216 (N_216,In_48,N_111);
and U217 (N_217,In_138,In_55);
or U218 (N_218,N_39,In_275);
or U219 (N_219,In_60,In_454);
and U220 (N_220,N_71,In_332);
xor U221 (N_221,In_45,N_55);
nor U222 (N_222,N_96,In_141);
nor U223 (N_223,In_273,In_238);
nor U224 (N_224,In_32,In_330);
nor U225 (N_225,N_87,N_28);
nor U226 (N_226,In_247,In_198);
or U227 (N_227,In_269,N_178);
nor U228 (N_228,N_151,N_83);
or U229 (N_229,In_495,In_158);
or U230 (N_230,In_182,N_79);
and U231 (N_231,N_175,In_430);
nand U232 (N_232,In_460,In_167);
nand U233 (N_233,N_220,N_205);
xnor U234 (N_234,N_123,N_176);
or U235 (N_235,N_199,N_149);
nor U236 (N_236,N_181,N_154);
or U237 (N_237,In_41,N_93);
and U238 (N_238,N_165,In_119);
nor U239 (N_239,N_170,N_140);
nor U240 (N_240,N_133,In_486);
nand U241 (N_241,N_197,N_61);
or U242 (N_242,N_167,In_181);
xor U243 (N_243,In_342,In_137);
nor U244 (N_244,N_174,N_116);
and U245 (N_245,N_157,N_60);
nor U246 (N_246,In_225,In_77);
and U247 (N_247,N_158,N_180);
xor U248 (N_248,N_37,In_423);
or U249 (N_249,In_36,In_433);
nor U250 (N_250,N_91,N_81);
or U251 (N_251,In_375,In_4);
xor U252 (N_252,N_84,In_11);
nand U253 (N_253,N_124,In_260);
and U254 (N_254,N_18,N_59);
or U255 (N_255,N_139,N_132);
nor U256 (N_256,N_211,N_145);
nor U257 (N_257,In_190,N_92);
and U258 (N_258,N_125,In_315);
and U259 (N_259,N_97,In_206);
and U260 (N_260,N_152,N_118);
nand U261 (N_261,In_271,In_318);
nand U262 (N_262,N_156,N_212);
nor U263 (N_263,In_337,N_215);
nand U264 (N_264,In_219,In_477);
nor U265 (N_265,In_255,N_224);
xnor U266 (N_266,N_200,N_90);
xnor U267 (N_267,N_213,N_219);
or U268 (N_268,N_131,N_41);
and U269 (N_269,In_192,In_487);
nor U270 (N_270,N_75,N_177);
nand U271 (N_271,In_435,In_434);
nand U272 (N_272,In_480,In_365);
or U273 (N_273,In_384,N_191);
xnor U274 (N_274,N_210,N_206);
nor U275 (N_275,In_376,N_56);
nand U276 (N_276,N_193,N_173);
xnor U277 (N_277,N_155,N_159);
nor U278 (N_278,N_223,N_153);
nor U279 (N_279,N_171,In_150);
nand U280 (N_280,In_71,N_29);
nand U281 (N_281,In_466,In_85);
nand U282 (N_282,In_402,In_463);
and U283 (N_283,In_154,N_218);
and U284 (N_284,N_190,In_319);
nand U285 (N_285,In_326,N_22);
and U286 (N_286,In_478,In_336);
and U287 (N_287,In_250,In_355);
nor U288 (N_288,N_160,N_146);
nor U289 (N_289,N_104,In_1);
xor U290 (N_290,N_24,In_185);
and U291 (N_291,N_189,N_8);
nand U292 (N_292,In_98,N_204);
and U293 (N_293,N_122,In_308);
nand U294 (N_294,N_166,In_441);
nor U295 (N_295,In_22,In_287);
nor U296 (N_296,N_10,In_459);
xnor U297 (N_297,N_11,In_2);
and U298 (N_298,In_146,In_393);
nand U299 (N_299,In_282,In_134);
and U300 (N_300,N_198,N_150);
and U301 (N_301,N_249,N_268);
or U302 (N_302,In_114,N_89);
and U303 (N_303,N_196,N_262);
or U304 (N_304,N_201,N_273);
and U305 (N_305,N_57,In_444);
nor U306 (N_306,N_287,N_186);
nor U307 (N_307,In_188,N_284);
xor U308 (N_308,In_214,N_117);
xor U309 (N_309,N_247,N_80);
nor U310 (N_310,N_192,N_242);
nand U311 (N_311,N_234,In_256);
and U312 (N_312,N_270,In_212);
and U313 (N_313,In_193,N_32);
nor U314 (N_314,N_194,N_246);
xnor U315 (N_315,N_230,N_278);
or U316 (N_316,In_127,In_338);
and U317 (N_317,In_494,N_290);
or U318 (N_318,N_235,N_269);
nand U319 (N_319,N_209,N_179);
and U320 (N_320,N_267,N_276);
xor U321 (N_321,N_188,In_358);
nor U322 (N_322,N_285,N_70);
and U323 (N_323,N_216,N_232);
or U324 (N_324,N_134,In_333);
xor U325 (N_325,In_120,N_208);
or U326 (N_326,N_107,In_314);
nand U327 (N_327,N_17,In_93);
or U328 (N_328,N_214,N_238);
and U329 (N_329,In_54,N_40);
and U330 (N_330,In_112,In_24);
nor U331 (N_331,N_251,N_299);
or U332 (N_332,In_75,In_16);
nor U333 (N_333,In_157,N_144);
or U334 (N_334,N_105,In_482);
xor U335 (N_335,N_282,N_172);
xor U336 (N_336,In_475,In_306);
xnor U337 (N_337,N_183,In_235);
or U338 (N_338,N_185,N_225);
nor U339 (N_339,In_320,N_236);
xnor U340 (N_340,N_277,In_86);
nor U341 (N_341,In_177,N_279);
and U342 (N_342,N_280,N_239);
nand U343 (N_343,N_95,N_20);
nand U344 (N_344,N_23,N_127);
and U345 (N_345,N_51,N_202);
and U346 (N_346,N_221,In_148);
nor U347 (N_347,N_257,In_171);
nand U348 (N_348,N_203,N_298);
nor U349 (N_349,N_254,In_175);
nor U350 (N_350,N_275,N_50);
nand U351 (N_351,N_207,N_294);
or U352 (N_352,N_237,In_344);
nand U353 (N_353,N_250,In_406);
and U354 (N_354,In_449,N_296);
xnor U355 (N_355,N_63,N_245);
nor U356 (N_356,N_163,N_147);
nand U357 (N_357,N_281,In_92);
and U358 (N_358,In_227,In_204);
nand U359 (N_359,N_297,N_115);
or U360 (N_360,N_291,In_259);
xor U361 (N_361,In_103,N_231);
xnor U362 (N_362,N_272,N_226);
nor U363 (N_363,N_266,N_240);
nor U364 (N_364,N_228,In_43);
xnor U365 (N_365,N_248,N_164);
nand U366 (N_366,N_2,N_99);
nand U367 (N_367,In_23,N_271);
or U368 (N_368,N_182,In_189);
xor U369 (N_369,In_467,N_108);
nand U370 (N_370,N_184,In_362);
and U371 (N_371,N_288,In_413);
nor U372 (N_372,N_169,In_97);
xnor U373 (N_373,In_383,N_187);
and U374 (N_374,N_243,In_272);
and U375 (N_375,N_103,N_233);
xnor U376 (N_376,In_416,N_321);
nor U377 (N_377,N_229,N_358);
nor U378 (N_378,N_307,N_313);
and U379 (N_379,N_333,N_304);
xnor U380 (N_380,N_365,N_295);
nand U381 (N_381,N_363,N_227);
xor U382 (N_382,N_372,N_258);
nand U383 (N_383,N_367,N_332);
nor U384 (N_384,N_315,N_373);
nor U385 (N_385,N_293,N_309);
and U386 (N_386,N_253,In_80);
nor U387 (N_387,N_252,In_373);
nand U388 (N_388,N_346,N_341);
xnor U389 (N_389,In_357,N_328);
or U390 (N_390,N_329,N_255);
nand U391 (N_391,N_318,N_286);
nor U392 (N_392,N_324,N_330);
and U393 (N_393,N_338,N_325);
and U394 (N_394,N_340,N_264);
nor U395 (N_395,N_359,N_303);
or U396 (N_396,N_265,In_386);
and U397 (N_397,N_310,In_244);
and U398 (N_398,N_292,N_371);
or U399 (N_399,In_327,N_162);
nand U400 (N_400,N_327,N_263);
xor U401 (N_401,N_317,N_195);
nor U402 (N_402,In_231,N_334);
nor U403 (N_403,N_316,N_161);
nor U404 (N_404,N_312,N_322);
or U405 (N_405,N_260,N_256);
and U406 (N_406,N_342,N_241);
nor U407 (N_407,N_351,In_437);
or U408 (N_408,N_336,N_311);
xnor U409 (N_409,N_348,N_305);
and U410 (N_410,N_259,In_396);
or U411 (N_411,In_490,N_357);
nand U412 (N_412,N_362,N_217);
xnor U413 (N_413,N_335,N_274);
xnor U414 (N_414,N_356,N_347);
and U415 (N_415,N_354,N_337);
and U416 (N_416,N_302,In_136);
nor U417 (N_417,In_296,In_122);
and U418 (N_418,N_364,N_343);
xnor U419 (N_419,N_350,N_355);
nand U420 (N_420,N_369,N_344);
xnor U421 (N_421,N_244,N_222);
and U422 (N_422,N_308,N_314);
and U423 (N_423,In_297,N_300);
xor U424 (N_424,N_301,N_88);
or U425 (N_425,N_306,N_360);
xnor U426 (N_426,N_261,In_316);
and U427 (N_427,N_168,N_339);
and U428 (N_428,N_345,N_114);
nand U429 (N_429,N_283,N_352);
or U430 (N_430,N_374,N_331);
nand U431 (N_431,N_353,N_370);
nor U432 (N_432,N_361,N_319);
and U433 (N_433,N_349,N_326);
and U434 (N_434,N_289,In_405);
nand U435 (N_435,N_323,N_368);
xor U436 (N_436,N_366,N_128);
or U437 (N_437,N_320,N_358);
and U438 (N_438,N_317,N_356);
nor U439 (N_439,N_333,N_367);
xnor U440 (N_440,N_229,N_333);
or U441 (N_441,N_309,In_136);
or U442 (N_442,N_364,N_354);
nand U443 (N_443,N_336,N_364);
and U444 (N_444,In_327,N_350);
xnor U445 (N_445,N_354,N_340);
xnor U446 (N_446,N_315,N_306);
xor U447 (N_447,N_342,N_368);
xnor U448 (N_448,N_347,N_258);
nand U449 (N_449,In_122,N_258);
xnor U450 (N_450,N_437,N_445);
or U451 (N_451,N_434,N_386);
nor U452 (N_452,N_448,N_442);
xor U453 (N_453,N_396,N_419);
nand U454 (N_454,N_376,N_401);
xor U455 (N_455,N_414,N_384);
or U456 (N_456,N_426,N_440);
xnor U457 (N_457,N_441,N_425);
or U458 (N_458,N_435,N_428);
nand U459 (N_459,N_413,N_397);
or U460 (N_460,N_411,N_392);
or U461 (N_461,N_421,N_377);
xnor U462 (N_462,N_429,N_449);
and U463 (N_463,N_424,N_389);
or U464 (N_464,N_410,N_408);
or U465 (N_465,N_394,N_409);
nor U466 (N_466,N_378,N_444);
xnor U467 (N_467,N_391,N_405);
and U468 (N_468,N_403,N_375);
nand U469 (N_469,N_400,N_422);
or U470 (N_470,N_438,N_431);
or U471 (N_471,N_380,N_447);
nor U472 (N_472,N_420,N_393);
or U473 (N_473,N_407,N_382);
nand U474 (N_474,N_446,N_387);
xor U475 (N_475,N_379,N_390);
nand U476 (N_476,N_388,N_416);
and U477 (N_477,N_398,N_417);
or U478 (N_478,N_436,N_432);
xnor U479 (N_479,N_423,N_383);
or U480 (N_480,N_418,N_430);
nor U481 (N_481,N_415,N_427);
nand U482 (N_482,N_433,N_439);
or U483 (N_483,N_443,N_381);
nor U484 (N_484,N_399,N_406);
nand U485 (N_485,N_395,N_385);
xnor U486 (N_486,N_412,N_404);
xor U487 (N_487,N_402,N_382);
and U488 (N_488,N_422,N_390);
nand U489 (N_489,N_387,N_441);
and U490 (N_490,N_430,N_388);
and U491 (N_491,N_429,N_396);
or U492 (N_492,N_395,N_412);
and U493 (N_493,N_383,N_441);
xnor U494 (N_494,N_376,N_398);
nand U495 (N_495,N_393,N_403);
nor U496 (N_496,N_434,N_376);
and U497 (N_497,N_447,N_428);
xor U498 (N_498,N_380,N_438);
nand U499 (N_499,N_439,N_411);
and U500 (N_500,N_435,N_382);
nand U501 (N_501,N_401,N_448);
and U502 (N_502,N_389,N_437);
or U503 (N_503,N_437,N_382);
xor U504 (N_504,N_400,N_419);
xnor U505 (N_505,N_387,N_416);
nand U506 (N_506,N_402,N_433);
nand U507 (N_507,N_431,N_412);
nand U508 (N_508,N_398,N_395);
nand U509 (N_509,N_391,N_399);
and U510 (N_510,N_422,N_375);
nand U511 (N_511,N_377,N_415);
or U512 (N_512,N_442,N_422);
nor U513 (N_513,N_406,N_449);
or U514 (N_514,N_391,N_388);
xor U515 (N_515,N_384,N_397);
or U516 (N_516,N_434,N_440);
nand U517 (N_517,N_431,N_441);
and U518 (N_518,N_437,N_420);
nor U519 (N_519,N_404,N_416);
xor U520 (N_520,N_430,N_422);
nand U521 (N_521,N_390,N_413);
nand U522 (N_522,N_443,N_442);
nor U523 (N_523,N_382,N_417);
nand U524 (N_524,N_428,N_444);
xnor U525 (N_525,N_455,N_493);
nor U526 (N_526,N_524,N_523);
xor U527 (N_527,N_520,N_506);
or U528 (N_528,N_467,N_484);
nor U529 (N_529,N_509,N_465);
nor U530 (N_530,N_480,N_472);
xor U531 (N_531,N_517,N_471);
and U532 (N_532,N_481,N_477);
xnor U533 (N_533,N_462,N_492);
or U534 (N_534,N_497,N_461);
nor U535 (N_535,N_512,N_504);
nand U536 (N_536,N_502,N_479);
and U537 (N_537,N_507,N_463);
and U538 (N_538,N_519,N_518);
or U539 (N_539,N_514,N_456);
or U540 (N_540,N_508,N_483);
or U541 (N_541,N_451,N_468);
nor U542 (N_542,N_500,N_495);
nor U543 (N_543,N_459,N_460);
and U544 (N_544,N_499,N_515);
xor U545 (N_545,N_513,N_450);
nand U546 (N_546,N_458,N_470);
xor U547 (N_547,N_454,N_473);
and U548 (N_548,N_511,N_486);
and U549 (N_549,N_490,N_474);
and U550 (N_550,N_453,N_487);
nor U551 (N_551,N_521,N_485);
nor U552 (N_552,N_482,N_494);
xor U553 (N_553,N_503,N_488);
xor U554 (N_554,N_452,N_478);
or U555 (N_555,N_510,N_466);
xnor U556 (N_556,N_522,N_491);
xnor U557 (N_557,N_489,N_501);
xor U558 (N_558,N_464,N_457);
xnor U559 (N_559,N_505,N_469);
nor U560 (N_560,N_516,N_496);
and U561 (N_561,N_475,N_498);
nor U562 (N_562,N_476,N_498);
xnor U563 (N_563,N_516,N_452);
nor U564 (N_564,N_507,N_504);
nor U565 (N_565,N_452,N_482);
nand U566 (N_566,N_497,N_523);
xnor U567 (N_567,N_481,N_460);
nand U568 (N_568,N_457,N_508);
or U569 (N_569,N_502,N_457);
or U570 (N_570,N_468,N_520);
nand U571 (N_571,N_516,N_465);
or U572 (N_572,N_476,N_505);
nor U573 (N_573,N_502,N_487);
and U574 (N_574,N_466,N_520);
and U575 (N_575,N_476,N_516);
xor U576 (N_576,N_474,N_489);
nand U577 (N_577,N_459,N_524);
or U578 (N_578,N_513,N_478);
nand U579 (N_579,N_467,N_470);
or U580 (N_580,N_505,N_455);
and U581 (N_581,N_488,N_502);
and U582 (N_582,N_504,N_474);
or U583 (N_583,N_450,N_493);
or U584 (N_584,N_510,N_517);
nor U585 (N_585,N_492,N_463);
nand U586 (N_586,N_480,N_488);
xnor U587 (N_587,N_491,N_515);
nand U588 (N_588,N_501,N_498);
nor U589 (N_589,N_469,N_487);
nand U590 (N_590,N_464,N_481);
or U591 (N_591,N_485,N_452);
nand U592 (N_592,N_523,N_450);
nor U593 (N_593,N_520,N_453);
and U594 (N_594,N_490,N_457);
and U595 (N_595,N_515,N_490);
and U596 (N_596,N_466,N_486);
xnor U597 (N_597,N_460,N_471);
or U598 (N_598,N_518,N_514);
nand U599 (N_599,N_475,N_502);
xor U600 (N_600,N_552,N_580);
nor U601 (N_601,N_597,N_599);
and U602 (N_602,N_584,N_572);
or U603 (N_603,N_563,N_542);
and U604 (N_604,N_585,N_587);
xnor U605 (N_605,N_548,N_537);
nand U606 (N_606,N_562,N_539);
nor U607 (N_607,N_568,N_594);
and U608 (N_608,N_543,N_531);
and U609 (N_609,N_554,N_574);
nand U610 (N_610,N_576,N_550);
xnor U611 (N_611,N_598,N_591);
nand U612 (N_612,N_545,N_564);
xnor U613 (N_613,N_535,N_556);
xnor U614 (N_614,N_527,N_561);
nand U615 (N_615,N_577,N_551);
xnor U616 (N_616,N_528,N_592);
nor U617 (N_617,N_532,N_579);
and U618 (N_618,N_553,N_525);
or U619 (N_619,N_566,N_544);
nand U620 (N_620,N_593,N_582);
and U621 (N_621,N_555,N_570);
xor U622 (N_622,N_573,N_583);
nor U623 (N_623,N_557,N_578);
or U624 (N_624,N_541,N_589);
nor U625 (N_625,N_586,N_526);
and U626 (N_626,N_595,N_558);
nand U627 (N_627,N_546,N_560);
or U628 (N_628,N_559,N_529);
and U629 (N_629,N_538,N_533);
xor U630 (N_630,N_567,N_596);
xnor U631 (N_631,N_569,N_575);
or U632 (N_632,N_530,N_540);
xor U633 (N_633,N_565,N_590);
nand U634 (N_634,N_547,N_549);
xor U635 (N_635,N_571,N_588);
or U636 (N_636,N_581,N_534);
and U637 (N_637,N_536,N_577);
or U638 (N_638,N_559,N_558);
and U639 (N_639,N_565,N_578);
or U640 (N_640,N_547,N_540);
nor U641 (N_641,N_530,N_579);
nor U642 (N_642,N_579,N_573);
xor U643 (N_643,N_526,N_542);
or U644 (N_644,N_560,N_549);
and U645 (N_645,N_572,N_585);
nor U646 (N_646,N_596,N_565);
nor U647 (N_647,N_551,N_549);
or U648 (N_648,N_561,N_552);
and U649 (N_649,N_592,N_593);
nand U650 (N_650,N_570,N_554);
nand U651 (N_651,N_561,N_545);
nor U652 (N_652,N_529,N_543);
nor U653 (N_653,N_530,N_599);
nor U654 (N_654,N_573,N_591);
nand U655 (N_655,N_571,N_590);
nand U656 (N_656,N_535,N_533);
and U657 (N_657,N_598,N_531);
and U658 (N_658,N_574,N_572);
and U659 (N_659,N_586,N_580);
xor U660 (N_660,N_571,N_527);
and U661 (N_661,N_593,N_539);
xor U662 (N_662,N_591,N_545);
or U663 (N_663,N_537,N_574);
nand U664 (N_664,N_547,N_539);
nand U665 (N_665,N_565,N_568);
nor U666 (N_666,N_570,N_553);
and U667 (N_667,N_550,N_535);
nor U668 (N_668,N_585,N_556);
nor U669 (N_669,N_544,N_538);
and U670 (N_670,N_557,N_551);
or U671 (N_671,N_594,N_562);
or U672 (N_672,N_594,N_550);
or U673 (N_673,N_557,N_558);
or U674 (N_674,N_528,N_583);
xnor U675 (N_675,N_616,N_661);
xnor U676 (N_676,N_649,N_653);
nor U677 (N_677,N_652,N_623);
nand U678 (N_678,N_646,N_626);
xor U679 (N_679,N_651,N_607);
and U680 (N_680,N_628,N_637);
nor U681 (N_681,N_604,N_617);
or U682 (N_682,N_610,N_638);
xor U683 (N_683,N_621,N_609);
or U684 (N_684,N_664,N_668);
xor U685 (N_685,N_656,N_658);
nand U686 (N_686,N_647,N_613);
or U687 (N_687,N_643,N_640);
nand U688 (N_688,N_650,N_670);
xnor U689 (N_689,N_615,N_618);
nand U690 (N_690,N_620,N_654);
nand U691 (N_691,N_659,N_612);
and U692 (N_692,N_672,N_632);
and U693 (N_693,N_603,N_600);
and U694 (N_694,N_619,N_641);
or U695 (N_695,N_669,N_630);
nand U696 (N_696,N_655,N_633);
nand U697 (N_697,N_660,N_673);
nand U698 (N_698,N_624,N_642);
or U699 (N_699,N_606,N_605);
nor U700 (N_700,N_627,N_635);
and U701 (N_701,N_601,N_665);
nand U702 (N_702,N_648,N_602);
nand U703 (N_703,N_663,N_636);
nand U704 (N_704,N_674,N_631);
nor U705 (N_705,N_622,N_634);
nor U706 (N_706,N_625,N_611);
nand U707 (N_707,N_671,N_657);
and U708 (N_708,N_608,N_667);
and U709 (N_709,N_662,N_629);
and U710 (N_710,N_666,N_644);
nor U711 (N_711,N_639,N_645);
xnor U712 (N_712,N_614,N_656);
and U713 (N_713,N_617,N_671);
xnor U714 (N_714,N_646,N_634);
and U715 (N_715,N_660,N_664);
nand U716 (N_716,N_614,N_647);
nand U717 (N_717,N_654,N_631);
xor U718 (N_718,N_641,N_600);
nand U719 (N_719,N_654,N_656);
or U720 (N_720,N_654,N_612);
xnor U721 (N_721,N_614,N_627);
nor U722 (N_722,N_658,N_655);
nor U723 (N_723,N_611,N_671);
or U724 (N_724,N_667,N_636);
nand U725 (N_725,N_656,N_666);
or U726 (N_726,N_643,N_661);
and U727 (N_727,N_616,N_669);
xnor U728 (N_728,N_606,N_619);
xor U729 (N_729,N_621,N_642);
nand U730 (N_730,N_665,N_667);
nand U731 (N_731,N_630,N_639);
and U732 (N_732,N_660,N_648);
nand U733 (N_733,N_626,N_667);
nand U734 (N_734,N_623,N_632);
nor U735 (N_735,N_618,N_628);
nand U736 (N_736,N_666,N_662);
xor U737 (N_737,N_632,N_665);
and U738 (N_738,N_667,N_646);
nor U739 (N_739,N_643,N_663);
or U740 (N_740,N_662,N_656);
xor U741 (N_741,N_610,N_606);
and U742 (N_742,N_617,N_660);
nor U743 (N_743,N_621,N_673);
nand U744 (N_744,N_630,N_622);
and U745 (N_745,N_656,N_635);
nor U746 (N_746,N_667,N_656);
or U747 (N_747,N_651,N_643);
nor U748 (N_748,N_647,N_661);
or U749 (N_749,N_664,N_619);
or U750 (N_750,N_676,N_693);
xor U751 (N_751,N_719,N_739);
nand U752 (N_752,N_721,N_708);
and U753 (N_753,N_731,N_701);
xor U754 (N_754,N_710,N_725);
nand U755 (N_755,N_684,N_738);
xnor U756 (N_756,N_730,N_727);
nor U757 (N_757,N_709,N_702);
xnor U758 (N_758,N_711,N_675);
nor U759 (N_759,N_740,N_677);
nand U760 (N_760,N_746,N_698);
nand U761 (N_761,N_722,N_712);
and U762 (N_762,N_682,N_742);
xor U763 (N_763,N_694,N_747);
or U764 (N_764,N_723,N_745);
or U765 (N_765,N_741,N_706);
and U766 (N_766,N_703,N_692);
or U767 (N_767,N_680,N_685);
nand U768 (N_768,N_687,N_716);
and U769 (N_769,N_696,N_724);
or U770 (N_770,N_733,N_715);
xor U771 (N_771,N_704,N_734);
xnor U772 (N_772,N_705,N_697);
and U773 (N_773,N_713,N_695);
or U774 (N_774,N_688,N_720);
xor U775 (N_775,N_735,N_744);
and U776 (N_776,N_690,N_678);
and U777 (N_777,N_686,N_726);
nand U778 (N_778,N_743,N_683);
and U779 (N_779,N_717,N_689);
and U780 (N_780,N_699,N_748);
xor U781 (N_781,N_718,N_679);
and U782 (N_782,N_729,N_732);
and U783 (N_783,N_700,N_691);
xor U784 (N_784,N_728,N_707);
nor U785 (N_785,N_737,N_714);
nor U786 (N_786,N_736,N_749);
or U787 (N_787,N_681,N_741);
xor U788 (N_788,N_735,N_737);
and U789 (N_789,N_685,N_708);
and U790 (N_790,N_736,N_678);
nand U791 (N_791,N_696,N_700);
or U792 (N_792,N_689,N_743);
nand U793 (N_793,N_732,N_685);
nand U794 (N_794,N_722,N_723);
or U795 (N_795,N_699,N_696);
nand U796 (N_796,N_714,N_745);
nand U797 (N_797,N_700,N_699);
or U798 (N_798,N_704,N_685);
xnor U799 (N_799,N_726,N_701);
and U800 (N_800,N_726,N_745);
nor U801 (N_801,N_735,N_717);
or U802 (N_802,N_700,N_704);
xor U803 (N_803,N_680,N_706);
nor U804 (N_804,N_739,N_730);
and U805 (N_805,N_726,N_718);
or U806 (N_806,N_713,N_732);
xnor U807 (N_807,N_736,N_732);
and U808 (N_808,N_693,N_708);
or U809 (N_809,N_742,N_741);
or U810 (N_810,N_746,N_697);
nor U811 (N_811,N_698,N_692);
nor U812 (N_812,N_737,N_688);
nor U813 (N_813,N_717,N_720);
xnor U814 (N_814,N_704,N_697);
xnor U815 (N_815,N_736,N_714);
nand U816 (N_816,N_696,N_732);
nor U817 (N_817,N_715,N_725);
nor U818 (N_818,N_713,N_733);
or U819 (N_819,N_736,N_685);
nor U820 (N_820,N_721,N_726);
nor U821 (N_821,N_723,N_729);
xor U822 (N_822,N_737,N_729);
nand U823 (N_823,N_717,N_746);
nor U824 (N_824,N_736,N_720);
xor U825 (N_825,N_798,N_751);
or U826 (N_826,N_782,N_822);
nor U827 (N_827,N_770,N_786);
and U828 (N_828,N_760,N_755);
and U829 (N_829,N_792,N_819);
xnor U830 (N_830,N_762,N_795);
and U831 (N_831,N_815,N_820);
xor U832 (N_832,N_750,N_775);
nand U833 (N_833,N_752,N_768);
nor U834 (N_834,N_804,N_773);
nor U835 (N_835,N_780,N_817);
nand U836 (N_836,N_808,N_806);
or U837 (N_837,N_754,N_794);
nor U838 (N_838,N_769,N_793);
nand U839 (N_839,N_805,N_783);
xor U840 (N_840,N_759,N_761);
or U841 (N_841,N_789,N_824);
nand U842 (N_842,N_778,N_799);
xor U843 (N_843,N_813,N_764);
nor U844 (N_844,N_818,N_814);
and U845 (N_845,N_756,N_801);
and U846 (N_846,N_785,N_800);
xnor U847 (N_847,N_781,N_758);
xor U848 (N_848,N_772,N_816);
nand U849 (N_849,N_776,N_753);
xnor U850 (N_850,N_763,N_796);
or U851 (N_851,N_757,N_790);
or U852 (N_852,N_787,N_807);
nor U853 (N_853,N_771,N_823);
nand U854 (N_854,N_812,N_777);
xnor U855 (N_855,N_784,N_810);
or U856 (N_856,N_809,N_797);
xor U857 (N_857,N_774,N_779);
nand U858 (N_858,N_802,N_791);
nand U859 (N_859,N_765,N_811);
nor U860 (N_860,N_803,N_767);
nor U861 (N_861,N_788,N_821);
nand U862 (N_862,N_766,N_780);
or U863 (N_863,N_823,N_812);
xnor U864 (N_864,N_794,N_786);
and U865 (N_865,N_824,N_791);
nand U866 (N_866,N_793,N_754);
nor U867 (N_867,N_773,N_781);
and U868 (N_868,N_752,N_805);
or U869 (N_869,N_765,N_780);
and U870 (N_870,N_759,N_778);
nor U871 (N_871,N_784,N_767);
or U872 (N_872,N_766,N_784);
and U873 (N_873,N_803,N_811);
and U874 (N_874,N_761,N_762);
or U875 (N_875,N_811,N_760);
nor U876 (N_876,N_790,N_797);
xor U877 (N_877,N_818,N_792);
nor U878 (N_878,N_801,N_817);
nand U879 (N_879,N_797,N_812);
nand U880 (N_880,N_785,N_765);
nand U881 (N_881,N_775,N_763);
and U882 (N_882,N_763,N_793);
or U883 (N_883,N_775,N_789);
or U884 (N_884,N_783,N_784);
xnor U885 (N_885,N_782,N_784);
nor U886 (N_886,N_787,N_755);
nor U887 (N_887,N_755,N_822);
nor U888 (N_888,N_820,N_775);
xnor U889 (N_889,N_761,N_782);
or U890 (N_890,N_777,N_809);
and U891 (N_891,N_759,N_790);
xor U892 (N_892,N_798,N_773);
xnor U893 (N_893,N_799,N_816);
nand U894 (N_894,N_755,N_786);
xnor U895 (N_895,N_813,N_793);
or U896 (N_896,N_820,N_813);
xnor U897 (N_897,N_797,N_788);
nand U898 (N_898,N_775,N_802);
nand U899 (N_899,N_757,N_755);
xnor U900 (N_900,N_860,N_899);
xor U901 (N_901,N_846,N_889);
and U902 (N_902,N_886,N_891);
and U903 (N_903,N_898,N_840);
nor U904 (N_904,N_895,N_838);
and U905 (N_905,N_867,N_848);
or U906 (N_906,N_873,N_883);
nand U907 (N_907,N_855,N_879);
xnor U908 (N_908,N_837,N_884);
nand U909 (N_909,N_835,N_826);
nor U910 (N_910,N_857,N_865);
xor U911 (N_911,N_874,N_872);
and U912 (N_912,N_869,N_849);
or U913 (N_913,N_829,N_853);
nand U914 (N_914,N_854,N_862);
or U915 (N_915,N_827,N_839);
nor U916 (N_916,N_871,N_893);
xnor U917 (N_917,N_866,N_864);
and U918 (N_918,N_887,N_842);
and U919 (N_919,N_845,N_897);
xor U920 (N_920,N_885,N_832);
and U921 (N_921,N_878,N_861);
nor U922 (N_922,N_847,N_831);
and U923 (N_923,N_859,N_841);
and U924 (N_924,N_888,N_833);
nor U925 (N_925,N_890,N_894);
nand U926 (N_926,N_896,N_876);
or U927 (N_927,N_843,N_830);
and U928 (N_928,N_892,N_870);
or U929 (N_929,N_852,N_880);
nor U930 (N_930,N_844,N_851);
and U931 (N_931,N_858,N_863);
nand U932 (N_932,N_881,N_875);
nand U933 (N_933,N_868,N_825);
or U934 (N_934,N_828,N_856);
nor U935 (N_935,N_836,N_850);
and U936 (N_936,N_877,N_882);
and U937 (N_937,N_834,N_835);
and U938 (N_938,N_867,N_855);
nor U939 (N_939,N_895,N_873);
or U940 (N_940,N_835,N_888);
xor U941 (N_941,N_872,N_831);
nor U942 (N_942,N_862,N_874);
nor U943 (N_943,N_896,N_864);
and U944 (N_944,N_849,N_876);
nor U945 (N_945,N_825,N_867);
xor U946 (N_946,N_849,N_891);
and U947 (N_947,N_879,N_841);
nand U948 (N_948,N_825,N_845);
xnor U949 (N_949,N_898,N_864);
and U950 (N_950,N_858,N_876);
nor U951 (N_951,N_890,N_881);
and U952 (N_952,N_856,N_831);
or U953 (N_953,N_887,N_859);
nor U954 (N_954,N_835,N_875);
nor U955 (N_955,N_886,N_894);
nand U956 (N_956,N_862,N_841);
nor U957 (N_957,N_871,N_876);
xor U958 (N_958,N_895,N_884);
or U959 (N_959,N_828,N_840);
or U960 (N_960,N_842,N_892);
nand U961 (N_961,N_881,N_876);
nand U962 (N_962,N_853,N_887);
xnor U963 (N_963,N_863,N_888);
or U964 (N_964,N_856,N_849);
and U965 (N_965,N_853,N_882);
or U966 (N_966,N_865,N_831);
or U967 (N_967,N_845,N_887);
nor U968 (N_968,N_886,N_846);
xnor U969 (N_969,N_848,N_845);
nor U970 (N_970,N_860,N_861);
or U971 (N_971,N_866,N_892);
nor U972 (N_972,N_897,N_863);
and U973 (N_973,N_868,N_867);
nand U974 (N_974,N_887,N_889);
and U975 (N_975,N_943,N_948);
xor U976 (N_976,N_921,N_970);
and U977 (N_977,N_922,N_936);
and U978 (N_978,N_967,N_949);
xor U979 (N_979,N_904,N_969);
or U980 (N_980,N_950,N_918);
xor U981 (N_981,N_944,N_947);
nor U982 (N_982,N_939,N_937);
xor U983 (N_983,N_928,N_910);
and U984 (N_984,N_938,N_905);
xor U985 (N_985,N_902,N_908);
xnor U986 (N_986,N_920,N_912);
nor U987 (N_987,N_966,N_946);
xor U988 (N_988,N_913,N_915);
nor U989 (N_989,N_907,N_951);
or U990 (N_990,N_952,N_960);
and U991 (N_991,N_926,N_903);
and U992 (N_992,N_914,N_933);
nor U993 (N_993,N_962,N_953);
xnor U994 (N_994,N_974,N_929);
nand U995 (N_995,N_942,N_924);
xnor U996 (N_996,N_963,N_935);
and U997 (N_997,N_956,N_911);
nand U998 (N_998,N_901,N_959);
xor U999 (N_999,N_954,N_934);
or U1000 (N_1000,N_916,N_925);
nand U1001 (N_1001,N_945,N_971);
xnor U1002 (N_1002,N_973,N_923);
and U1003 (N_1003,N_917,N_940);
xor U1004 (N_1004,N_927,N_909);
nand U1005 (N_1005,N_941,N_932);
or U1006 (N_1006,N_968,N_919);
xor U1007 (N_1007,N_972,N_958);
xor U1008 (N_1008,N_955,N_964);
xor U1009 (N_1009,N_900,N_961);
or U1010 (N_1010,N_906,N_965);
and U1011 (N_1011,N_931,N_957);
and U1012 (N_1012,N_930,N_970);
xnor U1013 (N_1013,N_900,N_920);
nor U1014 (N_1014,N_903,N_943);
nand U1015 (N_1015,N_939,N_941);
nand U1016 (N_1016,N_966,N_971);
and U1017 (N_1017,N_927,N_966);
nor U1018 (N_1018,N_928,N_946);
nor U1019 (N_1019,N_917,N_946);
xnor U1020 (N_1020,N_912,N_916);
nor U1021 (N_1021,N_921,N_972);
nand U1022 (N_1022,N_932,N_963);
xor U1023 (N_1023,N_951,N_908);
and U1024 (N_1024,N_961,N_956);
nor U1025 (N_1025,N_903,N_952);
or U1026 (N_1026,N_934,N_911);
and U1027 (N_1027,N_943,N_966);
xnor U1028 (N_1028,N_930,N_937);
and U1029 (N_1029,N_908,N_935);
nand U1030 (N_1030,N_903,N_908);
xor U1031 (N_1031,N_928,N_955);
or U1032 (N_1032,N_973,N_904);
nand U1033 (N_1033,N_914,N_968);
and U1034 (N_1034,N_911,N_932);
xnor U1035 (N_1035,N_918,N_919);
nand U1036 (N_1036,N_963,N_910);
nand U1037 (N_1037,N_940,N_971);
and U1038 (N_1038,N_930,N_955);
nand U1039 (N_1039,N_940,N_913);
nor U1040 (N_1040,N_900,N_918);
nand U1041 (N_1041,N_900,N_903);
xnor U1042 (N_1042,N_952,N_942);
and U1043 (N_1043,N_956,N_929);
xor U1044 (N_1044,N_927,N_940);
nand U1045 (N_1045,N_964,N_902);
xor U1046 (N_1046,N_931,N_904);
or U1047 (N_1047,N_940,N_901);
or U1048 (N_1048,N_919,N_958);
and U1049 (N_1049,N_959,N_952);
or U1050 (N_1050,N_1026,N_1019);
and U1051 (N_1051,N_992,N_1041);
xnor U1052 (N_1052,N_996,N_1037);
nor U1053 (N_1053,N_975,N_1033);
and U1054 (N_1054,N_1008,N_1040);
nor U1055 (N_1055,N_1016,N_1031);
and U1056 (N_1056,N_994,N_1021);
or U1057 (N_1057,N_1046,N_1004);
nor U1058 (N_1058,N_1017,N_989);
or U1059 (N_1059,N_980,N_995);
xnor U1060 (N_1060,N_1015,N_1042);
nor U1061 (N_1061,N_1035,N_1049);
and U1062 (N_1062,N_1047,N_1012);
nand U1063 (N_1063,N_979,N_986);
and U1064 (N_1064,N_1039,N_1036);
xor U1065 (N_1065,N_982,N_997);
nor U1066 (N_1066,N_1043,N_978);
xor U1067 (N_1067,N_1023,N_1025);
nor U1068 (N_1068,N_1007,N_1044);
and U1069 (N_1069,N_1032,N_998);
or U1070 (N_1070,N_1028,N_983);
nand U1071 (N_1071,N_981,N_1020);
and U1072 (N_1072,N_1009,N_984);
nand U1073 (N_1073,N_993,N_1048);
and U1074 (N_1074,N_1034,N_987);
and U1075 (N_1075,N_1024,N_1005);
nand U1076 (N_1076,N_1038,N_1001);
or U1077 (N_1077,N_977,N_1030);
nand U1078 (N_1078,N_1002,N_1022);
nand U1079 (N_1079,N_990,N_991);
or U1080 (N_1080,N_1003,N_1014);
and U1081 (N_1081,N_1000,N_988);
or U1082 (N_1082,N_1018,N_1045);
and U1083 (N_1083,N_1027,N_985);
xor U1084 (N_1084,N_999,N_1006);
and U1085 (N_1085,N_1029,N_1011);
nand U1086 (N_1086,N_1010,N_1013);
xor U1087 (N_1087,N_976,N_1031);
and U1088 (N_1088,N_1022,N_998);
nor U1089 (N_1089,N_1023,N_1002);
nand U1090 (N_1090,N_984,N_1011);
and U1091 (N_1091,N_985,N_1030);
or U1092 (N_1092,N_999,N_982);
nor U1093 (N_1093,N_993,N_1005);
or U1094 (N_1094,N_1039,N_1020);
nor U1095 (N_1095,N_1038,N_1008);
nor U1096 (N_1096,N_1006,N_1035);
nand U1097 (N_1097,N_1041,N_975);
nor U1098 (N_1098,N_979,N_976);
nand U1099 (N_1099,N_1011,N_1037);
nand U1100 (N_1100,N_1006,N_1021);
xnor U1101 (N_1101,N_979,N_999);
xnor U1102 (N_1102,N_985,N_1028);
or U1103 (N_1103,N_1037,N_1047);
and U1104 (N_1104,N_1031,N_987);
nor U1105 (N_1105,N_983,N_987);
or U1106 (N_1106,N_1031,N_1042);
nor U1107 (N_1107,N_992,N_1006);
or U1108 (N_1108,N_1037,N_1012);
xnor U1109 (N_1109,N_1017,N_982);
or U1110 (N_1110,N_991,N_1010);
nor U1111 (N_1111,N_1028,N_998);
nand U1112 (N_1112,N_1043,N_985);
xnor U1113 (N_1113,N_1043,N_1019);
or U1114 (N_1114,N_1003,N_1024);
and U1115 (N_1115,N_992,N_1011);
or U1116 (N_1116,N_997,N_1021);
and U1117 (N_1117,N_979,N_1014);
nand U1118 (N_1118,N_994,N_1000);
and U1119 (N_1119,N_1041,N_1008);
or U1120 (N_1120,N_1025,N_1003);
xnor U1121 (N_1121,N_1048,N_999);
nand U1122 (N_1122,N_1009,N_1020);
and U1123 (N_1123,N_1037,N_1014);
nand U1124 (N_1124,N_1001,N_1043);
nand U1125 (N_1125,N_1121,N_1061);
xor U1126 (N_1126,N_1103,N_1082);
or U1127 (N_1127,N_1102,N_1050);
nand U1128 (N_1128,N_1086,N_1119);
nor U1129 (N_1129,N_1088,N_1099);
nand U1130 (N_1130,N_1118,N_1078);
and U1131 (N_1131,N_1063,N_1053);
or U1132 (N_1132,N_1062,N_1092);
nor U1133 (N_1133,N_1066,N_1064);
nand U1134 (N_1134,N_1105,N_1090);
or U1135 (N_1135,N_1079,N_1055);
or U1136 (N_1136,N_1122,N_1070);
xor U1137 (N_1137,N_1104,N_1091);
nand U1138 (N_1138,N_1120,N_1112);
nand U1139 (N_1139,N_1089,N_1097);
nand U1140 (N_1140,N_1095,N_1074);
nand U1141 (N_1141,N_1116,N_1108);
nand U1142 (N_1142,N_1051,N_1100);
nor U1143 (N_1143,N_1060,N_1077);
xnor U1144 (N_1144,N_1107,N_1084);
nand U1145 (N_1145,N_1058,N_1081);
nor U1146 (N_1146,N_1071,N_1059);
xnor U1147 (N_1147,N_1073,N_1113);
nor U1148 (N_1148,N_1101,N_1124);
xor U1149 (N_1149,N_1111,N_1069);
nor U1150 (N_1150,N_1052,N_1106);
nor U1151 (N_1151,N_1072,N_1085);
nor U1152 (N_1152,N_1109,N_1083);
nand U1153 (N_1153,N_1067,N_1065);
or U1154 (N_1154,N_1068,N_1115);
xnor U1155 (N_1155,N_1123,N_1080);
and U1156 (N_1156,N_1110,N_1114);
nor U1157 (N_1157,N_1117,N_1054);
nor U1158 (N_1158,N_1096,N_1076);
nand U1159 (N_1159,N_1094,N_1098);
nor U1160 (N_1160,N_1075,N_1057);
or U1161 (N_1161,N_1056,N_1087);
and U1162 (N_1162,N_1093,N_1079);
xnor U1163 (N_1163,N_1120,N_1072);
xor U1164 (N_1164,N_1052,N_1082);
xor U1165 (N_1165,N_1102,N_1058);
xnor U1166 (N_1166,N_1078,N_1066);
xor U1167 (N_1167,N_1057,N_1051);
nor U1168 (N_1168,N_1067,N_1076);
xnor U1169 (N_1169,N_1064,N_1067);
xor U1170 (N_1170,N_1064,N_1084);
or U1171 (N_1171,N_1079,N_1074);
xnor U1172 (N_1172,N_1073,N_1078);
or U1173 (N_1173,N_1123,N_1065);
nor U1174 (N_1174,N_1099,N_1066);
nand U1175 (N_1175,N_1116,N_1078);
nand U1176 (N_1176,N_1121,N_1064);
nand U1177 (N_1177,N_1075,N_1119);
xnor U1178 (N_1178,N_1068,N_1060);
xor U1179 (N_1179,N_1060,N_1105);
nand U1180 (N_1180,N_1066,N_1056);
or U1181 (N_1181,N_1106,N_1095);
or U1182 (N_1182,N_1070,N_1124);
nor U1183 (N_1183,N_1102,N_1091);
nor U1184 (N_1184,N_1050,N_1068);
nor U1185 (N_1185,N_1076,N_1091);
nand U1186 (N_1186,N_1122,N_1068);
and U1187 (N_1187,N_1086,N_1050);
or U1188 (N_1188,N_1119,N_1089);
or U1189 (N_1189,N_1113,N_1090);
nor U1190 (N_1190,N_1079,N_1116);
nand U1191 (N_1191,N_1096,N_1109);
or U1192 (N_1192,N_1067,N_1086);
nor U1193 (N_1193,N_1060,N_1067);
nor U1194 (N_1194,N_1081,N_1097);
xor U1195 (N_1195,N_1052,N_1058);
nor U1196 (N_1196,N_1065,N_1087);
and U1197 (N_1197,N_1067,N_1113);
nor U1198 (N_1198,N_1110,N_1103);
nand U1199 (N_1199,N_1101,N_1102);
and U1200 (N_1200,N_1142,N_1180);
or U1201 (N_1201,N_1185,N_1189);
nand U1202 (N_1202,N_1195,N_1182);
nor U1203 (N_1203,N_1176,N_1199);
or U1204 (N_1204,N_1173,N_1145);
nand U1205 (N_1205,N_1193,N_1174);
xor U1206 (N_1206,N_1139,N_1163);
nor U1207 (N_1207,N_1156,N_1184);
and U1208 (N_1208,N_1164,N_1157);
nor U1209 (N_1209,N_1168,N_1147);
nand U1210 (N_1210,N_1167,N_1165);
nand U1211 (N_1211,N_1188,N_1136);
nand U1212 (N_1212,N_1170,N_1175);
or U1213 (N_1213,N_1190,N_1140);
xor U1214 (N_1214,N_1162,N_1192);
or U1215 (N_1215,N_1153,N_1178);
nand U1216 (N_1216,N_1135,N_1166);
nand U1217 (N_1217,N_1134,N_1172);
xor U1218 (N_1218,N_1197,N_1150);
and U1219 (N_1219,N_1160,N_1196);
or U1220 (N_1220,N_1128,N_1177);
or U1221 (N_1221,N_1138,N_1159);
xor U1222 (N_1222,N_1126,N_1194);
xor U1223 (N_1223,N_1141,N_1151);
xor U1224 (N_1224,N_1158,N_1169);
nand U1225 (N_1225,N_1144,N_1148);
nor U1226 (N_1226,N_1149,N_1132);
nand U1227 (N_1227,N_1146,N_1133);
nand U1228 (N_1228,N_1130,N_1171);
nand U1229 (N_1229,N_1129,N_1198);
xnor U1230 (N_1230,N_1181,N_1143);
nand U1231 (N_1231,N_1131,N_1187);
nor U1232 (N_1232,N_1155,N_1127);
or U1233 (N_1233,N_1137,N_1186);
xnor U1234 (N_1234,N_1152,N_1183);
nand U1235 (N_1235,N_1125,N_1154);
nand U1236 (N_1236,N_1191,N_1179);
or U1237 (N_1237,N_1161,N_1125);
nand U1238 (N_1238,N_1171,N_1149);
xnor U1239 (N_1239,N_1178,N_1156);
or U1240 (N_1240,N_1153,N_1143);
or U1241 (N_1241,N_1184,N_1181);
nand U1242 (N_1242,N_1136,N_1127);
nand U1243 (N_1243,N_1191,N_1168);
xor U1244 (N_1244,N_1125,N_1165);
or U1245 (N_1245,N_1158,N_1141);
nand U1246 (N_1246,N_1197,N_1185);
nor U1247 (N_1247,N_1157,N_1140);
nand U1248 (N_1248,N_1173,N_1170);
or U1249 (N_1249,N_1180,N_1159);
nand U1250 (N_1250,N_1161,N_1139);
and U1251 (N_1251,N_1167,N_1145);
xnor U1252 (N_1252,N_1140,N_1177);
nor U1253 (N_1253,N_1125,N_1170);
xor U1254 (N_1254,N_1128,N_1199);
nand U1255 (N_1255,N_1189,N_1180);
nor U1256 (N_1256,N_1188,N_1130);
nor U1257 (N_1257,N_1183,N_1184);
nor U1258 (N_1258,N_1138,N_1165);
and U1259 (N_1259,N_1193,N_1176);
nand U1260 (N_1260,N_1160,N_1135);
nor U1261 (N_1261,N_1146,N_1193);
or U1262 (N_1262,N_1192,N_1176);
xor U1263 (N_1263,N_1190,N_1164);
and U1264 (N_1264,N_1198,N_1157);
nand U1265 (N_1265,N_1165,N_1152);
xnor U1266 (N_1266,N_1151,N_1192);
nor U1267 (N_1267,N_1146,N_1150);
or U1268 (N_1268,N_1170,N_1130);
nor U1269 (N_1269,N_1148,N_1173);
or U1270 (N_1270,N_1174,N_1161);
nand U1271 (N_1271,N_1162,N_1172);
nor U1272 (N_1272,N_1134,N_1127);
or U1273 (N_1273,N_1132,N_1127);
and U1274 (N_1274,N_1152,N_1141);
and U1275 (N_1275,N_1244,N_1240);
nor U1276 (N_1276,N_1253,N_1201);
xor U1277 (N_1277,N_1265,N_1207);
nor U1278 (N_1278,N_1269,N_1235);
nand U1279 (N_1279,N_1214,N_1210);
or U1280 (N_1280,N_1229,N_1247);
xor U1281 (N_1281,N_1254,N_1242);
and U1282 (N_1282,N_1205,N_1225);
or U1283 (N_1283,N_1211,N_1206);
nor U1284 (N_1284,N_1264,N_1262);
nand U1285 (N_1285,N_1250,N_1217);
and U1286 (N_1286,N_1237,N_1226);
or U1287 (N_1287,N_1227,N_1238);
or U1288 (N_1288,N_1223,N_1224);
and U1289 (N_1289,N_1215,N_1231);
or U1290 (N_1290,N_1246,N_1274);
xor U1291 (N_1291,N_1266,N_1252);
xor U1292 (N_1292,N_1261,N_1221);
xnor U1293 (N_1293,N_1267,N_1218);
or U1294 (N_1294,N_1204,N_1232);
or U1295 (N_1295,N_1257,N_1216);
nand U1296 (N_1296,N_1270,N_1222);
nor U1297 (N_1297,N_1236,N_1209);
or U1298 (N_1298,N_1251,N_1203);
and U1299 (N_1299,N_1202,N_1256);
nand U1300 (N_1300,N_1248,N_1272);
and U1301 (N_1301,N_1271,N_1273);
or U1302 (N_1302,N_1239,N_1255);
nand U1303 (N_1303,N_1233,N_1230);
or U1304 (N_1304,N_1234,N_1228);
and U1305 (N_1305,N_1213,N_1249);
or U1306 (N_1306,N_1200,N_1243);
nor U1307 (N_1307,N_1241,N_1219);
or U1308 (N_1308,N_1208,N_1212);
xor U1309 (N_1309,N_1263,N_1268);
nor U1310 (N_1310,N_1245,N_1260);
or U1311 (N_1311,N_1259,N_1220);
nand U1312 (N_1312,N_1258,N_1237);
nor U1313 (N_1313,N_1223,N_1221);
nor U1314 (N_1314,N_1203,N_1246);
and U1315 (N_1315,N_1239,N_1234);
or U1316 (N_1316,N_1220,N_1212);
xnor U1317 (N_1317,N_1252,N_1208);
and U1318 (N_1318,N_1205,N_1212);
nor U1319 (N_1319,N_1249,N_1264);
or U1320 (N_1320,N_1252,N_1214);
or U1321 (N_1321,N_1272,N_1268);
xor U1322 (N_1322,N_1249,N_1238);
xnor U1323 (N_1323,N_1271,N_1203);
nand U1324 (N_1324,N_1267,N_1269);
and U1325 (N_1325,N_1231,N_1211);
nand U1326 (N_1326,N_1227,N_1211);
xor U1327 (N_1327,N_1223,N_1237);
xor U1328 (N_1328,N_1258,N_1261);
xor U1329 (N_1329,N_1267,N_1237);
and U1330 (N_1330,N_1209,N_1264);
or U1331 (N_1331,N_1217,N_1269);
nand U1332 (N_1332,N_1263,N_1236);
nand U1333 (N_1333,N_1222,N_1261);
or U1334 (N_1334,N_1215,N_1230);
nor U1335 (N_1335,N_1226,N_1206);
and U1336 (N_1336,N_1257,N_1242);
nor U1337 (N_1337,N_1222,N_1211);
xnor U1338 (N_1338,N_1255,N_1209);
nand U1339 (N_1339,N_1223,N_1235);
xnor U1340 (N_1340,N_1268,N_1262);
and U1341 (N_1341,N_1239,N_1236);
nand U1342 (N_1342,N_1265,N_1200);
nor U1343 (N_1343,N_1257,N_1205);
xor U1344 (N_1344,N_1205,N_1230);
and U1345 (N_1345,N_1201,N_1213);
nand U1346 (N_1346,N_1269,N_1258);
nor U1347 (N_1347,N_1222,N_1212);
nor U1348 (N_1348,N_1232,N_1200);
nor U1349 (N_1349,N_1232,N_1254);
and U1350 (N_1350,N_1343,N_1318);
nand U1351 (N_1351,N_1319,N_1309);
nor U1352 (N_1352,N_1307,N_1349);
nor U1353 (N_1353,N_1288,N_1314);
nand U1354 (N_1354,N_1315,N_1303);
or U1355 (N_1355,N_1332,N_1345);
nor U1356 (N_1356,N_1334,N_1284);
xor U1357 (N_1357,N_1336,N_1338);
xor U1358 (N_1358,N_1297,N_1323);
xnor U1359 (N_1359,N_1298,N_1324);
nand U1360 (N_1360,N_1335,N_1312);
xnor U1361 (N_1361,N_1329,N_1278);
and U1362 (N_1362,N_1341,N_1296);
nand U1363 (N_1363,N_1282,N_1285);
nor U1364 (N_1364,N_1287,N_1333);
or U1365 (N_1365,N_1313,N_1299);
and U1366 (N_1366,N_1306,N_1283);
nand U1367 (N_1367,N_1280,N_1279);
nand U1368 (N_1368,N_1286,N_1328);
nor U1369 (N_1369,N_1305,N_1304);
nor U1370 (N_1370,N_1275,N_1325);
or U1371 (N_1371,N_1308,N_1301);
nor U1372 (N_1372,N_1326,N_1316);
nor U1373 (N_1373,N_1348,N_1346);
xnor U1374 (N_1374,N_1289,N_1320);
nor U1375 (N_1375,N_1292,N_1276);
xor U1376 (N_1376,N_1322,N_1337);
nor U1377 (N_1377,N_1331,N_1327);
nor U1378 (N_1378,N_1293,N_1347);
and U1379 (N_1379,N_1294,N_1290);
xnor U1380 (N_1380,N_1339,N_1321);
nand U1381 (N_1381,N_1340,N_1311);
nand U1382 (N_1382,N_1295,N_1291);
or U1383 (N_1383,N_1342,N_1317);
or U1384 (N_1384,N_1310,N_1344);
or U1385 (N_1385,N_1302,N_1281);
nand U1386 (N_1386,N_1277,N_1330);
nor U1387 (N_1387,N_1300,N_1283);
xnor U1388 (N_1388,N_1318,N_1284);
nor U1389 (N_1389,N_1301,N_1311);
nand U1390 (N_1390,N_1277,N_1279);
xnor U1391 (N_1391,N_1319,N_1303);
or U1392 (N_1392,N_1317,N_1322);
nand U1393 (N_1393,N_1281,N_1296);
nor U1394 (N_1394,N_1333,N_1343);
xor U1395 (N_1395,N_1294,N_1318);
nand U1396 (N_1396,N_1285,N_1278);
nor U1397 (N_1397,N_1347,N_1332);
nand U1398 (N_1398,N_1323,N_1349);
and U1399 (N_1399,N_1324,N_1287);
nor U1400 (N_1400,N_1325,N_1285);
nand U1401 (N_1401,N_1279,N_1337);
and U1402 (N_1402,N_1324,N_1348);
xnor U1403 (N_1403,N_1328,N_1284);
nor U1404 (N_1404,N_1292,N_1328);
nand U1405 (N_1405,N_1282,N_1349);
or U1406 (N_1406,N_1326,N_1305);
nand U1407 (N_1407,N_1301,N_1285);
nor U1408 (N_1408,N_1318,N_1289);
and U1409 (N_1409,N_1302,N_1311);
nor U1410 (N_1410,N_1291,N_1304);
or U1411 (N_1411,N_1327,N_1339);
xor U1412 (N_1412,N_1330,N_1303);
or U1413 (N_1413,N_1314,N_1301);
or U1414 (N_1414,N_1349,N_1299);
nand U1415 (N_1415,N_1284,N_1306);
nor U1416 (N_1416,N_1345,N_1314);
xnor U1417 (N_1417,N_1332,N_1338);
and U1418 (N_1418,N_1320,N_1279);
nand U1419 (N_1419,N_1300,N_1320);
and U1420 (N_1420,N_1348,N_1292);
xor U1421 (N_1421,N_1337,N_1346);
xor U1422 (N_1422,N_1307,N_1286);
nor U1423 (N_1423,N_1300,N_1278);
or U1424 (N_1424,N_1285,N_1284);
and U1425 (N_1425,N_1363,N_1394);
nand U1426 (N_1426,N_1388,N_1376);
xor U1427 (N_1427,N_1362,N_1351);
and U1428 (N_1428,N_1379,N_1371);
nand U1429 (N_1429,N_1421,N_1420);
nor U1430 (N_1430,N_1360,N_1359);
nor U1431 (N_1431,N_1410,N_1390);
xor U1432 (N_1432,N_1422,N_1424);
nand U1433 (N_1433,N_1405,N_1383);
nand U1434 (N_1434,N_1396,N_1366);
nand U1435 (N_1435,N_1361,N_1423);
or U1436 (N_1436,N_1406,N_1399);
xnor U1437 (N_1437,N_1404,N_1403);
and U1438 (N_1438,N_1380,N_1395);
and U1439 (N_1439,N_1386,N_1353);
or U1440 (N_1440,N_1417,N_1365);
nand U1441 (N_1441,N_1384,N_1387);
or U1442 (N_1442,N_1382,N_1389);
nand U1443 (N_1443,N_1357,N_1354);
and U1444 (N_1444,N_1375,N_1358);
nor U1445 (N_1445,N_1377,N_1393);
nor U1446 (N_1446,N_1378,N_1415);
nand U1447 (N_1447,N_1397,N_1402);
nor U1448 (N_1448,N_1364,N_1352);
nor U1449 (N_1449,N_1408,N_1416);
nand U1450 (N_1450,N_1414,N_1381);
nor U1451 (N_1451,N_1385,N_1391);
or U1452 (N_1452,N_1373,N_1392);
xor U1453 (N_1453,N_1368,N_1401);
xor U1454 (N_1454,N_1374,N_1398);
nor U1455 (N_1455,N_1413,N_1356);
and U1456 (N_1456,N_1372,N_1419);
nor U1457 (N_1457,N_1409,N_1411);
nor U1458 (N_1458,N_1350,N_1412);
or U1459 (N_1459,N_1418,N_1400);
nand U1460 (N_1460,N_1407,N_1355);
nand U1461 (N_1461,N_1367,N_1370);
and U1462 (N_1462,N_1369,N_1373);
and U1463 (N_1463,N_1354,N_1401);
and U1464 (N_1464,N_1415,N_1396);
nand U1465 (N_1465,N_1392,N_1396);
xor U1466 (N_1466,N_1413,N_1353);
and U1467 (N_1467,N_1377,N_1422);
or U1468 (N_1468,N_1418,N_1382);
nor U1469 (N_1469,N_1414,N_1393);
xor U1470 (N_1470,N_1383,N_1361);
and U1471 (N_1471,N_1384,N_1352);
xor U1472 (N_1472,N_1359,N_1355);
nand U1473 (N_1473,N_1387,N_1405);
nand U1474 (N_1474,N_1353,N_1400);
or U1475 (N_1475,N_1357,N_1403);
and U1476 (N_1476,N_1407,N_1399);
nor U1477 (N_1477,N_1389,N_1358);
and U1478 (N_1478,N_1404,N_1390);
and U1479 (N_1479,N_1376,N_1422);
or U1480 (N_1480,N_1370,N_1361);
and U1481 (N_1481,N_1369,N_1354);
or U1482 (N_1482,N_1353,N_1420);
nor U1483 (N_1483,N_1351,N_1400);
or U1484 (N_1484,N_1355,N_1396);
or U1485 (N_1485,N_1419,N_1353);
or U1486 (N_1486,N_1361,N_1419);
or U1487 (N_1487,N_1404,N_1353);
nor U1488 (N_1488,N_1376,N_1350);
xnor U1489 (N_1489,N_1381,N_1396);
and U1490 (N_1490,N_1402,N_1351);
xor U1491 (N_1491,N_1421,N_1385);
xnor U1492 (N_1492,N_1418,N_1380);
or U1493 (N_1493,N_1351,N_1396);
and U1494 (N_1494,N_1419,N_1374);
or U1495 (N_1495,N_1387,N_1367);
nand U1496 (N_1496,N_1362,N_1353);
nor U1497 (N_1497,N_1382,N_1353);
nand U1498 (N_1498,N_1416,N_1360);
nor U1499 (N_1499,N_1402,N_1396);
xor U1500 (N_1500,N_1457,N_1461);
xnor U1501 (N_1501,N_1471,N_1466);
and U1502 (N_1502,N_1463,N_1432);
nor U1503 (N_1503,N_1486,N_1438);
and U1504 (N_1504,N_1441,N_1468);
nor U1505 (N_1505,N_1488,N_1456);
nor U1506 (N_1506,N_1450,N_1433);
nor U1507 (N_1507,N_1439,N_1453);
or U1508 (N_1508,N_1491,N_1490);
nand U1509 (N_1509,N_1464,N_1426);
nor U1510 (N_1510,N_1469,N_1448);
nand U1511 (N_1511,N_1436,N_1492);
or U1512 (N_1512,N_1489,N_1454);
nand U1513 (N_1513,N_1444,N_1427);
nor U1514 (N_1514,N_1478,N_1482);
nand U1515 (N_1515,N_1440,N_1496);
nor U1516 (N_1516,N_1449,N_1497);
and U1517 (N_1517,N_1475,N_1460);
or U1518 (N_1518,N_1446,N_1465);
nor U1519 (N_1519,N_1498,N_1476);
xnor U1520 (N_1520,N_1472,N_1442);
nand U1521 (N_1521,N_1479,N_1458);
and U1522 (N_1522,N_1451,N_1455);
and U1523 (N_1523,N_1470,N_1477);
nand U1524 (N_1524,N_1452,N_1462);
nor U1525 (N_1525,N_1493,N_1487);
or U1526 (N_1526,N_1480,N_1459);
nand U1527 (N_1527,N_1483,N_1429);
nor U1528 (N_1528,N_1428,N_1474);
xor U1529 (N_1529,N_1445,N_1499);
nor U1530 (N_1530,N_1481,N_1473);
nor U1531 (N_1531,N_1485,N_1484);
nor U1532 (N_1532,N_1425,N_1447);
and U1533 (N_1533,N_1430,N_1494);
xor U1534 (N_1534,N_1443,N_1495);
xnor U1535 (N_1535,N_1437,N_1434);
or U1536 (N_1536,N_1435,N_1431);
nand U1537 (N_1537,N_1467,N_1450);
or U1538 (N_1538,N_1483,N_1425);
nand U1539 (N_1539,N_1443,N_1493);
nand U1540 (N_1540,N_1493,N_1485);
xor U1541 (N_1541,N_1431,N_1491);
xor U1542 (N_1542,N_1437,N_1475);
xor U1543 (N_1543,N_1485,N_1433);
and U1544 (N_1544,N_1466,N_1458);
nor U1545 (N_1545,N_1438,N_1443);
nor U1546 (N_1546,N_1474,N_1445);
or U1547 (N_1547,N_1464,N_1436);
and U1548 (N_1548,N_1429,N_1450);
xor U1549 (N_1549,N_1444,N_1494);
or U1550 (N_1550,N_1432,N_1477);
nor U1551 (N_1551,N_1427,N_1431);
and U1552 (N_1552,N_1496,N_1485);
and U1553 (N_1553,N_1483,N_1433);
nor U1554 (N_1554,N_1454,N_1466);
or U1555 (N_1555,N_1485,N_1439);
nor U1556 (N_1556,N_1444,N_1476);
or U1557 (N_1557,N_1442,N_1459);
nand U1558 (N_1558,N_1453,N_1488);
nor U1559 (N_1559,N_1478,N_1499);
or U1560 (N_1560,N_1429,N_1497);
xor U1561 (N_1561,N_1469,N_1499);
nand U1562 (N_1562,N_1475,N_1447);
nor U1563 (N_1563,N_1486,N_1487);
or U1564 (N_1564,N_1474,N_1473);
or U1565 (N_1565,N_1452,N_1433);
and U1566 (N_1566,N_1480,N_1448);
nor U1567 (N_1567,N_1486,N_1451);
nand U1568 (N_1568,N_1463,N_1446);
nor U1569 (N_1569,N_1451,N_1468);
and U1570 (N_1570,N_1447,N_1429);
xor U1571 (N_1571,N_1431,N_1488);
or U1572 (N_1572,N_1487,N_1474);
nand U1573 (N_1573,N_1494,N_1485);
nor U1574 (N_1574,N_1482,N_1441);
nor U1575 (N_1575,N_1570,N_1523);
nand U1576 (N_1576,N_1541,N_1514);
nor U1577 (N_1577,N_1572,N_1567);
xnor U1578 (N_1578,N_1560,N_1528);
xor U1579 (N_1579,N_1546,N_1561);
or U1580 (N_1580,N_1535,N_1529);
xnor U1581 (N_1581,N_1538,N_1516);
nand U1582 (N_1582,N_1566,N_1506);
and U1583 (N_1583,N_1512,N_1547);
nor U1584 (N_1584,N_1574,N_1507);
and U1585 (N_1585,N_1534,N_1532);
nand U1586 (N_1586,N_1510,N_1520);
xnor U1587 (N_1587,N_1509,N_1525);
nand U1588 (N_1588,N_1521,N_1563);
nor U1589 (N_1589,N_1530,N_1522);
nor U1590 (N_1590,N_1504,N_1519);
and U1591 (N_1591,N_1501,N_1517);
nand U1592 (N_1592,N_1524,N_1550);
or U1593 (N_1593,N_1539,N_1537);
nand U1594 (N_1594,N_1559,N_1518);
or U1595 (N_1595,N_1531,N_1556);
xnor U1596 (N_1596,N_1571,N_1549);
xor U1597 (N_1597,N_1573,N_1543);
xnor U1598 (N_1598,N_1554,N_1500);
or U1599 (N_1599,N_1533,N_1515);
nor U1600 (N_1600,N_1568,N_1569);
nor U1601 (N_1601,N_1536,N_1548);
nor U1602 (N_1602,N_1526,N_1565);
xor U1603 (N_1603,N_1558,N_1557);
or U1604 (N_1604,N_1540,N_1542);
and U1605 (N_1605,N_1552,N_1555);
nand U1606 (N_1606,N_1562,N_1527);
and U1607 (N_1607,N_1545,N_1564);
nor U1608 (N_1608,N_1553,N_1551);
nand U1609 (N_1609,N_1544,N_1505);
nor U1610 (N_1610,N_1511,N_1502);
nand U1611 (N_1611,N_1503,N_1513);
nand U1612 (N_1612,N_1508,N_1530);
and U1613 (N_1613,N_1569,N_1541);
or U1614 (N_1614,N_1572,N_1547);
nand U1615 (N_1615,N_1559,N_1545);
nor U1616 (N_1616,N_1554,N_1533);
and U1617 (N_1617,N_1520,N_1535);
xor U1618 (N_1618,N_1531,N_1508);
and U1619 (N_1619,N_1567,N_1530);
nor U1620 (N_1620,N_1528,N_1557);
nor U1621 (N_1621,N_1523,N_1565);
nand U1622 (N_1622,N_1504,N_1536);
nand U1623 (N_1623,N_1551,N_1527);
nor U1624 (N_1624,N_1522,N_1525);
nand U1625 (N_1625,N_1545,N_1512);
xnor U1626 (N_1626,N_1541,N_1540);
nand U1627 (N_1627,N_1534,N_1528);
xnor U1628 (N_1628,N_1535,N_1574);
or U1629 (N_1629,N_1528,N_1521);
nor U1630 (N_1630,N_1510,N_1543);
and U1631 (N_1631,N_1539,N_1564);
nor U1632 (N_1632,N_1567,N_1562);
nor U1633 (N_1633,N_1555,N_1563);
xor U1634 (N_1634,N_1563,N_1562);
or U1635 (N_1635,N_1573,N_1512);
and U1636 (N_1636,N_1554,N_1560);
nor U1637 (N_1637,N_1532,N_1509);
xnor U1638 (N_1638,N_1573,N_1513);
nand U1639 (N_1639,N_1510,N_1548);
and U1640 (N_1640,N_1564,N_1527);
or U1641 (N_1641,N_1516,N_1530);
xor U1642 (N_1642,N_1570,N_1525);
or U1643 (N_1643,N_1510,N_1567);
xnor U1644 (N_1644,N_1547,N_1522);
nor U1645 (N_1645,N_1537,N_1540);
nor U1646 (N_1646,N_1504,N_1547);
nor U1647 (N_1647,N_1530,N_1566);
nand U1648 (N_1648,N_1546,N_1556);
nand U1649 (N_1649,N_1510,N_1530);
nor U1650 (N_1650,N_1633,N_1608);
xnor U1651 (N_1651,N_1629,N_1638);
and U1652 (N_1652,N_1601,N_1634);
nand U1653 (N_1653,N_1576,N_1612);
or U1654 (N_1654,N_1585,N_1609);
nor U1655 (N_1655,N_1588,N_1625);
or U1656 (N_1656,N_1610,N_1647);
xnor U1657 (N_1657,N_1595,N_1578);
nand U1658 (N_1658,N_1600,N_1641);
or U1659 (N_1659,N_1620,N_1632);
nor U1660 (N_1660,N_1596,N_1648);
xor U1661 (N_1661,N_1624,N_1640);
and U1662 (N_1662,N_1618,N_1605);
nor U1663 (N_1663,N_1619,N_1590);
and U1664 (N_1664,N_1603,N_1644);
nor U1665 (N_1665,N_1615,N_1611);
nand U1666 (N_1666,N_1622,N_1623);
xor U1667 (N_1667,N_1582,N_1583);
and U1668 (N_1668,N_1616,N_1602);
xor U1669 (N_1669,N_1581,N_1599);
and U1670 (N_1670,N_1630,N_1598);
xor U1671 (N_1671,N_1580,N_1642);
nand U1672 (N_1672,N_1607,N_1575);
and U1673 (N_1673,N_1646,N_1639);
or U1674 (N_1674,N_1636,N_1617);
xor U1675 (N_1675,N_1613,N_1591);
or U1676 (N_1676,N_1645,N_1589);
and U1677 (N_1677,N_1628,N_1597);
nor U1678 (N_1678,N_1592,N_1631);
and U1679 (N_1679,N_1621,N_1635);
and U1680 (N_1680,N_1649,N_1586);
or U1681 (N_1681,N_1584,N_1604);
xor U1682 (N_1682,N_1643,N_1627);
nand U1683 (N_1683,N_1637,N_1587);
xnor U1684 (N_1684,N_1626,N_1594);
or U1685 (N_1685,N_1614,N_1593);
xor U1686 (N_1686,N_1579,N_1577);
xnor U1687 (N_1687,N_1606,N_1575);
xnor U1688 (N_1688,N_1647,N_1586);
xor U1689 (N_1689,N_1614,N_1637);
and U1690 (N_1690,N_1648,N_1594);
and U1691 (N_1691,N_1591,N_1639);
xor U1692 (N_1692,N_1635,N_1576);
nor U1693 (N_1693,N_1648,N_1643);
nand U1694 (N_1694,N_1645,N_1598);
or U1695 (N_1695,N_1630,N_1595);
and U1696 (N_1696,N_1626,N_1577);
or U1697 (N_1697,N_1635,N_1619);
or U1698 (N_1698,N_1646,N_1624);
and U1699 (N_1699,N_1625,N_1617);
nand U1700 (N_1700,N_1640,N_1637);
or U1701 (N_1701,N_1641,N_1635);
or U1702 (N_1702,N_1629,N_1582);
nor U1703 (N_1703,N_1645,N_1637);
nand U1704 (N_1704,N_1589,N_1631);
nand U1705 (N_1705,N_1627,N_1585);
nand U1706 (N_1706,N_1610,N_1603);
and U1707 (N_1707,N_1616,N_1631);
xnor U1708 (N_1708,N_1599,N_1643);
nor U1709 (N_1709,N_1575,N_1586);
nor U1710 (N_1710,N_1616,N_1642);
nor U1711 (N_1711,N_1587,N_1576);
xnor U1712 (N_1712,N_1635,N_1605);
nor U1713 (N_1713,N_1616,N_1618);
and U1714 (N_1714,N_1598,N_1624);
nor U1715 (N_1715,N_1576,N_1596);
nand U1716 (N_1716,N_1627,N_1587);
nor U1717 (N_1717,N_1606,N_1611);
xnor U1718 (N_1718,N_1622,N_1633);
and U1719 (N_1719,N_1612,N_1577);
or U1720 (N_1720,N_1622,N_1585);
and U1721 (N_1721,N_1598,N_1593);
nor U1722 (N_1722,N_1604,N_1613);
and U1723 (N_1723,N_1608,N_1628);
and U1724 (N_1724,N_1577,N_1596);
or U1725 (N_1725,N_1718,N_1703);
and U1726 (N_1726,N_1660,N_1657);
or U1727 (N_1727,N_1673,N_1669);
nand U1728 (N_1728,N_1721,N_1711);
nor U1729 (N_1729,N_1707,N_1663);
nand U1730 (N_1730,N_1719,N_1700);
and U1731 (N_1731,N_1690,N_1691);
or U1732 (N_1732,N_1668,N_1684);
xor U1733 (N_1733,N_1723,N_1708);
and U1734 (N_1734,N_1722,N_1683);
and U1735 (N_1735,N_1677,N_1680);
or U1736 (N_1736,N_1685,N_1658);
nor U1737 (N_1737,N_1714,N_1713);
and U1738 (N_1738,N_1654,N_1662);
and U1739 (N_1739,N_1667,N_1653);
or U1740 (N_1740,N_1715,N_1720);
or U1741 (N_1741,N_1698,N_1717);
nand U1742 (N_1742,N_1687,N_1659);
or U1743 (N_1743,N_1699,N_1692);
xnor U1744 (N_1744,N_1702,N_1665);
xnor U1745 (N_1745,N_1693,N_1696);
or U1746 (N_1746,N_1678,N_1670);
nand U1747 (N_1747,N_1712,N_1666);
nor U1748 (N_1748,N_1686,N_1697);
nor U1749 (N_1749,N_1672,N_1689);
or U1750 (N_1750,N_1709,N_1650);
nand U1751 (N_1751,N_1704,N_1655);
and U1752 (N_1752,N_1675,N_1701);
or U1753 (N_1753,N_1674,N_1671);
or U1754 (N_1754,N_1694,N_1651);
nand U1755 (N_1755,N_1652,N_1664);
xnor U1756 (N_1756,N_1676,N_1679);
nor U1757 (N_1757,N_1710,N_1688);
or U1758 (N_1758,N_1695,N_1705);
nor U1759 (N_1759,N_1682,N_1724);
nand U1760 (N_1760,N_1716,N_1681);
or U1761 (N_1761,N_1706,N_1661);
and U1762 (N_1762,N_1656,N_1682);
or U1763 (N_1763,N_1672,N_1652);
xor U1764 (N_1764,N_1675,N_1650);
nand U1765 (N_1765,N_1724,N_1676);
and U1766 (N_1766,N_1718,N_1683);
nand U1767 (N_1767,N_1680,N_1717);
nor U1768 (N_1768,N_1696,N_1718);
xnor U1769 (N_1769,N_1663,N_1661);
or U1770 (N_1770,N_1656,N_1678);
and U1771 (N_1771,N_1694,N_1715);
nand U1772 (N_1772,N_1702,N_1656);
nand U1773 (N_1773,N_1682,N_1702);
xor U1774 (N_1774,N_1683,N_1673);
xnor U1775 (N_1775,N_1711,N_1679);
or U1776 (N_1776,N_1677,N_1675);
or U1777 (N_1777,N_1651,N_1722);
nand U1778 (N_1778,N_1671,N_1703);
nand U1779 (N_1779,N_1679,N_1667);
or U1780 (N_1780,N_1659,N_1702);
and U1781 (N_1781,N_1665,N_1685);
xor U1782 (N_1782,N_1668,N_1698);
nand U1783 (N_1783,N_1703,N_1657);
xor U1784 (N_1784,N_1699,N_1650);
nor U1785 (N_1785,N_1680,N_1660);
nor U1786 (N_1786,N_1692,N_1711);
xor U1787 (N_1787,N_1661,N_1698);
or U1788 (N_1788,N_1655,N_1685);
or U1789 (N_1789,N_1709,N_1693);
and U1790 (N_1790,N_1705,N_1693);
nand U1791 (N_1791,N_1690,N_1689);
nand U1792 (N_1792,N_1706,N_1705);
xor U1793 (N_1793,N_1723,N_1670);
nor U1794 (N_1794,N_1721,N_1653);
or U1795 (N_1795,N_1677,N_1664);
nand U1796 (N_1796,N_1661,N_1688);
and U1797 (N_1797,N_1663,N_1660);
nand U1798 (N_1798,N_1717,N_1694);
nor U1799 (N_1799,N_1691,N_1721);
nor U1800 (N_1800,N_1731,N_1792);
xor U1801 (N_1801,N_1743,N_1756);
nand U1802 (N_1802,N_1775,N_1746);
nand U1803 (N_1803,N_1755,N_1725);
nor U1804 (N_1804,N_1789,N_1738);
xor U1805 (N_1805,N_1773,N_1765);
and U1806 (N_1806,N_1770,N_1768);
nand U1807 (N_1807,N_1788,N_1794);
or U1808 (N_1808,N_1739,N_1733);
and U1809 (N_1809,N_1757,N_1769);
nor U1810 (N_1810,N_1730,N_1778);
nand U1811 (N_1811,N_1750,N_1786);
xnor U1812 (N_1812,N_1798,N_1785);
nor U1813 (N_1813,N_1780,N_1774);
nor U1814 (N_1814,N_1781,N_1753);
and U1815 (N_1815,N_1763,N_1735);
nor U1816 (N_1816,N_1751,N_1741);
and U1817 (N_1817,N_1759,N_1787);
or U1818 (N_1818,N_1777,N_1727);
nor U1819 (N_1819,N_1734,N_1793);
and U1820 (N_1820,N_1767,N_1799);
and U1821 (N_1821,N_1779,N_1762);
and U1822 (N_1822,N_1782,N_1776);
nor U1823 (N_1823,N_1795,N_1796);
or U1824 (N_1824,N_1732,N_1771);
nor U1825 (N_1825,N_1784,N_1740);
or U1826 (N_1826,N_1748,N_1744);
nand U1827 (N_1827,N_1760,N_1772);
nand U1828 (N_1828,N_1752,N_1754);
xor U1829 (N_1829,N_1758,N_1726);
nor U1830 (N_1830,N_1749,N_1747);
xnor U1831 (N_1831,N_1742,N_1764);
and U1832 (N_1832,N_1790,N_1766);
and U1833 (N_1833,N_1737,N_1745);
or U1834 (N_1834,N_1797,N_1791);
xnor U1835 (N_1835,N_1736,N_1783);
nor U1836 (N_1836,N_1728,N_1729);
nor U1837 (N_1837,N_1761,N_1784);
xor U1838 (N_1838,N_1734,N_1781);
and U1839 (N_1839,N_1768,N_1734);
or U1840 (N_1840,N_1794,N_1795);
nand U1841 (N_1841,N_1779,N_1748);
and U1842 (N_1842,N_1784,N_1730);
and U1843 (N_1843,N_1756,N_1764);
xor U1844 (N_1844,N_1778,N_1776);
xor U1845 (N_1845,N_1734,N_1787);
nand U1846 (N_1846,N_1776,N_1793);
nor U1847 (N_1847,N_1765,N_1753);
and U1848 (N_1848,N_1778,N_1742);
nor U1849 (N_1849,N_1779,N_1731);
nor U1850 (N_1850,N_1796,N_1750);
nand U1851 (N_1851,N_1735,N_1771);
nor U1852 (N_1852,N_1775,N_1776);
nor U1853 (N_1853,N_1769,N_1755);
xnor U1854 (N_1854,N_1750,N_1751);
xnor U1855 (N_1855,N_1771,N_1729);
nor U1856 (N_1856,N_1786,N_1736);
or U1857 (N_1857,N_1788,N_1783);
nand U1858 (N_1858,N_1747,N_1773);
nor U1859 (N_1859,N_1794,N_1744);
nand U1860 (N_1860,N_1728,N_1797);
and U1861 (N_1861,N_1741,N_1775);
and U1862 (N_1862,N_1786,N_1789);
xnor U1863 (N_1863,N_1760,N_1762);
and U1864 (N_1864,N_1751,N_1767);
and U1865 (N_1865,N_1742,N_1739);
xnor U1866 (N_1866,N_1730,N_1762);
or U1867 (N_1867,N_1736,N_1753);
xnor U1868 (N_1868,N_1739,N_1762);
nand U1869 (N_1869,N_1799,N_1749);
or U1870 (N_1870,N_1786,N_1740);
nand U1871 (N_1871,N_1730,N_1785);
nor U1872 (N_1872,N_1748,N_1784);
nor U1873 (N_1873,N_1796,N_1778);
or U1874 (N_1874,N_1760,N_1780);
and U1875 (N_1875,N_1823,N_1816);
nand U1876 (N_1876,N_1862,N_1810);
nor U1877 (N_1877,N_1855,N_1827);
and U1878 (N_1878,N_1806,N_1836);
or U1879 (N_1879,N_1824,N_1852);
nor U1880 (N_1880,N_1844,N_1809);
and U1881 (N_1881,N_1856,N_1868);
xnor U1882 (N_1882,N_1814,N_1858);
nor U1883 (N_1883,N_1839,N_1849);
nor U1884 (N_1884,N_1859,N_1861);
and U1885 (N_1885,N_1831,N_1867);
xor U1886 (N_1886,N_1845,N_1802);
and U1887 (N_1887,N_1846,N_1818);
and U1888 (N_1888,N_1820,N_1874);
and U1889 (N_1889,N_1860,N_1826);
nor U1890 (N_1890,N_1869,N_1822);
or U1891 (N_1891,N_1870,N_1837);
nand U1892 (N_1892,N_1873,N_1804);
nor U1893 (N_1893,N_1847,N_1813);
nor U1894 (N_1894,N_1865,N_1834);
nor U1895 (N_1895,N_1812,N_1841);
nand U1896 (N_1896,N_1808,N_1807);
and U1897 (N_1897,N_1821,N_1840);
or U1898 (N_1898,N_1842,N_1825);
nand U1899 (N_1899,N_1829,N_1848);
or U1900 (N_1900,N_1835,N_1800);
nor U1901 (N_1901,N_1830,N_1828);
nand U1902 (N_1902,N_1871,N_1817);
and U1903 (N_1903,N_1872,N_1811);
nand U1904 (N_1904,N_1833,N_1801);
xnor U1905 (N_1905,N_1857,N_1864);
and U1906 (N_1906,N_1832,N_1843);
nor U1907 (N_1907,N_1863,N_1866);
xor U1908 (N_1908,N_1803,N_1854);
and U1909 (N_1909,N_1805,N_1853);
nor U1910 (N_1910,N_1819,N_1850);
xnor U1911 (N_1911,N_1815,N_1851);
nor U1912 (N_1912,N_1838,N_1820);
nand U1913 (N_1913,N_1835,N_1864);
and U1914 (N_1914,N_1848,N_1806);
or U1915 (N_1915,N_1825,N_1815);
or U1916 (N_1916,N_1849,N_1834);
nand U1917 (N_1917,N_1810,N_1822);
xor U1918 (N_1918,N_1808,N_1833);
and U1919 (N_1919,N_1825,N_1810);
or U1920 (N_1920,N_1849,N_1853);
nand U1921 (N_1921,N_1838,N_1868);
xor U1922 (N_1922,N_1854,N_1872);
and U1923 (N_1923,N_1847,N_1800);
nor U1924 (N_1924,N_1873,N_1815);
or U1925 (N_1925,N_1840,N_1817);
or U1926 (N_1926,N_1867,N_1806);
and U1927 (N_1927,N_1805,N_1838);
nand U1928 (N_1928,N_1831,N_1870);
nor U1929 (N_1929,N_1829,N_1826);
nor U1930 (N_1930,N_1863,N_1801);
nor U1931 (N_1931,N_1853,N_1823);
nand U1932 (N_1932,N_1808,N_1801);
and U1933 (N_1933,N_1851,N_1812);
or U1934 (N_1934,N_1861,N_1801);
nor U1935 (N_1935,N_1820,N_1823);
xnor U1936 (N_1936,N_1846,N_1813);
and U1937 (N_1937,N_1830,N_1858);
nor U1938 (N_1938,N_1844,N_1870);
xor U1939 (N_1939,N_1814,N_1846);
or U1940 (N_1940,N_1805,N_1832);
nand U1941 (N_1941,N_1816,N_1804);
and U1942 (N_1942,N_1860,N_1853);
and U1943 (N_1943,N_1815,N_1871);
nor U1944 (N_1944,N_1842,N_1839);
nand U1945 (N_1945,N_1800,N_1801);
nand U1946 (N_1946,N_1850,N_1840);
and U1947 (N_1947,N_1852,N_1820);
and U1948 (N_1948,N_1846,N_1802);
or U1949 (N_1949,N_1833,N_1873);
or U1950 (N_1950,N_1926,N_1883);
or U1951 (N_1951,N_1875,N_1927);
nand U1952 (N_1952,N_1943,N_1907);
xor U1953 (N_1953,N_1880,N_1918);
or U1954 (N_1954,N_1902,N_1888);
xor U1955 (N_1955,N_1947,N_1936);
xnor U1956 (N_1956,N_1884,N_1895);
nand U1957 (N_1957,N_1900,N_1901);
xor U1958 (N_1958,N_1920,N_1881);
xor U1959 (N_1959,N_1882,N_1941);
and U1960 (N_1960,N_1878,N_1885);
or U1961 (N_1961,N_1929,N_1897);
and U1962 (N_1962,N_1937,N_1891);
nand U1963 (N_1963,N_1908,N_1894);
xnor U1964 (N_1964,N_1924,N_1914);
or U1965 (N_1965,N_1903,N_1949);
and U1966 (N_1966,N_1917,N_1877);
nor U1967 (N_1967,N_1879,N_1913);
nor U1968 (N_1968,N_1942,N_1889);
and U1969 (N_1969,N_1923,N_1928);
nand U1970 (N_1970,N_1898,N_1915);
nor U1971 (N_1971,N_1919,N_1945);
xor U1972 (N_1972,N_1899,N_1909);
nor U1973 (N_1973,N_1916,N_1896);
and U1974 (N_1974,N_1935,N_1876);
and U1975 (N_1975,N_1905,N_1946);
and U1976 (N_1976,N_1886,N_1948);
nor U1977 (N_1977,N_1910,N_1890);
xor U1978 (N_1978,N_1922,N_1939);
nor U1979 (N_1979,N_1912,N_1931);
xnor U1980 (N_1980,N_1940,N_1932);
nand U1981 (N_1981,N_1925,N_1893);
nor U1982 (N_1982,N_1944,N_1938);
xnor U1983 (N_1983,N_1887,N_1906);
and U1984 (N_1984,N_1933,N_1904);
or U1985 (N_1985,N_1934,N_1911);
nand U1986 (N_1986,N_1892,N_1921);
or U1987 (N_1987,N_1930,N_1927);
nand U1988 (N_1988,N_1929,N_1895);
nor U1989 (N_1989,N_1894,N_1902);
and U1990 (N_1990,N_1890,N_1881);
xor U1991 (N_1991,N_1944,N_1919);
xnor U1992 (N_1992,N_1942,N_1894);
nor U1993 (N_1993,N_1880,N_1942);
nor U1994 (N_1994,N_1921,N_1879);
nor U1995 (N_1995,N_1914,N_1902);
nand U1996 (N_1996,N_1891,N_1949);
nand U1997 (N_1997,N_1941,N_1935);
nand U1998 (N_1998,N_1905,N_1942);
nor U1999 (N_1999,N_1945,N_1914);
nand U2000 (N_2000,N_1940,N_1912);
xnor U2001 (N_2001,N_1923,N_1892);
xor U2002 (N_2002,N_1909,N_1923);
and U2003 (N_2003,N_1949,N_1900);
nand U2004 (N_2004,N_1906,N_1930);
nor U2005 (N_2005,N_1880,N_1945);
xor U2006 (N_2006,N_1900,N_1928);
nand U2007 (N_2007,N_1913,N_1937);
xnor U2008 (N_2008,N_1884,N_1901);
xor U2009 (N_2009,N_1903,N_1889);
xnor U2010 (N_2010,N_1913,N_1938);
or U2011 (N_2011,N_1939,N_1900);
or U2012 (N_2012,N_1932,N_1889);
and U2013 (N_2013,N_1943,N_1893);
and U2014 (N_2014,N_1917,N_1928);
and U2015 (N_2015,N_1931,N_1884);
nor U2016 (N_2016,N_1920,N_1890);
and U2017 (N_2017,N_1878,N_1935);
nand U2018 (N_2018,N_1880,N_1883);
and U2019 (N_2019,N_1936,N_1902);
xor U2020 (N_2020,N_1877,N_1919);
and U2021 (N_2021,N_1935,N_1891);
or U2022 (N_2022,N_1928,N_1913);
nand U2023 (N_2023,N_1886,N_1879);
or U2024 (N_2024,N_1901,N_1904);
and U2025 (N_2025,N_1998,N_1991);
nor U2026 (N_2026,N_2018,N_1955);
nand U2027 (N_2027,N_1957,N_2015);
nand U2028 (N_2028,N_1983,N_1990);
or U2029 (N_2029,N_1986,N_1968);
xor U2030 (N_2030,N_2016,N_1994);
nand U2031 (N_2031,N_1976,N_1958);
xor U2032 (N_2032,N_1964,N_2011);
or U2033 (N_2033,N_2006,N_2010);
and U2034 (N_2034,N_2023,N_1977);
nor U2035 (N_2035,N_2000,N_1979);
xnor U2036 (N_2036,N_2017,N_1971);
nand U2037 (N_2037,N_2022,N_1973);
nand U2038 (N_2038,N_1969,N_1975);
and U2039 (N_2039,N_1972,N_1995);
and U2040 (N_2040,N_1989,N_1988);
and U2041 (N_2041,N_2019,N_1993);
nand U2042 (N_2042,N_1956,N_1961);
xor U2043 (N_2043,N_1987,N_1952);
nand U2044 (N_2044,N_1951,N_1965);
or U2045 (N_2045,N_2005,N_1950);
and U2046 (N_2046,N_1984,N_1963);
nor U2047 (N_2047,N_1997,N_1970);
or U2048 (N_2048,N_1999,N_2013);
or U2049 (N_2049,N_1974,N_2014);
and U2050 (N_2050,N_1966,N_1996);
nand U2051 (N_2051,N_2020,N_2009);
or U2052 (N_2052,N_2007,N_1982);
and U2053 (N_2053,N_2024,N_1985);
or U2054 (N_2054,N_1992,N_2008);
nor U2055 (N_2055,N_1953,N_2004);
and U2056 (N_2056,N_1962,N_1981);
and U2057 (N_2057,N_2001,N_1978);
and U2058 (N_2058,N_1967,N_1960);
nor U2059 (N_2059,N_2003,N_2012);
or U2060 (N_2060,N_1954,N_1959);
and U2061 (N_2061,N_2002,N_1980);
and U2062 (N_2062,N_2021,N_1995);
xnor U2063 (N_2063,N_1975,N_1968);
and U2064 (N_2064,N_1967,N_2008);
nand U2065 (N_2065,N_1977,N_1992);
nand U2066 (N_2066,N_1979,N_1955);
nor U2067 (N_2067,N_1990,N_1968);
nor U2068 (N_2068,N_1987,N_1988);
xor U2069 (N_2069,N_2017,N_1954);
and U2070 (N_2070,N_1975,N_2019);
or U2071 (N_2071,N_2020,N_1954);
or U2072 (N_2072,N_1968,N_1977);
or U2073 (N_2073,N_2002,N_2018);
xnor U2074 (N_2074,N_2005,N_1993);
xnor U2075 (N_2075,N_2006,N_1979);
or U2076 (N_2076,N_2002,N_2023);
xnor U2077 (N_2077,N_2008,N_1989);
nand U2078 (N_2078,N_2017,N_2009);
or U2079 (N_2079,N_1982,N_1988);
nor U2080 (N_2080,N_1950,N_1993);
xor U2081 (N_2081,N_2001,N_1986);
and U2082 (N_2082,N_1985,N_1950);
nor U2083 (N_2083,N_1966,N_2015);
nand U2084 (N_2084,N_1986,N_2004);
and U2085 (N_2085,N_1981,N_1953);
or U2086 (N_2086,N_1952,N_1984);
and U2087 (N_2087,N_1975,N_1966);
nand U2088 (N_2088,N_1982,N_2004);
nor U2089 (N_2089,N_2000,N_1969);
or U2090 (N_2090,N_2023,N_2019);
or U2091 (N_2091,N_1984,N_1961);
or U2092 (N_2092,N_2010,N_2011);
nor U2093 (N_2093,N_1962,N_2005);
nor U2094 (N_2094,N_1996,N_1956);
or U2095 (N_2095,N_1958,N_1970);
or U2096 (N_2096,N_2003,N_1987);
nand U2097 (N_2097,N_1967,N_1954);
or U2098 (N_2098,N_1954,N_2021);
xnor U2099 (N_2099,N_2013,N_1990);
nor U2100 (N_2100,N_2068,N_2035);
xor U2101 (N_2101,N_2055,N_2037);
nor U2102 (N_2102,N_2044,N_2047);
nand U2103 (N_2103,N_2065,N_2071);
nor U2104 (N_2104,N_2030,N_2069);
nor U2105 (N_2105,N_2045,N_2040);
nand U2106 (N_2106,N_2082,N_2064);
or U2107 (N_2107,N_2085,N_2076);
nor U2108 (N_2108,N_2051,N_2089);
or U2109 (N_2109,N_2078,N_2099);
nor U2110 (N_2110,N_2087,N_2039);
nand U2111 (N_2111,N_2097,N_2056);
nor U2112 (N_2112,N_2077,N_2095);
and U2113 (N_2113,N_2049,N_2038);
or U2114 (N_2114,N_2062,N_2098);
nor U2115 (N_2115,N_2091,N_2066);
or U2116 (N_2116,N_2029,N_2033);
and U2117 (N_2117,N_2086,N_2088);
xnor U2118 (N_2118,N_2043,N_2060);
nor U2119 (N_2119,N_2048,N_2058);
xor U2120 (N_2120,N_2096,N_2059);
nor U2121 (N_2121,N_2025,N_2063);
and U2122 (N_2122,N_2026,N_2027);
and U2123 (N_2123,N_2074,N_2041);
xnor U2124 (N_2124,N_2032,N_2067);
nor U2125 (N_2125,N_2072,N_2094);
and U2126 (N_2126,N_2092,N_2075);
nor U2127 (N_2127,N_2034,N_2054);
and U2128 (N_2128,N_2046,N_2028);
and U2129 (N_2129,N_2053,N_2070);
or U2130 (N_2130,N_2052,N_2083);
and U2131 (N_2131,N_2036,N_2079);
nor U2132 (N_2132,N_2061,N_2050);
xor U2133 (N_2133,N_2081,N_2073);
or U2134 (N_2134,N_2093,N_2057);
or U2135 (N_2135,N_2090,N_2042);
xnor U2136 (N_2136,N_2084,N_2031);
or U2137 (N_2137,N_2080,N_2057);
nand U2138 (N_2138,N_2078,N_2079);
xor U2139 (N_2139,N_2042,N_2072);
and U2140 (N_2140,N_2086,N_2025);
or U2141 (N_2141,N_2027,N_2041);
or U2142 (N_2142,N_2056,N_2066);
nand U2143 (N_2143,N_2040,N_2031);
and U2144 (N_2144,N_2048,N_2075);
and U2145 (N_2145,N_2037,N_2079);
and U2146 (N_2146,N_2096,N_2075);
or U2147 (N_2147,N_2097,N_2042);
or U2148 (N_2148,N_2084,N_2078);
nand U2149 (N_2149,N_2092,N_2088);
nor U2150 (N_2150,N_2041,N_2082);
xor U2151 (N_2151,N_2082,N_2047);
xor U2152 (N_2152,N_2029,N_2063);
nand U2153 (N_2153,N_2031,N_2036);
nand U2154 (N_2154,N_2090,N_2026);
nand U2155 (N_2155,N_2073,N_2041);
xor U2156 (N_2156,N_2035,N_2080);
nor U2157 (N_2157,N_2042,N_2035);
or U2158 (N_2158,N_2098,N_2026);
nand U2159 (N_2159,N_2026,N_2028);
xnor U2160 (N_2160,N_2049,N_2062);
xor U2161 (N_2161,N_2067,N_2025);
or U2162 (N_2162,N_2085,N_2056);
nor U2163 (N_2163,N_2073,N_2074);
and U2164 (N_2164,N_2086,N_2060);
or U2165 (N_2165,N_2092,N_2043);
nor U2166 (N_2166,N_2030,N_2026);
xnor U2167 (N_2167,N_2045,N_2099);
and U2168 (N_2168,N_2061,N_2046);
or U2169 (N_2169,N_2063,N_2032);
and U2170 (N_2170,N_2072,N_2071);
and U2171 (N_2171,N_2081,N_2089);
nand U2172 (N_2172,N_2026,N_2071);
xor U2173 (N_2173,N_2060,N_2087);
nand U2174 (N_2174,N_2094,N_2077);
xor U2175 (N_2175,N_2161,N_2122);
and U2176 (N_2176,N_2110,N_2116);
nand U2177 (N_2177,N_2174,N_2163);
nand U2178 (N_2178,N_2155,N_2130);
or U2179 (N_2179,N_2133,N_2162);
nor U2180 (N_2180,N_2169,N_2146);
nand U2181 (N_2181,N_2100,N_2103);
or U2182 (N_2182,N_2135,N_2117);
nor U2183 (N_2183,N_2112,N_2111);
and U2184 (N_2184,N_2141,N_2173);
or U2185 (N_2185,N_2151,N_2102);
nand U2186 (N_2186,N_2106,N_2147);
and U2187 (N_2187,N_2160,N_2114);
xor U2188 (N_2188,N_2115,N_2104);
nand U2189 (N_2189,N_2123,N_2125);
nor U2190 (N_2190,N_2120,N_2157);
or U2191 (N_2191,N_2172,N_2109);
xnor U2192 (N_2192,N_2142,N_2134);
and U2193 (N_2193,N_2148,N_2136);
and U2194 (N_2194,N_2159,N_2121);
and U2195 (N_2195,N_2126,N_2101);
xor U2196 (N_2196,N_2153,N_2168);
or U2197 (N_2197,N_2165,N_2107);
and U2198 (N_2198,N_2164,N_2128);
xnor U2199 (N_2199,N_2144,N_2156);
xnor U2200 (N_2200,N_2124,N_2149);
xor U2201 (N_2201,N_2127,N_2143);
xnor U2202 (N_2202,N_2170,N_2119);
and U2203 (N_2203,N_2139,N_2140);
xor U2204 (N_2204,N_2152,N_2154);
nand U2205 (N_2205,N_2129,N_2113);
and U2206 (N_2206,N_2138,N_2137);
nand U2207 (N_2207,N_2105,N_2167);
nor U2208 (N_2208,N_2108,N_2131);
and U2209 (N_2209,N_2118,N_2150);
nand U2210 (N_2210,N_2132,N_2166);
nand U2211 (N_2211,N_2158,N_2145);
xor U2212 (N_2212,N_2171,N_2168);
and U2213 (N_2213,N_2102,N_2120);
and U2214 (N_2214,N_2171,N_2155);
and U2215 (N_2215,N_2139,N_2150);
and U2216 (N_2216,N_2107,N_2163);
or U2217 (N_2217,N_2170,N_2102);
nor U2218 (N_2218,N_2131,N_2152);
nor U2219 (N_2219,N_2138,N_2107);
xor U2220 (N_2220,N_2157,N_2139);
nand U2221 (N_2221,N_2108,N_2161);
nor U2222 (N_2222,N_2109,N_2105);
nor U2223 (N_2223,N_2158,N_2104);
nand U2224 (N_2224,N_2174,N_2107);
nand U2225 (N_2225,N_2103,N_2166);
or U2226 (N_2226,N_2118,N_2135);
xor U2227 (N_2227,N_2162,N_2124);
nor U2228 (N_2228,N_2108,N_2153);
and U2229 (N_2229,N_2155,N_2103);
nand U2230 (N_2230,N_2101,N_2149);
or U2231 (N_2231,N_2157,N_2163);
xnor U2232 (N_2232,N_2129,N_2110);
nand U2233 (N_2233,N_2128,N_2170);
nand U2234 (N_2234,N_2117,N_2102);
and U2235 (N_2235,N_2123,N_2141);
or U2236 (N_2236,N_2153,N_2115);
nand U2237 (N_2237,N_2140,N_2104);
nor U2238 (N_2238,N_2151,N_2174);
or U2239 (N_2239,N_2125,N_2152);
nand U2240 (N_2240,N_2111,N_2149);
xnor U2241 (N_2241,N_2161,N_2158);
nand U2242 (N_2242,N_2149,N_2161);
or U2243 (N_2243,N_2161,N_2159);
and U2244 (N_2244,N_2115,N_2145);
or U2245 (N_2245,N_2120,N_2126);
and U2246 (N_2246,N_2117,N_2150);
xor U2247 (N_2247,N_2128,N_2104);
nor U2248 (N_2248,N_2120,N_2155);
nor U2249 (N_2249,N_2143,N_2117);
or U2250 (N_2250,N_2239,N_2183);
and U2251 (N_2251,N_2197,N_2248);
or U2252 (N_2252,N_2178,N_2232);
nor U2253 (N_2253,N_2236,N_2217);
nand U2254 (N_2254,N_2247,N_2195);
nor U2255 (N_2255,N_2216,N_2226);
nand U2256 (N_2256,N_2219,N_2175);
or U2257 (N_2257,N_2198,N_2204);
and U2258 (N_2258,N_2209,N_2184);
nand U2259 (N_2259,N_2213,N_2194);
nor U2260 (N_2260,N_2210,N_2193);
and U2261 (N_2261,N_2203,N_2221);
nand U2262 (N_2262,N_2207,N_2233);
xnor U2263 (N_2263,N_2223,N_2230);
xor U2264 (N_2264,N_2218,N_2205);
or U2265 (N_2265,N_2245,N_2220);
or U2266 (N_2266,N_2225,N_2199);
or U2267 (N_2267,N_2235,N_2212);
and U2268 (N_2268,N_2215,N_2234);
nor U2269 (N_2269,N_2182,N_2224);
nand U2270 (N_2270,N_2229,N_2176);
xnor U2271 (N_2271,N_2191,N_2202);
nand U2272 (N_2272,N_2240,N_2181);
xnor U2273 (N_2273,N_2186,N_2188);
nand U2274 (N_2274,N_2206,N_2227);
and U2275 (N_2275,N_2196,N_2243);
xnor U2276 (N_2276,N_2177,N_2241);
nand U2277 (N_2277,N_2211,N_2214);
nor U2278 (N_2278,N_2249,N_2246);
xor U2279 (N_2279,N_2237,N_2192);
xor U2280 (N_2280,N_2244,N_2231);
nor U2281 (N_2281,N_2190,N_2200);
xnor U2282 (N_2282,N_2222,N_2238);
or U2283 (N_2283,N_2187,N_2185);
xnor U2284 (N_2284,N_2201,N_2180);
nand U2285 (N_2285,N_2179,N_2228);
nand U2286 (N_2286,N_2208,N_2189);
xor U2287 (N_2287,N_2242,N_2210);
and U2288 (N_2288,N_2235,N_2225);
xnor U2289 (N_2289,N_2192,N_2231);
or U2290 (N_2290,N_2194,N_2241);
xnor U2291 (N_2291,N_2245,N_2211);
nand U2292 (N_2292,N_2182,N_2207);
or U2293 (N_2293,N_2225,N_2236);
nor U2294 (N_2294,N_2188,N_2238);
or U2295 (N_2295,N_2194,N_2243);
and U2296 (N_2296,N_2228,N_2218);
and U2297 (N_2297,N_2233,N_2214);
or U2298 (N_2298,N_2217,N_2210);
or U2299 (N_2299,N_2221,N_2201);
nand U2300 (N_2300,N_2185,N_2199);
and U2301 (N_2301,N_2216,N_2202);
and U2302 (N_2302,N_2189,N_2211);
xnor U2303 (N_2303,N_2181,N_2218);
nand U2304 (N_2304,N_2204,N_2246);
nor U2305 (N_2305,N_2223,N_2236);
nor U2306 (N_2306,N_2237,N_2236);
or U2307 (N_2307,N_2176,N_2225);
xnor U2308 (N_2308,N_2235,N_2205);
and U2309 (N_2309,N_2194,N_2185);
or U2310 (N_2310,N_2185,N_2223);
nor U2311 (N_2311,N_2197,N_2189);
nor U2312 (N_2312,N_2189,N_2216);
or U2313 (N_2313,N_2176,N_2199);
nor U2314 (N_2314,N_2206,N_2240);
nor U2315 (N_2315,N_2194,N_2210);
nand U2316 (N_2316,N_2229,N_2211);
nand U2317 (N_2317,N_2221,N_2249);
nand U2318 (N_2318,N_2247,N_2248);
nand U2319 (N_2319,N_2242,N_2238);
xnor U2320 (N_2320,N_2222,N_2185);
or U2321 (N_2321,N_2210,N_2232);
nor U2322 (N_2322,N_2234,N_2175);
or U2323 (N_2323,N_2243,N_2176);
xor U2324 (N_2324,N_2208,N_2225);
xnor U2325 (N_2325,N_2315,N_2324);
xor U2326 (N_2326,N_2257,N_2268);
or U2327 (N_2327,N_2313,N_2263);
and U2328 (N_2328,N_2251,N_2278);
or U2329 (N_2329,N_2304,N_2293);
xor U2330 (N_2330,N_2297,N_2286);
and U2331 (N_2331,N_2308,N_2289);
xor U2332 (N_2332,N_2292,N_2294);
xnor U2333 (N_2333,N_2319,N_2266);
and U2334 (N_2334,N_2250,N_2274);
nor U2335 (N_2335,N_2253,N_2302);
or U2336 (N_2336,N_2320,N_2287);
nand U2337 (N_2337,N_2271,N_2279);
and U2338 (N_2338,N_2281,N_2273);
nand U2339 (N_2339,N_2322,N_2284);
and U2340 (N_2340,N_2312,N_2318);
nand U2341 (N_2341,N_2269,N_2306);
xor U2342 (N_2342,N_2288,N_2262);
nand U2343 (N_2343,N_2307,N_2280);
xor U2344 (N_2344,N_2317,N_2265);
or U2345 (N_2345,N_2277,N_2323);
and U2346 (N_2346,N_2252,N_2300);
and U2347 (N_2347,N_2285,N_2258);
nand U2348 (N_2348,N_2290,N_2256);
xor U2349 (N_2349,N_2303,N_2301);
or U2350 (N_2350,N_2255,N_2259);
nor U2351 (N_2351,N_2283,N_2316);
or U2352 (N_2352,N_2264,N_2260);
and U2353 (N_2353,N_2267,N_2314);
and U2354 (N_2354,N_2311,N_2270);
xnor U2355 (N_2355,N_2321,N_2254);
xor U2356 (N_2356,N_2291,N_2261);
xnor U2357 (N_2357,N_2298,N_2310);
nand U2358 (N_2358,N_2295,N_2276);
nand U2359 (N_2359,N_2305,N_2296);
nor U2360 (N_2360,N_2272,N_2282);
nor U2361 (N_2361,N_2299,N_2309);
nor U2362 (N_2362,N_2275,N_2302);
or U2363 (N_2363,N_2271,N_2305);
or U2364 (N_2364,N_2255,N_2295);
or U2365 (N_2365,N_2293,N_2303);
nand U2366 (N_2366,N_2285,N_2256);
xor U2367 (N_2367,N_2306,N_2297);
nor U2368 (N_2368,N_2313,N_2311);
nor U2369 (N_2369,N_2282,N_2296);
nand U2370 (N_2370,N_2311,N_2285);
or U2371 (N_2371,N_2260,N_2262);
and U2372 (N_2372,N_2299,N_2285);
and U2373 (N_2373,N_2266,N_2304);
nand U2374 (N_2374,N_2299,N_2316);
and U2375 (N_2375,N_2252,N_2279);
nor U2376 (N_2376,N_2264,N_2296);
nor U2377 (N_2377,N_2269,N_2253);
xor U2378 (N_2378,N_2296,N_2306);
or U2379 (N_2379,N_2266,N_2281);
or U2380 (N_2380,N_2270,N_2302);
or U2381 (N_2381,N_2314,N_2321);
and U2382 (N_2382,N_2294,N_2260);
nor U2383 (N_2383,N_2293,N_2297);
and U2384 (N_2384,N_2257,N_2310);
or U2385 (N_2385,N_2303,N_2267);
xor U2386 (N_2386,N_2302,N_2282);
or U2387 (N_2387,N_2303,N_2289);
and U2388 (N_2388,N_2272,N_2277);
or U2389 (N_2389,N_2274,N_2290);
and U2390 (N_2390,N_2310,N_2317);
nor U2391 (N_2391,N_2321,N_2320);
or U2392 (N_2392,N_2271,N_2298);
or U2393 (N_2393,N_2280,N_2304);
or U2394 (N_2394,N_2318,N_2280);
xnor U2395 (N_2395,N_2313,N_2269);
xnor U2396 (N_2396,N_2268,N_2308);
nor U2397 (N_2397,N_2277,N_2298);
or U2398 (N_2398,N_2315,N_2257);
or U2399 (N_2399,N_2267,N_2296);
xor U2400 (N_2400,N_2352,N_2359);
and U2401 (N_2401,N_2392,N_2335);
or U2402 (N_2402,N_2371,N_2381);
nand U2403 (N_2403,N_2349,N_2347);
and U2404 (N_2404,N_2330,N_2396);
or U2405 (N_2405,N_2399,N_2345);
xnor U2406 (N_2406,N_2386,N_2387);
or U2407 (N_2407,N_2336,N_2397);
nor U2408 (N_2408,N_2388,N_2383);
and U2409 (N_2409,N_2382,N_2325);
xnor U2410 (N_2410,N_2341,N_2384);
and U2411 (N_2411,N_2385,N_2367);
or U2412 (N_2412,N_2343,N_2373);
xor U2413 (N_2413,N_2334,N_2355);
and U2414 (N_2414,N_2368,N_2333);
and U2415 (N_2415,N_2332,N_2398);
or U2416 (N_2416,N_2357,N_2395);
and U2417 (N_2417,N_2365,N_2331);
xnor U2418 (N_2418,N_2358,N_2393);
nand U2419 (N_2419,N_2342,N_2361);
nor U2420 (N_2420,N_2394,N_2350);
xor U2421 (N_2421,N_2378,N_2391);
and U2422 (N_2422,N_2363,N_2379);
nor U2423 (N_2423,N_2338,N_2326);
xnor U2424 (N_2424,N_2362,N_2337);
xnor U2425 (N_2425,N_2353,N_2380);
nor U2426 (N_2426,N_2370,N_2376);
nor U2427 (N_2427,N_2389,N_2344);
or U2428 (N_2428,N_2372,N_2348);
nand U2429 (N_2429,N_2351,N_2366);
nand U2430 (N_2430,N_2328,N_2374);
nor U2431 (N_2431,N_2354,N_2364);
and U2432 (N_2432,N_2329,N_2360);
and U2433 (N_2433,N_2369,N_2377);
and U2434 (N_2434,N_2340,N_2390);
or U2435 (N_2435,N_2375,N_2346);
or U2436 (N_2436,N_2356,N_2339);
and U2437 (N_2437,N_2327,N_2371);
nand U2438 (N_2438,N_2366,N_2392);
or U2439 (N_2439,N_2366,N_2396);
nand U2440 (N_2440,N_2397,N_2369);
or U2441 (N_2441,N_2393,N_2353);
or U2442 (N_2442,N_2366,N_2325);
xor U2443 (N_2443,N_2370,N_2386);
and U2444 (N_2444,N_2335,N_2338);
or U2445 (N_2445,N_2399,N_2376);
or U2446 (N_2446,N_2340,N_2378);
xnor U2447 (N_2447,N_2333,N_2345);
and U2448 (N_2448,N_2397,N_2325);
nand U2449 (N_2449,N_2328,N_2394);
xor U2450 (N_2450,N_2381,N_2358);
and U2451 (N_2451,N_2334,N_2391);
or U2452 (N_2452,N_2378,N_2346);
nor U2453 (N_2453,N_2356,N_2386);
or U2454 (N_2454,N_2334,N_2383);
nand U2455 (N_2455,N_2370,N_2329);
xor U2456 (N_2456,N_2340,N_2375);
and U2457 (N_2457,N_2390,N_2382);
nand U2458 (N_2458,N_2370,N_2366);
or U2459 (N_2459,N_2355,N_2383);
and U2460 (N_2460,N_2338,N_2360);
nor U2461 (N_2461,N_2397,N_2349);
xnor U2462 (N_2462,N_2373,N_2382);
nor U2463 (N_2463,N_2358,N_2369);
nand U2464 (N_2464,N_2345,N_2366);
or U2465 (N_2465,N_2334,N_2375);
nand U2466 (N_2466,N_2355,N_2347);
or U2467 (N_2467,N_2359,N_2329);
nand U2468 (N_2468,N_2325,N_2372);
and U2469 (N_2469,N_2377,N_2386);
nor U2470 (N_2470,N_2333,N_2387);
and U2471 (N_2471,N_2382,N_2398);
xnor U2472 (N_2472,N_2397,N_2380);
and U2473 (N_2473,N_2376,N_2386);
nor U2474 (N_2474,N_2335,N_2399);
or U2475 (N_2475,N_2426,N_2469);
nand U2476 (N_2476,N_2421,N_2462);
nand U2477 (N_2477,N_2403,N_2430);
or U2478 (N_2478,N_2439,N_2400);
nor U2479 (N_2479,N_2445,N_2470);
nor U2480 (N_2480,N_2471,N_2465);
nor U2481 (N_2481,N_2412,N_2467);
nand U2482 (N_2482,N_2401,N_2436);
or U2483 (N_2483,N_2459,N_2418);
nor U2484 (N_2484,N_2438,N_2419);
nor U2485 (N_2485,N_2468,N_2433);
nand U2486 (N_2486,N_2455,N_2429);
nand U2487 (N_2487,N_2428,N_2464);
or U2488 (N_2488,N_2413,N_2406);
nand U2489 (N_2489,N_2417,N_2449);
nand U2490 (N_2490,N_2423,N_2404);
xor U2491 (N_2491,N_2450,N_2440);
nor U2492 (N_2492,N_2416,N_2473);
xor U2493 (N_2493,N_2454,N_2431);
nand U2494 (N_2494,N_2402,N_2466);
nand U2495 (N_2495,N_2407,N_2458);
or U2496 (N_2496,N_2432,N_2435);
nand U2497 (N_2497,N_2410,N_2442);
nand U2498 (N_2498,N_2456,N_2405);
nor U2499 (N_2499,N_2420,N_2425);
xnor U2500 (N_2500,N_2463,N_2414);
or U2501 (N_2501,N_2451,N_2452);
and U2502 (N_2502,N_2453,N_2408);
and U2503 (N_2503,N_2422,N_2460);
nand U2504 (N_2504,N_2461,N_2409);
xnor U2505 (N_2505,N_2437,N_2411);
xor U2506 (N_2506,N_2447,N_2457);
nor U2507 (N_2507,N_2434,N_2444);
nand U2508 (N_2508,N_2446,N_2443);
and U2509 (N_2509,N_2427,N_2474);
nor U2510 (N_2510,N_2441,N_2472);
nand U2511 (N_2511,N_2415,N_2424);
xor U2512 (N_2512,N_2448,N_2470);
and U2513 (N_2513,N_2436,N_2438);
and U2514 (N_2514,N_2406,N_2459);
xor U2515 (N_2515,N_2439,N_2432);
or U2516 (N_2516,N_2434,N_2427);
xnor U2517 (N_2517,N_2464,N_2445);
and U2518 (N_2518,N_2434,N_2430);
nor U2519 (N_2519,N_2430,N_2432);
nor U2520 (N_2520,N_2463,N_2436);
nor U2521 (N_2521,N_2447,N_2449);
nor U2522 (N_2522,N_2423,N_2470);
or U2523 (N_2523,N_2463,N_2459);
and U2524 (N_2524,N_2415,N_2456);
xnor U2525 (N_2525,N_2432,N_2438);
or U2526 (N_2526,N_2419,N_2460);
or U2527 (N_2527,N_2474,N_2469);
nand U2528 (N_2528,N_2433,N_2451);
or U2529 (N_2529,N_2412,N_2423);
nand U2530 (N_2530,N_2436,N_2450);
nand U2531 (N_2531,N_2429,N_2437);
or U2532 (N_2532,N_2446,N_2425);
xnor U2533 (N_2533,N_2443,N_2405);
nand U2534 (N_2534,N_2416,N_2460);
and U2535 (N_2535,N_2412,N_2455);
or U2536 (N_2536,N_2412,N_2473);
xnor U2537 (N_2537,N_2414,N_2452);
nand U2538 (N_2538,N_2401,N_2466);
nor U2539 (N_2539,N_2409,N_2446);
or U2540 (N_2540,N_2461,N_2438);
and U2541 (N_2541,N_2420,N_2427);
or U2542 (N_2542,N_2444,N_2454);
or U2543 (N_2543,N_2409,N_2449);
nor U2544 (N_2544,N_2422,N_2442);
and U2545 (N_2545,N_2403,N_2467);
nand U2546 (N_2546,N_2431,N_2411);
or U2547 (N_2547,N_2408,N_2449);
xnor U2548 (N_2548,N_2458,N_2467);
nand U2549 (N_2549,N_2407,N_2445);
or U2550 (N_2550,N_2478,N_2539);
or U2551 (N_2551,N_2506,N_2489);
nor U2552 (N_2552,N_2547,N_2494);
or U2553 (N_2553,N_2488,N_2502);
nor U2554 (N_2554,N_2479,N_2483);
xnor U2555 (N_2555,N_2533,N_2515);
or U2556 (N_2556,N_2517,N_2514);
and U2557 (N_2557,N_2480,N_2544);
xnor U2558 (N_2558,N_2500,N_2531);
nor U2559 (N_2559,N_2520,N_2496);
or U2560 (N_2560,N_2535,N_2513);
xnor U2561 (N_2561,N_2490,N_2542);
and U2562 (N_2562,N_2487,N_2532);
xor U2563 (N_2563,N_2485,N_2512);
nand U2564 (N_2564,N_2484,N_2525);
nand U2565 (N_2565,N_2497,N_2523);
or U2566 (N_2566,N_2522,N_2476);
and U2567 (N_2567,N_2495,N_2538);
or U2568 (N_2568,N_2499,N_2509);
xor U2569 (N_2569,N_2516,N_2508);
or U2570 (N_2570,N_2518,N_2503);
nor U2571 (N_2571,N_2545,N_2549);
nor U2572 (N_2572,N_2504,N_2537);
and U2573 (N_2573,N_2501,N_2548);
nand U2574 (N_2574,N_2486,N_2510);
and U2575 (N_2575,N_2505,N_2492);
nand U2576 (N_2576,N_2477,N_2530);
xor U2577 (N_2577,N_2475,N_2546);
nor U2578 (N_2578,N_2482,N_2507);
nand U2579 (N_2579,N_2528,N_2491);
xor U2580 (N_2580,N_2521,N_2541);
or U2581 (N_2581,N_2524,N_2534);
or U2582 (N_2582,N_2527,N_2526);
or U2583 (N_2583,N_2536,N_2529);
xor U2584 (N_2584,N_2543,N_2540);
nand U2585 (N_2585,N_2481,N_2498);
and U2586 (N_2586,N_2493,N_2519);
nand U2587 (N_2587,N_2511,N_2509);
nand U2588 (N_2588,N_2526,N_2494);
nand U2589 (N_2589,N_2479,N_2544);
and U2590 (N_2590,N_2525,N_2483);
and U2591 (N_2591,N_2520,N_2482);
nor U2592 (N_2592,N_2545,N_2486);
and U2593 (N_2593,N_2533,N_2535);
nor U2594 (N_2594,N_2522,N_2530);
nor U2595 (N_2595,N_2479,N_2543);
nand U2596 (N_2596,N_2531,N_2523);
nand U2597 (N_2597,N_2506,N_2538);
or U2598 (N_2598,N_2500,N_2543);
nor U2599 (N_2599,N_2480,N_2539);
nand U2600 (N_2600,N_2496,N_2544);
xnor U2601 (N_2601,N_2513,N_2520);
xor U2602 (N_2602,N_2495,N_2543);
nand U2603 (N_2603,N_2546,N_2542);
and U2604 (N_2604,N_2514,N_2511);
or U2605 (N_2605,N_2511,N_2512);
and U2606 (N_2606,N_2504,N_2517);
xor U2607 (N_2607,N_2499,N_2549);
or U2608 (N_2608,N_2535,N_2512);
nand U2609 (N_2609,N_2548,N_2483);
nor U2610 (N_2610,N_2496,N_2525);
and U2611 (N_2611,N_2515,N_2521);
or U2612 (N_2612,N_2480,N_2487);
and U2613 (N_2613,N_2542,N_2523);
xnor U2614 (N_2614,N_2544,N_2483);
xnor U2615 (N_2615,N_2541,N_2480);
nor U2616 (N_2616,N_2548,N_2484);
nand U2617 (N_2617,N_2514,N_2483);
nor U2618 (N_2618,N_2541,N_2495);
xnor U2619 (N_2619,N_2500,N_2525);
nand U2620 (N_2620,N_2485,N_2523);
xor U2621 (N_2621,N_2538,N_2535);
nand U2622 (N_2622,N_2534,N_2509);
or U2623 (N_2623,N_2525,N_2477);
nand U2624 (N_2624,N_2485,N_2479);
or U2625 (N_2625,N_2561,N_2576);
or U2626 (N_2626,N_2568,N_2559);
and U2627 (N_2627,N_2554,N_2571);
or U2628 (N_2628,N_2589,N_2622);
xnor U2629 (N_2629,N_2588,N_2621);
xnor U2630 (N_2630,N_2565,N_2581);
or U2631 (N_2631,N_2603,N_2607);
nand U2632 (N_2632,N_2585,N_2600);
nand U2633 (N_2633,N_2580,N_2557);
xnor U2634 (N_2634,N_2555,N_2587);
or U2635 (N_2635,N_2606,N_2601);
and U2636 (N_2636,N_2586,N_2579);
nand U2637 (N_2637,N_2550,N_2605);
nand U2638 (N_2638,N_2558,N_2623);
or U2639 (N_2639,N_2562,N_2611);
or U2640 (N_2640,N_2613,N_2567);
nor U2641 (N_2641,N_2598,N_2624);
nor U2642 (N_2642,N_2616,N_2596);
nand U2643 (N_2643,N_2612,N_2570);
or U2644 (N_2644,N_2617,N_2595);
xor U2645 (N_2645,N_2591,N_2597);
xor U2646 (N_2646,N_2594,N_2608);
nand U2647 (N_2647,N_2573,N_2556);
nand U2648 (N_2648,N_2574,N_2560);
xor U2649 (N_2649,N_2609,N_2590);
or U2650 (N_2650,N_2575,N_2614);
nand U2651 (N_2651,N_2582,N_2618);
xor U2652 (N_2652,N_2615,N_2577);
nor U2653 (N_2653,N_2583,N_2593);
xor U2654 (N_2654,N_2619,N_2592);
nand U2655 (N_2655,N_2553,N_2572);
xor U2656 (N_2656,N_2563,N_2604);
or U2657 (N_2657,N_2569,N_2610);
nand U2658 (N_2658,N_2566,N_2599);
and U2659 (N_2659,N_2564,N_2551);
nor U2660 (N_2660,N_2602,N_2620);
xor U2661 (N_2661,N_2552,N_2578);
or U2662 (N_2662,N_2584,N_2554);
xor U2663 (N_2663,N_2580,N_2560);
and U2664 (N_2664,N_2601,N_2573);
or U2665 (N_2665,N_2587,N_2597);
xnor U2666 (N_2666,N_2594,N_2592);
xnor U2667 (N_2667,N_2611,N_2624);
nor U2668 (N_2668,N_2561,N_2604);
or U2669 (N_2669,N_2613,N_2601);
nor U2670 (N_2670,N_2605,N_2593);
or U2671 (N_2671,N_2579,N_2612);
or U2672 (N_2672,N_2619,N_2601);
and U2673 (N_2673,N_2558,N_2567);
or U2674 (N_2674,N_2591,N_2616);
and U2675 (N_2675,N_2591,N_2596);
nand U2676 (N_2676,N_2569,N_2563);
xor U2677 (N_2677,N_2595,N_2612);
and U2678 (N_2678,N_2569,N_2576);
and U2679 (N_2679,N_2551,N_2578);
xor U2680 (N_2680,N_2611,N_2594);
and U2681 (N_2681,N_2594,N_2562);
or U2682 (N_2682,N_2615,N_2568);
nor U2683 (N_2683,N_2564,N_2569);
nor U2684 (N_2684,N_2614,N_2589);
nor U2685 (N_2685,N_2620,N_2619);
or U2686 (N_2686,N_2622,N_2605);
and U2687 (N_2687,N_2590,N_2558);
and U2688 (N_2688,N_2600,N_2616);
xnor U2689 (N_2689,N_2612,N_2567);
or U2690 (N_2690,N_2614,N_2553);
and U2691 (N_2691,N_2603,N_2571);
nor U2692 (N_2692,N_2590,N_2619);
xnor U2693 (N_2693,N_2617,N_2590);
nor U2694 (N_2694,N_2599,N_2570);
nand U2695 (N_2695,N_2585,N_2609);
nand U2696 (N_2696,N_2594,N_2581);
or U2697 (N_2697,N_2553,N_2623);
xnor U2698 (N_2698,N_2597,N_2613);
xor U2699 (N_2699,N_2619,N_2560);
xnor U2700 (N_2700,N_2689,N_2666);
or U2701 (N_2701,N_2667,N_2631);
and U2702 (N_2702,N_2641,N_2658);
or U2703 (N_2703,N_2688,N_2673);
nand U2704 (N_2704,N_2644,N_2678);
or U2705 (N_2705,N_2677,N_2634);
nand U2706 (N_2706,N_2640,N_2676);
or U2707 (N_2707,N_2661,N_2687);
xor U2708 (N_2708,N_2636,N_2649);
nor U2709 (N_2709,N_2680,N_2638);
and U2710 (N_2710,N_2628,N_2691);
nor U2711 (N_2711,N_2629,N_2665);
and U2712 (N_2712,N_2681,N_2692);
nand U2713 (N_2713,N_2682,N_2650);
nand U2714 (N_2714,N_2625,N_2693);
xnor U2715 (N_2715,N_2664,N_2651);
or U2716 (N_2716,N_2655,N_2659);
and U2717 (N_2717,N_2660,N_2685);
or U2718 (N_2718,N_2663,N_2647);
nor U2719 (N_2719,N_2646,N_2656);
or U2720 (N_2720,N_2639,N_2635);
xnor U2721 (N_2721,N_2697,N_2674);
xnor U2722 (N_2722,N_2698,N_2627);
nor U2723 (N_2723,N_2654,N_2679);
xor U2724 (N_2724,N_2652,N_2642);
nand U2725 (N_2725,N_2653,N_2645);
xor U2726 (N_2726,N_2696,N_2637);
or U2727 (N_2727,N_2668,N_2648);
or U2728 (N_2728,N_2675,N_2684);
nor U2729 (N_2729,N_2699,N_2672);
xnor U2730 (N_2730,N_2662,N_2686);
or U2731 (N_2731,N_2670,N_2630);
xnor U2732 (N_2732,N_2626,N_2671);
or U2733 (N_2733,N_2695,N_2669);
or U2734 (N_2734,N_2633,N_2657);
nand U2735 (N_2735,N_2643,N_2632);
and U2736 (N_2736,N_2683,N_2690);
and U2737 (N_2737,N_2694,N_2650);
xor U2738 (N_2738,N_2660,N_2647);
and U2739 (N_2739,N_2635,N_2680);
nor U2740 (N_2740,N_2687,N_2699);
nor U2741 (N_2741,N_2641,N_2650);
and U2742 (N_2742,N_2674,N_2678);
or U2743 (N_2743,N_2664,N_2674);
nand U2744 (N_2744,N_2660,N_2689);
or U2745 (N_2745,N_2696,N_2675);
nor U2746 (N_2746,N_2663,N_2634);
nand U2747 (N_2747,N_2666,N_2631);
and U2748 (N_2748,N_2684,N_2696);
nor U2749 (N_2749,N_2662,N_2630);
and U2750 (N_2750,N_2645,N_2677);
nor U2751 (N_2751,N_2626,N_2689);
nor U2752 (N_2752,N_2673,N_2689);
or U2753 (N_2753,N_2626,N_2659);
nor U2754 (N_2754,N_2699,N_2682);
nand U2755 (N_2755,N_2672,N_2636);
nor U2756 (N_2756,N_2696,N_2695);
xor U2757 (N_2757,N_2680,N_2684);
or U2758 (N_2758,N_2698,N_2645);
xnor U2759 (N_2759,N_2644,N_2690);
and U2760 (N_2760,N_2659,N_2674);
xnor U2761 (N_2761,N_2656,N_2637);
or U2762 (N_2762,N_2636,N_2657);
nand U2763 (N_2763,N_2656,N_2699);
xnor U2764 (N_2764,N_2688,N_2626);
and U2765 (N_2765,N_2643,N_2627);
xnor U2766 (N_2766,N_2639,N_2645);
or U2767 (N_2767,N_2650,N_2693);
or U2768 (N_2768,N_2663,N_2633);
or U2769 (N_2769,N_2697,N_2687);
xnor U2770 (N_2770,N_2640,N_2641);
nor U2771 (N_2771,N_2686,N_2652);
xnor U2772 (N_2772,N_2660,N_2639);
and U2773 (N_2773,N_2696,N_2655);
nand U2774 (N_2774,N_2642,N_2666);
xnor U2775 (N_2775,N_2764,N_2712);
nand U2776 (N_2776,N_2759,N_2721);
nor U2777 (N_2777,N_2718,N_2728);
and U2778 (N_2778,N_2773,N_2709);
and U2779 (N_2779,N_2719,N_2750);
and U2780 (N_2780,N_2770,N_2741);
nand U2781 (N_2781,N_2704,N_2761);
xnor U2782 (N_2782,N_2760,N_2742);
nand U2783 (N_2783,N_2722,N_2714);
or U2784 (N_2784,N_2735,N_2766);
and U2785 (N_2785,N_2702,N_2758);
xor U2786 (N_2786,N_2710,N_2754);
and U2787 (N_2787,N_2727,N_2767);
nand U2788 (N_2788,N_2752,N_2706);
nor U2789 (N_2789,N_2705,N_2734);
xor U2790 (N_2790,N_2716,N_2724);
and U2791 (N_2791,N_2771,N_2749);
or U2792 (N_2792,N_2723,N_2729);
or U2793 (N_2793,N_2739,N_2756);
or U2794 (N_2794,N_2748,N_2733);
nor U2795 (N_2795,N_2703,N_2726);
or U2796 (N_2796,N_2737,N_2700);
and U2797 (N_2797,N_2772,N_2715);
xnor U2798 (N_2798,N_2747,N_2725);
and U2799 (N_2799,N_2753,N_2740);
nor U2800 (N_2800,N_2701,N_2707);
nor U2801 (N_2801,N_2755,N_2738);
xor U2802 (N_2802,N_2731,N_2736);
or U2803 (N_2803,N_2743,N_2751);
xor U2804 (N_2804,N_2765,N_2713);
xnor U2805 (N_2805,N_2732,N_2757);
or U2806 (N_2806,N_2711,N_2768);
xor U2807 (N_2807,N_2762,N_2769);
or U2808 (N_2808,N_2774,N_2717);
nor U2809 (N_2809,N_2746,N_2720);
or U2810 (N_2810,N_2763,N_2730);
nor U2811 (N_2811,N_2745,N_2744);
or U2812 (N_2812,N_2708,N_2765);
xnor U2813 (N_2813,N_2764,N_2701);
nor U2814 (N_2814,N_2762,N_2730);
and U2815 (N_2815,N_2732,N_2718);
or U2816 (N_2816,N_2754,N_2749);
nand U2817 (N_2817,N_2748,N_2773);
and U2818 (N_2818,N_2702,N_2715);
nor U2819 (N_2819,N_2702,N_2769);
nor U2820 (N_2820,N_2726,N_2711);
nand U2821 (N_2821,N_2750,N_2772);
nor U2822 (N_2822,N_2744,N_2768);
and U2823 (N_2823,N_2703,N_2739);
xnor U2824 (N_2824,N_2711,N_2741);
or U2825 (N_2825,N_2744,N_2705);
nand U2826 (N_2826,N_2714,N_2713);
and U2827 (N_2827,N_2774,N_2732);
or U2828 (N_2828,N_2720,N_2741);
nor U2829 (N_2829,N_2721,N_2731);
nor U2830 (N_2830,N_2711,N_2727);
nand U2831 (N_2831,N_2762,N_2770);
nand U2832 (N_2832,N_2761,N_2721);
nor U2833 (N_2833,N_2700,N_2717);
nor U2834 (N_2834,N_2750,N_2735);
nand U2835 (N_2835,N_2710,N_2732);
or U2836 (N_2836,N_2753,N_2701);
nor U2837 (N_2837,N_2723,N_2770);
and U2838 (N_2838,N_2716,N_2714);
nand U2839 (N_2839,N_2758,N_2711);
nand U2840 (N_2840,N_2767,N_2745);
or U2841 (N_2841,N_2770,N_2763);
and U2842 (N_2842,N_2765,N_2700);
nor U2843 (N_2843,N_2701,N_2756);
nor U2844 (N_2844,N_2713,N_2736);
nor U2845 (N_2845,N_2714,N_2772);
nor U2846 (N_2846,N_2726,N_2759);
nand U2847 (N_2847,N_2740,N_2768);
nand U2848 (N_2848,N_2748,N_2702);
xor U2849 (N_2849,N_2711,N_2704);
nand U2850 (N_2850,N_2826,N_2809);
nor U2851 (N_2851,N_2791,N_2812);
nand U2852 (N_2852,N_2841,N_2831);
and U2853 (N_2853,N_2825,N_2847);
nor U2854 (N_2854,N_2793,N_2800);
xor U2855 (N_2855,N_2794,N_2790);
nor U2856 (N_2856,N_2846,N_2818);
or U2857 (N_2857,N_2781,N_2799);
nor U2858 (N_2858,N_2798,N_2807);
nor U2859 (N_2859,N_2777,N_2816);
nand U2860 (N_2860,N_2796,N_2786);
nor U2861 (N_2861,N_2849,N_2776);
and U2862 (N_2862,N_2815,N_2802);
or U2863 (N_2863,N_2819,N_2840);
and U2864 (N_2864,N_2834,N_2797);
nor U2865 (N_2865,N_2839,N_2820);
or U2866 (N_2866,N_2842,N_2824);
or U2867 (N_2867,N_2832,N_2845);
nand U2868 (N_2868,N_2835,N_2783);
or U2869 (N_2869,N_2789,N_2817);
nand U2870 (N_2870,N_2828,N_2801);
or U2871 (N_2871,N_2827,N_2813);
and U2872 (N_2872,N_2810,N_2804);
nor U2873 (N_2873,N_2829,N_2836);
xnor U2874 (N_2874,N_2795,N_2833);
nor U2875 (N_2875,N_2788,N_2787);
nand U2876 (N_2876,N_2821,N_2784);
nand U2877 (N_2877,N_2837,N_2808);
nand U2878 (N_2878,N_2805,N_2806);
xor U2879 (N_2879,N_2782,N_2803);
xnor U2880 (N_2880,N_2780,N_2838);
or U2881 (N_2881,N_2830,N_2848);
and U2882 (N_2882,N_2785,N_2814);
xor U2883 (N_2883,N_2811,N_2775);
or U2884 (N_2884,N_2823,N_2843);
nor U2885 (N_2885,N_2779,N_2844);
or U2886 (N_2886,N_2778,N_2822);
nand U2887 (N_2887,N_2792,N_2831);
xor U2888 (N_2888,N_2781,N_2844);
or U2889 (N_2889,N_2789,N_2814);
or U2890 (N_2890,N_2804,N_2842);
and U2891 (N_2891,N_2849,N_2810);
xor U2892 (N_2892,N_2799,N_2777);
or U2893 (N_2893,N_2806,N_2840);
or U2894 (N_2894,N_2802,N_2796);
xnor U2895 (N_2895,N_2818,N_2842);
and U2896 (N_2896,N_2780,N_2806);
and U2897 (N_2897,N_2787,N_2790);
and U2898 (N_2898,N_2846,N_2823);
nand U2899 (N_2899,N_2831,N_2838);
nand U2900 (N_2900,N_2777,N_2824);
nor U2901 (N_2901,N_2843,N_2798);
and U2902 (N_2902,N_2822,N_2820);
nand U2903 (N_2903,N_2838,N_2805);
xor U2904 (N_2904,N_2819,N_2794);
and U2905 (N_2905,N_2839,N_2803);
nor U2906 (N_2906,N_2823,N_2792);
and U2907 (N_2907,N_2783,N_2811);
xnor U2908 (N_2908,N_2787,N_2814);
nand U2909 (N_2909,N_2798,N_2818);
xor U2910 (N_2910,N_2814,N_2775);
nand U2911 (N_2911,N_2777,N_2791);
nand U2912 (N_2912,N_2819,N_2823);
and U2913 (N_2913,N_2787,N_2844);
nand U2914 (N_2914,N_2805,N_2804);
nand U2915 (N_2915,N_2824,N_2817);
or U2916 (N_2916,N_2816,N_2803);
xnor U2917 (N_2917,N_2780,N_2778);
xnor U2918 (N_2918,N_2820,N_2806);
nor U2919 (N_2919,N_2802,N_2806);
nor U2920 (N_2920,N_2791,N_2831);
nor U2921 (N_2921,N_2782,N_2800);
and U2922 (N_2922,N_2809,N_2802);
nor U2923 (N_2923,N_2790,N_2829);
nor U2924 (N_2924,N_2782,N_2832);
xor U2925 (N_2925,N_2902,N_2862);
xnor U2926 (N_2926,N_2896,N_2898);
and U2927 (N_2927,N_2911,N_2920);
or U2928 (N_2928,N_2913,N_2912);
or U2929 (N_2929,N_2894,N_2878);
nand U2930 (N_2930,N_2903,N_2866);
or U2931 (N_2931,N_2918,N_2871);
and U2932 (N_2932,N_2850,N_2917);
nand U2933 (N_2933,N_2895,N_2883);
nor U2934 (N_2934,N_2885,N_2857);
and U2935 (N_2935,N_2873,N_2916);
and U2936 (N_2936,N_2861,N_2859);
nand U2937 (N_2937,N_2900,N_2893);
or U2938 (N_2938,N_2910,N_2879);
nor U2939 (N_2939,N_2884,N_2867);
nor U2940 (N_2940,N_2909,N_2924);
nand U2941 (N_2941,N_2856,N_2858);
or U2942 (N_2942,N_2922,N_2921);
nor U2943 (N_2943,N_2881,N_2906);
nand U2944 (N_2944,N_2892,N_2880);
nand U2945 (N_2945,N_2890,N_2853);
nor U2946 (N_2946,N_2901,N_2872);
or U2947 (N_2947,N_2868,N_2907);
or U2948 (N_2948,N_2882,N_2869);
and U2949 (N_2949,N_2863,N_2886);
or U2950 (N_2950,N_2875,N_2852);
and U2951 (N_2951,N_2876,N_2855);
xor U2952 (N_2952,N_2915,N_2897);
nor U2953 (N_2953,N_2923,N_2887);
nand U2954 (N_2954,N_2874,N_2891);
nor U2955 (N_2955,N_2864,N_2877);
nor U2956 (N_2956,N_2860,N_2899);
and U2957 (N_2957,N_2905,N_2908);
or U2958 (N_2958,N_2854,N_2870);
and U2959 (N_2959,N_2851,N_2888);
or U2960 (N_2960,N_2865,N_2904);
or U2961 (N_2961,N_2914,N_2919);
nand U2962 (N_2962,N_2889,N_2911);
and U2963 (N_2963,N_2885,N_2915);
or U2964 (N_2964,N_2890,N_2897);
xnor U2965 (N_2965,N_2870,N_2889);
nor U2966 (N_2966,N_2896,N_2905);
or U2967 (N_2967,N_2875,N_2856);
nand U2968 (N_2968,N_2872,N_2875);
and U2969 (N_2969,N_2872,N_2921);
or U2970 (N_2970,N_2864,N_2904);
or U2971 (N_2971,N_2891,N_2855);
and U2972 (N_2972,N_2857,N_2854);
nand U2973 (N_2973,N_2874,N_2922);
nand U2974 (N_2974,N_2904,N_2879);
and U2975 (N_2975,N_2857,N_2909);
nand U2976 (N_2976,N_2853,N_2910);
nor U2977 (N_2977,N_2864,N_2916);
nor U2978 (N_2978,N_2872,N_2898);
xor U2979 (N_2979,N_2905,N_2882);
or U2980 (N_2980,N_2900,N_2890);
xor U2981 (N_2981,N_2868,N_2856);
xnor U2982 (N_2982,N_2858,N_2853);
nor U2983 (N_2983,N_2873,N_2897);
nand U2984 (N_2984,N_2893,N_2877);
nor U2985 (N_2985,N_2874,N_2887);
nor U2986 (N_2986,N_2918,N_2877);
or U2987 (N_2987,N_2894,N_2888);
nor U2988 (N_2988,N_2892,N_2885);
or U2989 (N_2989,N_2922,N_2886);
nand U2990 (N_2990,N_2871,N_2919);
nor U2991 (N_2991,N_2878,N_2880);
xnor U2992 (N_2992,N_2908,N_2864);
or U2993 (N_2993,N_2873,N_2882);
nand U2994 (N_2994,N_2906,N_2854);
or U2995 (N_2995,N_2862,N_2860);
xnor U2996 (N_2996,N_2911,N_2923);
or U2997 (N_2997,N_2911,N_2881);
nand U2998 (N_2998,N_2876,N_2872);
and U2999 (N_2999,N_2905,N_2871);
nand UO_0 (O_0,N_2958,N_2992);
or UO_1 (O_1,N_2964,N_2951);
nor UO_2 (O_2,N_2956,N_2945);
and UO_3 (O_3,N_2931,N_2952);
or UO_4 (O_4,N_2934,N_2962);
and UO_5 (O_5,N_2989,N_2981);
nor UO_6 (O_6,N_2959,N_2974);
xor UO_7 (O_7,N_2982,N_2999);
nand UO_8 (O_8,N_2939,N_2997);
nand UO_9 (O_9,N_2957,N_2947);
or UO_10 (O_10,N_2971,N_2984);
nand UO_11 (O_11,N_2938,N_2973);
or UO_12 (O_12,N_2978,N_2954);
xor UO_13 (O_13,N_2967,N_2980);
nand UO_14 (O_14,N_2936,N_2941);
and UO_15 (O_15,N_2942,N_2944);
nor UO_16 (O_16,N_2977,N_2927);
xor UO_17 (O_17,N_2937,N_2976);
nand UO_18 (O_18,N_2970,N_2943);
nand UO_19 (O_19,N_2991,N_2987);
nor UO_20 (O_20,N_2949,N_2928);
xnor UO_21 (O_21,N_2990,N_2950);
xnor UO_22 (O_22,N_2929,N_2986);
nor UO_23 (O_23,N_2926,N_2975);
and UO_24 (O_24,N_2994,N_2965);
nand UO_25 (O_25,N_2995,N_2979);
nor UO_26 (O_26,N_2948,N_2935);
nor UO_27 (O_27,N_2966,N_2968);
and UO_28 (O_28,N_2946,N_2953);
nand UO_29 (O_29,N_2983,N_2940);
nor UO_30 (O_30,N_2985,N_2932);
or UO_31 (O_31,N_2961,N_2969);
nand UO_32 (O_32,N_2993,N_2955);
or UO_33 (O_33,N_2933,N_2988);
nor UO_34 (O_34,N_2925,N_2996);
or UO_35 (O_35,N_2972,N_2930);
nor UO_36 (O_36,N_2998,N_2960);
nand UO_37 (O_37,N_2963,N_2937);
nand UO_38 (O_38,N_2939,N_2988);
xor UO_39 (O_39,N_2963,N_2926);
xor UO_40 (O_40,N_2983,N_2970);
and UO_41 (O_41,N_2952,N_2948);
and UO_42 (O_42,N_2962,N_2999);
or UO_43 (O_43,N_2940,N_2995);
and UO_44 (O_44,N_2962,N_2954);
nor UO_45 (O_45,N_2999,N_2973);
xor UO_46 (O_46,N_2995,N_2933);
nor UO_47 (O_47,N_2979,N_2972);
nand UO_48 (O_48,N_2926,N_2945);
nor UO_49 (O_49,N_2939,N_2999);
nor UO_50 (O_50,N_2984,N_2925);
nand UO_51 (O_51,N_2933,N_2949);
xor UO_52 (O_52,N_2928,N_2993);
nor UO_53 (O_53,N_2930,N_2974);
nand UO_54 (O_54,N_2967,N_2949);
nand UO_55 (O_55,N_2961,N_2926);
nand UO_56 (O_56,N_2947,N_2975);
or UO_57 (O_57,N_2925,N_2952);
and UO_58 (O_58,N_2978,N_2996);
nor UO_59 (O_59,N_2958,N_2998);
nor UO_60 (O_60,N_2995,N_2978);
nor UO_61 (O_61,N_2962,N_2953);
nand UO_62 (O_62,N_2989,N_2943);
nor UO_63 (O_63,N_2943,N_2952);
xnor UO_64 (O_64,N_2969,N_2978);
xor UO_65 (O_65,N_2956,N_2971);
or UO_66 (O_66,N_2942,N_2967);
nand UO_67 (O_67,N_2955,N_2965);
nor UO_68 (O_68,N_2963,N_2999);
xor UO_69 (O_69,N_2928,N_2957);
xnor UO_70 (O_70,N_2987,N_2982);
nand UO_71 (O_71,N_2947,N_2954);
nand UO_72 (O_72,N_2958,N_2959);
nor UO_73 (O_73,N_2971,N_2952);
and UO_74 (O_74,N_2939,N_2961);
or UO_75 (O_75,N_2962,N_2943);
xnor UO_76 (O_76,N_2972,N_2931);
nand UO_77 (O_77,N_2972,N_2995);
and UO_78 (O_78,N_2980,N_2932);
or UO_79 (O_79,N_2997,N_2990);
or UO_80 (O_80,N_2948,N_2981);
nand UO_81 (O_81,N_2996,N_2929);
xor UO_82 (O_82,N_2979,N_2968);
xor UO_83 (O_83,N_2934,N_2973);
xor UO_84 (O_84,N_2957,N_2976);
and UO_85 (O_85,N_2977,N_2969);
or UO_86 (O_86,N_2972,N_2984);
nand UO_87 (O_87,N_2945,N_2994);
or UO_88 (O_88,N_2931,N_2961);
nand UO_89 (O_89,N_2987,N_2931);
and UO_90 (O_90,N_2974,N_2958);
nand UO_91 (O_91,N_2942,N_2947);
or UO_92 (O_92,N_2959,N_2988);
nand UO_93 (O_93,N_2985,N_2957);
nand UO_94 (O_94,N_2970,N_2979);
nor UO_95 (O_95,N_2938,N_2958);
nor UO_96 (O_96,N_2941,N_2978);
nand UO_97 (O_97,N_2952,N_2946);
and UO_98 (O_98,N_2967,N_2954);
and UO_99 (O_99,N_2973,N_2941);
and UO_100 (O_100,N_2925,N_2941);
or UO_101 (O_101,N_2959,N_2994);
or UO_102 (O_102,N_2993,N_2937);
and UO_103 (O_103,N_2991,N_2989);
and UO_104 (O_104,N_2942,N_2986);
or UO_105 (O_105,N_2971,N_2959);
nand UO_106 (O_106,N_2974,N_2979);
nor UO_107 (O_107,N_2927,N_2954);
nand UO_108 (O_108,N_2962,N_2931);
and UO_109 (O_109,N_2973,N_2950);
nor UO_110 (O_110,N_2943,N_2991);
and UO_111 (O_111,N_2944,N_2931);
xnor UO_112 (O_112,N_2951,N_2931);
nand UO_113 (O_113,N_2984,N_2926);
nor UO_114 (O_114,N_2931,N_2997);
nor UO_115 (O_115,N_2995,N_2997);
nand UO_116 (O_116,N_2987,N_2960);
xor UO_117 (O_117,N_2928,N_2927);
nand UO_118 (O_118,N_2969,N_2956);
xor UO_119 (O_119,N_2936,N_2942);
xnor UO_120 (O_120,N_2958,N_2953);
and UO_121 (O_121,N_2972,N_2942);
xor UO_122 (O_122,N_2941,N_2949);
nor UO_123 (O_123,N_2996,N_2982);
nand UO_124 (O_124,N_2934,N_2942);
and UO_125 (O_125,N_2956,N_2941);
nor UO_126 (O_126,N_2928,N_2999);
and UO_127 (O_127,N_2974,N_2941);
and UO_128 (O_128,N_2989,N_2940);
nor UO_129 (O_129,N_2934,N_2978);
nor UO_130 (O_130,N_2971,N_2940);
xnor UO_131 (O_131,N_2933,N_2958);
nand UO_132 (O_132,N_2943,N_2998);
xor UO_133 (O_133,N_2934,N_2948);
and UO_134 (O_134,N_2944,N_2997);
or UO_135 (O_135,N_2934,N_2957);
nor UO_136 (O_136,N_2942,N_2991);
or UO_137 (O_137,N_2995,N_2929);
and UO_138 (O_138,N_2991,N_2927);
xnor UO_139 (O_139,N_2973,N_2991);
nand UO_140 (O_140,N_2949,N_2927);
nor UO_141 (O_141,N_2934,N_2965);
or UO_142 (O_142,N_2971,N_2978);
nor UO_143 (O_143,N_2988,N_2985);
nor UO_144 (O_144,N_2967,N_2984);
and UO_145 (O_145,N_2970,N_2990);
or UO_146 (O_146,N_2933,N_2960);
nand UO_147 (O_147,N_2944,N_2980);
nor UO_148 (O_148,N_2933,N_2926);
xor UO_149 (O_149,N_2957,N_2962);
nor UO_150 (O_150,N_2953,N_2965);
nor UO_151 (O_151,N_2945,N_2941);
xnor UO_152 (O_152,N_2935,N_2959);
nand UO_153 (O_153,N_2980,N_2997);
nor UO_154 (O_154,N_2965,N_2966);
nor UO_155 (O_155,N_2959,N_2925);
nand UO_156 (O_156,N_2985,N_2951);
nor UO_157 (O_157,N_2947,N_2989);
nor UO_158 (O_158,N_2933,N_2928);
nor UO_159 (O_159,N_2987,N_2932);
nand UO_160 (O_160,N_2979,N_2948);
or UO_161 (O_161,N_2949,N_2965);
or UO_162 (O_162,N_2932,N_2945);
and UO_163 (O_163,N_2965,N_2937);
and UO_164 (O_164,N_2947,N_2967);
nor UO_165 (O_165,N_2936,N_2947);
nand UO_166 (O_166,N_2981,N_2996);
or UO_167 (O_167,N_2942,N_2965);
xnor UO_168 (O_168,N_2955,N_2946);
and UO_169 (O_169,N_2933,N_2975);
and UO_170 (O_170,N_2995,N_2958);
or UO_171 (O_171,N_2993,N_2951);
nor UO_172 (O_172,N_2950,N_2948);
and UO_173 (O_173,N_2963,N_2928);
or UO_174 (O_174,N_2994,N_2949);
and UO_175 (O_175,N_2939,N_2950);
or UO_176 (O_176,N_2971,N_2993);
and UO_177 (O_177,N_2983,N_2941);
nand UO_178 (O_178,N_2935,N_2949);
xor UO_179 (O_179,N_2926,N_2937);
or UO_180 (O_180,N_2982,N_2962);
or UO_181 (O_181,N_2994,N_2975);
or UO_182 (O_182,N_2929,N_2971);
nand UO_183 (O_183,N_2974,N_2985);
or UO_184 (O_184,N_2973,N_2939);
xor UO_185 (O_185,N_2939,N_2956);
xor UO_186 (O_186,N_2988,N_2999);
nand UO_187 (O_187,N_2977,N_2978);
or UO_188 (O_188,N_2998,N_2938);
or UO_189 (O_189,N_2928,N_2998);
nor UO_190 (O_190,N_2944,N_2928);
and UO_191 (O_191,N_2971,N_2927);
and UO_192 (O_192,N_2961,N_2996);
nor UO_193 (O_193,N_2959,N_2997);
and UO_194 (O_194,N_2966,N_2932);
xnor UO_195 (O_195,N_2959,N_2998);
nor UO_196 (O_196,N_2954,N_2997);
or UO_197 (O_197,N_2999,N_2969);
nor UO_198 (O_198,N_2961,N_2997);
or UO_199 (O_199,N_2937,N_2947);
and UO_200 (O_200,N_2925,N_2966);
and UO_201 (O_201,N_2947,N_2994);
nand UO_202 (O_202,N_2963,N_2943);
xnor UO_203 (O_203,N_2995,N_2962);
nand UO_204 (O_204,N_2996,N_2948);
nand UO_205 (O_205,N_2938,N_2979);
nand UO_206 (O_206,N_2974,N_2926);
nand UO_207 (O_207,N_2956,N_2989);
nor UO_208 (O_208,N_2951,N_2927);
or UO_209 (O_209,N_2979,N_2930);
and UO_210 (O_210,N_2953,N_2943);
nor UO_211 (O_211,N_2943,N_2958);
nor UO_212 (O_212,N_2944,N_2967);
xnor UO_213 (O_213,N_2981,N_2990);
xnor UO_214 (O_214,N_2942,N_2993);
nor UO_215 (O_215,N_2990,N_2953);
nand UO_216 (O_216,N_2954,N_2970);
xnor UO_217 (O_217,N_2951,N_2925);
nand UO_218 (O_218,N_2942,N_2952);
xor UO_219 (O_219,N_2948,N_2997);
xor UO_220 (O_220,N_2934,N_2982);
and UO_221 (O_221,N_2982,N_2943);
or UO_222 (O_222,N_2967,N_2982);
and UO_223 (O_223,N_2952,N_2961);
and UO_224 (O_224,N_2984,N_2992);
nor UO_225 (O_225,N_2990,N_2979);
xnor UO_226 (O_226,N_2927,N_2948);
nand UO_227 (O_227,N_2940,N_2999);
and UO_228 (O_228,N_2970,N_2964);
xnor UO_229 (O_229,N_2996,N_2926);
xor UO_230 (O_230,N_2957,N_2986);
nand UO_231 (O_231,N_2978,N_2938);
and UO_232 (O_232,N_2929,N_2978);
and UO_233 (O_233,N_2958,N_2934);
nand UO_234 (O_234,N_2937,N_2954);
nor UO_235 (O_235,N_2938,N_2946);
nor UO_236 (O_236,N_2939,N_2928);
nand UO_237 (O_237,N_2965,N_2984);
or UO_238 (O_238,N_2928,N_2990);
xnor UO_239 (O_239,N_2925,N_2940);
and UO_240 (O_240,N_2948,N_2939);
and UO_241 (O_241,N_2925,N_2935);
xor UO_242 (O_242,N_2949,N_2999);
and UO_243 (O_243,N_2991,N_2960);
xnor UO_244 (O_244,N_2984,N_2999);
xnor UO_245 (O_245,N_2949,N_2977);
nor UO_246 (O_246,N_2951,N_2982);
nor UO_247 (O_247,N_2994,N_2974);
or UO_248 (O_248,N_2932,N_2934);
nand UO_249 (O_249,N_2959,N_2979);
xnor UO_250 (O_250,N_2967,N_2997);
or UO_251 (O_251,N_2950,N_2947);
xnor UO_252 (O_252,N_2997,N_2957);
and UO_253 (O_253,N_2988,N_2980);
xnor UO_254 (O_254,N_2946,N_2993);
or UO_255 (O_255,N_2943,N_2980);
or UO_256 (O_256,N_2970,N_2934);
nand UO_257 (O_257,N_2951,N_2957);
or UO_258 (O_258,N_2997,N_2969);
xor UO_259 (O_259,N_2957,N_2993);
xnor UO_260 (O_260,N_2954,N_2961);
xor UO_261 (O_261,N_2960,N_2957);
and UO_262 (O_262,N_2986,N_2963);
or UO_263 (O_263,N_2969,N_2974);
xor UO_264 (O_264,N_2999,N_2966);
xnor UO_265 (O_265,N_2998,N_2975);
and UO_266 (O_266,N_2988,N_2975);
and UO_267 (O_267,N_2936,N_2930);
nand UO_268 (O_268,N_2938,N_2991);
xnor UO_269 (O_269,N_2965,N_2970);
or UO_270 (O_270,N_2955,N_2942);
nor UO_271 (O_271,N_2955,N_2976);
and UO_272 (O_272,N_2983,N_2945);
nand UO_273 (O_273,N_2926,N_2936);
and UO_274 (O_274,N_2946,N_2984);
or UO_275 (O_275,N_2934,N_2987);
nand UO_276 (O_276,N_2972,N_2939);
xnor UO_277 (O_277,N_2938,N_2954);
xnor UO_278 (O_278,N_2956,N_2978);
xor UO_279 (O_279,N_2947,N_2952);
and UO_280 (O_280,N_2999,N_2975);
and UO_281 (O_281,N_2968,N_2932);
nor UO_282 (O_282,N_2969,N_2964);
or UO_283 (O_283,N_2937,N_2988);
nand UO_284 (O_284,N_2984,N_2935);
or UO_285 (O_285,N_2965,N_2987);
nand UO_286 (O_286,N_2948,N_2931);
nand UO_287 (O_287,N_2979,N_2954);
and UO_288 (O_288,N_2973,N_2967);
nand UO_289 (O_289,N_2941,N_2943);
or UO_290 (O_290,N_2942,N_2945);
or UO_291 (O_291,N_2955,N_2983);
and UO_292 (O_292,N_2944,N_2982);
nor UO_293 (O_293,N_2940,N_2936);
nor UO_294 (O_294,N_2964,N_2992);
nor UO_295 (O_295,N_2934,N_2997);
and UO_296 (O_296,N_2969,N_2992);
nand UO_297 (O_297,N_2972,N_2946);
or UO_298 (O_298,N_2998,N_2997);
or UO_299 (O_299,N_2966,N_2964);
or UO_300 (O_300,N_2952,N_2953);
nor UO_301 (O_301,N_2933,N_2956);
nor UO_302 (O_302,N_2970,N_2945);
nand UO_303 (O_303,N_2995,N_2938);
and UO_304 (O_304,N_2932,N_2941);
xor UO_305 (O_305,N_2996,N_2944);
and UO_306 (O_306,N_2936,N_2955);
nand UO_307 (O_307,N_2957,N_2936);
nor UO_308 (O_308,N_2930,N_2985);
or UO_309 (O_309,N_2966,N_2996);
and UO_310 (O_310,N_2939,N_2970);
and UO_311 (O_311,N_2992,N_2976);
or UO_312 (O_312,N_2935,N_2988);
and UO_313 (O_313,N_2961,N_2943);
or UO_314 (O_314,N_2991,N_2990);
or UO_315 (O_315,N_2994,N_2991);
nand UO_316 (O_316,N_2991,N_2983);
nand UO_317 (O_317,N_2974,N_2967);
nor UO_318 (O_318,N_2931,N_2955);
and UO_319 (O_319,N_2987,N_2988);
or UO_320 (O_320,N_2957,N_2992);
xor UO_321 (O_321,N_2941,N_2940);
nor UO_322 (O_322,N_2940,N_2990);
and UO_323 (O_323,N_2979,N_2961);
xnor UO_324 (O_324,N_2993,N_2934);
xor UO_325 (O_325,N_2966,N_2988);
or UO_326 (O_326,N_2994,N_2929);
or UO_327 (O_327,N_2940,N_2988);
and UO_328 (O_328,N_2942,N_2938);
xnor UO_329 (O_329,N_2961,N_2930);
xor UO_330 (O_330,N_2977,N_2982);
nand UO_331 (O_331,N_2954,N_2995);
xnor UO_332 (O_332,N_2932,N_2956);
or UO_333 (O_333,N_2950,N_2938);
or UO_334 (O_334,N_2960,N_2929);
xnor UO_335 (O_335,N_2966,N_2946);
and UO_336 (O_336,N_2975,N_2944);
and UO_337 (O_337,N_2947,N_2968);
xor UO_338 (O_338,N_2995,N_2973);
nand UO_339 (O_339,N_2943,N_2974);
nor UO_340 (O_340,N_2995,N_2990);
or UO_341 (O_341,N_2955,N_2925);
xnor UO_342 (O_342,N_2988,N_2932);
and UO_343 (O_343,N_2965,N_2991);
or UO_344 (O_344,N_2995,N_2930);
nand UO_345 (O_345,N_2999,N_2964);
nand UO_346 (O_346,N_2981,N_2999);
and UO_347 (O_347,N_2955,N_2954);
and UO_348 (O_348,N_2965,N_2945);
nor UO_349 (O_349,N_2999,N_2943);
xor UO_350 (O_350,N_2945,N_2950);
xnor UO_351 (O_351,N_2996,N_2958);
nor UO_352 (O_352,N_2979,N_2966);
xor UO_353 (O_353,N_2999,N_2934);
and UO_354 (O_354,N_2983,N_2951);
xor UO_355 (O_355,N_2951,N_2987);
or UO_356 (O_356,N_2944,N_2947);
xnor UO_357 (O_357,N_2998,N_2956);
or UO_358 (O_358,N_2950,N_2971);
nand UO_359 (O_359,N_2974,N_2957);
nand UO_360 (O_360,N_2963,N_2936);
or UO_361 (O_361,N_2959,N_2937);
xnor UO_362 (O_362,N_2988,N_2949);
or UO_363 (O_363,N_2999,N_2960);
and UO_364 (O_364,N_2957,N_2933);
xor UO_365 (O_365,N_2994,N_2943);
or UO_366 (O_366,N_2961,N_2972);
or UO_367 (O_367,N_2994,N_2961);
nor UO_368 (O_368,N_2947,N_2987);
or UO_369 (O_369,N_2984,N_2927);
or UO_370 (O_370,N_2929,N_2987);
xnor UO_371 (O_371,N_2945,N_2943);
or UO_372 (O_372,N_2943,N_2928);
or UO_373 (O_373,N_2960,N_2935);
or UO_374 (O_374,N_2953,N_2973);
xor UO_375 (O_375,N_2995,N_2993);
or UO_376 (O_376,N_2961,N_2944);
or UO_377 (O_377,N_2970,N_2992);
or UO_378 (O_378,N_2968,N_2931);
or UO_379 (O_379,N_2937,N_2953);
and UO_380 (O_380,N_2957,N_2975);
nor UO_381 (O_381,N_2977,N_2975);
and UO_382 (O_382,N_2940,N_2966);
or UO_383 (O_383,N_2966,N_2995);
nand UO_384 (O_384,N_2956,N_2954);
nor UO_385 (O_385,N_2930,N_2993);
nand UO_386 (O_386,N_2928,N_2982);
and UO_387 (O_387,N_2955,N_2953);
and UO_388 (O_388,N_2930,N_2938);
nor UO_389 (O_389,N_2933,N_2953);
nand UO_390 (O_390,N_2966,N_2959);
or UO_391 (O_391,N_2963,N_2982);
or UO_392 (O_392,N_2993,N_2984);
xnor UO_393 (O_393,N_2930,N_2998);
and UO_394 (O_394,N_2956,N_2942);
or UO_395 (O_395,N_2995,N_2985);
and UO_396 (O_396,N_2982,N_2981);
nor UO_397 (O_397,N_2969,N_2932);
or UO_398 (O_398,N_2935,N_2963);
and UO_399 (O_399,N_2941,N_2981);
or UO_400 (O_400,N_2969,N_2945);
or UO_401 (O_401,N_2975,N_2967);
nor UO_402 (O_402,N_2939,N_2998);
and UO_403 (O_403,N_2948,N_2998);
xor UO_404 (O_404,N_2975,N_2954);
and UO_405 (O_405,N_2935,N_2986);
and UO_406 (O_406,N_2947,N_2959);
xnor UO_407 (O_407,N_2927,N_2987);
xnor UO_408 (O_408,N_2942,N_2925);
nand UO_409 (O_409,N_2938,N_2929);
xnor UO_410 (O_410,N_2940,N_2982);
xor UO_411 (O_411,N_2936,N_2972);
or UO_412 (O_412,N_2958,N_2976);
or UO_413 (O_413,N_2985,N_2970);
and UO_414 (O_414,N_2959,N_2976);
nand UO_415 (O_415,N_2969,N_2944);
or UO_416 (O_416,N_2975,N_2973);
or UO_417 (O_417,N_2986,N_2984);
nor UO_418 (O_418,N_2953,N_2975);
nand UO_419 (O_419,N_2993,N_2987);
nand UO_420 (O_420,N_2975,N_2939);
or UO_421 (O_421,N_2962,N_2996);
xnor UO_422 (O_422,N_2940,N_2945);
and UO_423 (O_423,N_2997,N_2937);
xnor UO_424 (O_424,N_2957,N_2925);
or UO_425 (O_425,N_2938,N_2967);
xnor UO_426 (O_426,N_2941,N_2970);
xor UO_427 (O_427,N_2975,N_2986);
nand UO_428 (O_428,N_2996,N_2956);
or UO_429 (O_429,N_2963,N_2961);
or UO_430 (O_430,N_2993,N_2979);
xnor UO_431 (O_431,N_2933,N_2962);
and UO_432 (O_432,N_2950,N_2989);
and UO_433 (O_433,N_2986,N_2992);
nor UO_434 (O_434,N_2946,N_2951);
nor UO_435 (O_435,N_2937,N_2980);
and UO_436 (O_436,N_2932,N_2974);
and UO_437 (O_437,N_2964,N_2933);
or UO_438 (O_438,N_2948,N_2929);
and UO_439 (O_439,N_2992,N_2979);
nor UO_440 (O_440,N_2992,N_2935);
nor UO_441 (O_441,N_2962,N_2949);
nor UO_442 (O_442,N_2967,N_2950);
or UO_443 (O_443,N_2939,N_2932);
xnor UO_444 (O_444,N_2961,N_2982);
nor UO_445 (O_445,N_2938,N_2983);
nand UO_446 (O_446,N_2968,N_2952);
nand UO_447 (O_447,N_2950,N_2981);
nor UO_448 (O_448,N_2993,N_2944);
xnor UO_449 (O_449,N_2967,N_2953);
or UO_450 (O_450,N_2954,N_2933);
xnor UO_451 (O_451,N_2982,N_2988);
xnor UO_452 (O_452,N_2991,N_2948);
nand UO_453 (O_453,N_2931,N_2982);
or UO_454 (O_454,N_2981,N_2949);
nor UO_455 (O_455,N_2925,N_2988);
xnor UO_456 (O_456,N_2950,N_2943);
nor UO_457 (O_457,N_2968,N_2974);
nor UO_458 (O_458,N_2967,N_2961);
or UO_459 (O_459,N_2942,N_2960);
and UO_460 (O_460,N_2960,N_2993);
and UO_461 (O_461,N_2952,N_2991);
or UO_462 (O_462,N_2982,N_2989);
and UO_463 (O_463,N_2964,N_2959);
or UO_464 (O_464,N_2983,N_2943);
xnor UO_465 (O_465,N_2969,N_2947);
nor UO_466 (O_466,N_2945,N_2993);
or UO_467 (O_467,N_2951,N_2974);
nor UO_468 (O_468,N_2930,N_2966);
xor UO_469 (O_469,N_2936,N_2951);
nor UO_470 (O_470,N_2966,N_2973);
nor UO_471 (O_471,N_2947,N_2948);
nand UO_472 (O_472,N_2951,N_2965);
nand UO_473 (O_473,N_2937,N_2961);
xor UO_474 (O_474,N_2942,N_2999);
nor UO_475 (O_475,N_2981,N_2934);
nor UO_476 (O_476,N_2987,N_2985);
or UO_477 (O_477,N_2933,N_2977);
nand UO_478 (O_478,N_2971,N_2944);
nor UO_479 (O_479,N_2955,N_2985);
and UO_480 (O_480,N_2960,N_2977);
and UO_481 (O_481,N_2937,N_2998);
nand UO_482 (O_482,N_2999,N_2927);
or UO_483 (O_483,N_2978,N_2974);
and UO_484 (O_484,N_2967,N_2952);
nor UO_485 (O_485,N_2947,N_2981);
xnor UO_486 (O_486,N_2957,N_2994);
xor UO_487 (O_487,N_2980,N_2977);
nor UO_488 (O_488,N_2927,N_2980);
xor UO_489 (O_489,N_2935,N_2944);
or UO_490 (O_490,N_2995,N_2984);
or UO_491 (O_491,N_2935,N_2990);
xnor UO_492 (O_492,N_2926,N_2986);
xor UO_493 (O_493,N_2992,N_2946);
nand UO_494 (O_494,N_2964,N_2958);
nand UO_495 (O_495,N_2930,N_2941);
nor UO_496 (O_496,N_2969,N_2951);
xnor UO_497 (O_497,N_2941,N_2965);
xor UO_498 (O_498,N_2986,N_2971);
nor UO_499 (O_499,N_2973,N_2985);
endmodule