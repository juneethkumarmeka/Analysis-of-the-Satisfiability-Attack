module basic_500_3000_500_60_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_35,In_251);
nor U1 (N_1,In_357,In_9);
nor U2 (N_2,In_270,In_18);
and U3 (N_3,In_255,In_388);
and U4 (N_4,In_353,In_126);
nor U5 (N_5,In_90,In_33);
nor U6 (N_6,In_27,In_183);
or U7 (N_7,In_247,In_62);
nor U8 (N_8,In_449,In_193);
nand U9 (N_9,In_43,In_291);
or U10 (N_10,In_64,In_222);
xor U11 (N_11,In_82,In_481);
nand U12 (N_12,In_471,In_352);
and U13 (N_13,In_301,In_407);
nand U14 (N_14,In_215,In_25);
nor U15 (N_15,In_414,In_191);
nor U16 (N_16,In_254,In_29);
and U17 (N_17,In_166,In_52);
nand U18 (N_18,In_122,In_311);
or U19 (N_19,In_425,In_487);
or U20 (N_20,In_292,In_171);
nor U21 (N_21,In_63,In_77);
and U22 (N_22,In_307,In_235);
and U23 (N_23,In_323,In_7);
or U24 (N_24,In_361,In_66);
nand U25 (N_25,In_121,In_367);
nand U26 (N_26,In_169,In_279);
or U27 (N_27,In_170,In_34);
nand U28 (N_28,In_368,In_92);
nor U29 (N_29,In_376,In_54);
and U30 (N_30,In_349,In_480);
and U31 (N_31,In_435,In_369);
or U32 (N_32,In_356,In_145);
or U33 (N_33,In_103,In_30);
nand U34 (N_34,In_61,In_46);
nand U35 (N_35,In_19,In_337);
or U36 (N_36,In_115,In_111);
nor U37 (N_37,In_37,In_83);
and U38 (N_38,In_152,In_70);
nand U39 (N_39,In_155,In_58);
nor U40 (N_40,In_236,In_475);
and U41 (N_41,In_49,In_26);
or U42 (N_42,In_326,In_399);
or U43 (N_43,In_14,In_269);
and U44 (N_44,In_226,In_218);
nor U45 (N_45,In_404,In_396);
and U46 (N_46,In_392,In_462);
or U47 (N_47,In_478,In_79);
and U48 (N_48,In_452,In_119);
nand U49 (N_49,In_293,In_335);
nand U50 (N_50,In_24,In_371);
nand U51 (N_51,In_424,In_265);
and U52 (N_52,In_214,In_182);
nand U53 (N_53,In_281,In_477);
or U54 (N_54,In_472,In_428);
nand U55 (N_55,In_243,In_441);
nand U56 (N_56,In_437,N_16);
or U57 (N_57,In_344,In_482);
nor U58 (N_58,In_336,N_1);
nor U59 (N_59,In_302,In_375);
or U60 (N_60,In_387,In_186);
and U61 (N_61,In_467,In_248);
nand U62 (N_62,In_0,N_34);
nor U63 (N_63,In_310,In_355);
nand U64 (N_64,In_76,In_200);
nor U65 (N_65,In_130,In_59);
nor U66 (N_66,In_474,N_24);
or U67 (N_67,In_296,In_363);
or U68 (N_68,In_411,In_149);
nand U69 (N_69,In_427,N_18);
nand U70 (N_70,In_391,In_284);
nand U71 (N_71,In_495,In_57);
nand U72 (N_72,In_250,In_362);
nand U73 (N_73,In_298,In_370);
nor U74 (N_74,In_499,In_458);
and U75 (N_75,N_45,In_436);
nor U76 (N_76,In_394,N_11);
nor U77 (N_77,In_490,In_60);
nor U78 (N_78,In_319,In_275);
nor U79 (N_79,In_460,In_295);
or U80 (N_80,In_91,In_348);
xnor U81 (N_81,In_238,N_37);
nor U82 (N_82,In_290,In_160);
nor U83 (N_83,In_180,In_98);
and U84 (N_84,In_211,In_213);
or U85 (N_85,In_317,In_315);
nor U86 (N_86,In_448,In_93);
nand U87 (N_87,In_492,In_413);
nor U88 (N_88,In_320,In_278);
nor U89 (N_89,In_306,N_35);
nor U90 (N_90,In_162,In_453);
or U91 (N_91,In_339,In_38);
nand U92 (N_92,In_331,In_354);
or U93 (N_93,In_419,In_245);
nand U94 (N_94,In_165,In_114);
nor U95 (N_95,In_393,In_268);
and U96 (N_96,In_283,In_260);
nand U97 (N_97,N_15,In_289);
nand U98 (N_98,In_264,In_410);
nand U99 (N_99,In_68,N_7);
nor U100 (N_100,In_11,N_74);
nor U101 (N_101,N_73,N_77);
nor U102 (N_102,In_282,N_46);
or U103 (N_103,N_75,In_343);
and U104 (N_104,In_409,In_347);
or U105 (N_105,In_172,In_173);
and U106 (N_106,In_135,In_443);
and U107 (N_107,N_90,In_16);
and U108 (N_108,In_242,In_48);
or U109 (N_109,In_325,In_280);
xnor U110 (N_110,N_89,In_234);
nand U111 (N_111,In_142,N_97);
nor U112 (N_112,N_5,In_434);
or U113 (N_113,In_256,In_198);
or U114 (N_114,In_39,In_131);
nand U115 (N_115,In_440,In_322);
or U116 (N_116,In_312,In_384);
or U117 (N_117,In_288,In_318);
nand U118 (N_118,In_316,In_266);
nor U119 (N_119,In_476,In_415);
nand U120 (N_120,N_86,In_333);
nor U121 (N_121,In_395,N_19);
or U122 (N_122,In_385,In_176);
nand U123 (N_123,In_273,In_469);
or U124 (N_124,In_21,N_87);
nor U125 (N_125,In_456,In_313);
or U126 (N_126,In_342,In_13);
xor U127 (N_127,In_194,In_377);
and U128 (N_128,N_81,In_12);
nand U129 (N_129,In_457,In_340);
and U130 (N_130,In_168,In_154);
nor U131 (N_131,In_22,N_2);
or U132 (N_132,In_3,In_398);
or U133 (N_133,N_50,In_96);
nand U134 (N_134,In_277,In_224);
nand U135 (N_135,In_229,N_99);
or U136 (N_136,N_96,In_258);
or U137 (N_137,In_41,In_286);
nor U138 (N_138,In_403,In_178);
and U139 (N_139,N_61,In_167);
and U140 (N_140,In_8,In_221);
or U141 (N_141,In_459,In_105);
and U142 (N_142,In_416,In_207);
nand U143 (N_143,N_25,N_9);
and U144 (N_144,In_137,In_406);
nand U145 (N_145,N_68,N_91);
or U146 (N_146,In_204,In_464);
or U147 (N_147,In_496,In_153);
or U148 (N_148,N_8,In_146);
and U149 (N_149,In_484,N_49);
nor U150 (N_150,In_455,In_350);
and U151 (N_151,In_321,In_144);
nor U152 (N_152,In_241,N_105);
nand U153 (N_153,N_78,N_63);
nor U154 (N_154,In_240,In_157);
or U155 (N_155,N_98,N_116);
or U156 (N_156,In_116,N_148);
or U157 (N_157,In_239,N_129);
nand U158 (N_158,In_175,N_149);
nor U159 (N_159,In_5,N_64);
nand U160 (N_160,N_136,In_237);
and U161 (N_161,N_102,In_461);
and U162 (N_162,N_145,In_212);
nand U163 (N_163,In_303,In_179);
nor U164 (N_164,In_23,In_216);
nor U165 (N_165,N_126,In_285);
and U166 (N_166,N_32,In_104);
nand U167 (N_167,N_95,N_0);
nand U168 (N_168,N_72,N_62);
nand U169 (N_169,In_421,In_341);
nor U170 (N_170,N_69,In_328);
or U171 (N_171,N_33,N_54);
nand U172 (N_172,In_386,N_121);
nor U173 (N_173,In_101,In_156);
nand U174 (N_174,In_489,In_118);
xnor U175 (N_175,N_39,In_4);
and U176 (N_176,In_379,N_142);
nand U177 (N_177,In_259,In_364);
nand U178 (N_178,In_220,In_15);
nand U179 (N_179,In_205,N_14);
and U180 (N_180,In_89,N_135);
and U181 (N_181,N_23,In_124);
nand U182 (N_182,In_99,In_181);
nor U183 (N_183,N_144,In_188);
or U184 (N_184,In_51,In_494);
or U185 (N_185,N_125,In_465);
nor U186 (N_186,N_70,N_103);
or U187 (N_187,In_232,In_345);
or U188 (N_188,N_141,N_130);
and U189 (N_189,In_473,N_71);
xnor U190 (N_190,N_36,In_108);
nand U191 (N_191,In_133,In_327);
or U192 (N_192,In_246,In_113);
nand U193 (N_193,In_109,In_69);
and U194 (N_194,In_73,In_334);
nor U195 (N_195,N_52,In_192);
or U196 (N_196,N_85,N_10);
and U197 (N_197,In_134,N_104);
nand U198 (N_198,In_405,In_147);
or U199 (N_199,In_78,N_30);
or U200 (N_200,In_252,N_140);
and U201 (N_201,In_380,N_146);
and U202 (N_202,N_17,N_185);
and U203 (N_203,In_366,In_201);
and U204 (N_204,N_76,In_117);
or U205 (N_205,In_365,In_120);
and U206 (N_206,In_2,N_13);
nand U207 (N_207,N_177,N_107);
and U208 (N_208,In_329,N_26);
nand U209 (N_209,In_88,In_87);
nand U210 (N_210,N_12,In_136);
or U211 (N_211,In_276,In_378);
nor U212 (N_212,N_139,In_227);
nor U213 (N_213,In_206,N_199);
nor U214 (N_214,N_186,N_172);
and U215 (N_215,N_128,N_183);
and U216 (N_216,N_115,In_418);
or U217 (N_217,In_438,In_140);
nor U218 (N_218,N_188,In_44);
or U219 (N_219,N_154,In_223);
and U220 (N_220,N_40,In_497);
and U221 (N_221,In_479,In_228);
and U222 (N_222,In_219,In_129);
or U223 (N_223,In_300,In_360);
nand U224 (N_224,In_97,In_138);
or U225 (N_225,N_159,In_148);
nand U226 (N_226,In_84,In_485);
nand U227 (N_227,In_422,In_50);
or U228 (N_228,In_304,In_100);
or U229 (N_229,N_184,In_81);
or U230 (N_230,In_257,In_493);
nor U231 (N_231,In_95,N_127);
or U232 (N_232,In_470,In_151);
nor U233 (N_233,N_80,In_208);
and U234 (N_234,In_47,N_117);
or U235 (N_235,N_41,N_38);
and U236 (N_236,In_28,In_486);
and U237 (N_237,In_209,N_176);
and U238 (N_238,N_22,N_51);
nand U239 (N_239,N_189,In_190);
or U240 (N_240,In_324,In_445);
or U241 (N_241,In_230,In_261);
and U242 (N_242,N_28,In_491);
or U243 (N_243,N_181,In_346);
or U244 (N_244,N_124,N_173);
nor U245 (N_245,N_158,In_463);
nand U246 (N_246,In_139,N_113);
nand U247 (N_247,N_170,In_444);
and U248 (N_248,N_58,In_483);
or U249 (N_249,N_166,N_155);
or U250 (N_250,N_27,N_137);
or U251 (N_251,In_225,N_67);
xnor U252 (N_252,N_232,In_125);
and U253 (N_253,In_299,N_92);
nand U254 (N_254,N_100,In_432);
or U255 (N_255,N_48,In_309);
or U256 (N_256,In_210,N_60);
or U257 (N_257,In_159,In_203);
or U258 (N_258,N_204,In_372);
and U259 (N_259,N_198,In_294);
or U260 (N_260,N_4,N_168);
nor U261 (N_261,N_182,N_157);
nor U262 (N_262,N_209,In_158);
and U263 (N_263,N_163,In_196);
or U264 (N_264,N_245,In_127);
nor U265 (N_265,N_122,N_147);
or U266 (N_266,In_451,N_150);
or U267 (N_267,N_203,In_86);
or U268 (N_268,In_20,N_165);
nand U269 (N_269,N_47,In_429);
and U270 (N_270,In_263,In_297);
and U271 (N_271,N_195,In_233);
nor U272 (N_272,In_253,In_488);
or U273 (N_273,In_31,In_106);
xor U274 (N_274,In_163,In_189);
nand U275 (N_275,N_153,In_80);
nor U276 (N_276,N_21,In_217);
or U277 (N_277,N_242,N_57);
or U278 (N_278,N_119,In_272);
or U279 (N_279,In_195,In_132);
nor U280 (N_280,In_314,In_454);
nand U281 (N_281,N_240,N_132);
nand U282 (N_282,In_267,N_218);
or U283 (N_283,N_201,In_32);
nor U284 (N_284,N_123,N_179);
and U285 (N_285,In_143,In_164);
nand U286 (N_286,N_221,N_215);
and U287 (N_287,N_217,In_231);
and U288 (N_288,In_1,N_167);
nand U289 (N_289,In_358,N_223);
nand U290 (N_290,In_197,In_374);
nor U291 (N_291,N_233,In_262);
or U292 (N_292,In_412,N_212);
or U293 (N_293,N_202,In_184);
and U294 (N_294,N_214,N_227);
and U295 (N_295,In_401,In_433);
nor U296 (N_296,In_468,N_224);
or U297 (N_297,N_55,In_67);
and U298 (N_298,N_190,In_426);
nand U299 (N_299,In_10,N_120);
nand U300 (N_300,N_269,In_107);
and U301 (N_301,In_85,N_29);
or U302 (N_302,In_271,N_205);
and U303 (N_303,In_308,In_161);
or U304 (N_304,N_280,N_156);
and U305 (N_305,N_281,In_417);
nand U306 (N_306,N_275,N_261);
or U307 (N_307,N_152,N_151);
or U308 (N_308,N_110,In_373);
or U309 (N_309,N_171,In_498);
nand U310 (N_310,N_108,N_222);
and U311 (N_311,N_162,N_265);
nand U312 (N_312,N_208,N_274);
nand U313 (N_313,N_270,N_93);
and U314 (N_314,In_72,N_262);
and U315 (N_315,In_110,N_279);
nand U316 (N_316,In_408,N_295);
or U317 (N_317,N_289,N_79);
and U318 (N_318,N_138,In_150);
or U319 (N_319,N_213,In_141);
and U320 (N_320,N_109,N_247);
and U321 (N_321,In_185,N_299);
nor U322 (N_322,In_123,N_246);
and U323 (N_323,N_294,N_255);
nand U324 (N_324,N_206,In_74);
nand U325 (N_325,In_56,N_239);
xor U326 (N_326,N_219,In_359);
nand U327 (N_327,N_200,N_106);
and U328 (N_328,In_244,N_134);
or U329 (N_329,N_286,N_293);
nor U330 (N_330,N_263,In_442);
nor U331 (N_331,N_220,N_161);
or U332 (N_332,In_450,In_6);
or U333 (N_333,In_45,N_44);
nor U334 (N_334,In_397,N_131);
nor U335 (N_335,In_466,In_447);
and U336 (N_336,In_389,N_277);
xnor U337 (N_337,N_252,N_288);
or U338 (N_338,N_118,N_266);
or U339 (N_339,N_187,In_42);
nand U340 (N_340,N_175,N_160);
nand U341 (N_341,In_102,N_114);
and U342 (N_342,N_291,N_236);
or U343 (N_343,In_330,In_332);
and U344 (N_344,In_439,N_231);
or U345 (N_345,N_143,N_268);
nor U346 (N_346,In_17,N_282);
nand U347 (N_347,N_241,In_128);
nor U348 (N_348,In_65,In_305);
nand U349 (N_349,In_390,In_383);
nand U350 (N_350,N_348,N_178);
nor U351 (N_351,N_340,N_257);
nor U352 (N_352,N_344,N_31);
nor U353 (N_353,N_260,N_133);
or U354 (N_354,N_250,N_88);
nor U355 (N_355,N_328,N_243);
or U356 (N_356,N_301,N_66);
or U357 (N_357,N_307,N_229);
nor U358 (N_358,N_322,N_326);
and U359 (N_359,N_272,N_194);
nand U360 (N_360,N_287,In_174);
nor U361 (N_361,N_207,N_6);
nand U362 (N_362,N_53,N_169);
nand U363 (N_363,N_325,N_311);
or U364 (N_364,N_82,N_228);
and U365 (N_365,In_446,In_400);
nand U366 (N_366,N_235,N_341);
and U367 (N_367,N_284,N_290);
nor U368 (N_368,N_237,In_382);
and U369 (N_369,N_56,N_337);
or U370 (N_370,N_59,N_347);
nor U371 (N_371,N_310,N_336);
nand U372 (N_372,N_258,In_381);
nor U373 (N_373,N_343,N_327);
nand U374 (N_374,In_177,In_112);
nor U375 (N_375,N_278,N_312);
and U376 (N_376,N_285,N_321);
or U377 (N_377,N_248,N_94);
nor U378 (N_378,N_346,N_300);
nor U379 (N_379,In_55,In_431);
and U380 (N_380,In_338,N_324);
nand U381 (N_381,In_40,N_254);
or U382 (N_382,In_71,N_308);
nor U383 (N_383,In_187,N_234);
or U384 (N_384,N_238,N_244);
nand U385 (N_385,In_36,N_334);
nand U386 (N_386,N_332,N_319);
and U387 (N_387,N_43,In_94);
nor U388 (N_388,N_314,N_256);
or U389 (N_389,In_287,In_274);
nand U390 (N_390,N_349,N_329);
and U391 (N_391,N_320,N_292);
nor U392 (N_392,N_342,N_316);
nor U393 (N_393,In_351,N_230);
and U394 (N_394,N_112,N_226);
and U395 (N_395,N_297,N_111);
or U396 (N_396,N_216,In_202);
nand U397 (N_397,N_303,In_199);
nor U398 (N_398,N_315,N_264);
and U399 (N_399,N_164,N_271);
nor U400 (N_400,N_251,In_420);
and U401 (N_401,N_372,N_42);
nor U402 (N_402,N_358,In_75);
and U403 (N_403,N_65,N_389);
and U404 (N_404,N_225,N_197);
and U405 (N_405,N_335,N_374);
or U406 (N_406,N_354,N_353);
nor U407 (N_407,In_402,N_318);
or U408 (N_408,In_53,N_399);
nand U409 (N_409,N_373,N_330);
nand U410 (N_410,N_383,N_196);
xnor U411 (N_411,N_362,N_305);
nand U412 (N_412,N_364,N_317);
xor U413 (N_413,N_369,N_352);
nor U414 (N_414,N_376,N_339);
or U415 (N_415,N_385,N_302);
and U416 (N_416,N_396,N_345);
nor U417 (N_417,N_360,N_382);
nand U418 (N_418,N_386,N_367);
and U419 (N_419,N_180,N_366);
and U420 (N_420,N_333,N_391);
and U421 (N_421,N_381,N_192);
nand U422 (N_422,N_101,N_378);
or U423 (N_423,N_283,N_313);
nor U424 (N_424,N_377,N_84);
or U425 (N_425,N_331,N_375);
or U426 (N_426,N_191,N_253);
or U427 (N_427,N_276,N_361);
and U428 (N_428,N_363,N_397);
or U429 (N_429,N_296,N_83);
nor U430 (N_430,N_394,N_371);
nand U431 (N_431,N_384,N_249);
nor U432 (N_432,In_430,N_387);
nor U433 (N_433,N_174,N_359);
or U434 (N_434,N_338,N_210);
nor U435 (N_435,N_390,N_350);
nor U436 (N_436,N_267,N_259);
or U437 (N_437,N_392,N_365);
and U438 (N_438,N_304,N_323);
and U439 (N_439,N_298,N_273);
nor U440 (N_440,N_393,N_193);
nand U441 (N_441,N_379,N_370);
or U442 (N_442,N_356,N_306);
and U443 (N_443,N_380,N_398);
nor U444 (N_444,N_211,In_423);
and U445 (N_445,N_309,N_357);
and U446 (N_446,In_249,N_395);
or U447 (N_447,N_368,N_20);
and U448 (N_448,N_355,N_351);
or U449 (N_449,N_388,N_3);
nor U450 (N_450,N_424,N_401);
or U451 (N_451,N_431,N_403);
and U452 (N_452,N_404,N_409);
and U453 (N_453,N_430,N_432);
or U454 (N_454,N_446,N_405);
and U455 (N_455,N_443,N_437);
nor U456 (N_456,N_433,N_414);
nor U457 (N_457,N_442,N_400);
nand U458 (N_458,N_428,N_422);
or U459 (N_459,N_415,N_439);
and U460 (N_460,N_418,N_423);
nand U461 (N_461,N_426,N_448);
nor U462 (N_462,N_402,N_412);
nor U463 (N_463,N_425,N_436);
nand U464 (N_464,N_419,N_434);
and U465 (N_465,N_417,N_441);
nand U466 (N_466,N_444,N_413);
nor U467 (N_467,N_410,N_408);
nor U468 (N_468,N_445,N_407);
nor U469 (N_469,N_435,N_429);
nand U470 (N_470,N_421,N_420);
nor U471 (N_471,N_411,N_438);
and U472 (N_472,N_406,N_440);
xor U473 (N_473,N_447,N_416);
and U474 (N_474,N_449,N_427);
and U475 (N_475,N_419,N_447);
or U476 (N_476,N_419,N_412);
and U477 (N_477,N_441,N_429);
or U478 (N_478,N_402,N_417);
nor U479 (N_479,N_412,N_437);
or U480 (N_480,N_411,N_432);
or U481 (N_481,N_423,N_446);
or U482 (N_482,N_405,N_439);
and U483 (N_483,N_400,N_430);
xnor U484 (N_484,N_403,N_418);
nand U485 (N_485,N_447,N_432);
nand U486 (N_486,N_428,N_448);
nand U487 (N_487,N_427,N_407);
and U488 (N_488,N_432,N_416);
and U489 (N_489,N_410,N_414);
nor U490 (N_490,N_416,N_417);
or U491 (N_491,N_448,N_444);
xor U492 (N_492,N_407,N_419);
and U493 (N_493,N_414,N_443);
and U494 (N_494,N_429,N_414);
nor U495 (N_495,N_441,N_440);
or U496 (N_496,N_425,N_417);
nand U497 (N_497,N_403,N_410);
nor U498 (N_498,N_416,N_446);
nand U499 (N_499,N_435,N_422);
or U500 (N_500,N_456,N_497);
or U501 (N_501,N_451,N_461);
or U502 (N_502,N_489,N_494);
or U503 (N_503,N_466,N_457);
and U504 (N_504,N_499,N_477);
nand U505 (N_505,N_458,N_485);
nor U506 (N_506,N_479,N_488);
xnor U507 (N_507,N_453,N_468);
nor U508 (N_508,N_459,N_474);
nand U509 (N_509,N_470,N_476);
nor U510 (N_510,N_464,N_465);
nor U511 (N_511,N_455,N_486);
nor U512 (N_512,N_472,N_473);
and U513 (N_513,N_463,N_460);
nor U514 (N_514,N_491,N_469);
or U515 (N_515,N_483,N_493);
nor U516 (N_516,N_496,N_475);
and U517 (N_517,N_484,N_487);
nor U518 (N_518,N_462,N_498);
nand U519 (N_519,N_471,N_490);
and U520 (N_520,N_450,N_482);
nor U521 (N_521,N_478,N_495);
nor U522 (N_522,N_481,N_467);
nor U523 (N_523,N_492,N_452);
nand U524 (N_524,N_480,N_454);
nand U525 (N_525,N_471,N_479);
and U526 (N_526,N_468,N_499);
or U527 (N_527,N_466,N_493);
or U528 (N_528,N_485,N_497);
and U529 (N_529,N_457,N_464);
nor U530 (N_530,N_486,N_483);
nand U531 (N_531,N_488,N_497);
and U532 (N_532,N_459,N_489);
and U533 (N_533,N_484,N_479);
and U534 (N_534,N_467,N_456);
or U535 (N_535,N_451,N_458);
nor U536 (N_536,N_498,N_453);
nand U537 (N_537,N_451,N_466);
nor U538 (N_538,N_468,N_484);
nand U539 (N_539,N_467,N_492);
nand U540 (N_540,N_462,N_456);
or U541 (N_541,N_480,N_485);
and U542 (N_542,N_489,N_490);
and U543 (N_543,N_455,N_469);
nand U544 (N_544,N_458,N_480);
xor U545 (N_545,N_499,N_495);
nand U546 (N_546,N_497,N_474);
nand U547 (N_547,N_494,N_467);
nor U548 (N_548,N_478,N_455);
nor U549 (N_549,N_455,N_457);
and U550 (N_550,N_527,N_545);
and U551 (N_551,N_503,N_524);
nor U552 (N_552,N_521,N_514);
nor U553 (N_553,N_517,N_542);
or U554 (N_554,N_536,N_537);
and U555 (N_555,N_531,N_520);
and U556 (N_556,N_533,N_515);
nand U557 (N_557,N_513,N_509);
or U558 (N_558,N_522,N_504);
and U559 (N_559,N_502,N_511);
nor U560 (N_560,N_506,N_546);
nor U561 (N_561,N_501,N_535);
nand U562 (N_562,N_532,N_500);
nand U563 (N_563,N_507,N_534);
and U564 (N_564,N_510,N_544);
and U565 (N_565,N_538,N_548);
and U566 (N_566,N_526,N_529);
and U567 (N_567,N_519,N_549);
and U568 (N_568,N_516,N_523);
and U569 (N_569,N_540,N_528);
nand U570 (N_570,N_525,N_508);
nand U571 (N_571,N_518,N_505);
and U572 (N_572,N_547,N_543);
or U573 (N_573,N_539,N_512);
and U574 (N_574,N_541,N_530);
nand U575 (N_575,N_512,N_538);
nand U576 (N_576,N_524,N_523);
and U577 (N_577,N_519,N_543);
nand U578 (N_578,N_520,N_543);
nand U579 (N_579,N_512,N_536);
or U580 (N_580,N_542,N_524);
and U581 (N_581,N_510,N_500);
or U582 (N_582,N_529,N_501);
and U583 (N_583,N_502,N_531);
nor U584 (N_584,N_524,N_509);
or U585 (N_585,N_509,N_501);
nor U586 (N_586,N_541,N_527);
and U587 (N_587,N_529,N_518);
nor U588 (N_588,N_512,N_500);
nor U589 (N_589,N_529,N_548);
nand U590 (N_590,N_500,N_541);
nand U591 (N_591,N_546,N_536);
xnor U592 (N_592,N_533,N_527);
nor U593 (N_593,N_540,N_511);
or U594 (N_594,N_512,N_502);
or U595 (N_595,N_511,N_546);
nor U596 (N_596,N_503,N_537);
or U597 (N_597,N_510,N_511);
nor U598 (N_598,N_501,N_531);
nor U599 (N_599,N_518,N_524);
nand U600 (N_600,N_585,N_590);
or U601 (N_601,N_570,N_568);
nor U602 (N_602,N_583,N_567);
or U603 (N_603,N_554,N_576);
or U604 (N_604,N_562,N_595);
and U605 (N_605,N_555,N_592);
nor U606 (N_606,N_574,N_577);
nand U607 (N_607,N_586,N_558);
or U608 (N_608,N_572,N_566);
or U609 (N_609,N_598,N_551);
and U610 (N_610,N_563,N_561);
and U611 (N_611,N_559,N_569);
nand U612 (N_612,N_584,N_591);
nand U613 (N_613,N_552,N_560);
or U614 (N_614,N_553,N_564);
and U615 (N_615,N_571,N_593);
or U616 (N_616,N_582,N_599);
and U617 (N_617,N_578,N_556);
nor U618 (N_618,N_565,N_550);
nor U619 (N_619,N_589,N_594);
nand U620 (N_620,N_588,N_580);
nand U621 (N_621,N_596,N_587);
and U622 (N_622,N_579,N_557);
or U623 (N_623,N_597,N_581);
or U624 (N_624,N_573,N_575);
and U625 (N_625,N_552,N_576);
nand U626 (N_626,N_558,N_577);
nand U627 (N_627,N_588,N_599);
nand U628 (N_628,N_592,N_550);
and U629 (N_629,N_579,N_570);
nand U630 (N_630,N_550,N_589);
nand U631 (N_631,N_582,N_577);
xnor U632 (N_632,N_568,N_560);
or U633 (N_633,N_551,N_571);
or U634 (N_634,N_583,N_552);
nand U635 (N_635,N_586,N_575);
or U636 (N_636,N_555,N_599);
nor U637 (N_637,N_560,N_578);
and U638 (N_638,N_553,N_550);
and U639 (N_639,N_584,N_553);
nand U640 (N_640,N_591,N_555);
nand U641 (N_641,N_598,N_553);
nand U642 (N_642,N_581,N_554);
nor U643 (N_643,N_583,N_580);
or U644 (N_644,N_592,N_581);
or U645 (N_645,N_565,N_595);
xor U646 (N_646,N_577,N_563);
nor U647 (N_647,N_560,N_591);
nand U648 (N_648,N_577,N_565);
nand U649 (N_649,N_590,N_559);
nor U650 (N_650,N_632,N_603);
nor U651 (N_651,N_618,N_604);
or U652 (N_652,N_649,N_602);
and U653 (N_653,N_646,N_620);
nor U654 (N_654,N_623,N_600);
nor U655 (N_655,N_606,N_610);
and U656 (N_656,N_640,N_631);
nand U657 (N_657,N_637,N_641);
or U658 (N_658,N_630,N_607);
nand U659 (N_659,N_621,N_628);
nand U660 (N_660,N_622,N_643);
nor U661 (N_661,N_612,N_634);
and U662 (N_662,N_635,N_636);
nor U663 (N_663,N_645,N_639);
or U664 (N_664,N_609,N_619);
nand U665 (N_665,N_625,N_601);
nor U666 (N_666,N_642,N_611);
nand U667 (N_667,N_627,N_626);
nor U668 (N_668,N_633,N_614);
or U669 (N_669,N_605,N_613);
xnor U670 (N_670,N_616,N_608);
or U671 (N_671,N_647,N_644);
and U672 (N_672,N_629,N_648);
or U673 (N_673,N_615,N_617);
and U674 (N_674,N_624,N_638);
nand U675 (N_675,N_629,N_631);
nand U676 (N_676,N_627,N_639);
nor U677 (N_677,N_613,N_610);
nand U678 (N_678,N_603,N_615);
nand U679 (N_679,N_608,N_648);
or U680 (N_680,N_642,N_627);
nor U681 (N_681,N_616,N_640);
nand U682 (N_682,N_644,N_636);
nand U683 (N_683,N_604,N_634);
nor U684 (N_684,N_626,N_621);
and U685 (N_685,N_645,N_648);
and U686 (N_686,N_608,N_627);
nor U687 (N_687,N_633,N_624);
and U688 (N_688,N_631,N_608);
nand U689 (N_689,N_608,N_623);
and U690 (N_690,N_624,N_611);
xor U691 (N_691,N_629,N_605);
nand U692 (N_692,N_609,N_631);
nand U693 (N_693,N_608,N_602);
or U694 (N_694,N_612,N_645);
xor U695 (N_695,N_604,N_642);
nor U696 (N_696,N_635,N_643);
xor U697 (N_697,N_647,N_639);
and U698 (N_698,N_641,N_601);
or U699 (N_699,N_604,N_640);
nand U700 (N_700,N_672,N_669);
nor U701 (N_701,N_674,N_655);
or U702 (N_702,N_664,N_697);
and U703 (N_703,N_650,N_665);
nand U704 (N_704,N_666,N_660);
and U705 (N_705,N_696,N_698);
xnor U706 (N_706,N_673,N_657);
or U707 (N_707,N_653,N_679);
and U708 (N_708,N_685,N_651);
or U709 (N_709,N_694,N_677);
or U710 (N_710,N_695,N_662);
or U711 (N_711,N_656,N_663);
or U712 (N_712,N_678,N_699);
or U713 (N_713,N_686,N_676);
nand U714 (N_714,N_684,N_659);
or U715 (N_715,N_675,N_680);
or U716 (N_716,N_671,N_681);
nor U717 (N_717,N_692,N_654);
nor U718 (N_718,N_690,N_682);
nand U719 (N_719,N_689,N_683);
nand U720 (N_720,N_658,N_691);
nor U721 (N_721,N_652,N_661);
and U722 (N_722,N_670,N_693);
and U723 (N_723,N_688,N_668);
nand U724 (N_724,N_687,N_667);
nor U725 (N_725,N_675,N_670);
or U726 (N_726,N_650,N_687);
and U727 (N_727,N_654,N_696);
or U728 (N_728,N_694,N_680);
nor U729 (N_729,N_656,N_657);
or U730 (N_730,N_660,N_657);
or U731 (N_731,N_682,N_689);
nand U732 (N_732,N_678,N_687);
nor U733 (N_733,N_673,N_665);
nor U734 (N_734,N_672,N_650);
nor U735 (N_735,N_652,N_697);
nand U736 (N_736,N_680,N_685);
nand U737 (N_737,N_691,N_694);
or U738 (N_738,N_661,N_667);
and U739 (N_739,N_687,N_675);
nor U740 (N_740,N_651,N_668);
nor U741 (N_741,N_660,N_684);
or U742 (N_742,N_674,N_660);
nor U743 (N_743,N_693,N_650);
and U744 (N_744,N_676,N_677);
nand U745 (N_745,N_690,N_662);
or U746 (N_746,N_656,N_682);
nor U747 (N_747,N_689,N_670);
and U748 (N_748,N_685,N_690);
nor U749 (N_749,N_668,N_680);
nor U750 (N_750,N_747,N_718);
or U751 (N_751,N_731,N_723);
nor U752 (N_752,N_725,N_716);
and U753 (N_753,N_733,N_737);
or U754 (N_754,N_705,N_746);
and U755 (N_755,N_744,N_739);
or U756 (N_756,N_710,N_729);
nand U757 (N_757,N_713,N_743);
or U758 (N_758,N_709,N_748);
xor U759 (N_759,N_749,N_724);
nand U760 (N_760,N_728,N_736);
or U761 (N_761,N_726,N_721);
and U762 (N_762,N_732,N_703);
and U763 (N_763,N_708,N_707);
and U764 (N_764,N_740,N_712);
or U765 (N_765,N_734,N_727);
nand U766 (N_766,N_720,N_741);
and U767 (N_767,N_722,N_717);
and U768 (N_768,N_735,N_719);
or U769 (N_769,N_701,N_702);
nor U770 (N_770,N_700,N_738);
nand U771 (N_771,N_704,N_714);
and U772 (N_772,N_730,N_745);
nand U773 (N_773,N_711,N_715);
nand U774 (N_774,N_742,N_706);
nor U775 (N_775,N_722,N_747);
or U776 (N_776,N_718,N_744);
nand U777 (N_777,N_722,N_740);
and U778 (N_778,N_743,N_748);
nor U779 (N_779,N_732,N_714);
and U780 (N_780,N_732,N_711);
nor U781 (N_781,N_711,N_745);
nand U782 (N_782,N_711,N_729);
or U783 (N_783,N_749,N_741);
nand U784 (N_784,N_728,N_714);
nor U785 (N_785,N_705,N_703);
nor U786 (N_786,N_730,N_729);
nand U787 (N_787,N_717,N_705);
nor U788 (N_788,N_717,N_701);
nor U789 (N_789,N_740,N_703);
nand U790 (N_790,N_732,N_717);
and U791 (N_791,N_738,N_735);
or U792 (N_792,N_738,N_736);
or U793 (N_793,N_735,N_716);
and U794 (N_794,N_700,N_737);
or U795 (N_795,N_727,N_717);
nor U796 (N_796,N_710,N_732);
nor U797 (N_797,N_714,N_740);
and U798 (N_798,N_710,N_734);
and U799 (N_799,N_713,N_744);
and U800 (N_800,N_790,N_792);
nor U801 (N_801,N_796,N_769);
or U802 (N_802,N_755,N_768);
nand U803 (N_803,N_783,N_757);
and U804 (N_804,N_763,N_752);
nor U805 (N_805,N_776,N_779);
nand U806 (N_806,N_762,N_764);
and U807 (N_807,N_767,N_785);
or U808 (N_808,N_775,N_766);
or U809 (N_809,N_784,N_750);
or U810 (N_810,N_795,N_791);
or U811 (N_811,N_781,N_778);
or U812 (N_812,N_782,N_794);
xor U813 (N_813,N_789,N_774);
nor U814 (N_814,N_754,N_751);
nor U815 (N_815,N_756,N_780);
and U816 (N_816,N_773,N_777);
or U817 (N_817,N_772,N_787);
or U818 (N_818,N_797,N_760);
or U819 (N_819,N_761,N_753);
or U820 (N_820,N_771,N_793);
and U821 (N_821,N_765,N_759);
nor U822 (N_822,N_786,N_799);
nor U823 (N_823,N_758,N_798);
and U824 (N_824,N_788,N_770);
and U825 (N_825,N_782,N_752);
or U826 (N_826,N_770,N_773);
or U827 (N_827,N_769,N_767);
and U828 (N_828,N_760,N_795);
nor U829 (N_829,N_792,N_761);
nor U830 (N_830,N_792,N_797);
nand U831 (N_831,N_791,N_753);
nand U832 (N_832,N_774,N_777);
nor U833 (N_833,N_798,N_786);
nor U834 (N_834,N_768,N_790);
or U835 (N_835,N_784,N_768);
and U836 (N_836,N_755,N_774);
and U837 (N_837,N_751,N_780);
or U838 (N_838,N_787,N_764);
or U839 (N_839,N_765,N_769);
nand U840 (N_840,N_770,N_793);
nor U841 (N_841,N_798,N_780);
or U842 (N_842,N_774,N_750);
or U843 (N_843,N_767,N_776);
and U844 (N_844,N_783,N_763);
or U845 (N_845,N_757,N_767);
and U846 (N_846,N_777,N_769);
xor U847 (N_847,N_798,N_754);
nand U848 (N_848,N_766,N_767);
nand U849 (N_849,N_791,N_790);
nand U850 (N_850,N_824,N_818);
nand U851 (N_851,N_849,N_846);
nor U852 (N_852,N_813,N_806);
xnor U853 (N_853,N_819,N_834);
and U854 (N_854,N_825,N_838);
nor U855 (N_855,N_839,N_804);
and U856 (N_856,N_830,N_837);
nand U857 (N_857,N_814,N_842);
and U858 (N_858,N_815,N_843);
nand U859 (N_859,N_816,N_840);
or U860 (N_860,N_822,N_800);
or U861 (N_861,N_832,N_848);
or U862 (N_862,N_828,N_812);
nand U863 (N_863,N_831,N_841);
nand U864 (N_864,N_836,N_829);
nor U865 (N_865,N_809,N_844);
nand U866 (N_866,N_835,N_802);
and U867 (N_867,N_805,N_801);
or U868 (N_868,N_827,N_810);
nor U869 (N_869,N_811,N_821);
nor U870 (N_870,N_847,N_808);
and U871 (N_871,N_820,N_817);
and U872 (N_872,N_826,N_823);
and U873 (N_873,N_807,N_803);
nand U874 (N_874,N_845,N_833);
nor U875 (N_875,N_817,N_839);
nor U876 (N_876,N_808,N_843);
or U877 (N_877,N_824,N_816);
or U878 (N_878,N_805,N_827);
and U879 (N_879,N_849,N_845);
nor U880 (N_880,N_821,N_835);
and U881 (N_881,N_817,N_840);
or U882 (N_882,N_808,N_831);
nand U883 (N_883,N_836,N_803);
or U884 (N_884,N_813,N_819);
nor U885 (N_885,N_822,N_817);
nor U886 (N_886,N_840,N_805);
or U887 (N_887,N_808,N_810);
and U888 (N_888,N_809,N_800);
and U889 (N_889,N_845,N_817);
and U890 (N_890,N_843,N_845);
xnor U891 (N_891,N_831,N_840);
nand U892 (N_892,N_811,N_810);
or U893 (N_893,N_815,N_844);
and U894 (N_894,N_820,N_814);
xnor U895 (N_895,N_802,N_829);
or U896 (N_896,N_817,N_849);
or U897 (N_897,N_814,N_826);
nor U898 (N_898,N_817,N_805);
nand U899 (N_899,N_829,N_820);
or U900 (N_900,N_868,N_898);
and U901 (N_901,N_874,N_860);
or U902 (N_902,N_878,N_889);
xor U903 (N_903,N_873,N_852);
nand U904 (N_904,N_856,N_854);
nand U905 (N_905,N_876,N_851);
and U906 (N_906,N_885,N_853);
xnor U907 (N_907,N_867,N_869);
nor U908 (N_908,N_891,N_880);
nand U909 (N_909,N_897,N_872);
nand U910 (N_910,N_875,N_855);
nor U911 (N_911,N_882,N_879);
nor U912 (N_912,N_857,N_896);
nand U913 (N_913,N_864,N_859);
nand U914 (N_914,N_892,N_893);
nand U915 (N_915,N_850,N_884);
xor U916 (N_916,N_883,N_894);
and U917 (N_917,N_890,N_888);
or U918 (N_918,N_871,N_887);
nand U919 (N_919,N_865,N_895);
or U920 (N_920,N_866,N_886);
xor U921 (N_921,N_881,N_870);
or U922 (N_922,N_877,N_862);
nand U923 (N_923,N_899,N_863);
nand U924 (N_924,N_861,N_858);
or U925 (N_925,N_882,N_869);
nand U926 (N_926,N_886,N_856);
nor U927 (N_927,N_890,N_858);
nand U928 (N_928,N_888,N_858);
nand U929 (N_929,N_863,N_894);
nand U930 (N_930,N_881,N_863);
nor U931 (N_931,N_863,N_875);
nand U932 (N_932,N_898,N_860);
and U933 (N_933,N_861,N_864);
and U934 (N_934,N_899,N_851);
and U935 (N_935,N_892,N_861);
and U936 (N_936,N_896,N_852);
xnor U937 (N_937,N_881,N_878);
nand U938 (N_938,N_860,N_895);
or U939 (N_939,N_896,N_862);
or U940 (N_940,N_895,N_879);
nor U941 (N_941,N_852,N_886);
nand U942 (N_942,N_872,N_899);
nor U943 (N_943,N_878,N_865);
nor U944 (N_944,N_866,N_894);
or U945 (N_945,N_874,N_857);
xor U946 (N_946,N_860,N_859);
nand U947 (N_947,N_862,N_880);
nand U948 (N_948,N_865,N_867);
nand U949 (N_949,N_897,N_886);
nand U950 (N_950,N_905,N_926);
or U951 (N_951,N_921,N_910);
or U952 (N_952,N_919,N_918);
or U953 (N_953,N_920,N_936);
or U954 (N_954,N_931,N_914);
and U955 (N_955,N_906,N_938);
nand U956 (N_956,N_913,N_916);
and U957 (N_957,N_923,N_929);
or U958 (N_958,N_903,N_909);
nand U959 (N_959,N_922,N_901);
nand U960 (N_960,N_934,N_930);
nand U961 (N_961,N_935,N_900);
and U962 (N_962,N_902,N_949);
nand U963 (N_963,N_915,N_933);
or U964 (N_964,N_924,N_932);
nand U965 (N_965,N_917,N_908);
and U966 (N_966,N_942,N_928);
nand U967 (N_967,N_946,N_911);
or U968 (N_968,N_945,N_904);
or U969 (N_969,N_939,N_947);
and U970 (N_970,N_927,N_912);
and U971 (N_971,N_948,N_937);
and U972 (N_972,N_943,N_907);
nor U973 (N_973,N_940,N_941);
and U974 (N_974,N_944,N_925);
and U975 (N_975,N_924,N_943);
nor U976 (N_976,N_920,N_906);
nor U977 (N_977,N_926,N_942);
or U978 (N_978,N_940,N_938);
nand U979 (N_979,N_918,N_934);
nand U980 (N_980,N_936,N_901);
nor U981 (N_981,N_934,N_914);
and U982 (N_982,N_946,N_932);
and U983 (N_983,N_920,N_921);
nand U984 (N_984,N_939,N_937);
and U985 (N_985,N_948,N_939);
nand U986 (N_986,N_945,N_947);
or U987 (N_987,N_928,N_946);
or U988 (N_988,N_902,N_947);
or U989 (N_989,N_916,N_931);
nand U990 (N_990,N_905,N_903);
nor U991 (N_991,N_932,N_945);
or U992 (N_992,N_913,N_927);
and U993 (N_993,N_911,N_922);
nor U994 (N_994,N_915,N_936);
and U995 (N_995,N_949,N_919);
nor U996 (N_996,N_901,N_916);
nand U997 (N_997,N_904,N_906);
or U998 (N_998,N_940,N_904);
and U999 (N_999,N_922,N_903);
or U1000 (N_1000,N_988,N_990);
or U1001 (N_1001,N_989,N_966);
or U1002 (N_1002,N_972,N_977);
nand U1003 (N_1003,N_969,N_950);
nor U1004 (N_1004,N_964,N_974);
nand U1005 (N_1005,N_962,N_959);
or U1006 (N_1006,N_981,N_960);
or U1007 (N_1007,N_982,N_963);
or U1008 (N_1008,N_954,N_958);
or U1009 (N_1009,N_951,N_952);
and U1010 (N_1010,N_967,N_993);
nor U1011 (N_1011,N_985,N_961);
and U1012 (N_1012,N_973,N_965);
nand U1013 (N_1013,N_976,N_991);
nor U1014 (N_1014,N_979,N_998);
nor U1015 (N_1015,N_999,N_994);
nand U1016 (N_1016,N_996,N_983);
nand U1017 (N_1017,N_986,N_957);
nor U1018 (N_1018,N_978,N_953);
nor U1019 (N_1019,N_987,N_971);
nand U1020 (N_1020,N_970,N_968);
nor U1021 (N_1021,N_997,N_980);
nor U1022 (N_1022,N_956,N_984);
nor U1023 (N_1023,N_992,N_975);
and U1024 (N_1024,N_995,N_955);
nand U1025 (N_1025,N_990,N_956);
and U1026 (N_1026,N_958,N_965);
and U1027 (N_1027,N_993,N_959);
nor U1028 (N_1028,N_965,N_954);
nor U1029 (N_1029,N_989,N_993);
or U1030 (N_1030,N_956,N_962);
nor U1031 (N_1031,N_967,N_976);
and U1032 (N_1032,N_954,N_963);
nand U1033 (N_1033,N_961,N_954);
nand U1034 (N_1034,N_967,N_999);
and U1035 (N_1035,N_971,N_959);
or U1036 (N_1036,N_967,N_968);
nand U1037 (N_1037,N_992,N_953);
nand U1038 (N_1038,N_960,N_961);
and U1039 (N_1039,N_991,N_982);
nor U1040 (N_1040,N_953,N_966);
or U1041 (N_1041,N_988,N_998);
nand U1042 (N_1042,N_998,N_954);
or U1043 (N_1043,N_964,N_963);
and U1044 (N_1044,N_986,N_955);
nor U1045 (N_1045,N_970,N_993);
or U1046 (N_1046,N_967,N_982);
nand U1047 (N_1047,N_992,N_960);
nand U1048 (N_1048,N_972,N_995);
nor U1049 (N_1049,N_995,N_987);
nor U1050 (N_1050,N_1036,N_1008);
or U1051 (N_1051,N_1019,N_1022);
and U1052 (N_1052,N_1035,N_1018);
xor U1053 (N_1053,N_1009,N_1042);
and U1054 (N_1054,N_1031,N_1028);
or U1055 (N_1055,N_1040,N_1046);
and U1056 (N_1056,N_1010,N_1025);
nor U1057 (N_1057,N_1016,N_1000);
nor U1058 (N_1058,N_1004,N_1014);
and U1059 (N_1059,N_1015,N_1020);
and U1060 (N_1060,N_1002,N_1024);
nand U1061 (N_1061,N_1048,N_1013);
nand U1062 (N_1062,N_1001,N_1041);
and U1063 (N_1063,N_1047,N_1027);
or U1064 (N_1064,N_1045,N_1044);
or U1065 (N_1065,N_1007,N_1049);
and U1066 (N_1066,N_1043,N_1003);
and U1067 (N_1067,N_1030,N_1034);
and U1068 (N_1068,N_1037,N_1005);
xnor U1069 (N_1069,N_1011,N_1017);
nor U1070 (N_1070,N_1026,N_1029);
nor U1071 (N_1071,N_1032,N_1033);
or U1072 (N_1072,N_1039,N_1006);
nand U1073 (N_1073,N_1012,N_1038);
or U1074 (N_1074,N_1023,N_1021);
nor U1075 (N_1075,N_1006,N_1005);
nor U1076 (N_1076,N_1007,N_1006);
nand U1077 (N_1077,N_1015,N_1021);
or U1078 (N_1078,N_1041,N_1037);
nand U1079 (N_1079,N_1043,N_1012);
nor U1080 (N_1080,N_1008,N_1046);
nand U1081 (N_1081,N_1047,N_1015);
or U1082 (N_1082,N_1010,N_1019);
nand U1083 (N_1083,N_1009,N_1039);
nor U1084 (N_1084,N_1026,N_1012);
nor U1085 (N_1085,N_1006,N_1049);
nor U1086 (N_1086,N_1007,N_1037);
nor U1087 (N_1087,N_1033,N_1004);
xnor U1088 (N_1088,N_1016,N_1006);
and U1089 (N_1089,N_1028,N_1012);
and U1090 (N_1090,N_1044,N_1021);
nor U1091 (N_1091,N_1017,N_1013);
and U1092 (N_1092,N_1045,N_1047);
nand U1093 (N_1093,N_1034,N_1022);
and U1094 (N_1094,N_1044,N_1015);
and U1095 (N_1095,N_1043,N_1048);
and U1096 (N_1096,N_1037,N_1008);
nor U1097 (N_1097,N_1030,N_1019);
and U1098 (N_1098,N_1043,N_1016);
nor U1099 (N_1099,N_1023,N_1036);
nand U1100 (N_1100,N_1092,N_1098);
and U1101 (N_1101,N_1087,N_1054);
nor U1102 (N_1102,N_1082,N_1097);
or U1103 (N_1103,N_1061,N_1068);
nor U1104 (N_1104,N_1090,N_1091);
or U1105 (N_1105,N_1050,N_1069);
nor U1106 (N_1106,N_1065,N_1085);
nor U1107 (N_1107,N_1072,N_1053);
nor U1108 (N_1108,N_1058,N_1060);
or U1109 (N_1109,N_1096,N_1099);
nor U1110 (N_1110,N_1059,N_1076);
and U1111 (N_1111,N_1073,N_1062);
nand U1112 (N_1112,N_1055,N_1052);
nand U1113 (N_1113,N_1093,N_1056);
xor U1114 (N_1114,N_1079,N_1095);
nand U1115 (N_1115,N_1077,N_1063);
and U1116 (N_1116,N_1084,N_1080);
and U1117 (N_1117,N_1074,N_1081);
nor U1118 (N_1118,N_1051,N_1088);
or U1119 (N_1119,N_1071,N_1066);
nand U1120 (N_1120,N_1070,N_1094);
nand U1121 (N_1121,N_1075,N_1083);
and U1122 (N_1122,N_1086,N_1067);
nor U1123 (N_1123,N_1078,N_1089);
nand U1124 (N_1124,N_1057,N_1064);
xnor U1125 (N_1125,N_1096,N_1062);
nor U1126 (N_1126,N_1093,N_1095);
nor U1127 (N_1127,N_1050,N_1076);
nand U1128 (N_1128,N_1097,N_1063);
or U1129 (N_1129,N_1083,N_1060);
and U1130 (N_1130,N_1071,N_1061);
nor U1131 (N_1131,N_1065,N_1053);
nand U1132 (N_1132,N_1050,N_1070);
nor U1133 (N_1133,N_1069,N_1060);
and U1134 (N_1134,N_1099,N_1076);
or U1135 (N_1135,N_1074,N_1070);
or U1136 (N_1136,N_1089,N_1092);
nand U1137 (N_1137,N_1078,N_1075);
nand U1138 (N_1138,N_1053,N_1091);
nand U1139 (N_1139,N_1065,N_1079);
nor U1140 (N_1140,N_1064,N_1076);
nor U1141 (N_1141,N_1076,N_1074);
and U1142 (N_1142,N_1055,N_1062);
or U1143 (N_1143,N_1083,N_1064);
nor U1144 (N_1144,N_1063,N_1051);
and U1145 (N_1145,N_1062,N_1087);
or U1146 (N_1146,N_1069,N_1064);
and U1147 (N_1147,N_1094,N_1053);
nor U1148 (N_1148,N_1067,N_1081);
nand U1149 (N_1149,N_1077,N_1093);
nand U1150 (N_1150,N_1146,N_1103);
nand U1151 (N_1151,N_1140,N_1126);
nand U1152 (N_1152,N_1147,N_1134);
nor U1153 (N_1153,N_1106,N_1132);
or U1154 (N_1154,N_1124,N_1102);
and U1155 (N_1155,N_1111,N_1123);
and U1156 (N_1156,N_1125,N_1100);
and U1157 (N_1157,N_1105,N_1107);
nor U1158 (N_1158,N_1122,N_1104);
nor U1159 (N_1159,N_1130,N_1143);
and U1160 (N_1160,N_1117,N_1119);
nor U1161 (N_1161,N_1138,N_1101);
nor U1162 (N_1162,N_1109,N_1133);
or U1163 (N_1163,N_1137,N_1108);
and U1164 (N_1164,N_1112,N_1115);
and U1165 (N_1165,N_1144,N_1128);
nand U1166 (N_1166,N_1149,N_1141);
nor U1167 (N_1167,N_1127,N_1114);
or U1168 (N_1168,N_1110,N_1148);
nand U1169 (N_1169,N_1121,N_1120);
or U1170 (N_1170,N_1116,N_1129);
nand U1171 (N_1171,N_1142,N_1135);
nor U1172 (N_1172,N_1131,N_1113);
nand U1173 (N_1173,N_1139,N_1145);
nor U1174 (N_1174,N_1118,N_1136);
nand U1175 (N_1175,N_1102,N_1105);
xor U1176 (N_1176,N_1132,N_1131);
nand U1177 (N_1177,N_1125,N_1137);
nor U1178 (N_1178,N_1131,N_1122);
and U1179 (N_1179,N_1117,N_1104);
or U1180 (N_1180,N_1109,N_1140);
nand U1181 (N_1181,N_1105,N_1125);
nand U1182 (N_1182,N_1114,N_1136);
or U1183 (N_1183,N_1127,N_1138);
or U1184 (N_1184,N_1111,N_1130);
or U1185 (N_1185,N_1123,N_1119);
nand U1186 (N_1186,N_1143,N_1107);
and U1187 (N_1187,N_1117,N_1101);
or U1188 (N_1188,N_1119,N_1140);
xor U1189 (N_1189,N_1142,N_1113);
nor U1190 (N_1190,N_1143,N_1104);
or U1191 (N_1191,N_1108,N_1106);
nor U1192 (N_1192,N_1107,N_1111);
and U1193 (N_1193,N_1147,N_1145);
and U1194 (N_1194,N_1118,N_1131);
or U1195 (N_1195,N_1142,N_1146);
nand U1196 (N_1196,N_1147,N_1148);
nand U1197 (N_1197,N_1138,N_1133);
nor U1198 (N_1198,N_1147,N_1101);
nand U1199 (N_1199,N_1149,N_1130);
or U1200 (N_1200,N_1184,N_1192);
and U1201 (N_1201,N_1177,N_1199);
or U1202 (N_1202,N_1159,N_1162);
nand U1203 (N_1203,N_1163,N_1160);
and U1204 (N_1204,N_1191,N_1155);
or U1205 (N_1205,N_1195,N_1174);
nor U1206 (N_1206,N_1170,N_1193);
nor U1207 (N_1207,N_1166,N_1171);
nand U1208 (N_1208,N_1154,N_1179);
or U1209 (N_1209,N_1183,N_1167);
and U1210 (N_1210,N_1187,N_1165);
and U1211 (N_1211,N_1180,N_1190);
and U1212 (N_1212,N_1172,N_1157);
nand U1213 (N_1213,N_1151,N_1176);
nor U1214 (N_1214,N_1185,N_1173);
and U1215 (N_1215,N_1198,N_1158);
nor U1216 (N_1216,N_1175,N_1194);
and U1217 (N_1217,N_1181,N_1197);
nor U1218 (N_1218,N_1169,N_1186);
nor U1219 (N_1219,N_1156,N_1161);
nand U1220 (N_1220,N_1189,N_1188);
nand U1221 (N_1221,N_1153,N_1164);
and U1222 (N_1222,N_1150,N_1178);
nor U1223 (N_1223,N_1152,N_1168);
nor U1224 (N_1224,N_1182,N_1196);
and U1225 (N_1225,N_1188,N_1191);
and U1226 (N_1226,N_1166,N_1189);
or U1227 (N_1227,N_1174,N_1185);
and U1228 (N_1228,N_1179,N_1177);
nand U1229 (N_1229,N_1178,N_1177);
nand U1230 (N_1230,N_1167,N_1166);
nand U1231 (N_1231,N_1198,N_1153);
and U1232 (N_1232,N_1180,N_1155);
and U1233 (N_1233,N_1171,N_1151);
or U1234 (N_1234,N_1165,N_1151);
or U1235 (N_1235,N_1181,N_1176);
or U1236 (N_1236,N_1152,N_1181);
nand U1237 (N_1237,N_1161,N_1187);
xor U1238 (N_1238,N_1163,N_1189);
nand U1239 (N_1239,N_1190,N_1199);
or U1240 (N_1240,N_1186,N_1154);
nand U1241 (N_1241,N_1163,N_1172);
xnor U1242 (N_1242,N_1179,N_1190);
or U1243 (N_1243,N_1190,N_1172);
nor U1244 (N_1244,N_1187,N_1153);
and U1245 (N_1245,N_1154,N_1177);
nor U1246 (N_1246,N_1184,N_1188);
and U1247 (N_1247,N_1165,N_1157);
nand U1248 (N_1248,N_1160,N_1198);
nor U1249 (N_1249,N_1164,N_1169);
and U1250 (N_1250,N_1242,N_1207);
nor U1251 (N_1251,N_1247,N_1201);
nand U1252 (N_1252,N_1222,N_1245);
or U1253 (N_1253,N_1228,N_1238);
or U1254 (N_1254,N_1226,N_1235);
and U1255 (N_1255,N_1215,N_1229);
or U1256 (N_1256,N_1205,N_1206);
nor U1257 (N_1257,N_1211,N_1214);
nor U1258 (N_1258,N_1217,N_1223);
nand U1259 (N_1259,N_1237,N_1219);
or U1260 (N_1260,N_1244,N_1213);
and U1261 (N_1261,N_1227,N_1210);
or U1262 (N_1262,N_1203,N_1209);
or U1263 (N_1263,N_1246,N_1220);
or U1264 (N_1264,N_1232,N_1248);
or U1265 (N_1265,N_1202,N_1230);
and U1266 (N_1266,N_1243,N_1200);
or U1267 (N_1267,N_1204,N_1234);
and U1268 (N_1268,N_1249,N_1208);
and U1269 (N_1269,N_1221,N_1216);
nor U1270 (N_1270,N_1218,N_1212);
nand U1271 (N_1271,N_1231,N_1236);
or U1272 (N_1272,N_1224,N_1241);
nand U1273 (N_1273,N_1225,N_1233);
or U1274 (N_1274,N_1240,N_1239);
nand U1275 (N_1275,N_1223,N_1212);
and U1276 (N_1276,N_1217,N_1211);
nand U1277 (N_1277,N_1243,N_1203);
nand U1278 (N_1278,N_1230,N_1225);
nor U1279 (N_1279,N_1234,N_1219);
nor U1280 (N_1280,N_1210,N_1249);
nand U1281 (N_1281,N_1247,N_1224);
xor U1282 (N_1282,N_1244,N_1210);
nand U1283 (N_1283,N_1248,N_1242);
and U1284 (N_1284,N_1227,N_1205);
and U1285 (N_1285,N_1206,N_1234);
or U1286 (N_1286,N_1245,N_1201);
nor U1287 (N_1287,N_1217,N_1248);
nor U1288 (N_1288,N_1243,N_1221);
nor U1289 (N_1289,N_1214,N_1240);
and U1290 (N_1290,N_1218,N_1241);
and U1291 (N_1291,N_1212,N_1235);
nor U1292 (N_1292,N_1249,N_1246);
and U1293 (N_1293,N_1228,N_1243);
and U1294 (N_1294,N_1205,N_1210);
and U1295 (N_1295,N_1247,N_1236);
nor U1296 (N_1296,N_1248,N_1229);
nand U1297 (N_1297,N_1239,N_1216);
or U1298 (N_1298,N_1200,N_1207);
nand U1299 (N_1299,N_1241,N_1213);
nand U1300 (N_1300,N_1285,N_1287);
nand U1301 (N_1301,N_1273,N_1267);
or U1302 (N_1302,N_1264,N_1277);
nor U1303 (N_1303,N_1278,N_1282);
nor U1304 (N_1304,N_1288,N_1258);
and U1305 (N_1305,N_1291,N_1261);
or U1306 (N_1306,N_1284,N_1251);
and U1307 (N_1307,N_1252,N_1280);
nor U1308 (N_1308,N_1254,N_1257);
or U1309 (N_1309,N_1256,N_1299);
nand U1310 (N_1310,N_1297,N_1296);
or U1311 (N_1311,N_1265,N_1292);
nor U1312 (N_1312,N_1298,N_1281);
and U1313 (N_1313,N_1289,N_1271);
nor U1314 (N_1314,N_1262,N_1260);
nand U1315 (N_1315,N_1253,N_1294);
and U1316 (N_1316,N_1286,N_1263);
or U1317 (N_1317,N_1290,N_1255);
nand U1318 (N_1318,N_1272,N_1268);
nand U1319 (N_1319,N_1266,N_1270);
nand U1320 (N_1320,N_1259,N_1295);
and U1321 (N_1321,N_1293,N_1283);
nand U1322 (N_1322,N_1269,N_1274);
or U1323 (N_1323,N_1276,N_1279);
and U1324 (N_1324,N_1275,N_1250);
nor U1325 (N_1325,N_1272,N_1253);
and U1326 (N_1326,N_1261,N_1259);
nor U1327 (N_1327,N_1268,N_1289);
nor U1328 (N_1328,N_1254,N_1272);
nand U1329 (N_1329,N_1278,N_1262);
nand U1330 (N_1330,N_1283,N_1265);
nand U1331 (N_1331,N_1274,N_1289);
and U1332 (N_1332,N_1282,N_1286);
and U1333 (N_1333,N_1280,N_1266);
nor U1334 (N_1334,N_1255,N_1280);
nor U1335 (N_1335,N_1252,N_1295);
and U1336 (N_1336,N_1275,N_1291);
or U1337 (N_1337,N_1257,N_1253);
and U1338 (N_1338,N_1281,N_1253);
and U1339 (N_1339,N_1250,N_1286);
or U1340 (N_1340,N_1256,N_1287);
nand U1341 (N_1341,N_1298,N_1283);
nor U1342 (N_1342,N_1254,N_1268);
or U1343 (N_1343,N_1273,N_1292);
or U1344 (N_1344,N_1282,N_1273);
xnor U1345 (N_1345,N_1288,N_1298);
and U1346 (N_1346,N_1274,N_1298);
xor U1347 (N_1347,N_1267,N_1293);
nand U1348 (N_1348,N_1253,N_1258);
xnor U1349 (N_1349,N_1276,N_1284);
nand U1350 (N_1350,N_1340,N_1345);
and U1351 (N_1351,N_1335,N_1326);
nor U1352 (N_1352,N_1343,N_1301);
or U1353 (N_1353,N_1321,N_1346);
and U1354 (N_1354,N_1309,N_1304);
nand U1355 (N_1355,N_1312,N_1323);
nand U1356 (N_1356,N_1331,N_1322);
nand U1357 (N_1357,N_1316,N_1300);
nor U1358 (N_1358,N_1314,N_1307);
and U1359 (N_1359,N_1319,N_1349);
and U1360 (N_1360,N_1320,N_1339);
nor U1361 (N_1361,N_1329,N_1303);
nor U1362 (N_1362,N_1348,N_1341);
or U1363 (N_1363,N_1336,N_1306);
nor U1364 (N_1364,N_1317,N_1330);
or U1365 (N_1365,N_1313,N_1332);
and U1366 (N_1366,N_1342,N_1328);
nor U1367 (N_1367,N_1344,N_1308);
nor U1368 (N_1368,N_1337,N_1318);
nor U1369 (N_1369,N_1324,N_1333);
or U1370 (N_1370,N_1305,N_1327);
and U1371 (N_1371,N_1334,N_1315);
or U1372 (N_1372,N_1311,N_1338);
and U1373 (N_1373,N_1302,N_1347);
and U1374 (N_1374,N_1310,N_1325);
nor U1375 (N_1375,N_1343,N_1318);
and U1376 (N_1376,N_1332,N_1335);
or U1377 (N_1377,N_1316,N_1331);
nor U1378 (N_1378,N_1306,N_1342);
or U1379 (N_1379,N_1331,N_1317);
nand U1380 (N_1380,N_1335,N_1324);
nor U1381 (N_1381,N_1334,N_1303);
nand U1382 (N_1382,N_1325,N_1327);
or U1383 (N_1383,N_1305,N_1337);
and U1384 (N_1384,N_1335,N_1323);
nand U1385 (N_1385,N_1308,N_1336);
and U1386 (N_1386,N_1317,N_1301);
or U1387 (N_1387,N_1306,N_1330);
xor U1388 (N_1388,N_1329,N_1311);
or U1389 (N_1389,N_1340,N_1330);
nand U1390 (N_1390,N_1306,N_1327);
or U1391 (N_1391,N_1324,N_1309);
or U1392 (N_1392,N_1318,N_1338);
and U1393 (N_1393,N_1336,N_1302);
nand U1394 (N_1394,N_1343,N_1320);
nor U1395 (N_1395,N_1312,N_1342);
nand U1396 (N_1396,N_1325,N_1306);
nor U1397 (N_1397,N_1312,N_1314);
or U1398 (N_1398,N_1322,N_1302);
nor U1399 (N_1399,N_1326,N_1339);
nor U1400 (N_1400,N_1390,N_1366);
or U1401 (N_1401,N_1371,N_1394);
and U1402 (N_1402,N_1397,N_1370);
nor U1403 (N_1403,N_1398,N_1358);
or U1404 (N_1404,N_1374,N_1373);
nor U1405 (N_1405,N_1379,N_1386);
nand U1406 (N_1406,N_1372,N_1375);
nand U1407 (N_1407,N_1387,N_1380);
and U1408 (N_1408,N_1359,N_1383);
and U1409 (N_1409,N_1377,N_1354);
nand U1410 (N_1410,N_1388,N_1384);
nand U1411 (N_1411,N_1355,N_1352);
nor U1412 (N_1412,N_1376,N_1356);
or U1413 (N_1413,N_1382,N_1360);
nand U1414 (N_1414,N_1396,N_1362);
or U1415 (N_1415,N_1395,N_1367);
or U1416 (N_1416,N_1391,N_1353);
or U1417 (N_1417,N_1361,N_1351);
and U1418 (N_1418,N_1364,N_1369);
and U1419 (N_1419,N_1393,N_1381);
or U1420 (N_1420,N_1392,N_1368);
nand U1421 (N_1421,N_1357,N_1378);
and U1422 (N_1422,N_1350,N_1365);
nor U1423 (N_1423,N_1363,N_1399);
or U1424 (N_1424,N_1389,N_1385);
nand U1425 (N_1425,N_1363,N_1360);
and U1426 (N_1426,N_1358,N_1364);
nand U1427 (N_1427,N_1380,N_1396);
or U1428 (N_1428,N_1389,N_1383);
nand U1429 (N_1429,N_1380,N_1358);
nor U1430 (N_1430,N_1375,N_1355);
and U1431 (N_1431,N_1395,N_1376);
nor U1432 (N_1432,N_1367,N_1355);
or U1433 (N_1433,N_1398,N_1392);
xnor U1434 (N_1434,N_1361,N_1369);
nor U1435 (N_1435,N_1392,N_1372);
or U1436 (N_1436,N_1390,N_1370);
and U1437 (N_1437,N_1379,N_1360);
or U1438 (N_1438,N_1390,N_1399);
and U1439 (N_1439,N_1383,N_1382);
nand U1440 (N_1440,N_1360,N_1367);
and U1441 (N_1441,N_1380,N_1385);
and U1442 (N_1442,N_1392,N_1374);
or U1443 (N_1443,N_1374,N_1370);
nor U1444 (N_1444,N_1393,N_1377);
nor U1445 (N_1445,N_1373,N_1394);
and U1446 (N_1446,N_1351,N_1373);
nand U1447 (N_1447,N_1376,N_1394);
xnor U1448 (N_1448,N_1376,N_1390);
or U1449 (N_1449,N_1396,N_1391);
and U1450 (N_1450,N_1404,N_1415);
nand U1451 (N_1451,N_1444,N_1418);
or U1452 (N_1452,N_1416,N_1447);
and U1453 (N_1453,N_1420,N_1449);
nor U1454 (N_1454,N_1403,N_1445);
and U1455 (N_1455,N_1441,N_1402);
nor U1456 (N_1456,N_1412,N_1448);
or U1457 (N_1457,N_1426,N_1414);
nor U1458 (N_1458,N_1425,N_1400);
or U1459 (N_1459,N_1423,N_1428);
nor U1460 (N_1460,N_1439,N_1408);
or U1461 (N_1461,N_1422,N_1411);
nand U1462 (N_1462,N_1407,N_1438);
nand U1463 (N_1463,N_1436,N_1429);
nand U1464 (N_1464,N_1405,N_1409);
xor U1465 (N_1465,N_1442,N_1421);
or U1466 (N_1466,N_1430,N_1406);
nand U1467 (N_1467,N_1434,N_1437);
nor U1468 (N_1468,N_1424,N_1413);
nand U1469 (N_1469,N_1410,N_1427);
nor U1470 (N_1470,N_1433,N_1419);
or U1471 (N_1471,N_1446,N_1440);
nand U1472 (N_1472,N_1417,N_1401);
or U1473 (N_1473,N_1431,N_1432);
or U1474 (N_1474,N_1435,N_1443);
and U1475 (N_1475,N_1403,N_1426);
nand U1476 (N_1476,N_1409,N_1441);
nor U1477 (N_1477,N_1402,N_1443);
xor U1478 (N_1478,N_1434,N_1438);
nand U1479 (N_1479,N_1447,N_1408);
and U1480 (N_1480,N_1410,N_1430);
and U1481 (N_1481,N_1448,N_1443);
nand U1482 (N_1482,N_1444,N_1420);
and U1483 (N_1483,N_1416,N_1444);
nand U1484 (N_1484,N_1410,N_1437);
nand U1485 (N_1485,N_1400,N_1420);
nor U1486 (N_1486,N_1431,N_1437);
nor U1487 (N_1487,N_1441,N_1446);
or U1488 (N_1488,N_1413,N_1435);
nor U1489 (N_1489,N_1432,N_1436);
and U1490 (N_1490,N_1449,N_1438);
nand U1491 (N_1491,N_1409,N_1431);
or U1492 (N_1492,N_1445,N_1430);
and U1493 (N_1493,N_1433,N_1441);
and U1494 (N_1494,N_1433,N_1421);
nand U1495 (N_1495,N_1402,N_1442);
and U1496 (N_1496,N_1408,N_1449);
or U1497 (N_1497,N_1402,N_1406);
nor U1498 (N_1498,N_1421,N_1406);
and U1499 (N_1499,N_1405,N_1415);
nand U1500 (N_1500,N_1479,N_1471);
nor U1501 (N_1501,N_1469,N_1473);
nand U1502 (N_1502,N_1456,N_1470);
nand U1503 (N_1503,N_1451,N_1477);
and U1504 (N_1504,N_1468,N_1490);
and U1505 (N_1505,N_1478,N_1465);
nand U1506 (N_1506,N_1453,N_1499);
nor U1507 (N_1507,N_1450,N_1480);
or U1508 (N_1508,N_1498,N_1475);
and U1509 (N_1509,N_1457,N_1485);
nor U1510 (N_1510,N_1483,N_1464);
nand U1511 (N_1511,N_1496,N_1493);
nand U1512 (N_1512,N_1472,N_1458);
nor U1513 (N_1513,N_1497,N_1455);
and U1514 (N_1514,N_1494,N_1491);
and U1515 (N_1515,N_1463,N_1481);
or U1516 (N_1516,N_1495,N_1462);
xor U1517 (N_1517,N_1489,N_1476);
and U1518 (N_1518,N_1474,N_1460);
nor U1519 (N_1519,N_1488,N_1461);
or U1520 (N_1520,N_1487,N_1482);
nor U1521 (N_1521,N_1467,N_1459);
and U1522 (N_1522,N_1484,N_1454);
and U1523 (N_1523,N_1486,N_1452);
nor U1524 (N_1524,N_1466,N_1492);
nor U1525 (N_1525,N_1472,N_1455);
nor U1526 (N_1526,N_1494,N_1479);
nor U1527 (N_1527,N_1463,N_1455);
nor U1528 (N_1528,N_1491,N_1477);
or U1529 (N_1529,N_1482,N_1453);
and U1530 (N_1530,N_1454,N_1490);
and U1531 (N_1531,N_1460,N_1473);
and U1532 (N_1532,N_1485,N_1482);
nor U1533 (N_1533,N_1457,N_1458);
or U1534 (N_1534,N_1473,N_1488);
nand U1535 (N_1535,N_1480,N_1456);
or U1536 (N_1536,N_1458,N_1466);
and U1537 (N_1537,N_1452,N_1481);
nor U1538 (N_1538,N_1460,N_1492);
and U1539 (N_1539,N_1451,N_1484);
nor U1540 (N_1540,N_1465,N_1493);
or U1541 (N_1541,N_1453,N_1496);
nand U1542 (N_1542,N_1477,N_1450);
or U1543 (N_1543,N_1486,N_1461);
nand U1544 (N_1544,N_1482,N_1467);
or U1545 (N_1545,N_1451,N_1471);
nand U1546 (N_1546,N_1473,N_1478);
nand U1547 (N_1547,N_1450,N_1464);
nand U1548 (N_1548,N_1493,N_1490);
or U1549 (N_1549,N_1477,N_1473);
or U1550 (N_1550,N_1512,N_1515);
nand U1551 (N_1551,N_1516,N_1519);
or U1552 (N_1552,N_1526,N_1543);
nand U1553 (N_1553,N_1508,N_1520);
and U1554 (N_1554,N_1538,N_1523);
and U1555 (N_1555,N_1522,N_1547);
nor U1556 (N_1556,N_1502,N_1506);
or U1557 (N_1557,N_1527,N_1537);
nand U1558 (N_1558,N_1528,N_1535);
nor U1559 (N_1559,N_1511,N_1533);
or U1560 (N_1560,N_1534,N_1513);
or U1561 (N_1561,N_1549,N_1545);
or U1562 (N_1562,N_1509,N_1524);
nor U1563 (N_1563,N_1514,N_1544);
and U1564 (N_1564,N_1548,N_1531);
or U1565 (N_1565,N_1539,N_1536);
and U1566 (N_1566,N_1521,N_1525);
nand U1567 (N_1567,N_1542,N_1501);
nor U1568 (N_1568,N_1517,N_1546);
and U1569 (N_1569,N_1530,N_1529);
or U1570 (N_1570,N_1507,N_1503);
or U1571 (N_1571,N_1500,N_1505);
nor U1572 (N_1572,N_1518,N_1532);
and U1573 (N_1573,N_1504,N_1540);
and U1574 (N_1574,N_1510,N_1541);
nand U1575 (N_1575,N_1534,N_1501);
or U1576 (N_1576,N_1526,N_1544);
nor U1577 (N_1577,N_1542,N_1523);
and U1578 (N_1578,N_1514,N_1524);
nor U1579 (N_1579,N_1521,N_1542);
and U1580 (N_1580,N_1507,N_1533);
nor U1581 (N_1581,N_1523,N_1532);
or U1582 (N_1582,N_1502,N_1521);
and U1583 (N_1583,N_1509,N_1530);
or U1584 (N_1584,N_1519,N_1521);
nor U1585 (N_1585,N_1544,N_1538);
or U1586 (N_1586,N_1526,N_1538);
nor U1587 (N_1587,N_1519,N_1520);
or U1588 (N_1588,N_1548,N_1538);
or U1589 (N_1589,N_1545,N_1544);
nand U1590 (N_1590,N_1518,N_1513);
or U1591 (N_1591,N_1516,N_1534);
or U1592 (N_1592,N_1506,N_1513);
and U1593 (N_1593,N_1510,N_1529);
or U1594 (N_1594,N_1548,N_1530);
and U1595 (N_1595,N_1514,N_1500);
nand U1596 (N_1596,N_1519,N_1510);
nand U1597 (N_1597,N_1532,N_1540);
nor U1598 (N_1598,N_1543,N_1509);
nand U1599 (N_1599,N_1507,N_1529);
nor U1600 (N_1600,N_1570,N_1569);
nand U1601 (N_1601,N_1589,N_1566);
and U1602 (N_1602,N_1578,N_1573);
nor U1603 (N_1603,N_1581,N_1585);
nand U1604 (N_1604,N_1593,N_1565);
and U1605 (N_1605,N_1560,N_1556);
and U1606 (N_1606,N_1572,N_1597);
or U1607 (N_1607,N_1592,N_1580);
or U1608 (N_1608,N_1575,N_1553);
and U1609 (N_1609,N_1563,N_1587);
nor U1610 (N_1610,N_1584,N_1586);
nor U1611 (N_1611,N_1562,N_1576);
and U1612 (N_1612,N_1583,N_1571);
nand U1613 (N_1613,N_1574,N_1555);
or U1614 (N_1614,N_1550,N_1588);
nand U1615 (N_1615,N_1579,N_1552);
nand U1616 (N_1616,N_1567,N_1599);
and U1617 (N_1617,N_1591,N_1551);
and U1618 (N_1618,N_1554,N_1561);
or U1619 (N_1619,N_1557,N_1590);
nand U1620 (N_1620,N_1598,N_1577);
nand U1621 (N_1621,N_1558,N_1594);
and U1622 (N_1622,N_1564,N_1595);
and U1623 (N_1623,N_1582,N_1559);
and U1624 (N_1624,N_1568,N_1596);
or U1625 (N_1625,N_1587,N_1574);
and U1626 (N_1626,N_1559,N_1558);
and U1627 (N_1627,N_1573,N_1582);
nand U1628 (N_1628,N_1559,N_1593);
or U1629 (N_1629,N_1574,N_1582);
or U1630 (N_1630,N_1552,N_1585);
nor U1631 (N_1631,N_1551,N_1566);
or U1632 (N_1632,N_1581,N_1568);
or U1633 (N_1633,N_1563,N_1569);
and U1634 (N_1634,N_1580,N_1594);
nand U1635 (N_1635,N_1592,N_1563);
nor U1636 (N_1636,N_1581,N_1574);
nand U1637 (N_1637,N_1560,N_1574);
or U1638 (N_1638,N_1586,N_1551);
and U1639 (N_1639,N_1556,N_1558);
and U1640 (N_1640,N_1576,N_1568);
and U1641 (N_1641,N_1564,N_1573);
nor U1642 (N_1642,N_1574,N_1567);
xor U1643 (N_1643,N_1551,N_1572);
or U1644 (N_1644,N_1585,N_1562);
nor U1645 (N_1645,N_1572,N_1599);
and U1646 (N_1646,N_1563,N_1552);
nand U1647 (N_1647,N_1591,N_1563);
nand U1648 (N_1648,N_1593,N_1590);
nand U1649 (N_1649,N_1569,N_1584);
nor U1650 (N_1650,N_1607,N_1618);
or U1651 (N_1651,N_1616,N_1614);
and U1652 (N_1652,N_1619,N_1640);
xor U1653 (N_1653,N_1648,N_1632);
nand U1654 (N_1654,N_1615,N_1626);
nor U1655 (N_1655,N_1630,N_1647);
and U1656 (N_1656,N_1608,N_1603);
nor U1657 (N_1657,N_1645,N_1629);
or U1658 (N_1658,N_1605,N_1633);
xnor U1659 (N_1659,N_1601,N_1644);
nor U1660 (N_1660,N_1636,N_1631);
xor U1661 (N_1661,N_1627,N_1637);
nor U1662 (N_1662,N_1641,N_1634);
or U1663 (N_1663,N_1610,N_1611);
and U1664 (N_1664,N_1606,N_1639);
and U1665 (N_1665,N_1617,N_1621);
or U1666 (N_1666,N_1643,N_1628);
or U1667 (N_1667,N_1646,N_1604);
nand U1668 (N_1668,N_1649,N_1613);
nor U1669 (N_1669,N_1624,N_1642);
and U1670 (N_1670,N_1635,N_1623);
nand U1671 (N_1671,N_1600,N_1625);
nor U1672 (N_1672,N_1622,N_1602);
nand U1673 (N_1673,N_1609,N_1638);
nand U1674 (N_1674,N_1612,N_1620);
xnor U1675 (N_1675,N_1615,N_1611);
nor U1676 (N_1676,N_1614,N_1628);
and U1677 (N_1677,N_1604,N_1616);
or U1678 (N_1678,N_1627,N_1623);
or U1679 (N_1679,N_1609,N_1628);
and U1680 (N_1680,N_1624,N_1605);
or U1681 (N_1681,N_1615,N_1623);
nor U1682 (N_1682,N_1605,N_1608);
or U1683 (N_1683,N_1617,N_1614);
nand U1684 (N_1684,N_1604,N_1627);
nand U1685 (N_1685,N_1636,N_1640);
nand U1686 (N_1686,N_1641,N_1621);
or U1687 (N_1687,N_1646,N_1608);
or U1688 (N_1688,N_1646,N_1641);
and U1689 (N_1689,N_1621,N_1613);
and U1690 (N_1690,N_1642,N_1603);
nor U1691 (N_1691,N_1603,N_1617);
and U1692 (N_1692,N_1616,N_1646);
or U1693 (N_1693,N_1614,N_1641);
xor U1694 (N_1694,N_1641,N_1636);
nand U1695 (N_1695,N_1643,N_1648);
or U1696 (N_1696,N_1644,N_1600);
and U1697 (N_1697,N_1630,N_1629);
nor U1698 (N_1698,N_1640,N_1641);
xnor U1699 (N_1699,N_1630,N_1636);
or U1700 (N_1700,N_1698,N_1677);
nor U1701 (N_1701,N_1669,N_1654);
nor U1702 (N_1702,N_1663,N_1681);
xnor U1703 (N_1703,N_1655,N_1668);
and U1704 (N_1704,N_1678,N_1657);
nor U1705 (N_1705,N_1683,N_1665);
and U1706 (N_1706,N_1691,N_1673);
nor U1707 (N_1707,N_1684,N_1692);
nor U1708 (N_1708,N_1660,N_1690);
and U1709 (N_1709,N_1661,N_1662);
or U1710 (N_1710,N_1667,N_1679);
nor U1711 (N_1711,N_1672,N_1676);
nor U1712 (N_1712,N_1687,N_1680);
and U1713 (N_1713,N_1675,N_1696);
and U1714 (N_1714,N_1650,N_1671);
or U1715 (N_1715,N_1659,N_1666);
or U1716 (N_1716,N_1685,N_1653);
or U1717 (N_1717,N_1674,N_1682);
nor U1718 (N_1718,N_1670,N_1664);
or U1719 (N_1719,N_1693,N_1658);
or U1720 (N_1720,N_1697,N_1686);
nand U1721 (N_1721,N_1694,N_1656);
or U1722 (N_1722,N_1688,N_1699);
nand U1723 (N_1723,N_1652,N_1695);
or U1724 (N_1724,N_1689,N_1651);
or U1725 (N_1725,N_1695,N_1688);
nand U1726 (N_1726,N_1693,N_1684);
nand U1727 (N_1727,N_1672,N_1688);
nor U1728 (N_1728,N_1658,N_1678);
nand U1729 (N_1729,N_1687,N_1664);
or U1730 (N_1730,N_1650,N_1694);
or U1731 (N_1731,N_1651,N_1686);
or U1732 (N_1732,N_1691,N_1685);
and U1733 (N_1733,N_1679,N_1657);
nand U1734 (N_1734,N_1688,N_1656);
or U1735 (N_1735,N_1659,N_1679);
nand U1736 (N_1736,N_1692,N_1694);
nor U1737 (N_1737,N_1679,N_1693);
and U1738 (N_1738,N_1667,N_1675);
and U1739 (N_1739,N_1673,N_1657);
and U1740 (N_1740,N_1691,N_1696);
or U1741 (N_1741,N_1680,N_1655);
nor U1742 (N_1742,N_1696,N_1656);
or U1743 (N_1743,N_1654,N_1661);
and U1744 (N_1744,N_1656,N_1689);
nor U1745 (N_1745,N_1668,N_1691);
nand U1746 (N_1746,N_1650,N_1666);
or U1747 (N_1747,N_1656,N_1687);
nand U1748 (N_1748,N_1695,N_1677);
and U1749 (N_1749,N_1655,N_1682);
and U1750 (N_1750,N_1725,N_1708);
nor U1751 (N_1751,N_1706,N_1730);
and U1752 (N_1752,N_1736,N_1700);
and U1753 (N_1753,N_1735,N_1705);
or U1754 (N_1754,N_1743,N_1746);
nor U1755 (N_1755,N_1718,N_1702);
or U1756 (N_1756,N_1748,N_1749);
and U1757 (N_1757,N_1747,N_1716);
and U1758 (N_1758,N_1737,N_1724);
and U1759 (N_1759,N_1717,N_1728);
and U1760 (N_1760,N_1710,N_1739);
nand U1761 (N_1761,N_1721,N_1704);
nor U1762 (N_1762,N_1742,N_1740);
nor U1763 (N_1763,N_1745,N_1719);
nand U1764 (N_1764,N_1738,N_1707);
or U1765 (N_1765,N_1732,N_1731);
nand U1766 (N_1766,N_1727,N_1726);
nor U1767 (N_1767,N_1715,N_1744);
or U1768 (N_1768,N_1701,N_1709);
and U1769 (N_1769,N_1720,N_1711);
nor U1770 (N_1770,N_1713,N_1741);
and U1771 (N_1771,N_1734,N_1714);
or U1772 (N_1772,N_1729,N_1703);
xnor U1773 (N_1773,N_1723,N_1722);
and U1774 (N_1774,N_1733,N_1712);
nand U1775 (N_1775,N_1706,N_1719);
or U1776 (N_1776,N_1716,N_1743);
or U1777 (N_1777,N_1723,N_1746);
nor U1778 (N_1778,N_1727,N_1701);
nor U1779 (N_1779,N_1705,N_1703);
nor U1780 (N_1780,N_1739,N_1747);
and U1781 (N_1781,N_1735,N_1744);
nor U1782 (N_1782,N_1700,N_1710);
nand U1783 (N_1783,N_1726,N_1710);
nand U1784 (N_1784,N_1703,N_1735);
nand U1785 (N_1785,N_1721,N_1703);
nor U1786 (N_1786,N_1747,N_1746);
nand U1787 (N_1787,N_1732,N_1741);
nand U1788 (N_1788,N_1729,N_1715);
nand U1789 (N_1789,N_1726,N_1717);
nand U1790 (N_1790,N_1742,N_1747);
and U1791 (N_1791,N_1729,N_1739);
and U1792 (N_1792,N_1742,N_1717);
nand U1793 (N_1793,N_1710,N_1721);
or U1794 (N_1794,N_1721,N_1722);
nor U1795 (N_1795,N_1738,N_1702);
and U1796 (N_1796,N_1737,N_1733);
nand U1797 (N_1797,N_1713,N_1715);
xnor U1798 (N_1798,N_1745,N_1737);
nor U1799 (N_1799,N_1711,N_1717);
and U1800 (N_1800,N_1765,N_1795);
nand U1801 (N_1801,N_1754,N_1793);
nand U1802 (N_1802,N_1757,N_1779);
or U1803 (N_1803,N_1767,N_1755);
nor U1804 (N_1804,N_1776,N_1756);
nor U1805 (N_1805,N_1782,N_1787);
nor U1806 (N_1806,N_1771,N_1763);
or U1807 (N_1807,N_1766,N_1794);
xor U1808 (N_1808,N_1773,N_1768);
or U1809 (N_1809,N_1798,N_1750);
xnor U1810 (N_1810,N_1788,N_1772);
or U1811 (N_1811,N_1774,N_1760);
nand U1812 (N_1812,N_1777,N_1770);
and U1813 (N_1813,N_1790,N_1791);
nor U1814 (N_1814,N_1786,N_1751);
nand U1815 (N_1815,N_1762,N_1775);
or U1816 (N_1816,N_1764,N_1785);
or U1817 (N_1817,N_1781,N_1761);
and U1818 (N_1818,N_1789,N_1759);
or U1819 (N_1819,N_1784,N_1758);
nor U1820 (N_1820,N_1753,N_1752);
nand U1821 (N_1821,N_1783,N_1769);
or U1822 (N_1822,N_1780,N_1799);
and U1823 (N_1823,N_1778,N_1796);
nand U1824 (N_1824,N_1792,N_1797);
or U1825 (N_1825,N_1798,N_1758);
or U1826 (N_1826,N_1772,N_1773);
xnor U1827 (N_1827,N_1791,N_1781);
nor U1828 (N_1828,N_1757,N_1771);
and U1829 (N_1829,N_1792,N_1780);
and U1830 (N_1830,N_1776,N_1785);
and U1831 (N_1831,N_1796,N_1798);
and U1832 (N_1832,N_1759,N_1795);
nand U1833 (N_1833,N_1771,N_1761);
nand U1834 (N_1834,N_1779,N_1769);
and U1835 (N_1835,N_1786,N_1776);
nand U1836 (N_1836,N_1771,N_1792);
nor U1837 (N_1837,N_1763,N_1772);
and U1838 (N_1838,N_1757,N_1794);
nor U1839 (N_1839,N_1764,N_1780);
nand U1840 (N_1840,N_1759,N_1776);
or U1841 (N_1841,N_1795,N_1776);
nor U1842 (N_1842,N_1782,N_1781);
nor U1843 (N_1843,N_1798,N_1755);
and U1844 (N_1844,N_1794,N_1773);
and U1845 (N_1845,N_1792,N_1782);
nand U1846 (N_1846,N_1766,N_1774);
and U1847 (N_1847,N_1779,N_1776);
and U1848 (N_1848,N_1786,N_1764);
nand U1849 (N_1849,N_1755,N_1775);
and U1850 (N_1850,N_1811,N_1832);
nor U1851 (N_1851,N_1809,N_1840);
nand U1852 (N_1852,N_1838,N_1836);
nand U1853 (N_1853,N_1819,N_1806);
nor U1854 (N_1854,N_1843,N_1822);
and U1855 (N_1855,N_1803,N_1825);
nand U1856 (N_1856,N_1842,N_1828);
nand U1857 (N_1857,N_1826,N_1810);
and U1858 (N_1858,N_1800,N_1831);
nor U1859 (N_1859,N_1827,N_1833);
nand U1860 (N_1860,N_1815,N_1844);
nand U1861 (N_1861,N_1839,N_1820);
nand U1862 (N_1862,N_1834,N_1813);
or U1863 (N_1863,N_1823,N_1812);
nor U1864 (N_1864,N_1848,N_1847);
nor U1865 (N_1865,N_1802,N_1837);
and U1866 (N_1866,N_1849,N_1807);
or U1867 (N_1867,N_1821,N_1801);
or U1868 (N_1868,N_1816,N_1805);
or U1869 (N_1869,N_1817,N_1835);
nand U1870 (N_1870,N_1804,N_1814);
nor U1871 (N_1871,N_1845,N_1830);
nand U1872 (N_1872,N_1829,N_1818);
or U1873 (N_1873,N_1846,N_1808);
or U1874 (N_1874,N_1824,N_1841);
nor U1875 (N_1875,N_1842,N_1823);
or U1876 (N_1876,N_1839,N_1841);
or U1877 (N_1877,N_1804,N_1827);
nand U1878 (N_1878,N_1838,N_1824);
and U1879 (N_1879,N_1827,N_1847);
nand U1880 (N_1880,N_1811,N_1831);
and U1881 (N_1881,N_1818,N_1838);
nand U1882 (N_1882,N_1839,N_1814);
nand U1883 (N_1883,N_1823,N_1824);
nor U1884 (N_1884,N_1817,N_1826);
and U1885 (N_1885,N_1823,N_1827);
and U1886 (N_1886,N_1841,N_1821);
nand U1887 (N_1887,N_1800,N_1844);
nand U1888 (N_1888,N_1802,N_1818);
or U1889 (N_1889,N_1835,N_1807);
nand U1890 (N_1890,N_1822,N_1821);
and U1891 (N_1891,N_1823,N_1802);
and U1892 (N_1892,N_1814,N_1829);
or U1893 (N_1893,N_1818,N_1809);
nor U1894 (N_1894,N_1835,N_1831);
and U1895 (N_1895,N_1809,N_1811);
or U1896 (N_1896,N_1810,N_1800);
or U1897 (N_1897,N_1833,N_1844);
or U1898 (N_1898,N_1834,N_1848);
nand U1899 (N_1899,N_1819,N_1805);
or U1900 (N_1900,N_1887,N_1884);
nor U1901 (N_1901,N_1852,N_1862);
or U1902 (N_1902,N_1898,N_1869);
or U1903 (N_1903,N_1880,N_1867);
and U1904 (N_1904,N_1873,N_1878);
nor U1905 (N_1905,N_1856,N_1854);
nand U1906 (N_1906,N_1872,N_1851);
nand U1907 (N_1907,N_1883,N_1850);
nand U1908 (N_1908,N_1858,N_1882);
xor U1909 (N_1909,N_1875,N_1855);
or U1910 (N_1910,N_1865,N_1859);
nor U1911 (N_1911,N_1897,N_1861);
nand U1912 (N_1912,N_1896,N_1881);
or U1913 (N_1913,N_1870,N_1899);
nand U1914 (N_1914,N_1864,N_1894);
and U1915 (N_1915,N_1890,N_1879);
and U1916 (N_1916,N_1876,N_1868);
or U1917 (N_1917,N_1891,N_1866);
nor U1918 (N_1918,N_1853,N_1889);
or U1919 (N_1919,N_1863,N_1857);
and U1920 (N_1920,N_1871,N_1893);
or U1921 (N_1921,N_1895,N_1885);
or U1922 (N_1922,N_1874,N_1886);
xor U1923 (N_1923,N_1877,N_1892);
nand U1924 (N_1924,N_1860,N_1888);
nor U1925 (N_1925,N_1889,N_1872);
and U1926 (N_1926,N_1868,N_1859);
nand U1927 (N_1927,N_1860,N_1889);
and U1928 (N_1928,N_1886,N_1854);
nand U1929 (N_1929,N_1898,N_1871);
or U1930 (N_1930,N_1887,N_1894);
or U1931 (N_1931,N_1850,N_1862);
nor U1932 (N_1932,N_1898,N_1864);
nor U1933 (N_1933,N_1873,N_1893);
nor U1934 (N_1934,N_1861,N_1872);
nand U1935 (N_1935,N_1888,N_1871);
nand U1936 (N_1936,N_1874,N_1859);
nor U1937 (N_1937,N_1877,N_1899);
and U1938 (N_1938,N_1857,N_1858);
and U1939 (N_1939,N_1880,N_1888);
and U1940 (N_1940,N_1887,N_1897);
nand U1941 (N_1941,N_1899,N_1882);
nor U1942 (N_1942,N_1898,N_1853);
nand U1943 (N_1943,N_1854,N_1859);
or U1944 (N_1944,N_1889,N_1858);
or U1945 (N_1945,N_1882,N_1863);
and U1946 (N_1946,N_1868,N_1858);
and U1947 (N_1947,N_1851,N_1891);
nor U1948 (N_1948,N_1891,N_1887);
nand U1949 (N_1949,N_1886,N_1864);
and U1950 (N_1950,N_1929,N_1925);
and U1951 (N_1951,N_1918,N_1934);
or U1952 (N_1952,N_1900,N_1937);
nand U1953 (N_1953,N_1931,N_1924);
and U1954 (N_1954,N_1943,N_1917);
and U1955 (N_1955,N_1945,N_1906);
and U1956 (N_1956,N_1904,N_1944);
nor U1957 (N_1957,N_1923,N_1949);
nand U1958 (N_1958,N_1947,N_1941);
or U1959 (N_1959,N_1920,N_1905);
and U1960 (N_1960,N_1930,N_1908);
nor U1961 (N_1961,N_1933,N_1919);
and U1962 (N_1962,N_1948,N_1910);
nand U1963 (N_1963,N_1938,N_1909);
and U1964 (N_1964,N_1907,N_1932);
nor U1965 (N_1965,N_1916,N_1926);
or U1966 (N_1966,N_1902,N_1939);
nand U1967 (N_1967,N_1901,N_1946);
nor U1968 (N_1968,N_1912,N_1942);
or U1969 (N_1969,N_1911,N_1940);
and U1970 (N_1970,N_1915,N_1928);
nand U1971 (N_1971,N_1913,N_1914);
or U1972 (N_1972,N_1935,N_1903);
or U1973 (N_1973,N_1921,N_1922);
and U1974 (N_1974,N_1936,N_1927);
or U1975 (N_1975,N_1913,N_1920);
nand U1976 (N_1976,N_1941,N_1908);
or U1977 (N_1977,N_1907,N_1943);
nand U1978 (N_1978,N_1909,N_1907);
nand U1979 (N_1979,N_1906,N_1931);
nor U1980 (N_1980,N_1930,N_1927);
and U1981 (N_1981,N_1911,N_1910);
and U1982 (N_1982,N_1911,N_1902);
and U1983 (N_1983,N_1939,N_1915);
or U1984 (N_1984,N_1921,N_1942);
nand U1985 (N_1985,N_1918,N_1928);
nand U1986 (N_1986,N_1922,N_1937);
or U1987 (N_1987,N_1935,N_1924);
nor U1988 (N_1988,N_1948,N_1940);
and U1989 (N_1989,N_1922,N_1947);
or U1990 (N_1990,N_1910,N_1925);
xor U1991 (N_1991,N_1940,N_1932);
nor U1992 (N_1992,N_1942,N_1946);
nand U1993 (N_1993,N_1928,N_1924);
nor U1994 (N_1994,N_1932,N_1902);
nand U1995 (N_1995,N_1935,N_1910);
and U1996 (N_1996,N_1940,N_1943);
nor U1997 (N_1997,N_1918,N_1914);
or U1998 (N_1998,N_1919,N_1932);
nand U1999 (N_1999,N_1932,N_1948);
nor U2000 (N_2000,N_1973,N_1969);
nand U2001 (N_2001,N_1952,N_1982);
nand U2002 (N_2002,N_1964,N_1975);
and U2003 (N_2003,N_1954,N_1958);
nand U2004 (N_2004,N_1965,N_1986);
nor U2005 (N_2005,N_1990,N_1997);
nor U2006 (N_2006,N_1951,N_1981);
nand U2007 (N_2007,N_1978,N_1992);
or U2008 (N_2008,N_1974,N_1955);
and U2009 (N_2009,N_1961,N_1970);
and U2010 (N_2010,N_1963,N_1995);
nor U2011 (N_2011,N_1959,N_1971);
nor U2012 (N_2012,N_1979,N_1993);
or U2013 (N_2013,N_1980,N_1972);
nor U2014 (N_2014,N_1988,N_1950);
or U2015 (N_2015,N_1968,N_1956);
nand U2016 (N_2016,N_1994,N_1998);
or U2017 (N_2017,N_1976,N_1989);
and U2018 (N_2018,N_1996,N_1960);
nand U2019 (N_2019,N_1953,N_1967);
or U2020 (N_2020,N_1985,N_1962);
and U2021 (N_2021,N_1984,N_1987);
nor U2022 (N_2022,N_1983,N_1957);
nand U2023 (N_2023,N_1977,N_1966);
or U2024 (N_2024,N_1991,N_1999);
nand U2025 (N_2025,N_1962,N_1987);
nor U2026 (N_2026,N_1963,N_1952);
nand U2027 (N_2027,N_1979,N_1969);
and U2028 (N_2028,N_1970,N_1968);
xnor U2029 (N_2029,N_1964,N_1957);
nor U2030 (N_2030,N_1983,N_1982);
and U2031 (N_2031,N_1979,N_1974);
nor U2032 (N_2032,N_1971,N_1966);
or U2033 (N_2033,N_1972,N_1950);
nor U2034 (N_2034,N_1959,N_1987);
nor U2035 (N_2035,N_1977,N_1984);
or U2036 (N_2036,N_1963,N_1986);
nor U2037 (N_2037,N_1968,N_1979);
and U2038 (N_2038,N_1959,N_1984);
or U2039 (N_2039,N_1981,N_1959);
nand U2040 (N_2040,N_1953,N_1999);
or U2041 (N_2041,N_1996,N_1976);
and U2042 (N_2042,N_1975,N_1952);
nor U2043 (N_2043,N_1977,N_1967);
nand U2044 (N_2044,N_1983,N_1985);
nand U2045 (N_2045,N_1995,N_1967);
nand U2046 (N_2046,N_1978,N_1953);
nand U2047 (N_2047,N_1990,N_1982);
and U2048 (N_2048,N_1985,N_1999);
nor U2049 (N_2049,N_1996,N_1991);
and U2050 (N_2050,N_2041,N_2040);
and U2051 (N_2051,N_2010,N_2014);
or U2052 (N_2052,N_2002,N_2022);
or U2053 (N_2053,N_2009,N_2008);
nand U2054 (N_2054,N_2035,N_2037);
nor U2055 (N_2055,N_2016,N_2011);
nor U2056 (N_2056,N_2028,N_2017);
nand U2057 (N_2057,N_2026,N_2025);
nor U2058 (N_2058,N_2018,N_2043);
xnor U2059 (N_2059,N_2045,N_2046);
or U2060 (N_2060,N_2048,N_2042);
and U2061 (N_2061,N_2029,N_2015);
and U2062 (N_2062,N_2032,N_2012);
nor U2063 (N_2063,N_2033,N_2004);
nand U2064 (N_2064,N_2031,N_2039);
nor U2065 (N_2065,N_2036,N_2027);
and U2066 (N_2066,N_2003,N_2019);
or U2067 (N_2067,N_2030,N_2007);
and U2068 (N_2068,N_2047,N_2049);
nor U2069 (N_2069,N_2001,N_2005);
nor U2070 (N_2070,N_2044,N_2021);
xor U2071 (N_2071,N_2013,N_2023);
nand U2072 (N_2072,N_2020,N_2024);
nor U2073 (N_2073,N_2000,N_2034);
and U2074 (N_2074,N_2038,N_2006);
nand U2075 (N_2075,N_2028,N_2045);
and U2076 (N_2076,N_2041,N_2013);
or U2077 (N_2077,N_2021,N_2019);
nand U2078 (N_2078,N_2042,N_2047);
nor U2079 (N_2079,N_2005,N_2039);
nor U2080 (N_2080,N_2024,N_2036);
nor U2081 (N_2081,N_2008,N_2020);
nor U2082 (N_2082,N_2000,N_2007);
or U2083 (N_2083,N_2027,N_2044);
nand U2084 (N_2084,N_2012,N_2025);
nor U2085 (N_2085,N_2000,N_2006);
nor U2086 (N_2086,N_2035,N_2014);
nor U2087 (N_2087,N_2000,N_2030);
nand U2088 (N_2088,N_2040,N_2017);
and U2089 (N_2089,N_2019,N_2022);
nand U2090 (N_2090,N_2034,N_2010);
and U2091 (N_2091,N_2048,N_2002);
and U2092 (N_2092,N_2021,N_2001);
and U2093 (N_2093,N_2025,N_2005);
and U2094 (N_2094,N_2049,N_2042);
nand U2095 (N_2095,N_2046,N_2010);
nor U2096 (N_2096,N_2012,N_2009);
or U2097 (N_2097,N_2016,N_2000);
nor U2098 (N_2098,N_2036,N_2009);
nand U2099 (N_2099,N_2029,N_2019);
nand U2100 (N_2100,N_2087,N_2065);
or U2101 (N_2101,N_2075,N_2061);
nor U2102 (N_2102,N_2082,N_2073);
nand U2103 (N_2103,N_2052,N_2077);
and U2104 (N_2104,N_2069,N_2072);
and U2105 (N_2105,N_2090,N_2094);
nor U2106 (N_2106,N_2068,N_2058);
nand U2107 (N_2107,N_2051,N_2098);
or U2108 (N_2108,N_2060,N_2095);
nand U2109 (N_2109,N_2057,N_2080);
nor U2110 (N_2110,N_2078,N_2096);
nor U2111 (N_2111,N_2088,N_2091);
nor U2112 (N_2112,N_2064,N_2062);
nand U2113 (N_2113,N_2070,N_2099);
or U2114 (N_2114,N_2074,N_2059);
nand U2115 (N_2115,N_2079,N_2076);
and U2116 (N_2116,N_2092,N_2071);
nor U2117 (N_2117,N_2063,N_2086);
or U2118 (N_2118,N_2085,N_2084);
or U2119 (N_2119,N_2055,N_2050);
nor U2120 (N_2120,N_2056,N_2089);
and U2121 (N_2121,N_2093,N_2083);
nor U2122 (N_2122,N_2054,N_2053);
nand U2123 (N_2123,N_2067,N_2081);
nor U2124 (N_2124,N_2097,N_2066);
and U2125 (N_2125,N_2093,N_2096);
and U2126 (N_2126,N_2091,N_2096);
and U2127 (N_2127,N_2065,N_2090);
and U2128 (N_2128,N_2060,N_2064);
nand U2129 (N_2129,N_2087,N_2072);
or U2130 (N_2130,N_2075,N_2087);
nor U2131 (N_2131,N_2053,N_2099);
nor U2132 (N_2132,N_2056,N_2062);
and U2133 (N_2133,N_2079,N_2064);
and U2134 (N_2134,N_2078,N_2091);
nor U2135 (N_2135,N_2052,N_2060);
or U2136 (N_2136,N_2099,N_2067);
or U2137 (N_2137,N_2092,N_2069);
nor U2138 (N_2138,N_2071,N_2099);
nor U2139 (N_2139,N_2090,N_2080);
xor U2140 (N_2140,N_2060,N_2067);
and U2141 (N_2141,N_2076,N_2050);
nand U2142 (N_2142,N_2075,N_2079);
and U2143 (N_2143,N_2061,N_2094);
and U2144 (N_2144,N_2056,N_2079);
or U2145 (N_2145,N_2096,N_2074);
or U2146 (N_2146,N_2072,N_2052);
and U2147 (N_2147,N_2051,N_2088);
nand U2148 (N_2148,N_2064,N_2052);
nand U2149 (N_2149,N_2069,N_2067);
and U2150 (N_2150,N_2128,N_2107);
xor U2151 (N_2151,N_2112,N_2148);
nand U2152 (N_2152,N_2134,N_2138);
xnor U2153 (N_2153,N_2124,N_2136);
and U2154 (N_2154,N_2118,N_2137);
or U2155 (N_2155,N_2133,N_2146);
nand U2156 (N_2156,N_2106,N_2140);
or U2157 (N_2157,N_2139,N_2117);
or U2158 (N_2158,N_2120,N_2126);
nor U2159 (N_2159,N_2110,N_2145);
nand U2160 (N_2160,N_2127,N_2144);
nand U2161 (N_2161,N_2109,N_2141);
or U2162 (N_2162,N_2108,N_2119);
nor U2163 (N_2163,N_2135,N_2122);
nand U2164 (N_2164,N_2121,N_2147);
and U2165 (N_2165,N_2104,N_2142);
and U2166 (N_2166,N_2101,N_2103);
or U2167 (N_2167,N_2100,N_2131);
nand U2168 (N_2168,N_2125,N_2102);
or U2169 (N_2169,N_2130,N_2114);
nand U2170 (N_2170,N_2143,N_2132);
or U2171 (N_2171,N_2111,N_2113);
nor U2172 (N_2172,N_2115,N_2129);
nand U2173 (N_2173,N_2105,N_2149);
nand U2174 (N_2174,N_2116,N_2123);
nand U2175 (N_2175,N_2141,N_2112);
nand U2176 (N_2176,N_2121,N_2107);
nand U2177 (N_2177,N_2109,N_2149);
and U2178 (N_2178,N_2126,N_2117);
xnor U2179 (N_2179,N_2120,N_2114);
nor U2180 (N_2180,N_2143,N_2114);
and U2181 (N_2181,N_2137,N_2146);
nor U2182 (N_2182,N_2109,N_2136);
nor U2183 (N_2183,N_2139,N_2141);
nor U2184 (N_2184,N_2100,N_2137);
nand U2185 (N_2185,N_2113,N_2140);
nand U2186 (N_2186,N_2126,N_2123);
or U2187 (N_2187,N_2134,N_2126);
nand U2188 (N_2188,N_2143,N_2106);
nand U2189 (N_2189,N_2102,N_2134);
nand U2190 (N_2190,N_2132,N_2124);
nand U2191 (N_2191,N_2140,N_2118);
nand U2192 (N_2192,N_2133,N_2123);
and U2193 (N_2193,N_2130,N_2148);
or U2194 (N_2194,N_2114,N_2126);
or U2195 (N_2195,N_2137,N_2107);
nor U2196 (N_2196,N_2130,N_2120);
nand U2197 (N_2197,N_2129,N_2117);
nor U2198 (N_2198,N_2142,N_2117);
nand U2199 (N_2199,N_2124,N_2144);
nor U2200 (N_2200,N_2161,N_2195);
and U2201 (N_2201,N_2150,N_2171);
or U2202 (N_2202,N_2152,N_2198);
nor U2203 (N_2203,N_2160,N_2199);
or U2204 (N_2204,N_2189,N_2154);
or U2205 (N_2205,N_2155,N_2177);
nor U2206 (N_2206,N_2190,N_2159);
nand U2207 (N_2207,N_2188,N_2166);
and U2208 (N_2208,N_2194,N_2158);
or U2209 (N_2209,N_2181,N_2185);
nor U2210 (N_2210,N_2196,N_2187);
or U2211 (N_2211,N_2163,N_2169);
or U2212 (N_2212,N_2193,N_2184);
and U2213 (N_2213,N_2167,N_2175);
and U2214 (N_2214,N_2168,N_2170);
xor U2215 (N_2215,N_2179,N_2183);
nor U2216 (N_2216,N_2173,N_2182);
nor U2217 (N_2217,N_2197,N_2164);
and U2218 (N_2218,N_2157,N_2192);
nand U2219 (N_2219,N_2178,N_2180);
nand U2220 (N_2220,N_2151,N_2172);
or U2221 (N_2221,N_2156,N_2186);
and U2222 (N_2222,N_2191,N_2176);
nand U2223 (N_2223,N_2162,N_2153);
nor U2224 (N_2224,N_2165,N_2174);
nor U2225 (N_2225,N_2187,N_2183);
and U2226 (N_2226,N_2196,N_2179);
and U2227 (N_2227,N_2183,N_2178);
nor U2228 (N_2228,N_2172,N_2166);
and U2229 (N_2229,N_2187,N_2179);
nand U2230 (N_2230,N_2193,N_2158);
and U2231 (N_2231,N_2192,N_2159);
nor U2232 (N_2232,N_2194,N_2170);
nand U2233 (N_2233,N_2185,N_2177);
nor U2234 (N_2234,N_2153,N_2185);
and U2235 (N_2235,N_2192,N_2162);
and U2236 (N_2236,N_2161,N_2163);
and U2237 (N_2237,N_2162,N_2159);
nand U2238 (N_2238,N_2198,N_2163);
and U2239 (N_2239,N_2195,N_2176);
and U2240 (N_2240,N_2171,N_2179);
nor U2241 (N_2241,N_2150,N_2168);
nand U2242 (N_2242,N_2164,N_2192);
or U2243 (N_2243,N_2189,N_2156);
or U2244 (N_2244,N_2197,N_2153);
and U2245 (N_2245,N_2172,N_2188);
and U2246 (N_2246,N_2151,N_2179);
and U2247 (N_2247,N_2156,N_2176);
or U2248 (N_2248,N_2157,N_2185);
nor U2249 (N_2249,N_2179,N_2172);
or U2250 (N_2250,N_2244,N_2204);
nor U2251 (N_2251,N_2205,N_2229);
and U2252 (N_2252,N_2201,N_2247);
nor U2253 (N_2253,N_2239,N_2219);
or U2254 (N_2254,N_2208,N_2231);
xor U2255 (N_2255,N_2236,N_2212);
nor U2256 (N_2256,N_2238,N_2214);
nor U2257 (N_2257,N_2230,N_2249);
and U2258 (N_2258,N_2225,N_2248);
and U2259 (N_2259,N_2211,N_2207);
and U2260 (N_2260,N_2203,N_2215);
and U2261 (N_2261,N_2202,N_2235);
and U2262 (N_2262,N_2240,N_2209);
nor U2263 (N_2263,N_2223,N_2237);
nor U2264 (N_2264,N_2228,N_2232);
and U2265 (N_2265,N_2241,N_2222);
nand U2266 (N_2266,N_2245,N_2233);
nand U2267 (N_2267,N_2200,N_2227);
nor U2268 (N_2268,N_2206,N_2246);
xor U2269 (N_2269,N_2217,N_2234);
and U2270 (N_2270,N_2220,N_2213);
nand U2271 (N_2271,N_2218,N_2216);
nor U2272 (N_2272,N_2243,N_2221);
and U2273 (N_2273,N_2226,N_2242);
nand U2274 (N_2274,N_2210,N_2224);
and U2275 (N_2275,N_2212,N_2214);
nand U2276 (N_2276,N_2235,N_2238);
and U2277 (N_2277,N_2225,N_2220);
nand U2278 (N_2278,N_2229,N_2218);
and U2279 (N_2279,N_2229,N_2200);
nor U2280 (N_2280,N_2208,N_2225);
nor U2281 (N_2281,N_2248,N_2211);
nor U2282 (N_2282,N_2225,N_2205);
or U2283 (N_2283,N_2205,N_2201);
nand U2284 (N_2284,N_2248,N_2222);
and U2285 (N_2285,N_2234,N_2238);
nor U2286 (N_2286,N_2219,N_2235);
or U2287 (N_2287,N_2228,N_2236);
or U2288 (N_2288,N_2233,N_2239);
xnor U2289 (N_2289,N_2219,N_2207);
and U2290 (N_2290,N_2235,N_2232);
and U2291 (N_2291,N_2229,N_2244);
xor U2292 (N_2292,N_2206,N_2203);
nor U2293 (N_2293,N_2245,N_2212);
and U2294 (N_2294,N_2217,N_2218);
nand U2295 (N_2295,N_2204,N_2202);
or U2296 (N_2296,N_2240,N_2204);
and U2297 (N_2297,N_2206,N_2221);
nand U2298 (N_2298,N_2213,N_2226);
or U2299 (N_2299,N_2205,N_2238);
nor U2300 (N_2300,N_2281,N_2274);
nor U2301 (N_2301,N_2276,N_2261);
nand U2302 (N_2302,N_2271,N_2262);
and U2303 (N_2303,N_2279,N_2294);
nor U2304 (N_2304,N_2289,N_2256);
nand U2305 (N_2305,N_2253,N_2287);
or U2306 (N_2306,N_2292,N_2297);
nand U2307 (N_2307,N_2283,N_2286);
or U2308 (N_2308,N_2278,N_2293);
or U2309 (N_2309,N_2258,N_2252);
xnor U2310 (N_2310,N_2251,N_2280);
nor U2311 (N_2311,N_2285,N_2266);
nand U2312 (N_2312,N_2265,N_2288);
or U2313 (N_2313,N_2284,N_2264);
nand U2314 (N_2314,N_2277,N_2299);
nand U2315 (N_2315,N_2267,N_2272);
nor U2316 (N_2316,N_2257,N_2291);
and U2317 (N_2317,N_2250,N_2254);
nand U2318 (N_2318,N_2259,N_2275);
or U2319 (N_2319,N_2296,N_2268);
and U2320 (N_2320,N_2269,N_2255);
or U2321 (N_2321,N_2273,N_2270);
nor U2322 (N_2322,N_2260,N_2263);
and U2323 (N_2323,N_2298,N_2290);
and U2324 (N_2324,N_2295,N_2282);
nor U2325 (N_2325,N_2262,N_2250);
xnor U2326 (N_2326,N_2262,N_2269);
nor U2327 (N_2327,N_2254,N_2294);
nor U2328 (N_2328,N_2272,N_2250);
nand U2329 (N_2329,N_2293,N_2266);
and U2330 (N_2330,N_2259,N_2254);
or U2331 (N_2331,N_2277,N_2295);
nor U2332 (N_2332,N_2273,N_2274);
and U2333 (N_2333,N_2264,N_2274);
or U2334 (N_2334,N_2279,N_2277);
nor U2335 (N_2335,N_2290,N_2266);
nand U2336 (N_2336,N_2252,N_2266);
or U2337 (N_2337,N_2273,N_2262);
and U2338 (N_2338,N_2289,N_2277);
nand U2339 (N_2339,N_2282,N_2269);
and U2340 (N_2340,N_2298,N_2263);
or U2341 (N_2341,N_2277,N_2266);
nor U2342 (N_2342,N_2299,N_2266);
xnor U2343 (N_2343,N_2278,N_2286);
nand U2344 (N_2344,N_2255,N_2274);
nor U2345 (N_2345,N_2267,N_2260);
nor U2346 (N_2346,N_2261,N_2259);
nor U2347 (N_2347,N_2259,N_2295);
or U2348 (N_2348,N_2277,N_2255);
and U2349 (N_2349,N_2299,N_2290);
nand U2350 (N_2350,N_2319,N_2347);
or U2351 (N_2351,N_2335,N_2302);
nor U2352 (N_2352,N_2321,N_2325);
nand U2353 (N_2353,N_2349,N_2345);
or U2354 (N_2354,N_2315,N_2344);
and U2355 (N_2355,N_2308,N_2327);
nand U2356 (N_2356,N_2300,N_2317);
or U2357 (N_2357,N_2314,N_2316);
nand U2358 (N_2358,N_2337,N_2318);
or U2359 (N_2359,N_2322,N_2346);
or U2360 (N_2360,N_2343,N_2348);
nand U2361 (N_2361,N_2334,N_2305);
and U2362 (N_2362,N_2303,N_2332);
and U2363 (N_2363,N_2331,N_2328);
nor U2364 (N_2364,N_2323,N_2304);
nand U2365 (N_2365,N_2341,N_2340);
nand U2366 (N_2366,N_2312,N_2313);
and U2367 (N_2367,N_2311,N_2338);
or U2368 (N_2368,N_2339,N_2310);
and U2369 (N_2369,N_2324,N_2336);
and U2370 (N_2370,N_2307,N_2329);
nor U2371 (N_2371,N_2326,N_2309);
nor U2372 (N_2372,N_2342,N_2333);
nor U2373 (N_2373,N_2306,N_2301);
nor U2374 (N_2374,N_2330,N_2320);
and U2375 (N_2375,N_2307,N_2337);
nand U2376 (N_2376,N_2325,N_2333);
and U2377 (N_2377,N_2340,N_2306);
and U2378 (N_2378,N_2335,N_2334);
or U2379 (N_2379,N_2325,N_2324);
and U2380 (N_2380,N_2308,N_2320);
and U2381 (N_2381,N_2316,N_2308);
nor U2382 (N_2382,N_2334,N_2331);
or U2383 (N_2383,N_2324,N_2322);
nor U2384 (N_2384,N_2340,N_2318);
nand U2385 (N_2385,N_2313,N_2315);
and U2386 (N_2386,N_2331,N_2309);
nor U2387 (N_2387,N_2312,N_2306);
nor U2388 (N_2388,N_2349,N_2311);
or U2389 (N_2389,N_2340,N_2342);
nand U2390 (N_2390,N_2327,N_2302);
or U2391 (N_2391,N_2341,N_2332);
nand U2392 (N_2392,N_2332,N_2333);
and U2393 (N_2393,N_2333,N_2315);
and U2394 (N_2394,N_2334,N_2319);
nor U2395 (N_2395,N_2323,N_2300);
nand U2396 (N_2396,N_2319,N_2341);
nand U2397 (N_2397,N_2322,N_2341);
and U2398 (N_2398,N_2301,N_2342);
or U2399 (N_2399,N_2347,N_2349);
nor U2400 (N_2400,N_2366,N_2384);
or U2401 (N_2401,N_2359,N_2368);
and U2402 (N_2402,N_2367,N_2399);
and U2403 (N_2403,N_2396,N_2398);
xnor U2404 (N_2404,N_2389,N_2355);
and U2405 (N_2405,N_2387,N_2388);
nand U2406 (N_2406,N_2379,N_2358);
nor U2407 (N_2407,N_2361,N_2362);
nor U2408 (N_2408,N_2352,N_2385);
nand U2409 (N_2409,N_2394,N_2357);
nand U2410 (N_2410,N_2380,N_2354);
nor U2411 (N_2411,N_2372,N_2356);
or U2412 (N_2412,N_2397,N_2369);
and U2413 (N_2413,N_2383,N_2373);
and U2414 (N_2414,N_2391,N_2390);
and U2415 (N_2415,N_2375,N_2374);
or U2416 (N_2416,N_2377,N_2350);
nor U2417 (N_2417,N_2378,N_2376);
nor U2418 (N_2418,N_2386,N_2392);
and U2419 (N_2419,N_2363,N_2370);
and U2420 (N_2420,N_2353,N_2395);
nor U2421 (N_2421,N_2351,N_2381);
nor U2422 (N_2422,N_2360,N_2382);
or U2423 (N_2423,N_2365,N_2393);
or U2424 (N_2424,N_2364,N_2371);
nor U2425 (N_2425,N_2380,N_2364);
and U2426 (N_2426,N_2375,N_2396);
nand U2427 (N_2427,N_2364,N_2393);
nand U2428 (N_2428,N_2384,N_2396);
or U2429 (N_2429,N_2361,N_2360);
and U2430 (N_2430,N_2387,N_2369);
or U2431 (N_2431,N_2374,N_2377);
nand U2432 (N_2432,N_2364,N_2360);
or U2433 (N_2433,N_2397,N_2375);
nor U2434 (N_2434,N_2365,N_2399);
nor U2435 (N_2435,N_2358,N_2368);
nor U2436 (N_2436,N_2375,N_2355);
nand U2437 (N_2437,N_2391,N_2363);
or U2438 (N_2438,N_2396,N_2389);
nor U2439 (N_2439,N_2360,N_2393);
nand U2440 (N_2440,N_2387,N_2356);
nand U2441 (N_2441,N_2356,N_2360);
nor U2442 (N_2442,N_2384,N_2375);
nor U2443 (N_2443,N_2353,N_2364);
xnor U2444 (N_2444,N_2363,N_2368);
and U2445 (N_2445,N_2351,N_2397);
and U2446 (N_2446,N_2372,N_2364);
nand U2447 (N_2447,N_2368,N_2351);
nor U2448 (N_2448,N_2392,N_2383);
or U2449 (N_2449,N_2358,N_2378);
nand U2450 (N_2450,N_2445,N_2441);
nand U2451 (N_2451,N_2407,N_2438);
xor U2452 (N_2452,N_2439,N_2400);
nor U2453 (N_2453,N_2410,N_2406);
and U2454 (N_2454,N_2403,N_2415);
nand U2455 (N_2455,N_2433,N_2448);
or U2456 (N_2456,N_2419,N_2430);
and U2457 (N_2457,N_2425,N_2449);
nor U2458 (N_2458,N_2404,N_2440);
or U2459 (N_2459,N_2409,N_2416);
and U2460 (N_2460,N_2421,N_2401);
or U2461 (N_2461,N_2426,N_2432);
and U2462 (N_2462,N_2436,N_2424);
nor U2463 (N_2463,N_2434,N_2412);
nand U2464 (N_2464,N_2446,N_2408);
nand U2465 (N_2465,N_2422,N_2442);
or U2466 (N_2466,N_2429,N_2411);
or U2467 (N_2467,N_2437,N_2428);
and U2468 (N_2468,N_2414,N_2423);
nor U2469 (N_2469,N_2444,N_2427);
nand U2470 (N_2470,N_2447,N_2431);
nor U2471 (N_2471,N_2420,N_2417);
or U2472 (N_2472,N_2405,N_2402);
and U2473 (N_2473,N_2418,N_2413);
or U2474 (N_2474,N_2435,N_2443);
xnor U2475 (N_2475,N_2423,N_2444);
nor U2476 (N_2476,N_2411,N_2409);
and U2477 (N_2477,N_2424,N_2415);
nand U2478 (N_2478,N_2408,N_2444);
and U2479 (N_2479,N_2419,N_2440);
and U2480 (N_2480,N_2427,N_2439);
or U2481 (N_2481,N_2434,N_2436);
nand U2482 (N_2482,N_2432,N_2420);
nor U2483 (N_2483,N_2441,N_2405);
nand U2484 (N_2484,N_2411,N_2446);
nor U2485 (N_2485,N_2402,N_2415);
nand U2486 (N_2486,N_2405,N_2416);
nand U2487 (N_2487,N_2419,N_2414);
nor U2488 (N_2488,N_2433,N_2431);
or U2489 (N_2489,N_2425,N_2443);
nor U2490 (N_2490,N_2407,N_2443);
nor U2491 (N_2491,N_2444,N_2424);
or U2492 (N_2492,N_2427,N_2433);
or U2493 (N_2493,N_2438,N_2413);
nor U2494 (N_2494,N_2447,N_2426);
and U2495 (N_2495,N_2429,N_2405);
or U2496 (N_2496,N_2431,N_2445);
nor U2497 (N_2497,N_2423,N_2418);
nor U2498 (N_2498,N_2425,N_2402);
nor U2499 (N_2499,N_2428,N_2430);
and U2500 (N_2500,N_2454,N_2477);
nor U2501 (N_2501,N_2478,N_2489);
or U2502 (N_2502,N_2496,N_2479);
nor U2503 (N_2503,N_2460,N_2453);
or U2504 (N_2504,N_2487,N_2486);
nor U2505 (N_2505,N_2458,N_2463);
nor U2506 (N_2506,N_2473,N_2495);
and U2507 (N_2507,N_2459,N_2456);
or U2508 (N_2508,N_2499,N_2474);
or U2509 (N_2509,N_2465,N_2468);
or U2510 (N_2510,N_2467,N_2452);
and U2511 (N_2511,N_2482,N_2464);
nand U2512 (N_2512,N_2494,N_2466);
or U2513 (N_2513,N_2470,N_2471);
nor U2514 (N_2514,N_2455,N_2483);
and U2515 (N_2515,N_2492,N_2498);
xnor U2516 (N_2516,N_2461,N_2472);
xnor U2517 (N_2517,N_2491,N_2469);
or U2518 (N_2518,N_2484,N_2451);
and U2519 (N_2519,N_2462,N_2457);
nor U2520 (N_2520,N_2450,N_2480);
nor U2521 (N_2521,N_2488,N_2493);
nand U2522 (N_2522,N_2497,N_2485);
nand U2523 (N_2523,N_2481,N_2475);
nand U2524 (N_2524,N_2476,N_2490);
nand U2525 (N_2525,N_2453,N_2466);
nand U2526 (N_2526,N_2488,N_2477);
nand U2527 (N_2527,N_2496,N_2459);
nor U2528 (N_2528,N_2464,N_2465);
and U2529 (N_2529,N_2489,N_2462);
nor U2530 (N_2530,N_2477,N_2489);
or U2531 (N_2531,N_2485,N_2470);
and U2532 (N_2532,N_2464,N_2454);
nand U2533 (N_2533,N_2470,N_2476);
nand U2534 (N_2534,N_2495,N_2454);
nand U2535 (N_2535,N_2467,N_2451);
nor U2536 (N_2536,N_2497,N_2495);
and U2537 (N_2537,N_2458,N_2451);
nor U2538 (N_2538,N_2495,N_2484);
or U2539 (N_2539,N_2497,N_2490);
and U2540 (N_2540,N_2492,N_2475);
nand U2541 (N_2541,N_2451,N_2494);
or U2542 (N_2542,N_2495,N_2498);
nand U2543 (N_2543,N_2486,N_2469);
and U2544 (N_2544,N_2451,N_2465);
and U2545 (N_2545,N_2459,N_2458);
nand U2546 (N_2546,N_2499,N_2492);
and U2547 (N_2547,N_2462,N_2486);
and U2548 (N_2548,N_2466,N_2462);
nand U2549 (N_2549,N_2498,N_2482);
nor U2550 (N_2550,N_2548,N_2531);
nand U2551 (N_2551,N_2523,N_2517);
or U2552 (N_2552,N_2540,N_2542);
nor U2553 (N_2553,N_2518,N_2545);
nand U2554 (N_2554,N_2546,N_2526);
nor U2555 (N_2555,N_2524,N_2505);
nand U2556 (N_2556,N_2513,N_2516);
nand U2557 (N_2557,N_2514,N_2543);
nor U2558 (N_2558,N_2538,N_2507);
or U2559 (N_2559,N_2537,N_2549);
and U2560 (N_2560,N_2512,N_2519);
nor U2561 (N_2561,N_2520,N_2533);
nand U2562 (N_2562,N_2515,N_2541);
xor U2563 (N_2563,N_2532,N_2535);
nand U2564 (N_2564,N_2528,N_2500);
or U2565 (N_2565,N_2529,N_2530);
nor U2566 (N_2566,N_2525,N_2547);
and U2567 (N_2567,N_2522,N_2544);
and U2568 (N_2568,N_2539,N_2536);
nor U2569 (N_2569,N_2502,N_2501);
nand U2570 (N_2570,N_2504,N_2509);
nand U2571 (N_2571,N_2508,N_2527);
nand U2572 (N_2572,N_2521,N_2510);
or U2573 (N_2573,N_2534,N_2506);
nand U2574 (N_2574,N_2503,N_2511);
nand U2575 (N_2575,N_2545,N_2501);
nand U2576 (N_2576,N_2511,N_2520);
nor U2577 (N_2577,N_2516,N_2539);
nor U2578 (N_2578,N_2504,N_2537);
nor U2579 (N_2579,N_2518,N_2527);
nand U2580 (N_2580,N_2549,N_2520);
xnor U2581 (N_2581,N_2525,N_2545);
or U2582 (N_2582,N_2515,N_2531);
or U2583 (N_2583,N_2541,N_2512);
xor U2584 (N_2584,N_2517,N_2548);
nand U2585 (N_2585,N_2514,N_2548);
nand U2586 (N_2586,N_2522,N_2538);
and U2587 (N_2587,N_2546,N_2515);
and U2588 (N_2588,N_2519,N_2532);
nor U2589 (N_2589,N_2529,N_2543);
nand U2590 (N_2590,N_2510,N_2535);
nand U2591 (N_2591,N_2501,N_2547);
and U2592 (N_2592,N_2513,N_2537);
and U2593 (N_2593,N_2521,N_2518);
or U2594 (N_2594,N_2544,N_2505);
nor U2595 (N_2595,N_2530,N_2528);
nand U2596 (N_2596,N_2522,N_2520);
or U2597 (N_2597,N_2538,N_2505);
and U2598 (N_2598,N_2528,N_2521);
nand U2599 (N_2599,N_2529,N_2500);
nand U2600 (N_2600,N_2568,N_2598);
nor U2601 (N_2601,N_2583,N_2586);
or U2602 (N_2602,N_2591,N_2551);
nor U2603 (N_2603,N_2577,N_2560);
and U2604 (N_2604,N_2590,N_2584);
nor U2605 (N_2605,N_2593,N_2578);
nand U2606 (N_2606,N_2565,N_2595);
nor U2607 (N_2607,N_2553,N_2561);
xnor U2608 (N_2608,N_2564,N_2589);
or U2609 (N_2609,N_2588,N_2582);
nor U2610 (N_2610,N_2554,N_2563);
or U2611 (N_2611,N_2573,N_2571);
nor U2612 (N_2612,N_2570,N_2552);
and U2613 (N_2613,N_2585,N_2562);
or U2614 (N_2614,N_2579,N_2576);
nor U2615 (N_2615,N_2556,N_2575);
or U2616 (N_2616,N_2572,N_2555);
or U2617 (N_2617,N_2592,N_2557);
or U2618 (N_2618,N_2566,N_2594);
and U2619 (N_2619,N_2580,N_2569);
or U2620 (N_2620,N_2581,N_2574);
nor U2621 (N_2621,N_2596,N_2567);
nor U2622 (N_2622,N_2599,N_2559);
and U2623 (N_2623,N_2550,N_2587);
and U2624 (N_2624,N_2597,N_2558);
nor U2625 (N_2625,N_2573,N_2587);
or U2626 (N_2626,N_2557,N_2555);
or U2627 (N_2627,N_2594,N_2575);
nor U2628 (N_2628,N_2558,N_2563);
nand U2629 (N_2629,N_2556,N_2560);
xnor U2630 (N_2630,N_2570,N_2584);
nor U2631 (N_2631,N_2553,N_2589);
nor U2632 (N_2632,N_2574,N_2561);
or U2633 (N_2633,N_2551,N_2572);
nand U2634 (N_2634,N_2583,N_2552);
nor U2635 (N_2635,N_2563,N_2598);
nand U2636 (N_2636,N_2580,N_2581);
and U2637 (N_2637,N_2565,N_2555);
and U2638 (N_2638,N_2575,N_2568);
and U2639 (N_2639,N_2552,N_2592);
nor U2640 (N_2640,N_2557,N_2566);
and U2641 (N_2641,N_2596,N_2571);
nor U2642 (N_2642,N_2587,N_2552);
or U2643 (N_2643,N_2551,N_2590);
and U2644 (N_2644,N_2561,N_2571);
xnor U2645 (N_2645,N_2575,N_2561);
nor U2646 (N_2646,N_2582,N_2584);
or U2647 (N_2647,N_2596,N_2553);
nand U2648 (N_2648,N_2590,N_2582);
nand U2649 (N_2649,N_2580,N_2583);
nand U2650 (N_2650,N_2616,N_2628);
nand U2651 (N_2651,N_2615,N_2626);
xnor U2652 (N_2652,N_2621,N_2611);
or U2653 (N_2653,N_2605,N_2624);
nand U2654 (N_2654,N_2608,N_2601);
and U2655 (N_2655,N_2646,N_2640);
and U2656 (N_2656,N_2630,N_2600);
nand U2657 (N_2657,N_2643,N_2613);
nand U2658 (N_2658,N_2610,N_2607);
nand U2659 (N_2659,N_2645,N_2636);
nor U2660 (N_2660,N_2634,N_2629);
or U2661 (N_2661,N_2633,N_2638);
nand U2662 (N_2662,N_2625,N_2641);
nor U2663 (N_2663,N_2618,N_2644);
and U2664 (N_2664,N_2649,N_2637);
or U2665 (N_2665,N_2623,N_2604);
nor U2666 (N_2666,N_2647,N_2631);
and U2667 (N_2667,N_2639,N_2602);
nor U2668 (N_2668,N_2632,N_2606);
nand U2669 (N_2669,N_2617,N_2622);
nand U2670 (N_2670,N_2642,N_2603);
nand U2671 (N_2671,N_2619,N_2635);
and U2672 (N_2672,N_2620,N_2627);
nand U2673 (N_2673,N_2609,N_2614);
nor U2674 (N_2674,N_2648,N_2612);
nand U2675 (N_2675,N_2623,N_2614);
or U2676 (N_2676,N_2600,N_2641);
nand U2677 (N_2677,N_2640,N_2610);
and U2678 (N_2678,N_2617,N_2625);
nor U2679 (N_2679,N_2635,N_2639);
and U2680 (N_2680,N_2625,N_2647);
or U2681 (N_2681,N_2629,N_2644);
nor U2682 (N_2682,N_2622,N_2635);
or U2683 (N_2683,N_2648,N_2649);
nor U2684 (N_2684,N_2602,N_2624);
nor U2685 (N_2685,N_2612,N_2623);
xnor U2686 (N_2686,N_2646,N_2648);
nor U2687 (N_2687,N_2640,N_2606);
nor U2688 (N_2688,N_2642,N_2609);
nor U2689 (N_2689,N_2646,N_2608);
nor U2690 (N_2690,N_2629,N_2649);
and U2691 (N_2691,N_2625,N_2604);
nand U2692 (N_2692,N_2648,N_2630);
nor U2693 (N_2693,N_2643,N_2602);
nand U2694 (N_2694,N_2625,N_2632);
nand U2695 (N_2695,N_2628,N_2629);
nand U2696 (N_2696,N_2640,N_2607);
nand U2697 (N_2697,N_2625,N_2602);
nand U2698 (N_2698,N_2616,N_2604);
nor U2699 (N_2699,N_2624,N_2649);
or U2700 (N_2700,N_2650,N_2697);
nor U2701 (N_2701,N_2685,N_2674);
nor U2702 (N_2702,N_2671,N_2679);
or U2703 (N_2703,N_2693,N_2688);
nand U2704 (N_2704,N_2678,N_2699);
and U2705 (N_2705,N_2672,N_2651);
nor U2706 (N_2706,N_2663,N_2691);
and U2707 (N_2707,N_2670,N_2698);
nor U2708 (N_2708,N_2669,N_2683);
or U2709 (N_2709,N_2686,N_2653);
and U2710 (N_2710,N_2665,N_2680);
and U2711 (N_2711,N_2690,N_2682);
or U2712 (N_2712,N_2667,N_2656);
or U2713 (N_2713,N_2652,N_2668);
nor U2714 (N_2714,N_2657,N_2673);
or U2715 (N_2715,N_2681,N_2689);
nor U2716 (N_2716,N_2675,N_2692);
or U2717 (N_2717,N_2658,N_2684);
nor U2718 (N_2718,N_2655,N_2661);
and U2719 (N_2719,N_2654,N_2687);
or U2720 (N_2720,N_2694,N_2676);
nor U2721 (N_2721,N_2660,N_2659);
or U2722 (N_2722,N_2662,N_2677);
or U2723 (N_2723,N_2696,N_2695);
nand U2724 (N_2724,N_2666,N_2664);
and U2725 (N_2725,N_2674,N_2657);
and U2726 (N_2726,N_2650,N_2661);
or U2727 (N_2727,N_2658,N_2686);
nand U2728 (N_2728,N_2696,N_2684);
nor U2729 (N_2729,N_2696,N_2669);
nor U2730 (N_2730,N_2679,N_2675);
and U2731 (N_2731,N_2665,N_2658);
or U2732 (N_2732,N_2671,N_2699);
nand U2733 (N_2733,N_2690,N_2683);
nand U2734 (N_2734,N_2663,N_2654);
nor U2735 (N_2735,N_2677,N_2698);
nor U2736 (N_2736,N_2691,N_2680);
and U2737 (N_2737,N_2658,N_2659);
nand U2738 (N_2738,N_2685,N_2670);
and U2739 (N_2739,N_2652,N_2698);
nor U2740 (N_2740,N_2695,N_2650);
and U2741 (N_2741,N_2686,N_2650);
or U2742 (N_2742,N_2690,N_2673);
and U2743 (N_2743,N_2685,N_2678);
nand U2744 (N_2744,N_2676,N_2685);
and U2745 (N_2745,N_2651,N_2667);
nand U2746 (N_2746,N_2686,N_2685);
or U2747 (N_2747,N_2681,N_2698);
or U2748 (N_2748,N_2674,N_2675);
nand U2749 (N_2749,N_2679,N_2665);
and U2750 (N_2750,N_2712,N_2727);
and U2751 (N_2751,N_2710,N_2717);
or U2752 (N_2752,N_2713,N_2744);
and U2753 (N_2753,N_2738,N_2745);
and U2754 (N_2754,N_2718,N_2721);
nand U2755 (N_2755,N_2736,N_2728);
or U2756 (N_2756,N_2707,N_2743);
or U2757 (N_2757,N_2739,N_2716);
nand U2758 (N_2758,N_2723,N_2725);
nor U2759 (N_2759,N_2700,N_2734);
or U2760 (N_2760,N_2708,N_2735);
nor U2761 (N_2761,N_2737,N_2715);
nand U2762 (N_2762,N_2731,N_2733);
or U2763 (N_2763,N_2741,N_2701);
nor U2764 (N_2764,N_2719,N_2729);
nor U2765 (N_2765,N_2704,N_2742);
and U2766 (N_2766,N_2722,N_2711);
or U2767 (N_2767,N_2747,N_2732);
nor U2768 (N_2768,N_2709,N_2706);
nand U2769 (N_2769,N_2749,N_2705);
nor U2770 (N_2770,N_2714,N_2702);
and U2771 (N_2771,N_2740,N_2726);
nor U2772 (N_2772,N_2746,N_2730);
or U2773 (N_2773,N_2724,N_2703);
and U2774 (N_2774,N_2748,N_2720);
nor U2775 (N_2775,N_2735,N_2745);
or U2776 (N_2776,N_2741,N_2716);
nor U2777 (N_2777,N_2746,N_2719);
nor U2778 (N_2778,N_2718,N_2742);
nand U2779 (N_2779,N_2729,N_2735);
nor U2780 (N_2780,N_2729,N_2705);
nor U2781 (N_2781,N_2744,N_2719);
nor U2782 (N_2782,N_2727,N_2721);
nand U2783 (N_2783,N_2724,N_2737);
nor U2784 (N_2784,N_2741,N_2721);
and U2785 (N_2785,N_2736,N_2729);
nor U2786 (N_2786,N_2723,N_2707);
or U2787 (N_2787,N_2712,N_2741);
nand U2788 (N_2788,N_2740,N_2730);
nand U2789 (N_2789,N_2701,N_2704);
or U2790 (N_2790,N_2700,N_2702);
and U2791 (N_2791,N_2702,N_2736);
or U2792 (N_2792,N_2739,N_2741);
and U2793 (N_2793,N_2708,N_2744);
nor U2794 (N_2794,N_2726,N_2712);
xnor U2795 (N_2795,N_2718,N_2708);
or U2796 (N_2796,N_2702,N_2705);
nand U2797 (N_2797,N_2700,N_2737);
and U2798 (N_2798,N_2708,N_2737);
nor U2799 (N_2799,N_2719,N_2749);
nand U2800 (N_2800,N_2782,N_2795);
nand U2801 (N_2801,N_2792,N_2794);
and U2802 (N_2802,N_2751,N_2750);
or U2803 (N_2803,N_2796,N_2773);
nor U2804 (N_2804,N_2772,N_2754);
or U2805 (N_2805,N_2780,N_2769);
or U2806 (N_2806,N_2771,N_2784);
nor U2807 (N_2807,N_2783,N_2757);
nor U2808 (N_2808,N_2761,N_2766);
and U2809 (N_2809,N_2774,N_2787);
nor U2810 (N_2810,N_2793,N_2791);
or U2811 (N_2811,N_2785,N_2798);
nor U2812 (N_2812,N_2760,N_2762);
nand U2813 (N_2813,N_2770,N_2763);
nand U2814 (N_2814,N_2781,N_2758);
nor U2815 (N_2815,N_2786,N_2759);
nand U2816 (N_2816,N_2755,N_2799);
nand U2817 (N_2817,N_2776,N_2788);
and U2818 (N_2818,N_2764,N_2778);
or U2819 (N_2819,N_2789,N_2752);
and U2820 (N_2820,N_2756,N_2775);
or U2821 (N_2821,N_2767,N_2768);
nor U2822 (N_2822,N_2753,N_2790);
nand U2823 (N_2823,N_2765,N_2797);
nand U2824 (N_2824,N_2779,N_2777);
or U2825 (N_2825,N_2760,N_2777);
nor U2826 (N_2826,N_2762,N_2779);
or U2827 (N_2827,N_2751,N_2759);
nor U2828 (N_2828,N_2791,N_2768);
and U2829 (N_2829,N_2782,N_2770);
and U2830 (N_2830,N_2782,N_2790);
and U2831 (N_2831,N_2770,N_2760);
and U2832 (N_2832,N_2781,N_2754);
and U2833 (N_2833,N_2763,N_2795);
nand U2834 (N_2834,N_2788,N_2799);
nor U2835 (N_2835,N_2794,N_2765);
or U2836 (N_2836,N_2782,N_2759);
nor U2837 (N_2837,N_2795,N_2755);
nand U2838 (N_2838,N_2779,N_2781);
nor U2839 (N_2839,N_2794,N_2786);
or U2840 (N_2840,N_2761,N_2759);
nand U2841 (N_2841,N_2795,N_2779);
nand U2842 (N_2842,N_2778,N_2780);
and U2843 (N_2843,N_2756,N_2752);
or U2844 (N_2844,N_2797,N_2770);
and U2845 (N_2845,N_2795,N_2788);
or U2846 (N_2846,N_2784,N_2793);
or U2847 (N_2847,N_2792,N_2768);
and U2848 (N_2848,N_2767,N_2791);
nor U2849 (N_2849,N_2760,N_2795);
and U2850 (N_2850,N_2847,N_2825);
nand U2851 (N_2851,N_2803,N_2806);
nand U2852 (N_2852,N_2845,N_2832);
nand U2853 (N_2853,N_2823,N_2842);
or U2854 (N_2854,N_2801,N_2827);
xor U2855 (N_2855,N_2846,N_2811);
nand U2856 (N_2856,N_2841,N_2821);
and U2857 (N_2857,N_2819,N_2835);
and U2858 (N_2858,N_2834,N_2818);
nand U2859 (N_2859,N_2804,N_2830);
nand U2860 (N_2860,N_2807,N_2820);
nand U2861 (N_2861,N_2826,N_2849);
or U2862 (N_2862,N_2800,N_2815);
nor U2863 (N_2863,N_2838,N_2822);
nor U2864 (N_2864,N_2840,N_2814);
nand U2865 (N_2865,N_2833,N_2843);
nor U2866 (N_2866,N_2836,N_2831);
or U2867 (N_2867,N_2802,N_2816);
and U2868 (N_2868,N_2812,N_2808);
nand U2869 (N_2869,N_2828,N_2810);
or U2870 (N_2870,N_2809,N_2829);
or U2871 (N_2871,N_2848,N_2837);
or U2872 (N_2872,N_2805,N_2817);
nor U2873 (N_2873,N_2839,N_2813);
or U2874 (N_2874,N_2824,N_2844);
or U2875 (N_2875,N_2811,N_2807);
and U2876 (N_2876,N_2800,N_2845);
nand U2877 (N_2877,N_2832,N_2848);
or U2878 (N_2878,N_2820,N_2843);
nand U2879 (N_2879,N_2821,N_2830);
and U2880 (N_2880,N_2808,N_2843);
or U2881 (N_2881,N_2820,N_2838);
or U2882 (N_2882,N_2818,N_2808);
and U2883 (N_2883,N_2827,N_2821);
or U2884 (N_2884,N_2810,N_2803);
or U2885 (N_2885,N_2807,N_2821);
or U2886 (N_2886,N_2827,N_2813);
and U2887 (N_2887,N_2830,N_2824);
nor U2888 (N_2888,N_2829,N_2810);
and U2889 (N_2889,N_2821,N_2817);
nand U2890 (N_2890,N_2847,N_2826);
nand U2891 (N_2891,N_2822,N_2807);
or U2892 (N_2892,N_2818,N_2839);
and U2893 (N_2893,N_2811,N_2809);
nand U2894 (N_2894,N_2839,N_2802);
nand U2895 (N_2895,N_2834,N_2832);
nand U2896 (N_2896,N_2804,N_2849);
nand U2897 (N_2897,N_2834,N_2833);
nor U2898 (N_2898,N_2833,N_2809);
or U2899 (N_2899,N_2831,N_2809);
nand U2900 (N_2900,N_2889,N_2861);
nor U2901 (N_2901,N_2898,N_2864);
and U2902 (N_2902,N_2892,N_2881);
and U2903 (N_2903,N_2867,N_2872);
nand U2904 (N_2904,N_2860,N_2897);
nand U2905 (N_2905,N_2852,N_2862);
and U2906 (N_2906,N_2888,N_2869);
nor U2907 (N_2907,N_2858,N_2871);
nand U2908 (N_2908,N_2891,N_2857);
nand U2909 (N_2909,N_2895,N_2887);
and U2910 (N_2910,N_2859,N_2882);
nand U2911 (N_2911,N_2883,N_2878);
or U2912 (N_2912,N_2853,N_2863);
and U2913 (N_2913,N_2884,N_2893);
and U2914 (N_2914,N_2880,N_2885);
nand U2915 (N_2915,N_2850,N_2856);
nand U2916 (N_2916,N_2877,N_2870);
and U2917 (N_2917,N_2875,N_2890);
or U2918 (N_2918,N_2899,N_2866);
or U2919 (N_2919,N_2896,N_2854);
and U2920 (N_2920,N_2894,N_2879);
nand U2921 (N_2921,N_2851,N_2865);
and U2922 (N_2922,N_2855,N_2876);
and U2923 (N_2923,N_2874,N_2873);
nand U2924 (N_2924,N_2868,N_2886);
nor U2925 (N_2925,N_2881,N_2860);
and U2926 (N_2926,N_2857,N_2875);
nand U2927 (N_2927,N_2885,N_2855);
nand U2928 (N_2928,N_2857,N_2867);
or U2929 (N_2929,N_2860,N_2855);
nor U2930 (N_2930,N_2862,N_2856);
and U2931 (N_2931,N_2882,N_2870);
nand U2932 (N_2932,N_2894,N_2896);
xor U2933 (N_2933,N_2852,N_2853);
nand U2934 (N_2934,N_2864,N_2857);
or U2935 (N_2935,N_2850,N_2897);
nor U2936 (N_2936,N_2863,N_2884);
nand U2937 (N_2937,N_2894,N_2856);
and U2938 (N_2938,N_2864,N_2871);
nand U2939 (N_2939,N_2865,N_2875);
nand U2940 (N_2940,N_2875,N_2864);
nand U2941 (N_2941,N_2853,N_2871);
xor U2942 (N_2942,N_2879,N_2892);
or U2943 (N_2943,N_2857,N_2878);
or U2944 (N_2944,N_2864,N_2899);
and U2945 (N_2945,N_2871,N_2869);
nor U2946 (N_2946,N_2887,N_2873);
nor U2947 (N_2947,N_2857,N_2894);
and U2948 (N_2948,N_2898,N_2891);
nor U2949 (N_2949,N_2869,N_2896);
xnor U2950 (N_2950,N_2929,N_2946);
nand U2951 (N_2951,N_2931,N_2940);
or U2952 (N_2952,N_2910,N_2934);
or U2953 (N_2953,N_2937,N_2941);
and U2954 (N_2954,N_2913,N_2905);
or U2955 (N_2955,N_2935,N_2906);
and U2956 (N_2956,N_2949,N_2932);
or U2957 (N_2957,N_2924,N_2902);
and U2958 (N_2958,N_2919,N_2936);
or U2959 (N_2959,N_2914,N_2926);
nand U2960 (N_2960,N_2930,N_2928);
nand U2961 (N_2961,N_2912,N_2944);
xor U2962 (N_2962,N_2942,N_2901);
and U2963 (N_2963,N_2917,N_2939);
nor U2964 (N_2964,N_2904,N_2921);
or U2965 (N_2965,N_2909,N_2916);
nor U2966 (N_2966,N_2933,N_2903);
and U2967 (N_2967,N_2938,N_2911);
or U2968 (N_2968,N_2920,N_2943);
and U2969 (N_2969,N_2907,N_2948);
nand U2970 (N_2970,N_2908,N_2947);
and U2971 (N_2971,N_2927,N_2945);
and U2972 (N_2972,N_2915,N_2900);
nor U2973 (N_2973,N_2925,N_2923);
nor U2974 (N_2974,N_2918,N_2922);
or U2975 (N_2975,N_2923,N_2924);
and U2976 (N_2976,N_2943,N_2941);
and U2977 (N_2977,N_2911,N_2922);
nor U2978 (N_2978,N_2917,N_2904);
xor U2979 (N_2979,N_2927,N_2910);
nand U2980 (N_2980,N_2916,N_2923);
nand U2981 (N_2981,N_2911,N_2915);
or U2982 (N_2982,N_2947,N_2923);
nor U2983 (N_2983,N_2914,N_2939);
nand U2984 (N_2984,N_2937,N_2938);
nand U2985 (N_2985,N_2903,N_2932);
nand U2986 (N_2986,N_2944,N_2927);
or U2987 (N_2987,N_2935,N_2923);
nand U2988 (N_2988,N_2915,N_2919);
or U2989 (N_2989,N_2906,N_2943);
or U2990 (N_2990,N_2931,N_2901);
nor U2991 (N_2991,N_2948,N_2911);
nor U2992 (N_2992,N_2920,N_2924);
and U2993 (N_2993,N_2938,N_2936);
nor U2994 (N_2994,N_2906,N_2915);
nand U2995 (N_2995,N_2903,N_2936);
or U2996 (N_2996,N_2920,N_2946);
nor U2997 (N_2997,N_2948,N_2924);
nand U2998 (N_2998,N_2926,N_2945);
nor U2999 (N_2999,N_2924,N_2932);
nor UO_0 (O_0,N_2997,N_2983);
nand UO_1 (O_1,N_2984,N_2976);
or UO_2 (O_2,N_2982,N_2966);
and UO_3 (O_3,N_2964,N_2952);
nand UO_4 (O_4,N_2977,N_2988);
or UO_5 (O_5,N_2980,N_2981);
nor UO_6 (O_6,N_2968,N_2978);
or UO_7 (O_7,N_2961,N_2958);
or UO_8 (O_8,N_2990,N_2950);
or UO_9 (O_9,N_2965,N_2986);
nor UO_10 (O_10,N_2955,N_2959);
nand UO_11 (O_11,N_2957,N_2960);
and UO_12 (O_12,N_2973,N_2994);
or UO_13 (O_13,N_2975,N_2956);
nor UO_14 (O_14,N_2972,N_2951);
or UO_15 (O_15,N_2987,N_2954);
and UO_16 (O_16,N_2970,N_2999);
and UO_17 (O_17,N_2971,N_2995);
and UO_18 (O_18,N_2985,N_2967);
nor UO_19 (O_19,N_2953,N_2963);
or UO_20 (O_20,N_2974,N_2992);
or UO_21 (O_21,N_2993,N_2996);
and UO_22 (O_22,N_2991,N_2998);
or UO_23 (O_23,N_2979,N_2962);
or UO_24 (O_24,N_2969,N_2989);
nand UO_25 (O_25,N_2964,N_2969);
or UO_26 (O_26,N_2962,N_2995);
or UO_27 (O_27,N_2960,N_2950);
nand UO_28 (O_28,N_2978,N_2958);
nor UO_29 (O_29,N_2975,N_2977);
nand UO_30 (O_30,N_2973,N_2966);
nor UO_31 (O_31,N_2957,N_2951);
or UO_32 (O_32,N_2975,N_2987);
or UO_33 (O_33,N_2966,N_2959);
nand UO_34 (O_34,N_2962,N_2971);
and UO_35 (O_35,N_2958,N_2951);
or UO_36 (O_36,N_2955,N_2963);
nor UO_37 (O_37,N_2979,N_2953);
or UO_38 (O_38,N_2961,N_2967);
nor UO_39 (O_39,N_2969,N_2992);
nor UO_40 (O_40,N_2969,N_2950);
and UO_41 (O_41,N_2961,N_2962);
nand UO_42 (O_42,N_2993,N_2978);
nor UO_43 (O_43,N_2977,N_2996);
and UO_44 (O_44,N_2952,N_2972);
nor UO_45 (O_45,N_2952,N_2999);
nand UO_46 (O_46,N_2952,N_2968);
xor UO_47 (O_47,N_2970,N_2990);
nor UO_48 (O_48,N_2961,N_2984);
xnor UO_49 (O_49,N_2957,N_2998);
and UO_50 (O_50,N_2994,N_2952);
and UO_51 (O_51,N_2964,N_2999);
and UO_52 (O_52,N_2964,N_2957);
nand UO_53 (O_53,N_2970,N_2982);
nand UO_54 (O_54,N_2961,N_2980);
nand UO_55 (O_55,N_2986,N_2999);
nand UO_56 (O_56,N_2969,N_2953);
and UO_57 (O_57,N_2967,N_2981);
nor UO_58 (O_58,N_2974,N_2991);
nand UO_59 (O_59,N_2995,N_2952);
nor UO_60 (O_60,N_2986,N_2969);
xor UO_61 (O_61,N_2969,N_2952);
nand UO_62 (O_62,N_2951,N_2999);
or UO_63 (O_63,N_2973,N_2991);
and UO_64 (O_64,N_2995,N_2979);
nand UO_65 (O_65,N_2971,N_2976);
nor UO_66 (O_66,N_2987,N_2957);
nand UO_67 (O_67,N_2955,N_2998);
and UO_68 (O_68,N_2959,N_2981);
and UO_69 (O_69,N_2982,N_2961);
or UO_70 (O_70,N_2990,N_2955);
nor UO_71 (O_71,N_2956,N_2957);
and UO_72 (O_72,N_2968,N_2990);
or UO_73 (O_73,N_2998,N_2988);
or UO_74 (O_74,N_2961,N_2987);
nand UO_75 (O_75,N_2955,N_2996);
nor UO_76 (O_76,N_2974,N_2989);
and UO_77 (O_77,N_2982,N_2985);
or UO_78 (O_78,N_2964,N_2989);
nand UO_79 (O_79,N_2967,N_2955);
or UO_80 (O_80,N_2994,N_2980);
and UO_81 (O_81,N_2999,N_2979);
or UO_82 (O_82,N_2995,N_2950);
and UO_83 (O_83,N_2954,N_2962);
and UO_84 (O_84,N_2988,N_2978);
nand UO_85 (O_85,N_2976,N_2952);
nor UO_86 (O_86,N_2961,N_2977);
xor UO_87 (O_87,N_2988,N_2966);
nor UO_88 (O_88,N_2996,N_2995);
nor UO_89 (O_89,N_2998,N_2995);
or UO_90 (O_90,N_2965,N_2968);
nor UO_91 (O_91,N_2980,N_2952);
nand UO_92 (O_92,N_2950,N_2967);
or UO_93 (O_93,N_2973,N_2974);
or UO_94 (O_94,N_2994,N_2955);
or UO_95 (O_95,N_2960,N_2983);
nor UO_96 (O_96,N_2958,N_2986);
or UO_97 (O_97,N_2988,N_2952);
and UO_98 (O_98,N_2957,N_2984);
nand UO_99 (O_99,N_2951,N_2950);
nand UO_100 (O_100,N_2997,N_2999);
nand UO_101 (O_101,N_2952,N_2996);
nor UO_102 (O_102,N_2964,N_2995);
nor UO_103 (O_103,N_2976,N_2963);
or UO_104 (O_104,N_2984,N_2953);
or UO_105 (O_105,N_2971,N_2968);
or UO_106 (O_106,N_2981,N_2979);
nor UO_107 (O_107,N_2975,N_2952);
nor UO_108 (O_108,N_2986,N_2978);
or UO_109 (O_109,N_2989,N_2979);
nand UO_110 (O_110,N_2988,N_2990);
nand UO_111 (O_111,N_2965,N_2974);
nor UO_112 (O_112,N_2951,N_2989);
nand UO_113 (O_113,N_2957,N_2997);
nand UO_114 (O_114,N_2977,N_2985);
or UO_115 (O_115,N_2976,N_2961);
or UO_116 (O_116,N_2962,N_2984);
or UO_117 (O_117,N_2980,N_2996);
xnor UO_118 (O_118,N_2978,N_2950);
and UO_119 (O_119,N_2967,N_2972);
and UO_120 (O_120,N_2994,N_2964);
nor UO_121 (O_121,N_2988,N_2957);
and UO_122 (O_122,N_2979,N_2963);
nand UO_123 (O_123,N_2983,N_2956);
and UO_124 (O_124,N_2958,N_2992);
or UO_125 (O_125,N_2958,N_2988);
nand UO_126 (O_126,N_2998,N_2960);
or UO_127 (O_127,N_2999,N_2987);
or UO_128 (O_128,N_2962,N_2981);
or UO_129 (O_129,N_2986,N_2988);
nand UO_130 (O_130,N_2979,N_2984);
nand UO_131 (O_131,N_2957,N_2986);
nand UO_132 (O_132,N_2973,N_2977);
and UO_133 (O_133,N_2999,N_2957);
or UO_134 (O_134,N_2995,N_2988);
nand UO_135 (O_135,N_2985,N_2992);
or UO_136 (O_136,N_2994,N_2954);
or UO_137 (O_137,N_2991,N_2961);
nor UO_138 (O_138,N_2960,N_2962);
nand UO_139 (O_139,N_2968,N_2959);
nand UO_140 (O_140,N_2980,N_2965);
or UO_141 (O_141,N_2958,N_2977);
and UO_142 (O_142,N_2987,N_2959);
nand UO_143 (O_143,N_2978,N_2992);
nand UO_144 (O_144,N_2984,N_2999);
or UO_145 (O_145,N_2998,N_2992);
nand UO_146 (O_146,N_2969,N_2985);
nand UO_147 (O_147,N_2950,N_2966);
nor UO_148 (O_148,N_2952,N_2962);
nor UO_149 (O_149,N_2994,N_2976);
nor UO_150 (O_150,N_2980,N_2993);
nor UO_151 (O_151,N_2952,N_2974);
nor UO_152 (O_152,N_2970,N_2992);
and UO_153 (O_153,N_2998,N_2974);
xnor UO_154 (O_154,N_2978,N_2990);
and UO_155 (O_155,N_2995,N_2951);
or UO_156 (O_156,N_2987,N_2970);
or UO_157 (O_157,N_2950,N_2987);
nand UO_158 (O_158,N_2952,N_2966);
nor UO_159 (O_159,N_2996,N_2954);
nor UO_160 (O_160,N_2983,N_2986);
or UO_161 (O_161,N_2966,N_2996);
nor UO_162 (O_162,N_2959,N_2986);
and UO_163 (O_163,N_2991,N_2958);
and UO_164 (O_164,N_2992,N_2983);
or UO_165 (O_165,N_2976,N_2974);
or UO_166 (O_166,N_2985,N_2956);
nand UO_167 (O_167,N_2996,N_2991);
and UO_168 (O_168,N_2977,N_2950);
or UO_169 (O_169,N_2994,N_2991);
nand UO_170 (O_170,N_2961,N_2975);
and UO_171 (O_171,N_2955,N_2962);
and UO_172 (O_172,N_2997,N_2976);
or UO_173 (O_173,N_2965,N_2959);
nand UO_174 (O_174,N_2954,N_2977);
xor UO_175 (O_175,N_2959,N_2971);
nor UO_176 (O_176,N_2956,N_2955);
nand UO_177 (O_177,N_2993,N_2971);
xor UO_178 (O_178,N_2995,N_2997);
nand UO_179 (O_179,N_2996,N_2982);
nand UO_180 (O_180,N_2992,N_2959);
or UO_181 (O_181,N_2990,N_2965);
nand UO_182 (O_182,N_2964,N_2974);
nand UO_183 (O_183,N_2983,N_2970);
xnor UO_184 (O_184,N_2997,N_2984);
nand UO_185 (O_185,N_2980,N_2989);
nor UO_186 (O_186,N_2998,N_2982);
or UO_187 (O_187,N_2960,N_2953);
nor UO_188 (O_188,N_2960,N_2972);
and UO_189 (O_189,N_2980,N_2969);
nor UO_190 (O_190,N_2983,N_2964);
and UO_191 (O_191,N_2966,N_2992);
and UO_192 (O_192,N_2954,N_2951);
or UO_193 (O_193,N_2950,N_2974);
nand UO_194 (O_194,N_2987,N_2996);
and UO_195 (O_195,N_2950,N_2968);
or UO_196 (O_196,N_2972,N_2976);
nor UO_197 (O_197,N_2951,N_2968);
nand UO_198 (O_198,N_2990,N_2951);
nand UO_199 (O_199,N_2999,N_2969);
or UO_200 (O_200,N_2980,N_2958);
or UO_201 (O_201,N_2961,N_2969);
and UO_202 (O_202,N_2961,N_2956);
or UO_203 (O_203,N_2967,N_2959);
xnor UO_204 (O_204,N_2978,N_2956);
nor UO_205 (O_205,N_2983,N_2987);
or UO_206 (O_206,N_2954,N_2960);
and UO_207 (O_207,N_2952,N_2951);
nor UO_208 (O_208,N_2978,N_2977);
nor UO_209 (O_209,N_2973,N_2987);
nor UO_210 (O_210,N_2953,N_2993);
nor UO_211 (O_211,N_2997,N_2962);
or UO_212 (O_212,N_2985,N_2958);
nor UO_213 (O_213,N_2981,N_2992);
and UO_214 (O_214,N_2955,N_2992);
nand UO_215 (O_215,N_2981,N_2964);
and UO_216 (O_216,N_2989,N_2971);
nand UO_217 (O_217,N_2978,N_2997);
or UO_218 (O_218,N_2961,N_2964);
nor UO_219 (O_219,N_2958,N_2996);
or UO_220 (O_220,N_2971,N_2961);
nand UO_221 (O_221,N_2986,N_2966);
and UO_222 (O_222,N_2968,N_2999);
and UO_223 (O_223,N_2965,N_2953);
nor UO_224 (O_224,N_2986,N_2984);
nor UO_225 (O_225,N_2993,N_2961);
or UO_226 (O_226,N_2963,N_2990);
nand UO_227 (O_227,N_2974,N_2995);
nor UO_228 (O_228,N_2969,N_2954);
nor UO_229 (O_229,N_2977,N_2952);
and UO_230 (O_230,N_2983,N_2999);
and UO_231 (O_231,N_2954,N_2975);
or UO_232 (O_232,N_2974,N_2968);
or UO_233 (O_233,N_2958,N_2968);
nand UO_234 (O_234,N_2975,N_2965);
nor UO_235 (O_235,N_2979,N_2985);
nor UO_236 (O_236,N_2974,N_2997);
or UO_237 (O_237,N_2992,N_2962);
and UO_238 (O_238,N_2955,N_2972);
or UO_239 (O_239,N_2981,N_2988);
nand UO_240 (O_240,N_2986,N_2973);
or UO_241 (O_241,N_2980,N_2983);
nand UO_242 (O_242,N_2987,N_2960);
nor UO_243 (O_243,N_2960,N_2980);
or UO_244 (O_244,N_2979,N_2977);
nor UO_245 (O_245,N_2976,N_2999);
and UO_246 (O_246,N_2994,N_2959);
nor UO_247 (O_247,N_2955,N_2966);
and UO_248 (O_248,N_2983,N_2965);
nand UO_249 (O_249,N_2984,N_2955);
or UO_250 (O_250,N_2956,N_2976);
and UO_251 (O_251,N_2976,N_2959);
nor UO_252 (O_252,N_2990,N_2962);
nand UO_253 (O_253,N_2992,N_2999);
and UO_254 (O_254,N_2991,N_2951);
nor UO_255 (O_255,N_2998,N_2959);
nand UO_256 (O_256,N_2954,N_2999);
or UO_257 (O_257,N_2959,N_2984);
or UO_258 (O_258,N_2963,N_2958);
or UO_259 (O_259,N_2954,N_2973);
nor UO_260 (O_260,N_2958,N_2953);
nand UO_261 (O_261,N_2969,N_2979);
nand UO_262 (O_262,N_2971,N_2965);
or UO_263 (O_263,N_2993,N_2975);
or UO_264 (O_264,N_2977,N_2970);
or UO_265 (O_265,N_2976,N_2973);
and UO_266 (O_266,N_2971,N_2967);
or UO_267 (O_267,N_2953,N_2972);
nor UO_268 (O_268,N_2999,N_2991);
nor UO_269 (O_269,N_2981,N_2974);
nand UO_270 (O_270,N_2978,N_2994);
nor UO_271 (O_271,N_2997,N_2952);
nor UO_272 (O_272,N_2959,N_2970);
nand UO_273 (O_273,N_2951,N_2994);
nand UO_274 (O_274,N_2984,N_2964);
or UO_275 (O_275,N_2967,N_2952);
or UO_276 (O_276,N_2972,N_2983);
nor UO_277 (O_277,N_2987,N_2958);
and UO_278 (O_278,N_2974,N_2999);
nor UO_279 (O_279,N_2995,N_2985);
nand UO_280 (O_280,N_2955,N_2976);
or UO_281 (O_281,N_2986,N_2981);
nor UO_282 (O_282,N_2994,N_2990);
nor UO_283 (O_283,N_2956,N_2973);
nor UO_284 (O_284,N_2984,N_2968);
nor UO_285 (O_285,N_2967,N_2997);
or UO_286 (O_286,N_2977,N_2968);
and UO_287 (O_287,N_2950,N_2993);
nor UO_288 (O_288,N_2980,N_2976);
or UO_289 (O_289,N_2976,N_2967);
or UO_290 (O_290,N_2969,N_2972);
or UO_291 (O_291,N_2975,N_2973);
nand UO_292 (O_292,N_2969,N_2987);
nor UO_293 (O_293,N_2963,N_2982);
nand UO_294 (O_294,N_2968,N_2991);
or UO_295 (O_295,N_2963,N_2981);
nor UO_296 (O_296,N_2961,N_2953);
nand UO_297 (O_297,N_2992,N_2979);
nand UO_298 (O_298,N_2963,N_2971);
and UO_299 (O_299,N_2954,N_2957);
and UO_300 (O_300,N_2956,N_2979);
nor UO_301 (O_301,N_2994,N_2975);
nand UO_302 (O_302,N_2974,N_2993);
or UO_303 (O_303,N_2985,N_2960);
nor UO_304 (O_304,N_2987,N_2974);
nor UO_305 (O_305,N_2955,N_2985);
and UO_306 (O_306,N_2971,N_2973);
nand UO_307 (O_307,N_2957,N_2961);
and UO_308 (O_308,N_2967,N_2966);
nand UO_309 (O_309,N_2974,N_2979);
or UO_310 (O_310,N_2957,N_2975);
nor UO_311 (O_311,N_2958,N_2954);
nand UO_312 (O_312,N_2960,N_2959);
nor UO_313 (O_313,N_2994,N_2979);
nor UO_314 (O_314,N_2974,N_2958);
and UO_315 (O_315,N_2979,N_2996);
or UO_316 (O_316,N_2972,N_2958);
nor UO_317 (O_317,N_2982,N_2957);
and UO_318 (O_318,N_2956,N_2992);
and UO_319 (O_319,N_2997,N_2969);
and UO_320 (O_320,N_2983,N_2967);
and UO_321 (O_321,N_2998,N_2979);
nand UO_322 (O_322,N_2984,N_2973);
or UO_323 (O_323,N_2962,N_2998);
or UO_324 (O_324,N_2974,N_2961);
and UO_325 (O_325,N_2962,N_2950);
nand UO_326 (O_326,N_2998,N_2994);
or UO_327 (O_327,N_2985,N_2989);
or UO_328 (O_328,N_2974,N_2977);
nor UO_329 (O_329,N_2960,N_2994);
nor UO_330 (O_330,N_2952,N_2989);
and UO_331 (O_331,N_2966,N_2953);
nor UO_332 (O_332,N_2994,N_2961);
or UO_333 (O_333,N_2990,N_2958);
nor UO_334 (O_334,N_2990,N_2982);
and UO_335 (O_335,N_2961,N_2986);
and UO_336 (O_336,N_2953,N_2970);
or UO_337 (O_337,N_2966,N_2984);
nor UO_338 (O_338,N_2967,N_2988);
and UO_339 (O_339,N_2990,N_2961);
or UO_340 (O_340,N_2985,N_2999);
nand UO_341 (O_341,N_2962,N_2956);
nand UO_342 (O_342,N_2988,N_2989);
nor UO_343 (O_343,N_2953,N_2962);
and UO_344 (O_344,N_2973,N_2996);
nand UO_345 (O_345,N_2979,N_2978);
and UO_346 (O_346,N_2965,N_2962);
nand UO_347 (O_347,N_2997,N_2990);
xnor UO_348 (O_348,N_2984,N_2983);
nand UO_349 (O_349,N_2977,N_2953);
or UO_350 (O_350,N_2968,N_2980);
and UO_351 (O_351,N_2960,N_2966);
nand UO_352 (O_352,N_2981,N_2990);
nand UO_353 (O_353,N_2956,N_2995);
or UO_354 (O_354,N_2987,N_2992);
nor UO_355 (O_355,N_2977,N_2993);
or UO_356 (O_356,N_2982,N_2987);
or UO_357 (O_357,N_2953,N_2976);
and UO_358 (O_358,N_2967,N_2982);
nand UO_359 (O_359,N_2972,N_2995);
nor UO_360 (O_360,N_2997,N_2981);
nand UO_361 (O_361,N_2986,N_2967);
or UO_362 (O_362,N_2963,N_2969);
nor UO_363 (O_363,N_2983,N_2996);
or UO_364 (O_364,N_2977,N_2994);
nor UO_365 (O_365,N_2951,N_2983);
nor UO_366 (O_366,N_2963,N_2960);
and UO_367 (O_367,N_2997,N_2963);
or UO_368 (O_368,N_2954,N_2981);
nor UO_369 (O_369,N_2988,N_2976);
or UO_370 (O_370,N_2963,N_2966);
xnor UO_371 (O_371,N_2983,N_2989);
nand UO_372 (O_372,N_2994,N_2989);
nand UO_373 (O_373,N_2970,N_2971);
and UO_374 (O_374,N_2991,N_2971);
or UO_375 (O_375,N_2955,N_2986);
nand UO_376 (O_376,N_2997,N_2996);
and UO_377 (O_377,N_2996,N_2965);
and UO_378 (O_378,N_2984,N_2995);
or UO_379 (O_379,N_2995,N_2993);
or UO_380 (O_380,N_2988,N_2999);
nand UO_381 (O_381,N_2984,N_2980);
xnor UO_382 (O_382,N_2976,N_2992);
nor UO_383 (O_383,N_2956,N_2963);
nand UO_384 (O_384,N_2962,N_2999);
nor UO_385 (O_385,N_2982,N_2997);
or UO_386 (O_386,N_2983,N_2981);
nand UO_387 (O_387,N_2971,N_2952);
nand UO_388 (O_388,N_2969,N_2984);
xor UO_389 (O_389,N_2956,N_2966);
and UO_390 (O_390,N_2999,N_2955);
nor UO_391 (O_391,N_2951,N_2975);
nor UO_392 (O_392,N_2955,N_2973);
or UO_393 (O_393,N_2960,N_2990);
nor UO_394 (O_394,N_2962,N_2968);
or UO_395 (O_395,N_2981,N_2977);
and UO_396 (O_396,N_2956,N_2981);
and UO_397 (O_397,N_2993,N_2970);
nand UO_398 (O_398,N_2961,N_2965);
nor UO_399 (O_399,N_2978,N_2991);
nand UO_400 (O_400,N_2992,N_2960);
or UO_401 (O_401,N_2967,N_2956);
and UO_402 (O_402,N_2972,N_2971);
and UO_403 (O_403,N_2976,N_2989);
or UO_404 (O_404,N_2969,N_2990);
nor UO_405 (O_405,N_2987,N_2963);
nor UO_406 (O_406,N_2981,N_2968);
nor UO_407 (O_407,N_2961,N_2966);
and UO_408 (O_408,N_2992,N_2967);
and UO_409 (O_409,N_2954,N_2971);
or UO_410 (O_410,N_2972,N_2989);
and UO_411 (O_411,N_2979,N_2966);
nor UO_412 (O_412,N_2980,N_2954);
nand UO_413 (O_413,N_2995,N_2981);
or UO_414 (O_414,N_2976,N_2962);
or UO_415 (O_415,N_2997,N_2998);
nand UO_416 (O_416,N_2964,N_2962);
nand UO_417 (O_417,N_2950,N_2983);
nor UO_418 (O_418,N_2956,N_2971);
and UO_419 (O_419,N_2950,N_2964);
nor UO_420 (O_420,N_2956,N_2986);
nor UO_421 (O_421,N_2984,N_2994);
nor UO_422 (O_422,N_2992,N_2991);
or UO_423 (O_423,N_2955,N_2971);
and UO_424 (O_424,N_2968,N_2979);
or UO_425 (O_425,N_2985,N_2990);
and UO_426 (O_426,N_2952,N_2959);
nor UO_427 (O_427,N_2986,N_2968);
nor UO_428 (O_428,N_2983,N_2990);
or UO_429 (O_429,N_2956,N_2959);
nor UO_430 (O_430,N_2967,N_2973);
or UO_431 (O_431,N_2962,N_2966);
and UO_432 (O_432,N_2955,N_2995);
or UO_433 (O_433,N_2975,N_2998);
xor UO_434 (O_434,N_2986,N_2953);
nor UO_435 (O_435,N_2951,N_2973);
nand UO_436 (O_436,N_2967,N_2958);
nor UO_437 (O_437,N_2953,N_2955);
nor UO_438 (O_438,N_2978,N_2953);
or UO_439 (O_439,N_2970,N_2973);
and UO_440 (O_440,N_2960,N_2979);
xnor UO_441 (O_441,N_2970,N_2967);
nor UO_442 (O_442,N_2986,N_2996);
nand UO_443 (O_443,N_2992,N_2973);
or UO_444 (O_444,N_2966,N_2954);
or UO_445 (O_445,N_2998,N_2980);
nand UO_446 (O_446,N_2981,N_2953);
nor UO_447 (O_447,N_2974,N_2967);
and UO_448 (O_448,N_2950,N_2997);
and UO_449 (O_449,N_2953,N_2967);
nor UO_450 (O_450,N_2959,N_2983);
nor UO_451 (O_451,N_2951,N_2982);
or UO_452 (O_452,N_2986,N_2951);
or UO_453 (O_453,N_2974,N_2982);
nand UO_454 (O_454,N_2966,N_2970);
and UO_455 (O_455,N_2974,N_2994);
or UO_456 (O_456,N_2962,N_2951);
nand UO_457 (O_457,N_2999,N_2973);
xnor UO_458 (O_458,N_2970,N_2954);
and UO_459 (O_459,N_2993,N_2986);
nor UO_460 (O_460,N_2966,N_2994);
or UO_461 (O_461,N_2992,N_2968);
or UO_462 (O_462,N_2954,N_2965);
xor UO_463 (O_463,N_2962,N_2985);
or UO_464 (O_464,N_2990,N_2967);
nand UO_465 (O_465,N_2968,N_2954);
nor UO_466 (O_466,N_2990,N_2971);
nand UO_467 (O_467,N_2962,N_2963);
nand UO_468 (O_468,N_2950,N_2976);
or UO_469 (O_469,N_2955,N_2989);
nor UO_470 (O_470,N_2975,N_2984);
and UO_471 (O_471,N_2973,N_2989);
nor UO_472 (O_472,N_2964,N_2998);
or UO_473 (O_473,N_2953,N_2996);
nor UO_474 (O_474,N_2989,N_2960);
xnor UO_475 (O_475,N_2955,N_2975);
or UO_476 (O_476,N_2955,N_2997);
nor UO_477 (O_477,N_2963,N_2954);
nor UO_478 (O_478,N_2950,N_2952);
nand UO_479 (O_479,N_2968,N_2972);
nand UO_480 (O_480,N_2985,N_2981);
nand UO_481 (O_481,N_2997,N_2954);
and UO_482 (O_482,N_2982,N_2986);
nor UO_483 (O_483,N_2983,N_2993);
or UO_484 (O_484,N_2967,N_2962);
xnor UO_485 (O_485,N_2965,N_2998);
or UO_486 (O_486,N_2971,N_2983);
or UO_487 (O_487,N_2964,N_2967);
or UO_488 (O_488,N_2977,N_2986);
or UO_489 (O_489,N_2978,N_2980);
or UO_490 (O_490,N_2959,N_2979);
nor UO_491 (O_491,N_2972,N_2986);
or UO_492 (O_492,N_2955,N_2978);
or UO_493 (O_493,N_2958,N_2982);
or UO_494 (O_494,N_2970,N_2965);
nor UO_495 (O_495,N_2986,N_2992);
and UO_496 (O_496,N_2953,N_2974);
nor UO_497 (O_497,N_2958,N_2966);
and UO_498 (O_498,N_2988,N_2987);
or UO_499 (O_499,N_2995,N_2976);
endmodule