module basic_2500_25000_3000_8_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xnor U0 (N_0,In_143,In_423);
nand U1 (N_1,In_1430,In_1552);
and U2 (N_2,In_503,In_1568);
xor U3 (N_3,In_1629,In_1170);
nand U4 (N_4,In_1519,In_1817);
nor U5 (N_5,In_2128,In_615);
xnor U6 (N_6,In_657,In_1117);
xor U7 (N_7,In_1990,In_1722);
or U8 (N_8,In_231,In_1657);
xor U9 (N_9,In_1197,In_2148);
and U10 (N_10,In_263,In_1672);
xor U11 (N_11,In_2199,In_1499);
nor U12 (N_12,In_377,In_149);
or U13 (N_13,In_975,In_81);
nand U14 (N_14,In_361,In_485);
or U15 (N_15,In_1836,In_892);
nor U16 (N_16,In_1780,In_1653);
nor U17 (N_17,In_136,In_2481);
xor U18 (N_18,In_103,In_1193);
nand U19 (N_19,In_1700,In_1320);
xor U20 (N_20,In_148,In_1547);
xnor U21 (N_21,In_137,In_2390);
nand U22 (N_22,In_1309,In_2291);
xnor U23 (N_23,In_445,In_294);
nor U24 (N_24,In_1831,In_1219);
xor U25 (N_25,In_935,In_532);
and U26 (N_26,In_991,In_2020);
xnor U27 (N_27,In_1719,In_2005);
or U28 (N_28,In_2018,In_1962);
and U29 (N_29,In_934,In_446);
xnor U30 (N_30,In_2321,In_1821);
or U31 (N_31,In_1195,In_1559);
and U32 (N_32,In_1806,In_1603);
nand U33 (N_33,In_967,In_620);
and U34 (N_34,In_1776,In_781);
nand U35 (N_35,In_641,In_1937);
xnor U36 (N_36,In_1460,In_1261);
xnor U37 (N_37,In_1484,In_741);
xor U38 (N_38,In_2276,In_1079);
and U39 (N_39,In_910,In_875);
nand U40 (N_40,In_1730,In_379);
and U41 (N_41,In_1680,In_834);
and U42 (N_42,In_1216,In_1540);
and U43 (N_43,In_1929,In_307);
nor U44 (N_44,In_1704,In_1804);
nand U45 (N_45,In_683,In_971);
nand U46 (N_46,In_9,In_678);
and U47 (N_47,In_2361,In_1156);
nand U48 (N_48,In_2225,In_708);
xnor U49 (N_49,In_1126,In_255);
nor U50 (N_50,In_1186,In_576);
and U51 (N_51,In_1982,In_2324);
nor U52 (N_52,In_1556,In_2077);
and U53 (N_53,In_1297,In_504);
or U54 (N_54,In_780,In_2298);
or U55 (N_55,In_1744,In_1808);
xor U56 (N_56,In_2111,In_646);
nand U57 (N_57,In_367,In_1585);
xor U58 (N_58,In_162,In_2477);
nand U59 (N_59,In_1416,In_365);
nand U60 (N_60,In_61,In_2252);
nand U61 (N_61,In_755,In_2454);
nor U62 (N_62,In_1714,In_244);
xnor U63 (N_63,In_105,In_1157);
xor U64 (N_64,In_2320,In_617);
or U65 (N_65,In_2293,In_1686);
and U66 (N_66,In_2170,In_2141);
nor U67 (N_67,In_196,In_976);
and U68 (N_68,In_1949,In_596);
and U69 (N_69,In_1249,In_2081);
nand U70 (N_70,In_14,In_1662);
nor U71 (N_71,In_89,In_1671);
nor U72 (N_72,In_359,In_57);
xnor U73 (N_73,In_2061,In_2122);
nor U74 (N_74,In_321,In_1236);
or U75 (N_75,In_1,In_547);
nor U76 (N_76,In_2339,In_820);
xor U77 (N_77,In_1267,In_2112);
or U78 (N_78,In_2400,In_1592);
and U79 (N_79,In_2236,In_267);
or U80 (N_80,In_1119,In_749);
and U81 (N_81,In_878,In_1208);
xor U82 (N_82,In_1718,In_2188);
or U83 (N_83,In_165,In_1385);
or U84 (N_84,In_594,In_744);
nor U85 (N_85,In_145,In_1816);
and U86 (N_86,In_2427,In_1943);
nand U87 (N_87,In_872,In_1908);
xor U88 (N_88,In_1270,In_918);
nand U89 (N_89,In_1505,In_2340);
or U90 (N_90,In_658,In_2137);
nor U91 (N_91,In_649,In_2315);
and U92 (N_92,In_1665,In_1899);
and U93 (N_93,In_2443,In_1263);
xnor U94 (N_94,In_1098,In_2489);
or U95 (N_95,In_2003,In_17);
or U96 (N_96,In_524,In_1069);
nor U97 (N_97,In_1569,In_860);
xnor U98 (N_98,In_184,In_1842);
or U99 (N_99,In_1866,In_1476);
and U100 (N_100,In_1551,In_2255);
xor U101 (N_101,In_603,In_1077);
nand U102 (N_102,In_2186,In_2416);
xnor U103 (N_103,In_463,In_1223);
nand U104 (N_104,In_982,In_2384);
and U105 (N_105,In_358,In_1693);
or U106 (N_106,In_1595,In_684);
nor U107 (N_107,In_2375,In_1545);
and U108 (N_108,In_2224,In_1873);
xor U109 (N_109,In_917,In_602);
nor U110 (N_110,In_2373,In_1642);
or U111 (N_111,In_916,In_364);
nand U112 (N_112,In_554,In_447);
xor U113 (N_113,In_945,In_628);
nand U114 (N_114,In_1398,In_422);
and U115 (N_115,In_1896,In_1209);
xor U116 (N_116,In_2311,In_530);
nand U117 (N_117,In_1196,In_775);
and U118 (N_118,In_2129,In_2486);
and U119 (N_119,In_1262,In_1736);
nand U120 (N_120,In_369,In_1353);
nor U121 (N_121,In_200,In_2073);
nand U122 (N_122,In_689,In_1549);
or U123 (N_123,In_599,In_1888);
xnor U124 (N_124,In_1652,In_2260);
nand U125 (N_125,In_770,In_1845);
or U126 (N_126,In_2035,In_1521);
or U127 (N_127,In_1691,In_1107);
nand U128 (N_128,In_455,In_568);
nand U129 (N_129,In_521,In_42);
nand U130 (N_130,In_2187,In_2422);
or U131 (N_131,In_1684,In_2409);
nand U132 (N_132,In_331,In_693);
nor U133 (N_133,In_2149,In_798);
and U134 (N_134,In_2366,In_341);
nand U135 (N_135,In_1913,In_1354);
nor U136 (N_136,In_1052,In_2071);
and U137 (N_137,In_577,In_686);
nor U138 (N_138,In_2180,In_527);
nand U139 (N_139,In_1682,In_1846);
xor U140 (N_140,In_597,In_91);
nand U141 (N_141,In_2353,In_2494);
nand U142 (N_142,In_2197,In_1281);
nor U143 (N_143,In_2323,In_1100);
or U144 (N_144,In_1960,In_941);
xnor U145 (N_145,In_919,In_1633);
or U146 (N_146,In_2286,In_1989);
xor U147 (N_147,In_816,In_866);
nand U148 (N_148,In_1645,In_1073);
and U149 (N_149,In_519,In_893);
and U150 (N_150,In_213,In_1063);
and U151 (N_151,In_1362,In_2418);
and U152 (N_152,In_1455,In_1120);
xor U153 (N_153,In_484,In_1970);
nand U154 (N_154,In_1053,In_1474);
and U155 (N_155,In_2131,In_1066);
nor U156 (N_156,In_903,In_106);
xor U157 (N_157,In_64,In_2036);
nor U158 (N_158,In_842,In_1756);
xnor U159 (N_159,In_2176,In_1159);
and U160 (N_160,In_178,In_2302);
nand U161 (N_161,In_656,In_430);
xnor U162 (N_162,In_167,In_1106);
and U163 (N_163,In_397,In_762);
or U164 (N_164,In_2010,In_1811);
or U165 (N_165,In_2108,In_2239);
xor U166 (N_166,In_465,In_930);
nand U167 (N_167,In_1864,In_1016);
or U168 (N_168,In_2478,In_2341);
nand U169 (N_169,In_632,In_690);
or U170 (N_170,In_404,In_1560);
nand U171 (N_171,In_1390,In_352);
and U172 (N_172,In_2307,In_41);
nand U173 (N_173,In_2369,In_205);
nor U174 (N_174,In_822,In_135);
nand U175 (N_175,In_700,In_1952);
xor U176 (N_176,In_295,In_825);
nor U177 (N_177,In_1346,In_1173);
nand U178 (N_178,In_2192,In_957);
nor U179 (N_179,In_1885,In_697);
or U180 (N_180,In_2380,In_998);
nand U181 (N_181,In_1041,In_963);
nand U182 (N_182,In_300,In_996);
or U183 (N_183,In_1468,In_1858);
nand U184 (N_184,In_1648,In_886);
or U185 (N_185,In_507,In_898);
xor U186 (N_186,In_407,In_243);
and U187 (N_187,In_55,In_2483);
nor U188 (N_188,In_160,In_1646);
and U189 (N_189,In_1213,In_371);
and U190 (N_190,In_2113,In_1244);
nand U191 (N_191,In_1045,In_652);
xnor U192 (N_192,In_2475,In_1469);
xor U193 (N_193,In_1456,In_1789);
nor U194 (N_194,In_1465,In_662);
xnor U195 (N_195,In_20,In_1395);
or U196 (N_196,In_1210,In_328);
and U197 (N_197,In_1161,In_2110);
or U198 (N_198,In_2265,In_141);
and U199 (N_199,In_1902,In_843);
or U200 (N_200,In_174,In_647);
or U201 (N_201,In_1003,In_1214);
nand U202 (N_202,In_1936,In_1481);
and U203 (N_203,In_355,In_211);
and U204 (N_204,In_966,In_444);
and U205 (N_205,In_175,In_537);
nor U206 (N_206,In_2208,In_1500);
nor U207 (N_207,In_283,In_2305);
xnor U208 (N_208,In_1054,In_1876);
or U209 (N_209,In_1333,In_1670);
xor U210 (N_210,In_1594,In_409);
or U211 (N_211,In_1344,In_1278);
or U212 (N_212,In_1717,In_2026);
and U213 (N_213,In_1994,In_1993);
and U214 (N_214,In_1294,In_1254);
xnor U215 (N_215,In_185,In_310);
xor U216 (N_216,In_515,In_1538);
nor U217 (N_217,In_2356,In_606);
or U218 (N_218,In_1185,In_1938);
nor U219 (N_219,In_461,In_1525);
nand U220 (N_220,In_219,In_865);
xor U221 (N_221,In_2251,In_1364);
nand U222 (N_222,In_1823,In_2498);
xnor U223 (N_223,In_2370,In_436);
xnor U224 (N_224,In_150,In_1631);
and U225 (N_225,In_675,In_329);
nor U226 (N_226,In_2468,In_2145);
nand U227 (N_227,In_1421,In_1351);
nand U228 (N_228,In_78,In_1382);
and U229 (N_229,In_2266,In_1412);
and U230 (N_230,In_1392,In_2459);
and U231 (N_231,In_676,In_1737);
nand U232 (N_232,In_40,In_1690);
or U233 (N_233,In_1799,In_188);
nand U234 (N_234,In_2457,In_152);
nand U235 (N_235,In_1371,In_304);
nor U236 (N_236,In_588,In_2028);
nor U237 (N_237,In_2271,In_508);
xor U238 (N_238,In_1786,In_1009);
nand U239 (N_239,In_1508,In_1134);
or U240 (N_240,In_863,In_1383);
or U241 (N_241,In_1955,In_1643);
or U242 (N_242,In_642,In_1591);
nor U243 (N_243,In_1080,In_385);
nor U244 (N_244,In_2157,In_774);
nor U245 (N_245,In_2415,In_748);
nand U246 (N_246,In_129,In_1380);
or U247 (N_247,In_490,In_132);
or U248 (N_248,In_425,In_817);
and U249 (N_249,In_2177,In_284);
and U250 (N_250,In_846,In_1703);
and U251 (N_251,In_2181,In_1621);
and U252 (N_252,In_2058,In_2243);
or U253 (N_253,In_1164,In_1321);
nor U254 (N_254,In_1869,In_1745);
and U255 (N_255,In_1124,In_71);
nand U256 (N_256,In_1683,In_601);
and U257 (N_257,In_654,In_961);
xor U258 (N_258,In_1036,In_1588);
nor U259 (N_259,In_292,In_1599);
and U260 (N_260,In_1055,In_555);
and U261 (N_261,In_1659,In_1956);
xor U262 (N_262,In_1423,In_1890);
xor U263 (N_263,In_1749,In_1400);
and U264 (N_264,In_619,In_94);
or U265 (N_265,In_1087,In_349);
or U266 (N_266,In_711,In_831);
nand U267 (N_267,In_1613,In_122);
and U268 (N_268,In_1977,In_516);
and U269 (N_269,In_506,In_552);
or U270 (N_270,In_1367,In_1942);
xor U271 (N_271,In_1660,In_877);
and U272 (N_272,In_1168,In_2484);
or U273 (N_273,In_2487,In_2219);
nor U274 (N_274,In_27,In_1813);
or U275 (N_275,In_173,In_1338);
nor U276 (N_276,In_2413,In_66);
or U277 (N_277,In_1248,In_1975);
nor U278 (N_278,In_1513,In_2039);
nor U279 (N_279,In_1991,In_192);
or U280 (N_280,In_698,In_109);
xor U281 (N_281,In_626,In_1179);
nor U282 (N_282,In_335,In_1972);
nor U283 (N_283,In_906,In_2055);
nand U284 (N_284,In_142,In_37);
nand U285 (N_285,In_1735,In_881);
xnor U286 (N_286,In_1397,In_1494);
or U287 (N_287,In_1034,In_1868);
nor U288 (N_288,In_1352,In_1910);
nor U289 (N_289,In_853,In_2300);
or U290 (N_290,In_1905,In_2372);
xnor U291 (N_291,In_2068,In_1721);
nand U292 (N_292,In_2139,In_1002);
nor U293 (N_293,In_311,In_301);
nand U294 (N_294,In_25,In_50);
nor U295 (N_295,In_351,In_1753);
xor U296 (N_296,In_911,In_121);
xor U297 (N_297,In_1688,In_2059);
or U298 (N_298,In_1007,In_753);
and U299 (N_299,In_2294,In_2069);
nor U300 (N_300,In_207,In_2451);
and U301 (N_301,In_1641,In_1291);
nand U302 (N_302,In_685,In_977);
xnor U303 (N_303,In_1184,In_2253);
and U304 (N_304,In_882,In_2403);
xor U305 (N_305,In_2306,In_553);
and U306 (N_306,In_931,In_2445);
nand U307 (N_307,In_758,In_1129);
or U308 (N_308,In_2283,In_824);
nand U309 (N_309,In_456,In_2104);
or U310 (N_310,In_1096,In_2496);
nor U311 (N_311,In_69,In_8);
xnor U312 (N_312,In_2250,In_633);
and U313 (N_313,In_1325,In_1163);
or U314 (N_314,In_2327,In_2075);
xnor U315 (N_315,In_193,In_2309);
nor U316 (N_316,In_856,In_1764);
nand U317 (N_317,In_564,In_574);
or U318 (N_318,In_2034,In_709);
xor U319 (N_319,In_838,In_1527);
or U320 (N_320,In_155,In_2354);
and U321 (N_321,In_724,In_226);
nor U322 (N_322,In_1105,In_1862);
nor U323 (N_323,In_833,In_90);
nand U324 (N_324,In_728,In_453);
and U325 (N_325,In_1853,In_980);
xor U326 (N_326,In_5,In_320);
and U327 (N_327,In_1271,In_2203);
or U328 (N_328,In_117,In_2301);
nand U329 (N_329,In_1410,In_1289);
and U330 (N_330,In_542,In_1356);
and U331 (N_331,In_1807,In_1878);
nand U332 (N_332,In_1085,In_1812);
or U333 (N_333,In_73,In_1727);
nor U334 (N_334,In_2452,In_591);
nand U335 (N_335,In_1998,In_3);
nor U336 (N_336,In_478,In_67);
and U337 (N_337,In_1006,In_2395);
or U338 (N_338,In_1716,In_829);
or U339 (N_339,In_2226,In_1061);
xnor U340 (N_340,In_128,In_803);
nor U341 (N_341,In_1795,In_417);
or U342 (N_342,In_373,In_1487);
or U343 (N_343,In_2347,In_2116);
xnor U344 (N_344,In_1576,In_458);
nor U345 (N_345,In_2493,In_1572);
xnor U346 (N_346,In_2241,In_688);
nor U347 (N_347,In_565,In_1414);
and U348 (N_348,In_1429,In_1761);
and U349 (N_349,In_273,In_1194);
or U350 (N_350,In_1121,In_170);
xor U351 (N_351,In_2420,In_1983);
xnor U352 (N_352,In_260,In_1495);
xnor U353 (N_353,In_2019,In_545);
and U354 (N_354,In_290,In_1212);
nor U355 (N_355,In_2365,In_1507);
nor U356 (N_356,In_2138,In_2212);
nor U357 (N_357,In_2355,In_479);
nand U358 (N_358,In_1181,In_375);
nor U359 (N_359,In_237,In_2231);
xor U360 (N_360,In_238,In_274);
xnor U361 (N_361,In_2499,In_1402);
xor U362 (N_362,In_1292,In_1814);
and U363 (N_363,In_1930,In_1190);
nor U364 (N_364,In_1781,In_868);
or U365 (N_365,In_759,In_443);
nor U366 (N_366,In_637,In_1710);
nor U367 (N_367,In_1927,In_1755);
nor U368 (N_368,In_1706,In_2450);
nor U369 (N_369,In_792,In_901);
xnor U370 (N_370,In_1768,In_765);
nand U371 (N_371,In_922,In_1516);
or U372 (N_372,In_1228,In_248);
xnor U373 (N_373,In_433,In_393);
and U374 (N_374,In_10,In_948);
xor U375 (N_375,In_1895,In_1112);
or U376 (N_376,In_627,In_544);
and U377 (N_377,In_836,In_2277);
or U378 (N_378,In_1200,In_1115);
or U379 (N_379,In_1733,In_1747);
nand U380 (N_380,In_2325,In_392);
or U381 (N_381,In_1010,In_1189);
xor U382 (N_382,In_1987,In_1004);
nor U383 (N_383,In_2491,In_421);
xnor U384 (N_384,In_538,In_464);
or U385 (N_385,In_2134,In_1295);
or U386 (N_386,In_1488,In_650);
nor U387 (N_387,In_1360,In_2049);
and U388 (N_388,In_854,In_403);
nand U389 (N_389,In_206,In_2169);
or U390 (N_390,In_2168,In_288);
or U391 (N_391,In_1461,In_1825);
nand U392 (N_392,In_795,In_487);
nor U393 (N_393,In_2013,In_929);
nand U394 (N_394,In_197,In_794);
and U395 (N_395,In_1122,In_592);
and U396 (N_396,In_1422,In_1206);
xor U397 (N_397,In_1024,In_1413);
nand U398 (N_398,In_984,In_1779);
xnor U399 (N_399,In_286,In_883);
and U400 (N_400,In_1305,In_1600);
or U401 (N_401,In_93,In_1339);
nor U402 (N_402,In_1211,In_2067);
and U403 (N_403,In_1793,In_1841);
nand U404 (N_404,In_2407,In_983);
nor U405 (N_405,In_120,In_735);
nand U406 (N_406,In_876,In_925);
or U407 (N_407,In_1075,In_1537);
and U408 (N_408,In_1875,In_2431);
nor U409 (N_409,In_2453,In_1785);
nor U410 (N_410,In_442,In_2247);
xor U411 (N_411,In_413,In_2017);
and U412 (N_412,In_703,In_1911);
nor U413 (N_413,In_374,In_1791);
and U414 (N_414,In_449,In_1449);
nor U415 (N_415,In_52,In_1113);
xnor U416 (N_416,In_1090,In_182);
xnor U417 (N_417,In_191,In_102);
and U418 (N_418,In_810,In_2414);
and U419 (N_419,In_2002,In_43);
or U420 (N_420,In_1501,In_2357);
nand U421 (N_421,In_1019,In_2346);
xnor U422 (N_422,In_573,In_344);
and U423 (N_423,In_899,In_880);
xor U424 (N_424,In_805,In_635);
nor U425 (N_425,In_1300,In_651);
xor U426 (N_426,In_2095,In_823);
and U427 (N_427,In_797,In_1635);
nand U428 (N_428,In_1777,In_1137);
nor U429 (N_429,In_2497,In_2093);
or U430 (N_430,In_2490,In_895);
or U431 (N_431,In_1227,In_1546);
or U432 (N_432,In_879,In_604);
nor U433 (N_433,In_1614,In_1059);
nor U434 (N_434,In_1451,In_1229);
nand U435 (N_435,In_282,In_75);
or U436 (N_436,In_802,In_1459);
and U437 (N_437,In_1965,In_1247);
nor U438 (N_438,In_220,In_281);
xor U439 (N_439,In_240,In_2065);
or U440 (N_440,In_1114,In_97);
nand U441 (N_441,In_2485,In_2245);
nor U442 (N_442,In_1405,In_496);
xor U443 (N_443,In_955,In_887);
nand U444 (N_444,In_1550,In_1959);
or U445 (N_445,In_270,In_114);
or U446 (N_446,In_2359,In_681);
nand U447 (N_447,In_1389,In_1969);
or U448 (N_448,In_687,In_242);
and U449 (N_449,In_972,In_1441);
xor U450 (N_450,In_873,In_319);
nor U451 (N_451,In_1857,In_677);
xnor U452 (N_452,In_1180,In_1694);
nor U453 (N_453,In_1750,In_2173);
nand U454 (N_454,In_1759,In_2006);
nand U455 (N_455,In_2406,In_1057);
xor U456 (N_456,In_956,In_1832);
nand U457 (N_457,In_1819,In_707);
xor U458 (N_458,In_2393,In_2047);
nor U459 (N_459,In_1123,In_1796);
nand U460 (N_460,In_1192,In_1128);
nand U461 (N_461,In_2299,In_2052);
and U462 (N_462,In_2437,In_1666);
or U463 (N_463,In_2229,In_1043);
xnor U464 (N_464,In_845,In_1068);
nand U465 (N_465,In_1224,In_1801);
nor U466 (N_466,In_2201,In_648);
xnor U467 (N_467,In_1904,In_125);
and U468 (N_468,In_2230,In_1025);
xor U469 (N_469,In_1765,In_346);
or U470 (N_470,In_2469,In_2440);
xnor U471 (N_471,In_223,In_924);
xnor U472 (N_472,In_230,In_1084);
xor U473 (N_473,In_1529,In_1274);
nor U474 (N_474,In_1162,In_2417);
xnor U475 (N_475,In_2273,In_874);
or U476 (N_476,In_1770,In_1147);
nor U477 (N_477,In_153,In_1539);
or U478 (N_478,In_1177,In_2429);
and U479 (N_479,In_2473,In_1152);
and U480 (N_480,In_1350,In_287);
xor U481 (N_481,In_579,In_747);
nand U482 (N_482,In_1589,In_862);
xor U483 (N_483,In_891,In_1028);
xor U484 (N_484,In_1183,In_1205);
nor U485 (N_485,In_1676,In_101);
nand U486 (N_486,In_1239,In_1366);
nor U487 (N_487,In_2194,In_1883);
or U488 (N_488,In_1650,In_1536);
nand U489 (N_489,In_1404,In_1368);
and U490 (N_490,In_474,In_2408);
xnor U491 (N_491,In_1856,In_1681);
and U492 (N_492,In_428,In_2105);
or U493 (N_493,In_1399,In_2155);
or U494 (N_494,In_1361,In_1048);
xnor U495 (N_495,In_1088,In_1417);
xnor U496 (N_496,In_1583,In_1953);
nor U497 (N_497,In_978,In_2097);
xnor U498 (N_498,In_2434,In_398);
and U499 (N_499,In_246,In_357);
xnor U500 (N_500,In_1149,In_493);
or U501 (N_501,In_437,In_309);
nor U502 (N_502,In_1017,In_279);
or U503 (N_503,In_1654,In_1298);
or U504 (N_504,In_1941,In_1432);
and U505 (N_505,In_717,In_1323);
nand U506 (N_506,In_1784,In_1622);
or U507 (N_507,In_401,In_2183);
nand U508 (N_508,In_841,In_1995);
and U509 (N_509,In_2120,In_738);
nor U510 (N_510,In_83,In_1617);
or U511 (N_511,In_1518,In_1479);
nand U512 (N_512,In_1234,In_113);
and U513 (N_513,In_1932,In_1386);
or U514 (N_514,In_457,In_1407);
xnor U515 (N_515,In_750,In_2190);
and U516 (N_516,In_1877,In_811);
nand U517 (N_517,In_1237,In_531);
nand U518 (N_518,In_1601,In_2438);
xor U519 (N_519,In_1999,In_1935);
nand U520 (N_520,In_1669,In_2465);
and U521 (N_521,In_2057,In_1535);
or U522 (N_522,In_1701,In_1792);
nor U523 (N_523,In_1867,In_1109);
nand U524 (N_524,In_1299,In_2027);
nand U525 (N_525,In_1573,In_1304);
nand U526 (N_526,In_2444,In_847);
and U527 (N_527,In_1850,In_2023);
nand U528 (N_528,In_1698,In_222);
or U529 (N_529,In_1748,In_1306);
nor U530 (N_530,In_500,In_2433);
xnor U531 (N_531,In_2109,In_1317);
xnor U532 (N_532,In_187,In_2436);
and U533 (N_533,In_859,In_1901);
nor U534 (N_534,In_985,In_1453);
or U535 (N_535,In_1503,In_1463);
nor U536 (N_536,In_1245,In_1917);
nor U537 (N_537,In_607,In_1548);
nor U538 (N_538,In_1322,In_1616);
nor U539 (N_539,In_2410,In_1847);
nand U540 (N_540,In_2447,In_1153);
or U541 (N_541,In_696,In_462);
nand U542 (N_542,In_356,In_34);
nor U543 (N_543,In_827,In_1056);
or U544 (N_544,In_146,In_1387);
nor U545 (N_545,In_1921,In_68);
nor U546 (N_546,In_124,In_1944);
or U547 (N_547,In_1486,In_529);
and U548 (N_548,In_2303,In_1907);
or U549 (N_549,In_1437,In_1723);
and U550 (N_550,In_198,In_2078);
or U551 (N_551,In_2063,In_424);
nor U552 (N_552,In_2147,In_551);
nor U553 (N_553,In_2119,In_2151);
or U554 (N_554,In_960,In_24);
nor U555 (N_555,In_569,In_2043);
and U556 (N_556,In_2423,In_2064);
and U557 (N_557,In_826,In_1342);
xor U558 (N_558,In_2042,In_2238);
nand U559 (N_559,In_429,In_997);
xor U560 (N_560,In_1874,In_2313);
nor U561 (N_561,In_2421,In_721);
nor U562 (N_562,In_2174,In_1620);
or U563 (N_563,In_1011,In_345);
xor U564 (N_564,In_1757,In_2074);
nor U565 (N_565,In_119,In_885);
nand U566 (N_566,In_593,In_543);
and U567 (N_567,In_127,In_386);
nand U568 (N_568,In_1199,In_1467);
nand U569 (N_569,In_1715,In_2215);
xnor U570 (N_570,In_1071,In_302);
and U571 (N_571,In_889,In_1316);
nor U572 (N_572,In_2038,In_791);
nor U573 (N_573,In_1773,In_1070);
or U574 (N_574,In_1731,In_1464);
or U575 (N_575,In_2344,In_1751);
xor U576 (N_576,In_249,In_452);
xor U577 (N_577,In_2024,In_525);
or U578 (N_578,In_517,In_1427);
or U579 (N_579,In_567,In_1439);
nand U580 (N_580,In_927,In_308);
nand U581 (N_581,In_2011,In_271);
nor U582 (N_582,In_451,In_1624);
and U583 (N_583,In_154,In_1031);
nand U584 (N_584,In_1555,In_22);
nor U585 (N_585,In_1553,In_1489);
nand U586 (N_586,In_965,In_2285);
and U587 (N_587,In_742,In_1724);
nand U588 (N_588,In_376,In_840);
nor U589 (N_589,In_1575,In_1384);
xnor U590 (N_590,In_2084,In_858);
xnor U591 (N_591,In_951,In_183);
nand U592 (N_592,In_1512,In_118);
and U593 (N_593,In_315,In_618);
and U594 (N_594,In_1015,In_1668);
and U595 (N_595,In_566,In_180);
xnor U596 (N_596,In_1851,In_494);
nand U597 (N_597,In_2257,In_210);
xnor U598 (N_598,In_2470,In_1372);
or U599 (N_599,In_869,In_1490);
nand U600 (N_600,In_1457,In_1580);
and U601 (N_601,In_1340,In_256);
and U602 (N_602,In_1945,In_19);
and U603 (N_603,In_509,In_1782);
xor U604 (N_604,In_2256,In_589);
xnor U605 (N_605,In_2460,In_1363);
nor U606 (N_606,In_1720,In_1302);
or U607 (N_607,In_2371,In_1604);
nor U608 (N_608,In_1881,In_680);
and U609 (N_609,In_1844,In_1728);
and U610 (N_610,In_2331,In_253);
nand U611 (N_611,In_1805,In_2345);
xnor U612 (N_612,In_1951,In_1242);
xor U613 (N_613,In_303,In_1971);
xor U614 (N_614,In_2386,In_1510);
xor U615 (N_615,In_1732,In_785);
and U616 (N_616,In_992,In_1544);
nand U617 (N_617,In_2090,In_1058);
xnor U618 (N_618,In_1440,In_1794);
or U619 (N_619,In_655,In_756);
xnor U620 (N_620,In_147,In_2449);
and U621 (N_621,In_272,In_275);
nor U622 (N_622,In_161,In_549);
and U623 (N_623,In_2442,In_1283);
xnor U624 (N_624,In_432,In_2267);
and U625 (N_625,In_1886,In_1615);
nor U626 (N_626,In_2394,In_2363);
nor U627 (N_627,In_1145,In_914);
nor U628 (N_628,In_835,In_1810);
nor U629 (N_629,In_2448,In_2296);
xnor U630 (N_630,In_1477,In_2466);
and U631 (N_631,In_1837,In_766);
xor U632 (N_632,In_1606,In_2492);
nor U633 (N_633,In_2287,In_2349);
nor U634 (N_634,In_768,In_1130);
and U635 (N_635,In_1102,In_2016);
nor U636 (N_636,In_1158,In_2076);
xor U637 (N_637,In_861,In_1985);
xor U638 (N_638,In_1089,In_2009);
nor U639 (N_639,In_720,In_151);
nor U640 (N_640,In_340,In_959);
nand U641 (N_641,In_995,In_2144);
xor U642 (N_642,In_784,In_1980);
nand U643 (N_643,In_1377,In_1557);
xnor U644 (N_644,In_1127,In_408);
and U645 (N_645,In_1871,In_1638);
and U646 (N_646,In_1311,In_806);
and U647 (N_647,In_751,In_259);
xnor U648 (N_648,In_1605,In_1092);
xnor U649 (N_649,In_1329,In_399);
nand U650 (N_650,In_327,In_586);
and U651 (N_651,In_2040,In_130);
and U652 (N_652,In_614,In_2150);
xor U653 (N_653,In_177,In_1279);
nand U654 (N_654,In_1531,In_381);
or U655 (N_655,In_819,In_1923);
xor U656 (N_656,In_1151,In_1097);
xnor U657 (N_657,In_1740,In_366);
nand U658 (N_658,In_1963,In_695);
nand U659 (N_659,In_1636,In_1326);
and U660 (N_660,In_2439,In_608);
xor U661 (N_661,In_2153,In_2232);
nand U662 (N_662,In_715,In_634);
nor U663 (N_663,In_2278,In_1116);
xor U664 (N_664,In_1655,In_314);
or U665 (N_665,In_1296,In_2284);
nand U666 (N_666,In_1169,In_30);
nand U667 (N_667,In_782,In_2234);
or U668 (N_668,In_1238,In_434);
or U669 (N_669,In_1406,In_2261);
xnor U670 (N_670,In_664,In_1497);
nor U671 (N_671,In_1282,In_994);
nor U672 (N_672,In_333,In_1726);
and U673 (N_673,In_269,In_247);
nor U674 (N_674,In_1697,In_2166);
or U675 (N_675,In_2376,In_550);
xor U676 (N_676,In_1630,In_1778);
nand U677 (N_677,In_1649,In_216);
or U678 (N_678,In_1542,In_276);
or U679 (N_679,In_1696,In_1222);
xnor U680 (N_680,In_523,In_1754);
and U681 (N_681,In_779,In_737);
nor U682 (N_682,In_2136,In_2391);
xor U683 (N_683,In_1900,In_1394);
xor U684 (N_684,In_611,In_1976);
and U685 (N_685,In_1702,In_1050);
and U686 (N_686,In_1381,In_6);
or U687 (N_687,In_1915,In_419);
and U688 (N_688,In_337,In_754);
nor U689 (N_689,In_2279,In_84);
nand U690 (N_690,In_2242,In_1783);
and U691 (N_691,In_2101,In_813);
nand U692 (N_692,In_1752,In_80);
or U693 (N_693,In_1964,In_1897);
xor U694 (N_694,In_511,In_1496);
or U695 (N_695,In_76,In_268);
xnor U696 (N_696,In_1658,In_1452);
xor U697 (N_697,In_986,In_2062);
and U698 (N_698,In_1172,In_1632);
xnor U699 (N_699,In_1834,In_2085);
and U700 (N_700,In_414,In_2050);
nor U701 (N_701,In_2114,In_2319);
nor U702 (N_702,In_2246,In_2312);
nand U703 (N_703,In_1685,In_1835);
nand U704 (N_704,In_1664,In_2032);
xnor U705 (N_705,In_1515,In_2037);
and U706 (N_706,In_2079,In_2479);
nor U707 (N_707,In_204,In_2446);
or U708 (N_708,In_0,In_897);
and U709 (N_709,In_1928,In_1475);
and U710 (N_710,In_673,In_587);
nand U711 (N_711,In_2029,In_1524);
nor U712 (N_712,In_1428,In_790);
or U713 (N_713,In_1255,In_2220);
and U714 (N_714,In_1051,In_1091);
xnor U715 (N_715,In_1357,In_1712);
and U716 (N_716,In_2060,In_1358);
nand U717 (N_717,In_316,In_305);
xnor U718 (N_718,In_807,In_752);
or U719 (N_719,In_2015,In_1961);
xnor U720 (N_720,In_505,In_969);
or U721 (N_721,In_391,In_725);
or U722 (N_722,In_1454,In_1772);
nor U723 (N_723,In_388,In_653);
or U724 (N_724,In_2254,In_1922);
or U725 (N_725,In_2096,In_799);
xnor U726 (N_726,In_1619,In_2249);
or U727 (N_727,In_539,In_264);
and U728 (N_728,In_489,In_2412);
and U729 (N_729,In_2213,In_1000);
nand U730 (N_730,In_1391,In_1996);
nor U731 (N_731,In_659,In_1699);
nor U732 (N_732,In_1253,In_2160);
and U733 (N_733,In_1506,In_2046);
nor U734 (N_734,In_1865,In_426);
xnor U735 (N_735,In_131,In_1833);
xnor U736 (N_736,In_583,In_1286);
nor U737 (N_737,In_159,In_2218);
or U738 (N_738,In_1618,In_2329);
or U739 (N_739,In_1482,In_2143);
or U740 (N_740,In_1132,In_2171);
or U741 (N_741,In_1647,In_475);
or U742 (N_742,In_1891,In_1533);
and U743 (N_743,In_1528,In_2397);
and U744 (N_744,In_454,In_395);
nor U745 (N_745,In_258,In_1978);
or U746 (N_746,In_1374,In_450);
nand U747 (N_747,In_640,In_722);
and U748 (N_748,In_1403,In_410);
and U749 (N_749,In_1348,In_236);
or U750 (N_750,In_1215,In_1478);
and U751 (N_751,In_2159,In_1217);
or U752 (N_752,In_1378,In_39);
or U753 (N_753,In_353,In_1138);
and U754 (N_754,In_958,In_59);
and U755 (N_755,In_719,In_1656);
or U756 (N_756,In_1435,In_1256);
xor U757 (N_757,In_2126,In_1514);
xnor U758 (N_758,In_2031,In_1854);
or U759 (N_759,In_1230,In_1144);
xnor U760 (N_760,In_33,In_326);
and U761 (N_761,In_1135,In_763);
nor U762 (N_762,In_1424,In_2463);
xnor U763 (N_763,In_2411,In_942);
xnor U764 (N_764,In_1207,In_51);
xor U765 (N_765,In_907,In_418);
or U766 (N_766,In_126,In_2388);
nand U767 (N_767,In_2351,In_2185);
or U768 (N_768,In_1287,In_2041);
and U769 (N_769,In_1466,In_60);
and U770 (N_770,In_943,In_561);
nand U771 (N_771,In_767,In_849);
nor U772 (N_772,In_1520,In_28);
nand U773 (N_773,In_46,In_1046);
nand U774 (N_774,In_58,In_581);
or U775 (N_775,In_1674,In_1029);
nor U776 (N_776,In_266,In_317);
and U777 (N_777,In_2360,In_1852);
nand U778 (N_778,In_706,In_1027);
and U779 (N_779,In_100,In_909);
nand U780 (N_780,In_701,In_2);
or U781 (N_781,In_526,In_2217);
nand U782 (N_782,In_1558,In_1044);
nand U783 (N_783,In_336,In_2288);
nor U784 (N_784,In_427,In_1967);
nand U785 (N_785,In_714,In_221);
and U786 (N_786,In_1359,In_163);
and U787 (N_787,In_466,In_1957);
and U788 (N_788,In_2318,In_1760);
or U789 (N_789,In_2342,In_1349);
nand U790 (N_790,In_1082,In_548);
and U791 (N_791,In_1450,In_1554);
nor U792 (N_792,In_518,In_1203);
nand U793 (N_793,In_431,In_1142);
nor U794 (N_794,In_1771,In_1802);
or U795 (N_795,In_322,In_1252);
nand U796 (N_796,In_2401,In_1018);
or U797 (N_797,In_2044,In_343);
and U798 (N_798,In_1566,In_354);
nor U799 (N_799,In_482,In_535);
nand U800 (N_800,In_277,In_2207);
nand U801 (N_801,In_2399,In_1290);
or U802 (N_802,In_757,In_1925);
or U803 (N_803,In_2204,In_512);
and U804 (N_804,In_2182,In_1155);
xnor U805 (N_805,In_2263,In_469);
nand U806 (N_806,In_2382,In_2472);
xnor U807 (N_807,In_218,In_1882);
xor U808 (N_808,In_1692,In_718);
xnor U809 (N_809,In_2385,In_932);
nand U810 (N_810,In_1644,In_203);
nor U811 (N_811,In_1293,In_1912);
nor U812 (N_812,In_1918,In_1408);
nor U813 (N_813,In_674,In_783);
nor U814 (N_814,In_2198,In_402);
nand U815 (N_815,In_2383,In_514);
xnor U816 (N_816,In_2292,In_1218);
nor U817 (N_817,In_968,In_257);
xor U818 (N_818,In_86,In_1926);
and U819 (N_819,In_1341,In_495);
and U820 (N_820,In_2280,In_936);
nor U821 (N_821,In_2156,In_2165);
or U822 (N_822,In_1276,In_1979);
or U823 (N_823,In_852,In_1769);
nor U824 (N_824,In_533,In_1623);
nand U825 (N_825,In_1578,In_227);
and U826 (N_826,In_471,In_796);
or U827 (N_827,In_239,In_933);
and U828 (N_828,In_1889,In_855);
xor U829 (N_829,In_730,In_1187);
nand U830 (N_830,In_2124,In_1916);
nor U831 (N_831,In_2179,In_2348);
nand U832 (N_832,In_1275,In_172);
or U833 (N_833,In_1202,In_63);
nand U834 (N_834,In_743,In_1110);
and U835 (N_835,In_1729,In_1310);
xnor U836 (N_836,In_605,In_1365);
nand U837 (N_837,In_729,In_639);
nor U838 (N_838,In_1420,In_245);
nor U839 (N_839,In_476,In_1448);
and U840 (N_840,In_920,In_2387);
nor U841 (N_841,In_325,In_815);
nor U842 (N_842,In_2467,In_832);
xor U843 (N_843,In_1176,In_1790);
and U844 (N_844,In_1103,In_1442);
xor U845 (N_845,In_2163,In_2237);
and U846 (N_846,In_394,In_95);
and U847 (N_847,In_809,In_584);
xnor U848 (N_848,In_1787,In_104);
nand U849 (N_849,In_332,In_1948);
or U850 (N_850,In_734,In_1313);
and U851 (N_851,In_1331,In_2070);
xnor U852 (N_852,In_112,In_844);
or U853 (N_853,In_710,In_460);
nor U854 (N_854,In_1596,In_171);
nand U855 (N_855,In_1072,In_1264);
or U856 (N_856,In_1473,In_1860);
or U857 (N_857,In_1839,In_575);
and U858 (N_858,In_764,In_1436);
nor U859 (N_859,In_682,In_194);
and U860 (N_860,In_47,In_1014);
and U861 (N_861,In_771,In_1966);
and U862 (N_862,In_2200,In_926);
nand U863 (N_863,In_1893,In_1434);
xor U864 (N_864,In_625,In_179);
nand U865 (N_865,In_1005,In_987);
or U866 (N_866,In_1627,In_727);
xor U867 (N_867,In_2100,In_251);
nor U868 (N_868,In_777,In_699);
and U869 (N_869,In_472,In_435);
nand U870 (N_870,In_254,In_1492);
nand U871 (N_871,In_1301,In_1826);
nor U872 (N_872,In_1738,In_1037);
nor U873 (N_873,In_1861,In_139);
xnor U874 (N_874,In_1561,In_1243);
nand U875 (N_875,In_953,In_2336);
xor U876 (N_876,In_1064,In_339);
nor U877 (N_877,In_1954,In_1661);
or U878 (N_878,In_491,In_902);
nor U879 (N_879,In_1602,In_18);
nor U880 (N_880,In_2072,In_1968);
xor U881 (N_881,In_1023,In_1312);
nor U882 (N_882,In_1001,In_2310);
nor U883 (N_883,In_473,In_1033);
nand U884 (N_884,In_82,In_1133);
or U885 (N_885,In_1705,In_1268);
xor U886 (N_886,In_1446,In_140);
or U887 (N_887,In_2274,In_904);
nor U888 (N_888,In_1679,In_665);
and U889 (N_889,In_235,In_772);
or U890 (N_890,In_546,In_837);
or U891 (N_891,In_672,In_2014);
xor U892 (N_892,In_138,In_731);
or U893 (N_893,In_1260,In_420);
and U894 (N_894,In_2140,In_215);
or U895 (N_895,In_1369,In_2123);
xnor U896 (N_896,In_1415,In_440);
or U897 (N_897,In_778,In_974);
or U898 (N_898,In_1426,In_1742);
and U899 (N_899,In_952,In_1062);
nor U900 (N_900,In_1739,In_2425);
nand U901 (N_901,In_1809,In_1204);
nand U902 (N_902,In_857,In_691);
and U903 (N_903,In_1166,In_1711);
nand U904 (N_904,In_232,In_871);
and U905 (N_905,In_1458,In_629);
or U906 (N_906,In_1226,In_571);
nand U907 (N_907,In_610,In_1221);
and U908 (N_908,In_1610,In_1564);
nor U909 (N_909,In_480,In_199);
nor U910 (N_910,In_110,In_342);
nor U911 (N_911,In_1030,In_1065);
and U912 (N_912,In_580,In_1047);
nand U913 (N_913,In_1396,In_1509);
nand U914 (N_914,In_439,In_1272);
and U915 (N_915,In_733,In_2195);
or U916 (N_916,In_360,In_667);
nor U917 (N_917,In_2334,In_2317);
nand U918 (N_918,In_644,In_1178);
xnor U919 (N_919,In_801,In_488);
xnor U920 (N_920,In_928,In_2235);
or U921 (N_921,In_1040,In_2338);
xnor U922 (N_922,In_2398,In_800);
and U923 (N_923,In_2102,In_2088);
and U924 (N_924,In_1824,In_694);
and U925 (N_925,In_2080,In_2240);
or U926 (N_926,In_1020,In_704);
and U927 (N_927,In_609,In_2191);
nor U928 (N_928,In_1013,In_1143);
nand U929 (N_929,In_1502,In_2259);
or U930 (N_930,In_1689,In_528);
or U931 (N_931,In_2054,In_1541);
nand U932 (N_932,In_412,In_804);
and U933 (N_933,In_1843,In_1597);
and U934 (N_934,In_964,In_1708);
and U935 (N_935,In_534,In_168);
nand U936 (N_936,In_31,In_265);
nor U937 (N_937,In_2033,In_1154);
xnor U938 (N_938,In_1141,In_2089);
or U939 (N_939,In_1673,In_285);
or U940 (N_940,In_520,In_1574);
xor U941 (N_941,In_2456,In_212);
nor U942 (N_942,In_1829,In_1593);
or U943 (N_943,In_116,In_2332);
or U944 (N_944,In_1981,In_62);
or U945 (N_945,In_623,In_1042);
nor U946 (N_946,In_2424,In_1235);
nor U947 (N_947,In_821,In_1651);
or U948 (N_948,In_338,In_1388);
nor U949 (N_949,In_1988,In_828);
nand U950 (N_950,In_638,In_2053);
and U951 (N_951,In_947,In_1577);
or U952 (N_952,In_2189,In_1021);
nand U953 (N_953,In_1104,In_189);
or U954 (N_954,In_1447,In_1269);
nor U955 (N_955,In_1947,In_787);
nand U956 (N_956,In_590,In_912);
nand U957 (N_957,In_383,In_1131);
and U958 (N_958,In_2364,In_2295);
nor U959 (N_959,In_1225,In_598);
nor U960 (N_960,In_2161,In_250);
nand U961 (N_961,In_1148,In_888);
xor U962 (N_962,In_2099,In_2322);
nor U963 (N_963,In_2352,In_1892);
and U964 (N_964,In_1598,In_1584);
nor U965 (N_965,In_1146,In_380);
xnor U966 (N_966,In_1734,In_723);
xnor U967 (N_967,In_558,In_2094);
nor U968 (N_968,In_612,In_1774);
nor U969 (N_969,In_98,In_513);
and U970 (N_970,In_166,In_622);
or U971 (N_971,In_389,In_1167);
or U972 (N_972,In_56,In_670);
and U973 (N_973,In_1830,In_1863);
xnor U974 (N_974,In_72,In_390);
nand U975 (N_975,In_2214,In_2488);
and U976 (N_976,In_2127,In_108);
or U977 (N_977,In_1920,In_44);
nand U978 (N_978,In_908,In_467);
xor U979 (N_979,In_350,In_1797);
and U980 (N_980,In_900,In_201);
xor U981 (N_981,In_2103,In_2337);
or U982 (N_982,In_406,In_2012);
nand U983 (N_983,In_176,In_1590);
or U984 (N_984,In_378,In_228);
nor U985 (N_985,In_1343,In_870);
xor U986 (N_986,In_1160,In_382);
nand U987 (N_987,In_572,In_2227);
and U988 (N_988,In_2426,In_2184);
and U989 (N_989,In_1401,In_788);
nand U990 (N_990,In_745,In_1879);
nand U991 (N_991,In_2175,In_692);
nand U992 (N_992,In_2435,In_1887);
nand U993 (N_993,In_296,In_2378);
and U994 (N_994,In_950,In_864);
or U995 (N_995,In_363,In_1246);
nand U996 (N_996,In_1165,In_2392);
nand U997 (N_997,In_2381,In_2117);
and U998 (N_998,In_1675,In_702);
nor U999 (N_999,In_1438,In_1307);
nor U1000 (N_1000,In_1903,In_261);
nor U1001 (N_1001,In_1472,In_712);
and U1002 (N_1002,In_1498,In_289);
nand U1003 (N_1003,In_293,In_334);
or U1004 (N_1004,In_497,In_1511);
xnor U1005 (N_1005,In_2471,In_631);
and U1006 (N_1006,In_713,In_347);
or U1007 (N_1007,In_1946,In_23);
or U1008 (N_1008,In_1493,In_299);
nand U1009 (N_1009,In_1314,In_186);
xnor U1010 (N_1010,In_1251,In_45);
nand U1011 (N_1011,In_1480,In_217);
or U1012 (N_1012,In_1462,In_2428);
and U1013 (N_1013,In_1049,In_2222);
and U1014 (N_1014,In_368,In_416);
nand U1015 (N_1015,In_739,In_1335);
nor U1016 (N_1016,In_1931,In_35);
nand U1017 (N_1017,In_1327,In_1094);
xor U1018 (N_1018,In_1828,In_1108);
and U1019 (N_1019,In_2083,In_1827);
xor U1020 (N_1020,In_2262,In_208);
or U1021 (N_1021,In_448,In_793);
nor U1022 (N_1022,In_324,In_1445);
and U1023 (N_1023,In_1347,In_2001);
nor U1024 (N_1024,In_812,In_2164);
and U1025 (N_1025,In_760,In_2476);
nand U1026 (N_1026,In_1284,In_7);
nor U1027 (N_1027,In_195,In_2316);
nor U1028 (N_1028,In_2343,In_501);
nand U1029 (N_1029,In_1934,In_1880);
xor U1030 (N_1030,In_2281,In_123);
nand U1031 (N_1031,In_1280,In_158);
and U1032 (N_1032,In_560,In_1081);
xor U1033 (N_1033,In_536,In_2091);
xor U1034 (N_1034,In_15,In_2464);
or U1035 (N_1035,In_522,In_894);
or U1036 (N_1036,In_1330,In_492);
xor U1037 (N_1037,In_660,In_2000);
nor U1038 (N_1038,In_949,In_209);
and U1039 (N_1039,In_38,In_2223);
nand U1040 (N_1040,In_1093,In_2289);
nor U1041 (N_1041,In_1099,In_54);
and U1042 (N_1042,In_1678,In_1443);
xor U1043 (N_1043,In_570,In_541);
and U1044 (N_1044,In_1315,In_1587);
or U1045 (N_1045,In_306,In_1231);
and U1046 (N_1046,In_938,In_1111);
xnor U1047 (N_1047,In_278,In_2045);
nand U1048 (N_1048,In_441,In_1775);
xor U1049 (N_1049,In_921,In_915);
nand U1050 (N_1050,In_2130,In_1906);
xnor U1051 (N_1051,In_1820,In_666);
nor U1052 (N_1052,In_990,In_2121);
xnor U1053 (N_1053,In_1191,In_2167);
nand U1054 (N_1054,In_732,In_2106);
xor U1055 (N_1055,In_85,In_1840);
nor U1056 (N_1056,In_133,In_600);
nand U1057 (N_1057,In_2480,In_470);
xor U1058 (N_1058,In_2335,In_1285);
or U1059 (N_1059,In_1076,In_1884);
xor U1060 (N_1060,In_2367,In_318);
xor U1061 (N_1061,In_510,In_1379);
xnor U1062 (N_1062,In_1373,In_157);
xnor U1063 (N_1063,In_1266,In_1038);
nand U1064 (N_1064,In_2441,In_181);
nor U1065 (N_1065,In_1370,In_1914);
nand U1066 (N_1066,In_2098,In_1766);
xor U1067 (N_1067,In_1136,In_415);
nand U1068 (N_1068,In_99,In_2270);
and U1069 (N_1069,In_1709,In_1611);
xor U1070 (N_1070,In_939,In_2374);
nand U1071 (N_1071,In_2066,In_2202);
or U1072 (N_1072,In_77,In_1818);
or U1073 (N_1073,In_1265,In_2022);
nand U1074 (N_1074,In_624,In_1687);
xnor U1075 (N_1075,In_1083,In_1532);
xor U1076 (N_1076,In_1788,In_2154);
and U1077 (N_1077,In_1273,In_979);
and U1078 (N_1078,In_2082,In_233);
or U1079 (N_1079,In_164,In_1175);
xnor U1080 (N_1080,In_746,In_1798);
and U1081 (N_1081,In_2221,In_559);
nand U1082 (N_1082,In_1334,In_613);
xnor U1083 (N_1083,In_884,In_2377);
xor U1084 (N_1084,In_1713,In_1609);
and U1085 (N_1085,In_2304,In_585);
nor U1086 (N_1086,In_1530,In_2056);
xnor U1087 (N_1087,In_786,In_2402);
xor U1088 (N_1088,In_477,In_330);
and U1089 (N_1089,In_1958,In_769);
and U1090 (N_1090,In_2048,In_973);
nand U1091 (N_1091,In_252,In_1517);
xnor U1092 (N_1092,In_970,In_2405);
or U1093 (N_1093,In_2193,In_438);
or U1094 (N_1094,In_2087,In_1607);
xnor U1095 (N_1095,In_1319,In_313);
or U1096 (N_1096,In_1259,In_2362);
or U1097 (N_1097,In_1431,In_107);
and U1098 (N_1098,In_1419,In_26);
nor U1099 (N_1099,In_1355,In_2107);
nor U1100 (N_1100,In_2264,In_563);
xnor U1101 (N_1101,In_2172,In_663);
and U1102 (N_1102,In_2196,In_1411);
xor U1103 (N_1103,In_1523,In_2314);
nor U1104 (N_1104,In_578,In_2051);
nand U1105 (N_1105,In_1571,In_2482);
nand U1106 (N_1106,In_2419,In_115);
nor U1107 (N_1107,In_65,In_1425);
nor U1108 (N_1108,In_2210,In_11);
nand U1109 (N_1109,In_372,In_1565);
nand U1110 (N_1110,In_851,In_2396);
or U1111 (N_1111,In_1258,In_1232);
nor U1112 (N_1112,In_2233,In_70);
nor U1113 (N_1113,In_1626,In_323);
xor U1114 (N_1114,In_1337,In_671);
and U1115 (N_1115,In_1579,In_2474);
or U1116 (N_1116,In_1241,In_2205);
or U1117 (N_1117,In_2430,In_1336);
and U1118 (N_1118,In_1240,In_4);
xnor U1119 (N_1119,In_954,In_2248);
xor U1120 (N_1120,In_1008,In_2007);
xor U1121 (N_1121,In_616,In_1393);
and U1122 (N_1122,In_636,In_156);
nand U1123 (N_1123,In_36,In_1695);
xnor U1124 (N_1124,In_21,In_2333);
or U1125 (N_1125,In_1612,In_1257);
nand U1126 (N_1126,In_557,In_241);
nand U1127 (N_1127,In_705,In_1909);
xnor U1128 (N_1128,In_348,In_2021);
nor U1129 (N_1129,In_234,In_400);
or U1130 (N_1130,In_1188,In_1095);
and U1131 (N_1131,In_2118,In_1483);
nor U1132 (N_1132,In_1725,In_1220);
nand U1133 (N_1133,In_2228,In_2146);
and U1134 (N_1134,In_225,In_29);
nor U1135 (N_1135,In_12,In_1628);
nand U1136 (N_1136,In_1894,In_202);
and U1137 (N_1137,In_1940,In_483);
and U1138 (N_1138,In_2269,In_1986);
nand U1139 (N_1139,In_1032,In_229);
or U1140 (N_1140,In_1933,In_890);
and U1141 (N_1141,In_1471,In_92);
xor U1142 (N_1142,In_2086,In_773);
or U1143 (N_1143,In_2030,In_1086);
or U1144 (N_1144,In_1634,In_169);
and U1145 (N_1145,In_1800,In_1125);
nand U1146 (N_1146,In_944,In_1803);
nand U1147 (N_1147,In_481,In_1974);
nand U1148 (N_1148,In_1992,In_2158);
nand U1149 (N_1149,In_1444,In_1201);
nand U1150 (N_1150,In_2092,In_2495);
and U1151 (N_1151,In_1171,In_16);
nor U1152 (N_1152,In_630,In_669);
and U1153 (N_1153,In_1324,In_1586);
nor U1154 (N_1154,In_1677,In_1924);
nor U1155 (N_1155,In_1743,In_2244);
or U1156 (N_1156,In_297,In_2178);
nand U1157 (N_1157,In_1118,In_1526);
and U1158 (N_1158,In_387,In_1485);
xor U1159 (N_1159,In_867,In_1288);
and U1160 (N_1160,In_32,In_2368);
nor U1161 (N_1161,In_2432,In_224);
xor U1162 (N_1162,In_1815,In_362);
or U1163 (N_1163,In_53,In_1376);
and U1164 (N_1164,In_1303,In_2206);
xor U1165 (N_1165,In_74,In_1746);
xor U1166 (N_1166,In_2358,In_1308);
nand U1167 (N_1167,In_1640,In_1570);
and U1168 (N_1168,In_761,In_1898);
xnor U1169 (N_1169,In_1534,In_298);
nand U1170 (N_1170,In_1504,In_556);
xnor U1171 (N_1171,In_643,In_262);
nor U1172 (N_1172,In_818,In_726);
nand U1173 (N_1173,In_999,In_1182);
xnor U1174 (N_1174,In_1012,In_2135);
nor U1175 (N_1175,In_736,In_2142);
nor U1176 (N_1176,In_214,In_896);
xnor U1177 (N_1177,In_1973,In_993);
or U1178 (N_1178,In_1707,In_1637);
nor U1179 (N_1179,In_1433,In_96);
nand U1180 (N_1180,In_2379,In_280);
nand U1181 (N_1181,In_1039,In_2152);
nand U1182 (N_1182,In_1767,In_595);
or U1183 (N_1183,In_1563,In_1233);
and U1184 (N_1184,In_1939,In_2008);
nand U1185 (N_1185,In_946,In_1848);
nor U1186 (N_1186,In_1849,In_2290);
nor U1187 (N_1187,In_1139,In_937);
nor U1188 (N_1188,In_1984,In_582);
nor U1189 (N_1189,In_540,In_2308);
nor U1190 (N_1190,In_2216,In_1332);
or U1191 (N_1191,In_1250,In_1328);
and U1192 (N_1192,In_2297,In_981);
or U1193 (N_1193,In_498,In_1150);
nor U1194 (N_1194,In_940,In_1870);
nand U1195 (N_1195,In_1872,In_2458);
nor U1196 (N_1196,In_1859,In_716);
xor U1197 (N_1197,In_2115,In_923);
xnor U1198 (N_1198,In_1470,In_989);
xnor U1199 (N_1199,In_1277,In_370);
and U1200 (N_1200,In_499,In_1140);
or U1201 (N_1201,In_2125,In_1667);
xor U1202 (N_1202,In_459,In_1060);
nor U1203 (N_1203,In_2025,In_1026);
and U1204 (N_1204,In_486,In_2162);
and U1205 (N_1205,In_2462,In_1763);
and U1206 (N_1206,In_384,In_814);
nor U1207 (N_1207,In_645,In_405);
nor U1208 (N_1208,In_1822,In_621);
or U1209 (N_1209,In_789,In_144);
or U1210 (N_1210,In_291,In_679);
xnor U1211 (N_1211,In_2132,In_808);
xor U1212 (N_1212,In_2209,In_1198);
nand U1213 (N_1213,In_830,In_1491);
nand U1214 (N_1214,In_562,In_2133);
or U1215 (N_1215,In_190,In_411);
xnor U1216 (N_1216,In_2404,In_49);
xnor U1217 (N_1217,In_13,In_1762);
xnor U1218 (N_1218,In_1409,In_913);
nand U1219 (N_1219,In_1950,In_1067);
and U1220 (N_1220,In_2330,In_1562);
and U1221 (N_1221,In_962,In_2350);
or U1222 (N_1222,In_661,In_776);
nand U1223 (N_1223,In_1375,In_1174);
and U1224 (N_1224,In_1522,In_1919);
or U1225 (N_1225,In_1318,In_2282);
nand U1226 (N_1226,In_468,In_502);
and U1227 (N_1227,In_1543,In_740);
xnor U1228 (N_1228,In_848,In_1418);
and U1229 (N_1229,In_48,In_1741);
and U1230 (N_1230,In_988,In_2455);
or U1231 (N_1231,In_2268,In_1758);
and U1232 (N_1232,In_87,In_1035);
or U1233 (N_1233,In_1855,In_88);
xor U1234 (N_1234,In_1663,In_312);
and U1235 (N_1235,In_1582,In_396);
nor U1236 (N_1236,In_2328,In_2389);
nor U1237 (N_1237,In_1608,In_111);
or U1238 (N_1238,In_1838,In_1997);
xor U1239 (N_1239,In_2461,In_79);
and U1240 (N_1240,In_850,In_134);
and U1241 (N_1241,In_1625,In_1581);
nor U1242 (N_1242,In_668,In_1345);
xnor U1243 (N_1243,In_1101,In_1074);
nand U1244 (N_1244,In_2211,In_1567);
or U1245 (N_1245,In_1078,In_2272);
and U1246 (N_1246,In_2258,In_905);
nor U1247 (N_1247,In_2275,In_2326);
nand U1248 (N_1248,In_2004,In_1022);
nand U1249 (N_1249,In_839,In_1639);
and U1250 (N_1250,In_2464,In_2311);
and U1251 (N_1251,In_1992,In_2393);
nor U1252 (N_1252,In_1156,In_1209);
nor U1253 (N_1253,In_1134,In_370);
and U1254 (N_1254,In_2135,In_253);
nand U1255 (N_1255,In_1027,In_371);
xnor U1256 (N_1256,In_2318,In_392);
xnor U1257 (N_1257,In_788,In_1062);
or U1258 (N_1258,In_1057,In_2174);
xnor U1259 (N_1259,In_60,In_1070);
and U1260 (N_1260,In_357,In_1468);
and U1261 (N_1261,In_2356,In_2374);
nor U1262 (N_1262,In_395,In_2431);
nand U1263 (N_1263,In_1026,In_1620);
nor U1264 (N_1264,In_732,In_171);
or U1265 (N_1265,In_1006,In_1303);
or U1266 (N_1266,In_68,In_1657);
xor U1267 (N_1267,In_52,In_1740);
and U1268 (N_1268,In_2455,In_2429);
and U1269 (N_1269,In_549,In_1198);
nor U1270 (N_1270,In_549,In_540);
or U1271 (N_1271,In_1546,In_1072);
and U1272 (N_1272,In_1158,In_2072);
nor U1273 (N_1273,In_353,In_2435);
nor U1274 (N_1274,In_155,In_1301);
and U1275 (N_1275,In_495,In_1042);
or U1276 (N_1276,In_76,In_5);
xor U1277 (N_1277,In_437,In_1251);
nand U1278 (N_1278,In_2194,In_1995);
nand U1279 (N_1279,In_651,In_1027);
xnor U1280 (N_1280,In_108,In_2249);
nor U1281 (N_1281,In_1552,In_1742);
and U1282 (N_1282,In_1650,In_2361);
nor U1283 (N_1283,In_1652,In_1200);
nand U1284 (N_1284,In_1305,In_2001);
xnor U1285 (N_1285,In_1980,In_640);
nor U1286 (N_1286,In_2269,In_111);
nand U1287 (N_1287,In_1018,In_2336);
or U1288 (N_1288,In_1276,In_1023);
xnor U1289 (N_1289,In_1169,In_161);
nand U1290 (N_1290,In_469,In_505);
nor U1291 (N_1291,In_13,In_24);
and U1292 (N_1292,In_2431,In_1856);
nor U1293 (N_1293,In_696,In_1610);
nor U1294 (N_1294,In_1497,In_369);
xor U1295 (N_1295,In_1091,In_1113);
xnor U1296 (N_1296,In_1209,In_662);
nor U1297 (N_1297,In_1332,In_2324);
and U1298 (N_1298,In_2289,In_2129);
and U1299 (N_1299,In_447,In_1693);
nand U1300 (N_1300,In_2155,In_246);
nor U1301 (N_1301,In_2315,In_1515);
or U1302 (N_1302,In_935,In_2389);
and U1303 (N_1303,In_2073,In_2151);
and U1304 (N_1304,In_386,In_1423);
xor U1305 (N_1305,In_579,In_976);
and U1306 (N_1306,In_1890,In_1386);
and U1307 (N_1307,In_171,In_108);
or U1308 (N_1308,In_902,In_1145);
nand U1309 (N_1309,In_2032,In_820);
nand U1310 (N_1310,In_765,In_1264);
and U1311 (N_1311,In_784,In_1055);
and U1312 (N_1312,In_2075,In_1282);
nand U1313 (N_1313,In_97,In_1702);
xnor U1314 (N_1314,In_1226,In_481);
or U1315 (N_1315,In_2167,In_379);
nor U1316 (N_1316,In_2470,In_1350);
nand U1317 (N_1317,In_691,In_807);
xnor U1318 (N_1318,In_373,In_267);
or U1319 (N_1319,In_374,In_710);
and U1320 (N_1320,In_365,In_1994);
nor U1321 (N_1321,In_125,In_1013);
or U1322 (N_1322,In_1662,In_2219);
nand U1323 (N_1323,In_985,In_249);
and U1324 (N_1324,In_342,In_1579);
nor U1325 (N_1325,In_1530,In_382);
or U1326 (N_1326,In_78,In_1072);
nor U1327 (N_1327,In_457,In_1054);
xor U1328 (N_1328,In_1679,In_1733);
and U1329 (N_1329,In_983,In_1193);
xnor U1330 (N_1330,In_1802,In_2144);
xor U1331 (N_1331,In_2091,In_1860);
or U1332 (N_1332,In_963,In_848);
xnor U1333 (N_1333,In_816,In_1484);
nand U1334 (N_1334,In_2181,In_1472);
or U1335 (N_1335,In_1062,In_1586);
or U1336 (N_1336,In_2061,In_528);
or U1337 (N_1337,In_2044,In_412);
nor U1338 (N_1338,In_2200,In_2239);
and U1339 (N_1339,In_1297,In_1160);
or U1340 (N_1340,In_264,In_1712);
and U1341 (N_1341,In_2480,In_624);
and U1342 (N_1342,In_2041,In_526);
nor U1343 (N_1343,In_873,In_526);
xnor U1344 (N_1344,In_2141,In_1411);
and U1345 (N_1345,In_998,In_765);
xor U1346 (N_1346,In_1487,In_1686);
nor U1347 (N_1347,In_256,In_724);
nand U1348 (N_1348,In_899,In_1432);
or U1349 (N_1349,In_1424,In_1201);
xor U1350 (N_1350,In_2445,In_2327);
nand U1351 (N_1351,In_392,In_2405);
xor U1352 (N_1352,In_1626,In_2480);
nor U1353 (N_1353,In_1707,In_1693);
and U1354 (N_1354,In_521,In_1990);
and U1355 (N_1355,In_2044,In_219);
nand U1356 (N_1356,In_969,In_1945);
xnor U1357 (N_1357,In_1549,In_830);
nor U1358 (N_1358,In_922,In_250);
nand U1359 (N_1359,In_491,In_473);
nand U1360 (N_1360,In_1424,In_439);
nor U1361 (N_1361,In_2070,In_491);
or U1362 (N_1362,In_1196,In_120);
and U1363 (N_1363,In_511,In_1199);
xnor U1364 (N_1364,In_779,In_1043);
xnor U1365 (N_1365,In_1535,In_1531);
or U1366 (N_1366,In_1896,In_1926);
and U1367 (N_1367,In_878,In_2416);
and U1368 (N_1368,In_387,In_27);
nand U1369 (N_1369,In_296,In_782);
xnor U1370 (N_1370,In_563,In_238);
xnor U1371 (N_1371,In_2157,In_2275);
xor U1372 (N_1372,In_104,In_527);
and U1373 (N_1373,In_773,In_1895);
xor U1374 (N_1374,In_1274,In_1883);
xnor U1375 (N_1375,In_54,In_404);
or U1376 (N_1376,In_2329,In_836);
nor U1377 (N_1377,In_2126,In_1745);
nor U1378 (N_1378,In_1898,In_1906);
and U1379 (N_1379,In_178,In_489);
nor U1380 (N_1380,In_2337,In_2364);
nand U1381 (N_1381,In_1849,In_1314);
nand U1382 (N_1382,In_305,In_1368);
nand U1383 (N_1383,In_301,In_337);
and U1384 (N_1384,In_32,In_1430);
nor U1385 (N_1385,In_1725,In_125);
and U1386 (N_1386,In_1640,In_644);
or U1387 (N_1387,In_136,In_1258);
nor U1388 (N_1388,In_2253,In_1737);
nand U1389 (N_1389,In_686,In_408);
nand U1390 (N_1390,In_505,In_748);
nand U1391 (N_1391,In_1558,In_1772);
nand U1392 (N_1392,In_678,In_710);
nor U1393 (N_1393,In_1397,In_459);
nor U1394 (N_1394,In_1011,In_642);
nand U1395 (N_1395,In_179,In_50);
and U1396 (N_1396,In_828,In_388);
nand U1397 (N_1397,In_1131,In_1539);
or U1398 (N_1398,In_149,In_1790);
nor U1399 (N_1399,In_1779,In_845);
nand U1400 (N_1400,In_258,In_423);
or U1401 (N_1401,In_205,In_986);
or U1402 (N_1402,In_2273,In_2392);
nor U1403 (N_1403,In_1148,In_808);
and U1404 (N_1404,In_523,In_178);
nand U1405 (N_1405,In_2281,In_1070);
and U1406 (N_1406,In_2332,In_2368);
nor U1407 (N_1407,In_180,In_1571);
nand U1408 (N_1408,In_740,In_1526);
and U1409 (N_1409,In_865,In_1762);
xor U1410 (N_1410,In_1000,In_361);
nor U1411 (N_1411,In_1169,In_873);
xnor U1412 (N_1412,In_922,In_1104);
nor U1413 (N_1413,In_1168,In_232);
or U1414 (N_1414,In_634,In_1506);
nor U1415 (N_1415,In_1679,In_727);
or U1416 (N_1416,In_2197,In_1669);
or U1417 (N_1417,In_2037,In_802);
nor U1418 (N_1418,In_2379,In_2498);
nor U1419 (N_1419,In_726,In_2286);
nand U1420 (N_1420,In_1661,In_47);
or U1421 (N_1421,In_2273,In_51);
xnor U1422 (N_1422,In_1476,In_344);
or U1423 (N_1423,In_109,In_2059);
xnor U1424 (N_1424,In_1585,In_1715);
nand U1425 (N_1425,In_1654,In_1911);
nor U1426 (N_1426,In_1625,In_1281);
nand U1427 (N_1427,In_652,In_1375);
nand U1428 (N_1428,In_2354,In_1836);
nor U1429 (N_1429,In_554,In_1926);
xor U1430 (N_1430,In_1099,In_1780);
nor U1431 (N_1431,In_1994,In_2370);
xor U1432 (N_1432,In_587,In_1630);
and U1433 (N_1433,In_824,In_455);
nand U1434 (N_1434,In_1849,In_1880);
and U1435 (N_1435,In_1747,In_1406);
xor U1436 (N_1436,In_209,In_970);
nand U1437 (N_1437,In_1008,In_1604);
xnor U1438 (N_1438,In_4,In_349);
nor U1439 (N_1439,In_659,In_1103);
xnor U1440 (N_1440,In_2297,In_1556);
and U1441 (N_1441,In_696,In_23);
xnor U1442 (N_1442,In_2248,In_141);
xnor U1443 (N_1443,In_1974,In_1446);
nand U1444 (N_1444,In_59,In_1129);
nor U1445 (N_1445,In_1525,In_669);
nor U1446 (N_1446,In_1835,In_1518);
and U1447 (N_1447,In_711,In_2035);
and U1448 (N_1448,In_229,In_2264);
nand U1449 (N_1449,In_512,In_1388);
and U1450 (N_1450,In_1306,In_12);
nand U1451 (N_1451,In_1547,In_405);
and U1452 (N_1452,In_988,In_870);
xnor U1453 (N_1453,In_2036,In_1808);
or U1454 (N_1454,In_1633,In_1946);
nor U1455 (N_1455,In_2256,In_2482);
nor U1456 (N_1456,In_390,In_598);
or U1457 (N_1457,In_2167,In_1242);
nor U1458 (N_1458,In_1194,In_2349);
nor U1459 (N_1459,In_278,In_1287);
or U1460 (N_1460,In_624,In_217);
nand U1461 (N_1461,In_646,In_2318);
nor U1462 (N_1462,In_1486,In_1191);
nand U1463 (N_1463,In_2469,In_1034);
xor U1464 (N_1464,In_1390,In_584);
xor U1465 (N_1465,In_518,In_1334);
nor U1466 (N_1466,In_1745,In_643);
and U1467 (N_1467,In_2056,In_1926);
nand U1468 (N_1468,In_1426,In_2083);
or U1469 (N_1469,In_913,In_814);
or U1470 (N_1470,In_2458,In_538);
nor U1471 (N_1471,In_2191,In_655);
xnor U1472 (N_1472,In_529,In_1981);
xor U1473 (N_1473,In_369,In_1697);
xor U1474 (N_1474,In_670,In_1634);
xor U1475 (N_1475,In_1251,In_749);
or U1476 (N_1476,In_565,In_1970);
nand U1477 (N_1477,In_577,In_2291);
or U1478 (N_1478,In_1527,In_1837);
nand U1479 (N_1479,In_1058,In_2439);
and U1480 (N_1480,In_1054,In_1770);
or U1481 (N_1481,In_649,In_661);
or U1482 (N_1482,In_2390,In_1205);
and U1483 (N_1483,In_1845,In_1708);
or U1484 (N_1484,In_420,In_687);
nand U1485 (N_1485,In_2229,In_1298);
nor U1486 (N_1486,In_1608,In_798);
and U1487 (N_1487,In_424,In_44);
xnor U1488 (N_1488,In_513,In_669);
xnor U1489 (N_1489,In_112,In_1605);
nand U1490 (N_1490,In_348,In_443);
nor U1491 (N_1491,In_2206,In_1939);
or U1492 (N_1492,In_1511,In_816);
xor U1493 (N_1493,In_2205,In_1842);
and U1494 (N_1494,In_1572,In_803);
xnor U1495 (N_1495,In_534,In_1014);
and U1496 (N_1496,In_264,In_1690);
and U1497 (N_1497,In_21,In_2410);
or U1498 (N_1498,In_2339,In_2422);
nor U1499 (N_1499,In_2263,In_1123);
nand U1500 (N_1500,In_99,In_2027);
nand U1501 (N_1501,In_2308,In_1212);
nor U1502 (N_1502,In_95,In_805);
xnor U1503 (N_1503,In_478,In_341);
and U1504 (N_1504,In_1278,In_1838);
and U1505 (N_1505,In_2234,In_669);
and U1506 (N_1506,In_94,In_1082);
nor U1507 (N_1507,In_1686,In_820);
or U1508 (N_1508,In_297,In_2160);
nand U1509 (N_1509,In_420,In_142);
nand U1510 (N_1510,In_1801,In_972);
nor U1511 (N_1511,In_1709,In_121);
and U1512 (N_1512,In_1885,In_2045);
or U1513 (N_1513,In_998,In_491);
xor U1514 (N_1514,In_768,In_286);
nor U1515 (N_1515,In_1203,In_233);
nor U1516 (N_1516,In_681,In_1364);
or U1517 (N_1517,In_832,In_39);
and U1518 (N_1518,In_1602,In_1450);
nand U1519 (N_1519,In_2386,In_1317);
or U1520 (N_1520,In_855,In_2474);
or U1521 (N_1521,In_1966,In_1492);
and U1522 (N_1522,In_1700,In_988);
and U1523 (N_1523,In_1809,In_2059);
nor U1524 (N_1524,In_1955,In_177);
nand U1525 (N_1525,In_2176,In_1223);
nor U1526 (N_1526,In_1846,In_1330);
nor U1527 (N_1527,In_715,In_1563);
nand U1528 (N_1528,In_865,In_1072);
and U1529 (N_1529,In_321,In_2051);
or U1530 (N_1530,In_489,In_460);
nor U1531 (N_1531,In_1940,In_1211);
nand U1532 (N_1532,In_26,In_1679);
nand U1533 (N_1533,In_1936,In_2404);
or U1534 (N_1534,In_2223,In_2158);
xnor U1535 (N_1535,In_1674,In_1867);
nor U1536 (N_1536,In_1592,In_1995);
nor U1537 (N_1537,In_1355,In_2070);
nand U1538 (N_1538,In_1702,In_622);
nor U1539 (N_1539,In_1999,In_1828);
or U1540 (N_1540,In_582,In_756);
or U1541 (N_1541,In_1204,In_273);
or U1542 (N_1542,In_1384,In_1380);
nor U1543 (N_1543,In_1058,In_818);
and U1544 (N_1544,In_728,In_729);
nor U1545 (N_1545,In_432,In_589);
or U1546 (N_1546,In_388,In_357);
nand U1547 (N_1547,In_1685,In_45);
and U1548 (N_1548,In_1554,In_304);
nand U1549 (N_1549,In_55,In_97);
or U1550 (N_1550,In_1045,In_791);
nand U1551 (N_1551,In_157,In_1949);
and U1552 (N_1552,In_311,In_101);
and U1553 (N_1553,In_2446,In_2322);
nand U1554 (N_1554,In_1433,In_1083);
and U1555 (N_1555,In_1361,In_1811);
xnor U1556 (N_1556,In_1831,In_1986);
nand U1557 (N_1557,In_2430,In_1357);
nor U1558 (N_1558,In_1181,In_1821);
xor U1559 (N_1559,In_2437,In_827);
or U1560 (N_1560,In_540,In_2362);
nand U1561 (N_1561,In_1937,In_1279);
nand U1562 (N_1562,In_838,In_2328);
and U1563 (N_1563,In_1918,In_1481);
nand U1564 (N_1564,In_873,In_1845);
nor U1565 (N_1565,In_668,In_2133);
xnor U1566 (N_1566,In_2237,In_1748);
nor U1567 (N_1567,In_1850,In_2479);
and U1568 (N_1568,In_442,In_2427);
nand U1569 (N_1569,In_2187,In_1317);
or U1570 (N_1570,In_1716,In_916);
nor U1571 (N_1571,In_1404,In_440);
and U1572 (N_1572,In_2196,In_961);
nand U1573 (N_1573,In_1147,In_2408);
nor U1574 (N_1574,In_663,In_880);
nor U1575 (N_1575,In_2085,In_1003);
nand U1576 (N_1576,In_422,In_1925);
nor U1577 (N_1577,In_1410,In_1255);
or U1578 (N_1578,In_1289,In_2325);
or U1579 (N_1579,In_1098,In_34);
xor U1580 (N_1580,In_2381,In_2086);
nor U1581 (N_1581,In_1834,In_627);
nand U1582 (N_1582,In_1210,In_614);
xor U1583 (N_1583,In_1388,In_2286);
nand U1584 (N_1584,In_917,In_1073);
nor U1585 (N_1585,In_303,In_342);
nand U1586 (N_1586,In_1902,In_975);
xor U1587 (N_1587,In_2270,In_1455);
or U1588 (N_1588,In_1716,In_321);
and U1589 (N_1589,In_2176,In_1609);
nor U1590 (N_1590,In_1959,In_2484);
nor U1591 (N_1591,In_1223,In_438);
and U1592 (N_1592,In_2176,In_848);
and U1593 (N_1593,In_2122,In_1011);
xnor U1594 (N_1594,In_971,In_577);
or U1595 (N_1595,In_1815,In_270);
nand U1596 (N_1596,In_2272,In_1988);
nor U1597 (N_1597,In_1185,In_1020);
xor U1598 (N_1598,In_1401,In_439);
or U1599 (N_1599,In_1966,In_1190);
xnor U1600 (N_1600,In_1569,In_1198);
or U1601 (N_1601,In_1275,In_331);
xor U1602 (N_1602,In_851,In_694);
or U1603 (N_1603,In_2422,In_504);
and U1604 (N_1604,In_1337,In_341);
and U1605 (N_1605,In_1543,In_374);
and U1606 (N_1606,In_2438,In_427);
and U1607 (N_1607,In_1235,In_770);
or U1608 (N_1608,In_1163,In_2224);
nand U1609 (N_1609,In_2018,In_2384);
nor U1610 (N_1610,In_43,In_2198);
nor U1611 (N_1611,In_590,In_1415);
and U1612 (N_1612,In_2411,In_1686);
xnor U1613 (N_1613,In_4,In_995);
xnor U1614 (N_1614,In_1919,In_1067);
nand U1615 (N_1615,In_2191,In_473);
nand U1616 (N_1616,In_1618,In_1708);
xor U1617 (N_1617,In_236,In_1360);
xor U1618 (N_1618,In_1358,In_2389);
nand U1619 (N_1619,In_2210,In_767);
xor U1620 (N_1620,In_1456,In_2082);
nor U1621 (N_1621,In_1937,In_694);
nand U1622 (N_1622,In_1036,In_3);
xnor U1623 (N_1623,In_537,In_1244);
or U1624 (N_1624,In_1428,In_1828);
nand U1625 (N_1625,In_599,In_440);
xor U1626 (N_1626,In_743,In_775);
or U1627 (N_1627,In_864,In_913);
nor U1628 (N_1628,In_2182,In_578);
xor U1629 (N_1629,In_2276,In_2492);
and U1630 (N_1630,In_1573,In_1523);
xor U1631 (N_1631,In_1205,In_2469);
and U1632 (N_1632,In_1150,In_1593);
nand U1633 (N_1633,In_303,In_1986);
nand U1634 (N_1634,In_116,In_93);
nand U1635 (N_1635,In_1598,In_1964);
or U1636 (N_1636,In_949,In_635);
xnor U1637 (N_1637,In_549,In_1022);
nor U1638 (N_1638,In_765,In_1184);
nand U1639 (N_1639,In_1085,In_839);
and U1640 (N_1640,In_1320,In_1844);
nor U1641 (N_1641,In_1956,In_301);
or U1642 (N_1642,In_1195,In_1420);
nor U1643 (N_1643,In_1946,In_2493);
xnor U1644 (N_1644,In_371,In_2213);
nor U1645 (N_1645,In_2338,In_1979);
or U1646 (N_1646,In_787,In_1744);
xor U1647 (N_1647,In_1778,In_132);
nor U1648 (N_1648,In_2277,In_1244);
and U1649 (N_1649,In_1364,In_2487);
or U1650 (N_1650,In_1095,In_1285);
nor U1651 (N_1651,In_891,In_1695);
and U1652 (N_1652,In_1013,In_1715);
and U1653 (N_1653,In_1245,In_1294);
and U1654 (N_1654,In_375,In_2053);
or U1655 (N_1655,In_2110,In_5);
and U1656 (N_1656,In_448,In_1003);
nand U1657 (N_1657,In_561,In_552);
or U1658 (N_1658,In_1878,In_1897);
and U1659 (N_1659,In_652,In_1110);
nor U1660 (N_1660,In_2374,In_36);
nand U1661 (N_1661,In_126,In_1865);
xor U1662 (N_1662,In_671,In_1360);
nand U1663 (N_1663,In_465,In_1171);
xor U1664 (N_1664,In_400,In_35);
nor U1665 (N_1665,In_1239,In_2056);
or U1666 (N_1666,In_2277,In_1169);
xor U1667 (N_1667,In_2016,In_63);
or U1668 (N_1668,In_2483,In_992);
nor U1669 (N_1669,In_2448,In_1146);
or U1670 (N_1670,In_1427,In_742);
and U1671 (N_1671,In_826,In_1457);
or U1672 (N_1672,In_1764,In_2494);
or U1673 (N_1673,In_660,In_2393);
and U1674 (N_1674,In_561,In_393);
nand U1675 (N_1675,In_1975,In_1897);
and U1676 (N_1676,In_1063,In_364);
xnor U1677 (N_1677,In_1780,In_1546);
or U1678 (N_1678,In_871,In_1295);
xor U1679 (N_1679,In_1750,In_2108);
xor U1680 (N_1680,In_1028,In_1550);
nor U1681 (N_1681,In_1785,In_778);
or U1682 (N_1682,In_275,In_1976);
nor U1683 (N_1683,In_1211,In_453);
and U1684 (N_1684,In_1024,In_409);
or U1685 (N_1685,In_699,In_1033);
nand U1686 (N_1686,In_211,In_1768);
and U1687 (N_1687,In_1937,In_1362);
nor U1688 (N_1688,In_1980,In_537);
nand U1689 (N_1689,In_1780,In_1603);
xnor U1690 (N_1690,In_665,In_1404);
nor U1691 (N_1691,In_2477,In_1870);
nand U1692 (N_1692,In_2183,In_490);
nor U1693 (N_1693,In_671,In_2401);
nor U1694 (N_1694,In_392,In_1035);
nor U1695 (N_1695,In_1412,In_1555);
or U1696 (N_1696,In_1124,In_338);
xnor U1697 (N_1697,In_2006,In_742);
and U1698 (N_1698,In_2283,In_739);
nand U1699 (N_1699,In_667,In_79);
and U1700 (N_1700,In_2401,In_1205);
or U1701 (N_1701,In_167,In_2091);
nand U1702 (N_1702,In_635,In_163);
or U1703 (N_1703,In_2309,In_1901);
or U1704 (N_1704,In_1787,In_2243);
xor U1705 (N_1705,In_2020,In_1713);
xor U1706 (N_1706,In_674,In_1038);
and U1707 (N_1707,In_801,In_654);
nand U1708 (N_1708,In_2226,In_671);
and U1709 (N_1709,In_1855,In_1468);
nand U1710 (N_1710,In_819,In_2236);
nand U1711 (N_1711,In_1333,In_616);
or U1712 (N_1712,In_1305,In_2498);
nor U1713 (N_1713,In_698,In_1472);
nor U1714 (N_1714,In_2419,In_600);
xnor U1715 (N_1715,In_1207,In_1194);
nand U1716 (N_1716,In_1622,In_1583);
or U1717 (N_1717,In_2309,In_492);
and U1718 (N_1718,In_2047,In_702);
nand U1719 (N_1719,In_516,In_1710);
xor U1720 (N_1720,In_1346,In_1925);
or U1721 (N_1721,In_2213,In_1844);
and U1722 (N_1722,In_1458,In_2353);
xnor U1723 (N_1723,In_1180,In_184);
nand U1724 (N_1724,In_1335,In_667);
or U1725 (N_1725,In_1813,In_1507);
nand U1726 (N_1726,In_1380,In_1433);
nand U1727 (N_1727,In_2253,In_584);
and U1728 (N_1728,In_165,In_649);
xnor U1729 (N_1729,In_1182,In_1728);
nand U1730 (N_1730,In_554,In_911);
nand U1731 (N_1731,In_1829,In_2425);
and U1732 (N_1732,In_2484,In_1216);
xnor U1733 (N_1733,In_2110,In_1878);
or U1734 (N_1734,In_1998,In_2186);
xor U1735 (N_1735,In_1210,In_113);
or U1736 (N_1736,In_1638,In_1523);
nor U1737 (N_1737,In_1099,In_1055);
nor U1738 (N_1738,In_1596,In_94);
nand U1739 (N_1739,In_1237,In_1767);
and U1740 (N_1740,In_1205,In_1845);
or U1741 (N_1741,In_1155,In_1293);
nor U1742 (N_1742,In_2130,In_910);
xor U1743 (N_1743,In_37,In_900);
xor U1744 (N_1744,In_2442,In_711);
xor U1745 (N_1745,In_2178,In_1835);
nor U1746 (N_1746,In_2023,In_1794);
xor U1747 (N_1747,In_1505,In_2499);
or U1748 (N_1748,In_2494,In_1726);
or U1749 (N_1749,In_2498,In_2277);
nor U1750 (N_1750,In_822,In_834);
xor U1751 (N_1751,In_854,In_1477);
xnor U1752 (N_1752,In_1691,In_1896);
and U1753 (N_1753,In_2020,In_1788);
xor U1754 (N_1754,In_685,In_855);
xnor U1755 (N_1755,In_2040,In_1562);
or U1756 (N_1756,In_2473,In_2173);
nand U1757 (N_1757,In_830,In_820);
or U1758 (N_1758,In_2123,In_1588);
nand U1759 (N_1759,In_182,In_890);
or U1760 (N_1760,In_2143,In_2144);
or U1761 (N_1761,In_1242,In_1786);
nor U1762 (N_1762,In_1201,In_866);
xnor U1763 (N_1763,In_1577,In_2483);
xor U1764 (N_1764,In_910,In_761);
and U1765 (N_1765,In_1962,In_911);
xor U1766 (N_1766,In_866,In_2134);
nand U1767 (N_1767,In_1559,In_2066);
or U1768 (N_1768,In_1034,In_1838);
xor U1769 (N_1769,In_2411,In_112);
xor U1770 (N_1770,In_1571,In_1284);
nand U1771 (N_1771,In_112,In_961);
xnor U1772 (N_1772,In_924,In_1397);
or U1773 (N_1773,In_755,In_1020);
or U1774 (N_1774,In_1432,In_1992);
and U1775 (N_1775,In_358,In_2384);
and U1776 (N_1776,In_844,In_1415);
and U1777 (N_1777,In_1315,In_265);
nand U1778 (N_1778,In_1196,In_2341);
nand U1779 (N_1779,In_948,In_1265);
nand U1780 (N_1780,In_2183,In_2263);
nand U1781 (N_1781,In_2443,In_1239);
xor U1782 (N_1782,In_1226,In_2391);
nor U1783 (N_1783,In_2009,In_408);
or U1784 (N_1784,In_2291,In_843);
xor U1785 (N_1785,In_2091,In_1315);
xor U1786 (N_1786,In_1245,In_92);
nand U1787 (N_1787,In_390,In_2434);
or U1788 (N_1788,In_235,In_1707);
xor U1789 (N_1789,In_1873,In_1976);
xor U1790 (N_1790,In_672,In_1949);
or U1791 (N_1791,In_797,In_1274);
or U1792 (N_1792,In_1397,In_1510);
nor U1793 (N_1793,In_1400,In_859);
and U1794 (N_1794,In_1716,In_2072);
nor U1795 (N_1795,In_1565,In_1097);
nand U1796 (N_1796,In_1702,In_1274);
and U1797 (N_1797,In_108,In_742);
or U1798 (N_1798,In_1934,In_2357);
nand U1799 (N_1799,In_1818,In_709);
and U1800 (N_1800,In_276,In_2360);
or U1801 (N_1801,In_713,In_1086);
or U1802 (N_1802,In_1131,In_1561);
nand U1803 (N_1803,In_2060,In_902);
xnor U1804 (N_1804,In_419,In_2498);
and U1805 (N_1805,In_930,In_1339);
xor U1806 (N_1806,In_1593,In_1174);
nor U1807 (N_1807,In_909,In_46);
nor U1808 (N_1808,In_208,In_452);
nand U1809 (N_1809,In_1955,In_1624);
xor U1810 (N_1810,In_230,In_207);
nor U1811 (N_1811,In_2414,In_1877);
and U1812 (N_1812,In_1830,In_420);
nor U1813 (N_1813,In_2318,In_1289);
xnor U1814 (N_1814,In_844,In_691);
nand U1815 (N_1815,In_232,In_1355);
and U1816 (N_1816,In_2393,In_1152);
xnor U1817 (N_1817,In_2004,In_1932);
and U1818 (N_1818,In_528,In_1582);
and U1819 (N_1819,In_112,In_1611);
and U1820 (N_1820,In_942,In_1037);
and U1821 (N_1821,In_1089,In_593);
and U1822 (N_1822,In_1683,In_2128);
or U1823 (N_1823,In_1074,In_2283);
nor U1824 (N_1824,In_1595,In_2050);
or U1825 (N_1825,In_777,In_942);
and U1826 (N_1826,In_2207,In_153);
nor U1827 (N_1827,In_621,In_1462);
or U1828 (N_1828,In_35,In_733);
nand U1829 (N_1829,In_2293,In_280);
or U1830 (N_1830,In_2217,In_1881);
or U1831 (N_1831,In_369,In_289);
nor U1832 (N_1832,In_1638,In_953);
nand U1833 (N_1833,In_1462,In_2355);
nand U1834 (N_1834,In_2192,In_404);
and U1835 (N_1835,In_1620,In_2238);
and U1836 (N_1836,In_274,In_568);
nor U1837 (N_1837,In_798,In_667);
or U1838 (N_1838,In_1740,In_577);
and U1839 (N_1839,In_210,In_1379);
or U1840 (N_1840,In_1594,In_928);
nor U1841 (N_1841,In_1842,In_2061);
nor U1842 (N_1842,In_2167,In_666);
nor U1843 (N_1843,In_28,In_2198);
nand U1844 (N_1844,In_2405,In_598);
xnor U1845 (N_1845,In_412,In_289);
and U1846 (N_1846,In_48,In_729);
or U1847 (N_1847,In_618,In_1833);
or U1848 (N_1848,In_1229,In_2116);
nand U1849 (N_1849,In_846,In_1742);
or U1850 (N_1850,In_751,In_220);
xnor U1851 (N_1851,In_650,In_631);
nand U1852 (N_1852,In_2353,In_1535);
nor U1853 (N_1853,In_1502,In_1633);
and U1854 (N_1854,In_2304,In_991);
and U1855 (N_1855,In_1484,In_519);
nand U1856 (N_1856,In_1326,In_416);
nand U1857 (N_1857,In_2294,In_1497);
and U1858 (N_1858,In_2105,In_1308);
and U1859 (N_1859,In_1885,In_15);
nand U1860 (N_1860,In_1903,In_1658);
xnor U1861 (N_1861,In_1140,In_2214);
xnor U1862 (N_1862,In_193,In_696);
nor U1863 (N_1863,In_414,In_1118);
xnor U1864 (N_1864,In_1924,In_1926);
nand U1865 (N_1865,In_2482,In_1521);
or U1866 (N_1866,In_1374,In_1530);
or U1867 (N_1867,In_1978,In_752);
xnor U1868 (N_1868,In_1534,In_1664);
nor U1869 (N_1869,In_647,In_729);
nor U1870 (N_1870,In_533,In_880);
or U1871 (N_1871,In_766,In_1608);
nor U1872 (N_1872,In_939,In_1486);
and U1873 (N_1873,In_50,In_1179);
xor U1874 (N_1874,In_1584,In_1267);
and U1875 (N_1875,In_764,In_2324);
xor U1876 (N_1876,In_2176,In_1874);
or U1877 (N_1877,In_500,In_1026);
xnor U1878 (N_1878,In_2478,In_2479);
nor U1879 (N_1879,In_2382,In_933);
and U1880 (N_1880,In_919,In_1761);
or U1881 (N_1881,In_1953,In_148);
or U1882 (N_1882,In_253,In_2020);
nand U1883 (N_1883,In_1840,In_249);
xnor U1884 (N_1884,In_2139,In_1394);
or U1885 (N_1885,In_1259,In_883);
xor U1886 (N_1886,In_26,In_2027);
and U1887 (N_1887,In_623,In_696);
nand U1888 (N_1888,In_2351,In_1738);
nand U1889 (N_1889,In_1630,In_1621);
nor U1890 (N_1890,In_1187,In_2255);
nor U1891 (N_1891,In_810,In_1937);
or U1892 (N_1892,In_741,In_297);
nor U1893 (N_1893,In_1855,In_477);
or U1894 (N_1894,In_759,In_818);
or U1895 (N_1895,In_1407,In_2388);
and U1896 (N_1896,In_18,In_112);
and U1897 (N_1897,In_1378,In_1404);
xor U1898 (N_1898,In_871,In_1461);
nand U1899 (N_1899,In_224,In_1464);
nand U1900 (N_1900,In_2066,In_348);
nand U1901 (N_1901,In_2196,In_315);
nand U1902 (N_1902,In_2467,In_366);
and U1903 (N_1903,In_1620,In_2242);
nor U1904 (N_1904,In_1027,In_1070);
and U1905 (N_1905,In_2234,In_816);
nand U1906 (N_1906,In_2198,In_392);
nor U1907 (N_1907,In_1958,In_1662);
or U1908 (N_1908,In_2087,In_2454);
or U1909 (N_1909,In_946,In_2272);
and U1910 (N_1910,In_1027,In_2338);
xnor U1911 (N_1911,In_1657,In_1487);
nor U1912 (N_1912,In_304,In_2081);
nand U1913 (N_1913,In_425,In_1573);
xnor U1914 (N_1914,In_427,In_1970);
nand U1915 (N_1915,In_2155,In_1384);
nand U1916 (N_1916,In_1581,In_567);
or U1917 (N_1917,In_2323,In_144);
and U1918 (N_1918,In_974,In_1071);
or U1919 (N_1919,In_1909,In_1352);
and U1920 (N_1920,In_259,In_367);
and U1921 (N_1921,In_599,In_2121);
or U1922 (N_1922,In_1025,In_2446);
nor U1923 (N_1923,In_885,In_1822);
and U1924 (N_1924,In_576,In_1089);
or U1925 (N_1925,In_2252,In_74);
xnor U1926 (N_1926,In_1270,In_648);
xor U1927 (N_1927,In_2063,In_176);
nor U1928 (N_1928,In_1483,In_1246);
or U1929 (N_1929,In_980,In_2218);
nor U1930 (N_1930,In_732,In_936);
nor U1931 (N_1931,In_1030,In_2063);
nand U1932 (N_1932,In_1645,In_322);
or U1933 (N_1933,In_135,In_1606);
xor U1934 (N_1934,In_2229,In_342);
or U1935 (N_1935,In_773,In_1316);
nor U1936 (N_1936,In_998,In_1875);
xor U1937 (N_1937,In_783,In_1053);
xor U1938 (N_1938,In_1037,In_1698);
and U1939 (N_1939,In_927,In_2316);
xnor U1940 (N_1940,In_2347,In_1354);
nand U1941 (N_1941,In_1984,In_1398);
xnor U1942 (N_1942,In_949,In_1180);
and U1943 (N_1943,In_2003,In_2048);
or U1944 (N_1944,In_2303,In_1530);
xor U1945 (N_1945,In_734,In_323);
nor U1946 (N_1946,In_1440,In_1843);
or U1947 (N_1947,In_956,In_382);
nand U1948 (N_1948,In_1544,In_297);
nor U1949 (N_1949,In_1721,In_118);
and U1950 (N_1950,In_1689,In_530);
nor U1951 (N_1951,In_2497,In_531);
nor U1952 (N_1952,In_1419,In_1105);
and U1953 (N_1953,In_1711,In_589);
xnor U1954 (N_1954,In_524,In_286);
xnor U1955 (N_1955,In_1517,In_2391);
or U1956 (N_1956,In_2349,In_1475);
and U1957 (N_1957,In_494,In_2153);
xor U1958 (N_1958,In_2135,In_850);
and U1959 (N_1959,In_2139,In_1425);
nand U1960 (N_1960,In_448,In_1596);
nand U1961 (N_1961,In_698,In_2192);
xnor U1962 (N_1962,In_346,In_1133);
and U1963 (N_1963,In_2250,In_2175);
nand U1964 (N_1964,In_510,In_2256);
nor U1965 (N_1965,In_9,In_2200);
nand U1966 (N_1966,In_732,In_455);
and U1967 (N_1967,In_2458,In_1687);
nand U1968 (N_1968,In_427,In_1622);
or U1969 (N_1969,In_2358,In_227);
and U1970 (N_1970,In_1334,In_397);
nor U1971 (N_1971,In_1711,In_1262);
nand U1972 (N_1972,In_998,In_254);
xnor U1973 (N_1973,In_685,In_885);
or U1974 (N_1974,In_2057,In_2471);
nand U1975 (N_1975,In_1161,In_322);
xnor U1976 (N_1976,In_1248,In_1383);
or U1977 (N_1977,In_1568,In_946);
and U1978 (N_1978,In_134,In_1281);
xnor U1979 (N_1979,In_302,In_1908);
nand U1980 (N_1980,In_190,In_2184);
nor U1981 (N_1981,In_2163,In_1610);
nand U1982 (N_1982,In_995,In_1834);
nor U1983 (N_1983,In_1337,In_1964);
xor U1984 (N_1984,In_692,In_973);
or U1985 (N_1985,In_1238,In_1197);
xnor U1986 (N_1986,In_574,In_1242);
or U1987 (N_1987,In_133,In_630);
and U1988 (N_1988,In_1837,In_1277);
or U1989 (N_1989,In_2256,In_2413);
and U1990 (N_1990,In_289,In_2115);
and U1991 (N_1991,In_861,In_1971);
or U1992 (N_1992,In_165,In_201);
xnor U1993 (N_1993,In_711,In_748);
and U1994 (N_1994,In_438,In_1364);
nor U1995 (N_1995,In_2491,In_1487);
and U1996 (N_1996,In_248,In_50);
nand U1997 (N_1997,In_62,In_2246);
xnor U1998 (N_1998,In_1206,In_1819);
nor U1999 (N_1999,In_2168,In_2067);
or U2000 (N_2000,In_1,In_2482);
nand U2001 (N_2001,In_2498,In_998);
and U2002 (N_2002,In_106,In_1120);
nor U2003 (N_2003,In_651,In_2222);
nor U2004 (N_2004,In_1844,In_1036);
nand U2005 (N_2005,In_774,In_819);
or U2006 (N_2006,In_2264,In_1440);
nand U2007 (N_2007,In_2120,In_776);
nand U2008 (N_2008,In_1775,In_2022);
nand U2009 (N_2009,In_2379,In_171);
and U2010 (N_2010,In_2400,In_437);
xor U2011 (N_2011,In_11,In_1060);
nor U2012 (N_2012,In_562,In_692);
xnor U2013 (N_2013,In_1993,In_1803);
and U2014 (N_2014,In_2246,In_2146);
xnor U2015 (N_2015,In_1852,In_1293);
xnor U2016 (N_2016,In_459,In_2091);
xor U2017 (N_2017,In_339,In_243);
nor U2018 (N_2018,In_1295,In_1023);
or U2019 (N_2019,In_1630,In_586);
and U2020 (N_2020,In_2333,In_2210);
xor U2021 (N_2021,In_2162,In_1440);
nand U2022 (N_2022,In_1416,In_267);
xnor U2023 (N_2023,In_1185,In_1986);
xnor U2024 (N_2024,In_841,In_1412);
xor U2025 (N_2025,In_2261,In_1232);
and U2026 (N_2026,In_2487,In_909);
nor U2027 (N_2027,In_2070,In_1063);
nand U2028 (N_2028,In_1868,In_418);
xor U2029 (N_2029,In_1239,In_1920);
xor U2030 (N_2030,In_736,In_2380);
nor U2031 (N_2031,In_1336,In_1526);
xor U2032 (N_2032,In_446,In_2227);
and U2033 (N_2033,In_532,In_1056);
nand U2034 (N_2034,In_27,In_318);
xnor U2035 (N_2035,In_1445,In_1660);
or U2036 (N_2036,In_886,In_1383);
and U2037 (N_2037,In_2308,In_541);
nand U2038 (N_2038,In_1551,In_660);
nand U2039 (N_2039,In_1531,In_889);
or U2040 (N_2040,In_996,In_2432);
and U2041 (N_2041,In_387,In_2351);
xor U2042 (N_2042,In_769,In_1554);
xnor U2043 (N_2043,In_738,In_4);
and U2044 (N_2044,In_1032,In_1387);
and U2045 (N_2045,In_1602,In_687);
or U2046 (N_2046,In_2385,In_884);
nor U2047 (N_2047,In_2206,In_1287);
xnor U2048 (N_2048,In_493,In_1057);
nor U2049 (N_2049,In_94,In_1856);
xnor U2050 (N_2050,In_1547,In_1282);
xor U2051 (N_2051,In_76,In_445);
nor U2052 (N_2052,In_1818,In_2175);
xor U2053 (N_2053,In_1977,In_2297);
and U2054 (N_2054,In_2333,In_716);
nor U2055 (N_2055,In_847,In_2250);
nor U2056 (N_2056,In_1180,In_1719);
and U2057 (N_2057,In_621,In_709);
xnor U2058 (N_2058,In_922,In_856);
xor U2059 (N_2059,In_1541,In_880);
xnor U2060 (N_2060,In_1082,In_249);
nand U2061 (N_2061,In_879,In_2083);
nand U2062 (N_2062,In_553,In_87);
and U2063 (N_2063,In_1237,In_1545);
xor U2064 (N_2064,In_2252,In_1913);
nand U2065 (N_2065,In_2118,In_1585);
nand U2066 (N_2066,In_1695,In_1356);
or U2067 (N_2067,In_1655,In_2439);
or U2068 (N_2068,In_113,In_1541);
and U2069 (N_2069,In_1267,In_2430);
xor U2070 (N_2070,In_1501,In_1228);
nand U2071 (N_2071,In_435,In_1842);
nor U2072 (N_2072,In_703,In_2278);
and U2073 (N_2073,In_498,In_2332);
xor U2074 (N_2074,In_160,In_783);
xnor U2075 (N_2075,In_298,In_2150);
nand U2076 (N_2076,In_1055,In_2347);
nor U2077 (N_2077,In_2466,In_1761);
or U2078 (N_2078,In_934,In_2081);
and U2079 (N_2079,In_1754,In_78);
nand U2080 (N_2080,In_2282,In_185);
xor U2081 (N_2081,In_1169,In_1585);
xnor U2082 (N_2082,In_389,In_2179);
and U2083 (N_2083,In_496,In_1901);
xnor U2084 (N_2084,In_1577,In_1551);
nand U2085 (N_2085,In_1532,In_2117);
or U2086 (N_2086,In_250,In_713);
xor U2087 (N_2087,In_1979,In_1389);
or U2088 (N_2088,In_1120,In_223);
or U2089 (N_2089,In_1989,In_1392);
nor U2090 (N_2090,In_2014,In_1421);
xor U2091 (N_2091,In_319,In_2456);
and U2092 (N_2092,In_2392,In_1983);
nor U2093 (N_2093,In_2245,In_991);
or U2094 (N_2094,In_311,In_539);
nand U2095 (N_2095,In_1438,In_1644);
xnor U2096 (N_2096,In_47,In_215);
or U2097 (N_2097,In_2317,In_2247);
nand U2098 (N_2098,In_976,In_167);
and U2099 (N_2099,In_392,In_1871);
or U2100 (N_2100,In_37,In_1450);
xnor U2101 (N_2101,In_357,In_2223);
nor U2102 (N_2102,In_2080,In_64);
or U2103 (N_2103,In_2490,In_569);
and U2104 (N_2104,In_1069,In_1638);
or U2105 (N_2105,In_1603,In_800);
xnor U2106 (N_2106,In_63,In_587);
or U2107 (N_2107,In_66,In_2195);
and U2108 (N_2108,In_1438,In_1838);
nand U2109 (N_2109,In_975,In_1435);
and U2110 (N_2110,In_2343,In_1658);
nor U2111 (N_2111,In_2116,In_1738);
xor U2112 (N_2112,In_1878,In_910);
nor U2113 (N_2113,In_164,In_407);
nand U2114 (N_2114,In_946,In_1419);
nand U2115 (N_2115,In_141,In_1389);
or U2116 (N_2116,In_3,In_2425);
or U2117 (N_2117,In_950,In_1489);
nor U2118 (N_2118,In_338,In_1742);
nor U2119 (N_2119,In_1827,In_1822);
xnor U2120 (N_2120,In_2433,In_1030);
nand U2121 (N_2121,In_2381,In_1479);
and U2122 (N_2122,In_1200,In_34);
and U2123 (N_2123,In_789,In_704);
nand U2124 (N_2124,In_2161,In_638);
nor U2125 (N_2125,In_1661,In_1036);
or U2126 (N_2126,In_1233,In_1162);
nand U2127 (N_2127,In_689,In_1976);
or U2128 (N_2128,In_2406,In_128);
nor U2129 (N_2129,In_1084,In_2079);
nor U2130 (N_2130,In_2121,In_316);
nand U2131 (N_2131,In_1238,In_315);
and U2132 (N_2132,In_2496,In_2057);
nor U2133 (N_2133,In_1872,In_2256);
nor U2134 (N_2134,In_2433,In_1528);
or U2135 (N_2135,In_111,In_386);
and U2136 (N_2136,In_535,In_1785);
or U2137 (N_2137,In_1180,In_758);
nor U2138 (N_2138,In_2188,In_243);
or U2139 (N_2139,In_1347,In_1205);
xnor U2140 (N_2140,In_1693,In_1024);
or U2141 (N_2141,In_174,In_158);
nand U2142 (N_2142,In_1569,In_1674);
and U2143 (N_2143,In_1414,In_1667);
xor U2144 (N_2144,In_1778,In_1682);
and U2145 (N_2145,In_899,In_42);
xnor U2146 (N_2146,In_2172,In_1765);
nor U2147 (N_2147,In_2484,In_203);
xnor U2148 (N_2148,In_578,In_1493);
nor U2149 (N_2149,In_2221,In_1995);
and U2150 (N_2150,In_1155,In_1913);
and U2151 (N_2151,In_169,In_2250);
nor U2152 (N_2152,In_582,In_466);
xor U2153 (N_2153,In_287,In_1522);
nand U2154 (N_2154,In_1646,In_675);
or U2155 (N_2155,In_573,In_1333);
and U2156 (N_2156,In_810,In_194);
nand U2157 (N_2157,In_204,In_413);
or U2158 (N_2158,In_415,In_224);
and U2159 (N_2159,In_356,In_927);
and U2160 (N_2160,In_1441,In_804);
xor U2161 (N_2161,In_1803,In_831);
or U2162 (N_2162,In_2406,In_1346);
and U2163 (N_2163,In_1704,In_2041);
xnor U2164 (N_2164,In_771,In_1852);
and U2165 (N_2165,In_1687,In_2478);
or U2166 (N_2166,In_661,In_2019);
nand U2167 (N_2167,In_1909,In_2339);
and U2168 (N_2168,In_948,In_826);
nor U2169 (N_2169,In_902,In_1572);
xnor U2170 (N_2170,In_1547,In_1266);
nand U2171 (N_2171,In_1754,In_1951);
and U2172 (N_2172,In_1077,In_2072);
nand U2173 (N_2173,In_1464,In_2138);
or U2174 (N_2174,In_753,In_34);
xor U2175 (N_2175,In_565,In_1907);
nor U2176 (N_2176,In_290,In_1760);
nand U2177 (N_2177,In_2,In_1012);
xor U2178 (N_2178,In_2381,In_628);
or U2179 (N_2179,In_309,In_1857);
nor U2180 (N_2180,In_1396,In_1890);
xor U2181 (N_2181,In_869,In_1057);
nand U2182 (N_2182,In_2025,In_1505);
nand U2183 (N_2183,In_1389,In_2374);
or U2184 (N_2184,In_1014,In_676);
or U2185 (N_2185,In_703,In_1640);
or U2186 (N_2186,In_2227,In_1180);
nand U2187 (N_2187,In_1374,In_496);
and U2188 (N_2188,In_1968,In_517);
and U2189 (N_2189,In_2162,In_2264);
xor U2190 (N_2190,In_1184,In_1682);
xnor U2191 (N_2191,In_1317,In_2216);
and U2192 (N_2192,In_1379,In_320);
nand U2193 (N_2193,In_1767,In_498);
and U2194 (N_2194,In_1252,In_1313);
or U2195 (N_2195,In_321,In_161);
xnor U2196 (N_2196,In_890,In_1536);
nand U2197 (N_2197,In_1875,In_239);
and U2198 (N_2198,In_384,In_1924);
nand U2199 (N_2199,In_1822,In_521);
nand U2200 (N_2200,In_910,In_792);
and U2201 (N_2201,In_336,In_1646);
or U2202 (N_2202,In_1895,In_1946);
nand U2203 (N_2203,In_2035,In_97);
or U2204 (N_2204,In_492,In_1991);
and U2205 (N_2205,In_731,In_1310);
xnor U2206 (N_2206,In_742,In_1134);
and U2207 (N_2207,In_481,In_1295);
and U2208 (N_2208,In_1858,In_2157);
or U2209 (N_2209,In_1679,In_1022);
nor U2210 (N_2210,In_1938,In_553);
or U2211 (N_2211,In_307,In_1102);
xor U2212 (N_2212,In_2191,In_423);
xnor U2213 (N_2213,In_2233,In_2267);
xor U2214 (N_2214,In_1174,In_363);
or U2215 (N_2215,In_287,In_1150);
or U2216 (N_2216,In_2350,In_685);
nand U2217 (N_2217,In_1474,In_668);
nand U2218 (N_2218,In_1112,In_1864);
nand U2219 (N_2219,In_1728,In_785);
and U2220 (N_2220,In_147,In_2393);
and U2221 (N_2221,In_870,In_1708);
nor U2222 (N_2222,In_370,In_812);
nor U2223 (N_2223,In_992,In_1649);
nand U2224 (N_2224,In_797,In_1911);
nor U2225 (N_2225,In_1352,In_1800);
and U2226 (N_2226,In_1189,In_1029);
nor U2227 (N_2227,In_1249,In_1617);
and U2228 (N_2228,In_531,In_341);
nor U2229 (N_2229,In_1889,In_1609);
nand U2230 (N_2230,In_1633,In_851);
nand U2231 (N_2231,In_228,In_2415);
or U2232 (N_2232,In_7,In_1024);
xor U2233 (N_2233,In_1322,In_2365);
and U2234 (N_2234,In_382,In_2481);
xnor U2235 (N_2235,In_218,In_2309);
nand U2236 (N_2236,In_215,In_1750);
nand U2237 (N_2237,In_238,In_404);
xnor U2238 (N_2238,In_64,In_2350);
or U2239 (N_2239,In_1688,In_1012);
nor U2240 (N_2240,In_1039,In_1796);
xnor U2241 (N_2241,In_925,In_815);
or U2242 (N_2242,In_1868,In_503);
or U2243 (N_2243,In_1803,In_2453);
nor U2244 (N_2244,In_306,In_1902);
nor U2245 (N_2245,In_1405,In_1756);
and U2246 (N_2246,In_610,In_428);
xor U2247 (N_2247,In_2283,In_248);
nand U2248 (N_2248,In_1742,In_1075);
or U2249 (N_2249,In_2087,In_1311);
xnor U2250 (N_2250,In_600,In_1772);
or U2251 (N_2251,In_1019,In_843);
nor U2252 (N_2252,In_1216,In_672);
nor U2253 (N_2253,In_1638,In_2256);
and U2254 (N_2254,In_301,In_1576);
or U2255 (N_2255,In_2197,In_497);
nand U2256 (N_2256,In_1527,In_1587);
xnor U2257 (N_2257,In_2275,In_598);
and U2258 (N_2258,In_616,In_286);
xnor U2259 (N_2259,In_1247,In_70);
xor U2260 (N_2260,In_918,In_929);
and U2261 (N_2261,In_551,In_462);
xor U2262 (N_2262,In_1252,In_156);
nor U2263 (N_2263,In_1173,In_638);
nor U2264 (N_2264,In_1098,In_1683);
nor U2265 (N_2265,In_12,In_1456);
xnor U2266 (N_2266,In_1251,In_1423);
and U2267 (N_2267,In_1532,In_2221);
nand U2268 (N_2268,In_512,In_588);
nand U2269 (N_2269,In_1226,In_1276);
or U2270 (N_2270,In_1766,In_2374);
nor U2271 (N_2271,In_1122,In_132);
nand U2272 (N_2272,In_270,In_831);
nand U2273 (N_2273,In_384,In_1409);
or U2274 (N_2274,In_1018,In_351);
or U2275 (N_2275,In_2469,In_141);
and U2276 (N_2276,In_247,In_424);
nand U2277 (N_2277,In_94,In_1196);
nor U2278 (N_2278,In_1680,In_2213);
nor U2279 (N_2279,In_2462,In_1590);
xor U2280 (N_2280,In_147,In_2228);
nor U2281 (N_2281,In_1746,In_906);
nor U2282 (N_2282,In_2152,In_1324);
xor U2283 (N_2283,In_1288,In_2257);
and U2284 (N_2284,In_974,In_1937);
xor U2285 (N_2285,In_1867,In_1447);
nor U2286 (N_2286,In_177,In_2134);
nor U2287 (N_2287,In_1989,In_328);
or U2288 (N_2288,In_801,In_202);
nand U2289 (N_2289,In_2225,In_2128);
or U2290 (N_2290,In_401,In_765);
xnor U2291 (N_2291,In_315,In_1976);
nand U2292 (N_2292,In_1312,In_2049);
and U2293 (N_2293,In_1529,In_1893);
nor U2294 (N_2294,In_295,In_1089);
or U2295 (N_2295,In_1387,In_990);
or U2296 (N_2296,In_1023,In_2021);
xor U2297 (N_2297,In_2187,In_351);
nand U2298 (N_2298,In_19,In_679);
xor U2299 (N_2299,In_1232,In_1117);
nand U2300 (N_2300,In_531,In_1270);
xnor U2301 (N_2301,In_2080,In_710);
and U2302 (N_2302,In_1237,In_2239);
or U2303 (N_2303,In_1578,In_2043);
and U2304 (N_2304,In_2248,In_1842);
nor U2305 (N_2305,In_782,In_2209);
and U2306 (N_2306,In_2259,In_2328);
nor U2307 (N_2307,In_1598,In_2446);
and U2308 (N_2308,In_2199,In_1798);
xnor U2309 (N_2309,In_637,In_128);
and U2310 (N_2310,In_2406,In_1062);
xor U2311 (N_2311,In_311,In_1918);
nor U2312 (N_2312,In_1762,In_94);
xnor U2313 (N_2313,In_2303,In_2141);
nor U2314 (N_2314,In_2456,In_2012);
nor U2315 (N_2315,In_2273,In_850);
xor U2316 (N_2316,In_1139,In_281);
nor U2317 (N_2317,In_331,In_534);
and U2318 (N_2318,In_2211,In_2103);
and U2319 (N_2319,In_2433,In_924);
nand U2320 (N_2320,In_2265,In_958);
or U2321 (N_2321,In_2039,In_624);
xnor U2322 (N_2322,In_2126,In_1646);
and U2323 (N_2323,In_231,In_870);
xnor U2324 (N_2324,In_392,In_816);
nor U2325 (N_2325,In_468,In_1742);
and U2326 (N_2326,In_739,In_906);
xor U2327 (N_2327,In_1647,In_133);
nand U2328 (N_2328,In_562,In_119);
nor U2329 (N_2329,In_2478,In_529);
or U2330 (N_2330,In_1006,In_1392);
or U2331 (N_2331,In_103,In_2459);
nand U2332 (N_2332,In_1398,In_610);
nor U2333 (N_2333,In_1914,In_493);
nand U2334 (N_2334,In_2164,In_1603);
xor U2335 (N_2335,In_1772,In_984);
nor U2336 (N_2336,In_1860,In_1052);
nor U2337 (N_2337,In_916,In_1560);
and U2338 (N_2338,In_1590,In_913);
or U2339 (N_2339,In_1962,In_1339);
or U2340 (N_2340,In_974,In_2443);
xnor U2341 (N_2341,In_1954,In_527);
and U2342 (N_2342,In_1397,In_2054);
nor U2343 (N_2343,In_1092,In_1437);
nor U2344 (N_2344,In_726,In_1499);
xor U2345 (N_2345,In_510,In_1281);
nand U2346 (N_2346,In_1559,In_1006);
xor U2347 (N_2347,In_1259,In_777);
nand U2348 (N_2348,In_870,In_839);
nor U2349 (N_2349,In_175,In_1587);
nor U2350 (N_2350,In_2134,In_2140);
or U2351 (N_2351,In_1992,In_641);
nand U2352 (N_2352,In_1308,In_1855);
and U2353 (N_2353,In_1861,In_1654);
nor U2354 (N_2354,In_1382,In_3);
and U2355 (N_2355,In_1495,In_1428);
and U2356 (N_2356,In_1975,In_144);
or U2357 (N_2357,In_1000,In_1346);
xnor U2358 (N_2358,In_903,In_2200);
nor U2359 (N_2359,In_2092,In_2365);
nand U2360 (N_2360,In_211,In_1312);
and U2361 (N_2361,In_164,In_1920);
or U2362 (N_2362,In_340,In_316);
or U2363 (N_2363,In_1696,In_1215);
and U2364 (N_2364,In_2094,In_1311);
or U2365 (N_2365,In_1095,In_606);
nand U2366 (N_2366,In_1688,In_2463);
or U2367 (N_2367,In_961,In_926);
nand U2368 (N_2368,In_336,In_1506);
xor U2369 (N_2369,In_1182,In_1546);
or U2370 (N_2370,In_794,In_1520);
xor U2371 (N_2371,In_149,In_1913);
nand U2372 (N_2372,In_1128,In_170);
nor U2373 (N_2373,In_1196,In_182);
nor U2374 (N_2374,In_2486,In_569);
nor U2375 (N_2375,In_1959,In_1865);
nor U2376 (N_2376,In_1183,In_2483);
nor U2377 (N_2377,In_1053,In_2091);
or U2378 (N_2378,In_549,In_210);
and U2379 (N_2379,In_1479,In_1741);
and U2380 (N_2380,In_539,In_1234);
xnor U2381 (N_2381,In_623,In_2483);
xor U2382 (N_2382,In_186,In_1932);
or U2383 (N_2383,In_1704,In_556);
and U2384 (N_2384,In_1422,In_191);
nand U2385 (N_2385,In_2354,In_1106);
nor U2386 (N_2386,In_2096,In_586);
nand U2387 (N_2387,In_1763,In_787);
xor U2388 (N_2388,In_2070,In_2157);
nor U2389 (N_2389,In_1075,In_1366);
and U2390 (N_2390,In_1189,In_362);
or U2391 (N_2391,In_2330,In_2282);
nand U2392 (N_2392,In_920,In_1417);
and U2393 (N_2393,In_95,In_1530);
or U2394 (N_2394,In_436,In_1770);
and U2395 (N_2395,In_396,In_126);
nand U2396 (N_2396,In_1467,In_2124);
and U2397 (N_2397,In_505,In_2001);
nand U2398 (N_2398,In_960,In_2469);
nand U2399 (N_2399,In_229,In_688);
or U2400 (N_2400,In_1586,In_2473);
nor U2401 (N_2401,In_831,In_2202);
xor U2402 (N_2402,In_940,In_513);
nor U2403 (N_2403,In_2186,In_941);
and U2404 (N_2404,In_665,In_1354);
or U2405 (N_2405,In_1135,In_2425);
and U2406 (N_2406,In_1280,In_483);
or U2407 (N_2407,In_1722,In_1063);
and U2408 (N_2408,In_127,In_137);
xnor U2409 (N_2409,In_418,In_2056);
or U2410 (N_2410,In_486,In_1126);
nor U2411 (N_2411,In_2167,In_1966);
nand U2412 (N_2412,In_1882,In_39);
xor U2413 (N_2413,In_642,In_1);
and U2414 (N_2414,In_1773,In_1465);
or U2415 (N_2415,In_1004,In_1279);
xnor U2416 (N_2416,In_2011,In_1135);
xnor U2417 (N_2417,In_170,In_641);
nand U2418 (N_2418,In_1841,In_247);
nand U2419 (N_2419,In_2056,In_1659);
xor U2420 (N_2420,In_2243,In_2032);
xor U2421 (N_2421,In_218,In_375);
or U2422 (N_2422,In_1593,In_2447);
xnor U2423 (N_2423,In_827,In_309);
xor U2424 (N_2424,In_962,In_414);
xor U2425 (N_2425,In_1965,In_461);
or U2426 (N_2426,In_1413,In_2414);
nor U2427 (N_2427,In_2445,In_1506);
and U2428 (N_2428,In_1082,In_43);
nand U2429 (N_2429,In_307,In_2431);
and U2430 (N_2430,In_33,In_1215);
nor U2431 (N_2431,In_69,In_836);
nand U2432 (N_2432,In_1501,In_2012);
nand U2433 (N_2433,In_130,In_1469);
nor U2434 (N_2434,In_493,In_2307);
nand U2435 (N_2435,In_12,In_2216);
nor U2436 (N_2436,In_916,In_1818);
nor U2437 (N_2437,In_2410,In_1252);
nor U2438 (N_2438,In_963,In_1098);
or U2439 (N_2439,In_67,In_765);
and U2440 (N_2440,In_372,In_2362);
and U2441 (N_2441,In_1701,In_565);
nor U2442 (N_2442,In_637,In_1244);
nand U2443 (N_2443,In_2247,In_381);
xor U2444 (N_2444,In_875,In_2410);
nand U2445 (N_2445,In_2483,In_305);
nor U2446 (N_2446,In_1889,In_105);
nor U2447 (N_2447,In_2116,In_2282);
or U2448 (N_2448,In_445,In_2188);
xor U2449 (N_2449,In_1721,In_1180);
nor U2450 (N_2450,In_478,In_346);
xnor U2451 (N_2451,In_2025,In_317);
or U2452 (N_2452,In_1972,In_314);
nand U2453 (N_2453,In_1865,In_1638);
nor U2454 (N_2454,In_2208,In_1477);
nand U2455 (N_2455,In_345,In_942);
nor U2456 (N_2456,In_1287,In_2004);
or U2457 (N_2457,In_1765,In_194);
and U2458 (N_2458,In_2102,In_776);
xor U2459 (N_2459,In_2238,In_312);
and U2460 (N_2460,In_1147,In_2416);
and U2461 (N_2461,In_1621,In_322);
or U2462 (N_2462,In_648,In_2467);
nor U2463 (N_2463,In_1141,In_2237);
nor U2464 (N_2464,In_1744,In_882);
and U2465 (N_2465,In_1800,In_204);
or U2466 (N_2466,In_1889,In_1934);
nand U2467 (N_2467,In_1715,In_444);
nand U2468 (N_2468,In_2252,In_181);
nand U2469 (N_2469,In_1595,In_1627);
or U2470 (N_2470,In_1567,In_846);
and U2471 (N_2471,In_1138,In_1782);
or U2472 (N_2472,In_1428,In_1729);
xor U2473 (N_2473,In_2452,In_1773);
xnor U2474 (N_2474,In_235,In_1575);
or U2475 (N_2475,In_1190,In_2373);
and U2476 (N_2476,In_597,In_1978);
nand U2477 (N_2477,In_1213,In_2197);
and U2478 (N_2478,In_1024,In_921);
nand U2479 (N_2479,In_1116,In_1443);
nand U2480 (N_2480,In_1811,In_215);
nand U2481 (N_2481,In_41,In_1615);
or U2482 (N_2482,In_855,In_1764);
or U2483 (N_2483,In_2377,In_1177);
and U2484 (N_2484,In_2374,In_1360);
and U2485 (N_2485,In_649,In_828);
and U2486 (N_2486,In_539,In_2290);
xnor U2487 (N_2487,In_1938,In_1625);
nor U2488 (N_2488,In_1313,In_2453);
or U2489 (N_2489,In_951,In_770);
nand U2490 (N_2490,In_1371,In_812);
and U2491 (N_2491,In_1166,In_963);
or U2492 (N_2492,In_2264,In_833);
or U2493 (N_2493,In_1222,In_1130);
and U2494 (N_2494,In_1849,In_1418);
xor U2495 (N_2495,In_1806,In_2452);
nor U2496 (N_2496,In_1359,In_478);
or U2497 (N_2497,In_367,In_1785);
xnor U2498 (N_2498,In_511,In_1782);
or U2499 (N_2499,In_2328,In_1220);
nand U2500 (N_2500,In_1350,In_559);
nor U2501 (N_2501,In_2179,In_778);
or U2502 (N_2502,In_2023,In_1821);
or U2503 (N_2503,In_163,In_343);
or U2504 (N_2504,In_1431,In_264);
nor U2505 (N_2505,In_1192,In_181);
and U2506 (N_2506,In_105,In_1624);
nor U2507 (N_2507,In_1744,In_2406);
nor U2508 (N_2508,In_957,In_1767);
and U2509 (N_2509,In_418,In_1560);
and U2510 (N_2510,In_1875,In_1152);
nor U2511 (N_2511,In_1996,In_302);
nor U2512 (N_2512,In_1108,In_2452);
or U2513 (N_2513,In_924,In_971);
nor U2514 (N_2514,In_428,In_2275);
nand U2515 (N_2515,In_1933,In_1912);
nand U2516 (N_2516,In_1313,In_2105);
or U2517 (N_2517,In_34,In_246);
nand U2518 (N_2518,In_1835,In_112);
nand U2519 (N_2519,In_1856,In_1903);
and U2520 (N_2520,In_1702,In_1639);
or U2521 (N_2521,In_1726,In_1315);
and U2522 (N_2522,In_1915,In_500);
and U2523 (N_2523,In_2440,In_1149);
or U2524 (N_2524,In_1541,In_1206);
or U2525 (N_2525,In_287,In_2149);
or U2526 (N_2526,In_614,In_1519);
nor U2527 (N_2527,In_652,In_875);
or U2528 (N_2528,In_1843,In_381);
or U2529 (N_2529,In_2351,In_974);
nor U2530 (N_2530,In_2379,In_2051);
nand U2531 (N_2531,In_1490,In_2059);
nand U2532 (N_2532,In_198,In_1979);
nor U2533 (N_2533,In_1154,In_1294);
or U2534 (N_2534,In_841,In_2258);
and U2535 (N_2535,In_1208,In_188);
or U2536 (N_2536,In_249,In_2010);
nand U2537 (N_2537,In_1759,In_975);
nor U2538 (N_2538,In_483,In_1466);
xor U2539 (N_2539,In_2334,In_1037);
and U2540 (N_2540,In_1418,In_235);
or U2541 (N_2541,In_745,In_1222);
xor U2542 (N_2542,In_150,In_2294);
and U2543 (N_2543,In_867,In_1945);
or U2544 (N_2544,In_1461,In_275);
xnor U2545 (N_2545,In_1414,In_936);
and U2546 (N_2546,In_1176,In_2322);
xnor U2547 (N_2547,In_493,In_32);
nor U2548 (N_2548,In_853,In_2124);
or U2549 (N_2549,In_1911,In_1680);
or U2550 (N_2550,In_352,In_1915);
xor U2551 (N_2551,In_535,In_1928);
xor U2552 (N_2552,In_1479,In_1532);
or U2553 (N_2553,In_1163,In_435);
or U2554 (N_2554,In_1502,In_1084);
and U2555 (N_2555,In_322,In_1426);
or U2556 (N_2556,In_304,In_403);
nor U2557 (N_2557,In_1565,In_2287);
xnor U2558 (N_2558,In_1156,In_1370);
nand U2559 (N_2559,In_2277,In_1530);
and U2560 (N_2560,In_1751,In_2094);
and U2561 (N_2561,In_1749,In_1380);
and U2562 (N_2562,In_575,In_1816);
nor U2563 (N_2563,In_927,In_2484);
and U2564 (N_2564,In_173,In_446);
nand U2565 (N_2565,In_1281,In_535);
xnor U2566 (N_2566,In_851,In_1248);
nand U2567 (N_2567,In_2309,In_113);
or U2568 (N_2568,In_2255,In_2000);
and U2569 (N_2569,In_1498,In_916);
and U2570 (N_2570,In_519,In_32);
xnor U2571 (N_2571,In_251,In_2164);
and U2572 (N_2572,In_262,In_1293);
or U2573 (N_2573,In_230,In_1397);
and U2574 (N_2574,In_645,In_2216);
nand U2575 (N_2575,In_1952,In_267);
nand U2576 (N_2576,In_806,In_2429);
nand U2577 (N_2577,In_2177,In_227);
and U2578 (N_2578,In_605,In_88);
nor U2579 (N_2579,In_314,In_807);
nor U2580 (N_2580,In_1893,In_233);
nor U2581 (N_2581,In_439,In_560);
and U2582 (N_2582,In_2188,In_630);
and U2583 (N_2583,In_1535,In_198);
and U2584 (N_2584,In_901,In_1172);
and U2585 (N_2585,In_1367,In_329);
xor U2586 (N_2586,In_1528,In_571);
and U2587 (N_2587,In_1171,In_534);
xnor U2588 (N_2588,In_2167,In_1497);
or U2589 (N_2589,In_952,In_1571);
nand U2590 (N_2590,In_1325,In_1666);
nor U2591 (N_2591,In_1811,In_1182);
nand U2592 (N_2592,In_1474,In_2037);
xor U2593 (N_2593,In_2387,In_967);
xnor U2594 (N_2594,In_1210,In_2486);
or U2595 (N_2595,In_685,In_200);
nand U2596 (N_2596,In_1302,In_411);
nor U2597 (N_2597,In_2365,In_2203);
xnor U2598 (N_2598,In_1162,In_1150);
or U2599 (N_2599,In_662,In_611);
and U2600 (N_2600,In_1626,In_2306);
nand U2601 (N_2601,In_1571,In_1232);
and U2602 (N_2602,In_2096,In_680);
nor U2603 (N_2603,In_2433,In_2175);
nor U2604 (N_2604,In_568,In_1332);
nor U2605 (N_2605,In_2207,In_1994);
and U2606 (N_2606,In_2365,In_1210);
xnor U2607 (N_2607,In_1708,In_541);
xnor U2608 (N_2608,In_2239,In_1614);
or U2609 (N_2609,In_1799,In_223);
and U2610 (N_2610,In_707,In_1311);
xor U2611 (N_2611,In_661,In_2049);
or U2612 (N_2612,In_434,In_2132);
xor U2613 (N_2613,In_242,In_1486);
nand U2614 (N_2614,In_1592,In_2156);
nand U2615 (N_2615,In_1924,In_1455);
nor U2616 (N_2616,In_729,In_1610);
and U2617 (N_2617,In_96,In_1435);
and U2618 (N_2618,In_385,In_130);
or U2619 (N_2619,In_667,In_1880);
or U2620 (N_2620,In_1973,In_1932);
xor U2621 (N_2621,In_304,In_1472);
nor U2622 (N_2622,In_1189,In_1375);
or U2623 (N_2623,In_1573,In_2379);
nand U2624 (N_2624,In_666,In_273);
and U2625 (N_2625,In_406,In_2323);
nand U2626 (N_2626,In_1991,In_1);
xnor U2627 (N_2627,In_396,In_431);
or U2628 (N_2628,In_129,In_2393);
and U2629 (N_2629,In_1976,In_1557);
or U2630 (N_2630,In_310,In_2168);
or U2631 (N_2631,In_659,In_1672);
nor U2632 (N_2632,In_709,In_345);
or U2633 (N_2633,In_45,In_1265);
and U2634 (N_2634,In_341,In_1821);
xnor U2635 (N_2635,In_1722,In_234);
nor U2636 (N_2636,In_1192,In_2485);
xor U2637 (N_2637,In_32,In_1235);
or U2638 (N_2638,In_1432,In_114);
xnor U2639 (N_2639,In_2084,In_1106);
or U2640 (N_2640,In_1408,In_160);
or U2641 (N_2641,In_641,In_2364);
nor U2642 (N_2642,In_1713,In_210);
nand U2643 (N_2643,In_1276,In_1734);
or U2644 (N_2644,In_1340,In_1495);
xor U2645 (N_2645,In_1597,In_1391);
nor U2646 (N_2646,In_1603,In_1300);
nor U2647 (N_2647,In_1032,In_717);
xor U2648 (N_2648,In_2417,In_1755);
and U2649 (N_2649,In_1939,In_1783);
xor U2650 (N_2650,In_1724,In_2008);
nand U2651 (N_2651,In_1771,In_897);
xor U2652 (N_2652,In_790,In_1742);
or U2653 (N_2653,In_1845,In_430);
and U2654 (N_2654,In_486,In_728);
and U2655 (N_2655,In_2274,In_2079);
and U2656 (N_2656,In_1034,In_776);
nor U2657 (N_2657,In_1960,In_2119);
xnor U2658 (N_2658,In_724,In_2436);
and U2659 (N_2659,In_1626,In_1822);
nor U2660 (N_2660,In_869,In_1281);
nand U2661 (N_2661,In_917,In_2156);
xnor U2662 (N_2662,In_1027,In_2416);
xnor U2663 (N_2663,In_1598,In_2064);
xnor U2664 (N_2664,In_2170,In_1000);
nand U2665 (N_2665,In_1498,In_49);
or U2666 (N_2666,In_1518,In_2349);
and U2667 (N_2667,In_2215,In_1102);
and U2668 (N_2668,In_1930,In_127);
or U2669 (N_2669,In_2040,In_1631);
or U2670 (N_2670,In_161,In_1116);
xor U2671 (N_2671,In_2039,In_1428);
xor U2672 (N_2672,In_2035,In_1988);
and U2673 (N_2673,In_2447,In_561);
xor U2674 (N_2674,In_2483,In_2341);
xnor U2675 (N_2675,In_1004,In_2289);
nand U2676 (N_2676,In_2495,In_1601);
xnor U2677 (N_2677,In_1431,In_755);
xnor U2678 (N_2678,In_947,In_1224);
and U2679 (N_2679,In_603,In_1569);
or U2680 (N_2680,In_438,In_759);
nor U2681 (N_2681,In_1578,In_1323);
nand U2682 (N_2682,In_1409,In_2204);
xnor U2683 (N_2683,In_2484,In_2128);
nand U2684 (N_2684,In_547,In_936);
nor U2685 (N_2685,In_2111,In_280);
nor U2686 (N_2686,In_308,In_2063);
and U2687 (N_2687,In_2351,In_434);
nand U2688 (N_2688,In_740,In_1541);
or U2689 (N_2689,In_2239,In_1010);
nor U2690 (N_2690,In_1026,In_1435);
xnor U2691 (N_2691,In_129,In_753);
nand U2692 (N_2692,In_401,In_1716);
nand U2693 (N_2693,In_1417,In_2088);
and U2694 (N_2694,In_2182,In_2090);
nand U2695 (N_2695,In_623,In_846);
xor U2696 (N_2696,In_871,In_1848);
nor U2697 (N_2697,In_71,In_1466);
and U2698 (N_2698,In_1912,In_842);
nor U2699 (N_2699,In_2093,In_1501);
or U2700 (N_2700,In_1922,In_500);
and U2701 (N_2701,In_762,In_1319);
nor U2702 (N_2702,In_1481,In_50);
and U2703 (N_2703,In_1681,In_1554);
or U2704 (N_2704,In_411,In_205);
and U2705 (N_2705,In_2126,In_2420);
nand U2706 (N_2706,In_1113,In_607);
and U2707 (N_2707,In_2219,In_1202);
nor U2708 (N_2708,In_2055,In_1791);
and U2709 (N_2709,In_584,In_1678);
or U2710 (N_2710,In_1201,In_756);
nand U2711 (N_2711,In_1038,In_1231);
nand U2712 (N_2712,In_709,In_2002);
nand U2713 (N_2713,In_2090,In_2222);
xnor U2714 (N_2714,In_2183,In_573);
or U2715 (N_2715,In_126,In_745);
and U2716 (N_2716,In_1521,In_944);
xor U2717 (N_2717,In_1659,In_549);
or U2718 (N_2718,In_2093,In_1803);
or U2719 (N_2719,In_1638,In_221);
and U2720 (N_2720,In_1750,In_1320);
nor U2721 (N_2721,In_212,In_2146);
nor U2722 (N_2722,In_2054,In_1864);
xor U2723 (N_2723,In_1602,In_36);
nand U2724 (N_2724,In_2486,In_311);
nor U2725 (N_2725,In_1215,In_351);
or U2726 (N_2726,In_1518,In_359);
nand U2727 (N_2727,In_2030,In_1951);
and U2728 (N_2728,In_66,In_654);
and U2729 (N_2729,In_1045,In_493);
and U2730 (N_2730,In_597,In_966);
or U2731 (N_2731,In_959,In_1712);
nand U2732 (N_2732,In_1972,In_1963);
xnor U2733 (N_2733,In_68,In_1996);
xor U2734 (N_2734,In_2056,In_1030);
and U2735 (N_2735,In_1375,In_1617);
xnor U2736 (N_2736,In_1573,In_1849);
nor U2737 (N_2737,In_818,In_1156);
nor U2738 (N_2738,In_2183,In_1180);
xor U2739 (N_2739,In_1011,In_482);
and U2740 (N_2740,In_1211,In_54);
nor U2741 (N_2741,In_1571,In_442);
nor U2742 (N_2742,In_1801,In_1573);
or U2743 (N_2743,In_1517,In_873);
nand U2744 (N_2744,In_401,In_340);
or U2745 (N_2745,In_1120,In_73);
xor U2746 (N_2746,In_355,In_2004);
or U2747 (N_2747,In_468,In_351);
or U2748 (N_2748,In_1869,In_687);
nand U2749 (N_2749,In_2491,In_348);
nor U2750 (N_2750,In_1183,In_2035);
nor U2751 (N_2751,In_817,In_952);
and U2752 (N_2752,In_725,In_2485);
xnor U2753 (N_2753,In_1845,In_1991);
nand U2754 (N_2754,In_349,In_790);
and U2755 (N_2755,In_2292,In_1695);
nand U2756 (N_2756,In_1277,In_2062);
xor U2757 (N_2757,In_32,In_734);
nand U2758 (N_2758,In_1860,In_2378);
xor U2759 (N_2759,In_940,In_1151);
or U2760 (N_2760,In_230,In_527);
or U2761 (N_2761,In_1317,In_1047);
nor U2762 (N_2762,In_1411,In_476);
or U2763 (N_2763,In_376,In_2484);
or U2764 (N_2764,In_1279,In_231);
xnor U2765 (N_2765,In_283,In_137);
nand U2766 (N_2766,In_2029,In_741);
and U2767 (N_2767,In_83,In_327);
or U2768 (N_2768,In_707,In_1437);
nand U2769 (N_2769,In_302,In_2049);
nor U2770 (N_2770,In_2490,In_1376);
and U2771 (N_2771,In_2433,In_295);
and U2772 (N_2772,In_2281,In_356);
and U2773 (N_2773,In_3,In_1987);
nor U2774 (N_2774,In_325,In_1928);
nand U2775 (N_2775,In_2058,In_879);
or U2776 (N_2776,In_1219,In_2444);
nor U2777 (N_2777,In_64,In_1559);
nor U2778 (N_2778,In_2070,In_135);
xnor U2779 (N_2779,In_556,In_2130);
nor U2780 (N_2780,In_1724,In_2144);
nand U2781 (N_2781,In_32,In_2322);
and U2782 (N_2782,In_1661,In_866);
nor U2783 (N_2783,In_2050,In_583);
or U2784 (N_2784,In_964,In_2054);
nand U2785 (N_2785,In_2338,In_1129);
nand U2786 (N_2786,In_1514,In_292);
and U2787 (N_2787,In_1761,In_1266);
nand U2788 (N_2788,In_2256,In_1790);
or U2789 (N_2789,In_1374,In_7);
and U2790 (N_2790,In_660,In_263);
xnor U2791 (N_2791,In_1284,In_2261);
and U2792 (N_2792,In_1671,In_2286);
or U2793 (N_2793,In_2421,In_1117);
or U2794 (N_2794,In_2291,In_1023);
or U2795 (N_2795,In_1959,In_938);
nand U2796 (N_2796,In_2339,In_477);
or U2797 (N_2797,In_357,In_1830);
and U2798 (N_2798,In_2370,In_1234);
and U2799 (N_2799,In_1839,In_1710);
xor U2800 (N_2800,In_1783,In_557);
nand U2801 (N_2801,In_2483,In_1039);
nand U2802 (N_2802,In_2404,In_1486);
or U2803 (N_2803,In_1258,In_1335);
xnor U2804 (N_2804,In_740,In_732);
nand U2805 (N_2805,In_1672,In_556);
nor U2806 (N_2806,In_584,In_1254);
and U2807 (N_2807,In_2333,In_2277);
nand U2808 (N_2808,In_490,In_2020);
nor U2809 (N_2809,In_1809,In_2045);
nand U2810 (N_2810,In_2391,In_2480);
and U2811 (N_2811,In_1028,In_2488);
and U2812 (N_2812,In_2068,In_1618);
nand U2813 (N_2813,In_1764,In_838);
nor U2814 (N_2814,In_1225,In_1365);
xnor U2815 (N_2815,In_780,In_1377);
nand U2816 (N_2816,In_2461,In_2479);
or U2817 (N_2817,In_2231,In_21);
nor U2818 (N_2818,In_976,In_2368);
or U2819 (N_2819,In_668,In_215);
nand U2820 (N_2820,In_2457,In_1180);
and U2821 (N_2821,In_622,In_1592);
and U2822 (N_2822,In_2490,In_1788);
nor U2823 (N_2823,In_1027,In_1161);
xor U2824 (N_2824,In_68,In_20);
and U2825 (N_2825,In_319,In_784);
and U2826 (N_2826,In_32,In_1035);
and U2827 (N_2827,In_1394,In_6);
and U2828 (N_2828,In_110,In_1225);
and U2829 (N_2829,In_1214,In_503);
and U2830 (N_2830,In_1515,In_1598);
or U2831 (N_2831,In_757,In_912);
nand U2832 (N_2832,In_629,In_1139);
and U2833 (N_2833,In_1889,In_460);
xor U2834 (N_2834,In_2291,In_1643);
nor U2835 (N_2835,In_1399,In_1823);
nor U2836 (N_2836,In_874,In_674);
nand U2837 (N_2837,In_918,In_1806);
nand U2838 (N_2838,In_1479,In_2431);
or U2839 (N_2839,In_919,In_2253);
or U2840 (N_2840,In_1782,In_2388);
and U2841 (N_2841,In_2410,In_1505);
nand U2842 (N_2842,In_2446,In_1255);
and U2843 (N_2843,In_244,In_2102);
nor U2844 (N_2844,In_244,In_2292);
nor U2845 (N_2845,In_241,In_1974);
or U2846 (N_2846,In_901,In_2024);
and U2847 (N_2847,In_1642,In_171);
or U2848 (N_2848,In_1396,In_1004);
nand U2849 (N_2849,In_2233,In_1310);
xor U2850 (N_2850,In_781,In_820);
nor U2851 (N_2851,In_1310,In_2157);
xnor U2852 (N_2852,In_393,In_171);
nor U2853 (N_2853,In_2371,In_2155);
or U2854 (N_2854,In_1689,In_1314);
nor U2855 (N_2855,In_892,In_1389);
xor U2856 (N_2856,In_2151,In_2464);
and U2857 (N_2857,In_1540,In_739);
and U2858 (N_2858,In_2187,In_1446);
nand U2859 (N_2859,In_453,In_180);
or U2860 (N_2860,In_1374,In_513);
nand U2861 (N_2861,In_203,In_1997);
and U2862 (N_2862,In_365,In_356);
and U2863 (N_2863,In_912,In_1112);
nor U2864 (N_2864,In_1031,In_1887);
nor U2865 (N_2865,In_1074,In_98);
nand U2866 (N_2866,In_2495,In_2267);
nor U2867 (N_2867,In_1968,In_2059);
nor U2868 (N_2868,In_12,In_861);
and U2869 (N_2869,In_1533,In_483);
and U2870 (N_2870,In_1604,In_869);
nor U2871 (N_2871,In_993,In_69);
and U2872 (N_2872,In_358,In_91);
xnor U2873 (N_2873,In_1047,In_1921);
nand U2874 (N_2874,In_1013,In_24);
nor U2875 (N_2875,In_1749,In_1);
nor U2876 (N_2876,In_533,In_135);
nand U2877 (N_2877,In_1344,In_953);
and U2878 (N_2878,In_1644,In_132);
nor U2879 (N_2879,In_2082,In_2139);
nand U2880 (N_2880,In_1600,In_2351);
nand U2881 (N_2881,In_445,In_1513);
nor U2882 (N_2882,In_1693,In_1253);
nand U2883 (N_2883,In_2145,In_1821);
nand U2884 (N_2884,In_769,In_470);
nand U2885 (N_2885,In_2215,In_2153);
and U2886 (N_2886,In_587,In_1640);
nand U2887 (N_2887,In_2434,In_364);
nand U2888 (N_2888,In_1001,In_1970);
nand U2889 (N_2889,In_1335,In_2047);
xor U2890 (N_2890,In_1775,In_1222);
or U2891 (N_2891,In_1451,In_1894);
or U2892 (N_2892,In_1797,In_546);
or U2893 (N_2893,In_1337,In_249);
nor U2894 (N_2894,In_1931,In_651);
nand U2895 (N_2895,In_1314,In_1730);
nand U2896 (N_2896,In_1990,In_928);
and U2897 (N_2897,In_775,In_1362);
xor U2898 (N_2898,In_992,In_126);
and U2899 (N_2899,In_1577,In_379);
xor U2900 (N_2900,In_2261,In_1139);
or U2901 (N_2901,In_360,In_523);
xnor U2902 (N_2902,In_1594,In_674);
and U2903 (N_2903,In_1977,In_213);
xnor U2904 (N_2904,In_1225,In_1957);
and U2905 (N_2905,In_555,In_174);
xnor U2906 (N_2906,In_1575,In_2486);
nor U2907 (N_2907,In_385,In_2460);
or U2908 (N_2908,In_27,In_317);
nor U2909 (N_2909,In_2085,In_1798);
nand U2910 (N_2910,In_26,In_1450);
or U2911 (N_2911,In_1932,In_1155);
nor U2912 (N_2912,In_2224,In_1315);
nor U2913 (N_2913,In_1201,In_1160);
and U2914 (N_2914,In_1185,In_1737);
and U2915 (N_2915,In_9,In_1359);
nand U2916 (N_2916,In_473,In_2284);
and U2917 (N_2917,In_1976,In_1970);
nor U2918 (N_2918,In_953,In_2451);
or U2919 (N_2919,In_153,In_2122);
or U2920 (N_2920,In_121,In_894);
nand U2921 (N_2921,In_1071,In_359);
nand U2922 (N_2922,In_1055,In_2265);
xor U2923 (N_2923,In_1150,In_1293);
nor U2924 (N_2924,In_1337,In_280);
nor U2925 (N_2925,In_1857,In_579);
and U2926 (N_2926,In_1229,In_238);
or U2927 (N_2927,In_660,In_810);
nor U2928 (N_2928,In_2487,In_1481);
xor U2929 (N_2929,In_2169,In_2371);
nor U2930 (N_2930,In_2290,In_2167);
nor U2931 (N_2931,In_1750,In_744);
nor U2932 (N_2932,In_1200,In_1970);
nor U2933 (N_2933,In_2445,In_1798);
xor U2934 (N_2934,In_1519,In_1367);
and U2935 (N_2935,In_553,In_961);
xnor U2936 (N_2936,In_1165,In_1019);
nor U2937 (N_2937,In_2386,In_297);
or U2938 (N_2938,In_1117,In_2393);
and U2939 (N_2939,In_354,In_530);
nand U2940 (N_2940,In_1727,In_1640);
nand U2941 (N_2941,In_1322,In_1207);
nor U2942 (N_2942,In_1777,In_2322);
nand U2943 (N_2943,In_28,In_2149);
nand U2944 (N_2944,In_2442,In_1741);
and U2945 (N_2945,In_1039,In_1212);
or U2946 (N_2946,In_1014,In_403);
and U2947 (N_2947,In_1208,In_2365);
and U2948 (N_2948,In_1287,In_1713);
or U2949 (N_2949,In_493,In_2379);
nand U2950 (N_2950,In_1769,In_874);
or U2951 (N_2951,In_597,In_724);
and U2952 (N_2952,In_2421,In_753);
xor U2953 (N_2953,In_989,In_2142);
nand U2954 (N_2954,In_2490,In_1549);
xor U2955 (N_2955,In_135,In_1059);
nand U2956 (N_2956,In_931,In_682);
nor U2957 (N_2957,In_1767,In_1164);
nor U2958 (N_2958,In_1596,In_1406);
and U2959 (N_2959,In_733,In_2088);
and U2960 (N_2960,In_1982,In_426);
nand U2961 (N_2961,In_1909,In_22);
nor U2962 (N_2962,In_703,In_2375);
nor U2963 (N_2963,In_986,In_867);
xnor U2964 (N_2964,In_215,In_1792);
nand U2965 (N_2965,In_2362,In_860);
nand U2966 (N_2966,In_1789,In_601);
and U2967 (N_2967,In_2321,In_144);
nor U2968 (N_2968,In_387,In_369);
or U2969 (N_2969,In_2263,In_1641);
xor U2970 (N_2970,In_1119,In_575);
or U2971 (N_2971,In_709,In_475);
or U2972 (N_2972,In_1883,In_1754);
or U2973 (N_2973,In_297,In_1285);
and U2974 (N_2974,In_1569,In_352);
and U2975 (N_2975,In_1618,In_1296);
or U2976 (N_2976,In_678,In_2346);
xnor U2977 (N_2977,In_2378,In_681);
or U2978 (N_2978,In_2441,In_29);
or U2979 (N_2979,In_1276,In_1978);
nand U2980 (N_2980,In_785,In_507);
and U2981 (N_2981,In_1246,In_558);
or U2982 (N_2982,In_1775,In_2329);
and U2983 (N_2983,In_223,In_531);
or U2984 (N_2984,In_1543,In_2261);
xnor U2985 (N_2985,In_2437,In_1309);
xnor U2986 (N_2986,In_1593,In_396);
or U2987 (N_2987,In_1362,In_25);
and U2988 (N_2988,In_994,In_199);
nand U2989 (N_2989,In_90,In_111);
nand U2990 (N_2990,In_1626,In_630);
xnor U2991 (N_2991,In_103,In_1075);
or U2992 (N_2992,In_1500,In_2245);
nor U2993 (N_2993,In_137,In_1322);
xor U2994 (N_2994,In_126,In_342);
or U2995 (N_2995,In_2459,In_1809);
nor U2996 (N_2996,In_1977,In_813);
and U2997 (N_2997,In_907,In_2017);
xor U2998 (N_2998,In_1332,In_1929);
nor U2999 (N_2999,In_1499,In_109);
nor U3000 (N_3000,In_2232,In_1402);
and U3001 (N_3001,In_1947,In_2019);
nand U3002 (N_3002,In_1722,In_379);
nand U3003 (N_3003,In_1672,In_486);
or U3004 (N_3004,In_1786,In_1027);
or U3005 (N_3005,In_2206,In_477);
xnor U3006 (N_3006,In_1264,In_196);
and U3007 (N_3007,In_1660,In_81);
nor U3008 (N_3008,In_316,In_1374);
and U3009 (N_3009,In_834,In_413);
xor U3010 (N_3010,In_2345,In_1127);
nand U3011 (N_3011,In_1530,In_1287);
nand U3012 (N_3012,In_55,In_839);
or U3013 (N_3013,In_2119,In_255);
xor U3014 (N_3014,In_622,In_1540);
nor U3015 (N_3015,In_726,In_569);
nand U3016 (N_3016,In_1799,In_459);
and U3017 (N_3017,In_2302,In_1356);
nor U3018 (N_3018,In_1341,In_873);
or U3019 (N_3019,In_353,In_1044);
xnor U3020 (N_3020,In_2020,In_2470);
nor U3021 (N_3021,In_2311,In_1120);
xnor U3022 (N_3022,In_1032,In_2030);
nand U3023 (N_3023,In_327,In_922);
xnor U3024 (N_3024,In_2182,In_807);
xor U3025 (N_3025,In_1044,In_1719);
xnor U3026 (N_3026,In_1210,In_2288);
and U3027 (N_3027,In_1178,In_2321);
xnor U3028 (N_3028,In_2432,In_1820);
and U3029 (N_3029,In_513,In_373);
nor U3030 (N_3030,In_346,In_426);
nand U3031 (N_3031,In_1931,In_2390);
nand U3032 (N_3032,In_2366,In_155);
and U3033 (N_3033,In_500,In_2025);
nand U3034 (N_3034,In_431,In_933);
xor U3035 (N_3035,In_1891,In_1082);
and U3036 (N_3036,In_2259,In_1408);
or U3037 (N_3037,In_1637,In_177);
nand U3038 (N_3038,In_106,In_1252);
or U3039 (N_3039,In_1820,In_114);
or U3040 (N_3040,In_1228,In_1174);
nor U3041 (N_3041,In_1631,In_1130);
nor U3042 (N_3042,In_2155,In_1305);
nand U3043 (N_3043,In_2137,In_1824);
or U3044 (N_3044,In_1677,In_93);
xnor U3045 (N_3045,In_2464,In_1945);
nor U3046 (N_3046,In_1337,In_1430);
or U3047 (N_3047,In_879,In_2349);
nand U3048 (N_3048,In_1341,In_602);
nor U3049 (N_3049,In_270,In_1622);
and U3050 (N_3050,In_1253,In_972);
or U3051 (N_3051,In_1624,In_1842);
nand U3052 (N_3052,In_1121,In_2101);
and U3053 (N_3053,In_950,In_1472);
and U3054 (N_3054,In_775,In_2128);
xor U3055 (N_3055,In_2198,In_1671);
and U3056 (N_3056,In_1275,In_1226);
nor U3057 (N_3057,In_1677,In_1537);
or U3058 (N_3058,In_719,In_1273);
nand U3059 (N_3059,In_1674,In_2261);
xor U3060 (N_3060,In_1313,In_537);
nor U3061 (N_3061,In_401,In_2261);
and U3062 (N_3062,In_1711,In_2364);
xnor U3063 (N_3063,In_1375,In_46);
or U3064 (N_3064,In_600,In_2216);
xnor U3065 (N_3065,In_2274,In_1827);
nand U3066 (N_3066,In_1836,In_1409);
or U3067 (N_3067,In_1818,In_2071);
nor U3068 (N_3068,In_1673,In_2207);
or U3069 (N_3069,In_1648,In_806);
or U3070 (N_3070,In_980,In_1892);
or U3071 (N_3071,In_510,In_2426);
or U3072 (N_3072,In_222,In_2372);
xor U3073 (N_3073,In_1948,In_2361);
and U3074 (N_3074,In_787,In_637);
xor U3075 (N_3075,In_43,In_2046);
nand U3076 (N_3076,In_1838,In_2367);
and U3077 (N_3077,In_1165,In_2049);
or U3078 (N_3078,In_1422,In_1575);
xnor U3079 (N_3079,In_667,In_2347);
nand U3080 (N_3080,In_435,In_1645);
and U3081 (N_3081,In_2446,In_1996);
or U3082 (N_3082,In_2027,In_58);
xor U3083 (N_3083,In_436,In_1180);
or U3084 (N_3084,In_505,In_1618);
and U3085 (N_3085,In_1806,In_1717);
and U3086 (N_3086,In_1668,In_100);
or U3087 (N_3087,In_1516,In_297);
nor U3088 (N_3088,In_1190,In_1026);
nand U3089 (N_3089,In_788,In_1909);
nand U3090 (N_3090,In_1471,In_2010);
or U3091 (N_3091,In_1867,In_2399);
xor U3092 (N_3092,In_569,In_401);
nand U3093 (N_3093,In_1050,In_1776);
or U3094 (N_3094,In_853,In_466);
nor U3095 (N_3095,In_1503,In_465);
nor U3096 (N_3096,In_1180,In_930);
or U3097 (N_3097,In_582,In_1458);
or U3098 (N_3098,In_1101,In_618);
nand U3099 (N_3099,In_700,In_719);
or U3100 (N_3100,In_577,In_977);
nor U3101 (N_3101,In_2037,In_2092);
nand U3102 (N_3102,In_1430,In_2384);
and U3103 (N_3103,In_31,In_1777);
xor U3104 (N_3104,In_870,In_1609);
and U3105 (N_3105,In_89,In_1394);
nor U3106 (N_3106,In_584,In_706);
nor U3107 (N_3107,In_2456,In_1107);
xnor U3108 (N_3108,In_1944,In_1060);
nand U3109 (N_3109,In_798,In_264);
or U3110 (N_3110,In_47,In_2149);
xor U3111 (N_3111,In_2463,In_1955);
nand U3112 (N_3112,In_1965,In_1132);
nor U3113 (N_3113,In_738,In_877);
nand U3114 (N_3114,In_1309,In_757);
xnor U3115 (N_3115,In_1184,In_992);
or U3116 (N_3116,In_1205,In_1907);
nand U3117 (N_3117,In_1785,In_211);
xor U3118 (N_3118,In_434,In_2203);
and U3119 (N_3119,In_1832,In_195);
or U3120 (N_3120,In_1715,In_2471);
nand U3121 (N_3121,In_698,In_1088);
or U3122 (N_3122,In_1935,In_276);
nor U3123 (N_3123,In_1930,In_295);
nor U3124 (N_3124,In_2012,In_2029);
xor U3125 (N_3125,N_88,N_1390);
xor U3126 (N_3126,N_684,N_1268);
or U3127 (N_3127,N_2937,N_1104);
nand U3128 (N_3128,N_2758,N_1361);
nor U3129 (N_3129,N_359,N_1605);
nand U3130 (N_3130,N_53,N_609);
and U3131 (N_3131,N_294,N_534);
nor U3132 (N_3132,N_3067,N_2185);
or U3133 (N_3133,N_204,N_1915);
xor U3134 (N_3134,N_829,N_2754);
nor U3135 (N_3135,N_1671,N_1971);
nor U3136 (N_3136,N_437,N_1124);
xor U3137 (N_3137,N_1501,N_2112);
or U3138 (N_3138,N_645,N_1843);
xnor U3139 (N_3139,N_599,N_778);
or U3140 (N_3140,N_1591,N_1481);
and U3141 (N_3141,N_2459,N_1836);
nand U3142 (N_3142,N_1767,N_1326);
or U3143 (N_3143,N_2681,N_1386);
nand U3144 (N_3144,N_263,N_1012);
and U3145 (N_3145,N_1623,N_2542);
xnor U3146 (N_3146,N_2197,N_2016);
xnor U3147 (N_3147,N_535,N_2161);
and U3148 (N_3148,N_1822,N_668);
or U3149 (N_3149,N_3054,N_1788);
or U3150 (N_3150,N_2799,N_2828);
nor U3151 (N_3151,N_991,N_2104);
and U3152 (N_3152,N_488,N_944);
nand U3153 (N_3153,N_1436,N_107);
or U3154 (N_3154,N_981,N_949);
and U3155 (N_3155,N_2117,N_508);
xnor U3156 (N_3156,N_2254,N_2956);
nor U3157 (N_3157,N_281,N_2687);
and U3158 (N_3158,N_1205,N_186);
xnor U3159 (N_3159,N_2826,N_2794);
nand U3160 (N_3160,N_1022,N_1113);
nand U3161 (N_3161,N_2830,N_3089);
and U3162 (N_3162,N_142,N_2417);
and U3163 (N_3163,N_3092,N_293);
and U3164 (N_3164,N_1457,N_933);
and U3165 (N_3165,N_1450,N_1017);
or U3166 (N_3166,N_2227,N_2388);
and U3167 (N_3167,N_2684,N_966);
nor U3168 (N_3168,N_223,N_209);
xnor U3169 (N_3169,N_3064,N_1860);
or U3170 (N_3170,N_1429,N_2887);
xnor U3171 (N_3171,N_3005,N_1520);
nand U3172 (N_3172,N_2603,N_1564);
nand U3173 (N_3173,N_2389,N_737);
nor U3174 (N_3174,N_34,N_2840);
xnor U3175 (N_3175,N_1695,N_271);
and U3176 (N_3176,N_1459,N_208);
nor U3177 (N_3177,N_1762,N_4);
nand U3178 (N_3178,N_901,N_279);
and U3179 (N_3179,N_137,N_2962);
and U3180 (N_3180,N_2678,N_1280);
or U3181 (N_3181,N_1653,N_995);
nor U3182 (N_3182,N_3118,N_2636);
or U3183 (N_3183,N_2346,N_2610);
and U3184 (N_3184,N_2436,N_809);
nand U3185 (N_3185,N_2215,N_1829);
xnor U3186 (N_3186,N_986,N_2420);
nand U3187 (N_3187,N_461,N_1147);
nand U3188 (N_3188,N_2852,N_1743);
nand U3189 (N_3189,N_1899,N_1275);
and U3190 (N_3190,N_808,N_1406);
xnor U3191 (N_3191,N_554,N_18);
xor U3192 (N_3192,N_1435,N_1444);
nor U3193 (N_3193,N_1222,N_196);
nand U3194 (N_3194,N_2866,N_1865);
and U3195 (N_3195,N_1988,N_2409);
xor U3196 (N_3196,N_1905,N_1417);
nand U3197 (N_3197,N_699,N_1054);
xor U3198 (N_3198,N_1438,N_2317);
nand U3199 (N_3199,N_1560,N_1993);
xor U3200 (N_3200,N_487,N_2963);
nor U3201 (N_3201,N_2219,N_1688);
nand U3202 (N_3202,N_2570,N_265);
or U3203 (N_3203,N_1439,N_2623);
and U3204 (N_3204,N_1904,N_1981);
xnor U3205 (N_3205,N_185,N_1835);
nor U3206 (N_3206,N_1462,N_584);
or U3207 (N_3207,N_909,N_1954);
nor U3208 (N_3208,N_2070,N_568);
and U3209 (N_3209,N_2903,N_2045);
xnor U3210 (N_3210,N_2637,N_1402);
nor U3211 (N_3211,N_375,N_1344);
nor U3212 (N_3212,N_1534,N_2128);
and U3213 (N_3213,N_2474,N_2783);
xnor U3214 (N_3214,N_1952,N_15);
or U3215 (N_3215,N_3081,N_2911);
and U3216 (N_3216,N_1182,N_2562);
xor U3217 (N_3217,N_754,N_2785);
or U3218 (N_3218,N_2088,N_2546);
nand U3219 (N_3219,N_1109,N_1223);
and U3220 (N_3220,N_2941,N_1728);
and U3221 (N_3221,N_2976,N_3026);
nor U3222 (N_3222,N_3091,N_2527);
xnor U3223 (N_3223,N_1261,N_2136);
nor U3224 (N_3224,N_575,N_2156);
or U3225 (N_3225,N_1764,N_132);
and U3226 (N_3226,N_2931,N_2113);
nor U3227 (N_3227,N_750,N_150);
and U3228 (N_3228,N_2877,N_937);
nand U3229 (N_3229,N_2449,N_2705);
and U3230 (N_3230,N_963,N_2853);
or U3231 (N_3231,N_1946,N_2402);
and U3232 (N_3232,N_708,N_1136);
nand U3233 (N_3233,N_690,N_190);
xnor U3234 (N_3234,N_1575,N_2658);
nor U3235 (N_3235,N_1636,N_1755);
and U3236 (N_3236,N_540,N_2448);
nor U3237 (N_3237,N_2593,N_2737);
nor U3238 (N_3238,N_449,N_2279);
or U3239 (N_3239,N_1831,N_2103);
nor U3240 (N_3240,N_2429,N_1309);
nor U3241 (N_3241,N_1687,N_1141);
nand U3242 (N_3242,N_1121,N_2632);
xor U3243 (N_3243,N_510,N_358);
or U3244 (N_3244,N_2290,N_1974);
xnor U3245 (N_3245,N_843,N_1286);
and U3246 (N_3246,N_2578,N_1738);
and U3247 (N_3247,N_2564,N_1737);
xor U3248 (N_3248,N_2005,N_2200);
nor U3249 (N_3249,N_1046,N_1292);
nor U3250 (N_3250,N_2985,N_1067);
nand U3251 (N_3251,N_466,N_1320);
and U3252 (N_3252,N_173,N_2944);
xor U3253 (N_3253,N_946,N_2999);
nor U3254 (N_3254,N_2790,N_2524);
and U3255 (N_3255,N_739,N_1886);
nand U3256 (N_3256,N_1706,N_2888);
or U3257 (N_3257,N_1165,N_528);
or U3258 (N_3258,N_2968,N_112);
and U3259 (N_3259,N_861,N_194);
nand U3260 (N_3260,N_598,N_974);
and U3261 (N_3261,N_1805,N_2745);
nand U3262 (N_3262,N_2577,N_2349);
or U3263 (N_3263,N_1015,N_2509);
nor U3264 (N_3264,N_386,N_2867);
or U3265 (N_3265,N_1639,N_1630);
nor U3266 (N_3266,N_700,N_2195);
or U3267 (N_3267,N_2316,N_49);
nand U3268 (N_3268,N_2686,N_2833);
nor U3269 (N_3269,N_1563,N_2393);
and U3270 (N_3270,N_694,N_3053);
xnor U3271 (N_3271,N_2808,N_1152);
xor U3272 (N_3272,N_1503,N_2476);
nor U3273 (N_3273,N_727,N_845);
nand U3274 (N_3274,N_2299,N_311);
and U3275 (N_3275,N_893,N_1255);
nor U3276 (N_3276,N_1778,N_1224);
nor U3277 (N_3277,N_2364,N_2955);
and U3278 (N_3278,N_369,N_717);
and U3279 (N_3279,N_695,N_734);
or U3280 (N_3280,N_563,N_2077);
xnor U3281 (N_3281,N_2099,N_1019);
nand U3282 (N_3282,N_2120,N_3102);
nor U3283 (N_3283,N_2488,N_1812);
and U3284 (N_3284,N_116,N_1960);
xor U3285 (N_3285,N_570,N_309);
nand U3286 (N_3286,N_2276,N_2368);
nand U3287 (N_3287,N_2143,N_51);
or U3288 (N_3288,N_1134,N_2525);
and U3289 (N_3289,N_62,N_1279);
nor U3290 (N_3290,N_1799,N_2266);
or U3291 (N_3291,N_1139,N_2567);
or U3292 (N_3292,N_1098,N_240);
nor U3293 (N_3293,N_26,N_2454);
nand U3294 (N_3294,N_1825,N_3036);
nand U3295 (N_3295,N_2157,N_1162);
nand U3296 (N_3296,N_2190,N_2739);
nor U3297 (N_3297,N_644,N_926);
or U3298 (N_3298,N_280,N_2773);
nand U3299 (N_3299,N_1202,N_1685);
xor U3300 (N_3300,N_622,N_1794);
xor U3301 (N_3301,N_2089,N_1854);
xor U3302 (N_3302,N_648,N_1911);
nand U3303 (N_3303,N_2587,N_463);
nand U3304 (N_3304,N_658,N_2924);
xnor U3305 (N_3305,N_2897,N_2856);
nand U3306 (N_3306,N_1285,N_217);
nand U3307 (N_3307,N_1164,N_2443);
xnor U3308 (N_3308,N_678,N_191);
nor U3309 (N_3309,N_1416,N_2304);
and U3310 (N_3310,N_1317,N_1287);
nand U3311 (N_3311,N_2249,N_2093);
xnor U3312 (N_3312,N_958,N_3056);
nor U3313 (N_3313,N_1138,N_774);
nand U3314 (N_3314,N_121,N_1426);
nand U3315 (N_3315,N_2134,N_2118);
xnor U3316 (N_3316,N_682,N_2683);
and U3317 (N_3317,N_2600,N_101);
and U3318 (N_3318,N_925,N_2170);
or U3319 (N_3319,N_3079,N_788);
or U3320 (N_3320,N_670,N_1477);
nand U3321 (N_3321,N_3008,N_3070);
xnor U3322 (N_3322,N_1568,N_1909);
and U3323 (N_3323,N_1670,N_122);
xor U3324 (N_3324,N_1561,N_2614);
xnor U3325 (N_3325,N_1510,N_2321);
and U3326 (N_3326,N_1272,N_2064);
or U3327 (N_3327,N_701,N_274);
and U3328 (N_3328,N_206,N_1385);
and U3329 (N_3329,N_1025,N_2302);
xnor U3330 (N_3330,N_2895,N_2504);
nor U3331 (N_3331,N_1731,N_702);
xor U3332 (N_3332,N_485,N_1947);
and U3333 (N_3333,N_432,N_1919);
nor U3334 (N_3334,N_1972,N_5);
nor U3335 (N_3335,N_1772,N_400);
xnor U3336 (N_3336,N_1745,N_320);
nor U3337 (N_3337,N_533,N_1232);
nor U3338 (N_3338,N_1902,N_520);
or U3339 (N_3339,N_591,N_1966);
nor U3340 (N_3340,N_3060,N_1316);
xnor U3341 (N_3341,N_742,N_2668);
or U3342 (N_3342,N_1662,N_356);
or U3343 (N_3343,N_833,N_2966);
and U3344 (N_3344,N_3065,N_2996);
nand U3345 (N_3345,N_525,N_831);
nand U3346 (N_3346,N_2286,N_1199);
nand U3347 (N_3347,N_2141,N_342);
nand U3348 (N_3348,N_1242,N_257);
nand U3349 (N_3349,N_420,N_1415);
nor U3350 (N_3350,N_667,N_1346);
and U3351 (N_3351,N_3093,N_2814);
xnor U3352 (N_3352,N_2182,N_2842);
nand U3353 (N_3353,N_1618,N_59);
nor U3354 (N_3354,N_1768,N_354);
and U3355 (N_3355,N_1890,N_552);
xnor U3356 (N_3356,N_43,N_847);
xor U3357 (N_3357,N_1424,N_1403);
xnor U3358 (N_3358,N_2152,N_2601);
nand U3359 (N_3359,N_1075,N_2169);
nand U3360 (N_3360,N_2029,N_1889);
xor U3361 (N_3361,N_2934,N_2554);
xor U3362 (N_3362,N_1719,N_814);
and U3363 (N_3363,N_1625,N_556);
nand U3364 (N_3364,N_1254,N_1684);
or U3365 (N_3365,N_177,N_429);
or U3366 (N_3366,N_1296,N_1480);
xnor U3367 (N_3367,N_1330,N_1715);
nor U3368 (N_3368,N_2072,N_2948);
xor U3369 (N_3369,N_785,N_797);
nand U3370 (N_3370,N_617,N_2083);
or U3371 (N_3371,N_923,N_221);
nand U3372 (N_3372,N_2631,N_2718);
nor U3373 (N_3373,N_2694,N_2869);
or U3374 (N_3374,N_868,N_2752);
nand U3375 (N_3375,N_2438,N_1053);
nor U3376 (N_3376,N_2451,N_1203);
nor U3377 (N_3377,N_1391,N_45);
and U3378 (N_3378,N_943,N_1641);
xnor U3379 (N_3379,N_2859,N_1442);
nand U3380 (N_3380,N_1431,N_1632);
nor U3381 (N_3381,N_1950,N_1600);
xnor U3382 (N_3382,N_394,N_2063);
or U3383 (N_3383,N_300,N_21);
nor U3384 (N_3384,N_1983,N_284);
xor U3385 (N_3385,N_823,N_1358);
nor U3386 (N_3386,N_2810,N_1441);
or U3387 (N_3387,N_2557,N_1991);
xnor U3388 (N_3388,N_2708,N_1702);
xor U3389 (N_3389,N_2091,N_1542);
or U3390 (N_3390,N_1577,N_2303);
nor U3391 (N_3391,N_626,N_2384);
or U3392 (N_3392,N_2971,N_1711);
nand U3393 (N_3393,N_1980,N_1935);
xor U3394 (N_3394,N_757,N_292);
and U3395 (N_3395,N_1530,N_2160);
nand U3396 (N_3396,N_2677,N_1445);
xnor U3397 (N_3397,N_1814,N_3087);
or U3398 (N_3398,N_2282,N_2483);
nand U3399 (N_3399,N_1452,N_2750);
xnor U3400 (N_3400,N_524,N_1877);
and U3401 (N_3401,N_2165,N_2928);
nor U3402 (N_3402,N_817,N_3052);
xnor U3403 (N_3403,N_2981,N_1876);
nand U3404 (N_3404,N_3015,N_414);
or U3405 (N_3405,N_1273,N_806);
nor U3406 (N_3406,N_1258,N_1644);
and U3407 (N_3407,N_1428,N_1566);
nand U3408 (N_3408,N_1389,N_2522);
nand U3409 (N_3409,N_3028,N_2820);
and U3410 (N_3410,N_1661,N_32);
nand U3411 (N_3411,N_161,N_1884);
xor U3412 (N_3412,N_1156,N_1225);
and U3413 (N_3413,N_1796,N_1107);
nor U3414 (N_3414,N_2635,N_2967);
nand U3415 (N_3415,N_2571,N_1864);
nand U3416 (N_3416,N_481,N_580);
or U3417 (N_3417,N_2854,N_2943);
xor U3418 (N_3418,N_2111,N_2183);
or U3419 (N_3419,N_2293,N_2115);
nor U3420 (N_3420,N_384,N_2753);
nor U3421 (N_3421,N_2439,N_1354);
xnor U3422 (N_3422,N_764,N_2689);
nand U3423 (N_3423,N_1837,N_1968);
nor U3424 (N_3424,N_2847,N_2994);
and U3425 (N_3425,N_44,N_2776);
nor U3426 (N_3426,N_786,N_2904);
and U3427 (N_3427,N_1553,N_721);
and U3428 (N_3428,N_1663,N_1739);
nand U3429 (N_3429,N_2767,N_1364);
and U3430 (N_3430,N_1185,N_800);
and U3431 (N_3431,N_422,N_766);
nand U3432 (N_3432,N_2717,N_140);
nand U3433 (N_3433,N_882,N_2068);
nor U3434 (N_3434,N_3062,N_1126);
nand U3435 (N_3435,N_476,N_2883);
nand U3436 (N_3436,N_33,N_357);
and U3437 (N_3437,N_1473,N_2919);
nor U3438 (N_3438,N_2851,N_1698);
nand U3439 (N_3439,N_82,N_50);
nor U3440 (N_3440,N_2611,N_2478);
xor U3441 (N_3441,N_2145,N_732);
or U3442 (N_3442,N_1874,N_705);
xnor U3443 (N_3443,N_2258,N_455);
nand U3444 (N_3444,N_984,N_1106);
nor U3445 (N_3445,N_1891,N_1454);
and U3446 (N_3446,N_1064,N_2263);
or U3447 (N_3447,N_1052,N_1448);
nand U3448 (N_3448,N_1730,N_2127);
nand U3449 (N_3449,N_1013,N_363);
nor U3450 (N_3450,N_2138,N_1859);
nor U3451 (N_3451,N_1782,N_366);
xor U3452 (N_3452,N_1040,N_2836);
and U3453 (N_3453,N_1423,N_825);
nor U3454 (N_3454,N_589,N_2837);
or U3455 (N_3455,N_339,N_2645);
nand U3456 (N_3456,N_1949,N_147);
or U3457 (N_3457,N_1602,N_887);
or U3458 (N_3458,N_881,N_319);
nor U3459 (N_3459,N_1253,N_315);
or U3460 (N_3460,N_2844,N_755);
nor U3461 (N_3461,N_336,N_2764);
nand U3462 (N_3462,N_1434,N_2756);
nor U3463 (N_3463,N_1074,N_912);
or U3464 (N_3464,N_3096,N_2308);
and U3465 (N_3465,N_3120,N_2347);
xnor U3466 (N_3466,N_215,N_2080);
nand U3467 (N_3467,N_2982,N_1154);
nand U3468 (N_3468,N_1992,N_3021);
nor U3469 (N_3469,N_1592,N_1734);
nor U3470 (N_3470,N_3097,N_553);
nand U3471 (N_3471,N_496,N_2873);
or U3472 (N_3472,N_1844,N_1505);
xnor U3473 (N_3473,N_776,N_1102);
and U3474 (N_3474,N_582,N_1009);
nand U3475 (N_3475,N_1117,N_1725);
nand U3476 (N_3476,N_2806,N_2561);
or U3477 (N_3477,N_962,N_1616);
xnor U3478 (N_3478,N_2426,N_2101);
xnor U3479 (N_3479,N_1601,N_2591);
nor U3480 (N_3480,N_1907,N_685);
and U3481 (N_3481,N_3111,N_2235);
or U3482 (N_3482,N_1249,N_178);
xnor U3483 (N_3483,N_1845,N_1137);
nand U3484 (N_3484,N_1771,N_1676);
xor U3485 (N_3485,N_1395,N_261);
nand U3486 (N_3486,N_2144,N_2709);
nor U3487 (N_3487,N_2445,N_398);
and U3488 (N_3488,N_2898,N_379);
xor U3489 (N_3489,N_1783,N_3082);
xor U3490 (N_3490,N_2017,N_1748);
xnor U3491 (N_3491,N_2301,N_1823);
nor U3492 (N_3492,N_457,N_1540);
and U3493 (N_3493,N_2733,N_1525);
nand U3494 (N_3494,N_1063,N_174);
nor U3495 (N_3495,N_1100,N_1780);
and U3496 (N_3496,N_16,N_2619);
nand U3497 (N_3497,N_143,N_910);
or U3498 (N_3498,N_841,N_2995);
nor U3499 (N_3499,N_3116,N_1882);
nand U3500 (N_3500,N_3041,N_1245);
xor U3501 (N_3501,N_1797,N_188);
or U3502 (N_3502,N_581,N_1155);
xor U3503 (N_3503,N_2654,N_1500);
nor U3504 (N_3504,N_1016,N_2046);
or U3505 (N_3505,N_1627,N_2122);
or U3506 (N_3506,N_1712,N_1161);
nand U3507 (N_3507,N_2085,N_3023);
or U3508 (N_3508,N_9,N_1490);
nand U3509 (N_3509,N_406,N_54);
xnor U3510 (N_3510,N_166,N_2218);
or U3511 (N_3511,N_975,N_3078);
or U3512 (N_3512,N_515,N_1701);
nand U3513 (N_3513,N_692,N_688);
nor U3514 (N_3514,N_1437,N_2899);
xnor U3515 (N_3515,N_2918,N_1190);
xnor U3516 (N_3516,N_1682,N_2914);
nor U3517 (N_3517,N_2908,N_1924);
or U3518 (N_3518,N_664,N_155);
nor U3519 (N_3519,N_2876,N_22);
and U3520 (N_3520,N_839,N_2628);
xor U3521 (N_3521,N_1871,N_1422);
and U3522 (N_3522,N_574,N_2788);
or U3523 (N_3523,N_815,N_97);
nand U3524 (N_3524,N_1214,N_1328);
or U3525 (N_3525,N_1370,N_896);
and U3526 (N_3526,N_3004,N_1956);
xor U3527 (N_3527,N_511,N_1321);
nor U3528 (N_3528,N_2180,N_430);
or U3529 (N_3529,N_973,N_2087);
and U3530 (N_3530,N_865,N_2255);
nor U3531 (N_3531,N_335,N_289);
and U3532 (N_3532,N_2625,N_2413);
nand U3533 (N_3533,N_3071,N_693);
xor U3534 (N_3534,N_2580,N_1580);
and U3535 (N_3535,N_947,N_518);
nand U3536 (N_3536,N_1244,N_703);
or U3537 (N_3537,N_1832,N_1917);
nor U3538 (N_3538,N_426,N_2675);
or U3539 (N_3539,N_1150,N_451);
nand U3540 (N_3540,N_743,N_1629);
nor U3541 (N_3541,N_965,N_1140);
nor U3542 (N_3542,N_2855,N_713);
or U3543 (N_3543,N_2378,N_583);
nand U3544 (N_3544,N_1869,N_182);
nand U3545 (N_3545,N_2174,N_2444);
and U3546 (N_3546,N_63,N_940);
and U3547 (N_3547,N_2435,N_205);
nand U3548 (N_3548,N_1918,N_2274);
nor U3549 (N_3549,N_1948,N_850);
nor U3550 (N_3550,N_578,N_2366);
nand U3551 (N_3551,N_1290,N_244);
xor U3552 (N_3552,N_2599,N_250);
nor U3553 (N_3553,N_2606,N_1800);
xnor U3554 (N_3554,N_2595,N_314);
nor U3555 (N_3555,N_1509,N_2618);
xnor U3556 (N_3556,N_1614,N_2671);
and U3557 (N_3557,N_1953,N_1951);
and U3558 (N_3558,N_863,N_7);
xor U3559 (N_3559,N_1791,N_276);
xnor U3560 (N_3560,N_1099,N_862);
or U3561 (N_3561,N_1329,N_842);
nand U3562 (N_3562,N_820,N_1331);
nor U3563 (N_3563,N_1848,N_197);
nand U3564 (N_3564,N_2437,N_1872);
xnor U3565 (N_3565,N_832,N_1754);
or U3566 (N_3566,N_397,N_1733);
nor U3567 (N_3567,N_1545,N_2412);
nor U3568 (N_3568,N_2375,N_768);
xor U3569 (N_3569,N_1759,N_2511);
or U3570 (N_3570,N_2804,N_3080);
nand U3571 (N_3571,N_2358,N_412);
and U3572 (N_3572,N_548,N_1518);
xnor U3573 (N_3573,N_2786,N_2862);
nor U3574 (N_3574,N_2335,N_564);
xnor U3575 (N_3575,N_2140,N_784);
nand U3576 (N_3576,N_1359,N_2596);
nand U3577 (N_3577,N_1377,N_1234);
or U3578 (N_3578,N_3045,N_2265);
or U3579 (N_3579,N_2617,N_1830);
or U3580 (N_3580,N_1908,N_1861);
nor U3581 (N_3581,N_2433,N_2231);
nor U3582 (N_3582,N_38,N_1041);
xnor U3583 (N_3583,N_2012,N_1210);
and U3584 (N_3584,N_25,N_2958);
nand U3585 (N_3585,N_1938,N_1945);
xor U3586 (N_3586,N_2835,N_472);
xor U3587 (N_3587,N_1557,N_1893);
nand U3588 (N_3588,N_828,N_2359);
xnor U3589 (N_3589,N_1963,N_1315);
or U3590 (N_3590,N_927,N_2704);
and U3591 (N_3591,N_2015,N_399);
nand U3592 (N_3592,N_1095,N_931);
nor U3593 (N_3593,N_616,N_1192);
and U3594 (N_3594,N_2629,N_623);
nor U3595 (N_3595,N_3039,N_2442);
xnor U3596 (N_3596,N_2177,N_1875);
nand U3597 (N_3597,N_2053,N_268);
or U3598 (N_3598,N_1420,N_2990);
nor U3599 (N_3599,N_990,N_2295);
or U3600 (N_3600,N_1471,N_2333);
xor U3601 (N_3601,N_1648,N_1114);
xor U3602 (N_3602,N_23,N_2228);
and U3603 (N_3603,N_1982,N_911);
xnor U3604 (N_3604,N_1880,N_2465);
nor U3605 (N_3605,N_2748,N_483);
and U3606 (N_3606,N_1351,N_2233);
or U3607 (N_3607,N_352,N_1282);
nor U3608 (N_3608,N_1519,N_40);
and U3609 (N_3609,N_2408,N_630);
nor U3610 (N_3610,N_2864,N_1958);
xor U3611 (N_3611,N_2207,N_1200);
and U3612 (N_3612,N_2076,N_1236);
nand U3613 (N_3613,N_2229,N_1355);
xor U3614 (N_3614,N_2801,N_607);
nand U3615 (N_3615,N_720,N_1786);
nor U3616 (N_3616,N_480,N_770);
or U3617 (N_3617,N_2734,N_1957);
nor U3618 (N_3618,N_291,N_663);
nand U3619 (N_3619,N_1342,N_1115);
nor U3620 (N_3620,N_2616,N_1174);
and U3621 (N_3621,N_2882,N_913);
or U3622 (N_3622,N_1717,N_1596);
or U3623 (N_3623,N_1892,N_1611);
nor U3624 (N_3624,N_930,N_407);
or U3625 (N_3625,N_456,N_453);
nor U3626 (N_3626,N_164,N_2781);
xor U3627 (N_3627,N_1578,N_1476);
nand U3628 (N_3628,N_1045,N_641);
xor U3629 (N_3629,N_2418,N_3099);
nor U3630 (N_3630,N_2774,N_920);
nand U3631 (N_3631,N_3088,N_2498);
nand U3632 (N_3632,N_1504,N_138);
or U3633 (N_3633,N_2468,N_2150);
nand U3634 (N_3634,N_3090,N_2322);
xnor U3635 (N_3635,N_1923,N_1129);
nor U3636 (N_3636,N_902,N_2807);
nand U3637 (N_3637,N_1427,N_473);
or U3638 (N_3638,N_718,N_1247);
nor U3639 (N_3639,N_1533,N_1726);
nand U3640 (N_3640,N_2749,N_1319);
and U3641 (N_3641,N_1493,N_710);
nand U3642 (N_3642,N_1043,N_301);
nor U3643 (N_3643,N_2540,N_2812);
nand U3644 (N_3644,N_1460,N_1570);
and U3645 (N_3645,N_2309,N_2428);
or U3646 (N_3646,N_596,N_37);
nor U3647 (N_3647,N_199,N_1218);
nor U3648 (N_3648,N_129,N_2641);
and U3649 (N_3649,N_450,N_816);
nand U3650 (N_3650,N_1667,N_633);
and U3651 (N_3651,N_1350,N_118);
or U3652 (N_3652,N_1037,N_922);
xor U3653 (N_3653,N_2779,N_2455);
or U3654 (N_3654,N_780,N_2380);
or U3655 (N_3655,N_2738,N_489);
or U3656 (N_3656,N_2706,N_2666);
nand U3657 (N_3657,N_1101,N_1967);
and U3658 (N_3658,N_2487,N_2818);
nor U3659 (N_3659,N_3051,N_748);
and U3660 (N_3660,N_572,N_1191);
nand U3661 (N_3661,N_1850,N_202);
nor U3662 (N_3662,N_1686,N_945);
xnor U3663 (N_3663,N_1603,N_1527);
xor U3664 (N_3664,N_1252,N_948);
or U3665 (N_3665,N_1487,N_2946);
nand U3666 (N_3666,N_2761,N_689);
and U3667 (N_3667,N_2431,N_1118);
nand U3668 (N_3668,N_2890,N_2823);
nor U3669 (N_3669,N_327,N_2208);
nand U3670 (N_3670,N_2952,N_2473);
or U3671 (N_3671,N_68,N_275);
or U3672 (N_3672,N_2660,N_758);
or U3673 (N_3673,N_2860,N_796);
xor U3674 (N_3674,N_2298,N_1231);
nand U3675 (N_3675,N_904,N_2798);
nand U3676 (N_3676,N_2612,N_2397);
nor U3677 (N_3677,N_2372,N_2288);
nor U3678 (N_3678,N_2777,N_1365);
and U3679 (N_3679,N_497,N_3072);
xnor U3680 (N_3680,N_1628,N_762);
and U3681 (N_3681,N_1011,N_1607);
and U3682 (N_3682,N_1581,N_2555);
and U3683 (N_3683,N_640,N_2519);
xnor U3684 (N_3684,N_2332,N_340);
and U3685 (N_3685,N_2021,N_2998);
or U3686 (N_3686,N_1149,N_2551);
and U3687 (N_3687,N_193,N_3123);
xor U3688 (N_3688,N_2663,N_310);
nor U3689 (N_3689,N_248,N_544);
or U3690 (N_3690,N_539,N_638);
nand U3691 (N_3691,N_334,N_2422);
xor U3692 (N_3692,N_1289,N_1562);
or U3693 (N_3693,N_566,N_370);
and U3694 (N_3694,N_1400,N_959);
nor U3695 (N_3695,N_2537,N_1397);
nor U3696 (N_3696,N_592,N_1680);
or U3697 (N_3697,N_1322,N_3057);
or U3698 (N_3698,N_2661,N_871);
nand U3699 (N_3699,N_2827,N_2740);
nor U3700 (N_3700,N_2874,N_1709);
and U3701 (N_3701,N_254,N_2116);
xor U3702 (N_3702,N_730,N_2633);
nand U3703 (N_3703,N_2881,N_1595);
nand U3704 (N_3704,N_1023,N_728);
and U3705 (N_3705,N_2163,N_2392);
xnor U3706 (N_3706,N_2896,N_345);
and U3707 (N_3707,N_2283,N_228);
nand U3708 (N_3708,N_2023,N_2868);
nand U3709 (N_3709,N_318,N_649);
nand U3710 (N_3710,N_2699,N_1057);
nor U3711 (N_3711,N_794,N_752);
nor U3712 (N_3712,N_2547,N_586);
nand U3713 (N_3713,N_1307,N_2188);
nor U3714 (N_3714,N_2351,N_3086);
nand U3715 (N_3715,N_368,N_113);
and U3716 (N_3716,N_1120,N_287);
nand U3717 (N_3717,N_1820,N_1668);
xnor U3718 (N_3718,N_1828,N_170);
xnor U3719 (N_3719,N_1070,N_1511);
or U3720 (N_3720,N_2220,N_2760);
xor U3721 (N_3721,N_1146,N_64);
nand U3722 (N_3722,N_2137,N_526);
nand U3723 (N_3723,N_2172,N_1018);
nor U3724 (N_3724,N_1461,N_1325);
nor U3725 (N_3725,N_2075,N_2710);
or U3726 (N_3726,N_928,N_1105);
nand U3727 (N_3727,N_30,N_2736);
and U3728 (N_3728,N_2135,N_423);
nor U3729 (N_3729,N_12,N_19);
xor U3730 (N_3730,N_2497,N_337);
nand U3731 (N_3731,N_636,N_1821);
and U3732 (N_3732,N_151,N_988);
or U3733 (N_3733,N_821,N_1903);
xor U3734 (N_3734,N_2313,N_2712);
nor U3735 (N_3735,N_1897,N_978);
nor U3736 (N_3736,N_341,N_2314);
or U3737 (N_3737,N_2843,N_478);
nand U3738 (N_3738,N_2634,N_2037);
or U3739 (N_3739,N_1001,N_1656);
xnor U3740 (N_3740,N_3018,N_3050);
and U3741 (N_3741,N_1744,N_672);
nor U3742 (N_3742,N_1973,N_2598);
nand U3743 (N_3743,N_3104,N_2884);
or U3744 (N_3744,N_646,N_2797);
nand U3745 (N_3745,N_1683,N_210);
xor U3746 (N_3746,N_2535,N_1246);
nand U3747 (N_3747,N_2545,N_2379);
or U3748 (N_3748,N_216,N_2421);
and U3749 (N_3749,N_1337,N_479);
and U3750 (N_3750,N_2722,N_2825);
xor U3751 (N_3751,N_1213,N_2583);
nand U3752 (N_3752,N_1004,N_2484);
xor U3753 (N_3753,N_2132,N_2939);
xnor U3754 (N_3754,N_1116,N_1765);
and U3755 (N_3755,N_2977,N_3069);
and U3756 (N_3756,N_1896,N_441);
or U3757 (N_3757,N_2337,N_1887);
nand U3758 (N_3758,N_2667,N_1716);
xor U3759 (N_3759,N_421,N_2893);
nand U3760 (N_3760,N_1763,N_1250);
and U3761 (N_3761,N_704,N_783);
nor U3762 (N_3762,N_792,N_1606);
nand U3763 (N_3763,N_1048,N_560);
and U3764 (N_3764,N_2416,N_647);
xor U3765 (N_3765,N_1732,N_1274);
xnor U3766 (N_3766,N_2942,N_1776);
nor U3767 (N_3767,N_1555,N_1610);
nand U3768 (N_3768,N_2153,N_84);
or U3769 (N_3769,N_2167,N_1546);
and U3770 (N_3770,N_2932,N_537);
or U3771 (N_3771,N_2441,N_2399);
xor U3772 (N_3772,N_1489,N_2044);
nand U3773 (N_3773,N_2028,N_74);
xnor U3774 (N_3774,N_1166,N_857);
xnor U3775 (N_3775,N_2008,N_1007);
nor U3776 (N_3776,N_983,N_2850);
and U3777 (N_3777,N_719,N_477);
nor U3778 (N_3778,N_587,N_2791);
nand U3779 (N_3779,N_1804,N_2324);
nor U3780 (N_3780,N_2490,N_3);
or U3781 (N_3781,N_2613,N_434);
or U3782 (N_3782,N_756,N_2621);
and U3783 (N_3783,N_3084,N_1209);
nand U3784 (N_3784,N_152,N_2772);
nor U3785 (N_3785,N_3014,N_1270);
nand U3786 (N_3786,N_262,N_1005);
and U3787 (N_3787,N_2503,N_100);
or U3788 (N_3788,N_3094,N_36);
or U3789 (N_3789,N_1271,N_1827);
or U3790 (N_3790,N_2463,N_836);
or U3791 (N_3791,N_624,N_2539);
nand U3792 (N_3792,N_2902,N_2275);
nand U3793 (N_3793,N_2329,N_2682);
or U3794 (N_3794,N_594,N_2030);
and U3795 (N_3795,N_749,N_2056);
nor U3796 (N_3796,N_1132,N_621);
nand U3797 (N_3797,N_908,N_2261);
nor U3798 (N_3798,N_2566,N_490);
or U3799 (N_3799,N_117,N_1368);
nor U3800 (N_3800,N_1008,N_1241);
nor U3801 (N_3801,N_1846,N_391);
xnor U3802 (N_3802,N_3124,N_848);
and U3803 (N_3803,N_869,N_459);
or U3804 (N_3804,N_2202,N_76);
and U3805 (N_3805,N_1652,N_1620);
or U3806 (N_3806,N_2000,N_529);
and U3807 (N_3807,N_2650,N_2584);
nor U3808 (N_3808,N_2920,N_835);
or U3809 (N_3809,N_2510,N_1879);
nor U3810 (N_3810,N_1,N_725);
and U3811 (N_3811,N_1310,N_2848);
and U3812 (N_3812,N_2742,N_1649);
nand U3813 (N_3813,N_3083,N_231);
xnor U3814 (N_3814,N_1781,N_2370);
or U3815 (N_3815,N_2789,N_2496);
xnor U3816 (N_3816,N_2154,N_1729);
or U3817 (N_3817,N_2615,N_2560);
and U3818 (N_3818,N_2590,N_2086);
and U3819 (N_3819,N_789,N_1027);
and U3820 (N_3820,N_822,N_2194);
nor U3821 (N_3821,N_2373,N_380);
and U3822 (N_3822,N_1145,N_66);
nand U3823 (N_3823,N_2714,N_329);
nand U3824 (N_3824,N_2252,N_2575);
nor U3825 (N_3825,N_2011,N_2327);
xnor U3826 (N_3826,N_1412,N_298);
xnor U3827 (N_3827,N_259,N_2338);
and U3828 (N_3828,N_723,N_1708);
xor U3829 (N_3829,N_433,N_1779);
nand U3830 (N_3830,N_1293,N_2209);
nor U3831 (N_3831,N_1816,N_2270);
or U3832 (N_3832,N_1467,N_771);
or U3833 (N_3833,N_1179,N_1089);
xnor U3834 (N_3834,N_1554,N_3016);
and U3835 (N_3835,N_891,N_2815);
and U3836 (N_3836,N_1160,N_503);
xnor U3837 (N_3837,N_2186,N_2953);
or U3838 (N_3838,N_1151,N_1408);
or U3839 (N_3839,N_819,N_2082);
xor U3840 (N_3840,N_3003,N_154);
xor U3841 (N_3841,N_2205,N_2989);
nor U3842 (N_3842,N_2257,N_2688);
nand U3843 (N_3843,N_242,N_545);
nand U3844 (N_3844,N_2148,N_629);
xor U3845 (N_3845,N_39,N_964);
and U3846 (N_3846,N_258,N_3020);
xnor U3847 (N_3847,N_2236,N_998);
or U3848 (N_3848,N_2954,N_220);
nand U3849 (N_3849,N_219,N_58);
nor U3850 (N_3850,N_86,N_2224);
nor U3851 (N_3851,N_1483,N_48);
nand U3852 (N_3852,N_2656,N_1932);
xor U3853 (N_3853,N_494,N_3119);
and U3854 (N_3854,N_1032,N_2763);
nand U3855 (N_3855,N_2702,N_110);
nor U3856 (N_3856,N_347,N_120);
xnor U3857 (N_3857,N_1760,N_290);
nor U3858 (N_3858,N_953,N_42);
nand U3859 (N_3859,N_996,N_655);
and U3860 (N_3860,N_1758,N_2264);
nor U3861 (N_3861,N_3085,N_364);
or U3862 (N_3862,N_2244,N_1901);
or U3863 (N_3863,N_697,N_1123);
or U3864 (N_3864,N_1604,N_1793);
or U3865 (N_3865,N_2532,N_2526);
or U3866 (N_3866,N_805,N_712);
and U3867 (N_3867,N_1002,N_1086);
and U3868 (N_3868,N_1175,N_390);
nor U3869 (N_3869,N_2374,N_2466);
nand U3870 (N_3870,N_1718,N_2222);
xor U3871 (N_3871,N_2906,N_810);
or U3872 (N_3872,N_2731,N_388);
xor U3873 (N_3873,N_1507,N_1108);
and U3874 (N_3874,N_2960,N_2732);
nand U3875 (N_3875,N_1921,N_2315);
and U3876 (N_3876,N_2912,N_707);
nand U3877 (N_3877,N_1998,N_2917);
xor U3878 (N_3878,N_1589,N_1303);
xnor U3879 (N_3879,N_410,N_1650);
nand U3880 (N_3880,N_2940,N_1305);
or U3881 (N_3881,N_1978,N_813);
nor U3882 (N_3882,N_157,N_1065);
xnor U3883 (N_3883,N_844,N_306);
nand U3884 (N_3884,N_2446,N_1608);
or U3885 (N_3885,N_1194,N_2081);
and U3886 (N_3886,N_999,N_2430);
and U3887 (N_3887,N_2394,N_504);
nor U3888 (N_3888,N_2711,N_3095);
or U3889 (N_3889,N_392,N_2991);
nor U3890 (N_3890,N_232,N_2588);
or U3891 (N_3891,N_2052,N_2589);
and U3892 (N_3892,N_361,N_1721);
nor U3893 (N_3893,N_233,N_1425);
nand U3894 (N_3894,N_1163,N_971);
nor U3895 (N_3895,N_1934,N_2665);
nand U3896 (N_3896,N_360,N_2250);
nor U3897 (N_3897,N_2771,N_2980);
or U3898 (N_3898,N_585,N_1692);
nand U3899 (N_3899,N_1311,N_929);
xor U3900 (N_3900,N_2659,N_2004);
and U3901 (N_3901,N_543,N_1528);
nand U3902 (N_3902,N_3031,N_1069);
or U3903 (N_3903,N_127,N_1582);
xnor U3904 (N_3904,N_374,N_1637);
and U3905 (N_3905,N_735,N_2929);
or U3906 (N_3906,N_2947,N_2096);
or U3907 (N_3907,N_2355,N_2649);
nand U3908 (N_3908,N_2467,N_2834);
xor U3909 (N_3909,N_1984,N_2938);
and U3910 (N_3910,N_2701,N_2363);
xnor U3911 (N_3911,N_351,N_35);
or U3912 (N_3912,N_2067,N_2670);
or U3913 (N_3913,N_114,N_1088);
nor U3914 (N_3914,N_1288,N_299);
xor U3915 (N_3915,N_2513,N_1750);
nor U3916 (N_3916,N_1583,N_2997);
nor U3917 (N_3917,N_562,N_802);
and U3918 (N_3918,N_2987,N_94);
or U3919 (N_3919,N_1634,N_837);
and U3920 (N_3920,N_818,N_1376);
and U3921 (N_3921,N_2574,N_2969);
nand U3922 (N_3922,N_1299,N_2573);
nor U3923 (N_3923,N_1281,N_1111);
xnor U3924 (N_3924,N_2719,N_2604);
and U3925 (N_3925,N_1599,N_3046);
xnor U3926 (N_3926,N_2006,N_126);
nor U3927 (N_3927,N_2744,N_1349);
nand U3928 (N_3928,N_2729,N_1979);
nand U3929 (N_3929,N_2271,N_425);
nand U3930 (N_3930,N_2925,N_2543);
and U3931 (N_3931,N_1514,N_2090);
xor U3932 (N_3932,N_1997,N_1183);
nand U3933 (N_3933,N_1345,N_746);
nor U3934 (N_3934,N_2212,N_2406);
nor U3935 (N_3935,N_2273,N_1535);
nand U3936 (N_3936,N_1690,N_527);
or U3937 (N_3937,N_1380,N_1927);
nor U3938 (N_3938,N_2369,N_227);
and U3939 (N_3939,N_516,N_2272);
nor U3940 (N_3940,N_864,N_870);
and U3941 (N_3941,N_2770,N_1675);
and U3942 (N_3942,N_2927,N_1078);
nor U3943 (N_3943,N_2149,N_2909);
nand U3944 (N_3944,N_2470,N_2125);
nor U3945 (N_3945,N_377,N_2973);
nand U3946 (N_3946,N_2559,N_1588);
or U3947 (N_3947,N_2849,N_2891);
nor U3948 (N_3948,N_980,N_1168);
nor U3949 (N_3949,N_3049,N_1906);
xor U3950 (N_3950,N_13,N_236);
and U3951 (N_3951,N_866,N_2155);
and U3952 (N_3952,N_2690,N_716);
and U3953 (N_3953,N_46,N_1515);
and U3954 (N_3954,N_781,N_2162);
nor U3955 (N_3955,N_2010,N_2905);
xor U3956 (N_3956,N_83,N_3009);
and U3957 (N_3957,N_251,N_1752);
xnor U3958 (N_3958,N_2107,N_1833);
nor U3959 (N_3959,N_2320,N_2460);
and U3960 (N_3960,N_1735,N_2813);
or U3961 (N_3961,N_2300,N_546);
or U3962 (N_3962,N_1055,N_2766);
nor U3963 (N_3963,N_1849,N_2034);
nor U3964 (N_3964,N_1072,N_326);
xnor U3965 (N_3965,N_2092,N_415);
nor U3966 (N_3966,N_2472,N_977);
and U3967 (N_3967,N_1333,N_2401);
xnor U3968 (N_3968,N_2398,N_1196);
nand U3969 (N_3969,N_1727,N_1839);
xor U3970 (N_3970,N_1677,N_2858);
or U3971 (N_3971,N_2669,N_2432);
nand U3972 (N_3972,N_1167,N_47);
nor U3973 (N_3973,N_1014,N_2074);
nor U3974 (N_3974,N_2568,N_3109);
nor U3975 (N_3975,N_1153,N_634);
or U3976 (N_3976,N_2387,N_1856);
or U3977 (N_3977,N_2325,N_1478);
or U3978 (N_3978,N_2494,N_2974);
nand U3979 (N_3979,N_851,N_2031);
nand U3980 (N_3980,N_264,N_950);
or U3981 (N_3981,N_777,N_2395);
xor U3982 (N_3982,N_1083,N_373);
nor U3983 (N_3983,N_662,N_131);
nor U3984 (N_3984,N_2949,N_1257);
nor U3985 (N_3985,N_1537,N_1558);
nand U3986 (N_3986,N_181,N_1176);
or U3987 (N_3987,N_994,N_2486);
xnor U3988 (N_3988,N_1593,N_115);
and U3989 (N_3989,N_2130,N_2889);
xnor U3990 (N_3990,N_2979,N_652);
or U3991 (N_3991,N_2886,N_253);
nor U3992 (N_3992,N_601,N_125);
nor U3993 (N_3993,N_333,N_2558);
nand U3994 (N_3994,N_614,N_2735);
and U3995 (N_3995,N_1999,N_1853);
xnor U3996 (N_3996,N_1399,N_1995);
and U3997 (N_3997,N_1170,N_1736);
nor U3998 (N_3998,N_2725,N_1382);
nand U3999 (N_3999,N_2723,N_2585);
or U4000 (N_4000,N_283,N_2550);
and U4001 (N_4001,N_657,N_803);
nand U4002 (N_4002,N_1878,N_2396);
nor U4003 (N_4003,N_2841,N_1366);
and U4004 (N_4004,N_1312,N_1749);
nand U4005 (N_4005,N_2383,N_163);
or U4006 (N_4006,N_2326,N_1549);
nor U4007 (N_4007,N_2515,N_2097);
or U4008 (N_4008,N_2608,N_1042);
xnor U4009 (N_4009,N_939,N_635);
xor U4010 (N_4010,N_2253,N_1393);
and U4011 (N_4011,N_1085,N_2696);
nand U4012 (N_4012,N_2523,N_2533);
nor U4013 (N_4013,N_405,N_438);
or U4014 (N_4014,N_3002,N_2691);
and U4015 (N_4015,N_1010,N_2479);
nor U4016 (N_4016,N_1226,N_1747);
nor U4017 (N_4017,N_1785,N_895);
nand U4018 (N_4018,N_502,N_2102);
xor U4019 (N_4019,N_2334,N_1928);
nor U4020 (N_4020,N_698,N_799);
or U4021 (N_4021,N_1657,N_10);
xor U4022 (N_4022,N_2377,N_2013);
nor U4023 (N_4023,N_2247,N_2549);
nor U4024 (N_4024,N_637,N_1722);
nor U4025 (N_4025,N_763,N_2210);
nor U4026 (N_4026,N_1324,N_1418);
nand U4027 (N_4027,N_597,N_2318);
or U4028 (N_4028,N_1694,N_1339);
and U4029 (N_4029,N_979,N_350);
nand U4030 (N_4030,N_2312,N_650);
xnor U4031 (N_4031,N_396,N_168);
and U4032 (N_4032,N_222,N_691);
or U4033 (N_4033,N_1097,N_2341);
and U4034 (N_4034,N_2036,N_1789);
nand U4035 (N_4035,N_2189,N_1761);
nor U4036 (N_4036,N_1187,N_27);
nor U4037 (N_4037,N_613,N_951);
or U4038 (N_4038,N_3011,N_639);
xor U4039 (N_4039,N_71,N_2697);
nand U4040 (N_4040,N_2400,N_2305);
xnor U4041 (N_4041,N_60,N_753);
xor U4042 (N_4042,N_1082,N_2576);
or U4043 (N_4043,N_1506,N_1030);
or U4044 (N_4044,N_2381,N_1939);
nand U4045 (N_4045,N_2246,N_2181);
or U4046 (N_4046,N_2331,N_1713);
or U4047 (N_4047,N_95,N_1148);
nor U4048 (N_4048,N_907,N_2819);
xor U4049 (N_4049,N_714,N_1029);
or U4050 (N_4050,N_1409,N_256);
nand U4051 (N_4051,N_2992,N_2651);
nor U4052 (N_4052,N_1237,N_404);
and U4053 (N_4053,N_2453,N_3037);
nor U4054 (N_4054,N_296,N_1633);
and U4055 (N_4055,N_2700,N_1443);
and U4056 (N_4056,N_1857,N_2693);
xnor U4057 (N_4057,N_346,N_1819);
or U4058 (N_4058,N_444,N_1913);
and U4059 (N_4059,N_1774,N_1681);
nand U4060 (N_4060,N_3076,N_3113);
xnor U4061 (N_4061,N_550,N_499);
and U4062 (N_4062,N_134,N_2323);
nor U4063 (N_4063,N_602,N_1916);
xnor U4064 (N_4064,N_2643,N_2390);
xnor U4065 (N_4065,N_2071,N_849);
or U4066 (N_4066,N_3061,N_522);
nor U4067 (N_4067,N_1810,N_2586);
nor U4068 (N_4068,N_760,N_3058);
nand U4069 (N_4069,N_1851,N_612);
or U4070 (N_4070,N_3075,N_2597);
and U4071 (N_4071,N_569,N_1216);
or U4072 (N_4072,N_89,N_2730);
and U4073 (N_4073,N_2951,N_1621);
nand U4074 (N_4074,N_1195,N_2106);
or U4075 (N_4075,N_1091,N_69);
xor U4076 (N_4076,N_493,N_1215);
xnor U4077 (N_4077,N_2512,N_523);
nand U4078 (N_4078,N_162,N_2936);
nand U4079 (N_4079,N_1497,N_332);
or U4080 (N_4080,N_2447,N_317);
nand U4081 (N_4081,N_2114,N_1334);
xnor U4082 (N_4082,N_1598,N_956);
or U4083 (N_4083,N_2243,N_2664);
xor U4084 (N_4084,N_559,N_2289);
and U4085 (N_4085,N_903,N_793);
nor U4086 (N_4086,N_952,N_2720);
xor U4087 (N_4087,N_2223,N_610);
or U4088 (N_4088,N_2307,N_1551);
or U4089 (N_4089,N_1327,N_1679);
xor U4090 (N_4090,N_2237,N_653);
nand U4091 (N_4091,N_2009,N_874);
nand U4092 (N_4092,N_671,N_1741);
or U4093 (N_4093,N_2060,N_180);
or U4094 (N_4094,N_214,N_509);
nand U4095 (N_4095,N_1469,N_3038);
and U4096 (N_4096,N_1597,N_2986);
nor U4097 (N_4097,N_2592,N_452);
xor U4098 (N_4098,N_1294,N_970);
nor U4099 (N_4099,N_761,N_2362);
nor U4100 (N_4100,N_3013,N_158);
and U4101 (N_4101,N_1494,N_2050);
nand U4102 (N_4102,N_1306,N_1484);
xnor U4103 (N_4103,N_1658,N_2507);
xor U4104 (N_4104,N_877,N_1813);
or U4105 (N_4105,N_376,N_2024);
or U4106 (N_4106,N_1586,N_1447);
nand U4107 (N_4107,N_3098,N_2707);
nand U4108 (N_4108,N_1912,N_2199);
nor U4109 (N_4109,N_270,N_323);
or U4110 (N_4110,N_2646,N_967);
xor U4111 (N_4111,N_2469,N_2501);
xnor U4112 (N_4112,N_3025,N_2095);
xnor U4113 (N_4113,N_175,N_2073);
or U4114 (N_4114,N_1798,N_827);
nor U4115 (N_4115,N_372,N_779);
and U4116 (N_4116,N_498,N_798);
or U4117 (N_4117,N_2225,N_724);
and U4118 (N_4118,N_1543,N_1576);
nand U4119 (N_4119,N_136,N_2726);
or U4120 (N_4120,N_3112,N_2424);
and U4121 (N_4121,N_2245,N_1302);
xor U4122 (N_4122,N_941,N_892);
xor U4123 (N_4123,N_2240,N_1049);
nor U4124 (N_4124,N_1523,N_2935);
nand U4125 (N_4125,N_1375,N_660);
and U4126 (N_4126,N_1976,N_1532);
and U4127 (N_4127,N_2175,N_241);
or U4128 (N_4128,N_1169,N_2239);
and U4129 (N_4129,N_2213,N_2211);
xnor U4130 (N_4130,N_2269,N_1556);
and U4131 (N_4131,N_1449,N_1298);
nor U4132 (N_4132,N_1341,N_295);
nor U4133 (N_4133,N_1807,N_1584);
nand U4134 (N_4134,N_2014,N_312);
nor U4135 (N_4135,N_611,N_1340);
and U4136 (N_4136,N_2796,N_2471);
nand U4137 (N_4137,N_1524,N_3027);
and U4138 (N_4138,N_2795,N_916);
or U4139 (N_4139,N_2146,N_2350);
nor U4140 (N_4140,N_1955,N_876);
and U4141 (N_4141,N_2672,N_1517);
and U4142 (N_4142,N_1381,N_1077);
or U4143 (N_4143,N_989,N_1548);
or U4144 (N_4144,N_2280,N_447);
or U4145 (N_4145,N_1240,N_1486);
or U4146 (N_4146,N_385,N_1646);
nor U4147 (N_4147,N_1496,N_2232);
nor U4148 (N_4148,N_765,N_772);
xor U4149 (N_4149,N_1977,N_245);
nor U4150 (N_4150,N_2001,N_343);
nand U4151 (N_4151,N_458,N_1314);
xor U4152 (N_4152,N_2800,N_2961);
or U4153 (N_4153,N_1348,N_1544);
nand U4154 (N_4154,N_2662,N_2983);
nand U4155 (N_4155,N_378,N_3077);
nor U4156 (N_4156,N_1699,N_3019);
or U4157 (N_4157,N_1229,N_200);
nor U4158 (N_4158,N_595,N_1619);
xor U4159 (N_4159,N_1941,N_353);
or U4160 (N_4160,N_1446,N_3114);
xor U4161 (N_4161,N_484,N_2129);
nor U4162 (N_4162,N_73,N_2035);
or U4163 (N_4163,N_782,N_1177);
xnor U4164 (N_4164,N_211,N_542);
and U4165 (N_4165,N_715,N_555);
nor U4166 (N_4166,N_2724,N_557);
xnor U4167 (N_4167,N_2787,N_1357);
nor U4168 (N_4168,N_1451,N_2198);
and U4169 (N_4169,N_2988,N_1463);
nor U4170 (N_4170,N_1453,N_1970);
or U4171 (N_4171,N_2267,N_440);
or U4172 (N_4172,N_2630,N_1301);
and U4173 (N_4173,N_906,N_2556);
xor U4174 (N_4174,N_1659,N_2784);
or U4175 (N_4175,N_683,N_418);
xnor U4176 (N_4176,N_500,N_2489);
nand U4177 (N_4177,N_2747,N_2530);
or U4178 (N_4178,N_826,N_1895);
or U4179 (N_4179,N_3105,N_3048);
or U4180 (N_4180,N_2845,N_1883);
and U4181 (N_4181,N_1056,N_1826);
xnor U4182 (N_4182,N_1824,N_1531);
nor U4183 (N_4183,N_2022,N_2792);
xnor U4184 (N_4184,N_856,N_2328);
nor U4185 (N_4185,N_2880,N_1539);
nor U4186 (N_4186,N_224,N_179);
xor U4187 (N_4187,N_460,N_2802);
nor U4188 (N_4188,N_631,N_675);
nand U4189 (N_4189,N_736,N_3122);
and U4190 (N_4190,N_389,N_1474);
and U4191 (N_4191,N_3066,N_1547);
or U4192 (N_4192,N_2514,N_330);
and U4193 (N_4193,N_1021,N_1959);
xnor U4194 (N_4194,N_917,N_1071);
nor U4195 (N_4195,N_1757,N_1470);
xnor U4196 (N_4196,N_3000,N_1724);
or U4197 (N_4197,N_1297,N_801);
nor U4198 (N_4198,N_2529,N_2500);
nand U4199 (N_4199,N_1678,N_2970);
or U4200 (N_4200,N_3068,N_2480);
xnor U4201 (N_4201,N_1076,N_1922);
and U4202 (N_4202,N_1567,N_1405);
xnor U4203 (N_4203,N_184,N_1673);
or U4204 (N_4204,N_70,N_273);
nor U4205 (N_4205,N_1080,N_2032);
nand U4206 (N_4206,N_2356,N_618);
nand U4207 (N_4207,N_1172,N_1491);
and U4208 (N_4208,N_1094,N_600);
nand U4209 (N_4209,N_775,N_769);
and U4210 (N_4210,N_2018,N_3063);
nor U4211 (N_4211,N_55,N_81);
nand U4212 (N_4212,N_2196,N_2047);
nand U4213 (N_4213,N_1613,N_888);
and U4214 (N_4214,N_1624,N_2078);
and U4215 (N_4215,N_2782,N_1259);
xnor U4216 (N_4216,N_1300,N_1746);
or U4217 (N_4217,N_1792,N_3034);
nand U4218 (N_4218,N_2685,N_468);
and U4219 (N_4219,N_2191,N_1842);
or U4220 (N_4220,N_192,N_1863);
nand U4221 (N_4221,N_1204,N_1228);
xor U4222 (N_4222,N_1508,N_2340);
and U4223 (N_4223,N_2506,N_934);
nor U4224 (N_4224,N_883,N_2057);
xor U4225 (N_4225,N_321,N_1221);
nand U4226 (N_4226,N_2054,N_878);
nor U4227 (N_4227,N_237,N_17);
nand U4228 (N_4228,N_119,N_680);
or U4229 (N_4229,N_1660,N_1466);
xnor U4230 (N_4230,N_20,N_1087);
or U4231 (N_4231,N_324,N_2809);
xnor U4232 (N_4232,N_2405,N_1193);
xnor U4233 (N_4233,N_212,N_514);
nand U4234 (N_4234,N_530,N_2582);
nor U4235 (N_4235,N_665,N_632);
or U4236 (N_4236,N_2038,N_67);
nor U4237 (N_4237,N_2456,N_3017);
nor U4238 (N_4238,N_1888,N_954);
nor U4239 (N_4239,N_2870,N_2972);
nand U4240 (N_4240,N_2201,N_1407);
or U4241 (N_4241,N_924,N_1189);
nand U4242 (N_4242,N_867,N_2040);
nor U4243 (N_4243,N_1855,N_2492);
or U4244 (N_4244,N_1638,N_1024);
nand U4245 (N_4245,N_2262,N_767);
nand U4246 (N_4246,N_1211,N_2673);
and U4247 (N_4247,N_2142,N_2450);
nand U4248 (N_4248,N_2464,N_656);
and U4249 (N_4249,N_1465,N_1171);
xnor U4250 (N_4250,N_1128,N_3074);
nand U4251 (N_4251,N_759,N_371);
and U4252 (N_4252,N_1371,N_2775);
nor U4253 (N_4253,N_2759,N_2493);
nor U4254 (N_4254,N_1674,N_2780);
xnor U4255 (N_4255,N_3110,N_532);
or U4256 (N_4256,N_2565,N_676);
and U4257 (N_4257,N_465,N_565);
and U4258 (N_4258,N_679,N_2345);
or U4259 (N_4259,N_2915,N_1847);
or U4260 (N_4260,N_3006,N_521);
nor U4261 (N_4261,N_146,N_2344);
nand U4262 (N_4262,N_2193,N_1870);
nand U4263 (N_4263,N_2655,N_1513);
nor U4264 (N_4264,N_448,N_1217);
or U4265 (N_4265,N_1233,N_1937);
xnor U4266 (N_4266,N_1267,N_2049);
xnor U4267 (N_4267,N_2124,N_879);
or U4268 (N_4268,N_2226,N_286);
or U4269 (N_4269,N_838,N_2768);
nor U4270 (N_4270,N_551,N_2921);
nor U4271 (N_4271,N_2292,N_2105);
or U4272 (N_4272,N_787,N_2910);
nor U4273 (N_4273,N_282,N_85);
xnor U4274 (N_4274,N_2538,N_1051);
or U4275 (N_4275,N_2916,N_1262);
xnor U4276 (N_4276,N_1651,N_409);
and U4277 (N_4277,N_606,N_957);
nand U4278 (N_4278,N_1622,N_1868);
xnor U4279 (N_4279,N_111,N_2838);
nor U4280 (N_4280,N_304,N_169);
xor U4281 (N_4281,N_2354,N_1512);
nand U4282 (N_4282,N_79,N_2268);
or U4283 (N_4283,N_3101,N_328);
or U4284 (N_4284,N_619,N_2260);
and U4285 (N_4285,N_860,N_96);
nand U4286 (N_4286,N_135,N_3030);
and U4287 (N_4287,N_729,N_302);
nor U4288 (N_4288,N_1521,N_1092);
or U4289 (N_4289,N_1419,N_1044);
nor U4290 (N_4290,N_2336,N_2386);
or U4291 (N_4291,N_674,N_272);
or U4292 (N_4292,N_961,N_128);
and U4293 (N_4293,N_1464,N_897);
nor U4294 (N_4294,N_1784,N_935);
or U4295 (N_4295,N_1986,N_2572);
nand U4296 (N_4296,N_873,N_1440);
xnor U4297 (N_4297,N_1020,N_1336);
and U4298 (N_4298,N_1455,N_2811);
or U4299 (N_4299,N_884,N_393);
and U4300 (N_4300,N_915,N_1643);
and U4301 (N_4301,N_28,N_1144);
or U4302 (N_4302,N_285,N_2728);
nand U4303 (N_4303,N_2410,N_91);
and U4304 (N_4304,N_501,N_149);
xnor U4305 (N_4305,N_2640,N_1084);
nor U4306 (N_4306,N_408,N_2306);
nor U4307 (N_4307,N_29,N_3106);
xnor U4308 (N_4308,N_2234,N_1769);
nand U4309 (N_4309,N_834,N_1468);
and U4310 (N_4310,N_3121,N_2755);
xor U4311 (N_4311,N_2965,N_2894);
and U4312 (N_4312,N_1373,N_588);
and U4313 (N_4313,N_2769,N_1353);
or U4314 (N_4314,N_1867,N_3055);
xor U4315 (N_4315,N_1157,N_1615);
xnor U4316 (N_4316,N_247,N_905);
or U4317 (N_4317,N_1996,N_1647);
xnor U4318 (N_4318,N_1664,N_2100);
and U4319 (N_4319,N_102,N_2319);
nor U4320 (N_4320,N_854,N_2458);
or U4321 (N_4321,N_2713,N_454);
or U4322 (N_4322,N_1394,N_57);
or U4323 (N_4323,N_1178,N_277);
nand U4324 (N_4324,N_362,N_2178);
or U4325 (N_4325,N_431,N_852);
nor U4326 (N_4326,N_1975,N_1383);
nand U4327 (N_4327,N_1392,N_1372);
or U4328 (N_4328,N_1790,N_2741);
and U4329 (N_4329,N_2622,N_1817);
and U4330 (N_4330,N_1742,N_2743);
nand U4331 (N_4331,N_1432,N_2281);
nor U4332 (N_4332,N_218,N_2367);
nand U4333 (N_4333,N_1323,N_1093);
or U4334 (N_4334,N_1265,N_1989);
xor U4335 (N_4335,N_1264,N_2647);
or U4336 (N_4336,N_1482,N_141);
or U4337 (N_4337,N_462,N_1206);
nor U4338 (N_4338,N_2457,N_1714);
nor U4339 (N_4339,N_1964,N_3100);
nor U4340 (N_4340,N_1343,N_1038);
nor U4341 (N_4341,N_2901,N_1363);
xnor U4342 (N_4342,N_106,N_1404);
and U4343 (N_4343,N_148,N_2624);
xor U4344 (N_4344,N_2861,N_1655);
or U4345 (N_4345,N_2277,N_1858);
nor U4346 (N_4346,N_1188,N_932);
xor U4347 (N_4347,N_2371,N_666);
and U4348 (N_4348,N_2863,N_2019);
and U4349 (N_4349,N_383,N_2757);
and U4350 (N_4350,N_1263,N_2605);
nor U4351 (N_4351,N_495,N_2027);
or U4352 (N_4352,N_416,N_858);
and U4353 (N_4353,N_2123,N_1219);
nor U4354 (N_4354,N_187,N_1276);
xnor U4355 (N_4355,N_1081,N_2964);
and U4356 (N_4356,N_1672,N_513);
nand U4357 (N_4357,N_2805,N_1456);
nor U4358 (N_4358,N_938,N_278);
nor U4359 (N_4359,N_2033,N_1942);
and U4360 (N_4360,N_1207,N_367);
nand U4361 (N_4361,N_1645,N_2217);
and U4362 (N_4362,N_1693,N_1180);
nand U4363 (N_4363,N_1866,N_1617);
nand U4364 (N_4364,N_969,N_1283);
nor U4365 (N_4365,N_1006,N_1697);
and U4366 (N_4366,N_741,N_2339);
xnor U4367 (N_4367,N_1173,N_411);
nand U4368 (N_4368,N_997,N_252);
and U4369 (N_4369,N_1720,N_2648);
nor U4370 (N_4370,N_2168,N_561);
xor U4371 (N_4371,N_1929,N_2166);
xnor U4372 (N_4372,N_2505,N_2481);
nand U4373 (N_4373,N_1430,N_2176);
nand U4374 (N_4374,N_1186,N_2098);
and U4375 (N_4375,N_1936,N_2391);
nor U4376 (N_4376,N_2822,N_226);
xnor U4377 (N_4377,N_1498,N_436);
nand U4378 (N_4378,N_2,N_3024);
and U4379 (N_4379,N_976,N_307);
nor U4380 (N_4380,N_1352,N_2121);
and U4381 (N_4381,N_1809,N_2216);
or U4382 (N_4382,N_1926,N_1808);
xor U4383 (N_4383,N_1838,N_914);
nand U4384 (N_4384,N_2978,N_1707);
xnor U4385 (N_4385,N_2872,N_403);
or U4386 (N_4386,N_1061,N_1526);
nand U4387 (N_4387,N_322,N_439);
and U4388 (N_4388,N_1495,N_686);
and U4389 (N_4389,N_2119,N_1852);
xor U4390 (N_4390,N_1931,N_1110);
nor U4391 (N_4391,N_2495,N_14);
nand U4392 (N_4392,N_1818,N_824);
xnor U4393 (N_4393,N_2462,N_795);
nand U4394 (N_4394,N_1135,N_2491);
or U4395 (N_4395,N_1488,N_31);
nand U4396 (N_4396,N_2043,N_2594);
or U4397 (N_4397,N_1787,N_855);
xor U4398 (N_4398,N_677,N_1803);
or U4399 (N_4399,N_2287,N_1378);
xnor U4400 (N_4400,N_2680,N_2926);
nor U4401 (N_4401,N_2502,N_1654);
or U4402 (N_4402,N_918,N_2541);
xor U4403 (N_4403,N_625,N_139);
nand U4404 (N_4404,N_2657,N_471);
nand U4405 (N_4405,N_24,N_1840);
or U4406 (N_4406,N_1332,N_547);
nor U4407 (N_4407,N_604,N_1401);
or U4408 (N_4408,N_972,N_747);
or U4409 (N_4409,N_1529,N_2065);
or U4410 (N_4410,N_1198,N_577);
xnor U4411 (N_4411,N_3033,N_2900);
and U4412 (N_4412,N_2248,N_2816);
or U4413 (N_4413,N_99,N_2039);
xnor U4414 (N_4414,N_942,N_1961);
or U4415 (N_4415,N_2147,N_176);
and U4416 (N_4416,N_2411,N_1220);
and U4417 (N_4417,N_2579,N_1235);
and U4418 (N_4418,N_2626,N_1388);
and U4419 (N_4419,N_1421,N_2865);
nand U4420 (N_4420,N_608,N_1184);
nor U4421 (N_4421,N_1131,N_2126);
and U4422 (N_4422,N_1212,N_1569);
xnor U4423 (N_4423,N_93,N_108);
nor U4424 (N_4424,N_1571,N_872);
xnor U4425 (N_4425,N_90,N_1295);
and U4426 (N_4426,N_853,N_2055);
xnor U4427 (N_4427,N_443,N_3042);
xor U4428 (N_4428,N_2950,N_56);
xnor U4429 (N_4429,N_744,N_1112);
or U4430 (N_4430,N_1777,N_153);
xor U4431 (N_4431,N_642,N_1881);
nor U4432 (N_4432,N_401,N_2528);
nor U4433 (N_4433,N_2187,N_1740);
and U4434 (N_4434,N_2609,N_2569);
nand U4435 (N_4435,N_2676,N_1050);
nor U4436 (N_4436,N_1775,N_2581);
and U4437 (N_4437,N_2343,N_2878);
nor U4438 (N_4438,N_1035,N_1642);
nand U4439 (N_4439,N_1873,N_1594);
or U4440 (N_4440,N_3022,N_2051);
and U4441 (N_4441,N_1379,N_1090);
and U4442 (N_4442,N_2652,N_687);
and U4443 (N_4443,N_1230,N_260);
xor U4444 (N_4444,N_2984,N_2285);
nor U4445 (N_4445,N_1944,N_2242);
nor U4446 (N_4446,N_615,N_538);
or U4447 (N_4447,N_1269,N_1609);
or U4448 (N_4448,N_2913,N_541);
and U4449 (N_4449,N_885,N_2727);
or U4450 (N_4450,N_435,N_1550);
nand U4451 (N_4451,N_2173,N_2534);
xor U4452 (N_4452,N_3035,N_75);
nand U4453 (N_4453,N_1631,N_348);
or U4454 (N_4454,N_1079,N_144);
nor U4455 (N_4455,N_2922,N_1208);
and U4456 (N_4456,N_1585,N_2642);
xor U4457 (N_4457,N_886,N_519);
and U4458 (N_4458,N_2831,N_1885);
and U4459 (N_4459,N_1387,N_1073);
nand U4460 (N_4460,N_269,N_446);
and U4461 (N_4461,N_593,N_1834);
nand U4462 (N_4462,N_982,N_993);
xor U4463 (N_4463,N_738,N_3059);
nand U4464 (N_4464,N_382,N_2762);
xnor U4465 (N_4465,N_2907,N_77);
or U4466 (N_4466,N_238,N_2159);
or U4467 (N_4467,N_2007,N_344);
xor U4468 (N_4468,N_571,N_3043);
xnor U4469 (N_4469,N_2003,N_413);
xor U4470 (N_4470,N_2531,N_1723);
and U4471 (N_4471,N_2499,N_1028);
and U4472 (N_4472,N_2518,N_1806);
nor U4473 (N_4473,N_2817,N_2241);
nor U4474 (N_4474,N_2108,N_1753);
and U4475 (N_4475,N_2310,N_643);
and U4476 (N_4476,N_325,N_1384);
xor U4477 (N_4477,N_2674,N_2061);
and U4478 (N_4478,N_1238,N_2296);
nand U4479 (N_4479,N_65,N_1920);
or U4480 (N_4480,N_2376,N_899);
xor U4481 (N_4481,N_2821,N_1335);
nor U4482 (N_4482,N_159,N_1369);
or U4483 (N_4483,N_2875,N_2251);
and U4484 (N_4484,N_673,N_1304);
or U4485 (N_4485,N_1696,N_2508);
or U4486 (N_4486,N_791,N_1338);
and U4487 (N_4487,N_145,N_2548);
and U4488 (N_4488,N_1256,N_1410);
and U4489 (N_4489,N_11,N_417);
or U4490 (N_4490,N_1396,N_2026);
or U4491 (N_4491,N_512,N_573);
nor U4492 (N_4492,N_894,N_427);
or U4493 (N_4493,N_428,N_2692);
nand U4494 (N_4494,N_381,N_1367);
or U4495 (N_4495,N_2832,N_790);
nor U4496 (N_4496,N_2923,N_2353);
xor U4497 (N_4497,N_2765,N_2041);
nand U4498 (N_4498,N_651,N_711);
nor U4499 (N_4499,N_531,N_2602);
xor U4500 (N_4500,N_1587,N_1574);
and U4501 (N_4501,N_124,N_1239);
nand U4502 (N_4502,N_239,N_98);
and U4503 (N_4503,N_1266,N_213);
xor U4504 (N_4504,N_2330,N_2020);
and U4505 (N_4505,N_2427,N_442);
xnor U4506 (N_4506,N_2214,N_2482);
or U4507 (N_4507,N_2793,N_2829);
nand U4508 (N_4508,N_859,N_576);
or U4509 (N_4509,N_2164,N_2259);
or U4510 (N_4510,N_2094,N_1770);
or U4511 (N_4511,N_1590,N_3012);
or U4512 (N_4512,N_2256,N_1914);
nor U4513 (N_4513,N_1414,N_2404);
xnor U4514 (N_4514,N_243,N_2485);
and U4515 (N_4515,N_1036,N_2879);
and U4516 (N_4516,N_773,N_195);
and U4517 (N_4517,N_804,N_921);
nand U4518 (N_4518,N_1499,N_2993);
nand U4519 (N_4519,N_955,N_2885);
nand U4520 (N_4520,N_1700,N_1068);
and U4521 (N_4521,N_745,N_2434);
and U4522 (N_4522,N_1766,N_1047);
nand U4523 (N_4523,N_2002,N_445);
and U4524 (N_4524,N_41,N_3044);
or U4525 (N_4525,N_1987,N_338);
or U4526 (N_4526,N_1248,N_1122);
nor U4527 (N_4527,N_627,N_1990);
and U4528 (N_4528,N_78,N_3108);
xor U4529 (N_4529,N_419,N_2297);
or U4530 (N_4530,N_492,N_183);
or U4531 (N_4531,N_2945,N_160);
nand U4532 (N_4532,N_2698,N_1704);
nand U4533 (N_4533,N_2520,N_1612);
or U4534 (N_4534,N_1538,N_1969);
nor U4535 (N_4535,N_1096,N_740);
xor U4536 (N_4536,N_880,N_1201);
or U4537 (N_4537,N_1572,N_1691);
xor U4538 (N_4538,N_2348,N_2109);
and U4539 (N_4539,N_2110,N_985);
and U4540 (N_4540,N_2839,N_1278);
nor U4541 (N_4541,N_1492,N_2062);
nand U4542 (N_4542,N_3047,N_1033);
xor U4543 (N_4543,N_288,N_661);
xnor U4544 (N_4544,N_1894,N_1066);
nor U4545 (N_4545,N_109,N_133);
or U4546 (N_4546,N_467,N_1475);
and U4547 (N_4547,N_156,N_919);
nor U4548 (N_4548,N_3007,N_2357);
xnor U4549 (N_4549,N_1943,N_1965);
and U4550 (N_4550,N_1143,N_669);
nand U4551 (N_4551,N_2563,N_3115);
or U4552 (N_4552,N_105,N_1502);
xor U4553 (N_4553,N_2352,N_2516);
or U4554 (N_4554,N_2803,N_2221);
nor U4555 (N_4555,N_1318,N_2553);
nand U4556 (N_4556,N_230,N_2419);
nand U4557 (N_4557,N_2203,N_104);
or U4558 (N_4558,N_1243,N_305);
and U4559 (N_4559,N_297,N_1898);
nor U4560 (N_4560,N_2184,N_470);
nor U4561 (N_4561,N_1411,N_266);
or U4562 (N_4562,N_1994,N_80);
nand U4563 (N_4563,N_2360,N_696);
nor U4564 (N_4564,N_840,N_87);
nor U4565 (N_4565,N_1479,N_2385);
nand U4566 (N_4566,N_92,N_812);
and U4567 (N_4567,N_1127,N_890);
or U4568 (N_4568,N_1516,N_2620);
nor U4569 (N_4569,N_3029,N_2475);
or U4570 (N_4570,N_830,N_1795);
nand U4571 (N_4571,N_1669,N_2048);
and U4572 (N_4572,N_1125,N_1000);
nand U4573 (N_4573,N_1119,N_1398);
nand U4574 (N_4574,N_2423,N_2311);
xnor U4575 (N_4575,N_731,N_491);
nor U4576 (N_4576,N_1308,N_1756);
nand U4577 (N_4577,N_52,N_2975);
and U4578 (N_4578,N_1635,N_1284);
nor U4579 (N_4579,N_960,N_579);
nand U4580 (N_4580,N_2365,N_1522);
or U4581 (N_4581,N_2415,N_6);
nor U4582 (N_4582,N_198,N_3010);
nand U4583 (N_4583,N_2171,N_130);
and U4584 (N_4584,N_61,N_1039);
xnor U4585 (N_4585,N_2452,N_2607);
xnor U4586 (N_4586,N_203,N_469);
nand U4587 (N_4587,N_1579,N_2933);
or U4588 (N_4588,N_249,N_2824);
nor U4589 (N_4589,N_1703,N_172);
nor U4590 (N_4590,N_2959,N_2069);
xnor U4591 (N_4591,N_1142,N_1559);
and U4592 (N_4592,N_424,N_2414);
nand U4593 (N_4593,N_2957,N_1666);
and U4594 (N_4594,N_1811,N_2192);
xnor U4595 (N_4595,N_2552,N_1933);
xor U4596 (N_4596,N_2751,N_2627);
nand U4597 (N_4597,N_605,N_1060);
and U4598 (N_4598,N_659,N_992);
nand U4599 (N_4599,N_8,N_722);
nor U4600 (N_4600,N_402,N_1034);
nor U4601 (N_4601,N_474,N_2284);
nor U4602 (N_4602,N_1930,N_1841);
or U4603 (N_4603,N_1815,N_1640);
nor U4604 (N_4604,N_165,N_3032);
nand U4605 (N_4605,N_2846,N_2059);
nand U4606 (N_4606,N_875,N_900);
nand U4607 (N_4607,N_2079,N_255);
nand U4608 (N_4608,N_1689,N_2536);
or U4609 (N_4609,N_2179,N_2084);
xor U4610 (N_4610,N_1573,N_1472);
or U4611 (N_4611,N_1940,N_733);
nand U4612 (N_4612,N_2703,N_171);
and U4613 (N_4613,N_486,N_506);
nand U4614 (N_4614,N_1251,N_2230);
xor U4615 (N_4615,N_3107,N_1900);
or U4616 (N_4616,N_1003,N_267);
and U4617 (N_4617,N_1159,N_1541);
nand U4618 (N_4618,N_1031,N_603);
xnor U4619 (N_4619,N_3117,N_1802);
and U4620 (N_4620,N_2206,N_308);
nor U4621 (N_4621,N_2204,N_726);
xnor U4622 (N_4622,N_1962,N_1552);
or U4623 (N_4623,N_1197,N_3103);
nand U4624 (N_4624,N_620,N_681);
nand U4625 (N_4625,N_355,N_2425);
nand U4626 (N_4626,N_1158,N_1751);
or U4627 (N_4627,N_1059,N_505);
nor U4628 (N_4628,N_807,N_2695);
or U4629 (N_4629,N_2131,N_1277);
and U4630 (N_4630,N_303,N_2407);
nand U4631 (N_4631,N_2066,N_2644);
xnor U4632 (N_4632,N_1026,N_0);
and U4633 (N_4633,N_365,N_2679);
xnor U4634 (N_4634,N_2058,N_549);
nor U4635 (N_4635,N_2440,N_2930);
xnor U4636 (N_4636,N_2892,N_987);
nand U4637 (N_4637,N_1801,N_2477);
xnor U4638 (N_4638,N_2291,N_1058);
nand U4639 (N_4639,N_3001,N_225);
xor U4640 (N_4640,N_811,N_1433);
nand U4641 (N_4641,N_1536,N_207);
nor U4642 (N_4642,N_2517,N_1862);
and U4643 (N_4643,N_1485,N_2653);
or U4644 (N_4644,N_313,N_1710);
nand U4645 (N_4645,N_2871,N_1626);
or U4646 (N_4646,N_2342,N_2403);
and U4647 (N_4647,N_2639,N_1705);
nand U4648 (N_4648,N_1347,N_517);
nand U4649 (N_4649,N_1565,N_889);
xnor U4650 (N_4650,N_246,N_968);
nand U4651 (N_4651,N_1362,N_2716);
nand U4652 (N_4652,N_2294,N_2746);
or U4653 (N_4653,N_2158,N_2361);
nand U4654 (N_4654,N_936,N_2382);
xnor U4655 (N_4655,N_229,N_628);
or U4656 (N_4656,N_475,N_316);
xnor U4657 (N_4657,N_536,N_2721);
nor U4658 (N_4658,N_507,N_1062);
nand U4659 (N_4659,N_2238,N_2278);
xor U4660 (N_4660,N_1413,N_2857);
nor U4661 (N_4661,N_1360,N_1985);
or U4662 (N_4662,N_2025,N_2521);
nor U4663 (N_4663,N_167,N_2042);
xor U4664 (N_4664,N_1458,N_1374);
nand U4665 (N_4665,N_1103,N_567);
and U4666 (N_4666,N_1130,N_72);
nor U4667 (N_4667,N_2715,N_2461);
and U4668 (N_4668,N_464,N_898);
or U4669 (N_4669,N_1260,N_846);
nor U4670 (N_4670,N_482,N_709);
or U4671 (N_4671,N_3073,N_349);
xor U4672 (N_4672,N_1313,N_1133);
nand U4673 (N_4673,N_2139,N_706);
and U4674 (N_4674,N_2151,N_201);
xor U4675 (N_4675,N_1910,N_1773);
xnor U4676 (N_4676,N_751,N_2133);
and U4677 (N_4677,N_558,N_2544);
nand U4678 (N_4678,N_2778,N_235);
nand U4679 (N_4679,N_1227,N_331);
or U4680 (N_4680,N_1356,N_1925);
or U4681 (N_4681,N_654,N_103);
and U4682 (N_4682,N_590,N_123);
and U4683 (N_4683,N_3040,N_234);
nand U4684 (N_4684,N_189,N_2638);
nand U4685 (N_4685,N_1665,N_1181);
nor U4686 (N_4686,N_387,N_395);
xor U4687 (N_4687,N_1291,N_1258);
and U4688 (N_4688,N_3076,N_2150);
or U4689 (N_4689,N_93,N_707);
xor U4690 (N_4690,N_2478,N_2502);
or U4691 (N_4691,N_1693,N_2228);
nor U4692 (N_4692,N_3021,N_710);
nor U4693 (N_4693,N_1832,N_2400);
or U4694 (N_4694,N_560,N_387);
nand U4695 (N_4695,N_87,N_2257);
or U4696 (N_4696,N_989,N_1015);
xor U4697 (N_4697,N_250,N_873);
and U4698 (N_4698,N_1498,N_61);
and U4699 (N_4699,N_1248,N_1881);
nor U4700 (N_4700,N_2319,N_2431);
and U4701 (N_4701,N_2723,N_884);
and U4702 (N_4702,N_3083,N_1818);
xor U4703 (N_4703,N_1107,N_2185);
xnor U4704 (N_4704,N_2149,N_1981);
nor U4705 (N_4705,N_2385,N_2375);
nor U4706 (N_4706,N_811,N_580);
or U4707 (N_4707,N_1546,N_564);
nor U4708 (N_4708,N_191,N_2417);
and U4709 (N_4709,N_1157,N_508);
and U4710 (N_4710,N_415,N_140);
nor U4711 (N_4711,N_426,N_257);
and U4712 (N_4712,N_953,N_2554);
nand U4713 (N_4713,N_1970,N_2997);
and U4714 (N_4714,N_311,N_1786);
xnor U4715 (N_4715,N_1618,N_696);
and U4716 (N_4716,N_698,N_2089);
xor U4717 (N_4717,N_1096,N_2438);
nand U4718 (N_4718,N_1058,N_820);
xor U4719 (N_4719,N_365,N_1240);
and U4720 (N_4720,N_2254,N_2911);
or U4721 (N_4721,N_236,N_2652);
or U4722 (N_4722,N_430,N_1323);
nand U4723 (N_4723,N_2403,N_2449);
or U4724 (N_4724,N_1910,N_933);
and U4725 (N_4725,N_2274,N_330);
xnor U4726 (N_4726,N_3089,N_2372);
and U4727 (N_4727,N_1413,N_940);
nand U4728 (N_4728,N_2704,N_427);
and U4729 (N_4729,N_675,N_3033);
or U4730 (N_4730,N_2373,N_245);
nor U4731 (N_4731,N_2012,N_510);
and U4732 (N_4732,N_94,N_1651);
nor U4733 (N_4733,N_2381,N_15);
xnor U4734 (N_4734,N_2359,N_295);
nand U4735 (N_4735,N_2745,N_151);
nand U4736 (N_4736,N_2020,N_802);
or U4737 (N_4737,N_1869,N_918);
or U4738 (N_4738,N_2370,N_437);
nor U4739 (N_4739,N_2904,N_979);
and U4740 (N_4740,N_620,N_600);
xor U4741 (N_4741,N_2171,N_2503);
or U4742 (N_4742,N_3024,N_584);
or U4743 (N_4743,N_2634,N_2314);
xor U4744 (N_4744,N_2518,N_2555);
and U4745 (N_4745,N_2404,N_976);
nand U4746 (N_4746,N_1289,N_2398);
nor U4747 (N_4747,N_1013,N_1485);
nor U4748 (N_4748,N_90,N_2776);
or U4749 (N_4749,N_432,N_2626);
or U4750 (N_4750,N_1906,N_686);
nand U4751 (N_4751,N_2577,N_792);
xnor U4752 (N_4752,N_1591,N_1845);
nand U4753 (N_4753,N_2404,N_2017);
xor U4754 (N_4754,N_2251,N_964);
and U4755 (N_4755,N_416,N_2733);
nand U4756 (N_4756,N_34,N_2889);
and U4757 (N_4757,N_2998,N_573);
or U4758 (N_4758,N_2414,N_609);
nand U4759 (N_4759,N_3103,N_667);
xnor U4760 (N_4760,N_1972,N_2743);
nand U4761 (N_4761,N_620,N_411);
nand U4762 (N_4762,N_1431,N_209);
nor U4763 (N_4763,N_1590,N_1549);
or U4764 (N_4764,N_287,N_1762);
xor U4765 (N_4765,N_785,N_1291);
nand U4766 (N_4766,N_2672,N_2248);
and U4767 (N_4767,N_2937,N_2592);
xor U4768 (N_4768,N_2839,N_1909);
nor U4769 (N_4769,N_2608,N_2535);
xor U4770 (N_4770,N_685,N_1886);
xor U4771 (N_4771,N_2396,N_865);
or U4772 (N_4772,N_1276,N_1241);
nor U4773 (N_4773,N_2638,N_755);
nor U4774 (N_4774,N_398,N_1149);
or U4775 (N_4775,N_375,N_1673);
xnor U4776 (N_4776,N_1869,N_2961);
and U4777 (N_4777,N_395,N_2614);
xnor U4778 (N_4778,N_2606,N_2926);
or U4779 (N_4779,N_2364,N_934);
and U4780 (N_4780,N_1475,N_1269);
xor U4781 (N_4781,N_1826,N_236);
xor U4782 (N_4782,N_1090,N_1687);
nand U4783 (N_4783,N_3088,N_2353);
or U4784 (N_4784,N_593,N_2440);
xor U4785 (N_4785,N_1347,N_1223);
or U4786 (N_4786,N_786,N_660);
and U4787 (N_4787,N_1108,N_221);
xor U4788 (N_4788,N_1226,N_1515);
xnor U4789 (N_4789,N_755,N_2024);
or U4790 (N_4790,N_296,N_2539);
and U4791 (N_4791,N_1535,N_2817);
and U4792 (N_4792,N_3045,N_1189);
xnor U4793 (N_4793,N_822,N_2823);
nor U4794 (N_4794,N_2091,N_2932);
or U4795 (N_4795,N_628,N_2712);
nor U4796 (N_4796,N_432,N_3043);
nand U4797 (N_4797,N_1553,N_911);
xor U4798 (N_4798,N_2479,N_2878);
xor U4799 (N_4799,N_337,N_601);
xnor U4800 (N_4800,N_2198,N_2139);
nand U4801 (N_4801,N_1680,N_520);
nor U4802 (N_4802,N_2775,N_1344);
or U4803 (N_4803,N_1716,N_2857);
and U4804 (N_4804,N_608,N_94);
or U4805 (N_4805,N_629,N_1161);
nand U4806 (N_4806,N_452,N_259);
nor U4807 (N_4807,N_440,N_2435);
nor U4808 (N_4808,N_2487,N_1712);
and U4809 (N_4809,N_361,N_953);
xor U4810 (N_4810,N_1599,N_3049);
or U4811 (N_4811,N_684,N_1003);
or U4812 (N_4812,N_2881,N_771);
and U4813 (N_4813,N_3016,N_2161);
nand U4814 (N_4814,N_802,N_1172);
and U4815 (N_4815,N_2401,N_2276);
nand U4816 (N_4816,N_1086,N_940);
and U4817 (N_4817,N_1952,N_1911);
and U4818 (N_4818,N_1930,N_2041);
or U4819 (N_4819,N_928,N_2318);
nor U4820 (N_4820,N_338,N_3032);
nor U4821 (N_4821,N_633,N_933);
nand U4822 (N_4822,N_143,N_1551);
and U4823 (N_4823,N_1355,N_1811);
nand U4824 (N_4824,N_1094,N_948);
or U4825 (N_4825,N_79,N_2955);
nand U4826 (N_4826,N_2185,N_822);
nor U4827 (N_4827,N_2376,N_1639);
xnor U4828 (N_4828,N_228,N_602);
nor U4829 (N_4829,N_2524,N_2642);
and U4830 (N_4830,N_370,N_2942);
nor U4831 (N_4831,N_355,N_2095);
nor U4832 (N_4832,N_2755,N_773);
and U4833 (N_4833,N_680,N_1174);
nor U4834 (N_4834,N_1216,N_1197);
and U4835 (N_4835,N_1082,N_1103);
nand U4836 (N_4836,N_2993,N_996);
or U4837 (N_4837,N_2540,N_709);
nor U4838 (N_4838,N_1436,N_153);
or U4839 (N_4839,N_701,N_2630);
nand U4840 (N_4840,N_2541,N_1421);
nor U4841 (N_4841,N_2278,N_2590);
xnor U4842 (N_4842,N_1803,N_70);
nand U4843 (N_4843,N_200,N_2543);
and U4844 (N_4844,N_959,N_1682);
nor U4845 (N_4845,N_731,N_1453);
and U4846 (N_4846,N_1483,N_69);
and U4847 (N_4847,N_1101,N_1225);
or U4848 (N_4848,N_1521,N_3054);
or U4849 (N_4849,N_2033,N_3010);
nand U4850 (N_4850,N_129,N_799);
and U4851 (N_4851,N_1027,N_585);
nor U4852 (N_4852,N_2862,N_2447);
nor U4853 (N_4853,N_1509,N_183);
xnor U4854 (N_4854,N_1381,N_614);
and U4855 (N_4855,N_800,N_1938);
and U4856 (N_4856,N_2505,N_2796);
nor U4857 (N_4857,N_1633,N_461);
and U4858 (N_4858,N_505,N_2651);
or U4859 (N_4859,N_508,N_1501);
xnor U4860 (N_4860,N_2601,N_2433);
xnor U4861 (N_4861,N_2371,N_1884);
and U4862 (N_4862,N_59,N_2805);
nor U4863 (N_4863,N_2726,N_1570);
or U4864 (N_4864,N_402,N_135);
nand U4865 (N_4865,N_2065,N_1189);
nand U4866 (N_4866,N_122,N_1869);
nor U4867 (N_4867,N_1931,N_1182);
and U4868 (N_4868,N_644,N_526);
nand U4869 (N_4869,N_768,N_3061);
nand U4870 (N_4870,N_2817,N_25);
or U4871 (N_4871,N_335,N_639);
nor U4872 (N_4872,N_1850,N_1157);
and U4873 (N_4873,N_3009,N_1561);
xnor U4874 (N_4874,N_1042,N_731);
xor U4875 (N_4875,N_2947,N_965);
xor U4876 (N_4876,N_2889,N_1145);
or U4877 (N_4877,N_854,N_2069);
or U4878 (N_4878,N_1881,N_2305);
or U4879 (N_4879,N_1994,N_2241);
and U4880 (N_4880,N_1783,N_662);
nand U4881 (N_4881,N_1924,N_69);
nand U4882 (N_4882,N_1886,N_466);
nor U4883 (N_4883,N_2339,N_1909);
nand U4884 (N_4884,N_2932,N_1754);
nand U4885 (N_4885,N_175,N_903);
and U4886 (N_4886,N_2982,N_2612);
nand U4887 (N_4887,N_1486,N_2180);
nand U4888 (N_4888,N_1826,N_2568);
nand U4889 (N_4889,N_1890,N_2137);
nand U4890 (N_4890,N_377,N_48);
nand U4891 (N_4891,N_144,N_1060);
nand U4892 (N_4892,N_1400,N_2643);
xnor U4893 (N_4893,N_2847,N_1919);
nor U4894 (N_4894,N_2404,N_739);
nor U4895 (N_4895,N_2487,N_2486);
or U4896 (N_4896,N_2038,N_2938);
or U4897 (N_4897,N_2774,N_2507);
and U4898 (N_4898,N_800,N_1784);
nand U4899 (N_4899,N_2237,N_2904);
xor U4900 (N_4900,N_2978,N_2450);
or U4901 (N_4901,N_2684,N_2273);
nand U4902 (N_4902,N_930,N_1543);
xor U4903 (N_4903,N_11,N_2246);
nor U4904 (N_4904,N_2683,N_3049);
or U4905 (N_4905,N_2734,N_1018);
or U4906 (N_4906,N_913,N_1259);
and U4907 (N_4907,N_868,N_2824);
or U4908 (N_4908,N_2354,N_41);
or U4909 (N_4909,N_3001,N_2697);
nor U4910 (N_4910,N_1321,N_1410);
nor U4911 (N_4911,N_76,N_469);
and U4912 (N_4912,N_2605,N_2572);
xor U4913 (N_4913,N_1316,N_2554);
or U4914 (N_4914,N_1845,N_2725);
nand U4915 (N_4915,N_1262,N_1733);
or U4916 (N_4916,N_2864,N_852);
nand U4917 (N_4917,N_2248,N_2778);
nand U4918 (N_4918,N_2148,N_1564);
xor U4919 (N_4919,N_369,N_1153);
nor U4920 (N_4920,N_933,N_879);
nand U4921 (N_4921,N_811,N_812);
nor U4922 (N_4922,N_430,N_2690);
and U4923 (N_4923,N_1924,N_1607);
or U4924 (N_4924,N_2110,N_2021);
or U4925 (N_4925,N_1603,N_2134);
or U4926 (N_4926,N_951,N_1985);
and U4927 (N_4927,N_909,N_1955);
nand U4928 (N_4928,N_2392,N_1145);
nand U4929 (N_4929,N_1167,N_740);
or U4930 (N_4930,N_2764,N_2563);
and U4931 (N_4931,N_334,N_2292);
and U4932 (N_4932,N_4,N_2344);
xnor U4933 (N_4933,N_1894,N_1351);
nor U4934 (N_4934,N_2986,N_1847);
or U4935 (N_4935,N_677,N_917);
nor U4936 (N_4936,N_1646,N_121);
or U4937 (N_4937,N_616,N_2770);
nand U4938 (N_4938,N_2012,N_1378);
and U4939 (N_4939,N_1676,N_2619);
and U4940 (N_4940,N_871,N_1573);
nand U4941 (N_4941,N_1544,N_967);
nand U4942 (N_4942,N_1940,N_1567);
nor U4943 (N_4943,N_1251,N_1106);
xnor U4944 (N_4944,N_2148,N_1459);
xnor U4945 (N_4945,N_1179,N_2100);
nand U4946 (N_4946,N_794,N_2954);
nor U4947 (N_4947,N_3085,N_2247);
nand U4948 (N_4948,N_758,N_2652);
nor U4949 (N_4949,N_1162,N_512);
and U4950 (N_4950,N_42,N_227);
xnor U4951 (N_4951,N_1088,N_451);
nor U4952 (N_4952,N_2455,N_2244);
nor U4953 (N_4953,N_2441,N_295);
nand U4954 (N_4954,N_1967,N_1122);
or U4955 (N_4955,N_2454,N_2061);
or U4956 (N_4956,N_621,N_2626);
nor U4957 (N_4957,N_1607,N_255);
nand U4958 (N_4958,N_2285,N_2728);
nand U4959 (N_4959,N_2103,N_3082);
or U4960 (N_4960,N_2535,N_445);
xor U4961 (N_4961,N_2519,N_2731);
nand U4962 (N_4962,N_1858,N_2538);
and U4963 (N_4963,N_938,N_1544);
and U4964 (N_4964,N_2767,N_2703);
nand U4965 (N_4965,N_1121,N_2224);
nor U4966 (N_4966,N_2962,N_2464);
nor U4967 (N_4967,N_864,N_1174);
or U4968 (N_4968,N_3011,N_81);
nor U4969 (N_4969,N_1961,N_2022);
nor U4970 (N_4970,N_2828,N_325);
xnor U4971 (N_4971,N_847,N_1555);
or U4972 (N_4972,N_513,N_158);
nor U4973 (N_4973,N_2189,N_1093);
nand U4974 (N_4974,N_2192,N_2549);
nor U4975 (N_4975,N_2082,N_477);
or U4976 (N_4976,N_534,N_1314);
and U4977 (N_4977,N_69,N_2209);
or U4978 (N_4978,N_3107,N_479);
xor U4979 (N_4979,N_228,N_2951);
or U4980 (N_4980,N_2748,N_996);
nand U4981 (N_4981,N_14,N_2157);
nand U4982 (N_4982,N_1818,N_2473);
xnor U4983 (N_4983,N_2026,N_595);
or U4984 (N_4984,N_2999,N_2618);
nand U4985 (N_4985,N_2208,N_987);
nor U4986 (N_4986,N_2023,N_1372);
and U4987 (N_4987,N_1309,N_732);
and U4988 (N_4988,N_908,N_2819);
or U4989 (N_4989,N_1659,N_1252);
nand U4990 (N_4990,N_2785,N_889);
and U4991 (N_4991,N_1240,N_1617);
and U4992 (N_4992,N_1305,N_1572);
or U4993 (N_4993,N_36,N_768);
xor U4994 (N_4994,N_910,N_1142);
and U4995 (N_4995,N_939,N_892);
nand U4996 (N_4996,N_2989,N_2244);
nor U4997 (N_4997,N_1350,N_670);
xnor U4998 (N_4998,N_272,N_3039);
and U4999 (N_4999,N_363,N_2005);
nand U5000 (N_5000,N_2640,N_2792);
nand U5001 (N_5001,N_2396,N_1931);
nand U5002 (N_5002,N_570,N_1509);
nand U5003 (N_5003,N_97,N_206);
and U5004 (N_5004,N_1697,N_1509);
nand U5005 (N_5005,N_1470,N_1675);
nor U5006 (N_5006,N_746,N_1973);
nor U5007 (N_5007,N_824,N_1746);
nand U5008 (N_5008,N_384,N_931);
nor U5009 (N_5009,N_48,N_2713);
nor U5010 (N_5010,N_2432,N_2549);
or U5011 (N_5011,N_2032,N_2817);
and U5012 (N_5012,N_1658,N_2044);
or U5013 (N_5013,N_767,N_2457);
nand U5014 (N_5014,N_538,N_1992);
or U5015 (N_5015,N_76,N_105);
or U5016 (N_5016,N_1807,N_2537);
or U5017 (N_5017,N_105,N_3049);
and U5018 (N_5018,N_593,N_2843);
nand U5019 (N_5019,N_1995,N_1016);
and U5020 (N_5020,N_859,N_1931);
xnor U5021 (N_5021,N_929,N_22);
nand U5022 (N_5022,N_2881,N_955);
and U5023 (N_5023,N_2151,N_2853);
xnor U5024 (N_5024,N_1229,N_2693);
and U5025 (N_5025,N_1284,N_2370);
and U5026 (N_5026,N_165,N_2457);
or U5027 (N_5027,N_2425,N_3041);
nand U5028 (N_5028,N_3103,N_690);
xnor U5029 (N_5029,N_1964,N_1072);
or U5030 (N_5030,N_1256,N_2783);
nor U5031 (N_5031,N_2675,N_31);
nand U5032 (N_5032,N_1523,N_1677);
and U5033 (N_5033,N_2670,N_2444);
or U5034 (N_5034,N_1839,N_527);
xnor U5035 (N_5035,N_2010,N_2814);
nand U5036 (N_5036,N_2886,N_1309);
or U5037 (N_5037,N_535,N_2798);
nand U5038 (N_5038,N_1176,N_2687);
or U5039 (N_5039,N_2068,N_2543);
or U5040 (N_5040,N_1054,N_2586);
nand U5041 (N_5041,N_1930,N_208);
nor U5042 (N_5042,N_608,N_1567);
nor U5043 (N_5043,N_1858,N_2573);
nor U5044 (N_5044,N_2679,N_2773);
nand U5045 (N_5045,N_1644,N_1026);
xnor U5046 (N_5046,N_2178,N_1188);
and U5047 (N_5047,N_1442,N_728);
or U5048 (N_5048,N_3021,N_1308);
nor U5049 (N_5049,N_351,N_2455);
nand U5050 (N_5050,N_1453,N_2493);
xor U5051 (N_5051,N_1331,N_2478);
and U5052 (N_5052,N_1590,N_2167);
xnor U5053 (N_5053,N_2899,N_350);
xor U5054 (N_5054,N_3048,N_50);
and U5055 (N_5055,N_2369,N_1877);
nand U5056 (N_5056,N_1979,N_2709);
or U5057 (N_5057,N_579,N_610);
nor U5058 (N_5058,N_2991,N_1435);
and U5059 (N_5059,N_411,N_2829);
and U5060 (N_5060,N_36,N_196);
and U5061 (N_5061,N_464,N_1767);
xnor U5062 (N_5062,N_2526,N_447);
xor U5063 (N_5063,N_688,N_3000);
nand U5064 (N_5064,N_796,N_313);
or U5065 (N_5065,N_843,N_221);
and U5066 (N_5066,N_2952,N_1599);
nand U5067 (N_5067,N_1894,N_1999);
or U5068 (N_5068,N_2647,N_2331);
nor U5069 (N_5069,N_1041,N_1452);
or U5070 (N_5070,N_818,N_1835);
nand U5071 (N_5071,N_674,N_459);
nor U5072 (N_5072,N_324,N_364);
nand U5073 (N_5073,N_2734,N_2320);
xor U5074 (N_5074,N_249,N_419);
nand U5075 (N_5075,N_1516,N_3065);
and U5076 (N_5076,N_2273,N_747);
nand U5077 (N_5077,N_727,N_2263);
or U5078 (N_5078,N_2965,N_1019);
xor U5079 (N_5079,N_404,N_3084);
or U5080 (N_5080,N_2780,N_1189);
nor U5081 (N_5081,N_2167,N_1099);
or U5082 (N_5082,N_1257,N_1849);
and U5083 (N_5083,N_735,N_987);
or U5084 (N_5084,N_2467,N_1198);
or U5085 (N_5085,N_2005,N_1907);
and U5086 (N_5086,N_2105,N_1782);
nand U5087 (N_5087,N_205,N_2310);
xor U5088 (N_5088,N_780,N_2275);
nor U5089 (N_5089,N_1000,N_899);
or U5090 (N_5090,N_1355,N_2678);
xor U5091 (N_5091,N_950,N_1221);
and U5092 (N_5092,N_1756,N_2444);
nand U5093 (N_5093,N_2435,N_1713);
xnor U5094 (N_5094,N_942,N_545);
xnor U5095 (N_5095,N_3006,N_2948);
nor U5096 (N_5096,N_680,N_2650);
or U5097 (N_5097,N_3006,N_1050);
and U5098 (N_5098,N_1028,N_2384);
nand U5099 (N_5099,N_1288,N_646);
xnor U5100 (N_5100,N_873,N_2356);
or U5101 (N_5101,N_2222,N_396);
or U5102 (N_5102,N_2814,N_2684);
xnor U5103 (N_5103,N_2374,N_3046);
xnor U5104 (N_5104,N_104,N_208);
or U5105 (N_5105,N_2662,N_1778);
or U5106 (N_5106,N_2788,N_2521);
nand U5107 (N_5107,N_1894,N_2321);
and U5108 (N_5108,N_2752,N_2101);
nand U5109 (N_5109,N_2711,N_528);
or U5110 (N_5110,N_2520,N_2352);
and U5111 (N_5111,N_2913,N_2450);
or U5112 (N_5112,N_262,N_1419);
nand U5113 (N_5113,N_591,N_604);
and U5114 (N_5114,N_1665,N_1182);
nand U5115 (N_5115,N_487,N_776);
xor U5116 (N_5116,N_339,N_2494);
or U5117 (N_5117,N_416,N_2581);
or U5118 (N_5118,N_2920,N_2346);
or U5119 (N_5119,N_3028,N_2947);
or U5120 (N_5120,N_867,N_3043);
nand U5121 (N_5121,N_1747,N_18);
nand U5122 (N_5122,N_536,N_686);
and U5123 (N_5123,N_676,N_2210);
nor U5124 (N_5124,N_1810,N_712);
nor U5125 (N_5125,N_1805,N_939);
or U5126 (N_5126,N_2977,N_2022);
or U5127 (N_5127,N_2329,N_1387);
or U5128 (N_5128,N_1788,N_1464);
and U5129 (N_5129,N_1748,N_288);
nand U5130 (N_5130,N_2736,N_1336);
xor U5131 (N_5131,N_3113,N_991);
nand U5132 (N_5132,N_1707,N_2348);
or U5133 (N_5133,N_867,N_285);
or U5134 (N_5134,N_2902,N_1367);
and U5135 (N_5135,N_2549,N_2543);
nand U5136 (N_5136,N_1082,N_1284);
nand U5137 (N_5137,N_2820,N_1189);
or U5138 (N_5138,N_467,N_3119);
nand U5139 (N_5139,N_72,N_1990);
or U5140 (N_5140,N_3029,N_254);
and U5141 (N_5141,N_1658,N_983);
nand U5142 (N_5142,N_3026,N_3009);
or U5143 (N_5143,N_2952,N_170);
or U5144 (N_5144,N_2919,N_2159);
and U5145 (N_5145,N_533,N_783);
xor U5146 (N_5146,N_2915,N_3016);
xnor U5147 (N_5147,N_931,N_591);
nor U5148 (N_5148,N_1585,N_1359);
or U5149 (N_5149,N_2506,N_2657);
nor U5150 (N_5150,N_386,N_3043);
and U5151 (N_5151,N_789,N_2376);
nand U5152 (N_5152,N_2340,N_1386);
or U5153 (N_5153,N_201,N_1195);
nor U5154 (N_5154,N_1696,N_1128);
and U5155 (N_5155,N_2352,N_543);
nand U5156 (N_5156,N_2586,N_2878);
xor U5157 (N_5157,N_2692,N_135);
nand U5158 (N_5158,N_539,N_2755);
and U5159 (N_5159,N_2785,N_1452);
nand U5160 (N_5160,N_2039,N_779);
and U5161 (N_5161,N_2719,N_2844);
nand U5162 (N_5162,N_1676,N_1379);
nand U5163 (N_5163,N_2243,N_2268);
xor U5164 (N_5164,N_266,N_390);
nand U5165 (N_5165,N_3093,N_2494);
xnor U5166 (N_5166,N_2588,N_1146);
and U5167 (N_5167,N_2219,N_557);
nor U5168 (N_5168,N_1066,N_2209);
nand U5169 (N_5169,N_1020,N_85);
nor U5170 (N_5170,N_987,N_749);
or U5171 (N_5171,N_2912,N_416);
and U5172 (N_5172,N_2616,N_1207);
or U5173 (N_5173,N_975,N_1197);
or U5174 (N_5174,N_795,N_2963);
or U5175 (N_5175,N_3051,N_2665);
xor U5176 (N_5176,N_164,N_1442);
xor U5177 (N_5177,N_550,N_827);
and U5178 (N_5178,N_2347,N_46);
or U5179 (N_5179,N_2657,N_1691);
nand U5180 (N_5180,N_3071,N_775);
and U5181 (N_5181,N_1945,N_84);
or U5182 (N_5182,N_263,N_1392);
xnor U5183 (N_5183,N_2311,N_1949);
nand U5184 (N_5184,N_775,N_751);
nor U5185 (N_5185,N_1419,N_404);
nand U5186 (N_5186,N_825,N_1563);
or U5187 (N_5187,N_2846,N_2466);
and U5188 (N_5188,N_2375,N_444);
and U5189 (N_5189,N_101,N_2743);
nand U5190 (N_5190,N_2758,N_930);
nand U5191 (N_5191,N_2811,N_3032);
and U5192 (N_5192,N_2458,N_2668);
xor U5193 (N_5193,N_161,N_3108);
and U5194 (N_5194,N_878,N_2026);
xor U5195 (N_5195,N_2780,N_209);
or U5196 (N_5196,N_3078,N_2562);
and U5197 (N_5197,N_2727,N_1914);
or U5198 (N_5198,N_2896,N_3067);
and U5199 (N_5199,N_2852,N_1136);
or U5200 (N_5200,N_2060,N_2249);
nor U5201 (N_5201,N_730,N_1005);
or U5202 (N_5202,N_1736,N_2293);
nand U5203 (N_5203,N_329,N_3112);
and U5204 (N_5204,N_624,N_891);
xor U5205 (N_5205,N_708,N_1065);
nor U5206 (N_5206,N_479,N_1683);
nand U5207 (N_5207,N_3043,N_2569);
or U5208 (N_5208,N_1399,N_355);
xnor U5209 (N_5209,N_2357,N_1496);
xor U5210 (N_5210,N_1095,N_2987);
nand U5211 (N_5211,N_969,N_1191);
nor U5212 (N_5212,N_122,N_2014);
or U5213 (N_5213,N_657,N_3123);
and U5214 (N_5214,N_431,N_21);
and U5215 (N_5215,N_1874,N_2581);
or U5216 (N_5216,N_3052,N_1101);
or U5217 (N_5217,N_8,N_1433);
or U5218 (N_5218,N_2857,N_1935);
or U5219 (N_5219,N_246,N_2531);
xnor U5220 (N_5220,N_1832,N_1482);
or U5221 (N_5221,N_2618,N_2514);
or U5222 (N_5222,N_2641,N_564);
nor U5223 (N_5223,N_1817,N_533);
nand U5224 (N_5224,N_901,N_438);
nor U5225 (N_5225,N_2908,N_2081);
nand U5226 (N_5226,N_1217,N_1236);
or U5227 (N_5227,N_1983,N_1396);
nand U5228 (N_5228,N_2823,N_714);
nor U5229 (N_5229,N_1863,N_2704);
nor U5230 (N_5230,N_344,N_2379);
nor U5231 (N_5231,N_1050,N_1787);
nor U5232 (N_5232,N_1599,N_1964);
nor U5233 (N_5233,N_2950,N_2545);
or U5234 (N_5234,N_2520,N_1776);
and U5235 (N_5235,N_1567,N_2586);
nand U5236 (N_5236,N_2902,N_2749);
xor U5237 (N_5237,N_543,N_226);
nand U5238 (N_5238,N_1382,N_1453);
nand U5239 (N_5239,N_428,N_630);
xnor U5240 (N_5240,N_3087,N_1419);
xnor U5241 (N_5241,N_229,N_867);
nor U5242 (N_5242,N_323,N_228);
or U5243 (N_5243,N_2888,N_863);
nand U5244 (N_5244,N_326,N_2761);
and U5245 (N_5245,N_587,N_408);
and U5246 (N_5246,N_1537,N_2727);
nand U5247 (N_5247,N_1101,N_2276);
or U5248 (N_5248,N_1727,N_544);
xnor U5249 (N_5249,N_1383,N_279);
nand U5250 (N_5250,N_2907,N_2135);
and U5251 (N_5251,N_1991,N_1349);
nand U5252 (N_5252,N_1305,N_493);
nand U5253 (N_5253,N_856,N_657);
nand U5254 (N_5254,N_2618,N_926);
nor U5255 (N_5255,N_1970,N_2032);
and U5256 (N_5256,N_2889,N_1846);
and U5257 (N_5257,N_2645,N_1322);
nor U5258 (N_5258,N_2672,N_1877);
and U5259 (N_5259,N_2063,N_2009);
nor U5260 (N_5260,N_2572,N_1506);
or U5261 (N_5261,N_1296,N_872);
and U5262 (N_5262,N_2237,N_2611);
nand U5263 (N_5263,N_1556,N_2629);
or U5264 (N_5264,N_906,N_2700);
or U5265 (N_5265,N_2248,N_2978);
xor U5266 (N_5266,N_2888,N_1631);
xnor U5267 (N_5267,N_2012,N_153);
nand U5268 (N_5268,N_2098,N_440);
or U5269 (N_5269,N_5,N_836);
nor U5270 (N_5270,N_2804,N_366);
nand U5271 (N_5271,N_1094,N_1837);
or U5272 (N_5272,N_1779,N_709);
and U5273 (N_5273,N_77,N_2174);
nand U5274 (N_5274,N_2560,N_1804);
and U5275 (N_5275,N_1753,N_6);
and U5276 (N_5276,N_584,N_601);
or U5277 (N_5277,N_3079,N_710);
and U5278 (N_5278,N_2085,N_1103);
nor U5279 (N_5279,N_2098,N_461);
or U5280 (N_5280,N_1568,N_2134);
nor U5281 (N_5281,N_132,N_2254);
xnor U5282 (N_5282,N_1286,N_299);
nand U5283 (N_5283,N_2008,N_1288);
nand U5284 (N_5284,N_116,N_1569);
nand U5285 (N_5285,N_198,N_889);
or U5286 (N_5286,N_2614,N_355);
nor U5287 (N_5287,N_2930,N_542);
or U5288 (N_5288,N_3088,N_2386);
and U5289 (N_5289,N_169,N_1503);
nor U5290 (N_5290,N_1338,N_2408);
and U5291 (N_5291,N_2381,N_2252);
nor U5292 (N_5292,N_1950,N_4);
or U5293 (N_5293,N_2496,N_2229);
nor U5294 (N_5294,N_1418,N_2895);
and U5295 (N_5295,N_3044,N_2977);
and U5296 (N_5296,N_757,N_1105);
and U5297 (N_5297,N_1267,N_520);
and U5298 (N_5298,N_2981,N_915);
nand U5299 (N_5299,N_863,N_2363);
or U5300 (N_5300,N_1622,N_1397);
xor U5301 (N_5301,N_1987,N_2702);
xnor U5302 (N_5302,N_855,N_2324);
nand U5303 (N_5303,N_733,N_1287);
xor U5304 (N_5304,N_1040,N_579);
nand U5305 (N_5305,N_1660,N_1412);
nor U5306 (N_5306,N_2326,N_1717);
or U5307 (N_5307,N_1665,N_2471);
nand U5308 (N_5308,N_825,N_1079);
xnor U5309 (N_5309,N_588,N_2989);
nor U5310 (N_5310,N_2439,N_2569);
or U5311 (N_5311,N_211,N_32);
nand U5312 (N_5312,N_2291,N_449);
or U5313 (N_5313,N_2367,N_1256);
or U5314 (N_5314,N_2005,N_1033);
nand U5315 (N_5315,N_477,N_184);
xor U5316 (N_5316,N_1293,N_973);
nand U5317 (N_5317,N_2929,N_95);
xor U5318 (N_5318,N_2214,N_2906);
nor U5319 (N_5319,N_2332,N_2798);
xnor U5320 (N_5320,N_1736,N_1537);
or U5321 (N_5321,N_1715,N_1523);
nor U5322 (N_5322,N_2066,N_220);
nor U5323 (N_5323,N_1609,N_404);
nand U5324 (N_5324,N_2328,N_1820);
xnor U5325 (N_5325,N_1243,N_1519);
and U5326 (N_5326,N_1269,N_433);
xnor U5327 (N_5327,N_2108,N_1957);
nand U5328 (N_5328,N_1367,N_500);
and U5329 (N_5329,N_3018,N_1527);
nand U5330 (N_5330,N_781,N_402);
and U5331 (N_5331,N_2493,N_295);
xor U5332 (N_5332,N_3111,N_1010);
xnor U5333 (N_5333,N_2048,N_1273);
nand U5334 (N_5334,N_2190,N_974);
xor U5335 (N_5335,N_1068,N_2850);
nor U5336 (N_5336,N_87,N_1476);
and U5337 (N_5337,N_689,N_801);
and U5338 (N_5338,N_2942,N_450);
or U5339 (N_5339,N_1712,N_1703);
and U5340 (N_5340,N_889,N_1951);
xor U5341 (N_5341,N_1351,N_1467);
nor U5342 (N_5342,N_560,N_2380);
and U5343 (N_5343,N_1386,N_3038);
nand U5344 (N_5344,N_1301,N_1677);
nand U5345 (N_5345,N_980,N_1795);
xnor U5346 (N_5346,N_1218,N_441);
nor U5347 (N_5347,N_2101,N_2240);
nor U5348 (N_5348,N_2479,N_2141);
nand U5349 (N_5349,N_2312,N_1772);
nor U5350 (N_5350,N_2805,N_1832);
and U5351 (N_5351,N_2720,N_2864);
and U5352 (N_5352,N_612,N_2134);
nor U5353 (N_5353,N_2967,N_2869);
or U5354 (N_5354,N_37,N_3044);
xnor U5355 (N_5355,N_972,N_2817);
xnor U5356 (N_5356,N_482,N_989);
nand U5357 (N_5357,N_116,N_2294);
and U5358 (N_5358,N_3043,N_250);
or U5359 (N_5359,N_2188,N_389);
or U5360 (N_5360,N_1680,N_2294);
nand U5361 (N_5361,N_1656,N_491);
xnor U5362 (N_5362,N_1467,N_1216);
nor U5363 (N_5363,N_350,N_2483);
nand U5364 (N_5364,N_496,N_2812);
and U5365 (N_5365,N_1645,N_1846);
and U5366 (N_5366,N_1410,N_2491);
or U5367 (N_5367,N_1032,N_906);
and U5368 (N_5368,N_2312,N_2419);
nand U5369 (N_5369,N_1406,N_45);
or U5370 (N_5370,N_908,N_1702);
or U5371 (N_5371,N_146,N_1459);
nor U5372 (N_5372,N_883,N_804);
nor U5373 (N_5373,N_2405,N_2328);
nand U5374 (N_5374,N_965,N_1485);
and U5375 (N_5375,N_2854,N_2547);
nand U5376 (N_5376,N_1763,N_2262);
nor U5377 (N_5377,N_1657,N_1041);
and U5378 (N_5378,N_2615,N_1526);
or U5379 (N_5379,N_1899,N_3063);
xnor U5380 (N_5380,N_424,N_2038);
nand U5381 (N_5381,N_2479,N_410);
or U5382 (N_5382,N_2475,N_255);
or U5383 (N_5383,N_1800,N_1806);
nand U5384 (N_5384,N_2796,N_1527);
nand U5385 (N_5385,N_1100,N_1244);
xnor U5386 (N_5386,N_967,N_1824);
and U5387 (N_5387,N_879,N_2659);
or U5388 (N_5388,N_2375,N_3029);
or U5389 (N_5389,N_144,N_3089);
xnor U5390 (N_5390,N_2333,N_3100);
and U5391 (N_5391,N_2472,N_2507);
nand U5392 (N_5392,N_1320,N_808);
xnor U5393 (N_5393,N_1589,N_1083);
nand U5394 (N_5394,N_73,N_1914);
nand U5395 (N_5395,N_1333,N_1366);
nor U5396 (N_5396,N_2580,N_2649);
and U5397 (N_5397,N_1258,N_1743);
xnor U5398 (N_5398,N_362,N_282);
or U5399 (N_5399,N_2674,N_704);
xor U5400 (N_5400,N_954,N_2537);
nand U5401 (N_5401,N_2669,N_1306);
xnor U5402 (N_5402,N_10,N_2000);
nor U5403 (N_5403,N_1253,N_1927);
nand U5404 (N_5404,N_117,N_835);
or U5405 (N_5405,N_1831,N_2096);
xnor U5406 (N_5406,N_488,N_1477);
and U5407 (N_5407,N_306,N_522);
or U5408 (N_5408,N_518,N_1500);
and U5409 (N_5409,N_1419,N_2072);
xnor U5410 (N_5410,N_1733,N_256);
xor U5411 (N_5411,N_1547,N_1020);
or U5412 (N_5412,N_1373,N_249);
or U5413 (N_5413,N_896,N_2735);
and U5414 (N_5414,N_637,N_2139);
or U5415 (N_5415,N_2447,N_1873);
xnor U5416 (N_5416,N_2796,N_894);
nand U5417 (N_5417,N_953,N_437);
or U5418 (N_5418,N_1713,N_194);
nor U5419 (N_5419,N_1012,N_1880);
nand U5420 (N_5420,N_2698,N_193);
xor U5421 (N_5421,N_1292,N_697);
or U5422 (N_5422,N_829,N_762);
nor U5423 (N_5423,N_634,N_2673);
nor U5424 (N_5424,N_2349,N_1838);
nand U5425 (N_5425,N_303,N_3021);
nor U5426 (N_5426,N_2369,N_1274);
nand U5427 (N_5427,N_337,N_2779);
xor U5428 (N_5428,N_1467,N_1461);
or U5429 (N_5429,N_1512,N_512);
and U5430 (N_5430,N_969,N_2347);
nor U5431 (N_5431,N_1493,N_1047);
nand U5432 (N_5432,N_2815,N_2305);
nor U5433 (N_5433,N_2235,N_1147);
and U5434 (N_5434,N_2545,N_3021);
nand U5435 (N_5435,N_122,N_2087);
nor U5436 (N_5436,N_261,N_2781);
nor U5437 (N_5437,N_935,N_430);
and U5438 (N_5438,N_532,N_233);
or U5439 (N_5439,N_620,N_1226);
nand U5440 (N_5440,N_42,N_1530);
or U5441 (N_5441,N_2668,N_8);
nand U5442 (N_5442,N_2847,N_1569);
nor U5443 (N_5443,N_1475,N_3001);
xnor U5444 (N_5444,N_2898,N_1612);
and U5445 (N_5445,N_2331,N_1831);
nand U5446 (N_5446,N_1663,N_2693);
xnor U5447 (N_5447,N_625,N_1983);
nor U5448 (N_5448,N_683,N_831);
xnor U5449 (N_5449,N_2214,N_97);
nand U5450 (N_5450,N_22,N_2253);
nor U5451 (N_5451,N_1368,N_1789);
xor U5452 (N_5452,N_703,N_2812);
nor U5453 (N_5453,N_911,N_1251);
nor U5454 (N_5454,N_1849,N_2128);
nor U5455 (N_5455,N_3100,N_318);
and U5456 (N_5456,N_2385,N_1843);
and U5457 (N_5457,N_606,N_132);
xnor U5458 (N_5458,N_2070,N_2029);
or U5459 (N_5459,N_391,N_2337);
nor U5460 (N_5460,N_2628,N_2379);
nand U5461 (N_5461,N_2333,N_1484);
xor U5462 (N_5462,N_1239,N_56);
or U5463 (N_5463,N_1222,N_2929);
xor U5464 (N_5464,N_1391,N_1890);
nor U5465 (N_5465,N_2734,N_2645);
or U5466 (N_5466,N_2574,N_36);
xor U5467 (N_5467,N_1974,N_219);
nand U5468 (N_5468,N_2586,N_1700);
xor U5469 (N_5469,N_2727,N_1511);
nand U5470 (N_5470,N_830,N_921);
xor U5471 (N_5471,N_1710,N_2013);
nor U5472 (N_5472,N_1964,N_931);
and U5473 (N_5473,N_2734,N_2866);
nor U5474 (N_5474,N_422,N_843);
nand U5475 (N_5475,N_2077,N_535);
or U5476 (N_5476,N_2179,N_543);
nand U5477 (N_5477,N_991,N_2227);
and U5478 (N_5478,N_695,N_1817);
nor U5479 (N_5479,N_756,N_2722);
or U5480 (N_5480,N_2899,N_1596);
nand U5481 (N_5481,N_862,N_856);
nand U5482 (N_5482,N_138,N_1444);
xnor U5483 (N_5483,N_417,N_2061);
xor U5484 (N_5484,N_1996,N_1769);
nor U5485 (N_5485,N_1608,N_2104);
or U5486 (N_5486,N_2075,N_2739);
and U5487 (N_5487,N_2381,N_2803);
nand U5488 (N_5488,N_387,N_1028);
nand U5489 (N_5489,N_2750,N_1052);
xor U5490 (N_5490,N_1795,N_1998);
xnor U5491 (N_5491,N_392,N_1092);
xor U5492 (N_5492,N_2771,N_2845);
nor U5493 (N_5493,N_1745,N_1663);
and U5494 (N_5494,N_1598,N_1453);
nor U5495 (N_5495,N_2328,N_753);
xor U5496 (N_5496,N_612,N_475);
nand U5497 (N_5497,N_2245,N_1347);
nor U5498 (N_5498,N_2321,N_957);
nand U5499 (N_5499,N_171,N_2012);
nand U5500 (N_5500,N_2202,N_1041);
xor U5501 (N_5501,N_2879,N_2701);
or U5502 (N_5502,N_289,N_2955);
nor U5503 (N_5503,N_2166,N_1677);
or U5504 (N_5504,N_701,N_2172);
xor U5505 (N_5505,N_82,N_1741);
nand U5506 (N_5506,N_1303,N_2879);
xnor U5507 (N_5507,N_2633,N_1099);
and U5508 (N_5508,N_1123,N_1915);
and U5509 (N_5509,N_3021,N_2601);
nand U5510 (N_5510,N_704,N_1588);
and U5511 (N_5511,N_1845,N_1740);
xnor U5512 (N_5512,N_2854,N_1950);
and U5513 (N_5513,N_1838,N_419);
or U5514 (N_5514,N_304,N_916);
nor U5515 (N_5515,N_25,N_2369);
nor U5516 (N_5516,N_183,N_600);
and U5517 (N_5517,N_1535,N_1926);
and U5518 (N_5518,N_101,N_2);
or U5519 (N_5519,N_2602,N_704);
and U5520 (N_5520,N_2651,N_2748);
or U5521 (N_5521,N_2650,N_2243);
nand U5522 (N_5522,N_764,N_1592);
nor U5523 (N_5523,N_2720,N_500);
nor U5524 (N_5524,N_1101,N_96);
nand U5525 (N_5525,N_571,N_2128);
xor U5526 (N_5526,N_2552,N_2512);
xnor U5527 (N_5527,N_1556,N_1983);
and U5528 (N_5528,N_1544,N_803);
or U5529 (N_5529,N_2461,N_1018);
nor U5530 (N_5530,N_2758,N_1699);
xnor U5531 (N_5531,N_954,N_2926);
nand U5532 (N_5532,N_730,N_378);
and U5533 (N_5533,N_432,N_1212);
nor U5534 (N_5534,N_359,N_865);
xnor U5535 (N_5535,N_1027,N_2503);
xor U5536 (N_5536,N_1108,N_3066);
xnor U5537 (N_5537,N_1562,N_992);
xor U5538 (N_5538,N_590,N_2058);
and U5539 (N_5539,N_1116,N_964);
xnor U5540 (N_5540,N_229,N_1998);
or U5541 (N_5541,N_2191,N_680);
nor U5542 (N_5542,N_937,N_581);
xnor U5543 (N_5543,N_2035,N_1493);
nor U5544 (N_5544,N_2269,N_1049);
nand U5545 (N_5545,N_55,N_1652);
nor U5546 (N_5546,N_2783,N_1802);
or U5547 (N_5547,N_3040,N_1309);
and U5548 (N_5548,N_900,N_1617);
xnor U5549 (N_5549,N_466,N_941);
nor U5550 (N_5550,N_71,N_1013);
nor U5551 (N_5551,N_2301,N_71);
nand U5552 (N_5552,N_1778,N_2375);
nor U5553 (N_5553,N_1029,N_2942);
nor U5554 (N_5554,N_561,N_840);
nand U5555 (N_5555,N_1529,N_2373);
or U5556 (N_5556,N_1605,N_3082);
nor U5557 (N_5557,N_2988,N_2752);
or U5558 (N_5558,N_2167,N_1467);
and U5559 (N_5559,N_976,N_865);
xor U5560 (N_5560,N_2266,N_3026);
nand U5561 (N_5561,N_1862,N_2657);
nor U5562 (N_5562,N_66,N_2513);
and U5563 (N_5563,N_855,N_968);
xnor U5564 (N_5564,N_208,N_2095);
and U5565 (N_5565,N_582,N_2896);
nor U5566 (N_5566,N_2693,N_2086);
nand U5567 (N_5567,N_1577,N_1948);
or U5568 (N_5568,N_935,N_2711);
or U5569 (N_5569,N_2370,N_466);
nand U5570 (N_5570,N_1362,N_851);
nor U5571 (N_5571,N_216,N_2836);
xnor U5572 (N_5572,N_15,N_1943);
nor U5573 (N_5573,N_1566,N_658);
or U5574 (N_5574,N_1709,N_2850);
xnor U5575 (N_5575,N_1364,N_1401);
xor U5576 (N_5576,N_2756,N_2225);
and U5577 (N_5577,N_1796,N_1127);
or U5578 (N_5578,N_2134,N_1695);
xnor U5579 (N_5579,N_1479,N_1039);
xnor U5580 (N_5580,N_906,N_497);
nor U5581 (N_5581,N_1732,N_785);
xor U5582 (N_5582,N_638,N_587);
nor U5583 (N_5583,N_71,N_1052);
and U5584 (N_5584,N_1861,N_831);
nor U5585 (N_5585,N_439,N_1415);
and U5586 (N_5586,N_795,N_1108);
nand U5587 (N_5587,N_1419,N_3115);
xor U5588 (N_5588,N_353,N_205);
and U5589 (N_5589,N_1892,N_168);
or U5590 (N_5590,N_2805,N_391);
nand U5591 (N_5591,N_2754,N_2595);
or U5592 (N_5592,N_2538,N_1802);
nor U5593 (N_5593,N_2049,N_1536);
nor U5594 (N_5594,N_799,N_1347);
nor U5595 (N_5595,N_2279,N_1608);
xor U5596 (N_5596,N_2032,N_2249);
or U5597 (N_5597,N_2494,N_2908);
xnor U5598 (N_5598,N_1997,N_97);
nor U5599 (N_5599,N_1341,N_1682);
nand U5600 (N_5600,N_2178,N_2909);
xor U5601 (N_5601,N_3109,N_811);
nand U5602 (N_5602,N_1548,N_1571);
nor U5603 (N_5603,N_2180,N_383);
xnor U5604 (N_5604,N_1452,N_469);
or U5605 (N_5605,N_2035,N_2905);
xnor U5606 (N_5606,N_1705,N_1046);
and U5607 (N_5607,N_1385,N_2552);
nor U5608 (N_5608,N_1527,N_1587);
xnor U5609 (N_5609,N_1945,N_2068);
nor U5610 (N_5610,N_419,N_1410);
or U5611 (N_5611,N_1136,N_545);
nor U5612 (N_5612,N_2851,N_3033);
nor U5613 (N_5613,N_823,N_2667);
or U5614 (N_5614,N_2381,N_735);
xnor U5615 (N_5615,N_3122,N_2388);
or U5616 (N_5616,N_2945,N_1934);
nor U5617 (N_5617,N_142,N_2685);
xnor U5618 (N_5618,N_2580,N_511);
and U5619 (N_5619,N_2543,N_794);
and U5620 (N_5620,N_1354,N_791);
and U5621 (N_5621,N_135,N_1956);
xnor U5622 (N_5622,N_3000,N_2883);
xnor U5623 (N_5623,N_1120,N_111);
nand U5624 (N_5624,N_101,N_2708);
and U5625 (N_5625,N_42,N_556);
nor U5626 (N_5626,N_1725,N_3090);
nand U5627 (N_5627,N_224,N_55);
nand U5628 (N_5628,N_922,N_792);
and U5629 (N_5629,N_3081,N_983);
nor U5630 (N_5630,N_2115,N_1259);
nand U5631 (N_5631,N_1620,N_1426);
xnor U5632 (N_5632,N_2196,N_1835);
and U5633 (N_5633,N_2626,N_328);
xor U5634 (N_5634,N_1216,N_168);
xor U5635 (N_5635,N_1135,N_2165);
nand U5636 (N_5636,N_2162,N_2447);
and U5637 (N_5637,N_1248,N_2429);
xor U5638 (N_5638,N_2410,N_1172);
nand U5639 (N_5639,N_2548,N_2234);
or U5640 (N_5640,N_3013,N_209);
xnor U5641 (N_5641,N_31,N_1407);
nor U5642 (N_5642,N_3071,N_1809);
or U5643 (N_5643,N_1401,N_969);
nor U5644 (N_5644,N_748,N_1772);
or U5645 (N_5645,N_27,N_1498);
nand U5646 (N_5646,N_1029,N_2078);
or U5647 (N_5647,N_2149,N_2773);
or U5648 (N_5648,N_955,N_311);
and U5649 (N_5649,N_606,N_229);
or U5650 (N_5650,N_779,N_61);
or U5651 (N_5651,N_3051,N_162);
and U5652 (N_5652,N_1599,N_1096);
or U5653 (N_5653,N_41,N_648);
or U5654 (N_5654,N_1794,N_2898);
nor U5655 (N_5655,N_905,N_1256);
and U5656 (N_5656,N_2298,N_1840);
nand U5657 (N_5657,N_2990,N_1717);
nor U5658 (N_5658,N_1034,N_1264);
nand U5659 (N_5659,N_1844,N_2612);
xnor U5660 (N_5660,N_1887,N_2888);
nand U5661 (N_5661,N_1193,N_23);
or U5662 (N_5662,N_624,N_2052);
xor U5663 (N_5663,N_1007,N_2552);
nor U5664 (N_5664,N_2798,N_536);
nand U5665 (N_5665,N_511,N_3046);
xnor U5666 (N_5666,N_1576,N_1530);
nor U5667 (N_5667,N_1107,N_2636);
and U5668 (N_5668,N_665,N_2149);
nor U5669 (N_5669,N_3051,N_1134);
nor U5670 (N_5670,N_2129,N_2234);
xor U5671 (N_5671,N_2256,N_2176);
nor U5672 (N_5672,N_2943,N_1727);
nor U5673 (N_5673,N_2397,N_266);
nand U5674 (N_5674,N_592,N_1928);
nor U5675 (N_5675,N_2746,N_375);
and U5676 (N_5676,N_2514,N_352);
xnor U5677 (N_5677,N_2259,N_645);
nand U5678 (N_5678,N_1288,N_267);
xnor U5679 (N_5679,N_1326,N_2531);
nor U5680 (N_5680,N_2465,N_21);
nor U5681 (N_5681,N_2309,N_1277);
nand U5682 (N_5682,N_203,N_1933);
or U5683 (N_5683,N_1385,N_621);
or U5684 (N_5684,N_2620,N_1635);
xnor U5685 (N_5685,N_1301,N_516);
nor U5686 (N_5686,N_2123,N_492);
or U5687 (N_5687,N_1610,N_2988);
xnor U5688 (N_5688,N_1353,N_2468);
and U5689 (N_5689,N_2178,N_239);
and U5690 (N_5690,N_3034,N_2733);
nand U5691 (N_5691,N_775,N_1975);
xnor U5692 (N_5692,N_573,N_667);
xor U5693 (N_5693,N_812,N_2959);
or U5694 (N_5694,N_234,N_2265);
xor U5695 (N_5695,N_2740,N_3049);
nand U5696 (N_5696,N_275,N_2070);
and U5697 (N_5697,N_1470,N_391);
nand U5698 (N_5698,N_104,N_3110);
or U5699 (N_5699,N_326,N_883);
nand U5700 (N_5700,N_2193,N_1502);
xor U5701 (N_5701,N_1556,N_267);
nor U5702 (N_5702,N_1572,N_3014);
or U5703 (N_5703,N_19,N_1053);
or U5704 (N_5704,N_867,N_1340);
or U5705 (N_5705,N_2585,N_128);
xnor U5706 (N_5706,N_724,N_2514);
and U5707 (N_5707,N_3056,N_2938);
nand U5708 (N_5708,N_2472,N_624);
nand U5709 (N_5709,N_1059,N_2027);
and U5710 (N_5710,N_772,N_1307);
nand U5711 (N_5711,N_1662,N_1961);
and U5712 (N_5712,N_2610,N_1440);
xor U5713 (N_5713,N_283,N_1919);
and U5714 (N_5714,N_136,N_244);
or U5715 (N_5715,N_1718,N_885);
xnor U5716 (N_5716,N_1827,N_1973);
nand U5717 (N_5717,N_2477,N_1602);
xnor U5718 (N_5718,N_2396,N_1463);
nor U5719 (N_5719,N_1778,N_2733);
xnor U5720 (N_5720,N_899,N_1899);
nor U5721 (N_5721,N_1469,N_2516);
and U5722 (N_5722,N_1659,N_1639);
xnor U5723 (N_5723,N_1056,N_3071);
or U5724 (N_5724,N_1172,N_2004);
and U5725 (N_5725,N_1473,N_1439);
or U5726 (N_5726,N_1885,N_2972);
nand U5727 (N_5727,N_1376,N_1665);
nor U5728 (N_5728,N_2662,N_637);
or U5729 (N_5729,N_2913,N_1322);
and U5730 (N_5730,N_915,N_1308);
nand U5731 (N_5731,N_2041,N_462);
xor U5732 (N_5732,N_922,N_3);
nand U5733 (N_5733,N_1199,N_835);
or U5734 (N_5734,N_244,N_1521);
and U5735 (N_5735,N_2692,N_475);
xnor U5736 (N_5736,N_2104,N_1954);
nand U5737 (N_5737,N_1730,N_377);
xor U5738 (N_5738,N_3072,N_2721);
xor U5739 (N_5739,N_1467,N_1752);
xor U5740 (N_5740,N_1662,N_2309);
or U5741 (N_5741,N_2287,N_2741);
or U5742 (N_5742,N_1608,N_2567);
and U5743 (N_5743,N_2610,N_1433);
xnor U5744 (N_5744,N_286,N_2797);
nand U5745 (N_5745,N_139,N_2620);
or U5746 (N_5746,N_1139,N_2270);
xor U5747 (N_5747,N_1746,N_2697);
or U5748 (N_5748,N_2495,N_328);
or U5749 (N_5749,N_2003,N_749);
xnor U5750 (N_5750,N_2479,N_2126);
nand U5751 (N_5751,N_2408,N_1721);
xnor U5752 (N_5752,N_98,N_1086);
nand U5753 (N_5753,N_1489,N_2556);
nor U5754 (N_5754,N_1532,N_1944);
and U5755 (N_5755,N_2825,N_2546);
or U5756 (N_5756,N_731,N_2469);
nand U5757 (N_5757,N_923,N_2948);
nand U5758 (N_5758,N_283,N_1092);
nand U5759 (N_5759,N_1259,N_2984);
nand U5760 (N_5760,N_1792,N_31);
nand U5761 (N_5761,N_2005,N_1238);
or U5762 (N_5762,N_2535,N_2514);
and U5763 (N_5763,N_134,N_2101);
xnor U5764 (N_5764,N_472,N_3029);
nor U5765 (N_5765,N_1908,N_2274);
nor U5766 (N_5766,N_1990,N_1790);
and U5767 (N_5767,N_1041,N_2987);
or U5768 (N_5768,N_1007,N_1478);
nor U5769 (N_5769,N_1156,N_286);
xor U5770 (N_5770,N_2860,N_1253);
or U5771 (N_5771,N_1682,N_1233);
or U5772 (N_5772,N_1055,N_484);
nand U5773 (N_5773,N_1191,N_2171);
nor U5774 (N_5774,N_489,N_1120);
nand U5775 (N_5775,N_2318,N_331);
or U5776 (N_5776,N_1364,N_1061);
nor U5777 (N_5777,N_342,N_2812);
xnor U5778 (N_5778,N_1923,N_1351);
nor U5779 (N_5779,N_826,N_2285);
nor U5780 (N_5780,N_1138,N_489);
xnor U5781 (N_5781,N_2265,N_2273);
and U5782 (N_5782,N_2861,N_1013);
xnor U5783 (N_5783,N_142,N_1097);
or U5784 (N_5784,N_1243,N_2661);
nor U5785 (N_5785,N_2863,N_1614);
and U5786 (N_5786,N_1337,N_157);
xor U5787 (N_5787,N_2560,N_535);
nand U5788 (N_5788,N_2125,N_1556);
or U5789 (N_5789,N_1521,N_750);
nand U5790 (N_5790,N_2713,N_699);
and U5791 (N_5791,N_2173,N_2600);
or U5792 (N_5792,N_1842,N_3041);
nor U5793 (N_5793,N_1086,N_331);
or U5794 (N_5794,N_2587,N_2300);
or U5795 (N_5795,N_390,N_1037);
nor U5796 (N_5796,N_1590,N_1401);
xor U5797 (N_5797,N_1992,N_1474);
nor U5798 (N_5798,N_2039,N_2431);
and U5799 (N_5799,N_1856,N_2295);
and U5800 (N_5800,N_1768,N_1067);
and U5801 (N_5801,N_3031,N_2658);
nor U5802 (N_5802,N_276,N_2245);
or U5803 (N_5803,N_2120,N_2345);
and U5804 (N_5804,N_2872,N_3101);
nor U5805 (N_5805,N_1893,N_1383);
nand U5806 (N_5806,N_900,N_2703);
or U5807 (N_5807,N_109,N_298);
or U5808 (N_5808,N_2542,N_1626);
nor U5809 (N_5809,N_2514,N_711);
nand U5810 (N_5810,N_2478,N_1562);
or U5811 (N_5811,N_1722,N_740);
nand U5812 (N_5812,N_2697,N_11);
nand U5813 (N_5813,N_479,N_1020);
xor U5814 (N_5814,N_1360,N_204);
and U5815 (N_5815,N_2777,N_1659);
nor U5816 (N_5816,N_333,N_1324);
nand U5817 (N_5817,N_195,N_1850);
and U5818 (N_5818,N_776,N_2349);
nand U5819 (N_5819,N_1675,N_1225);
xnor U5820 (N_5820,N_356,N_2073);
xor U5821 (N_5821,N_770,N_164);
nor U5822 (N_5822,N_330,N_1080);
and U5823 (N_5823,N_2304,N_2675);
or U5824 (N_5824,N_1055,N_673);
nand U5825 (N_5825,N_302,N_1856);
and U5826 (N_5826,N_954,N_1252);
or U5827 (N_5827,N_1366,N_1248);
nand U5828 (N_5828,N_460,N_2422);
nor U5829 (N_5829,N_422,N_3036);
and U5830 (N_5830,N_1525,N_178);
nor U5831 (N_5831,N_1327,N_265);
and U5832 (N_5832,N_1033,N_285);
or U5833 (N_5833,N_1450,N_2135);
nor U5834 (N_5834,N_601,N_741);
xor U5835 (N_5835,N_2656,N_2337);
and U5836 (N_5836,N_848,N_69);
xnor U5837 (N_5837,N_885,N_152);
nand U5838 (N_5838,N_2272,N_1683);
and U5839 (N_5839,N_3050,N_2495);
nor U5840 (N_5840,N_749,N_635);
nand U5841 (N_5841,N_2684,N_280);
nor U5842 (N_5842,N_1662,N_873);
and U5843 (N_5843,N_1655,N_3009);
nand U5844 (N_5844,N_1325,N_88);
nand U5845 (N_5845,N_337,N_1582);
or U5846 (N_5846,N_1050,N_2698);
or U5847 (N_5847,N_1311,N_2305);
or U5848 (N_5848,N_856,N_2819);
or U5849 (N_5849,N_1398,N_1245);
and U5850 (N_5850,N_2782,N_1201);
or U5851 (N_5851,N_2858,N_2199);
nor U5852 (N_5852,N_1989,N_252);
or U5853 (N_5853,N_2276,N_84);
or U5854 (N_5854,N_2813,N_1948);
xor U5855 (N_5855,N_2590,N_1932);
or U5856 (N_5856,N_1330,N_2525);
nand U5857 (N_5857,N_451,N_311);
or U5858 (N_5858,N_1421,N_1726);
nor U5859 (N_5859,N_1186,N_3086);
and U5860 (N_5860,N_1620,N_2064);
nor U5861 (N_5861,N_1131,N_785);
or U5862 (N_5862,N_115,N_698);
nor U5863 (N_5863,N_687,N_464);
nor U5864 (N_5864,N_768,N_785);
xor U5865 (N_5865,N_3049,N_1634);
nor U5866 (N_5866,N_945,N_1280);
nor U5867 (N_5867,N_161,N_1407);
and U5868 (N_5868,N_2673,N_2938);
nor U5869 (N_5869,N_203,N_1009);
nand U5870 (N_5870,N_297,N_1506);
nor U5871 (N_5871,N_450,N_2524);
xor U5872 (N_5872,N_2570,N_968);
nor U5873 (N_5873,N_929,N_940);
and U5874 (N_5874,N_2068,N_1961);
xnor U5875 (N_5875,N_532,N_1076);
and U5876 (N_5876,N_2743,N_426);
xnor U5877 (N_5877,N_2365,N_625);
xor U5878 (N_5878,N_2632,N_1561);
and U5879 (N_5879,N_2048,N_2971);
nor U5880 (N_5880,N_292,N_1545);
xnor U5881 (N_5881,N_1354,N_1436);
xnor U5882 (N_5882,N_942,N_1943);
nor U5883 (N_5883,N_3017,N_2025);
or U5884 (N_5884,N_2511,N_2818);
or U5885 (N_5885,N_2607,N_524);
nor U5886 (N_5886,N_407,N_23);
nor U5887 (N_5887,N_420,N_1123);
and U5888 (N_5888,N_2540,N_2065);
nor U5889 (N_5889,N_1218,N_1988);
nand U5890 (N_5890,N_905,N_2311);
xor U5891 (N_5891,N_1205,N_76);
and U5892 (N_5892,N_199,N_1512);
and U5893 (N_5893,N_40,N_1767);
nand U5894 (N_5894,N_426,N_2223);
xor U5895 (N_5895,N_2644,N_2178);
xnor U5896 (N_5896,N_421,N_1627);
xnor U5897 (N_5897,N_350,N_3003);
nor U5898 (N_5898,N_2628,N_11);
and U5899 (N_5899,N_3046,N_1115);
nand U5900 (N_5900,N_368,N_1749);
nand U5901 (N_5901,N_96,N_267);
xnor U5902 (N_5902,N_2633,N_431);
nor U5903 (N_5903,N_423,N_242);
and U5904 (N_5904,N_637,N_2958);
and U5905 (N_5905,N_2976,N_482);
xnor U5906 (N_5906,N_1657,N_436);
xor U5907 (N_5907,N_217,N_3113);
or U5908 (N_5908,N_2753,N_254);
nor U5909 (N_5909,N_501,N_1545);
or U5910 (N_5910,N_1616,N_558);
and U5911 (N_5911,N_2913,N_1670);
or U5912 (N_5912,N_2979,N_1636);
xnor U5913 (N_5913,N_973,N_50);
nand U5914 (N_5914,N_1609,N_1157);
nand U5915 (N_5915,N_2878,N_678);
xnor U5916 (N_5916,N_630,N_1637);
and U5917 (N_5917,N_1465,N_644);
nor U5918 (N_5918,N_1581,N_338);
xnor U5919 (N_5919,N_345,N_2343);
nand U5920 (N_5920,N_1841,N_3122);
xnor U5921 (N_5921,N_126,N_2424);
nor U5922 (N_5922,N_1397,N_1436);
and U5923 (N_5923,N_674,N_936);
xor U5924 (N_5924,N_117,N_1109);
nand U5925 (N_5925,N_2844,N_2046);
xor U5926 (N_5926,N_364,N_1388);
or U5927 (N_5927,N_778,N_1119);
nand U5928 (N_5928,N_1979,N_2453);
xnor U5929 (N_5929,N_1502,N_360);
nand U5930 (N_5930,N_1001,N_2715);
and U5931 (N_5931,N_2549,N_773);
nand U5932 (N_5932,N_1634,N_2534);
nor U5933 (N_5933,N_39,N_2854);
nor U5934 (N_5934,N_372,N_1883);
or U5935 (N_5935,N_604,N_1719);
and U5936 (N_5936,N_2501,N_2618);
or U5937 (N_5937,N_1691,N_1558);
or U5938 (N_5938,N_2784,N_1474);
xnor U5939 (N_5939,N_1856,N_561);
xnor U5940 (N_5940,N_412,N_3099);
nor U5941 (N_5941,N_2518,N_731);
nor U5942 (N_5942,N_1724,N_1339);
xor U5943 (N_5943,N_125,N_2672);
nor U5944 (N_5944,N_64,N_1029);
or U5945 (N_5945,N_1943,N_1984);
xnor U5946 (N_5946,N_870,N_1710);
or U5947 (N_5947,N_1939,N_1224);
or U5948 (N_5948,N_1473,N_1941);
nand U5949 (N_5949,N_2726,N_575);
and U5950 (N_5950,N_3042,N_2805);
nor U5951 (N_5951,N_1826,N_424);
nor U5952 (N_5952,N_1218,N_1412);
xor U5953 (N_5953,N_1340,N_801);
nand U5954 (N_5954,N_1606,N_922);
nand U5955 (N_5955,N_452,N_1059);
xnor U5956 (N_5956,N_461,N_2588);
and U5957 (N_5957,N_2633,N_2655);
or U5958 (N_5958,N_1159,N_250);
nand U5959 (N_5959,N_159,N_1937);
and U5960 (N_5960,N_1098,N_3052);
or U5961 (N_5961,N_919,N_604);
and U5962 (N_5962,N_3084,N_761);
and U5963 (N_5963,N_1373,N_253);
xnor U5964 (N_5964,N_1905,N_1552);
xor U5965 (N_5965,N_1829,N_1253);
or U5966 (N_5966,N_284,N_2294);
or U5967 (N_5967,N_3111,N_211);
nor U5968 (N_5968,N_651,N_3105);
xnor U5969 (N_5969,N_39,N_654);
nor U5970 (N_5970,N_2207,N_92);
xnor U5971 (N_5971,N_324,N_2013);
or U5972 (N_5972,N_740,N_1150);
and U5973 (N_5973,N_725,N_1365);
and U5974 (N_5974,N_957,N_1887);
nand U5975 (N_5975,N_2553,N_2576);
xor U5976 (N_5976,N_1274,N_732);
nand U5977 (N_5977,N_1301,N_2772);
or U5978 (N_5978,N_2739,N_2526);
or U5979 (N_5979,N_855,N_391);
or U5980 (N_5980,N_189,N_1051);
and U5981 (N_5981,N_2559,N_2098);
nand U5982 (N_5982,N_1478,N_2087);
or U5983 (N_5983,N_1689,N_59);
nor U5984 (N_5984,N_1386,N_1367);
or U5985 (N_5985,N_1222,N_1245);
xor U5986 (N_5986,N_2278,N_2193);
nand U5987 (N_5987,N_509,N_63);
nor U5988 (N_5988,N_1854,N_1303);
nor U5989 (N_5989,N_2582,N_1650);
xor U5990 (N_5990,N_2114,N_181);
nor U5991 (N_5991,N_2747,N_18);
or U5992 (N_5992,N_1188,N_1798);
nand U5993 (N_5993,N_2933,N_2567);
and U5994 (N_5994,N_1949,N_366);
or U5995 (N_5995,N_2066,N_1739);
nand U5996 (N_5996,N_421,N_2601);
xor U5997 (N_5997,N_920,N_1102);
nor U5998 (N_5998,N_798,N_378);
and U5999 (N_5999,N_868,N_813);
or U6000 (N_6000,N_1442,N_533);
nor U6001 (N_6001,N_1709,N_1964);
nand U6002 (N_6002,N_3030,N_1868);
and U6003 (N_6003,N_2919,N_2645);
nand U6004 (N_6004,N_300,N_412);
nand U6005 (N_6005,N_546,N_2061);
nor U6006 (N_6006,N_610,N_1394);
nand U6007 (N_6007,N_39,N_428);
nand U6008 (N_6008,N_1660,N_2361);
and U6009 (N_6009,N_1275,N_2335);
and U6010 (N_6010,N_530,N_550);
or U6011 (N_6011,N_696,N_2605);
nand U6012 (N_6012,N_1415,N_481);
xnor U6013 (N_6013,N_1149,N_746);
nor U6014 (N_6014,N_274,N_2980);
nand U6015 (N_6015,N_864,N_3006);
or U6016 (N_6016,N_373,N_2824);
and U6017 (N_6017,N_2137,N_264);
nand U6018 (N_6018,N_1017,N_121);
or U6019 (N_6019,N_1235,N_1266);
or U6020 (N_6020,N_1564,N_1879);
xor U6021 (N_6021,N_2633,N_1950);
and U6022 (N_6022,N_2561,N_326);
nor U6023 (N_6023,N_2087,N_533);
and U6024 (N_6024,N_143,N_1853);
nor U6025 (N_6025,N_3055,N_1170);
xnor U6026 (N_6026,N_1688,N_1115);
and U6027 (N_6027,N_2899,N_2507);
xnor U6028 (N_6028,N_279,N_2436);
or U6029 (N_6029,N_840,N_2247);
nand U6030 (N_6030,N_1564,N_2967);
and U6031 (N_6031,N_2871,N_3069);
xnor U6032 (N_6032,N_1800,N_2971);
nor U6033 (N_6033,N_2467,N_2067);
or U6034 (N_6034,N_2411,N_1811);
xor U6035 (N_6035,N_48,N_949);
xnor U6036 (N_6036,N_355,N_2522);
or U6037 (N_6037,N_2302,N_2675);
nor U6038 (N_6038,N_967,N_2464);
or U6039 (N_6039,N_1867,N_841);
and U6040 (N_6040,N_2059,N_1287);
xnor U6041 (N_6041,N_1560,N_3095);
or U6042 (N_6042,N_48,N_2722);
or U6043 (N_6043,N_1557,N_1655);
nand U6044 (N_6044,N_203,N_187);
or U6045 (N_6045,N_868,N_2397);
nand U6046 (N_6046,N_627,N_1214);
xor U6047 (N_6047,N_2512,N_288);
xnor U6048 (N_6048,N_2288,N_335);
and U6049 (N_6049,N_2243,N_1285);
xor U6050 (N_6050,N_605,N_2826);
and U6051 (N_6051,N_2427,N_1838);
nor U6052 (N_6052,N_1416,N_2644);
nand U6053 (N_6053,N_134,N_2192);
nor U6054 (N_6054,N_26,N_732);
or U6055 (N_6055,N_1349,N_1389);
or U6056 (N_6056,N_816,N_1204);
nand U6057 (N_6057,N_2611,N_2729);
xor U6058 (N_6058,N_2580,N_406);
nand U6059 (N_6059,N_2917,N_1743);
nor U6060 (N_6060,N_1219,N_7);
and U6061 (N_6061,N_1284,N_2941);
nor U6062 (N_6062,N_1248,N_899);
nor U6063 (N_6063,N_1705,N_1323);
and U6064 (N_6064,N_2078,N_1469);
nor U6065 (N_6065,N_2759,N_1557);
and U6066 (N_6066,N_1838,N_2369);
and U6067 (N_6067,N_794,N_2771);
or U6068 (N_6068,N_524,N_520);
nand U6069 (N_6069,N_2417,N_1665);
or U6070 (N_6070,N_2170,N_3069);
and U6071 (N_6071,N_1643,N_2755);
nand U6072 (N_6072,N_785,N_1104);
and U6073 (N_6073,N_2366,N_1549);
and U6074 (N_6074,N_2351,N_3104);
and U6075 (N_6075,N_2735,N_1834);
or U6076 (N_6076,N_442,N_1950);
or U6077 (N_6077,N_1709,N_1812);
and U6078 (N_6078,N_491,N_2074);
xnor U6079 (N_6079,N_2887,N_2650);
xor U6080 (N_6080,N_2304,N_1976);
and U6081 (N_6081,N_191,N_110);
or U6082 (N_6082,N_1275,N_1451);
and U6083 (N_6083,N_1140,N_2829);
or U6084 (N_6084,N_1982,N_687);
nor U6085 (N_6085,N_1799,N_2540);
xor U6086 (N_6086,N_1859,N_2782);
nand U6087 (N_6087,N_2804,N_1284);
nand U6088 (N_6088,N_1949,N_504);
nand U6089 (N_6089,N_22,N_811);
xor U6090 (N_6090,N_1665,N_328);
nor U6091 (N_6091,N_2792,N_2507);
nor U6092 (N_6092,N_1636,N_338);
xor U6093 (N_6093,N_2466,N_3063);
or U6094 (N_6094,N_653,N_271);
nand U6095 (N_6095,N_132,N_1967);
nor U6096 (N_6096,N_1693,N_1188);
nand U6097 (N_6097,N_331,N_873);
xnor U6098 (N_6098,N_2645,N_2167);
nand U6099 (N_6099,N_491,N_1164);
and U6100 (N_6100,N_3041,N_2854);
and U6101 (N_6101,N_1259,N_2997);
or U6102 (N_6102,N_1708,N_73);
xor U6103 (N_6103,N_2605,N_289);
nor U6104 (N_6104,N_1538,N_2064);
and U6105 (N_6105,N_2517,N_2908);
nor U6106 (N_6106,N_1964,N_2094);
xor U6107 (N_6107,N_192,N_537);
nand U6108 (N_6108,N_2833,N_2036);
nor U6109 (N_6109,N_320,N_3102);
and U6110 (N_6110,N_2067,N_1161);
nor U6111 (N_6111,N_2293,N_1216);
xor U6112 (N_6112,N_2212,N_1463);
or U6113 (N_6113,N_347,N_1248);
nand U6114 (N_6114,N_3100,N_348);
nand U6115 (N_6115,N_1635,N_2172);
nand U6116 (N_6116,N_2335,N_754);
xnor U6117 (N_6117,N_366,N_666);
nor U6118 (N_6118,N_2699,N_2862);
and U6119 (N_6119,N_180,N_854);
nor U6120 (N_6120,N_2192,N_2740);
nor U6121 (N_6121,N_2558,N_2052);
nor U6122 (N_6122,N_1247,N_2380);
xor U6123 (N_6123,N_2544,N_2989);
xnor U6124 (N_6124,N_1716,N_1172);
and U6125 (N_6125,N_615,N_16);
or U6126 (N_6126,N_2829,N_2596);
and U6127 (N_6127,N_1545,N_1739);
nand U6128 (N_6128,N_1593,N_133);
nand U6129 (N_6129,N_2168,N_1792);
nor U6130 (N_6130,N_2473,N_298);
or U6131 (N_6131,N_2119,N_1869);
nor U6132 (N_6132,N_1346,N_1543);
xnor U6133 (N_6133,N_1624,N_1617);
and U6134 (N_6134,N_1836,N_2727);
nor U6135 (N_6135,N_328,N_1507);
nand U6136 (N_6136,N_116,N_2010);
and U6137 (N_6137,N_2171,N_283);
xor U6138 (N_6138,N_1038,N_268);
and U6139 (N_6139,N_779,N_377);
xnor U6140 (N_6140,N_1709,N_1451);
nand U6141 (N_6141,N_707,N_1190);
nor U6142 (N_6142,N_3093,N_612);
or U6143 (N_6143,N_1278,N_2117);
and U6144 (N_6144,N_2462,N_267);
xor U6145 (N_6145,N_200,N_1715);
nor U6146 (N_6146,N_2537,N_2911);
xnor U6147 (N_6147,N_310,N_1758);
xnor U6148 (N_6148,N_2361,N_30);
nand U6149 (N_6149,N_1247,N_1376);
nand U6150 (N_6150,N_909,N_1898);
nand U6151 (N_6151,N_1756,N_1063);
nor U6152 (N_6152,N_1285,N_485);
nor U6153 (N_6153,N_2962,N_86);
nor U6154 (N_6154,N_521,N_1331);
and U6155 (N_6155,N_122,N_2266);
or U6156 (N_6156,N_2028,N_11);
or U6157 (N_6157,N_1631,N_10);
xnor U6158 (N_6158,N_2806,N_2084);
xor U6159 (N_6159,N_278,N_2708);
xnor U6160 (N_6160,N_2305,N_498);
and U6161 (N_6161,N_2124,N_1403);
xor U6162 (N_6162,N_2944,N_2717);
or U6163 (N_6163,N_85,N_1262);
xor U6164 (N_6164,N_2786,N_1205);
nand U6165 (N_6165,N_2041,N_37);
nor U6166 (N_6166,N_252,N_1655);
nor U6167 (N_6167,N_1789,N_910);
nand U6168 (N_6168,N_1596,N_895);
or U6169 (N_6169,N_896,N_2438);
nand U6170 (N_6170,N_1760,N_2437);
and U6171 (N_6171,N_2787,N_2460);
or U6172 (N_6172,N_1468,N_195);
and U6173 (N_6173,N_1668,N_2204);
or U6174 (N_6174,N_802,N_2593);
nor U6175 (N_6175,N_711,N_3069);
nand U6176 (N_6176,N_320,N_1065);
nand U6177 (N_6177,N_2395,N_2518);
xor U6178 (N_6178,N_2170,N_744);
and U6179 (N_6179,N_3091,N_2007);
and U6180 (N_6180,N_1327,N_2443);
and U6181 (N_6181,N_2541,N_779);
or U6182 (N_6182,N_2503,N_1917);
or U6183 (N_6183,N_1902,N_2042);
or U6184 (N_6184,N_671,N_3023);
nand U6185 (N_6185,N_2337,N_2360);
xnor U6186 (N_6186,N_1264,N_498);
xor U6187 (N_6187,N_2185,N_1236);
xor U6188 (N_6188,N_1589,N_2338);
and U6189 (N_6189,N_694,N_736);
xor U6190 (N_6190,N_1900,N_394);
xnor U6191 (N_6191,N_193,N_1601);
and U6192 (N_6192,N_1954,N_852);
nor U6193 (N_6193,N_69,N_2246);
and U6194 (N_6194,N_3039,N_926);
nor U6195 (N_6195,N_932,N_1407);
nand U6196 (N_6196,N_687,N_801);
or U6197 (N_6197,N_226,N_236);
nand U6198 (N_6198,N_2985,N_1074);
and U6199 (N_6199,N_1001,N_2068);
nand U6200 (N_6200,N_1543,N_2836);
nor U6201 (N_6201,N_2263,N_1288);
and U6202 (N_6202,N_1301,N_1010);
nor U6203 (N_6203,N_1838,N_1970);
and U6204 (N_6204,N_2435,N_518);
nand U6205 (N_6205,N_1298,N_2752);
or U6206 (N_6206,N_760,N_2836);
or U6207 (N_6207,N_814,N_1397);
xor U6208 (N_6208,N_1079,N_1948);
and U6209 (N_6209,N_211,N_1736);
or U6210 (N_6210,N_1007,N_1911);
nand U6211 (N_6211,N_2947,N_2807);
nor U6212 (N_6212,N_2182,N_2239);
nand U6213 (N_6213,N_1322,N_2671);
xnor U6214 (N_6214,N_2410,N_866);
nand U6215 (N_6215,N_1894,N_1244);
or U6216 (N_6216,N_588,N_371);
or U6217 (N_6217,N_2898,N_1684);
nand U6218 (N_6218,N_1143,N_223);
xnor U6219 (N_6219,N_269,N_1474);
and U6220 (N_6220,N_801,N_1997);
xor U6221 (N_6221,N_2144,N_1190);
and U6222 (N_6222,N_2080,N_3119);
nand U6223 (N_6223,N_905,N_1468);
xnor U6224 (N_6224,N_1287,N_2428);
xor U6225 (N_6225,N_368,N_2361);
and U6226 (N_6226,N_2773,N_1744);
nor U6227 (N_6227,N_493,N_1793);
xnor U6228 (N_6228,N_3005,N_2432);
xor U6229 (N_6229,N_1256,N_5);
nor U6230 (N_6230,N_3005,N_3076);
xor U6231 (N_6231,N_2307,N_191);
nand U6232 (N_6232,N_2134,N_432);
nor U6233 (N_6233,N_1979,N_859);
and U6234 (N_6234,N_2733,N_2133);
nand U6235 (N_6235,N_729,N_680);
nand U6236 (N_6236,N_2363,N_2598);
nand U6237 (N_6237,N_1884,N_2883);
xnor U6238 (N_6238,N_262,N_3074);
xor U6239 (N_6239,N_1211,N_2066);
or U6240 (N_6240,N_3036,N_73);
nand U6241 (N_6241,N_2404,N_1101);
or U6242 (N_6242,N_1732,N_1464);
and U6243 (N_6243,N_2823,N_1461);
nor U6244 (N_6244,N_1351,N_1631);
or U6245 (N_6245,N_426,N_302);
nor U6246 (N_6246,N_3004,N_1971);
or U6247 (N_6247,N_861,N_76);
or U6248 (N_6248,N_2079,N_1975);
and U6249 (N_6249,N_1710,N_2497);
nor U6250 (N_6250,N_6229,N_4573);
nand U6251 (N_6251,N_4970,N_3619);
and U6252 (N_6252,N_4154,N_4467);
nor U6253 (N_6253,N_4853,N_5187);
xnor U6254 (N_6254,N_6101,N_4267);
nor U6255 (N_6255,N_3436,N_4872);
nor U6256 (N_6256,N_6136,N_3267);
nand U6257 (N_6257,N_3477,N_4379);
or U6258 (N_6258,N_4475,N_6019);
nand U6259 (N_6259,N_5133,N_5425);
or U6260 (N_6260,N_3419,N_4942);
and U6261 (N_6261,N_4733,N_3379);
nand U6262 (N_6262,N_6082,N_3246);
or U6263 (N_6263,N_3826,N_5209);
nor U6264 (N_6264,N_4882,N_5967);
nor U6265 (N_6265,N_3220,N_3644);
xor U6266 (N_6266,N_4114,N_5252);
and U6267 (N_6267,N_5927,N_6005);
nor U6268 (N_6268,N_5994,N_3707);
and U6269 (N_6269,N_6248,N_4779);
nand U6270 (N_6270,N_6026,N_3897);
nand U6271 (N_6271,N_6111,N_5582);
nand U6272 (N_6272,N_4259,N_5703);
and U6273 (N_6273,N_5917,N_3584);
and U6274 (N_6274,N_3806,N_5388);
and U6275 (N_6275,N_4108,N_5657);
nand U6276 (N_6276,N_3961,N_4222);
nand U6277 (N_6277,N_4753,N_4807);
nor U6278 (N_6278,N_3333,N_4959);
or U6279 (N_6279,N_6132,N_4177);
nor U6280 (N_6280,N_5830,N_3621);
and U6281 (N_6281,N_4889,N_5982);
or U6282 (N_6282,N_3256,N_6080);
nand U6283 (N_6283,N_4274,N_5717);
nor U6284 (N_6284,N_3132,N_5054);
nand U6285 (N_6285,N_5873,N_5642);
nand U6286 (N_6286,N_3561,N_4275);
nor U6287 (N_6287,N_5958,N_4436);
xor U6288 (N_6288,N_3176,N_3473);
xor U6289 (N_6289,N_5608,N_5814);
and U6290 (N_6290,N_4271,N_6023);
and U6291 (N_6291,N_5036,N_5130);
nand U6292 (N_6292,N_6104,N_5449);
nand U6293 (N_6293,N_5651,N_6220);
and U6294 (N_6294,N_3783,N_4496);
xor U6295 (N_6295,N_4273,N_3986);
or U6296 (N_6296,N_3348,N_3878);
nor U6297 (N_6297,N_4375,N_5047);
or U6298 (N_6298,N_4845,N_5355);
and U6299 (N_6299,N_5021,N_5874);
or U6300 (N_6300,N_6095,N_5416);
xor U6301 (N_6301,N_4893,N_4639);
xor U6302 (N_6302,N_5278,N_5617);
nand U6303 (N_6303,N_5628,N_5989);
and U6304 (N_6304,N_4456,N_4182);
and U6305 (N_6305,N_4416,N_5174);
and U6306 (N_6306,N_4127,N_4524);
nand U6307 (N_6307,N_5434,N_6207);
nand U6308 (N_6308,N_3574,N_3192);
nand U6309 (N_6309,N_5883,N_4877);
and U6310 (N_6310,N_5087,N_5141);
nor U6311 (N_6311,N_3834,N_3932);
nor U6312 (N_6312,N_4233,N_5094);
nor U6313 (N_6313,N_5501,N_4253);
and U6314 (N_6314,N_5713,N_5599);
xor U6315 (N_6315,N_5892,N_5399);
xnor U6316 (N_6316,N_3851,N_3388);
xor U6317 (N_6317,N_5264,N_5287);
xnor U6318 (N_6318,N_5083,N_4794);
nand U6319 (N_6319,N_3470,N_6179);
nand U6320 (N_6320,N_3260,N_4796);
and U6321 (N_6321,N_4378,N_5148);
xor U6322 (N_6322,N_5891,N_3965);
nand U6323 (N_6323,N_3616,N_4509);
and U6324 (N_6324,N_5186,N_3772);
and U6325 (N_6325,N_5670,N_4764);
nand U6326 (N_6326,N_3642,N_4937);
or U6327 (N_6327,N_4552,N_5333);
xnor U6328 (N_6328,N_4837,N_6202);
and U6329 (N_6329,N_3758,N_5732);
nand U6330 (N_6330,N_4815,N_3552);
and U6331 (N_6331,N_3865,N_3342);
and U6332 (N_6332,N_4590,N_4355);
and U6333 (N_6333,N_5941,N_3404);
nand U6334 (N_6334,N_5219,N_4068);
or U6335 (N_6335,N_4195,N_5409);
and U6336 (N_6336,N_5680,N_4351);
nor U6337 (N_6337,N_5869,N_4011);
or U6338 (N_6338,N_3815,N_5415);
and U6339 (N_6339,N_3202,N_4498);
or U6340 (N_6340,N_4157,N_4608);
and U6341 (N_6341,N_3341,N_5168);
nand U6342 (N_6342,N_3276,N_4574);
nor U6343 (N_6343,N_5284,N_3372);
nor U6344 (N_6344,N_4085,N_5022);
nand U6345 (N_6345,N_4503,N_5421);
and U6346 (N_6346,N_4756,N_5953);
or U6347 (N_6347,N_4159,N_6230);
nand U6348 (N_6348,N_4583,N_3273);
xor U6349 (N_6349,N_3374,N_3645);
and U6350 (N_6350,N_3723,N_5337);
nor U6351 (N_6351,N_6119,N_4001);
and U6352 (N_6352,N_3781,N_4603);
nor U6353 (N_6353,N_3973,N_3957);
xnor U6354 (N_6354,N_4985,N_5787);
nand U6355 (N_6355,N_4909,N_5178);
nand U6356 (N_6356,N_5442,N_5798);
nor U6357 (N_6357,N_3871,N_4582);
and U6358 (N_6358,N_4060,N_4399);
nor U6359 (N_6359,N_4955,N_4013);
xor U6360 (N_6360,N_5411,N_5214);
and U6361 (N_6361,N_5330,N_3441);
and U6362 (N_6362,N_4938,N_4530);
or U6363 (N_6363,N_4111,N_6043);
nor U6364 (N_6364,N_5556,N_4914);
xnor U6365 (N_6365,N_4719,N_3731);
nor U6366 (N_6366,N_6182,N_4268);
or U6367 (N_6367,N_5068,N_5108);
or U6368 (N_6368,N_3422,N_5461);
and U6369 (N_6369,N_5277,N_6091);
and U6370 (N_6370,N_5827,N_6145);
nand U6371 (N_6371,N_4553,N_3194);
and U6372 (N_6372,N_5946,N_4358);
nor U6373 (N_6373,N_3775,N_3369);
and U6374 (N_6374,N_3668,N_4960);
nor U6375 (N_6375,N_4606,N_3590);
and U6376 (N_6376,N_3523,N_4286);
and U6377 (N_6377,N_5822,N_3667);
nor U6378 (N_6378,N_4365,N_4096);
nand U6379 (N_6379,N_4414,N_5389);
xor U6380 (N_6380,N_5612,N_3627);
or U6381 (N_6381,N_3825,N_4121);
xnor U6382 (N_6382,N_5655,N_4324);
or U6383 (N_6383,N_3917,N_6064);
nand U6384 (N_6384,N_4663,N_4122);
nor U6385 (N_6385,N_5720,N_6083);
nand U6386 (N_6386,N_4835,N_4556);
nor U6387 (N_6387,N_4935,N_3448);
and U6388 (N_6388,N_3201,N_3634);
and U6389 (N_6389,N_3617,N_5926);
and U6390 (N_6390,N_5302,N_6167);
and U6391 (N_6391,N_3437,N_4287);
nand U6392 (N_6392,N_3160,N_6129);
and U6393 (N_6393,N_3340,N_4734);
and U6394 (N_6394,N_5244,N_3860);
nand U6395 (N_6395,N_5771,N_5895);
nor U6396 (N_6396,N_3290,N_5945);
xnor U6397 (N_6397,N_5886,N_3170);
xor U6398 (N_6398,N_3829,N_5129);
nand U6399 (N_6399,N_4843,N_6141);
nand U6400 (N_6400,N_6086,N_4161);
nor U6401 (N_6401,N_3647,N_5066);
xor U6402 (N_6402,N_4366,N_3942);
or U6403 (N_6403,N_4666,N_4097);
nand U6404 (N_6404,N_4501,N_6186);
nor U6405 (N_6405,N_4674,N_3258);
nor U6406 (N_6406,N_4795,N_4131);
nand U6407 (N_6407,N_6108,N_5654);
nand U6408 (N_6408,N_3182,N_4838);
and U6409 (N_6409,N_3925,N_3586);
xor U6410 (N_6410,N_3676,N_3930);
nand U6411 (N_6411,N_3518,N_3266);
or U6412 (N_6412,N_4851,N_3423);
nor U6413 (N_6413,N_5024,N_5254);
and U6414 (N_6414,N_4381,N_5290);
xnor U6415 (N_6415,N_6049,N_5076);
or U6416 (N_6416,N_3835,N_4419);
nand U6417 (N_6417,N_5731,N_3728);
nor U6418 (N_6418,N_4479,N_5759);
and U6419 (N_6419,N_6185,N_5908);
nand U6420 (N_6420,N_4057,N_5593);
or U6421 (N_6421,N_6050,N_5709);
and U6422 (N_6422,N_4242,N_5301);
and U6423 (N_6423,N_5041,N_6213);
nand U6424 (N_6424,N_3317,N_5951);
nand U6425 (N_6425,N_4304,N_5331);
nor U6426 (N_6426,N_5548,N_5096);
and U6427 (N_6427,N_6174,N_3820);
or U6428 (N_6428,N_4842,N_3777);
xnor U6429 (N_6429,N_6094,N_5524);
or U6430 (N_6430,N_3883,N_3169);
nor U6431 (N_6431,N_3785,N_5766);
or U6432 (N_6432,N_3329,N_3721);
nor U6433 (N_6433,N_3507,N_4782);
and U6434 (N_6434,N_3275,N_5398);
nor U6435 (N_6435,N_4083,N_3531);
and U6436 (N_6436,N_3370,N_4326);
and U6437 (N_6437,N_3792,N_5812);
xor U6438 (N_6438,N_6201,N_3277);
nor U6439 (N_6439,N_4035,N_4732);
or U6440 (N_6440,N_3771,N_4124);
nor U6441 (N_6441,N_4071,N_5183);
nor U6442 (N_6442,N_6062,N_5327);
xnor U6443 (N_6443,N_6238,N_6243);
nand U6444 (N_6444,N_4393,N_5393);
nor U6445 (N_6445,N_5833,N_4137);
or U6446 (N_6446,N_5013,N_5966);
and U6447 (N_6447,N_4327,N_4526);
nand U6448 (N_6448,N_4095,N_3378);
nand U6449 (N_6449,N_3803,N_6240);
and U6450 (N_6450,N_3732,N_4291);
and U6451 (N_6451,N_5577,N_4610);
and U6452 (N_6452,N_5899,N_5243);
xnor U6453 (N_6453,N_4979,N_5255);
or U6454 (N_6454,N_3940,N_3375);
xor U6455 (N_6455,N_5610,N_4962);
xor U6456 (N_6456,N_3754,N_5227);
xnor U6457 (N_6457,N_4369,N_5954);
or U6458 (N_6458,N_5669,N_4925);
or U6459 (N_6459,N_4688,N_5746);
nor U6460 (N_6460,N_3278,N_3136);
or U6461 (N_6461,N_4107,N_5520);
xor U6462 (N_6462,N_4755,N_4003);
and U6463 (N_6463,N_3671,N_3532);
nor U6464 (N_6464,N_4638,N_5157);
and U6465 (N_6465,N_5180,N_4328);
xor U6466 (N_6466,N_6098,N_3666);
and U6467 (N_6467,N_6002,N_5602);
and U6468 (N_6468,N_5872,N_4039);
or U6469 (N_6469,N_4309,N_3601);
nor U6470 (N_6470,N_4312,N_4836);
or U6471 (N_6471,N_3332,N_3528);
and U6472 (N_6472,N_4940,N_5781);
nor U6473 (N_6473,N_5795,N_4828);
xnor U6474 (N_6474,N_5631,N_5395);
or U6475 (N_6475,N_5205,N_4264);
nand U6476 (N_6476,N_5619,N_4272);
or U6477 (N_6477,N_5643,N_4991);
or U6478 (N_6478,N_5344,N_6116);
and U6479 (N_6479,N_3135,N_3742);
or U6480 (N_6480,N_4420,N_5860);
nand U6481 (N_6481,N_3364,N_3580);
nor U6482 (N_6482,N_4063,N_4873);
and U6483 (N_6483,N_4849,N_3499);
nand U6484 (N_6484,N_5796,N_3630);
nor U6485 (N_6485,N_4857,N_5320);
nor U6486 (N_6486,N_3365,N_5810);
or U6487 (N_6487,N_6096,N_4693);
xnor U6488 (N_6488,N_6017,N_3813);
xnor U6489 (N_6489,N_5073,N_5868);
xnor U6490 (N_6490,N_4100,N_3226);
and U6491 (N_6491,N_3740,N_3356);
or U6492 (N_6492,N_5028,N_5229);
nor U6493 (N_6493,N_4504,N_4440);
and U6494 (N_6494,N_3782,N_4752);
nor U6495 (N_6495,N_5218,N_4981);
nor U6496 (N_6496,N_3500,N_4657);
nand U6497 (N_6497,N_3347,N_3431);
and U6498 (N_6498,N_3884,N_5630);
or U6499 (N_6499,N_5295,N_5764);
and U6500 (N_6500,N_5986,N_4581);
nand U6501 (N_6501,N_5910,N_4319);
xor U6502 (N_6502,N_3307,N_5852);
or U6503 (N_6503,N_3377,N_3670);
and U6504 (N_6504,N_5894,N_4076);
nor U6505 (N_6505,N_3636,N_3309);
nand U6506 (N_6506,N_3190,N_3455);
nand U6507 (N_6507,N_3748,N_6100);
xor U6508 (N_6508,N_5907,N_4196);
and U6509 (N_6509,N_5478,N_3325);
nor U6510 (N_6510,N_5088,N_5674);
nor U6511 (N_6511,N_5864,N_6033);
or U6512 (N_6512,N_5134,N_4106);
nand U6513 (N_6513,N_4531,N_5314);
nand U6514 (N_6514,N_6221,N_3506);
or U6515 (N_6515,N_5271,N_6169);
xor U6516 (N_6516,N_3784,N_6006);
and U6517 (N_6517,N_3400,N_4026);
xnor U6518 (N_6518,N_4586,N_4936);
nor U6519 (N_6519,N_3461,N_5267);
nand U6520 (N_6520,N_4947,N_4762);
nand U6521 (N_6521,N_4249,N_3952);
nand U6522 (N_6522,N_6142,N_5974);
and U6523 (N_6523,N_4469,N_3412);
xnor U6524 (N_6524,N_6113,N_3494);
xnor U6525 (N_6525,N_3409,N_3217);
nand U6526 (N_6526,N_5127,N_4950);
or U6527 (N_6527,N_3738,N_3692);
or U6528 (N_6528,N_5361,N_3765);
and U6529 (N_6529,N_3373,N_3827);
or U6530 (N_6530,N_4700,N_3950);
nand U6531 (N_6531,N_6196,N_6237);
nand U6532 (N_6532,N_5420,N_3538);
xnor U6533 (N_6533,N_6135,N_5505);
nor U6534 (N_6534,N_4874,N_4783);
nand U6535 (N_6535,N_3969,N_6194);
and U6536 (N_6536,N_4450,N_6107);
xor U6537 (N_6537,N_3664,N_4775);
nor U6538 (N_6538,N_4799,N_3193);
or U6539 (N_6539,N_5211,N_4120);
nand U6540 (N_6540,N_5265,N_5740);
nand U6541 (N_6541,N_5542,N_5905);
nand U6542 (N_6542,N_4330,N_3480);
or U6543 (N_6543,N_4726,N_5242);
xor U6544 (N_6544,N_3222,N_3126);
xor U6545 (N_6545,N_5800,N_4622);
nand U6546 (N_6546,N_3594,N_3891);
and U6547 (N_6547,N_4356,N_5235);
nor U6548 (N_6548,N_4855,N_3174);
and U6549 (N_6549,N_5513,N_3401);
nor U6550 (N_6550,N_4844,N_4992);
nand U6551 (N_6551,N_4104,N_5568);
nor U6552 (N_6552,N_6037,N_5773);
and U6553 (N_6553,N_5611,N_6071);
xnor U6554 (N_6554,N_5203,N_4594);
nor U6555 (N_6555,N_3312,N_4896);
and U6556 (N_6556,N_4146,N_5431);
nand U6557 (N_6557,N_6151,N_6247);
nand U6558 (N_6558,N_3212,N_3888);
and U6559 (N_6559,N_3872,N_5526);
and U6560 (N_6560,N_5115,N_5418);
xor U6561 (N_6561,N_4801,N_6159);
or U6562 (N_6562,N_3467,N_4335);
xnor U6563 (N_6563,N_5373,N_3505);
xor U6564 (N_6564,N_4833,N_5805);
nor U6565 (N_6565,N_4141,N_4653);
nor U6566 (N_6566,N_6146,N_4256);
and U6567 (N_6567,N_4579,N_4702);
xor U6568 (N_6568,N_5516,N_4648);
or U6569 (N_6569,N_3191,N_3289);
nor U6570 (N_6570,N_3287,N_5444);
xnor U6571 (N_6571,N_5898,N_3795);
xnor U6572 (N_6572,N_4099,N_3900);
nand U6573 (N_6573,N_5109,N_5098);
and U6574 (N_6574,N_3614,N_5164);
nand U6575 (N_6575,N_3944,N_5086);
xnor U6576 (N_6576,N_4978,N_3776);
or U6577 (N_6577,N_5483,N_3894);
or U6578 (N_6578,N_3682,N_4205);
and U6579 (N_6579,N_4332,N_3547);
nand U6580 (N_6580,N_3301,N_6242);
and U6581 (N_6581,N_5341,N_5467);
nand U6582 (N_6582,N_5722,N_5554);
xor U6583 (N_6583,N_4892,N_5126);
and U6584 (N_6584,N_5138,N_4072);
nand U6585 (N_6585,N_4213,N_5043);
and U6586 (N_6586,N_6003,N_3546);
xnor U6587 (N_6587,N_3343,N_4093);
nand U6588 (N_6588,N_5595,N_6092);
and U6589 (N_6589,N_5909,N_5896);
or U6590 (N_6590,N_5716,N_3430);
or U6591 (N_6591,N_5633,N_3207);
nor U6592 (N_6592,N_5867,N_3241);
and U6593 (N_6593,N_4245,N_3306);
xnor U6594 (N_6594,N_3632,N_4187);
nor U6595 (N_6595,N_3922,N_4262);
nand U6596 (N_6596,N_4313,N_6183);
nor U6597 (N_6597,N_3846,N_5832);
and U6598 (N_6598,N_4193,N_3519);
xor U6599 (N_6599,N_5775,N_4422);
nor U6600 (N_6600,N_5348,N_5075);
xnor U6601 (N_6601,N_3658,N_4034);
xor U6602 (N_6602,N_5008,N_4966);
xnor U6603 (N_6603,N_5499,N_4151);
xnor U6604 (N_6604,N_4596,N_4727);
xor U6605 (N_6605,N_3495,N_5437);
xnor U6606 (N_6606,N_5564,N_4015);
nand U6607 (N_6607,N_4018,N_4510);
nand U6608 (N_6608,N_5809,N_4269);
or U6609 (N_6609,N_4659,N_3209);
and U6610 (N_6610,N_4441,N_4317);
nor U6611 (N_6611,N_3701,N_4618);
nor U6612 (N_6612,N_4051,N_5544);
nand U6613 (N_6613,N_5646,N_4410);
or U6614 (N_6614,N_4155,N_3439);
xor U6615 (N_6615,N_4718,N_6189);
nor U6616 (N_6616,N_5045,N_5104);
xor U6617 (N_6617,N_5707,N_5197);
nand U6618 (N_6618,N_4261,N_5149);
or U6619 (N_6619,N_3315,N_5534);
xor U6620 (N_6620,N_3533,N_3768);
nor U6621 (N_6621,N_3727,N_5458);
xnor U6622 (N_6622,N_4944,N_5491);
and U6623 (N_6623,N_5515,N_5057);
xor U6624 (N_6624,N_5377,N_3735);
nor U6625 (N_6625,N_4518,N_3992);
and U6626 (N_6626,N_3432,N_4406);
and U6627 (N_6627,N_4200,N_3831);
nor U6628 (N_6628,N_5317,N_4777);
and U6629 (N_6629,N_4360,N_4706);
and U6630 (N_6630,N_6227,N_4160);
xor U6631 (N_6631,N_5182,N_5792);
or U6632 (N_6632,N_5189,N_6231);
xor U6633 (N_6633,N_4126,N_5807);
nand U6634 (N_6634,N_4325,N_3296);
nor U6635 (N_6635,N_5351,N_5804);
or U6636 (N_6636,N_3935,N_3770);
nand U6637 (N_6637,N_3255,N_3767);
nand U6638 (N_6638,N_4624,N_5741);
nor U6639 (N_6639,N_3261,N_5500);
nand U6640 (N_6640,N_4294,N_4398);
nor U6641 (N_6641,N_5837,N_4387);
nor U6642 (N_6642,N_3639,N_5546);
or U6643 (N_6643,N_5046,N_5998);
and U6644 (N_6644,N_5503,N_4643);
nor U6645 (N_6645,N_4507,N_4823);
xor U6646 (N_6646,N_6035,N_5755);
and U6647 (N_6647,N_4280,N_4725);
xnor U6648 (N_6648,N_5213,N_3462);
and U6649 (N_6649,N_6154,N_5885);
or U6650 (N_6650,N_4152,N_5349);
nor U6651 (N_6651,N_5545,N_5492);
xnor U6652 (N_6652,N_4683,N_4293);
or U6653 (N_6653,N_4241,N_5992);
nor U6654 (N_6654,N_3737,N_3887);
and U6655 (N_6655,N_3648,N_5845);
nand U6656 (N_6656,N_3691,N_4982);
xor U6657 (N_6657,N_4595,N_3137);
nand U6658 (N_6658,N_5594,N_5884);
nor U6659 (N_6659,N_3128,N_4623);
or U6660 (N_6660,N_3408,N_5266);
or U6661 (N_6661,N_5813,N_6034);
xor U6662 (N_6662,N_4668,N_5914);
or U6663 (N_6663,N_3200,N_5676);
nand U6664 (N_6664,N_5817,N_5407);
nor U6665 (N_6665,N_5865,N_6022);
nor U6666 (N_6666,N_4932,N_4780);
and U6667 (N_6667,N_6015,N_3763);
nand U6668 (N_6668,N_5123,N_5258);
or U6669 (N_6669,N_6204,N_3282);
xor U6670 (N_6670,N_4729,N_6168);
or U6671 (N_6671,N_4132,N_4631);
xnor U6672 (N_6672,N_5942,N_4158);
nor U6673 (N_6673,N_5690,N_5721);
and U6674 (N_6674,N_3857,N_3281);
and U6675 (N_6675,N_3357,N_4862);
nand U6676 (N_6676,N_4118,N_3328);
nand U6677 (N_6677,N_3974,N_3310);
and U6678 (N_6678,N_4773,N_5701);
nor U6679 (N_6679,N_5962,N_3206);
nand U6680 (N_6680,N_3213,N_5163);
xor U6681 (N_6681,N_4956,N_4390);
or U6682 (N_6682,N_4585,N_4870);
nand U6683 (N_6683,N_4539,N_4993);
nand U6684 (N_6684,N_5818,N_4227);
xor U6685 (N_6685,N_5949,N_4066);
and U6686 (N_6686,N_3869,N_5750);
or U6687 (N_6687,N_4407,N_4776);
nand U6688 (N_6688,N_4391,N_5025);
xor U6689 (N_6689,N_3990,N_5626);
nor U6690 (N_6690,N_3384,N_5576);
nand U6691 (N_6691,N_3945,N_5144);
xnor U6692 (N_6692,N_4964,N_6027);
or U6693 (N_6693,N_6193,N_5777);
or U6694 (N_6694,N_5575,N_5705);
nor U6695 (N_6695,N_3355,N_3868);
nand U6696 (N_6696,N_4029,N_4611);
or U6697 (N_6697,N_4995,N_6233);
and U6698 (N_6698,N_5359,N_4565);
or U6699 (N_6699,N_5973,N_5502);
nor U6700 (N_6700,N_5439,N_5450);
xor U6701 (N_6701,N_4329,N_3510);
or U6702 (N_6702,N_5313,N_6122);
nand U6703 (N_6703,N_5085,N_3566);
or U6704 (N_6704,N_3149,N_4785);
nor U6705 (N_6705,N_3716,N_5596);
xor U6706 (N_6706,N_5736,N_4299);
or U6707 (N_6707,N_3497,N_3243);
nor U6708 (N_6708,N_5932,N_3620);
xor U6709 (N_6709,N_3535,N_5930);
xor U6710 (N_6710,N_4921,N_3219);
or U6711 (N_6711,N_4605,N_4528);
nand U6712 (N_6712,N_3605,N_3841);
nor U6713 (N_6713,N_5535,N_3956);
nand U6714 (N_6714,N_3840,N_3705);
or U6715 (N_6715,N_3324,N_5256);
and U6716 (N_6716,N_5991,N_3215);
xnor U6717 (N_6717,N_4832,N_4901);
nor U6718 (N_6718,N_5304,N_3877);
and U6719 (N_6719,N_5152,N_4554);
nand U6720 (N_6720,N_5143,N_3819);
nor U6721 (N_6721,N_4640,N_5474);
or U6722 (N_6722,N_4879,N_4613);
or U6723 (N_6723,N_3483,N_3873);
xor U6724 (N_6724,N_6025,N_4142);
and U6725 (N_6725,N_5275,N_4404);
xor U6726 (N_6726,N_6018,N_6188);
nand U6727 (N_6727,N_4426,N_4850);
or U6728 (N_6728,N_4316,N_5708);
xor U6729 (N_6729,N_4385,N_5414);
nand U6730 (N_6730,N_5291,N_4677);
nand U6731 (N_6731,N_3830,N_3623);
nand U6732 (N_6732,N_3934,N_5857);
and U6733 (N_6733,N_5298,N_3165);
and U6734 (N_6734,N_5090,N_5325);
xor U6735 (N_6735,N_4566,N_5072);
xor U6736 (N_6736,N_3527,N_4711);
or U6737 (N_6737,N_4545,N_5059);
xnor U6738 (N_6738,N_3263,N_5100);
nand U6739 (N_6739,N_3139,N_3903);
or U6740 (N_6740,N_5489,N_5011);
or U6741 (N_6741,N_3663,N_5462);
or U6742 (N_6742,N_3453,N_3832);
or U6743 (N_6743,N_5185,N_3780);
or U6744 (N_6744,N_5959,N_4564);
and U6745 (N_6745,N_3643,N_3850);
nand U6746 (N_6746,N_5099,N_4408);
xor U6747 (N_6747,N_5558,N_3380);
and U6748 (N_6748,N_5627,N_6051);
and U6749 (N_6749,N_3351,N_3606);
nor U6750 (N_6750,N_5841,N_4172);
and U6751 (N_6751,N_5172,N_3560);
nor U6752 (N_6752,N_4401,N_3635);
xor U6753 (N_6753,N_5221,N_4344);
nand U6754 (N_6754,N_4447,N_4339);
nand U6755 (N_6755,N_5368,N_4522);
xnor U6756 (N_6756,N_5251,N_3674);
or U6757 (N_6757,N_3793,N_3802);
or U6758 (N_6758,N_4221,N_4119);
and U6759 (N_6759,N_5641,N_3700);
xnor U6760 (N_6760,N_5177,N_3876);
nor U6761 (N_6761,N_4601,N_3719);
or U6762 (N_6762,N_4170,N_5062);
or U6763 (N_6763,N_4054,N_3913);
and U6764 (N_6764,N_4588,N_4954);
nand U6765 (N_6765,N_3294,N_4642);
xor U6766 (N_6766,N_6052,N_5681);
nand U6767 (N_6767,N_4786,N_5020);
xnor U6768 (N_6768,N_5581,N_4207);
nand U6769 (N_6769,N_4023,N_5481);
xor U6770 (N_6770,N_5385,N_3694);
xnor U6771 (N_6771,N_4058,N_3336);
nor U6772 (N_6772,N_3144,N_5523);
nand U6773 (N_6773,N_3382,N_4252);
xor U6774 (N_6774,N_5983,N_5977);
or U6775 (N_6775,N_3427,N_3853);
or U6776 (N_6776,N_5531,N_4499);
xnor U6777 (N_6777,N_4856,N_3308);
and U6778 (N_6778,N_4434,N_3446);
nor U6779 (N_6779,N_5122,N_3487);
nor U6780 (N_6780,N_3807,N_3843);
xnor U6781 (N_6781,N_5735,N_3173);
xnor U6782 (N_6782,N_5223,N_5055);
nor U6783 (N_6783,N_4968,N_3303);
or U6784 (N_6784,N_4140,N_5639);
nand U6785 (N_6785,N_3743,N_4690);
xor U6786 (N_6786,N_4548,N_4235);
nor U6787 (N_6787,N_3757,N_5934);
or U6788 (N_6788,N_5679,N_3710);
nor U6789 (N_6789,N_3762,N_4681);
nor U6790 (N_6790,N_5270,N_3895);
or U6791 (N_6791,N_4165,N_5620);
nor U6792 (N_6792,N_5370,N_4423);
nor U6793 (N_6793,N_5706,N_3822);
and U6794 (N_6794,N_5200,N_4383);
and U6795 (N_6795,N_3858,N_3541);
nor U6796 (N_6796,N_3141,N_5406);
xnor U6797 (N_6797,N_3958,N_4276);
and U6798 (N_6798,N_4922,N_4990);
or U6799 (N_6799,N_4377,N_6236);
xnor U6800 (N_6800,N_4634,N_5063);
xor U6801 (N_6801,N_3695,N_3394);
nand U6802 (N_6802,N_5527,N_4766);
and U6803 (N_6803,N_4130,N_5944);
nand U6804 (N_6804,N_3955,N_4951);
and U6805 (N_6805,N_5009,N_4948);
and U6806 (N_6806,N_4745,N_5756);
and U6807 (N_6807,N_4770,N_4115);
xnor U6808 (N_6808,N_6187,N_5533);
nor U6809 (N_6809,N_3808,N_6197);
nor U6810 (N_6810,N_5472,N_5035);
or U6811 (N_6811,N_6103,N_4769);
and U6812 (N_6812,N_3204,N_4074);
or U6813 (N_6813,N_5723,N_3398);
or U6814 (N_6814,N_4334,N_4396);
xor U6815 (N_6815,N_5195,N_5039);
nand U6816 (N_6816,N_4816,N_3970);
and U6817 (N_6817,N_3501,N_5136);
or U6818 (N_6818,N_6138,N_3524);
nor U6819 (N_6819,N_5618,N_4980);
xnor U6820 (N_6820,N_6115,N_3300);
nand U6821 (N_6821,N_4445,N_4656);
xnor U6822 (N_6822,N_3486,N_4350);
and U6823 (N_6823,N_3870,N_3655);
nor U6824 (N_6824,N_4513,N_3714);
nor U6825 (N_6825,N_5065,N_6061);
and U6826 (N_6826,N_5215,N_5422);
nor U6827 (N_6827,N_5662,N_3545);
nand U6828 (N_6828,N_4136,N_3690);
nand U6829 (N_6829,N_3800,N_3633);
and U6830 (N_6830,N_4989,N_3657);
nor U6831 (N_6831,N_4215,N_6065);
and U6832 (N_6832,N_5560,N_3319);
and U6833 (N_6833,N_6013,N_3572);
or U6834 (N_6834,N_5604,N_4219);
and U6835 (N_6835,N_4452,N_4340);
and U6836 (N_6836,N_5352,N_5786);
xor U6837 (N_6837,N_4535,N_4216);
nand U6838 (N_6838,N_3138,N_3228);
and U6839 (N_6839,N_4675,N_4139);
nor U6840 (N_6840,N_3752,N_3556);
nand U6841 (N_6841,N_4202,N_4813);
nand U6842 (N_6842,N_5002,N_5176);
nor U6843 (N_6843,N_5192,N_3517);
and U6844 (N_6844,N_5820,N_4555);
nor U6845 (N_6845,N_4515,N_4028);
nand U6846 (N_6846,N_4612,N_5345);
xnor U6847 (N_6847,N_3515,N_5372);
nand U6848 (N_6848,N_4863,N_4492);
or U6849 (N_6849,N_3167,N_5609);
nor U6850 (N_6850,N_3428,N_4143);
or U6851 (N_6851,N_3334,N_3660);
and U6852 (N_6852,N_5184,N_5774);
nand U6853 (N_6853,N_4374,N_4930);
or U6854 (N_6854,N_5167,N_3989);
or U6855 (N_6855,N_5485,N_4860);
xor U6856 (N_6856,N_5217,N_5844);
or U6857 (N_6857,N_3525,N_5162);
and U6858 (N_6858,N_3218,N_3665);
or U6859 (N_6859,N_4285,N_5603);
xor U6860 (N_6860,N_5836,N_3371);
or U6861 (N_6861,N_3361,N_4191);
nor U6862 (N_6862,N_3656,N_6024);
or U6863 (N_6863,N_4461,N_5871);
and U6864 (N_6864,N_4720,N_3549);
nor U6865 (N_6865,N_6218,N_5487);
xor U6866 (N_6866,N_3321,N_4288);
xor U6867 (N_6867,N_5715,N_6149);
nor U6868 (N_6868,N_5950,N_3235);
nand U6869 (N_6869,N_5069,N_6158);
and U6870 (N_6870,N_4997,N_3749);
xor U6871 (N_6871,N_5965,N_5346);
xor U6872 (N_6872,N_3753,N_4485);
xnor U6873 (N_6873,N_3905,N_5403);
nor U6874 (N_6874,N_3987,N_4210);
nand U6875 (N_6875,N_3567,N_5433);
xnor U6876 (N_6876,N_4232,N_4793);
xor U6877 (N_6877,N_4895,N_4791);
xnor U6878 (N_6878,N_5296,N_6172);
nand U6879 (N_6879,N_3330,N_5234);
or U6880 (N_6880,N_4084,N_5607);
xor U6881 (N_6881,N_3352,N_5095);
xnor U6882 (N_6882,N_4376,N_4866);
or U6883 (N_6883,N_5606,N_3286);
nor U6884 (N_6884,N_5634,N_3504);
or U6885 (N_6885,N_3946,N_5691);
and U6886 (N_6886,N_5017,N_4254);
xnor U6887 (N_6887,N_4800,N_3578);
nand U6888 (N_6888,N_3972,N_4091);
nor U6889 (N_6889,N_3976,N_3713);
xor U6890 (N_6890,N_5007,N_4435);
nor U6891 (N_6891,N_5825,N_4112);
nor U6892 (N_6892,N_4025,N_4443);
nand U6893 (N_6893,N_6073,N_3514);
xor U6894 (N_6894,N_4894,N_5142);
and U6895 (N_6895,N_5463,N_3562);
or U6896 (N_6896,N_5644,N_5369);
nand U6897 (N_6897,N_3415,N_4031);
nand U6898 (N_6898,N_4881,N_4069);
or U6899 (N_6899,N_5347,N_5240);
or U6900 (N_6900,N_4840,N_4967);
nor U6901 (N_6901,N_4803,N_5537);
nand U6902 (N_6902,N_6088,N_5719);
xor U6903 (N_6903,N_3725,N_4053);
xor U6904 (N_6904,N_5412,N_3469);
or U6905 (N_6905,N_5358,N_4508);
xnor U6906 (N_6906,N_5931,N_3910);
nand U6907 (N_6907,N_3456,N_5511);
xor U6908 (N_6908,N_5309,N_4713);
and U6909 (N_6909,N_3444,N_3602);
and U6910 (N_6910,N_5323,N_5725);
and U6911 (N_6911,N_3508,N_4953);
and U6912 (N_6912,N_3387,N_6045);
nand U6913 (N_6913,N_3610,N_5078);
or U6914 (N_6914,N_3845,N_5216);
and U6915 (N_6915,N_3180,N_3573);
nor U6916 (N_6916,N_4203,N_5689);
nand U6917 (N_6917,N_5056,N_3733);
or U6918 (N_6918,N_4250,N_6085);
nor U6919 (N_6919,N_5307,N_5044);
xor U6920 (N_6920,N_5292,N_3471);
and U6921 (N_6921,N_6016,N_5424);
or U6922 (N_6922,N_3199,N_3530);
nand U6923 (N_6923,N_3810,N_3151);
nand U6924 (N_6924,N_6001,N_5664);
or U6925 (N_6925,N_4336,N_5739);
nand U6926 (N_6926,N_3833,N_4739);
and U6927 (N_6927,N_4476,N_4346);
nand U6928 (N_6928,N_4297,N_5519);
or U6929 (N_6929,N_4497,N_5887);
or U6930 (N_6930,N_5427,N_5536);
nor U6931 (N_6931,N_5498,N_4214);
and U6932 (N_6932,N_4022,N_3592);
nand U6933 (N_6933,N_6114,N_5111);
or U6934 (N_6934,N_5324,N_4303);
or U6935 (N_6935,N_4045,N_4050);
or U6936 (N_6936,N_3434,N_3177);
nand U6937 (N_6937,N_3251,N_3809);
nor U6938 (N_6938,N_4077,N_3451);
or U6939 (N_6939,N_3607,N_4502);
and U6940 (N_6940,N_4934,N_4212);
nor U6941 (N_6941,N_5181,N_3236);
nand U6942 (N_6942,N_4987,N_5000);
or U6943 (N_6943,N_3280,N_3337);
xnor U6944 (N_6944,N_5367,N_4144);
nand U6945 (N_6945,N_3718,N_4321);
nand U6946 (N_6946,N_4352,N_4712);
nor U6947 (N_6947,N_5566,N_4048);
nand U6948 (N_6948,N_5394,N_4279);
or U6949 (N_6949,N_4103,N_4710);
nor U6950 (N_6950,N_3411,N_6177);
xnor U6951 (N_6951,N_4004,N_4886);
nor U6952 (N_6952,N_4629,N_5652);
nand U6953 (N_6953,N_4692,N_5808);
or U6954 (N_6954,N_4183,N_4699);
nand U6955 (N_6955,N_4614,N_4821);
or U6956 (N_6956,N_5935,N_5471);
xor U6957 (N_6957,N_4958,N_3159);
xnor U6958 (N_6958,N_5589,N_6044);
or U6959 (N_6959,N_4709,N_5636);
and U6960 (N_6960,N_3252,N_5274);
nor U6961 (N_6961,N_5879,N_3818);
or U6962 (N_6962,N_5473,N_3326);
xnor U6963 (N_6963,N_3929,N_3238);
nand U6964 (N_6964,N_3178,N_4283);
nand U6965 (N_6965,N_5699,N_5661);
xor U6966 (N_6966,N_6148,N_4086);
nor U6967 (N_6967,N_5006,N_4024);
and U6968 (N_6968,N_5048,N_6214);
nor U6969 (N_6969,N_3396,N_5312);
or U6970 (N_6970,N_5089,N_5768);
xor U6971 (N_6971,N_4721,N_5952);
xnor U6972 (N_6972,N_5482,N_5033);
xor U6973 (N_6973,N_5540,N_4455);
nor U6974 (N_6974,N_5955,N_3896);
xnor U6975 (N_6975,N_5030,N_4523);
and U6976 (N_6976,N_4741,N_5451);
nand U6977 (N_6977,N_5316,N_4749);
and U6978 (N_6978,N_4282,N_5976);
or U6979 (N_6979,N_5190,N_4189);
nor U6980 (N_6980,N_3168,N_3147);
nand U6981 (N_6981,N_6042,N_4201);
or U6982 (N_6982,N_5169,N_3516);
nor U6983 (N_6983,N_6060,N_4661);
nor U6984 (N_6984,N_4912,N_4395);
nand U6985 (N_6985,N_4305,N_3997);
nor U6986 (N_6986,N_4148,N_6057);
or U6987 (N_6987,N_4728,N_5012);
xnor U6988 (N_6988,N_5097,N_3397);
or U6989 (N_6989,N_4694,N_5876);
and U6990 (N_6990,N_4430,N_5118);
nand U6991 (N_6991,N_5999,N_4010);
nor U6992 (N_6992,N_5790,N_4149);
xnor U6993 (N_6993,N_5175,N_3916);
or U6994 (N_6994,N_5729,N_5226);
xnor U6995 (N_6995,N_6081,N_5261);
xor U6996 (N_6996,N_5692,N_6077);
and U6997 (N_6997,N_3175,N_5635);
nor U6998 (N_6998,N_5925,N_5245);
nor U6999 (N_6999,N_3271,N_5281);
and U7000 (N_7000,N_4134,N_6031);
and U7001 (N_7001,N_4907,N_6139);
xnor U7002 (N_7002,N_3588,N_5529);
xnor U7003 (N_7003,N_5788,N_5114);
and U7004 (N_7004,N_3225,N_3669);
and U7005 (N_7005,N_3249,N_5854);
or U7006 (N_7006,N_5052,N_3975);
nor U7007 (N_7007,N_4342,N_5426);
nand U7008 (N_7008,N_4705,N_5077);
and U7009 (N_7009,N_5615,N_4617);
and U7010 (N_7010,N_5658,N_5423);
and U7011 (N_7011,N_3927,N_3653);
or U7012 (N_7012,N_3652,N_5921);
nand U7013 (N_7013,N_5851,N_3570);
xnor U7014 (N_7014,N_4761,N_4179);
nor U7015 (N_7015,N_4314,N_5125);
nor U7016 (N_7016,N_4067,N_5488);
or U7017 (N_7017,N_3881,N_4021);
or U7018 (N_7018,N_5697,N_3982);
or U7019 (N_7019,N_3205,N_5561);
nand U7020 (N_7020,N_3231,N_4943);
or U7021 (N_7021,N_4707,N_3227);
or U7022 (N_7022,N_5366,N_5273);
xnor U7023 (N_7023,N_5567,N_4230);
or U7024 (N_7024,N_4918,N_4037);
xnor U7025 (N_7025,N_4432,N_5678);
nand U7026 (N_7026,N_5730,N_5528);
xor U7027 (N_7027,N_4743,N_6014);
nand U7028 (N_7028,N_5042,N_4880);
and U7029 (N_7029,N_3454,N_3479);
or U7030 (N_7030,N_4302,N_4908);
nand U7031 (N_7031,N_4903,N_5495);
xnor U7032 (N_7032,N_4372,N_4972);
nor U7033 (N_7033,N_3909,N_3320);
nand U7034 (N_7034,N_5794,N_4527);
or U7035 (N_7035,N_4965,N_5549);
nand U7036 (N_7036,N_5318,N_5948);
nand U7037 (N_7037,N_3814,N_3405);
nor U7038 (N_7038,N_5574,N_4983);
nor U7039 (N_7039,N_3734,N_4861);
xnor U7040 (N_7040,N_3198,N_4087);
nor U7041 (N_7041,N_3366,N_5738);
xnor U7042 (N_7042,N_5881,N_5849);
xnor U7043 (N_7043,N_4658,N_5454);
xnor U7044 (N_7044,N_5856,N_3880);
and U7045 (N_7045,N_5222,N_3403);
nand U7046 (N_7046,N_3521,N_4575);
and U7047 (N_7047,N_5672,N_5956);
or U7048 (N_7048,N_3335,N_4110);
or U7049 (N_7049,N_3376,N_4353);
nor U7050 (N_7050,N_5308,N_4505);
xor U7051 (N_7051,N_6021,N_5996);
or U7052 (N_7052,N_3902,N_5465);
xnor U7053 (N_7053,N_5508,N_5975);
nor U7054 (N_7054,N_3150,N_3582);
nand U7055 (N_7055,N_6164,N_5668);
and U7056 (N_7056,N_5819,N_3216);
nor U7057 (N_7057,N_4695,N_5419);
xor U7058 (N_7058,N_3678,N_4778);
and U7059 (N_7059,N_4331,N_6171);
nor U7060 (N_7060,N_5893,N_4005);
and U7061 (N_7061,N_4754,N_4409);
and U7062 (N_7062,N_3924,N_3787);
xor U7063 (N_7063,N_5649,N_5339);
nor U7064 (N_7064,N_4364,N_6178);
and U7065 (N_7065,N_5147,N_5547);
xor U7066 (N_7066,N_4412,N_4036);
xnor U7067 (N_7067,N_3688,N_3156);
nor U7068 (N_7068,N_4194,N_5405);
xor U7069 (N_7069,N_5645,N_4869);
or U7070 (N_7070,N_5532,N_3600);
xor U7071 (N_7071,N_5632,N_5023);
and U7072 (N_7072,N_4570,N_4345);
nor U7073 (N_7073,N_3338,N_5647);
nand U7074 (N_7074,N_3158,N_3912);
or U7075 (N_7075,N_5441,N_6184);
or U7076 (N_7076,N_3465,N_4102);
and U7077 (N_7077,N_3603,N_4760);
and U7078 (N_7078,N_5336,N_3904);
nor U7079 (N_7079,N_4865,N_3864);
or U7080 (N_7080,N_3583,N_3680);
nand U7081 (N_7081,N_4092,N_5802);
nand U7082 (N_7082,N_3661,N_4628);
nand U7083 (N_7083,N_5614,N_6165);
nand U7084 (N_7084,N_4389,N_3659);
and U7085 (N_7085,N_4883,N_3491);
nand U7086 (N_7086,N_4748,N_5300);
or U7087 (N_7087,N_4580,N_3548);
xor U7088 (N_7088,N_3390,N_4486);
and U7089 (N_7089,N_5479,N_3730);
nor U7090 (N_7090,N_4931,N_4751);
nor U7091 (N_7091,N_4175,N_5797);
xor U7092 (N_7092,N_4147,N_5922);
nand U7093 (N_7093,N_3270,N_3980);
or U7094 (N_7094,N_3188,N_5928);
or U7095 (N_7095,N_4625,N_3414);
nand U7096 (N_7096,N_5154,N_5460);
and U7097 (N_7097,N_3646,N_6239);
xnor U7098 (N_7098,N_4192,N_3629);
xor U7099 (N_7099,N_4225,N_5019);
nor U7100 (N_7100,N_3613,N_3746);
xor U7101 (N_7101,N_4589,N_3571);
nor U7102 (N_7102,N_4493,N_3130);
and U7103 (N_7103,N_3413,N_4236);
xnor U7104 (N_7104,N_6222,N_4569);
or U7105 (N_7105,N_3268,N_4027);
or U7106 (N_7106,N_3179,N_3611);
or U7107 (N_7107,N_4081,N_5987);
xor U7108 (N_7108,N_3741,N_3689);
xnor U7109 (N_7109,N_5246,N_6152);
nor U7110 (N_7110,N_5093,N_5663);
nor U7111 (N_7111,N_3847,N_5783);
xor U7112 (N_7112,N_5747,N_5082);
nor U7113 (N_7113,N_5897,N_5212);
or U7114 (N_7114,N_5834,N_3314);
xor U7115 (N_7115,N_4884,N_3994);
nand U7116 (N_7116,N_5693,N_5504);
nor U7117 (N_7117,N_5404,N_3859);
or U7118 (N_7118,N_6228,N_3421);
xor U7119 (N_7119,N_6123,N_4424);
and U7120 (N_7120,N_5137,N_4949);
and U7121 (N_7121,N_4265,N_4000);
nand U7122 (N_7122,N_4680,N_3146);
and U7123 (N_7123,N_4163,N_5963);
nand U7124 (N_7124,N_3890,N_5050);
or U7125 (N_7125,N_3196,N_6245);
xnor U7126 (N_7126,N_4697,N_5260);
nor U7127 (N_7127,N_4669,N_3797);
nor U7128 (N_7128,N_4717,N_3715);
nand U7129 (N_7129,N_3534,N_6216);
and U7130 (N_7130,N_4349,N_3596);
nand U7131 (N_7131,N_4229,N_4592);
nor U7132 (N_7132,N_4772,N_5824);
xnor U7133 (N_7133,N_3879,N_3766);
and U7134 (N_7134,N_3291,N_4808);
xor U7135 (N_7135,N_5294,N_4007);
or U7136 (N_7136,N_4576,N_4386);
nand U7137 (N_7137,N_3391,N_5677);
or U7138 (N_7138,N_3673,N_5113);
or U7139 (N_7139,N_5912,N_3893);
xnor U7140 (N_7140,N_5889,N_5410);
and U7141 (N_7141,N_4464,N_3631);
nor U7142 (N_7142,N_5829,N_3612);
xnor U7143 (N_7143,N_6203,N_3239);
and U7144 (N_7144,N_3512,N_6010);
nand U7145 (N_7145,N_4491,N_3615);
xor U7146 (N_7146,N_5381,N_3392);
nor U7147 (N_7147,N_3724,N_3755);
and U7148 (N_7148,N_5592,N_4337);
xor U7149 (N_7149,N_4627,N_4593);
nor U7150 (N_7150,N_5918,N_3699);
nand U7151 (N_7151,N_5064,N_4621);
xor U7152 (N_7152,N_4630,N_4824);
nor U7153 (N_7153,N_3624,N_6093);
and U7154 (N_7154,N_6223,N_6192);
and U7155 (N_7155,N_5588,N_5597);
and U7156 (N_7156,N_3224,N_5428);
xor U7157 (N_7157,N_3540,N_4070);
nand U7158 (N_7158,N_4549,N_4781);
nand U7159 (N_7159,N_5571,N_5900);
xor U7160 (N_7160,N_5408,N_4805);
nand U7161 (N_7161,N_3711,N_4238);
or U7162 (N_7162,N_4591,N_5239);
and U7163 (N_7163,N_5480,N_5838);
nor U7164 (N_7164,N_5605,N_5387);
or U7165 (N_7165,N_5058,N_3171);
and U7166 (N_7166,N_3208,N_3747);
and U7167 (N_7167,N_4234,N_3316);
nand U7168 (N_7168,N_6166,N_6190);
and U7169 (N_7169,N_5332,N_4354);
nor U7170 (N_7170,N_6075,N_6105);
xor U7171 (N_7171,N_5704,N_5029);
nor U7172 (N_7172,N_4308,N_6036);
nor U7173 (N_7173,N_3259,N_3554);
and U7174 (N_7174,N_4587,N_4758);
or U7175 (N_7175,N_3164,N_3157);
nor U7176 (N_7176,N_5842,N_5282);
nand U7177 (N_7177,N_4927,N_3242);
and U7178 (N_7178,N_3745,N_4164);
or U7179 (N_7179,N_4008,N_5758);
and U7180 (N_7180,N_6225,N_5683);
or U7181 (N_7181,N_4089,N_4059);
and U7182 (N_7182,N_3402,N_5193);
or U7183 (N_7183,N_5160,N_5230);
xor U7184 (N_7184,N_3778,N_4040);
xnor U7185 (N_7185,N_5916,N_4817);
or U7186 (N_7186,N_6070,N_5074);
nor U7187 (N_7187,N_4633,N_3297);
xnor U7188 (N_7188,N_5040,N_3686);
xnor U7189 (N_7189,N_4062,N_4292);
or U7190 (N_7190,N_5350,N_3311);
nor U7191 (N_7191,N_3195,N_6137);
nand U7192 (N_7192,N_5613,N_5380);
and U7193 (N_7193,N_3418,N_6038);
and U7194 (N_7194,N_3651,N_5196);
xnor U7195 (N_7195,N_5401,N_3416);
and U7196 (N_7196,N_3988,N_4536);
and U7197 (N_7197,N_3794,N_5194);
and U7198 (N_7198,N_4049,N_4890);
xor U7199 (N_7199,N_5507,N_3127);
nor U7200 (N_7200,N_3536,N_4599);
nor U7201 (N_7201,N_5080,N_5694);
nand U7202 (N_7202,N_4033,N_6124);
nor U7203 (N_7203,N_5943,N_5413);
xor U7204 (N_7204,N_5890,N_5671);
nor U7205 (N_7205,N_5468,N_4532);
nor U7206 (N_7206,N_3677,N_5329);
xnor U7207 (N_7207,N_5687,N_3223);
xnor U7208 (N_7208,N_3163,N_3589);
nand U7209 (N_7209,N_3717,N_5171);
xor U7210 (N_7210,N_4454,N_5456);
xnor U7211 (N_7211,N_3339,N_5303);
xor U7212 (N_7212,N_4446,N_3305);
nor U7213 (N_7213,N_5778,N_3520);
nand U7214 (N_7214,N_3722,N_4472);
nor U7215 (N_7215,N_5598,N_4906);
nor U7216 (N_7216,N_4012,N_5135);
or U7217 (N_7217,N_5362,N_4065);
xnor U7218 (N_7218,N_5855,N_4371);
nand U7219 (N_7219,N_5579,N_4277);
xnor U7220 (N_7220,N_4673,N_3229);
and U7221 (N_7221,N_6161,N_3816);
nand U7222 (N_7222,N_4812,N_5861);
xor U7223 (N_7223,N_5391,N_6039);
nand U7224 (N_7224,N_4723,N_5241);
nor U7225 (N_7225,N_4963,N_4730);
or U7226 (N_7226,N_5263,N_3964);
nand U7227 (N_7227,N_4998,N_3210);
nand U7228 (N_7228,N_5364,N_5521);
nand U7229 (N_7229,N_4670,N_5600);
nand U7230 (N_7230,N_5980,N_5710);
nand U7231 (N_7231,N_5131,N_3773);
and U7232 (N_7232,N_4363,N_4898);
or U7233 (N_7233,N_3604,N_5001);
nor U7234 (N_7234,N_4607,N_5475);
nor U7235 (N_7235,N_3662,N_3608);
nand U7236 (N_7236,N_5685,N_4402);
and U7237 (N_7237,N_3628,N_4228);
and U7238 (N_7238,N_5220,N_6128);
and U7239 (N_7239,N_6226,N_3492);
or U7240 (N_7240,N_4171,N_4318);
xnor U7241 (N_7241,N_4258,N_3595);
and U7242 (N_7242,N_5585,N_5018);
and U7243 (N_7243,N_5913,N_3466);
xor U7244 (N_7244,N_5911,N_5101);
nand U7245 (N_7245,N_5853,N_3443);
or U7246 (N_7246,N_3576,N_3654);
and U7247 (N_7247,N_3920,N_4902);
or U7248 (N_7248,N_6072,N_4218);
nand U7249 (N_7249,N_4248,N_4641);
nor U7250 (N_7250,N_5382,N_4296);
nor U7251 (N_7251,N_4417,N_5522);
xor U7252 (N_7252,N_4809,N_6191);
xor U7253 (N_7253,N_5660,N_4471);
xor U7254 (N_7254,N_3936,N_4686);
nor U7255 (N_7255,N_4854,N_5538);
nor U7256 (N_7256,N_6063,N_4572);
nand U7257 (N_7257,N_3640,N_5616);
nand U7258 (N_7258,N_6054,N_5859);
nor U7259 (N_7259,N_4125,N_6118);
nor U7260 (N_7260,N_3385,N_5343);
or U7261 (N_7261,N_4602,N_4016);
or U7262 (N_7262,N_5799,N_4541);
nand U7263 (N_7263,N_3726,N_4442);
or U7264 (N_7264,N_5601,N_3933);
and U7265 (N_7265,N_3323,N_5971);
xor U7266 (N_7266,N_5580,N_5675);
and U7267 (N_7267,N_3440,N_3230);
nor U7268 (N_7268,N_4109,N_6099);
and U7269 (N_7269,N_4433,N_3779);
and U7270 (N_7270,N_5995,N_3221);
or U7271 (N_7271,N_5640,N_3265);
nor U7272 (N_7272,N_4520,N_5079);
nand U7273 (N_7273,N_5803,N_3302);
nor U7274 (N_7274,N_6140,N_4765);
or U7275 (N_7275,N_5776,N_4788);
nor U7276 (N_7276,N_5762,N_4636);
nor U7277 (N_7277,N_4190,N_3801);
and U7278 (N_7278,N_3447,N_3962);
nand U7279 (N_7279,N_4976,N_4771);
xnor U7280 (N_7280,N_3899,N_4186);
or U7281 (N_7281,N_3346,N_5003);
nand U7282 (N_7282,N_4826,N_4660);
nand U7283 (N_7283,N_3452,N_5754);
nor U7284 (N_7284,N_4540,N_4534);
xor U7285 (N_7285,N_4437,N_4682);
nand U7286 (N_7286,N_3349,N_5402);
xnor U7287 (N_7287,N_5761,N_4952);
nand U7288 (N_7288,N_5637,N_4263);
or U7289 (N_7289,N_3796,N_3399);
nor U7290 (N_7290,N_3438,N_4584);
nor U7291 (N_7291,N_3503,N_3597);
or U7292 (N_7292,N_5552,N_5656);
nor U7293 (N_7293,N_5156,N_4078);
and U7294 (N_7294,N_3285,N_5638);
and U7295 (N_7295,N_5166,N_3798);
nor U7296 (N_7296,N_5979,N_4768);
nand U7297 (N_7297,N_3675,N_4347);
or U7298 (N_7298,N_5236,N_6032);
nor U7299 (N_7299,N_3183,N_5476);
or U7300 (N_7300,N_5466,N_4046);
and U7301 (N_7301,N_4767,N_4135);
and U7302 (N_7302,N_3283,N_5543);
nand U7303 (N_7303,N_5107,N_3756);
or U7304 (N_7304,N_4537,N_5117);
nor U7305 (N_7305,N_3907,N_3788);
or U7306 (N_7306,N_5334,N_6210);
nor U7307 (N_7307,N_4635,N_3248);
xor U7308 (N_7308,N_3790,N_3712);
nand U7309 (N_7309,N_6181,N_5026);
or U7310 (N_7310,N_4544,N_4382);
nor U7311 (N_7311,N_5015,N_5365);
or U7312 (N_7312,N_4338,N_4822);
and U7313 (N_7313,N_4735,N_3609);
nor U7314 (N_7314,N_3626,N_5306);
or U7315 (N_7315,N_5737,N_5625);
and U7316 (N_7316,N_3823,N_4484);
and U7317 (N_7317,N_5201,N_5743);
nor U7318 (N_7318,N_4370,N_4671);
and U7319 (N_7319,N_3187,N_6199);
nand U7320 (N_7320,N_3697,N_4480);
nand U7321 (N_7321,N_3886,N_5005);
and U7322 (N_7322,N_4620,N_4792);
nor U7323 (N_7323,N_4483,N_5623);
xor U7324 (N_7324,N_5497,N_4237);
nand U7325 (N_7325,N_4664,N_3482);
and U7326 (N_7326,N_4098,N_4133);
nor U7327 (N_7327,N_6170,N_4397);
xor U7328 (N_7328,N_5968,N_6089);
or U7329 (N_7329,N_5110,N_4521);
xor U7330 (N_7330,N_4787,N_5828);
nand U7331 (N_7331,N_3125,N_5964);
nand U7332 (N_7332,N_4487,N_5557);
or U7333 (N_7333,N_5753,N_4239);
xor U7334 (N_7334,N_5031,N_5121);
nor U7335 (N_7335,N_4834,N_4206);
nor U7336 (N_7336,N_4646,N_3919);
or U7337 (N_7337,N_5902,N_3761);
xor U7338 (N_7338,N_4094,N_3269);
nor U7339 (N_7339,N_4101,N_5342);
xnor U7340 (N_7340,N_3906,N_6028);
xor U7341 (N_7341,N_3331,N_4897);
xor U7342 (N_7342,N_4079,N_5988);
nor U7343 (N_7343,N_4551,N_5400);
or U7344 (N_7344,N_4105,N_5165);
nand U7345 (N_7345,N_6150,N_4310);
nor U7346 (N_7346,N_6011,N_5688);
nand U7347 (N_7347,N_5490,N_5877);
xor U7348 (N_7348,N_3789,N_4891);
xnor U7349 (N_7349,N_5459,N_3464);
and U7350 (N_7350,N_4244,N_5551);
nor U7351 (N_7351,N_3949,N_4055);
nand U7352 (N_7352,N_5622,N_5711);
xnor U7353 (N_7353,N_4240,N_3708);
nor U7354 (N_7354,N_5933,N_6121);
or U7355 (N_7355,N_5027,N_4413);
nor U7356 (N_7356,N_6206,N_6008);
or U7357 (N_7357,N_3926,N_3889);
and U7358 (N_7358,N_5248,N_3838);
or U7359 (N_7359,N_3383,N_3979);
nor U7360 (N_7360,N_6110,N_6000);
or U7361 (N_7361,N_3683,N_3485);
nand U7362 (N_7362,N_3824,N_3154);
nor U7363 (N_7363,N_5326,N_5283);
or U7364 (N_7364,N_3129,N_3953);
nor U7365 (N_7365,N_4810,N_4858);
and U7366 (N_7366,N_6109,N_4637);
nand U7367 (N_7367,N_3685,N_3849);
and U7368 (N_7368,N_4933,N_4211);
or U7369 (N_7369,N_6163,N_5440);
and U7370 (N_7370,N_4392,N_3426);
xnor U7371 (N_7371,N_4679,N_5360);
nor U7372 (N_7372,N_3599,N_4373);
nand U7373 (N_7373,N_3577,N_3698);
xnor U7374 (N_7374,N_5570,N_4284);
and U7375 (N_7375,N_4973,N_5880);
nor U7376 (N_7376,N_5696,N_4223);
and U7377 (N_7377,N_6058,N_5319);
or U7378 (N_7378,N_6102,N_4789);
nand U7379 (N_7379,N_3898,N_4859);
or U7380 (N_7380,N_4724,N_6041);
nor U7381 (N_7381,N_3564,N_3553);
nor U7382 (N_7382,N_4198,N_5765);
or U7383 (N_7383,N_4871,N_6126);
and U7384 (N_7384,N_5496,N_3978);
nor U7385 (N_7385,N_5684,N_5749);
nand U7386 (N_7386,N_6079,N_5791);
xor U7387 (N_7387,N_4500,N_5037);
nor U7388 (N_7388,N_3148,N_3232);
nand U7389 (N_7389,N_4672,N_3460);
xor U7390 (N_7390,N_6212,N_5470);
nand U7391 (N_7391,N_4563,N_6234);
xnor U7392 (N_7392,N_4868,N_4550);
and U7393 (N_7393,N_3184,N_3542);
nor U7394 (N_7394,N_5972,N_5038);
nand U7395 (N_7395,N_5923,N_6056);
nor U7396 (N_7396,N_6059,N_3429);
xnor U7397 (N_7397,N_4348,N_4208);
and U7398 (N_7398,N_4744,N_4829);
or U7399 (N_7399,N_3817,N_5882);
and U7400 (N_7400,N_5839,N_6160);
nor U7401 (N_7401,N_5961,N_6156);
or U7402 (N_7402,N_5555,N_3344);
nor U7403 (N_7403,N_5539,N_3579);
or U7404 (N_7404,N_3410,N_3923);
or U7405 (N_7405,N_5780,N_5666);
and U7406 (N_7406,N_5060,N_3569);
xor U7407 (N_7407,N_3197,N_3234);
or U7408 (N_7408,N_3943,N_3702);
xor U7409 (N_7409,N_6211,N_3172);
xor U7410 (N_7410,N_3954,N_6069);
or U7411 (N_7411,N_3472,N_5293);
nor U7412 (N_7412,N_5734,N_6097);
or U7413 (N_7413,N_6205,N_6112);
nor U7414 (N_7414,N_3509,N_5793);
or U7415 (N_7415,N_6106,N_5578);
and U7416 (N_7416,N_3529,N_4665);
xor U7417 (N_7417,N_3852,N_3358);
or U7418 (N_7418,N_4511,N_3996);
nand U7419 (N_7419,N_5782,N_4619);
nand U7420 (N_7420,N_4246,N_4002);
nand U7421 (N_7421,N_4425,N_3951);
nor U7422 (N_7422,N_6130,N_4802);
nand U7423 (N_7423,N_3736,N_3993);
xnor U7424 (N_7424,N_5997,N_3250);
nand U7425 (N_7425,N_4774,N_3966);
or U7426 (N_7426,N_4220,N_6224);
xnor U7427 (N_7427,N_3947,N_5335);
xnor U7428 (N_7428,N_5821,N_5228);
and U7429 (N_7429,N_4923,N_4061);
and U7430 (N_7430,N_5034,N_4052);
xor U7431 (N_7431,N_5384,N_5464);
or U7432 (N_7432,N_4514,N_5204);
and U7433 (N_7433,N_5469,N_5378);
or U7434 (N_7434,N_4696,N_4281);
nand U7435 (N_7435,N_5940,N_3551);
xor U7436 (N_7436,N_4919,N_5870);
nor U7437 (N_7437,N_5806,N_5700);
xnor U7438 (N_7438,N_3750,N_5363);
nor U7439 (N_7439,N_4905,N_4138);
nand U7440 (N_7440,N_3568,N_5202);
xnor U7441 (N_7441,N_5102,N_4655);
xnor U7442 (N_7442,N_4928,N_5748);
xnor U7443 (N_7443,N_4662,N_6241);
and U7444 (N_7444,N_3995,N_5586);
or U7445 (N_7445,N_5843,N_6215);
and U7446 (N_7446,N_6147,N_5151);
nor U7447 (N_7447,N_5863,N_3288);
xnor U7448 (N_7448,N_4568,N_5233);
xor U7449 (N_7449,N_5390,N_3575);
or U7450 (N_7450,N_4156,N_4831);
nand U7451 (N_7451,N_4295,N_3511);
or U7452 (N_7452,N_3587,N_6029);
nand U7453 (N_7453,N_3967,N_3550);
nor U7454 (N_7454,N_4559,N_3960);
nor U7455 (N_7455,N_5016,N_3759);
xor U7456 (N_7456,N_4615,N_4519);
nor U7457 (N_7457,N_3393,N_5231);
nor U7458 (N_7458,N_4512,N_5051);
xnor U7459 (N_7459,N_3293,N_4266);
or U7460 (N_7460,N_5665,N_3585);
and U7461 (N_7461,N_5155,N_4394);
and U7462 (N_7462,N_4459,N_4009);
xnor U7463 (N_7463,N_4438,N_4790);
nand U7464 (N_7464,N_4848,N_3882);
and U7465 (N_7465,N_5158,N_5702);
and U7466 (N_7466,N_5297,N_4988);
nand U7467 (N_7467,N_4030,N_3313);
nor U7468 (N_7468,N_5004,N_6157);
nand U7469 (N_7469,N_4428,N_4911);
xnor U7470 (N_7470,N_5315,N_3435);
and U7471 (N_7471,N_6125,N_5591);
xor U7472 (N_7472,N_4014,N_4431);
nand U7473 (N_7473,N_6134,N_3769);
nand U7474 (N_7474,N_6053,N_4969);
or U7475 (N_7475,N_5446,N_3650);
or U7476 (N_7476,N_5067,N_4494);
nand U7477 (N_7477,N_5150,N_6020);
nand U7478 (N_7478,N_5624,N_4204);
or U7479 (N_7479,N_3984,N_5170);
nand U7480 (N_7480,N_4926,N_3837);
or U7481 (N_7481,N_4341,N_4384);
nand U7482 (N_7482,N_4867,N_5493);
or U7483 (N_7483,N_5846,N_4561);
xor U7484 (N_7484,N_4311,N_5159);
or U7485 (N_7485,N_3679,N_3867);
nor U7486 (N_7486,N_3362,N_4080);
or U7487 (N_7487,N_5929,N_4738);
xnor U7488 (N_7488,N_4506,N_4517);
and U7489 (N_7489,N_5767,N_3140);
nand U7490 (N_7490,N_3921,N_5695);
nor U7491 (N_7491,N_3638,N_3963);
nand U7492 (N_7492,N_3999,N_4557);
or U7493 (N_7493,N_4231,N_5801);
or U7494 (N_7494,N_5733,N_4737);
nand U7495 (N_7495,N_4270,N_6040);
nor U7496 (N_7496,N_3848,N_3433);
xor U7497 (N_7497,N_5712,N_4448);
nand U7498 (N_7498,N_3490,N_5698);
nor U7499 (N_7499,N_5206,N_4626);
and U7500 (N_7500,N_4473,N_5924);
xnor U7501 (N_7501,N_4917,N_6219);
nand U7502 (N_7502,N_6153,N_3295);
nand U7503 (N_7503,N_5299,N_5569);
and U7504 (N_7504,N_4714,N_6074);
nor U7505 (N_7505,N_5310,N_6246);
nor U7506 (N_7506,N_4994,N_3812);
or U7507 (N_7507,N_4961,N_3693);
xnor U7508 (N_7508,N_5375,N_4247);
nand U7509 (N_7509,N_3622,N_5727);
nor U7510 (N_7510,N_3928,N_5779);
or U7511 (N_7511,N_4913,N_5587);
nand U7512 (N_7512,N_6155,N_5562);
and U7513 (N_7513,N_5573,N_3458);
xor U7514 (N_7514,N_3493,N_4463);
nor U7515 (N_7515,N_4468,N_4255);
nand U7516 (N_7516,N_4343,N_4043);
xor U7517 (N_7517,N_4759,N_4533);
or U7518 (N_7518,N_6009,N_4088);
nor U7519 (N_7519,N_5448,N_3914);
or U7520 (N_7520,N_4920,N_4481);
and U7521 (N_7521,N_3240,N_3475);
nor U7522 (N_7522,N_4538,N_3214);
nor U7523 (N_7523,N_4260,N_3791);
nor U7524 (N_7524,N_3544,N_3417);
or U7525 (N_7525,N_4439,N_4600);
or U7526 (N_7526,N_4176,N_5901);
nor U7527 (N_7527,N_5760,N_3424);
or U7528 (N_7528,N_3598,N_5288);
nand U7529 (N_7529,N_5014,N_5584);
and U7530 (N_7530,N_3875,N_4676);
nand U7531 (N_7531,N_4529,N_5259);
nor U7532 (N_7532,N_4684,N_4567);
or U7533 (N_7533,N_4558,N_3526);
nor U7534 (N_7534,N_5374,N_3977);
and U7535 (N_7535,N_4017,N_4731);
nor U7536 (N_7536,N_3406,N_4169);
nor U7537 (N_7537,N_3828,N_4747);
and U7538 (N_7538,N_5396,N_5957);
xnor U7539 (N_7539,N_4691,N_4453);
or U7540 (N_7540,N_3253,N_4703);
nand U7541 (N_7541,N_5866,N_3703);
or U7542 (N_7542,N_4181,N_6090);
nor U7543 (N_7543,N_5937,N_5583);
nand U7544 (N_7544,N_4543,N_4916);
or U7545 (N_7545,N_5112,N_5984);
nor U7546 (N_7546,N_5272,N_3359);
nor U7547 (N_7547,N_5509,N_3322);
nor U7548 (N_7548,N_6200,N_5457);
nor U7549 (N_7549,N_4746,N_4546);
and U7550 (N_7550,N_4166,N_3998);
and U7551 (N_7551,N_5140,N_6162);
or U7552 (N_7552,N_5659,N_4019);
and U7553 (N_7553,N_4887,N_3593);
nand U7554 (N_7554,N_4278,N_3720);
nand U7555 (N_7555,N_4300,N_5970);
nor U7556 (N_7556,N_5338,N_5161);
nand U7557 (N_7557,N_6046,N_5435);
or U7558 (N_7558,N_3211,N_5084);
nand U7559 (N_7559,N_4167,N_4560);
nand U7560 (N_7560,N_5438,N_5772);
or U7561 (N_7561,N_3672,N_4904);
nor U7562 (N_7562,N_3189,N_3637);
xor U7563 (N_7563,N_5276,N_5826);
nor U7564 (N_7564,N_3939,N_4929);
nor U7565 (N_7565,N_6144,N_3618);
and U7566 (N_7566,N_6209,N_3641);
nor U7567 (N_7567,N_4806,N_4818);
xnor U7568 (N_7568,N_3892,N_5443);
and U7569 (N_7569,N_5198,N_4457);
nand U7570 (N_7570,N_4489,N_3185);
and U7571 (N_7571,N_4449,N_3937);
and U7572 (N_7572,N_4090,N_4722);
xor U7573 (N_7573,N_4116,N_5386);
or U7574 (N_7574,N_3537,N_4041);
nand U7575 (N_7575,N_4403,N_3774);
nor U7576 (N_7576,N_3704,N_3751);
nor U7577 (N_7577,N_3459,N_4830);
and U7578 (N_7578,N_4975,N_5506);
or U7579 (N_7579,N_4827,N_3557);
nor U7580 (N_7580,N_5145,N_3181);
nor U7581 (N_7581,N_3363,N_5831);
nor U7582 (N_7582,N_3318,N_5947);
nor U7583 (N_7583,N_4650,N_5432);
nor U7584 (N_7584,N_4864,N_3555);
nand U7585 (N_7585,N_5541,N_5081);
nor U7586 (N_7586,N_6131,N_3245);
nand U7587 (N_7587,N_5904,N_5990);
or U7588 (N_7588,N_5120,N_4939);
nand U7589 (N_7589,N_3991,N_4571);
xor U7590 (N_7590,N_4689,N_4128);
and U7591 (N_7591,N_3968,N_5146);
and U7592 (N_7592,N_3799,N_3476);
and U7593 (N_7593,N_6249,N_5848);
nor U7594 (N_7594,N_5888,N_3327);
nand U7595 (N_7595,N_4482,N_5285);
nor U7596 (N_7596,N_5518,N_4323);
xnor U7597 (N_7597,N_3866,N_6084);
nand U7598 (N_7598,N_5340,N_4451);
xnor U7599 (N_7599,N_3681,N_5477);
or U7600 (N_7600,N_5268,N_5321);
nand U7601 (N_7601,N_5572,N_5279);
nand U7602 (N_7602,N_4380,N_3360);
nand U7603 (N_7603,N_3489,N_5789);
or U7604 (N_7604,N_5686,N_5010);
nand U7605 (N_7605,N_4361,N_5116);
or U7606 (N_7606,N_5960,N_5286);
xnor U7607 (N_7607,N_4458,N_4290);
nand U7608 (N_7608,N_6175,N_4162);
or U7609 (N_7609,N_5835,N_3463);
or U7610 (N_7610,N_4357,N_4117);
or U7611 (N_7611,N_5862,N_3367);
nor U7612 (N_7612,N_3166,N_5728);
nand U7613 (N_7613,N_4400,N_5514);
and U7614 (N_7614,N_5550,N_4477);
or U7615 (N_7615,N_6244,N_4974);
nor U7616 (N_7616,N_6232,N_4075);
nand U7617 (N_7617,N_5745,N_4852);
xnor U7618 (N_7618,N_5430,N_6208);
xor U7619 (N_7619,N_3563,N_4444);
and U7620 (N_7620,N_5981,N_4150);
nand U7621 (N_7621,N_5621,N_4547);
or U7622 (N_7622,N_4708,N_3706);
and U7623 (N_7623,N_4129,N_5199);
xor U7624 (N_7624,N_4819,N_5191);
nand U7625 (N_7625,N_4184,N_5969);
nor U7626 (N_7626,N_4632,N_4876);
nor U7627 (N_7627,N_4044,N_6087);
nor U7628 (N_7628,N_3805,N_4495);
or U7629 (N_7629,N_6217,N_5071);
xnor U7630 (N_7630,N_6055,N_3985);
nand U7631 (N_7631,N_5070,N_4811);
and U7632 (N_7632,N_5253,N_5305);
nor U7633 (N_7633,N_3407,N_5173);
and U7634 (N_7634,N_4224,N_6078);
or U7635 (N_7635,N_3284,N_4797);
nor U7636 (N_7636,N_5132,N_4465);
and U7637 (N_7637,N_4847,N_5128);
nor U7638 (N_7638,N_3948,N_4957);
xnor U7639 (N_7639,N_5978,N_4888);
xnor U7640 (N_7640,N_4999,N_4687);
nor U7641 (N_7641,N_4032,N_4123);
xnor U7642 (N_7642,N_4715,N_4427);
or U7643 (N_7643,N_3911,N_4047);
or U7644 (N_7644,N_4885,N_3591);
or U7645 (N_7645,N_4814,N_5565);
and U7646 (N_7646,N_3445,N_6004);
nor U7647 (N_7647,N_6127,N_6012);
and U7648 (N_7648,N_4945,N_6198);
and U7649 (N_7649,N_5757,N_4006);
or U7650 (N_7650,N_3468,N_5494);
nand U7651 (N_7651,N_5847,N_6180);
and U7652 (N_7652,N_3299,N_4578);
and U7653 (N_7653,N_5850,N_4804);
xor U7654 (N_7654,N_6066,N_5938);
or U7655 (N_7655,N_5770,N_4678);
xor U7656 (N_7656,N_4388,N_5563);
nor U7657 (N_7657,N_3729,N_4362);
or U7658 (N_7658,N_5650,N_5486);
nand U7659 (N_7659,N_4525,N_4073);
or U7660 (N_7660,N_4020,N_4616);
nand U7661 (N_7661,N_4704,N_3162);
xor U7662 (N_7662,N_5353,N_5225);
and U7663 (N_7663,N_4307,N_5993);
xnor U7664 (N_7664,N_5322,N_5667);
nor U7665 (N_7665,N_3836,N_5262);
nand U7666 (N_7666,N_3292,N_3498);
or U7667 (N_7667,N_5744,N_3861);
nor U7668 (N_7668,N_4243,N_4298);
nand U7669 (N_7669,N_5257,N_4429);
and U7670 (N_7670,N_4460,N_3395);
or U7671 (N_7671,N_3145,N_3131);
nor U7672 (N_7672,N_3983,N_5673);
xor U7673 (N_7673,N_5208,N_3442);
nand U7674 (N_7674,N_3565,N_6068);
nor U7675 (N_7675,N_4333,N_4742);
xnor U7676 (N_7676,N_3474,N_4209);
and U7677 (N_7677,N_4082,N_5920);
xor U7678 (N_7678,N_6076,N_3760);
nand U7679 (N_7679,N_4784,N_4598);
nand U7680 (N_7680,N_3959,N_4359);
nor U7681 (N_7681,N_3821,N_3696);
nor U7682 (N_7682,N_5357,N_5238);
and U7683 (N_7683,N_5179,N_4185);
nor U7684 (N_7684,N_4421,N_5106);
xor U7685 (N_7685,N_3420,N_3739);
or U7686 (N_7686,N_4644,N_5653);
xnor U7687 (N_7687,N_3496,N_5119);
and U7688 (N_7688,N_4320,N_3203);
nor U7689 (N_7689,N_5250,N_4846);
nor U7690 (N_7690,N_4197,N_3938);
and U7691 (N_7691,N_5429,N_5525);
xor U7692 (N_7692,N_5328,N_5224);
nand U7693 (N_7693,N_4597,N_4466);
nor U7694 (N_7694,N_5752,N_3354);
and U7695 (N_7695,N_4667,N_5445);
nor U7696 (N_7696,N_5858,N_5092);
or U7697 (N_7697,N_5379,N_4289);
nand U7698 (N_7698,N_3522,N_6007);
or U7699 (N_7699,N_3244,N_3345);
and U7700 (N_7700,N_4900,N_6133);
and U7701 (N_7701,N_5371,N_3457);
xnor U7702 (N_7702,N_5455,N_4645);
nor U7703 (N_7703,N_3449,N_5875);
xnor U7704 (N_7704,N_3481,N_3581);
nor U7705 (N_7705,N_3862,N_3839);
nor U7706 (N_7706,N_6030,N_4038);
and U7707 (N_7707,N_3186,N_4145);
nor U7708 (N_7708,N_3152,N_5816);
nand U7709 (N_7709,N_3257,N_3298);
or U7710 (N_7710,N_5397,N_4405);
or U7711 (N_7711,N_5453,N_4226);
and U7712 (N_7712,N_5718,N_3133);
or U7713 (N_7713,N_3687,N_4415);
nand U7714 (N_7714,N_4217,N_3237);
xnor U7715 (N_7715,N_5648,N_3350);
and U7716 (N_7716,N_4652,N_6048);
nor U7717 (N_7717,N_5510,N_6176);
or U7718 (N_7718,N_3559,N_3901);
nand U7719 (N_7719,N_4875,N_5061);
nor U7720 (N_7720,N_5232,N_4971);
and U7721 (N_7721,N_6235,N_3425);
and U7722 (N_7722,N_4798,N_3279);
nand U7723 (N_7723,N_4367,N_4474);
nand U7724 (N_7724,N_4251,N_3543);
or U7725 (N_7725,N_4478,N_4174);
nand U7726 (N_7726,N_3625,N_4946);
and U7727 (N_7727,N_5985,N_5280);
xnor U7728 (N_7728,N_5512,N_4168);
nor U7729 (N_7729,N_5553,N_5237);
and U7730 (N_7730,N_3513,N_4986);
and U7731 (N_7731,N_4841,N_4180);
nor U7732 (N_7732,N_3161,N_4820);
xor U7733 (N_7733,N_5247,N_3874);
xor U7734 (N_7734,N_3941,N_5311);
nand U7735 (N_7735,N_3885,N_4763);
nand U7736 (N_7736,N_3272,N_5785);
nand U7737 (N_7737,N_3262,N_4470);
xor U7738 (N_7738,N_3155,N_5417);
xnor U7739 (N_7739,N_5188,N_3353);
or U7740 (N_7740,N_5124,N_4418);
xnor U7741 (N_7741,N_5249,N_5919);
and U7742 (N_7742,N_4757,N_5207);
xor U7743 (N_7743,N_4322,N_4516);
nand U7744 (N_7744,N_3478,N_5815);
nor U7745 (N_7745,N_3386,N_3381);
nor U7746 (N_7746,N_4698,N_5354);
nand U7747 (N_7747,N_4064,N_3684);
or U7748 (N_7748,N_5903,N_3908);
nor U7749 (N_7749,N_4042,N_4941);
nor U7750 (N_7750,N_4490,N_4178);
xnor U7751 (N_7751,N_4736,N_5936);
and U7752 (N_7752,N_5742,N_4647);
nand U7753 (N_7753,N_6120,N_3488);
or U7754 (N_7754,N_5091,N_5769);
nor U7755 (N_7755,N_3844,N_4199);
xnor U7756 (N_7756,N_3450,N_3981);
xnor U7757 (N_7757,N_5906,N_4306);
nor U7758 (N_7758,N_3502,N_6067);
or U7759 (N_7759,N_3254,N_5724);
nand U7760 (N_7760,N_4609,N_3484);
nor U7761 (N_7761,N_5629,N_5139);
nand U7762 (N_7762,N_4649,N_4542);
xor U7763 (N_7763,N_3709,N_3804);
xor U7764 (N_7764,N_5153,N_4701);
or U7765 (N_7765,N_3142,N_5447);
or U7766 (N_7766,N_5823,N_3304);
and U7767 (N_7767,N_4654,N_5915);
and U7768 (N_7768,N_4188,N_4315);
nand U7769 (N_7769,N_5269,N_3811);
nand U7770 (N_7770,N_6143,N_5517);
and U7771 (N_7771,N_3931,N_5210);
nand U7772 (N_7772,N_4924,N_5049);
nand U7773 (N_7773,N_4910,N_3842);
nand U7774 (N_7774,N_4899,N_3134);
nor U7775 (N_7775,N_3143,N_5590);
nor U7776 (N_7776,N_4878,N_6173);
xor U7777 (N_7777,N_5105,N_4577);
or U7778 (N_7778,N_3855,N_5714);
or U7779 (N_7779,N_4825,N_4740);
and U7780 (N_7780,N_3539,N_5530);
and U7781 (N_7781,N_3153,N_5452);
and U7782 (N_7782,N_3971,N_6117);
and U7783 (N_7783,N_4604,N_3856);
xor U7784 (N_7784,N_4685,N_4462);
nand U7785 (N_7785,N_3786,N_4257);
nand U7786 (N_7786,N_5103,N_4984);
or U7787 (N_7787,N_3558,N_4173);
or U7788 (N_7788,N_3918,N_4996);
xor U7789 (N_7789,N_5811,N_3915);
nand U7790 (N_7790,N_4750,N_5383);
xnor U7791 (N_7791,N_3264,N_6047);
and U7792 (N_7792,N_4651,N_3233);
or U7793 (N_7793,N_3744,N_4839);
xnor U7794 (N_7794,N_4977,N_5436);
nor U7795 (N_7795,N_5392,N_4915);
and U7796 (N_7796,N_4153,N_5840);
nand U7797 (N_7797,N_4716,N_5289);
nor U7798 (N_7798,N_3247,N_5726);
and U7799 (N_7799,N_4056,N_5484);
nor U7800 (N_7800,N_4368,N_5751);
xor U7801 (N_7801,N_4301,N_5376);
and U7802 (N_7802,N_5784,N_3389);
nand U7803 (N_7803,N_3863,N_6195);
or U7804 (N_7804,N_4488,N_5763);
and U7805 (N_7805,N_3274,N_3649);
nand U7806 (N_7806,N_5053,N_3368);
nor U7807 (N_7807,N_5682,N_3764);
xor U7808 (N_7808,N_5878,N_5939);
nor U7809 (N_7809,N_5559,N_4411);
nor U7810 (N_7810,N_4562,N_4113);
nor U7811 (N_7811,N_5032,N_5356);
and U7812 (N_7812,N_3854,N_3947);
nor U7813 (N_7813,N_4763,N_5556);
nand U7814 (N_7814,N_5131,N_6012);
nand U7815 (N_7815,N_3318,N_4467);
nor U7816 (N_7816,N_4993,N_4538);
and U7817 (N_7817,N_5692,N_3136);
or U7818 (N_7818,N_4599,N_3510);
nand U7819 (N_7819,N_4646,N_5153);
nand U7820 (N_7820,N_5885,N_3565);
or U7821 (N_7821,N_5762,N_3894);
or U7822 (N_7822,N_4936,N_3548);
or U7823 (N_7823,N_4688,N_4283);
nand U7824 (N_7824,N_4986,N_4705);
nand U7825 (N_7825,N_5346,N_3165);
nand U7826 (N_7826,N_3366,N_4382);
or U7827 (N_7827,N_6161,N_6052);
xnor U7828 (N_7828,N_3439,N_6242);
and U7829 (N_7829,N_3381,N_4463);
xnor U7830 (N_7830,N_5047,N_4578);
and U7831 (N_7831,N_6083,N_3880);
or U7832 (N_7832,N_6242,N_4023);
nor U7833 (N_7833,N_5680,N_4927);
nor U7834 (N_7834,N_6165,N_4462);
and U7835 (N_7835,N_3507,N_3804);
or U7836 (N_7836,N_3844,N_4922);
and U7837 (N_7837,N_4090,N_4318);
xor U7838 (N_7838,N_5633,N_3554);
nor U7839 (N_7839,N_5714,N_5438);
or U7840 (N_7840,N_5048,N_6027);
nor U7841 (N_7841,N_3945,N_5073);
and U7842 (N_7842,N_4272,N_5586);
or U7843 (N_7843,N_4013,N_5887);
xnor U7844 (N_7844,N_3452,N_3571);
and U7845 (N_7845,N_4804,N_4243);
and U7846 (N_7846,N_4168,N_6076);
and U7847 (N_7847,N_5706,N_6012);
and U7848 (N_7848,N_6062,N_4014);
nand U7849 (N_7849,N_3442,N_3665);
nand U7850 (N_7850,N_6076,N_4373);
xor U7851 (N_7851,N_4763,N_4271);
xor U7852 (N_7852,N_5345,N_3603);
and U7853 (N_7853,N_6103,N_3300);
and U7854 (N_7854,N_6131,N_6051);
nor U7855 (N_7855,N_4920,N_5503);
or U7856 (N_7856,N_4577,N_5367);
or U7857 (N_7857,N_5607,N_5739);
nand U7858 (N_7858,N_4796,N_6134);
or U7859 (N_7859,N_5599,N_5190);
or U7860 (N_7860,N_3150,N_3680);
or U7861 (N_7861,N_4739,N_5781);
nand U7862 (N_7862,N_4984,N_6092);
nand U7863 (N_7863,N_5292,N_5631);
and U7864 (N_7864,N_4688,N_4715);
or U7865 (N_7865,N_3944,N_3793);
xor U7866 (N_7866,N_5458,N_6215);
nand U7867 (N_7867,N_6010,N_4000);
xor U7868 (N_7868,N_3549,N_5852);
xor U7869 (N_7869,N_5554,N_4551);
nand U7870 (N_7870,N_5604,N_5281);
xnor U7871 (N_7871,N_4844,N_4225);
or U7872 (N_7872,N_3423,N_3820);
xnor U7873 (N_7873,N_3171,N_5399);
nand U7874 (N_7874,N_4462,N_3794);
and U7875 (N_7875,N_4668,N_4295);
nand U7876 (N_7876,N_3439,N_4363);
nand U7877 (N_7877,N_3991,N_4513);
nand U7878 (N_7878,N_5133,N_6011);
nand U7879 (N_7879,N_3167,N_4353);
nand U7880 (N_7880,N_4060,N_5872);
and U7881 (N_7881,N_6100,N_5025);
or U7882 (N_7882,N_5176,N_6043);
or U7883 (N_7883,N_3798,N_3502);
or U7884 (N_7884,N_3839,N_4335);
or U7885 (N_7885,N_6130,N_3966);
nor U7886 (N_7886,N_6186,N_4495);
nand U7887 (N_7887,N_4062,N_4268);
nor U7888 (N_7888,N_5106,N_6103);
and U7889 (N_7889,N_3766,N_5010);
nor U7890 (N_7890,N_4558,N_4993);
nor U7891 (N_7891,N_5435,N_5641);
xnor U7892 (N_7892,N_3915,N_3732);
and U7893 (N_7893,N_4148,N_3763);
and U7894 (N_7894,N_3299,N_4854);
xnor U7895 (N_7895,N_4358,N_5636);
xnor U7896 (N_7896,N_5799,N_3696);
xor U7897 (N_7897,N_4341,N_5979);
and U7898 (N_7898,N_5796,N_5065);
nor U7899 (N_7899,N_6081,N_5427);
and U7900 (N_7900,N_4232,N_4704);
and U7901 (N_7901,N_5242,N_4002);
and U7902 (N_7902,N_6171,N_4428);
nor U7903 (N_7903,N_6167,N_3322);
or U7904 (N_7904,N_4799,N_5748);
nand U7905 (N_7905,N_4359,N_4934);
or U7906 (N_7906,N_3380,N_5938);
nor U7907 (N_7907,N_3643,N_5311);
or U7908 (N_7908,N_4426,N_5675);
nand U7909 (N_7909,N_4958,N_5541);
or U7910 (N_7910,N_5347,N_4312);
or U7911 (N_7911,N_3293,N_4208);
xnor U7912 (N_7912,N_3791,N_4736);
nor U7913 (N_7913,N_5517,N_5961);
or U7914 (N_7914,N_6155,N_3588);
nor U7915 (N_7915,N_4716,N_5701);
and U7916 (N_7916,N_5668,N_5268);
or U7917 (N_7917,N_4746,N_3632);
or U7918 (N_7918,N_3941,N_5355);
or U7919 (N_7919,N_4415,N_3555);
nand U7920 (N_7920,N_5532,N_5807);
nor U7921 (N_7921,N_5178,N_4311);
or U7922 (N_7922,N_3912,N_5280);
nand U7923 (N_7923,N_4053,N_6031);
or U7924 (N_7924,N_6053,N_3288);
nor U7925 (N_7925,N_4186,N_4579);
or U7926 (N_7926,N_3691,N_5199);
nor U7927 (N_7927,N_4612,N_5676);
or U7928 (N_7928,N_5860,N_5527);
and U7929 (N_7929,N_5409,N_4847);
or U7930 (N_7930,N_6041,N_4623);
nor U7931 (N_7931,N_4017,N_4891);
nand U7932 (N_7932,N_5974,N_5955);
xor U7933 (N_7933,N_4392,N_5795);
nand U7934 (N_7934,N_5799,N_3299);
and U7935 (N_7935,N_5324,N_5635);
or U7936 (N_7936,N_4479,N_6218);
nor U7937 (N_7937,N_5558,N_4352);
nand U7938 (N_7938,N_5117,N_6133);
nor U7939 (N_7939,N_4820,N_4006);
xnor U7940 (N_7940,N_4249,N_3936);
or U7941 (N_7941,N_5524,N_3821);
xnor U7942 (N_7942,N_3577,N_5159);
xor U7943 (N_7943,N_5881,N_3383);
or U7944 (N_7944,N_5586,N_4863);
nor U7945 (N_7945,N_6024,N_4154);
or U7946 (N_7946,N_5637,N_5186);
nor U7947 (N_7947,N_6015,N_3263);
nand U7948 (N_7948,N_4161,N_5289);
nand U7949 (N_7949,N_4140,N_4778);
xor U7950 (N_7950,N_3315,N_5883);
and U7951 (N_7951,N_3934,N_5280);
and U7952 (N_7952,N_4060,N_5731);
and U7953 (N_7953,N_4069,N_4671);
nor U7954 (N_7954,N_4577,N_4915);
and U7955 (N_7955,N_4601,N_5185);
nor U7956 (N_7956,N_6009,N_6223);
nor U7957 (N_7957,N_5804,N_5142);
or U7958 (N_7958,N_4779,N_5300);
and U7959 (N_7959,N_3969,N_3854);
nor U7960 (N_7960,N_6064,N_5581);
nand U7961 (N_7961,N_4498,N_4927);
xor U7962 (N_7962,N_5773,N_4560);
or U7963 (N_7963,N_4823,N_6005);
nand U7964 (N_7964,N_4950,N_3934);
xor U7965 (N_7965,N_3978,N_5461);
nor U7966 (N_7966,N_3554,N_5627);
nand U7967 (N_7967,N_3176,N_4772);
and U7968 (N_7968,N_3710,N_3980);
xor U7969 (N_7969,N_4117,N_3993);
xnor U7970 (N_7970,N_3371,N_3612);
or U7971 (N_7971,N_3854,N_5344);
xnor U7972 (N_7972,N_3526,N_3976);
nand U7973 (N_7973,N_3811,N_3752);
and U7974 (N_7974,N_5446,N_4325);
nand U7975 (N_7975,N_4584,N_5104);
nor U7976 (N_7976,N_5834,N_3188);
or U7977 (N_7977,N_3305,N_4040);
nor U7978 (N_7978,N_5870,N_5149);
nand U7979 (N_7979,N_5624,N_3268);
nand U7980 (N_7980,N_3829,N_6008);
xnor U7981 (N_7981,N_4756,N_5767);
or U7982 (N_7982,N_3272,N_3447);
xnor U7983 (N_7983,N_4897,N_6154);
nand U7984 (N_7984,N_5443,N_3638);
and U7985 (N_7985,N_5345,N_5229);
xnor U7986 (N_7986,N_4534,N_4641);
nand U7987 (N_7987,N_4663,N_5003);
or U7988 (N_7988,N_5806,N_3129);
nor U7989 (N_7989,N_3191,N_3484);
and U7990 (N_7990,N_3211,N_4784);
nand U7991 (N_7991,N_3512,N_5919);
nand U7992 (N_7992,N_5903,N_4191);
xor U7993 (N_7993,N_6005,N_3864);
xor U7994 (N_7994,N_4691,N_4680);
and U7995 (N_7995,N_3379,N_4721);
and U7996 (N_7996,N_5105,N_4636);
nor U7997 (N_7997,N_4400,N_5321);
and U7998 (N_7998,N_3315,N_5989);
nor U7999 (N_7999,N_5510,N_4000);
xor U8000 (N_8000,N_3616,N_6035);
or U8001 (N_8001,N_4985,N_4654);
or U8002 (N_8002,N_5418,N_5252);
xor U8003 (N_8003,N_4254,N_5063);
and U8004 (N_8004,N_5345,N_4990);
nor U8005 (N_8005,N_6151,N_3715);
or U8006 (N_8006,N_5092,N_4007);
nor U8007 (N_8007,N_4567,N_4634);
and U8008 (N_8008,N_4072,N_6056);
or U8009 (N_8009,N_4011,N_5973);
and U8010 (N_8010,N_3501,N_5506);
nor U8011 (N_8011,N_4189,N_5571);
and U8012 (N_8012,N_3165,N_5180);
and U8013 (N_8013,N_5827,N_4444);
nor U8014 (N_8014,N_3657,N_5126);
and U8015 (N_8015,N_4173,N_5630);
and U8016 (N_8016,N_3206,N_4478);
and U8017 (N_8017,N_4054,N_5255);
nand U8018 (N_8018,N_3803,N_6231);
nor U8019 (N_8019,N_4141,N_3982);
nand U8020 (N_8020,N_5907,N_4329);
or U8021 (N_8021,N_4471,N_3878);
xnor U8022 (N_8022,N_4208,N_5016);
xor U8023 (N_8023,N_5136,N_5313);
and U8024 (N_8024,N_5892,N_4770);
nand U8025 (N_8025,N_5985,N_3710);
xnor U8026 (N_8026,N_3709,N_3263);
nor U8027 (N_8027,N_5110,N_4480);
or U8028 (N_8028,N_4794,N_5289);
xor U8029 (N_8029,N_4782,N_5208);
nor U8030 (N_8030,N_4983,N_5317);
nand U8031 (N_8031,N_5361,N_4254);
nand U8032 (N_8032,N_3334,N_3893);
and U8033 (N_8033,N_4816,N_3813);
nand U8034 (N_8034,N_4135,N_4655);
nand U8035 (N_8035,N_3708,N_4826);
xor U8036 (N_8036,N_5110,N_4277);
xnor U8037 (N_8037,N_4761,N_5847);
xnor U8038 (N_8038,N_6023,N_5988);
nand U8039 (N_8039,N_5764,N_5959);
nor U8040 (N_8040,N_3272,N_5786);
and U8041 (N_8041,N_5532,N_6052);
xor U8042 (N_8042,N_6174,N_3995);
nand U8043 (N_8043,N_3972,N_3448);
and U8044 (N_8044,N_6030,N_4410);
nor U8045 (N_8045,N_4806,N_5387);
nor U8046 (N_8046,N_3654,N_4274);
or U8047 (N_8047,N_5626,N_3911);
nor U8048 (N_8048,N_3881,N_4104);
xnor U8049 (N_8049,N_3687,N_5571);
or U8050 (N_8050,N_6094,N_4571);
and U8051 (N_8051,N_4333,N_3785);
nand U8052 (N_8052,N_3966,N_3272);
nor U8053 (N_8053,N_4824,N_3374);
and U8054 (N_8054,N_3680,N_3571);
or U8055 (N_8055,N_3842,N_6183);
and U8056 (N_8056,N_5415,N_6081);
xnor U8057 (N_8057,N_3599,N_4275);
xnor U8058 (N_8058,N_3810,N_4037);
nand U8059 (N_8059,N_3663,N_3910);
nor U8060 (N_8060,N_5406,N_5322);
xnor U8061 (N_8061,N_6132,N_3498);
xor U8062 (N_8062,N_3409,N_4940);
nor U8063 (N_8063,N_6041,N_4635);
or U8064 (N_8064,N_4621,N_4107);
and U8065 (N_8065,N_4342,N_4637);
nand U8066 (N_8066,N_6065,N_4730);
and U8067 (N_8067,N_4955,N_5951);
nor U8068 (N_8068,N_5732,N_4134);
nor U8069 (N_8069,N_5735,N_4557);
nand U8070 (N_8070,N_5370,N_3936);
nand U8071 (N_8071,N_3198,N_5519);
and U8072 (N_8072,N_5054,N_3702);
nand U8073 (N_8073,N_3525,N_5253);
nor U8074 (N_8074,N_3784,N_5941);
nand U8075 (N_8075,N_4334,N_4955);
nor U8076 (N_8076,N_4829,N_5194);
nor U8077 (N_8077,N_5353,N_4325);
xor U8078 (N_8078,N_3127,N_4895);
nand U8079 (N_8079,N_4630,N_4476);
nor U8080 (N_8080,N_5165,N_3991);
xor U8081 (N_8081,N_4182,N_3844);
or U8082 (N_8082,N_4013,N_3904);
and U8083 (N_8083,N_4235,N_4019);
nor U8084 (N_8084,N_4796,N_3347);
nand U8085 (N_8085,N_4811,N_5593);
or U8086 (N_8086,N_3177,N_5000);
xor U8087 (N_8087,N_4359,N_3593);
and U8088 (N_8088,N_5133,N_4706);
or U8089 (N_8089,N_5056,N_4143);
xnor U8090 (N_8090,N_3425,N_5230);
nor U8091 (N_8091,N_4938,N_4758);
nand U8092 (N_8092,N_5042,N_5143);
or U8093 (N_8093,N_5225,N_3240);
nor U8094 (N_8094,N_3380,N_6200);
and U8095 (N_8095,N_4645,N_6098);
nor U8096 (N_8096,N_4286,N_4389);
xor U8097 (N_8097,N_4088,N_3234);
nand U8098 (N_8098,N_3950,N_5921);
and U8099 (N_8099,N_4321,N_5960);
or U8100 (N_8100,N_5568,N_3432);
or U8101 (N_8101,N_4165,N_3194);
nand U8102 (N_8102,N_5665,N_3460);
xnor U8103 (N_8103,N_6224,N_5650);
and U8104 (N_8104,N_4738,N_4826);
or U8105 (N_8105,N_5316,N_3630);
xnor U8106 (N_8106,N_4515,N_6247);
xor U8107 (N_8107,N_4856,N_5325);
and U8108 (N_8108,N_5210,N_5949);
xor U8109 (N_8109,N_5691,N_5230);
xor U8110 (N_8110,N_5507,N_5657);
nand U8111 (N_8111,N_3255,N_4942);
nor U8112 (N_8112,N_5255,N_5100);
or U8113 (N_8113,N_3221,N_5301);
and U8114 (N_8114,N_6032,N_5718);
xnor U8115 (N_8115,N_3573,N_5834);
nand U8116 (N_8116,N_5808,N_4574);
nor U8117 (N_8117,N_5736,N_4449);
and U8118 (N_8118,N_6038,N_5565);
or U8119 (N_8119,N_5432,N_4668);
and U8120 (N_8120,N_4916,N_5219);
nand U8121 (N_8121,N_5039,N_3411);
or U8122 (N_8122,N_6169,N_4397);
or U8123 (N_8123,N_4148,N_5451);
xnor U8124 (N_8124,N_4880,N_3814);
or U8125 (N_8125,N_5467,N_5906);
and U8126 (N_8126,N_3301,N_3805);
and U8127 (N_8127,N_3479,N_3331);
xnor U8128 (N_8128,N_4023,N_5322);
nor U8129 (N_8129,N_4776,N_5235);
and U8130 (N_8130,N_5069,N_5922);
xnor U8131 (N_8131,N_3716,N_3556);
and U8132 (N_8132,N_5458,N_3752);
nor U8133 (N_8133,N_5804,N_4048);
and U8134 (N_8134,N_5644,N_4460);
xnor U8135 (N_8135,N_5646,N_5804);
nor U8136 (N_8136,N_5941,N_3282);
or U8137 (N_8137,N_5962,N_3156);
or U8138 (N_8138,N_5683,N_4877);
nand U8139 (N_8139,N_3282,N_4536);
nor U8140 (N_8140,N_5046,N_6219);
or U8141 (N_8141,N_4768,N_4580);
or U8142 (N_8142,N_5010,N_3833);
and U8143 (N_8143,N_5924,N_5858);
nand U8144 (N_8144,N_3489,N_4772);
xor U8145 (N_8145,N_5455,N_5115);
and U8146 (N_8146,N_3459,N_5249);
or U8147 (N_8147,N_4850,N_3427);
and U8148 (N_8148,N_3570,N_4583);
xnor U8149 (N_8149,N_5081,N_4778);
or U8150 (N_8150,N_5390,N_5202);
nand U8151 (N_8151,N_4592,N_5707);
or U8152 (N_8152,N_4165,N_6190);
and U8153 (N_8153,N_5174,N_3127);
nand U8154 (N_8154,N_3845,N_6013);
or U8155 (N_8155,N_3805,N_4660);
or U8156 (N_8156,N_3324,N_3153);
and U8157 (N_8157,N_4033,N_4733);
nor U8158 (N_8158,N_3696,N_4573);
or U8159 (N_8159,N_4311,N_4251);
xor U8160 (N_8160,N_5187,N_5191);
nor U8161 (N_8161,N_6117,N_5673);
nor U8162 (N_8162,N_4342,N_5047);
nand U8163 (N_8163,N_3492,N_5988);
xor U8164 (N_8164,N_5073,N_3303);
nand U8165 (N_8165,N_3266,N_3653);
nor U8166 (N_8166,N_4773,N_3495);
nor U8167 (N_8167,N_4816,N_5432);
or U8168 (N_8168,N_5200,N_5940);
and U8169 (N_8169,N_4822,N_3510);
nor U8170 (N_8170,N_3663,N_5068);
nor U8171 (N_8171,N_3634,N_5346);
nor U8172 (N_8172,N_5924,N_5218);
and U8173 (N_8173,N_5512,N_5903);
nor U8174 (N_8174,N_3517,N_5815);
nand U8175 (N_8175,N_4991,N_4452);
and U8176 (N_8176,N_3531,N_4386);
or U8177 (N_8177,N_5751,N_3805);
or U8178 (N_8178,N_3288,N_4519);
and U8179 (N_8179,N_5853,N_6020);
nand U8180 (N_8180,N_5822,N_5900);
xor U8181 (N_8181,N_3913,N_4443);
xor U8182 (N_8182,N_4756,N_4628);
nor U8183 (N_8183,N_6089,N_3756);
nand U8184 (N_8184,N_5493,N_4526);
xnor U8185 (N_8185,N_3442,N_5245);
and U8186 (N_8186,N_6138,N_6035);
xor U8187 (N_8187,N_3364,N_5064);
nand U8188 (N_8188,N_5509,N_3982);
xnor U8189 (N_8189,N_3933,N_4725);
nand U8190 (N_8190,N_6217,N_5083);
xor U8191 (N_8191,N_4993,N_5625);
nor U8192 (N_8192,N_5583,N_5495);
nand U8193 (N_8193,N_4747,N_3760);
nand U8194 (N_8194,N_5893,N_3852);
nor U8195 (N_8195,N_3514,N_5222);
nor U8196 (N_8196,N_5899,N_3888);
nor U8197 (N_8197,N_5135,N_4174);
nand U8198 (N_8198,N_4023,N_5736);
and U8199 (N_8199,N_6177,N_5750);
or U8200 (N_8200,N_6064,N_5583);
or U8201 (N_8201,N_4344,N_4895);
and U8202 (N_8202,N_4078,N_4127);
or U8203 (N_8203,N_3468,N_4865);
xnor U8204 (N_8204,N_3648,N_5643);
xor U8205 (N_8205,N_4145,N_5943);
nor U8206 (N_8206,N_3275,N_4666);
nand U8207 (N_8207,N_3477,N_5087);
nand U8208 (N_8208,N_5026,N_3229);
nor U8209 (N_8209,N_3617,N_3299);
nand U8210 (N_8210,N_5836,N_5453);
nor U8211 (N_8211,N_3404,N_3416);
and U8212 (N_8212,N_6116,N_4013);
nand U8213 (N_8213,N_3588,N_4318);
and U8214 (N_8214,N_4753,N_4761);
nor U8215 (N_8215,N_4646,N_4215);
xor U8216 (N_8216,N_4372,N_4672);
or U8217 (N_8217,N_3409,N_4700);
xnor U8218 (N_8218,N_5696,N_5024);
and U8219 (N_8219,N_6117,N_6013);
nor U8220 (N_8220,N_3444,N_5347);
or U8221 (N_8221,N_5147,N_5371);
nor U8222 (N_8222,N_5099,N_6049);
nand U8223 (N_8223,N_5357,N_4417);
and U8224 (N_8224,N_4031,N_3308);
nor U8225 (N_8225,N_4236,N_4196);
or U8226 (N_8226,N_5010,N_5857);
and U8227 (N_8227,N_5801,N_4654);
xor U8228 (N_8228,N_5041,N_5445);
nor U8229 (N_8229,N_5801,N_6126);
and U8230 (N_8230,N_3297,N_3676);
and U8231 (N_8231,N_5710,N_3874);
xnor U8232 (N_8232,N_3207,N_6163);
xor U8233 (N_8233,N_5792,N_3268);
or U8234 (N_8234,N_4558,N_4050);
or U8235 (N_8235,N_5545,N_6205);
or U8236 (N_8236,N_3990,N_4384);
and U8237 (N_8237,N_5878,N_4565);
nor U8238 (N_8238,N_4836,N_3935);
or U8239 (N_8239,N_5231,N_6212);
or U8240 (N_8240,N_5386,N_3925);
xor U8241 (N_8241,N_3403,N_5750);
nor U8242 (N_8242,N_5181,N_5038);
xor U8243 (N_8243,N_3846,N_5142);
nor U8244 (N_8244,N_5480,N_3293);
or U8245 (N_8245,N_3435,N_5720);
or U8246 (N_8246,N_4258,N_5880);
xor U8247 (N_8247,N_3750,N_3260);
nand U8248 (N_8248,N_4609,N_5737);
or U8249 (N_8249,N_3814,N_3324);
and U8250 (N_8250,N_6043,N_5490);
nand U8251 (N_8251,N_5090,N_4041);
nand U8252 (N_8252,N_5374,N_5611);
nor U8253 (N_8253,N_4756,N_5378);
nor U8254 (N_8254,N_4573,N_5821);
nand U8255 (N_8255,N_5952,N_4473);
and U8256 (N_8256,N_5735,N_3188);
xnor U8257 (N_8257,N_3390,N_4099);
xnor U8258 (N_8258,N_4474,N_4630);
nand U8259 (N_8259,N_4797,N_5230);
xor U8260 (N_8260,N_4718,N_5982);
nor U8261 (N_8261,N_5780,N_4308);
or U8262 (N_8262,N_4657,N_5811);
nor U8263 (N_8263,N_5083,N_5122);
xor U8264 (N_8264,N_4947,N_5937);
and U8265 (N_8265,N_6096,N_4606);
or U8266 (N_8266,N_3663,N_4821);
or U8267 (N_8267,N_4055,N_5031);
and U8268 (N_8268,N_3337,N_5351);
or U8269 (N_8269,N_3132,N_3242);
nand U8270 (N_8270,N_3491,N_6240);
nor U8271 (N_8271,N_5538,N_3138);
nor U8272 (N_8272,N_3698,N_5577);
or U8273 (N_8273,N_6196,N_5549);
or U8274 (N_8274,N_4651,N_4481);
and U8275 (N_8275,N_6024,N_6167);
nand U8276 (N_8276,N_6191,N_4154);
or U8277 (N_8277,N_4291,N_3723);
nand U8278 (N_8278,N_3777,N_6070);
nand U8279 (N_8279,N_6102,N_4067);
xnor U8280 (N_8280,N_6043,N_4311);
or U8281 (N_8281,N_4328,N_3738);
or U8282 (N_8282,N_6199,N_5871);
xor U8283 (N_8283,N_4600,N_4113);
or U8284 (N_8284,N_5793,N_5150);
and U8285 (N_8285,N_5698,N_4133);
xor U8286 (N_8286,N_4164,N_4057);
xnor U8287 (N_8287,N_4895,N_5624);
and U8288 (N_8288,N_5337,N_5853);
and U8289 (N_8289,N_4308,N_4221);
or U8290 (N_8290,N_4432,N_3738);
and U8291 (N_8291,N_4234,N_5189);
nand U8292 (N_8292,N_3856,N_3894);
or U8293 (N_8293,N_5063,N_4807);
or U8294 (N_8294,N_4288,N_3518);
nand U8295 (N_8295,N_3462,N_5614);
nor U8296 (N_8296,N_3283,N_6239);
and U8297 (N_8297,N_5920,N_5762);
and U8298 (N_8298,N_4512,N_3968);
and U8299 (N_8299,N_4541,N_3285);
nor U8300 (N_8300,N_5176,N_3666);
nand U8301 (N_8301,N_4646,N_3489);
nor U8302 (N_8302,N_3960,N_6215);
nand U8303 (N_8303,N_3157,N_3150);
and U8304 (N_8304,N_4000,N_4896);
nor U8305 (N_8305,N_5034,N_5143);
xor U8306 (N_8306,N_5092,N_5048);
nand U8307 (N_8307,N_5527,N_5094);
or U8308 (N_8308,N_4938,N_5883);
xnor U8309 (N_8309,N_5067,N_5924);
nor U8310 (N_8310,N_4024,N_4711);
or U8311 (N_8311,N_5438,N_3404);
or U8312 (N_8312,N_3233,N_5724);
nor U8313 (N_8313,N_6211,N_5037);
nor U8314 (N_8314,N_3195,N_4568);
nand U8315 (N_8315,N_5863,N_5924);
nand U8316 (N_8316,N_5866,N_3164);
or U8317 (N_8317,N_5533,N_4356);
xor U8318 (N_8318,N_5141,N_5211);
or U8319 (N_8319,N_3476,N_4337);
or U8320 (N_8320,N_5170,N_3480);
and U8321 (N_8321,N_3790,N_5570);
and U8322 (N_8322,N_4730,N_4518);
xnor U8323 (N_8323,N_3265,N_5317);
xor U8324 (N_8324,N_4251,N_5396);
or U8325 (N_8325,N_4070,N_4303);
and U8326 (N_8326,N_3506,N_5735);
xor U8327 (N_8327,N_3784,N_3630);
and U8328 (N_8328,N_4293,N_4280);
nor U8329 (N_8329,N_5537,N_6195);
nor U8330 (N_8330,N_6117,N_4253);
or U8331 (N_8331,N_4571,N_4331);
and U8332 (N_8332,N_5475,N_5499);
or U8333 (N_8333,N_5620,N_3659);
or U8334 (N_8334,N_5101,N_5488);
and U8335 (N_8335,N_3340,N_5482);
nand U8336 (N_8336,N_5711,N_3244);
nor U8337 (N_8337,N_5384,N_5326);
and U8338 (N_8338,N_6168,N_3975);
xnor U8339 (N_8339,N_3844,N_4429);
or U8340 (N_8340,N_5298,N_5549);
xnor U8341 (N_8341,N_3690,N_3722);
or U8342 (N_8342,N_3244,N_3929);
nand U8343 (N_8343,N_5910,N_6195);
nand U8344 (N_8344,N_3278,N_3695);
xor U8345 (N_8345,N_6164,N_3327);
xnor U8346 (N_8346,N_3426,N_5202);
nor U8347 (N_8347,N_6088,N_3850);
or U8348 (N_8348,N_4905,N_3863);
nand U8349 (N_8349,N_3163,N_5896);
nor U8350 (N_8350,N_5184,N_3141);
xor U8351 (N_8351,N_4365,N_5796);
and U8352 (N_8352,N_4739,N_4531);
and U8353 (N_8353,N_6030,N_5990);
xnor U8354 (N_8354,N_5925,N_5089);
or U8355 (N_8355,N_4140,N_3432);
nand U8356 (N_8356,N_4436,N_4498);
nor U8357 (N_8357,N_4870,N_5002);
xnor U8358 (N_8358,N_3466,N_3605);
xor U8359 (N_8359,N_3447,N_3424);
nor U8360 (N_8360,N_3524,N_3968);
nor U8361 (N_8361,N_5285,N_3910);
and U8362 (N_8362,N_5936,N_5809);
and U8363 (N_8363,N_4153,N_5804);
xor U8364 (N_8364,N_5148,N_4772);
xor U8365 (N_8365,N_4995,N_5690);
nor U8366 (N_8366,N_3950,N_4788);
xnor U8367 (N_8367,N_3459,N_5871);
xnor U8368 (N_8368,N_5481,N_4327);
and U8369 (N_8369,N_6062,N_5125);
and U8370 (N_8370,N_4192,N_5979);
nor U8371 (N_8371,N_4069,N_4464);
nand U8372 (N_8372,N_4958,N_3965);
or U8373 (N_8373,N_5741,N_3959);
or U8374 (N_8374,N_4145,N_5399);
and U8375 (N_8375,N_5662,N_3854);
nor U8376 (N_8376,N_4810,N_4055);
nand U8377 (N_8377,N_3323,N_3840);
nand U8378 (N_8378,N_5388,N_3952);
and U8379 (N_8379,N_4807,N_4833);
nor U8380 (N_8380,N_4185,N_3844);
xnor U8381 (N_8381,N_4236,N_4869);
and U8382 (N_8382,N_3958,N_5707);
nand U8383 (N_8383,N_5713,N_5931);
nor U8384 (N_8384,N_3918,N_4478);
nor U8385 (N_8385,N_6100,N_5344);
nor U8386 (N_8386,N_5079,N_3553);
or U8387 (N_8387,N_5060,N_6197);
nand U8388 (N_8388,N_3925,N_3131);
and U8389 (N_8389,N_3714,N_5413);
nor U8390 (N_8390,N_3370,N_4575);
or U8391 (N_8391,N_3518,N_4417);
and U8392 (N_8392,N_4357,N_3487);
and U8393 (N_8393,N_5485,N_5612);
and U8394 (N_8394,N_6096,N_3173);
or U8395 (N_8395,N_3515,N_3411);
nor U8396 (N_8396,N_5849,N_5876);
and U8397 (N_8397,N_3590,N_5623);
and U8398 (N_8398,N_3906,N_3681);
nor U8399 (N_8399,N_5498,N_5558);
xnor U8400 (N_8400,N_5061,N_5869);
nor U8401 (N_8401,N_5170,N_5368);
or U8402 (N_8402,N_4701,N_3150);
and U8403 (N_8403,N_4048,N_3360);
and U8404 (N_8404,N_3819,N_5624);
or U8405 (N_8405,N_6082,N_3662);
and U8406 (N_8406,N_3218,N_4534);
and U8407 (N_8407,N_5152,N_3618);
nand U8408 (N_8408,N_5909,N_4989);
or U8409 (N_8409,N_4175,N_4062);
nand U8410 (N_8410,N_3729,N_6223);
nand U8411 (N_8411,N_5694,N_5093);
nand U8412 (N_8412,N_3268,N_3169);
nor U8413 (N_8413,N_4054,N_4536);
nand U8414 (N_8414,N_5811,N_4270);
and U8415 (N_8415,N_3354,N_5172);
nand U8416 (N_8416,N_5178,N_4182);
nand U8417 (N_8417,N_3156,N_4295);
or U8418 (N_8418,N_4667,N_4181);
nor U8419 (N_8419,N_5983,N_4697);
xor U8420 (N_8420,N_4204,N_5871);
or U8421 (N_8421,N_5419,N_4965);
nand U8422 (N_8422,N_3708,N_5256);
or U8423 (N_8423,N_6044,N_4108);
nor U8424 (N_8424,N_5597,N_5497);
xnor U8425 (N_8425,N_4442,N_5617);
or U8426 (N_8426,N_4052,N_5272);
nand U8427 (N_8427,N_3185,N_4759);
xor U8428 (N_8428,N_6051,N_4749);
and U8429 (N_8429,N_3579,N_6082);
nand U8430 (N_8430,N_3219,N_3769);
or U8431 (N_8431,N_5856,N_4627);
and U8432 (N_8432,N_3685,N_5680);
nand U8433 (N_8433,N_5649,N_3768);
and U8434 (N_8434,N_5128,N_5066);
xor U8435 (N_8435,N_5386,N_4987);
and U8436 (N_8436,N_3453,N_4780);
and U8437 (N_8437,N_5072,N_5875);
and U8438 (N_8438,N_3217,N_4561);
nor U8439 (N_8439,N_6166,N_3386);
or U8440 (N_8440,N_3828,N_5022);
nor U8441 (N_8441,N_5847,N_5568);
and U8442 (N_8442,N_6164,N_3133);
or U8443 (N_8443,N_5002,N_4778);
nor U8444 (N_8444,N_5878,N_4475);
nand U8445 (N_8445,N_5059,N_6205);
nor U8446 (N_8446,N_3906,N_5290);
and U8447 (N_8447,N_4729,N_4470);
or U8448 (N_8448,N_4642,N_3358);
or U8449 (N_8449,N_4832,N_4385);
nor U8450 (N_8450,N_6003,N_4993);
nand U8451 (N_8451,N_3192,N_3198);
nand U8452 (N_8452,N_3670,N_5822);
and U8453 (N_8453,N_3291,N_5461);
and U8454 (N_8454,N_4591,N_4128);
or U8455 (N_8455,N_4340,N_4033);
nor U8456 (N_8456,N_4298,N_5140);
nand U8457 (N_8457,N_5289,N_3381);
or U8458 (N_8458,N_3586,N_4241);
xnor U8459 (N_8459,N_5256,N_6078);
and U8460 (N_8460,N_3530,N_3588);
or U8461 (N_8461,N_4283,N_4473);
xor U8462 (N_8462,N_3630,N_3351);
and U8463 (N_8463,N_3919,N_4842);
and U8464 (N_8464,N_5133,N_3649);
nand U8465 (N_8465,N_5948,N_4579);
xor U8466 (N_8466,N_4079,N_3553);
or U8467 (N_8467,N_4530,N_5459);
nand U8468 (N_8468,N_5854,N_4986);
xnor U8469 (N_8469,N_6211,N_3497);
and U8470 (N_8470,N_4504,N_5015);
nand U8471 (N_8471,N_4811,N_3485);
nor U8472 (N_8472,N_4789,N_5319);
nor U8473 (N_8473,N_4071,N_3538);
or U8474 (N_8474,N_6096,N_3932);
and U8475 (N_8475,N_5547,N_4134);
nand U8476 (N_8476,N_4855,N_4249);
nor U8477 (N_8477,N_4902,N_3476);
nor U8478 (N_8478,N_5005,N_4180);
or U8479 (N_8479,N_6104,N_5486);
nor U8480 (N_8480,N_5142,N_5475);
or U8481 (N_8481,N_5754,N_6024);
xnor U8482 (N_8482,N_3520,N_4178);
xor U8483 (N_8483,N_4354,N_5808);
or U8484 (N_8484,N_5511,N_6181);
nand U8485 (N_8485,N_5396,N_5037);
nor U8486 (N_8486,N_3578,N_4469);
xor U8487 (N_8487,N_5442,N_3184);
xnor U8488 (N_8488,N_3447,N_3857);
nand U8489 (N_8489,N_5198,N_3243);
nand U8490 (N_8490,N_4039,N_6067);
nor U8491 (N_8491,N_5264,N_3186);
and U8492 (N_8492,N_4257,N_4184);
nand U8493 (N_8493,N_6004,N_5447);
nand U8494 (N_8494,N_5260,N_5487);
xnor U8495 (N_8495,N_5557,N_4427);
xor U8496 (N_8496,N_5467,N_5786);
or U8497 (N_8497,N_3207,N_5899);
nor U8498 (N_8498,N_3740,N_5277);
nand U8499 (N_8499,N_5788,N_4474);
xor U8500 (N_8500,N_5389,N_3939);
xnor U8501 (N_8501,N_5298,N_3687);
nor U8502 (N_8502,N_5880,N_4675);
nor U8503 (N_8503,N_4527,N_4150);
or U8504 (N_8504,N_5395,N_3202);
xor U8505 (N_8505,N_4811,N_3793);
nor U8506 (N_8506,N_3566,N_4077);
xor U8507 (N_8507,N_5565,N_6215);
nor U8508 (N_8508,N_4565,N_3653);
nand U8509 (N_8509,N_6034,N_6007);
nand U8510 (N_8510,N_6017,N_3366);
nand U8511 (N_8511,N_5726,N_4517);
xor U8512 (N_8512,N_3781,N_5782);
xnor U8513 (N_8513,N_4016,N_5951);
nor U8514 (N_8514,N_5113,N_4199);
xor U8515 (N_8515,N_3935,N_3516);
nand U8516 (N_8516,N_5203,N_5513);
xor U8517 (N_8517,N_3834,N_3682);
xor U8518 (N_8518,N_3391,N_5230);
nor U8519 (N_8519,N_4936,N_3838);
and U8520 (N_8520,N_5739,N_3146);
nor U8521 (N_8521,N_4384,N_5363);
nor U8522 (N_8522,N_5299,N_5480);
nand U8523 (N_8523,N_6046,N_4418);
or U8524 (N_8524,N_5397,N_5931);
nand U8525 (N_8525,N_3459,N_5677);
xor U8526 (N_8526,N_3801,N_5837);
nor U8527 (N_8527,N_4867,N_4570);
nor U8528 (N_8528,N_6104,N_3147);
and U8529 (N_8529,N_3338,N_5637);
or U8530 (N_8530,N_4780,N_3801);
xor U8531 (N_8531,N_3588,N_4385);
and U8532 (N_8532,N_6017,N_3960);
xor U8533 (N_8533,N_5082,N_3792);
xor U8534 (N_8534,N_3257,N_5367);
nor U8535 (N_8535,N_3949,N_4907);
and U8536 (N_8536,N_5588,N_4677);
and U8537 (N_8537,N_3682,N_6249);
or U8538 (N_8538,N_4363,N_4235);
or U8539 (N_8539,N_4102,N_3765);
or U8540 (N_8540,N_3520,N_3780);
or U8541 (N_8541,N_5594,N_4063);
nand U8542 (N_8542,N_3172,N_3237);
nor U8543 (N_8543,N_4472,N_3279);
xnor U8544 (N_8544,N_4120,N_4162);
nor U8545 (N_8545,N_5946,N_4735);
nor U8546 (N_8546,N_5002,N_5564);
nand U8547 (N_8547,N_5606,N_3915);
xor U8548 (N_8548,N_4976,N_3222);
nor U8549 (N_8549,N_4763,N_4307);
or U8550 (N_8550,N_3155,N_5533);
xor U8551 (N_8551,N_4915,N_3464);
or U8552 (N_8552,N_5181,N_3722);
nor U8553 (N_8553,N_4447,N_6087);
nor U8554 (N_8554,N_3431,N_4439);
or U8555 (N_8555,N_4579,N_3534);
or U8556 (N_8556,N_4619,N_3554);
and U8557 (N_8557,N_3613,N_5623);
or U8558 (N_8558,N_4589,N_4211);
or U8559 (N_8559,N_4641,N_5600);
or U8560 (N_8560,N_3663,N_5324);
nand U8561 (N_8561,N_6184,N_3377);
xnor U8562 (N_8562,N_5325,N_5419);
or U8563 (N_8563,N_5011,N_4971);
xnor U8564 (N_8564,N_4126,N_4673);
or U8565 (N_8565,N_5603,N_3332);
or U8566 (N_8566,N_3222,N_5736);
nand U8567 (N_8567,N_5222,N_4814);
and U8568 (N_8568,N_5074,N_5629);
nor U8569 (N_8569,N_4133,N_4100);
xnor U8570 (N_8570,N_3405,N_6226);
xnor U8571 (N_8571,N_5622,N_5432);
nor U8572 (N_8572,N_3990,N_6005);
and U8573 (N_8573,N_6121,N_5106);
and U8574 (N_8574,N_3868,N_4115);
xor U8575 (N_8575,N_3460,N_5944);
nand U8576 (N_8576,N_3521,N_3501);
nand U8577 (N_8577,N_3343,N_4131);
or U8578 (N_8578,N_3202,N_4235);
or U8579 (N_8579,N_5972,N_3912);
or U8580 (N_8580,N_5381,N_5602);
and U8581 (N_8581,N_3666,N_4107);
nand U8582 (N_8582,N_5646,N_5165);
or U8583 (N_8583,N_3585,N_4896);
nand U8584 (N_8584,N_4518,N_4111);
nand U8585 (N_8585,N_3881,N_5820);
and U8586 (N_8586,N_5588,N_3471);
or U8587 (N_8587,N_5185,N_5601);
and U8588 (N_8588,N_4918,N_6051);
nand U8589 (N_8589,N_4852,N_5448);
xnor U8590 (N_8590,N_3922,N_4320);
nand U8591 (N_8591,N_4880,N_4273);
nor U8592 (N_8592,N_5886,N_5392);
nand U8593 (N_8593,N_5911,N_3164);
or U8594 (N_8594,N_4568,N_4957);
or U8595 (N_8595,N_4938,N_3895);
nor U8596 (N_8596,N_4218,N_3231);
nor U8597 (N_8597,N_3293,N_5277);
nor U8598 (N_8598,N_6040,N_3377);
and U8599 (N_8599,N_3719,N_5018);
xnor U8600 (N_8600,N_5367,N_4411);
xnor U8601 (N_8601,N_4304,N_6004);
xnor U8602 (N_8602,N_3602,N_5045);
nor U8603 (N_8603,N_4172,N_3409);
xor U8604 (N_8604,N_5065,N_4881);
xnor U8605 (N_8605,N_3711,N_5461);
and U8606 (N_8606,N_3663,N_3474);
xnor U8607 (N_8607,N_5616,N_4797);
and U8608 (N_8608,N_3866,N_4580);
nor U8609 (N_8609,N_4630,N_4482);
and U8610 (N_8610,N_4208,N_5410);
and U8611 (N_8611,N_4412,N_6019);
and U8612 (N_8612,N_4185,N_4256);
or U8613 (N_8613,N_5315,N_3519);
nand U8614 (N_8614,N_4099,N_5552);
or U8615 (N_8615,N_4246,N_5146);
nor U8616 (N_8616,N_5289,N_3781);
nand U8617 (N_8617,N_3198,N_4304);
and U8618 (N_8618,N_4700,N_4302);
xor U8619 (N_8619,N_3996,N_4097);
nor U8620 (N_8620,N_4472,N_4554);
and U8621 (N_8621,N_5463,N_3286);
xor U8622 (N_8622,N_5753,N_3921);
xor U8623 (N_8623,N_4056,N_4259);
nor U8624 (N_8624,N_6149,N_6010);
nor U8625 (N_8625,N_3224,N_3600);
or U8626 (N_8626,N_4399,N_4360);
and U8627 (N_8627,N_3919,N_5529);
nor U8628 (N_8628,N_3364,N_3469);
nand U8629 (N_8629,N_5896,N_5840);
or U8630 (N_8630,N_6093,N_3220);
nor U8631 (N_8631,N_3951,N_4443);
xnor U8632 (N_8632,N_5728,N_3536);
xnor U8633 (N_8633,N_4433,N_4835);
and U8634 (N_8634,N_3326,N_4811);
nand U8635 (N_8635,N_3747,N_4256);
nand U8636 (N_8636,N_5934,N_3861);
nand U8637 (N_8637,N_5445,N_3457);
xor U8638 (N_8638,N_3318,N_4120);
or U8639 (N_8639,N_3308,N_5333);
xor U8640 (N_8640,N_4591,N_3318);
nand U8641 (N_8641,N_5319,N_4172);
nor U8642 (N_8642,N_5825,N_4601);
and U8643 (N_8643,N_3191,N_5810);
nand U8644 (N_8644,N_3370,N_4363);
and U8645 (N_8645,N_5753,N_4632);
nand U8646 (N_8646,N_3602,N_5337);
nor U8647 (N_8647,N_3934,N_3440);
and U8648 (N_8648,N_5389,N_5340);
or U8649 (N_8649,N_5608,N_5282);
and U8650 (N_8650,N_4694,N_3280);
or U8651 (N_8651,N_6160,N_5767);
nor U8652 (N_8652,N_5882,N_4428);
and U8653 (N_8653,N_5010,N_3672);
nand U8654 (N_8654,N_3442,N_4128);
nand U8655 (N_8655,N_6069,N_5308);
xor U8656 (N_8656,N_4805,N_4347);
or U8657 (N_8657,N_3207,N_3601);
xor U8658 (N_8658,N_4856,N_4848);
or U8659 (N_8659,N_5810,N_4669);
nand U8660 (N_8660,N_5605,N_3875);
xor U8661 (N_8661,N_4091,N_4904);
nor U8662 (N_8662,N_4823,N_5253);
nand U8663 (N_8663,N_5278,N_4276);
and U8664 (N_8664,N_4009,N_5573);
nor U8665 (N_8665,N_6074,N_4194);
or U8666 (N_8666,N_6024,N_4944);
or U8667 (N_8667,N_4852,N_5110);
or U8668 (N_8668,N_6215,N_4023);
or U8669 (N_8669,N_3715,N_5805);
and U8670 (N_8670,N_4462,N_3954);
nand U8671 (N_8671,N_5589,N_5778);
and U8672 (N_8672,N_3510,N_3152);
nand U8673 (N_8673,N_3397,N_4339);
nand U8674 (N_8674,N_3918,N_4581);
or U8675 (N_8675,N_3400,N_5174);
nand U8676 (N_8676,N_6123,N_4903);
or U8677 (N_8677,N_5010,N_4189);
xnor U8678 (N_8678,N_4217,N_4043);
nand U8679 (N_8679,N_5035,N_4291);
and U8680 (N_8680,N_5252,N_5296);
or U8681 (N_8681,N_5552,N_5570);
or U8682 (N_8682,N_4683,N_3715);
xnor U8683 (N_8683,N_5624,N_4606);
nand U8684 (N_8684,N_5544,N_6052);
nor U8685 (N_8685,N_4008,N_4767);
xnor U8686 (N_8686,N_5508,N_4114);
or U8687 (N_8687,N_4457,N_4198);
xor U8688 (N_8688,N_5837,N_4707);
and U8689 (N_8689,N_4249,N_5593);
xor U8690 (N_8690,N_4376,N_4157);
nand U8691 (N_8691,N_3626,N_3991);
and U8692 (N_8692,N_4328,N_4343);
or U8693 (N_8693,N_4095,N_4856);
or U8694 (N_8694,N_3567,N_3655);
or U8695 (N_8695,N_4651,N_5360);
or U8696 (N_8696,N_3306,N_3201);
nand U8697 (N_8697,N_5809,N_4057);
nand U8698 (N_8698,N_3591,N_5687);
nand U8699 (N_8699,N_5162,N_3928);
xor U8700 (N_8700,N_4714,N_3949);
nand U8701 (N_8701,N_5593,N_5077);
nor U8702 (N_8702,N_3429,N_4764);
and U8703 (N_8703,N_3438,N_3824);
or U8704 (N_8704,N_4751,N_4349);
and U8705 (N_8705,N_5768,N_3651);
and U8706 (N_8706,N_5319,N_5523);
xor U8707 (N_8707,N_4914,N_5987);
xor U8708 (N_8708,N_3272,N_4633);
nor U8709 (N_8709,N_4573,N_4818);
and U8710 (N_8710,N_4492,N_4290);
xnor U8711 (N_8711,N_5347,N_3813);
and U8712 (N_8712,N_5540,N_3372);
nand U8713 (N_8713,N_5708,N_3502);
nor U8714 (N_8714,N_4915,N_6150);
or U8715 (N_8715,N_5308,N_5746);
or U8716 (N_8716,N_4126,N_3996);
nor U8717 (N_8717,N_5958,N_3526);
xnor U8718 (N_8718,N_4747,N_4211);
or U8719 (N_8719,N_3377,N_3816);
and U8720 (N_8720,N_5324,N_5362);
xor U8721 (N_8721,N_3762,N_3229);
nor U8722 (N_8722,N_5500,N_3635);
xor U8723 (N_8723,N_3619,N_5897);
or U8724 (N_8724,N_5497,N_3581);
nor U8725 (N_8725,N_4778,N_4020);
nand U8726 (N_8726,N_4093,N_3217);
xnor U8727 (N_8727,N_5213,N_4671);
or U8728 (N_8728,N_4375,N_4502);
nand U8729 (N_8729,N_3704,N_4896);
or U8730 (N_8730,N_5222,N_5028);
nor U8731 (N_8731,N_6116,N_6169);
and U8732 (N_8732,N_3487,N_6223);
nand U8733 (N_8733,N_5258,N_3450);
and U8734 (N_8734,N_4135,N_4502);
xnor U8735 (N_8735,N_4290,N_5061);
xnor U8736 (N_8736,N_5197,N_3614);
nand U8737 (N_8737,N_6218,N_6210);
nor U8738 (N_8738,N_5067,N_4885);
and U8739 (N_8739,N_5040,N_5250);
nor U8740 (N_8740,N_4976,N_4975);
and U8741 (N_8741,N_4741,N_3769);
nor U8742 (N_8742,N_5094,N_5771);
xnor U8743 (N_8743,N_5886,N_5193);
and U8744 (N_8744,N_6112,N_4768);
and U8745 (N_8745,N_3462,N_3664);
or U8746 (N_8746,N_3327,N_4720);
and U8747 (N_8747,N_5744,N_5641);
nor U8748 (N_8748,N_3964,N_5372);
or U8749 (N_8749,N_4339,N_4517);
nor U8750 (N_8750,N_4604,N_5706);
or U8751 (N_8751,N_4840,N_6116);
nor U8752 (N_8752,N_3799,N_5278);
xor U8753 (N_8753,N_3158,N_6019);
xor U8754 (N_8754,N_4243,N_4273);
and U8755 (N_8755,N_3986,N_4172);
nor U8756 (N_8756,N_4181,N_5686);
nand U8757 (N_8757,N_4253,N_5243);
nor U8758 (N_8758,N_4010,N_5937);
nor U8759 (N_8759,N_4627,N_3701);
nor U8760 (N_8760,N_5803,N_3137);
nand U8761 (N_8761,N_6068,N_4344);
and U8762 (N_8762,N_5026,N_6012);
or U8763 (N_8763,N_4835,N_3972);
or U8764 (N_8764,N_4671,N_3202);
and U8765 (N_8765,N_4331,N_5030);
nor U8766 (N_8766,N_5023,N_4819);
and U8767 (N_8767,N_6009,N_6203);
nor U8768 (N_8768,N_3489,N_4109);
and U8769 (N_8769,N_4411,N_3433);
nor U8770 (N_8770,N_4006,N_4984);
nor U8771 (N_8771,N_5183,N_4451);
nand U8772 (N_8772,N_5015,N_4273);
or U8773 (N_8773,N_4035,N_5947);
and U8774 (N_8774,N_5965,N_4051);
and U8775 (N_8775,N_5632,N_4919);
nand U8776 (N_8776,N_5123,N_5980);
xnor U8777 (N_8777,N_3530,N_3487);
or U8778 (N_8778,N_3659,N_4167);
and U8779 (N_8779,N_4711,N_5632);
nor U8780 (N_8780,N_3173,N_4443);
nand U8781 (N_8781,N_4001,N_5999);
nand U8782 (N_8782,N_6182,N_3408);
and U8783 (N_8783,N_4987,N_5875);
nor U8784 (N_8784,N_6183,N_4664);
and U8785 (N_8785,N_4551,N_4391);
and U8786 (N_8786,N_4836,N_4359);
nand U8787 (N_8787,N_6169,N_3926);
and U8788 (N_8788,N_5863,N_4093);
xor U8789 (N_8789,N_4675,N_3404);
xnor U8790 (N_8790,N_5625,N_5343);
and U8791 (N_8791,N_6042,N_5431);
and U8792 (N_8792,N_3780,N_3988);
or U8793 (N_8793,N_5867,N_5265);
xnor U8794 (N_8794,N_5150,N_3682);
xor U8795 (N_8795,N_5364,N_3786);
or U8796 (N_8796,N_5899,N_3694);
nand U8797 (N_8797,N_3233,N_4136);
nor U8798 (N_8798,N_4902,N_5024);
xnor U8799 (N_8799,N_4349,N_3937);
or U8800 (N_8800,N_4252,N_4376);
nand U8801 (N_8801,N_3626,N_5809);
nand U8802 (N_8802,N_5592,N_5629);
and U8803 (N_8803,N_5925,N_5172);
xor U8804 (N_8804,N_5270,N_5596);
xor U8805 (N_8805,N_5753,N_6163);
nand U8806 (N_8806,N_5415,N_4676);
xor U8807 (N_8807,N_4861,N_6014);
or U8808 (N_8808,N_6045,N_5815);
xnor U8809 (N_8809,N_4291,N_4683);
xor U8810 (N_8810,N_3884,N_4109);
or U8811 (N_8811,N_3616,N_5645);
or U8812 (N_8812,N_4387,N_6100);
or U8813 (N_8813,N_5296,N_5544);
nor U8814 (N_8814,N_4059,N_3856);
nor U8815 (N_8815,N_4067,N_3444);
or U8816 (N_8816,N_4669,N_4113);
xnor U8817 (N_8817,N_3704,N_3769);
and U8818 (N_8818,N_5351,N_4176);
nor U8819 (N_8819,N_6181,N_3194);
nor U8820 (N_8820,N_4418,N_3280);
nand U8821 (N_8821,N_5798,N_3511);
nand U8822 (N_8822,N_6054,N_3823);
or U8823 (N_8823,N_4277,N_4982);
nand U8824 (N_8824,N_5979,N_5230);
nand U8825 (N_8825,N_6192,N_6164);
xnor U8826 (N_8826,N_5630,N_6165);
or U8827 (N_8827,N_4317,N_5429);
and U8828 (N_8828,N_5053,N_4934);
nand U8829 (N_8829,N_4131,N_6234);
or U8830 (N_8830,N_6015,N_3624);
nor U8831 (N_8831,N_4604,N_5772);
xnor U8832 (N_8832,N_5625,N_4683);
and U8833 (N_8833,N_5737,N_5118);
xor U8834 (N_8834,N_3400,N_4950);
nor U8835 (N_8835,N_3967,N_3957);
nor U8836 (N_8836,N_5633,N_5939);
xnor U8837 (N_8837,N_4520,N_6073);
xor U8838 (N_8838,N_4350,N_3624);
nor U8839 (N_8839,N_5810,N_4489);
and U8840 (N_8840,N_3213,N_3822);
or U8841 (N_8841,N_6167,N_5440);
or U8842 (N_8842,N_4474,N_3814);
nand U8843 (N_8843,N_5013,N_3818);
xnor U8844 (N_8844,N_5576,N_5540);
xor U8845 (N_8845,N_5625,N_4287);
nand U8846 (N_8846,N_4088,N_5423);
or U8847 (N_8847,N_5148,N_3658);
nor U8848 (N_8848,N_4750,N_5319);
or U8849 (N_8849,N_5768,N_3154);
xnor U8850 (N_8850,N_3597,N_5388);
nor U8851 (N_8851,N_3228,N_3828);
nand U8852 (N_8852,N_4876,N_5657);
nor U8853 (N_8853,N_4302,N_4558);
nand U8854 (N_8854,N_5094,N_4804);
or U8855 (N_8855,N_5483,N_3900);
nand U8856 (N_8856,N_3442,N_5378);
nor U8857 (N_8857,N_5861,N_4645);
nand U8858 (N_8858,N_3843,N_4417);
and U8859 (N_8859,N_4039,N_5492);
and U8860 (N_8860,N_3896,N_5551);
xnor U8861 (N_8861,N_5581,N_3916);
xnor U8862 (N_8862,N_5827,N_4182);
xor U8863 (N_8863,N_5713,N_4411);
or U8864 (N_8864,N_5602,N_6164);
nand U8865 (N_8865,N_4140,N_4320);
or U8866 (N_8866,N_5159,N_5821);
nand U8867 (N_8867,N_5997,N_5370);
nand U8868 (N_8868,N_4820,N_5786);
xor U8869 (N_8869,N_3602,N_3543);
nand U8870 (N_8870,N_3347,N_4708);
xor U8871 (N_8871,N_5854,N_4434);
xnor U8872 (N_8872,N_5849,N_4050);
and U8873 (N_8873,N_5070,N_4696);
nand U8874 (N_8874,N_5766,N_6033);
nor U8875 (N_8875,N_5381,N_3879);
nand U8876 (N_8876,N_4668,N_5412);
nand U8877 (N_8877,N_3917,N_3832);
xnor U8878 (N_8878,N_4094,N_5181);
or U8879 (N_8879,N_3275,N_5389);
xor U8880 (N_8880,N_4440,N_5246);
nand U8881 (N_8881,N_4887,N_3997);
xor U8882 (N_8882,N_3936,N_4121);
nand U8883 (N_8883,N_3759,N_4123);
nand U8884 (N_8884,N_3719,N_4668);
or U8885 (N_8885,N_4459,N_4534);
nand U8886 (N_8886,N_4373,N_5168);
nand U8887 (N_8887,N_6077,N_3883);
or U8888 (N_8888,N_6191,N_5506);
xor U8889 (N_8889,N_4899,N_5182);
nand U8890 (N_8890,N_4970,N_6019);
and U8891 (N_8891,N_5270,N_4412);
and U8892 (N_8892,N_4024,N_3991);
nor U8893 (N_8893,N_5041,N_4215);
and U8894 (N_8894,N_5355,N_6217);
or U8895 (N_8895,N_4857,N_4469);
and U8896 (N_8896,N_4601,N_5756);
xor U8897 (N_8897,N_3153,N_4424);
nand U8898 (N_8898,N_5131,N_5648);
or U8899 (N_8899,N_3213,N_3150);
nand U8900 (N_8900,N_5459,N_5877);
nor U8901 (N_8901,N_4883,N_3509);
nor U8902 (N_8902,N_5398,N_4689);
nor U8903 (N_8903,N_5490,N_5021);
nor U8904 (N_8904,N_4227,N_3464);
or U8905 (N_8905,N_5022,N_3813);
nand U8906 (N_8906,N_4028,N_3941);
or U8907 (N_8907,N_5379,N_4566);
nor U8908 (N_8908,N_5478,N_5207);
nor U8909 (N_8909,N_4024,N_5283);
nand U8910 (N_8910,N_4251,N_4915);
and U8911 (N_8911,N_4236,N_5356);
and U8912 (N_8912,N_5681,N_6000);
or U8913 (N_8913,N_5769,N_6142);
nor U8914 (N_8914,N_3878,N_5407);
xnor U8915 (N_8915,N_4273,N_6027);
nand U8916 (N_8916,N_3831,N_3357);
xor U8917 (N_8917,N_5332,N_3967);
or U8918 (N_8918,N_6135,N_5000);
and U8919 (N_8919,N_5639,N_4756);
nor U8920 (N_8920,N_4054,N_5648);
nand U8921 (N_8921,N_4748,N_5198);
and U8922 (N_8922,N_5048,N_3472);
xor U8923 (N_8923,N_5344,N_4588);
and U8924 (N_8924,N_5160,N_4911);
nor U8925 (N_8925,N_5108,N_4686);
xnor U8926 (N_8926,N_4231,N_5000);
xnor U8927 (N_8927,N_3569,N_3183);
nor U8928 (N_8928,N_6245,N_3588);
and U8929 (N_8929,N_4419,N_4146);
nor U8930 (N_8930,N_4106,N_4809);
and U8931 (N_8931,N_3977,N_5271);
and U8932 (N_8932,N_5860,N_5593);
nor U8933 (N_8933,N_5527,N_5148);
nand U8934 (N_8934,N_4932,N_4219);
or U8935 (N_8935,N_5089,N_4815);
nor U8936 (N_8936,N_5256,N_4365);
nor U8937 (N_8937,N_6124,N_3716);
nor U8938 (N_8938,N_5004,N_4277);
and U8939 (N_8939,N_5968,N_3927);
and U8940 (N_8940,N_4496,N_5901);
and U8941 (N_8941,N_3841,N_4954);
or U8942 (N_8942,N_3391,N_6156);
xor U8943 (N_8943,N_4716,N_4900);
or U8944 (N_8944,N_6144,N_3354);
xor U8945 (N_8945,N_5992,N_4506);
and U8946 (N_8946,N_4323,N_3646);
nor U8947 (N_8947,N_5599,N_3838);
and U8948 (N_8948,N_4779,N_6028);
nor U8949 (N_8949,N_6230,N_6048);
or U8950 (N_8950,N_3936,N_4560);
and U8951 (N_8951,N_5571,N_5991);
or U8952 (N_8952,N_5292,N_4667);
nand U8953 (N_8953,N_3333,N_3293);
or U8954 (N_8954,N_3721,N_4477);
or U8955 (N_8955,N_3261,N_4364);
xnor U8956 (N_8956,N_4875,N_5961);
nand U8957 (N_8957,N_4879,N_4461);
xor U8958 (N_8958,N_4767,N_4353);
nand U8959 (N_8959,N_5339,N_5536);
nand U8960 (N_8960,N_3395,N_6012);
and U8961 (N_8961,N_4273,N_4513);
nand U8962 (N_8962,N_5314,N_5860);
and U8963 (N_8963,N_5707,N_3842);
xor U8964 (N_8964,N_3290,N_6061);
nor U8965 (N_8965,N_5779,N_4193);
and U8966 (N_8966,N_3474,N_3551);
or U8967 (N_8967,N_5733,N_6011);
and U8968 (N_8968,N_4752,N_4469);
nor U8969 (N_8969,N_4484,N_6197);
or U8970 (N_8970,N_3352,N_4343);
nor U8971 (N_8971,N_4556,N_4333);
nand U8972 (N_8972,N_5128,N_3230);
nand U8973 (N_8973,N_5095,N_5111);
nor U8974 (N_8974,N_5129,N_5993);
xor U8975 (N_8975,N_3267,N_5035);
or U8976 (N_8976,N_5303,N_4829);
xor U8977 (N_8977,N_4696,N_5960);
or U8978 (N_8978,N_4085,N_5290);
or U8979 (N_8979,N_5381,N_5902);
or U8980 (N_8980,N_6050,N_4858);
nor U8981 (N_8981,N_4251,N_5520);
and U8982 (N_8982,N_3605,N_6135);
and U8983 (N_8983,N_5580,N_4346);
nand U8984 (N_8984,N_4549,N_6205);
or U8985 (N_8985,N_3807,N_4044);
nor U8986 (N_8986,N_6015,N_3404);
and U8987 (N_8987,N_4459,N_5067);
or U8988 (N_8988,N_5768,N_4229);
xnor U8989 (N_8989,N_5229,N_3622);
nor U8990 (N_8990,N_5269,N_3558);
xnor U8991 (N_8991,N_3230,N_6249);
and U8992 (N_8992,N_5438,N_3445);
nand U8993 (N_8993,N_4318,N_4928);
nand U8994 (N_8994,N_3935,N_5273);
nand U8995 (N_8995,N_3437,N_4599);
or U8996 (N_8996,N_4969,N_5414);
xor U8997 (N_8997,N_5714,N_6232);
nor U8998 (N_8998,N_4101,N_6121);
nand U8999 (N_8999,N_3516,N_3898);
nor U9000 (N_9000,N_5760,N_3128);
or U9001 (N_9001,N_6241,N_4366);
nand U9002 (N_9002,N_3475,N_5868);
nor U9003 (N_9003,N_4548,N_3715);
or U9004 (N_9004,N_4165,N_4117);
or U9005 (N_9005,N_5573,N_5698);
nand U9006 (N_9006,N_5585,N_5573);
xnor U9007 (N_9007,N_4302,N_4980);
nor U9008 (N_9008,N_5487,N_6219);
xnor U9009 (N_9009,N_4383,N_3370);
xnor U9010 (N_9010,N_4420,N_5419);
or U9011 (N_9011,N_6170,N_4547);
nor U9012 (N_9012,N_4188,N_5637);
nand U9013 (N_9013,N_5140,N_4446);
and U9014 (N_9014,N_4569,N_3150);
or U9015 (N_9015,N_5796,N_3674);
nor U9016 (N_9016,N_3448,N_3815);
or U9017 (N_9017,N_6081,N_5235);
or U9018 (N_9018,N_5029,N_4985);
nand U9019 (N_9019,N_5417,N_4684);
nor U9020 (N_9020,N_3232,N_3352);
and U9021 (N_9021,N_3291,N_5025);
or U9022 (N_9022,N_3988,N_5254);
nand U9023 (N_9023,N_3329,N_5743);
and U9024 (N_9024,N_4358,N_4366);
nand U9025 (N_9025,N_5776,N_4141);
nand U9026 (N_9026,N_5627,N_3597);
xor U9027 (N_9027,N_4558,N_5433);
and U9028 (N_9028,N_5830,N_6072);
nand U9029 (N_9029,N_5883,N_4116);
and U9030 (N_9030,N_5761,N_5400);
and U9031 (N_9031,N_3840,N_3222);
and U9032 (N_9032,N_4291,N_3918);
or U9033 (N_9033,N_3466,N_3435);
and U9034 (N_9034,N_5997,N_3687);
and U9035 (N_9035,N_5621,N_3908);
nor U9036 (N_9036,N_3394,N_4046);
nand U9037 (N_9037,N_3186,N_3146);
and U9038 (N_9038,N_4541,N_5561);
nor U9039 (N_9039,N_5748,N_4745);
and U9040 (N_9040,N_6220,N_3248);
and U9041 (N_9041,N_5825,N_3167);
or U9042 (N_9042,N_6054,N_3585);
nor U9043 (N_9043,N_4870,N_6005);
nand U9044 (N_9044,N_5868,N_3768);
nand U9045 (N_9045,N_3359,N_4051);
and U9046 (N_9046,N_4856,N_4134);
or U9047 (N_9047,N_5770,N_5163);
nand U9048 (N_9048,N_4464,N_4904);
and U9049 (N_9049,N_5705,N_5537);
and U9050 (N_9050,N_5827,N_3289);
nand U9051 (N_9051,N_6070,N_4415);
nand U9052 (N_9052,N_4561,N_4625);
and U9053 (N_9053,N_3415,N_5020);
and U9054 (N_9054,N_5458,N_6196);
xnor U9055 (N_9055,N_5914,N_5873);
nand U9056 (N_9056,N_4582,N_3962);
or U9057 (N_9057,N_3721,N_5711);
or U9058 (N_9058,N_5334,N_5769);
nand U9059 (N_9059,N_5899,N_3693);
xnor U9060 (N_9060,N_3805,N_4886);
or U9061 (N_9061,N_3705,N_4915);
xnor U9062 (N_9062,N_3278,N_4855);
xor U9063 (N_9063,N_4421,N_5810);
nand U9064 (N_9064,N_4531,N_3676);
nand U9065 (N_9065,N_5372,N_5341);
nand U9066 (N_9066,N_5055,N_5291);
or U9067 (N_9067,N_3205,N_4180);
nand U9068 (N_9068,N_5391,N_5162);
nand U9069 (N_9069,N_4282,N_4622);
and U9070 (N_9070,N_3884,N_5753);
xnor U9071 (N_9071,N_6082,N_5826);
nor U9072 (N_9072,N_4782,N_3676);
xor U9073 (N_9073,N_6012,N_3949);
xor U9074 (N_9074,N_4340,N_5930);
and U9075 (N_9075,N_4932,N_5325);
nand U9076 (N_9076,N_5158,N_3757);
nor U9077 (N_9077,N_6238,N_3741);
xor U9078 (N_9078,N_3667,N_5043);
nand U9079 (N_9079,N_3407,N_5113);
or U9080 (N_9080,N_4621,N_3361);
and U9081 (N_9081,N_5605,N_4196);
and U9082 (N_9082,N_5668,N_6008);
or U9083 (N_9083,N_5384,N_6078);
nor U9084 (N_9084,N_6230,N_4679);
nor U9085 (N_9085,N_5786,N_4928);
nand U9086 (N_9086,N_5249,N_5363);
or U9087 (N_9087,N_5173,N_4597);
and U9088 (N_9088,N_5265,N_4686);
or U9089 (N_9089,N_3438,N_4156);
and U9090 (N_9090,N_3192,N_4632);
nand U9091 (N_9091,N_3228,N_4875);
nor U9092 (N_9092,N_3210,N_4528);
nor U9093 (N_9093,N_3916,N_3168);
and U9094 (N_9094,N_3651,N_3952);
nand U9095 (N_9095,N_3382,N_3320);
or U9096 (N_9096,N_5598,N_4825);
nor U9097 (N_9097,N_5050,N_5091);
or U9098 (N_9098,N_5655,N_4605);
or U9099 (N_9099,N_5028,N_3834);
xnor U9100 (N_9100,N_5900,N_5638);
and U9101 (N_9101,N_3631,N_4390);
nor U9102 (N_9102,N_5173,N_6073);
xor U9103 (N_9103,N_6209,N_4395);
nand U9104 (N_9104,N_5337,N_3598);
nand U9105 (N_9105,N_5075,N_4561);
nand U9106 (N_9106,N_6042,N_5206);
or U9107 (N_9107,N_4336,N_3490);
nand U9108 (N_9108,N_5817,N_5689);
or U9109 (N_9109,N_4657,N_4631);
nand U9110 (N_9110,N_6203,N_4471);
and U9111 (N_9111,N_6078,N_5803);
nor U9112 (N_9112,N_3772,N_4816);
and U9113 (N_9113,N_5590,N_3415);
or U9114 (N_9114,N_3293,N_5015);
or U9115 (N_9115,N_4324,N_5699);
nor U9116 (N_9116,N_4054,N_3696);
nor U9117 (N_9117,N_4038,N_3941);
or U9118 (N_9118,N_5024,N_3538);
xor U9119 (N_9119,N_4424,N_5988);
nor U9120 (N_9120,N_3336,N_5786);
or U9121 (N_9121,N_5771,N_4412);
nor U9122 (N_9122,N_3631,N_5694);
or U9123 (N_9123,N_5538,N_4280);
nor U9124 (N_9124,N_3142,N_3778);
and U9125 (N_9125,N_3202,N_3284);
nand U9126 (N_9126,N_4073,N_3656);
and U9127 (N_9127,N_3493,N_5118);
nor U9128 (N_9128,N_3496,N_4504);
and U9129 (N_9129,N_4515,N_5522);
xor U9130 (N_9130,N_3670,N_4411);
or U9131 (N_9131,N_3606,N_5748);
nand U9132 (N_9132,N_6204,N_3719);
or U9133 (N_9133,N_3485,N_5968);
nand U9134 (N_9134,N_4606,N_3356);
and U9135 (N_9135,N_5073,N_3528);
nand U9136 (N_9136,N_3566,N_4822);
or U9137 (N_9137,N_5539,N_3808);
and U9138 (N_9138,N_3261,N_3503);
or U9139 (N_9139,N_5006,N_5340);
nor U9140 (N_9140,N_4862,N_3547);
nor U9141 (N_9141,N_3467,N_5094);
xnor U9142 (N_9142,N_4591,N_5377);
nand U9143 (N_9143,N_6166,N_4684);
nor U9144 (N_9144,N_5442,N_3724);
nor U9145 (N_9145,N_3349,N_3955);
xnor U9146 (N_9146,N_4863,N_3992);
or U9147 (N_9147,N_6203,N_5583);
nand U9148 (N_9148,N_3319,N_5864);
and U9149 (N_9149,N_5492,N_4714);
nand U9150 (N_9150,N_4486,N_3604);
and U9151 (N_9151,N_5922,N_4875);
nor U9152 (N_9152,N_4284,N_5153);
nor U9153 (N_9153,N_6043,N_3784);
nor U9154 (N_9154,N_5804,N_4319);
and U9155 (N_9155,N_4407,N_6016);
or U9156 (N_9156,N_4957,N_5717);
nor U9157 (N_9157,N_3137,N_6173);
or U9158 (N_9158,N_5358,N_5882);
nor U9159 (N_9159,N_3693,N_4618);
or U9160 (N_9160,N_4673,N_3252);
or U9161 (N_9161,N_4448,N_3171);
xor U9162 (N_9162,N_3969,N_4137);
nor U9163 (N_9163,N_4700,N_5385);
nor U9164 (N_9164,N_3137,N_6227);
nor U9165 (N_9165,N_4668,N_5419);
xor U9166 (N_9166,N_3366,N_6210);
nand U9167 (N_9167,N_4987,N_4231);
and U9168 (N_9168,N_5040,N_5518);
and U9169 (N_9169,N_5467,N_5283);
nor U9170 (N_9170,N_3837,N_5352);
and U9171 (N_9171,N_6208,N_5778);
xnor U9172 (N_9172,N_5945,N_3722);
nand U9173 (N_9173,N_5280,N_3538);
or U9174 (N_9174,N_3530,N_5533);
xnor U9175 (N_9175,N_5810,N_6173);
or U9176 (N_9176,N_5673,N_3827);
xor U9177 (N_9177,N_3721,N_5851);
nor U9178 (N_9178,N_3127,N_5336);
or U9179 (N_9179,N_3972,N_6082);
nor U9180 (N_9180,N_5454,N_3670);
nor U9181 (N_9181,N_5148,N_4131);
xnor U9182 (N_9182,N_4035,N_3653);
and U9183 (N_9183,N_5295,N_5769);
nor U9184 (N_9184,N_4962,N_5604);
nand U9185 (N_9185,N_3165,N_5728);
xnor U9186 (N_9186,N_5750,N_3198);
nand U9187 (N_9187,N_5367,N_3812);
nand U9188 (N_9188,N_4235,N_3486);
nor U9189 (N_9189,N_4593,N_4182);
or U9190 (N_9190,N_4412,N_3676);
nand U9191 (N_9191,N_3512,N_4739);
xnor U9192 (N_9192,N_5880,N_3877);
or U9193 (N_9193,N_5563,N_4947);
nand U9194 (N_9194,N_5637,N_4303);
nor U9195 (N_9195,N_4118,N_4932);
and U9196 (N_9196,N_6078,N_5493);
nor U9197 (N_9197,N_5798,N_3209);
nand U9198 (N_9198,N_5033,N_4941);
and U9199 (N_9199,N_6111,N_5988);
nand U9200 (N_9200,N_5431,N_5317);
nand U9201 (N_9201,N_4277,N_5591);
and U9202 (N_9202,N_4552,N_5857);
nor U9203 (N_9203,N_3963,N_4944);
xnor U9204 (N_9204,N_3137,N_4728);
and U9205 (N_9205,N_4406,N_5864);
and U9206 (N_9206,N_5796,N_5320);
or U9207 (N_9207,N_4258,N_6238);
nor U9208 (N_9208,N_3712,N_3367);
nand U9209 (N_9209,N_3715,N_5051);
or U9210 (N_9210,N_3217,N_4041);
nor U9211 (N_9211,N_3460,N_4958);
nand U9212 (N_9212,N_3561,N_5236);
nor U9213 (N_9213,N_4949,N_3665);
and U9214 (N_9214,N_3959,N_5078);
or U9215 (N_9215,N_5166,N_4828);
and U9216 (N_9216,N_5022,N_3359);
xor U9217 (N_9217,N_3353,N_3714);
or U9218 (N_9218,N_4125,N_3494);
and U9219 (N_9219,N_3536,N_4469);
nor U9220 (N_9220,N_5650,N_3171);
or U9221 (N_9221,N_4811,N_3569);
xor U9222 (N_9222,N_4464,N_5772);
nor U9223 (N_9223,N_3598,N_4851);
nor U9224 (N_9224,N_3431,N_4865);
and U9225 (N_9225,N_3572,N_5061);
nand U9226 (N_9226,N_5758,N_3953);
or U9227 (N_9227,N_5066,N_3352);
xor U9228 (N_9228,N_5693,N_5323);
xnor U9229 (N_9229,N_3629,N_5408);
nand U9230 (N_9230,N_4554,N_3399);
nand U9231 (N_9231,N_4153,N_5214);
xnor U9232 (N_9232,N_5713,N_5754);
nand U9233 (N_9233,N_4129,N_4853);
and U9234 (N_9234,N_3414,N_3338);
nor U9235 (N_9235,N_4338,N_4325);
xnor U9236 (N_9236,N_3713,N_5762);
xor U9237 (N_9237,N_4102,N_6094);
nor U9238 (N_9238,N_6166,N_5424);
or U9239 (N_9239,N_3732,N_3697);
nand U9240 (N_9240,N_5745,N_4288);
nor U9241 (N_9241,N_4238,N_6209);
xor U9242 (N_9242,N_4985,N_4565);
and U9243 (N_9243,N_3459,N_4454);
or U9244 (N_9244,N_5990,N_3341);
or U9245 (N_9245,N_4731,N_5303);
or U9246 (N_9246,N_5615,N_4644);
nand U9247 (N_9247,N_6193,N_5616);
and U9248 (N_9248,N_5604,N_3621);
nand U9249 (N_9249,N_4866,N_5272);
and U9250 (N_9250,N_3128,N_4249);
and U9251 (N_9251,N_5574,N_4505);
nor U9252 (N_9252,N_6034,N_3333);
nand U9253 (N_9253,N_4317,N_3550);
and U9254 (N_9254,N_5362,N_4538);
and U9255 (N_9255,N_3746,N_4729);
or U9256 (N_9256,N_4895,N_4277);
nand U9257 (N_9257,N_4954,N_5063);
nor U9258 (N_9258,N_3469,N_4781);
nand U9259 (N_9259,N_3427,N_5346);
nor U9260 (N_9260,N_4477,N_5968);
nor U9261 (N_9261,N_4819,N_4426);
and U9262 (N_9262,N_3636,N_3848);
or U9263 (N_9263,N_3912,N_5739);
or U9264 (N_9264,N_3169,N_5601);
and U9265 (N_9265,N_5524,N_4431);
nand U9266 (N_9266,N_5535,N_5375);
and U9267 (N_9267,N_3146,N_5881);
nand U9268 (N_9268,N_5259,N_4773);
nand U9269 (N_9269,N_4766,N_4500);
nor U9270 (N_9270,N_5603,N_5099);
nand U9271 (N_9271,N_3705,N_4635);
and U9272 (N_9272,N_3186,N_5739);
xor U9273 (N_9273,N_3893,N_3168);
xnor U9274 (N_9274,N_4931,N_4514);
xor U9275 (N_9275,N_4688,N_3368);
xnor U9276 (N_9276,N_3581,N_3643);
and U9277 (N_9277,N_3496,N_5275);
xnor U9278 (N_9278,N_3301,N_5807);
xnor U9279 (N_9279,N_3353,N_5287);
nor U9280 (N_9280,N_3238,N_5591);
and U9281 (N_9281,N_3996,N_5277);
and U9282 (N_9282,N_3690,N_4250);
and U9283 (N_9283,N_4907,N_4902);
or U9284 (N_9284,N_3247,N_5321);
nor U9285 (N_9285,N_4334,N_5119);
and U9286 (N_9286,N_5670,N_3834);
nand U9287 (N_9287,N_3151,N_5751);
and U9288 (N_9288,N_5393,N_3518);
xnor U9289 (N_9289,N_3731,N_3656);
nor U9290 (N_9290,N_6125,N_5210);
or U9291 (N_9291,N_5819,N_5083);
nand U9292 (N_9292,N_3897,N_4491);
xnor U9293 (N_9293,N_4758,N_3469);
xor U9294 (N_9294,N_4299,N_3346);
or U9295 (N_9295,N_4147,N_5528);
nand U9296 (N_9296,N_4288,N_5977);
xor U9297 (N_9297,N_5392,N_5635);
nand U9298 (N_9298,N_3308,N_5160);
xnor U9299 (N_9299,N_5366,N_4368);
nor U9300 (N_9300,N_5083,N_4332);
and U9301 (N_9301,N_5876,N_5337);
or U9302 (N_9302,N_3453,N_5299);
nor U9303 (N_9303,N_3746,N_5126);
nand U9304 (N_9304,N_5535,N_3665);
and U9305 (N_9305,N_5718,N_5928);
or U9306 (N_9306,N_4345,N_5300);
nand U9307 (N_9307,N_3691,N_4285);
nand U9308 (N_9308,N_4876,N_5645);
nand U9309 (N_9309,N_4389,N_5877);
nand U9310 (N_9310,N_5099,N_5394);
nor U9311 (N_9311,N_4910,N_3771);
nor U9312 (N_9312,N_5863,N_4354);
nor U9313 (N_9313,N_4821,N_6031);
nand U9314 (N_9314,N_4089,N_3359);
or U9315 (N_9315,N_5964,N_4746);
nor U9316 (N_9316,N_5551,N_4422);
and U9317 (N_9317,N_4488,N_6196);
nor U9318 (N_9318,N_4896,N_5618);
nor U9319 (N_9319,N_5231,N_3725);
and U9320 (N_9320,N_4587,N_3386);
nand U9321 (N_9321,N_3708,N_4138);
and U9322 (N_9322,N_4936,N_4673);
nor U9323 (N_9323,N_6028,N_4078);
nor U9324 (N_9324,N_4040,N_5177);
nand U9325 (N_9325,N_4506,N_3494);
and U9326 (N_9326,N_5506,N_4877);
nor U9327 (N_9327,N_6000,N_4083);
nand U9328 (N_9328,N_6181,N_6170);
nor U9329 (N_9329,N_3711,N_5330);
nor U9330 (N_9330,N_5203,N_4170);
and U9331 (N_9331,N_5046,N_5686);
nor U9332 (N_9332,N_4123,N_4566);
nor U9333 (N_9333,N_3938,N_3348);
nand U9334 (N_9334,N_4739,N_5862);
nand U9335 (N_9335,N_4613,N_6168);
xnor U9336 (N_9336,N_5124,N_4333);
nor U9337 (N_9337,N_4186,N_5165);
and U9338 (N_9338,N_4147,N_4701);
and U9339 (N_9339,N_4467,N_6050);
and U9340 (N_9340,N_3334,N_4621);
and U9341 (N_9341,N_3613,N_5896);
xnor U9342 (N_9342,N_5178,N_3788);
nand U9343 (N_9343,N_6151,N_3597);
xnor U9344 (N_9344,N_5465,N_3761);
nor U9345 (N_9345,N_4441,N_4505);
nor U9346 (N_9346,N_4243,N_4193);
xnor U9347 (N_9347,N_3367,N_5474);
xor U9348 (N_9348,N_6127,N_3240);
xnor U9349 (N_9349,N_5426,N_5144);
nand U9350 (N_9350,N_5971,N_5729);
and U9351 (N_9351,N_4694,N_5442);
nand U9352 (N_9352,N_5018,N_5860);
nand U9353 (N_9353,N_4422,N_5772);
nor U9354 (N_9354,N_3343,N_5998);
and U9355 (N_9355,N_4067,N_6129);
nor U9356 (N_9356,N_4104,N_4473);
nor U9357 (N_9357,N_5259,N_3945);
xnor U9358 (N_9358,N_6062,N_4012);
and U9359 (N_9359,N_3746,N_5590);
or U9360 (N_9360,N_4973,N_5546);
and U9361 (N_9361,N_4558,N_6172);
or U9362 (N_9362,N_3895,N_4329);
xor U9363 (N_9363,N_3279,N_5033);
xor U9364 (N_9364,N_3289,N_4365);
nand U9365 (N_9365,N_4557,N_5704);
nor U9366 (N_9366,N_5849,N_6002);
xnor U9367 (N_9367,N_6228,N_6041);
and U9368 (N_9368,N_3849,N_3812);
nor U9369 (N_9369,N_5188,N_4766);
xnor U9370 (N_9370,N_5659,N_3738);
xor U9371 (N_9371,N_3820,N_3556);
nand U9372 (N_9372,N_4037,N_4298);
or U9373 (N_9373,N_5571,N_5012);
nor U9374 (N_9374,N_5645,N_3589);
nor U9375 (N_9375,N_8309,N_6320);
or U9376 (N_9376,N_8540,N_8234);
nand U9377 (N_9377,N_8488,N_8889);
xor U9378 (N_9378,N_7832,N_6401);
xor U9379 (N_9379,N_7964,N_7392);
xor U9380 (N_9380,N_8909,N_6912);
nand U9381 (N_9381,N_7359,N_6334);
xnor U9382 (N_9382,N_7292,N_7354);
xor U9383 (N_9383,N_7011,N_8830);
or U9384 (N_9384,N_9233,N_7929);
xor U9385 (N_9385,N_9132,N_7989);
xor U9386 (N_9386,N_7312,N_8794);
xor U9387 (N_9387,N_6498,N_6885);
and U9388 (N_9388,N_8948,N_6790);
nand U9389 (N_9389,N_8829,N_6412);
and U9390 (N_9390,N_8766,N_9116);
nand U9391 (N_9391,N_7881,N_6992);
nor U9392 (N_9392,N_9046,N_6581);
nor U9393 (N_9393,N_8161,N_7251);
nand U9394 (N_9394,N_6668,N_7051);
and U9395 (N_9395,N_7517,N_8220);
or U9396 (N_9396,N_9028,N_8658);
or U9397 (N_9397,N_6374,N_6687);
xnor U9398 (N_9398,N_8086,N_8823);
xor U9399 (N_9399,N_9018,N_8386);
nand U9400 (N_9400,N_7775,N_8742);
nand U9401 (N_9401,N_6847,N_6643);
nor U9402 (N_9402,N_8724,N_8831);
or U9403 (N_9403,N_7304,N_7306);
nand U9404 (N_9404,N_6641,N_6487);
or U9405 (N_9405,N_7424,N_7639);
nor U9406 (N_9406,N_6659,N_6984);
xnor U9407 (N_9407,N_7633,N_6400);
or U9408 (N_9408,N_7166,N_8906);
nor U9409 (N_9409,N_8270,N_8033);
or U9410 (N_9410,N_7048,N_8355);
xor U9411 (N_9411,N_7740,N_8013);
nor U9412 (N_9412,N_7549,N_6416);
xnor U9413 (N_9413,N_7710,N_8068);
nand U9414 (N_9414,N_7723,N_7965);
and U9415 (N_9415,N_6467,N_6597);
nand U9416 (N_9416,N_7461,N_6373);
nand U9417 (N_9417,N_7445,N_6479);
and U9418 (N_9418,N_6795,N_7782);
and U9419 (N_9419,N_8390,N_9324);
nand U9420 (N_9420,N_7285,N_6389);
nor U9421 (N_9421,N_7010,N_8555);
and U9422 (N_9422,N_8259,N_6519);
xnor U9423 (N_9423,N_7019,N_8059);
nor U9424 (N_9424,N_7788,N_6300);
xnor U9425 (N_9425,N_7704,N_6989);
and U9426 (N_9426,N_6665,N_7045);
xnor U9427 (N_9427,N_8789,N_8773);
nor U9428 (N_9428,N_6741,N_8515);
xnor U9429 (N_9429,N_8801,N_8570);
or U9430 (N_9430,N_8617,N_7442);
or U9431 (N_9431,N_6252,N_7018);
xnor U9432 (N_9432,N_8980,N_7142);
xor U9433 (N_9433,N_8656,N_8004);
and U9434 (N_9434,N_9038,N_7602);
nor U9435 (N_9435,N_7590,N_7760);
nor U9436 (N_9436,N_6406,N_8181);
and U9437 (N_9437,N_7800,N_7819);
nor U9438 (N_9438,N_6644,N_9045);
or U9439 (N_9439,N_8786,N_7657);
xor U9440 (N_9440,N_7987,N_7844);
nand U9441 (N_9441,N_8535,N_9175);
xor U9442 (N_9442,N_7626,N_9230);
nand U9443 (N_9443,N_8592,N_6936);
nor U9444 (N_9444,N_9300,N_9353);
nand U9445 (N_9445,N_9053,N_8979);
nor U9446 (N_9446,N_7267,N_8659);
nor U9447 (N_9447,N_6906,N_8827);
xnor U9448 (N_9448,N_6635,N_9000);
xnor U9449 (N_9449,N_6716,N_8958);
nand U9450 (N_9450,N_8095,N_7500);
nand U9451 (N_9451,N_7315,N_8444);
nor U9452 (N_9452,N_8356,N_7383);
nand U9453 (N_9453,N_7348,N_6625);
or U9454 (N_9454,N_7257,N_8833);
nand U9455 (N_9455,N_8426,N_8728);
xnor U9456 (N_9456,N_9075,N_9192);
and U9457 (N_9457,N_7191,N_6604);
xnor U9458 (N_9458,N_8790,N_7105);
nor U9459 (N_9459,N_7938,N_9246);
nand U9460 (N_9460,N_8951,N_7574);
and U9461 (N_9461,N_8195,N_9281);
or U9462 (N_9462,N_8429,N_7095);
nor U9463 (N_9463,N_8674,N_6933);
nand U9464 (N_9464,N_8991,N_9225);
and U9465 (N_9465,N_7956,N_8969);
nand U9466 (N_9466,N_8915,N_7622);
nand U9467 (N_9467,N_9264,N_6398);
nand U9468 (N_9468,N_7181,N_8720);
nand U9469 (N_9469,N_8273,N_6305);
xor U9470 (N_9470,N_8248,N_7571);
and U9471 (N_9471,N_8424,N_7290);
or U9472 (N_9472,N_7620,N_8159);
nor U9473 (N_9473,N_6541,N_7401);
and U9474 (N_9474,N_7263,N_7414);
nor U9475 (N_9475,N_6911,N_6612);
nor U9476 (N_9476,N_6708,N_8895);
nor U9477 (N_9477,N_9009,N_7999);
or U9478 (N_9478,N_6454,N_6350);
nand U9479 (N_9479,N_8230,N_8137);
xor U9480 (N_9480,N_8636,N_7446);
nor U9481 (N_9481,N_6402,N_7258);
or U9482 (N_9482,N_8036,N_8443);
nor U9483 (N_9483,N_6471,N_7103);
nand U9484 (N_9484,N_8152,N_6421);
or U9485 (N_9485,N_9089,N_9207);
or U9486 (N_9486,N_8723,N_8372);
or U9487 (N_9487,N_8471,N_8306);
nand U9488 (N_9488,N_7836,N_8520);
and U9489 (N_9489,N_7222,N_8884);
nor U9490 (N_9490,N_8162,N_6673);
nand U9491 (N_9491,N_6792,N_7243);
and U9492 (N_9492,N_6803,N_9027);
nor U9493 (N_9493,N_7253,N_6898);
nand U9494 (N_9494,N_6493,N_8127);
or U9495 (N_9495,N_7785,N_9173);
nand U9496 (N_9496,N_7572,N_8898);
or U9497 (N_9497,N_8623,N_9163);
nor U9498 (N_9498,N_9321,N_7848);
nand U9499 (N_9499,N_9236,N_7884);
nor U9500 (N_9500,N_7066,N_7365);
xnor U9501 (N_9501,N_8870,N_8070);
xor U9502 (N_9502,N_9272,N_8029);
or U9503 (N_9503,N_8874,N_6411);
and U9504 (N_9504,N_7256,N_6821);
nand U9505 (N_9505,N_8041,N_7773);
or U9506 (N_9506,N_8154,N_9365);
nand U9507 (N_9507,N_9049,N_7981);
nor U9508 (N_9508,N_7717,N_7169);
xnor U9509 (N_9509,N_8448,N_6806);
nand U9510 (N_9510,N_7220,N_8650);
or U9511 (N_9511,N_6379,N_7658);
or U9512 (N_9512,N_9267,N_7289);
or U9513 (N_9513,N_7484,N_7711);
nor U9514 (N_9514,N_8584,N_6520);
and U9515 (N_9515,N_7847,N_6731);
or U9516 (N_9516,N_6796,N_7950);
nand U9517 (N_9517,N_8096,N_8813);
nand U9518 (N_9518,N_6399,N_7300);
and U9519 (N_9519,N_8964,N_8314);
nand U9520 (N_9520,N_6606,N_6884);
nand U9521 (N_9521,N_6955,N_8350);
nor U9522 (N_9522,N_9366,N_7694);
xor U9523 (N_9523,N_7806,N_7208);
or U9524 (N_9524,N_7079,N_6871);
or U9525 (N_9525,N_9087,N_6605);
nor U9526 (N_9526,N_7078,N_8917);
nand U9527 (N_9527,N_8064,N_6337);
nand U9528 (N_9528,N_7230,N_7369);
nand U9529 (N_9529,N_6969,N_8900);
xnor U9530 (N_9530,N_6981,N_7899);
nor U9531 (N_9531,N_7183,N_8608);
or U9532 (N_9532,N_7871,N_7867);
nand U9533 (N_9533,N_9188,N_7521);
nand U9534 (N_9534,N_8896,N_8912);
xnor U9535 (N_9535,N_8366,N_7933);
xnor U9536 (N_9536,N_8179,N_7404);
xnor U9537 (N_9537,N_8688,N_6284);
xnor U9538 (N_9538,N_8304,N_9251);
nor U9539 (N_9539,N_9187,N_6723);
and U9540 (N_9540,N_8691,N_9326);
nor U9541 (N_9541,N_7979,N_6367);
xnor U9542 (N_9542,N_8639,N_7842);
xor U9543 (N_9543,N_9364,N_7917);
or U9544 (N_9544,N_7088,N_6778);
nand U9545 (N_9545,N_8475,N_7813);
or U9546 (N_9546,N_8125,N_6995);
nand U9547 (N_9547,N_8452,N_7612);
and U9548 (N_9548,N_7543,N_7128);
nor U9549 (N_9549,N_8897,N_8343);
nor U9550 (N_9550,N_7471,N_6940);
nand U9551 (N_9551,N_8785,N_8307);
or U9552 (N_9552,N_8435,N_7207);
and U9553 (N_9553,N_6501,N_6975);
or U9554 (N_9554,N_6307,N_6596);
or U9555 (N_9555,N_9114,N_7408);
or U9556 (N_9556,N_8341,N_8732);
and U9557 (N_9557,N_9209,N_8959);
nand U9558 (N_9558,N_9243,N_7238);
and U9559 (N_9559,N_6346,N_6982);
or U9560 (N_9560,N_6507,N_8115);
xor U9561 (N_9561,N_9111,N_8677);
nand U9562 (N_9562,N_6967,N_7943);
nor U9563 (N_9563,N_8046,N_7619);
or U9564 (N_9564,N_8557,N_7156);
or U9565 (N_9565,N_9170,N_9128);
nor U9566 (N_9566,N_8297,N_7497);
nor U9567 (N_9567,N_8453,N_6461);
nor U9568 (N_9568,N_9304,N_6965);
and U9569 (N_9569,N_8071,N_9309);
or U9570 (N_9570,N_6922,N_6321);
or U9571 (N_9571,N_7994,N_6712);
and U9572 (N_9572,N_8178,N_8873);
or U9573 (N_9573,N_8971,N_7250);
nor U9574 (N_9574,N_6774,N_6862);
or U9575 (N_9575,N_9041,N_8147);
and U9576 (N_9576,N_8292,N_7162);
nand U9577 (N_9577,N_6525,N_6697);
nand U9578 (N_9578,N_6896,N_9021);
nand U9579 (N_9579,N_8202,N_8295);
xor U9580 (N_9580,N_7475,N_6759);
nand U9581 (N_9581,N_7034,N_8200);
and U9582 (N_9582,N_8711,N_6483);
xnor U9583 (N_9583,N_7921,N_8803);
nand U9584 (N_9584,N_6286,N_8301);
nor U9585 (N_9585,N_6433,N_6894);
nand U9586 (N_9586,N_8715,N_7457);
xnor U9587 (N_9587,N_9091,N_7685);
or U9588 (N_9588,N_6345,N_8845);
or U9589 (N_9589,N_8963,N_7124);
xnor U9590 (N_9590,N_6571,N_7108);
and U9591 (N_9591,N_8726,N_8903);
and U9592 (N_9592,N_8910,N_8411);
xor U9593 (N_9593,N_7906,N_9210);
or U9594 (N_9594,N_6527,N_7014);
nand U9595 (N_9595,N_8293,N_7254);
or U9596 (N_9596,N_9360,N_8467);
nand U9597 (N_9597,N_8911,N_8837);
nor U9598 (N_9598,N_7515,N_7623);
nand U9599 (N_9599,N_8970,N_7167);
xor U9600 (N_9600,N_9019,N_7866);
or U9601 (N_9601,N_7826,N_8373);
nor U9602 (N_9602,N_6856,N_7377);
or U9603 (N_9603,N_7667,N_7038);
nor U9604 (N_9604,N_6667,N_6876);
and U9605 (N_9605,N_7393,N_8529);
and U9606 (N_9606,N_7789,N_7485);
nor U9607 (N_9607,N_9219,N_8001);
nor U9608 (N_9608,N_7864,N_6424);
nand U9609 (N_9609,N_6548,N_6468);
nand U9610 (N_9610,N_9084,N_8354);
nand U9611 (N_9611,N_9354,N_9314);
nor U9612 (N_9612,N_6757,N_6623);
and U9613 (N_9613,N_8423,N_7883);
nor U9614 (N_9614,N_7988,N_8579);
nor U9615 (N_9615,N_7777,N_7216);
or U9616 (N_9616,N_7926,N_8439);
nor U9617 (N_9617,N_8569,N_7265);
or U9618 (N_9618,N_6572,N_6877);
nand U9619 (N_9619,N_7960,N_6892);
nor U9620 (N_9620,N_6480,N_6458);
or U9621 (N_9621,N_9013,N_6655);
nand U9622 (N_9622,N_8709,N_6509);
nor U9623 (N_9623,N_8264,N_8937);
nor U9624 (N_9624,N_8414,N_8985);
and U9625 (N_9625,N_8016,N_6949);
and U9626 (N_9626,N_6575,N_7287);
nor U9627 (N_9627,N_7647,N_7570);
xor U9628 (N_9628,N_7621,N_7232);
nand U9629 (N_9629,N_7770,N_6829);
nor U9630 (N_9630,N_7488,N_9295);
and U9631 (N_9631,N_7118,N_8308);
and U9632 (N_9632,N_7294,N_8591);
or U9633 (N_9633,N_6749,N_9277);
and U9634 (N_9634,N_6545,N_8408);
xor U9635 (N_9635,N_8278,N_8363);
nor U9636 (N_9636,N_9164,N_6564);
and U9637 (N_9637,N_8318,N_7396);
or U9638 (N_9638,N_7828,N_8498);
or U9639 (N_9639,N_8929,N_7990);
nor U9640 (N_9640,N_8242,N_7086);
nor U9641 (N_9641,N_6407,N_8196);
or U9642 (N_9642,N_7610,N_8327);
or U9643 (N_9643,N_8818,N_6423);
xnor U9644 (N_9644,N_8999,N_8719);
and U9645 (N_9645,N_6584,N_7525);
or U9646 (N_9646,N_6743,N_6409);
xnor U9647 (N_9647,N_7690,N_6392);
or U9648 (N_9648,N_8565,N_7060);
and U9649 (N_9649,N_7781,N_7052);
nand U9650 (N_9650,N_9216,N_7439);
xor U9651 (N_9651,N_6561,N_8871);
or U9652 (N_9652,N_6784,N_8641);
nor U9653 (N_9653,N_9303,N_7652);
or U9654 (N_9654,N_8085,N_7918);
or U9655 (N_9655,N_8705,N_7855);
and U9656 (N_9656,N_6262,N_6253);
xnor U9657 (N_9657,N_8702,N_8208);
or U9658 (N_9658,N_7040,N_8129);
nand U9659 (N_9659,N_7131,N_9115);
or U9660 (N_9660,N_7920,N_8133);
nand U9661 (N_9661,N_7930,N_7947);
nand U9662 (N_9662,N_7178,N_8776);
or U9663 (N_9663,N_9217,N_8024);
nand U9664 (N_9664,N_7958,N_8673);
nor U9665 (N_9665,N_7210,N_9103);
nor U9666 (N_9666,N_6628,N_7474);
nand U9667 (N_9667,N_7101,N_8167);
or U9668 (N_9668,N_8795,N_9190);
nor U9669 (N_9669,N_7767,N_7957);
nor U9670 (N_9670,N_7399,N_8023);
and U9671 (N_9671,N_6730,N_7391);
or U9672 (N_9672,N_7952,N_8245);
and U9673 (N_9673,N_8268,N_7159);
or U9674 (N_9674,N_7875,N_7235);
and U9675 (N_9675,N_7577,N_7636);
xor U9676 (N_9676,N_9288,N_6266);
nand U9677 (N_9677,N_7309,N_9048);
or U9678 (N_9678,N_8582,N_7675);
or U9679 (N_9679,N_7153,N_9339);
or U9680 (N_9680,N_6474,N_7659);
or U9681 (N_9681,N_6742,N_8485);
nor U9682 (N_9682,N_7043,N_6557);
and U9683 (N_9683,N_6717,N_7218);
nand U9684 (N_9684,N_8014,N_6931);
nor U9685 (N_9685,N_7948,N_7498);
xnor U9686 (N_9686,N_7878,N_9061);
xor U9687 (N_9687,N_8775,N_6325);
or U9688 (N_9688,N_6558,N_8566);
and U9689 (N_9689,N_9335,N_8735);
and U9690 (N_9690,N_7506,N_8274);
and U9691 (N_9691,N_6811,N_9119);
nor U9692 (N_9692,N_7523,N_7384);
or U9693 (N_9693,N_6593,N_8380);
and U9694 (N_9694,N_8788,N_6376);
and U9695 (N_9695,N_7106,N_7793);
and U9696 (N_9696,N_7469,N_7027);
nor U9697 (N_9697,N_8396,N_7737);
or U9698 (N_9698,N_7379,N_9244);
or U9699 (N_9699,N_6278,N_7650);
nor U9700 (N_9700,N_8457,N_6858);
xnor U9701 (N_9701,N_6848,N_6343);
and U9702 (N_9702,N_7597,N_7064);
and U9703 (N_9703,N_6588,N_7479);
nor U9704 (N_9704,N_9051,N_9313);
nor U9705 (N_9705,N_9249,N_6466);
nand U9706 (N_9706,N_7601,N_8104);
nand U9707 (N_9707,N_8962,N_7234);
nand U9708 (N_9708,N_8523,N_7795);
nor U9709 (N_9709,N_8215,N_7431);
xnor U9710 (N_9710,N_7198,N_8784);
and U9711 (N_9711,N_7606,N_8932);
nand U9712 (N_9712,N_9117,N_9350);
xor U9713 (N_9713,N_9323,N_7464);
or U9714 (N_9714,N_6491,N_8561);
and U9715 (N_9715,N_7308,N_8404);
or U9716 (N_9716,N_6941,N_6580);
and U9717 (N_9717,N_7538,N_7288);
xnor U9718 (N_9718,N_8822,N_8627);
xor U9719 (N_9719,N_7729,N_7302);
nand U9720 (N_9720,N_8984,N_6720);
or U9721 (N_9721,N_8696,N_7527);
nand U9722 (N_9722,N_7319,N_7629);
nor U9723 (N_9723,N_7746,N_7205);
and U9724 (N_9724,N_8533,N_6359);
xor U9725 (N_9725,N_8432,N_7037);
nand U9726 (N_9726,N_8568,N_8083);
and U9727 (N_9727,N_8412,N_6381);
nor U9728 (N_9728,N_9302,N_7858);
and U9729 (N_9729,N_9224,N_7651);
xor U9730 (N_9730,N_6878,N_6469);
or U9731 (N_9731,N_6622,N_9227);
xor U9732 (N_9732,N_8840,N_8849);
nor U9733 (N_9733,N_8155,N_7966);
nand U9734 (N_9734,N_6448,N_7024);
xor U9735 (N_9735,N_8060,N_6434);
xnor U9736 (N_9736,N_8119,N_7046);
nand U9737 (N_9737,N_7357,N_8619);
nand U9738 (N_9738,N_8043,N_9002);
xnor U9739 (N_9739,N_7055,N_6304);
nand U9740 (N_9740,N_9139,N_7152);
or U9741 (N_9741,N_9158,N_6642);
or U9742 (N_9742,N_6630,N_8197);
and U9743 (N_9743,N_6485,N_7587);
xnor U9744 (N_9744,N_9343,N_6762);
or U9745 (N_9745,N_7646,N_7366);
nor U9746 (N_9746,N_8078,N_7067);
and U9747 (N_9747,N_7708,N_6875);
and U9748 (N_9748,N_7790,N_7049);
or U9749 (N_9749,N_6926,N_6393);
or U9750 (N_9750,N_6983,N_7876);
or U9751 (N_9751,N_8280,N_8166);
nor U9752 (N_9752,N_6577,N_9130);
nor U9753 (N_9753,N_8713,N_6427);
nand U9754 (N_9754,N_8881,N_6355);
or U9755 (N_9755,N_9361,N_8493);
xnor U9756 (N_9756,N_8762,N_8516);
or U9757 (N_9757,N_7411,N_8668);
and U9758 (N_9758,N_7534,N_8199);
and U9759 (N_9759,N_6522,N_8755);
xor U9760 (N_9760,N_7008,N_8267);
nor U9761 (N_9761,N_8205,N_8872);
and U9762 (N_9762,N_8111,N_6654);
xnor U9763 (N_9763,N_7036,N_6768);
and U9764 (N_9764,N_6499,N_6861);
xnor U9765 (N_9765,N_7077,N_7147);
xnor U9766 (N_9766,N_7170,N_6935);
xor U9767 (N_9767,N_7430,N_8558);
or U9768 (N_9768,N_8997,N_8342);
or U9769 (N_9769,N_7664,N_6649);
nand U9770 (N_9770,N_8624,N_7532);
or U9771 (N_9771,N_7645,N_7598);
or U9772 (N_9772,N_6658,N_7042);
and U9773 (N_9773,N_8554,N_8758);
nand U9774 (N_9774,N_9297,N_8291);
nand U9775 (N_9775,N_6375,N_7419);
xor U9776 (N_9776,N_6349,N_8644);
nand U9777 (N_9777,N_8814,N_7451);
xor U9778 (N_9778,N_8940,N_6455);
xnor U9779 (N_9779,N_7341,N_8545);
or U9780 (N_9780,N_7363,N_9273);
or U9781 (N_9781,N_7890,N_7324);
nand U9782 (N_9782,N_7346,N_8358);
and U9783 (N_9783,N_9214,N_8103);
or U9784 (N_9784,N_6739,N_9341);
and U9785 (N_9785,N_7172,N_7127);
nor U9786 (N_9786,N_8028,N_6993);
xor U9787 (N_9787,N_8235,N_7565);
nor U9788 (N_9788,N_6497,N_7148);
nand U9789 (N_9789,N_8074,N_8421);
nand U9790 (N_9790,N_6978,N_7749);
or U9791 (N_9791,N_7436,N_9065);
and U9792 (N_9792,N_8954,N_9200);
or U9793 (N_9793,N_9133,N_7507);
nor U9794 (N_9794,N_7576,N_9247);
nand U9795 (N_9795,N_9104,N_7678);
and U9796 (N_9796,N_8527,N_8804);
nand U9797 (N_9797,N_7089,N_8405);
and U9798 (N_9798,N_7168,N_7528);
nand U9799 (N_9799,N_7386,N_9182);
nor U9800 (N_9800,N_8986,N_7703);
xor U9801 (N_9801,N_6808,N_8779);
nand U9802 (N_9802,N_8681,N_8106);
or U9803 (N_9803,N_8797,N_6533);
nand U9804 (N_9804,N_7279,N_7735);
and U9805 (N_9805,N_7882,N_9149);
nand U9806 (N_9806,N_9305,N_6396);
nor U9807 (N_9807,N_7797,N_7483);
and U9808 (N_9808,N_7119,N_6590);
nor U9809 (N_9809,N_8337,N_8393);
nor U9810 (N_9810,N_7231,N_8740);
nor U9811 (N_9811,N_7245,N_6728);
and U9812 (N_9812,N_7397,N_8721);
or U9813 (N_9813,N_6369,N_7900);
or U9814 (N_9814,N_6903,N_7677);
and U9815 (N_9815,N_8328,N_6939);
and U9816 (N_9816,N_7718,N_7504);
nand U9817 (N_9817,N_9318,N_8003);
or U9818 (N_9818,N_8759,N_7149);
xor U9819 (N_9819,N_8972,N_7083);
or U9820 (N_9820,N_8503,N_6329);
nor U9821 (N_9821,N_6394,N_8771);
nand U9822 (N_9822,N_7155,N_6341);
or U9823 (N_9823,N_8602,N_8838);
nor U9824 (N_9824,N_7996,N_8102);
and U9825 (N_9825,N_8645,N_6645);
xnor U9826 (N_9826,N_7567,N_8254);
nand U9827 (N_9827,N_8620,N_6705);
nor U9828 (N_9828,N_8654,N_8808);
and U9829 (N_9829,N_7827,N_8333);
and U9830 (N_9830,N_8231,N_8302);
and U9831 (N_9831,N_9107,N_6948);
xor U9832 (N_9832,N_7143,N_7100);
nand U9833 (N_9833,N_8692,N_6816);
nand U9834 (N_9834,N_9024,N_8596);
xnor U9835 (N_9835,N_8148,N_7846);
xor U9836 (N_9836,N_6290,N_9059);
or U9837 (N_9837,N_9369,N_8781);
and U9838 (N_9838,N_7811,N_7144);
nor U9839 (N_9839,N_8228,N_9081);
and U9840 (N_9840,N_6704,N_7531);
xnor U9841 (N_9841,N_8010,N_7971);
and U9842 (N_9842,N_8055,N_8743);
and U9843 (N_9843,N_7068,N_8441);
xnor U9844 (N_9844,N_8796,N_6632);
nand U9845 (N_9845,N_9261,N_6974);
xor U9846 (N_9846,N_9189,N_7969);
or U9847 (N_9847,N_7420,N_8073);
or U9848 (N_9848,N_8415,N_7801);
or U9849 (N_9849,N_9008,N_6333);
or U9850 (N_9850,N_8395,N_7164);
xor U9851 (N_9851,N_9319,N_6870);
nand U9852 (N_9852,N_8015,N_8279);
xor U9853 (N_9853,N_8360,N_8576);
or U9854 (N_9854,N_7841,N_8953);
and U9855 (N_9855,N_8683,N_6805);
nor U9856 (N_9856,N_8581,N_7542);
nand U9857 (N_9857,N_7074,N_8930);
and U9858 (N_9858,N_8486,N_6377);
nor U9859 (N_9859,N_8011,N_9242);
nand U9860 (N_9860,N_7829,N_8418);
and U9861 (N_9861,N_6494,N_9358);
or U9862 (N_9862,N_7266,N_6299);
xnor U9863 (N_9863,N_7936,N_6954);
or U9864 (N_9864,N_8760,N_8543);
nor U9865 (N_9865,N_8611,N_8300);
nand U9866 (N_9866,N_6651,N_6609);
and U9867 (N_9867,N_7277,N_7237);
xor U9868 (N_9868,N_8739,N_6823);
and U9869 (N_9869,N_6490,N_6279);
and U9870 (N_9870,N_6797,N_8989);
nor U9871 (N_9871,N_6582,N_8470);
nand U9872 (N_9872,N_6313,N_9290);
or U9873 (N_9873,N_8651,N_9085);
or U9874 (N_9874,N_6452,N_9262);
nand U9875 (N_9875,N_6288,N_7478);
nor U9876 (N_9876,N_7214,N_8922);
or U9877 (N_9877,N_7810,N_8116);
or U9878 (N_9878,N_8587,N_7177);
or U9879 (N_9879,N_7575,N_9152);
xnor U9880 (N_9880,N_7705,N_9289);
nand U9881 (N_9881,N_8560,N_6255);
nand U9882 (N_9882,N_7395,N_9347);
and U9883 (N_9883,N_7697,N_6924);
and U9884 (N_9884,N_8142,N_7454);
xnor U9885 (N_9885,N_8761,N_6351);
xnor U9886 (N_9886,N_8857,N_9362);
nor U9887 (N_9887,N_8737,N_6827);
xor U9888 (N_9888,N_8902,N_8577);
nor U9889 (N_9889,N_6842,N_9346);
xnor U9890 (N_9890,N_7186,N_7189);
or U9891 (N_9891,N_9368,N_6734);
and U9892 (N_9892,N_7752,N_8667);
and U9893 (N_9893,N_8745,N_7759);
nor U9894 (N_9894,N_7213,N_6419);
or U9895 (N_9895,N_7325,N_8050);
and U9896 (N_9896,N_7713,N_9222);
nand U9897 (N_9897,N_8381,N_9179);
nor U9898 (N_9898,N_7944,N_8539);
nand U9899 (N_9899,N_8512,N_8479);
nand U9900 (N_9900,N_7856,N_8661);
and U9901 (N_9901,N_6834,N_8921);
xnor U9902 (N_9902,N_6457,N_6624);
and U9903 (N_9903,N_8334,N_9078);
nor U9904 (N_9904,N_8362,N_8311);
and U9905 (N_9905,N_9331,N_8082);
xor U9906 (N_9906,N_7671,N_8826);
nand U9907 (N_9907,N_9235,N_7002);
or U9908 (N_9908,N_8262,N_9287);
or U9909 (N_9909,N_8916,N_8933);
nor U9910 (N_9910,N_9240,N_8186);
nand U9911 (N_9911,N_6947,N_8752);
nor U9912 (N_9912,N_7092,N_8614);
and U9913 (N_9913,N_8224,N_6793);
and U9914 (N_9914,N_7000,N_7734);
nor U9915 (N_9915,N_6570,N_7140);
xor U9916 (N_9916,N_7228,N_6388);
nor U9917 (N_9917,N_8514,N_8955);
nand U9918 (N_9918,N_8144,N_8975);
and U9919 (N_9919,N_7323,N_9333);
or U9920 (N_9920,N_6611,N_6818);
xnor U9921 (N_9921,N_7295,N_6781);
and U9922 (N_9922,N_8397,N_8714);
nand U9923 (N_9923,N_8239,N_9180);
and U9924 (N_9924,N_6976,N_7762);
nand U9925 (N_9925,N_8009,N_7683);
and U9926 (N_9926,N_8383,N_7780);
nor U9927 (N_9927,N_9142,N_7805);
and U9928 (N_9928,N_8810,N_6315);
nor U9929 (N_9929,N_8253,N_8047);
or U9930 (N_9930,N_8678,N_9094);
or U9931 (N_9931,N_6319,N_7047);
nand U9932 (N_9932,N_7426,N_7953);
nor U9933 (N_9933,N_7466,N_6985);
nand U9934 (N_9934,N_8243,N_7284);
or U9935 (N_9935,N_8156,N_8690);
nand U9936 (N_9936,N_8824,N_8710);
xor U9937 (N_9937,N_7955,N_8689);
nor U9938 (N_9938,N_7353,N_8131);
and U9939 (N_9939,N_7229,N_6602);
nor U9940 (N_9940,N_8496,N_8266);
and U9941 (N_9941,N_8244,N_8192);
and U9942 (N_9942,N_6257,N_7986);
xnor U9943 (N_9943,N_8981,N_7910);
xnor U9944 (N_9944,N_7462,N_8176);
or U9945 (N_9945,N_7865,N_7908);
or U9946 (N_9946,N_6357,N_9263);
nand U9947 (N_9947,N_7098,N_7702);
nor U9948 (N_9948,N_8031,N_6962);
and U9949 (N_9949,N_7480,N_6271);
xor U9950 (N_9950,N_7834,N_7879);
xnor U9951 (N_9951,N_6456,N_7932);
and U9952 (N_9952,N_7050,N_8330);
nand U9953 (N_9953,N_7916,N_7540);
nand U9954 (N_9954,N_7432,N_6820);
xor U9955 (N_9955,N_6966,N_6559);
xnor U9956 (N_9956,N_8583,N_6785);
nand U9957 (N_9957,N_9283,N_6599);
or U9958 (N_9958,N_6258,N_7361);
nand U9959 (N_9959,N_6619,N_8361);
xnor U9960 (N_9960,N_7467,N_8815);
nor U9961 (N_9961,N_8864,N_7907);
xor U9962 (N_9962,N_9102,N_7406);
nand U9963 (N_9963,N_9312,N_6486);
xor U9964 (N_9964,N_7758,N_6874);
nor U9965 (N_9965,N_6414,N_7894);
nand U9966 (N_9966,N_9015,N_6715);
and U9967 (N_9967,N_8382,N_9023);
nor U9968 (N_9968,N_7580,N_6740);
xnor U9969 (N_9969,N_9030,N_9159);
nor U9970 (N_9970,N_8855,N_9032);
xor U9971 (N_9971,N_6335,N_6869);
nand U9972 (N_9972,N_7812,N_9156);
and U9973 (N_9973,N_8780,N_7513);
or U9974 (N_9974,N_7934,N_7299);
xor U9975 (N_9975,N_8151,N_9168);
or U9976 (N_9976,N_7925,N_8676);
and U9977 (N_9977,N_6798,N_7796);
xnor U9978 (N_9978,N_7495,N_7692);
and U9979 (N_9979,N_7555,N_7364);
and U9980 (N_9980,N_8532,N_9035);
and U9981 (N_9981,N_8216,N_8035);
xor U9982 (N_9982,N_6987,N_8030);
nor U9983 (N_9983,N_8012,N_7338);
and U9984 (N_9984,N_9017,N_6565);
nand U9985 (N_9985,N_7129,N_8860);
and U9986 (N_9986,N_8778,N_7020);
nor U9987 (N_9987,N_8474,N_7732);
or U9988 (N_9988,N_7814,N_6640);
xnor U9989 (N_9989,N_8092,N_6825);
or U9990 (N_9990,N_7840,N_7502);
nor U9991 (N_9991,N_8489,N_7271);
or U9992 (N_9992,N_6621,N_9183);
nand U9993 (N_9993,N_9184,N_6365);
nor U9994 (N_9994,N_8447,N_9074);
nor U9995 (N_9995,N_8777,N_6857);
nor U9996 (N_9996,N_8173,N_9334);
nand U9997 (N_9997,N_8550,N_7317);
or U9998 (N_9998,N_8919,N_9201);
nand U9999 (N_9999,N_6953,N_6574);
or U10000 (N_10000,N_9037,N_8521);
xnor U10001 (N_10001,N_7815,N_7779);
or U10002 (N_10002,N_8883,N_7490);
and U10003 (N_10003,N_7154,N_9076);
and U10004 (N_10004,N_6316,N_7374);
nor U10005 (N_10005,N_7044,N_9160);
nand U10006 (N_10006,N_9072,N_9073);
and U10007 (N_10007,N_7766,N_8339);
nand U10008 (N_10008,N_7830,N_6724);
xor U10009 (N_10009,N_6372,N_8770);
or U10010 (N_10010,N_6826,N_7311);
nand U10011 (N_10011,N_7816,N_7056);
nor U10012 (N_10012,N_7187,N_8206);
or U10013 (N_10013,N_9204,N_9213);
and U10014 (N_10014,N_7026,N_6817);
xnor U10015 (N_10015,N_7672,N_6745);
and U10016 (N_10016,N_8237,N_9134);
nand U10017 (N_10017,N_8700,N_8646);
and U10018 (N_10018,N_8240,N_8947);
and U10019 (N_10019,N_9329,N_7298);
or U10020 (N_10020,N_8221,N_6804);
or U10021 (N_10021,N_6370,N_9113);
nor U10022 (N_10022,N_9100,N_7594);
or U10023 (N_10023,N_7013,N_8213);
xor U10024 (N_10024,N_7141,N_7526);
nand U10025 (N_10025,N_9348,N_8886);
nor U10026 (N_10026,N_8572,N_7967);
nand U10027 (N_10027,N_7371,N_6542);
xnor U10028 (N_10028,N_8296,N_7337);
nor U10029 (N_10029,N_7477,N_8519);
nand U10030 (N_10030,N_9291,N_6505);
nor U10031 (N_10031,N_8499,N_6900);
nor U10032 (N_10032,N_9255,N_8893);
and U10033 (N_10033,N_8157,N_7850);
and U10034 (N_10034,N_9036,N_9174);
or U10035 (N_10035,N_6569,N_7902);
or U10036 (N_10036,N_8580,N_6292);
xnor U10037 (N_10037,N_9055,N_8665);
and U10038 (N_10038,N_7945,N_7763);
xor U10039 (N_10039,N_6475,N_8034);
xor U10040 (N_10040,N_7617,N_9373);
nor U10041 (N_10041,N_9006,N_8251);
nor U10042 (N_10042,N_6986,N_8635);
and U10043 (N_10043,N_6354,N_8787);
nor U10044 (N_10044,N_8288,N_8392);
nor U10045 (N_10045,N_6838,N_7973);
or U10046 (N_10046,N_9274,N_9259);
nor U10047 (N_10047,N_9282,N_8663);
and U10048 (N_10048,N_8836,N_9062);
xnor U10049 (N_10049,N_8946,N_6528);
and U10050 (N_10050,N_8163,N_6907);
xnor U10051 (N_10051,N_6958,N_7328);
and U10052 (N_10052,N_8571,N_6405);
nor U10053 (N_10053,N_6783,N_6666);
nor U10054 (N_10054,N_9294,N_8349);
and U10055 (N_10055,N_6537,N_7138);
and U10056 (N_10056,N_6694,N_9203);
and U10057 (N_10057,N_8536,N_8615);
nand U10058 (N_10058,N_7197,N_7334);
nor U10059 (N_10059,N_7259,N_8445);
nor U10060 (N_10060,N_7915,N_6617);
nand U10061 (N_10061,N_7756,N_9197);
nand U10062 (N_10062,N_9260,N_8120);
nor U10063 (N_10063,N_8169,N_7370);
or U10064 (N_10064,N_7211,N_6945);
xnor U10065 (N_10065,N_7030,N_8391);
and U10066 (N_10066,N_7712,N_7557);
xnor U10067 (N_10067,N_8260,N_6314);
xor U10068 (N_10068,N_9101,N_8194);
and U10069 (N_10069,N_8212,N_8388);
nor U10070 (N_10070,N_8590,N_6689);
and U10071 (N_10071,N_9060,N_8487);
xnor U10072 (N_10072,N_6352,N_8145);
or U10073 (N_10073,N_9344,N_7928);
nor U10074 (N_10074,N_8124,N_7496);
xnor U10075 (N_10075,N_7435,N_7347);
nand U10076 (N_10076,N_6729,N_7449);
nor U10077 (N_10077,N_8126,N_7247);
and U10078 (N_10078,N_9181,N_8828);
xor U10079 (N_10079,N_7784,N_8706);
or U10080 (N_10080,N_7333,N_7799);
or U10081 (N_10081,N_6899,N_9371);
xor U10082 (N_10082,N_7120,N_6779);
and U10083 (N_10083,N_9337,N_6883);
and U10084 (N_10084,N_7453,N_8629);
nand U10085 (N_10085,N_8704,N_6988);
nand U10086 (N_10086,N_8846,N_6770);
xnor U10087 (N_10087,N_7403,N_7520);
xnor U10088 (N_10088,N_6767,N_6344);
and U10089 (N_10089,N_6855,N_7798);
xnor U10090 (N_10090,N_8338,N_6330);
nor U10091 (N_10091,N_9058,N_7774);
and U10092 (N_10092,N_7772,N_8918);
nand U10093 (N_10093,N_8305,N_7778);
nand U10094 (N_10094,N_6317,N_7503);
or U10095 (N_10095,N_6713,N_7874);
or U10096 (N_10096,N_6629,N_8730);
xnor U10097 (N_10097,N_8000,N_8416);
nand U10098 (N_10098,N_7997,N_8522);
xor U10099 (N_10099,N_8633,N_6880);
nor U10100 (N_10100,N_8121,N_7891);
nand U10101 (N_10101,N_7429,N_7058);
nor U10102 (N_10102,N_7951,N_7217);
or U10103 (N_10103,N_9338,N_7561);
and U10104 (N_10104,N_8364,N_7360);
xor U10105 (N_10105,N_8812,N_7742);
nand U10106 (N_10106,N_7508,N_7427);
or U10107 (N_10107,N_6618,N_6444);
xnor U10108 (N_10108,N_6553,N_8850);
xnor U10109 (N_10109,N_7402,N_6693);
nor U10110 (N_10110,N_8226,N_8741);
nand U10111 (N_10111,N_8854,N_7530);
and U10112 (N_10112,N_7085,N_6309);
nand U10113 (N_10113,N_9284,N_7946);
nor U10114 (N_10114,N_6919,N_9092);
nor U10115 (N_10115,N_6991,N_8025);
or U10116 (N_10116,N_6752,N_8128);
or U10117 (N_10117,N_7904,N_7838);
nand U10118 (N_10118,N_6523,N_8269);
or U10119 (N_10119,N_8171,N_9252);
and U10120 (N_10120,N_7861,N_8621);
or U10121 (N_10121,N_7887,N_8298);
nand U10122 (N_10122,N_6386,N_8585);
nand U10123 (N_10123,N_8865,N_6518);
and U10124 (N_10124,N_6589,N_7771);
xnor U10125 (N_10125,N_8482,N_7573);
or U10126 (N_10126,N_7698,N_7725);
xnor U10127 (N_10127,N_7145,N_7588);
or U10128 (N_10128,N_7303,N_7741);
nor U10129 (N_10129,N_7322,N_8575);
or U10130 (N_10130,N_8506,N_6657);
xnor U10131 (N_10131,N_7632,N_7161);
nand U10132 (N_10132,N_8105,N_7959);
or U10133 (N_10133,N_9178,N_8626);
xor U10134 (N_10134,N_8807,N_9218);
or U10135 (N_10135,N_7291,N_7150);
xnor U10136 (N_10136,N_6539,N_8227);
or U10137 (N_10137,N_8223,N_7362);
nand U10138 (N_10138,N_7889,N_7489);
and U10139 (N_10139,N_9278,N_6680);
or U10140 (N_10140,N_7059,N_9223);
and U10141 (N_10141,N_7073,N_8336);
xnor U10142 (N_10142,N_7417,N_7727);
and U10143 (N_10143,N_7977,N_7133);
xor U10144 (N_10144,N_8122,N_7722);
and U10145 (N_10145,N_7356,N_7716);
xnor U10146 (N_10146,N_6637,N_6994);
and U10147 (N_10147,N_9315,N_7991);
nand U10148 (N_10148,N_9016,N_7927);
xor U10149 (N_10149,N_6727,N_9025);
or U10150 (N_10150,N_8722,N_8492);
nand U10151 (N_10151,N_7367,N_6633);
and U10152 (N_10152,N_6272,N_8538);
xor U10153 (N_10153,N_8401,N_8477);
xor U10154 (N_10154,N_6601,N_6773);
xor U10155 (N_10155,N_6718,N_6476);
or U10156 (N_10156,N_9003,N_8738);
xor U10157 (N_10157,N_7548,N_7888);
xor U10158 (N_10158,N_9285,N_8282);
or U10159 (N_10159,N_8748,N_9150);
nor U10160 (N_10160,N_7082,N_6442);
or U10161 (N_10161,N_8344,N_8861);
xor U10162 (N_10162,N_7157,N_7335);
xnor U10163 (N_10163,N_8184,N_7553);
xor U10164 (N_10164,N_7822,N_8544);
nor U10165 (N_10165,N_8089,N_6824);
or U10166 (N_10166,N_6613,N_9239);
or U10167 (N_10167,N_8772,N_6746);
and U10168 (N_10168,N_8057,N_7736);
xnor U10169 (N_10169,N_8021,N_7663);
xor U10170 (N_10170,N_8586,N_7151);
nor U10171 (N_10171,N_8613,N_7007);
xnor U10172 (N_10172,N_7615,N_7857);
nor U10173 (N_10173,N_8019,N_7400);
nand U10174 (N_10174,N_6810,N_8075);
xor U10175 (N_10175,N_7137,N_9050);
nor U10176 (N_10176,N_8058,N_6780);
or U10177 (N_10177,N_7195,N_8394);
xor U10178 (N_10178,N_7352,N_8859);
nand U10179 (N_10179,N_8842,N_9144);
or U10180 (N_10180,N_6653,N_8791);
nor U10181 (N_10181,N_8261,N_7116);
and U10182 (N_10182,N_7776,N_8802);
and U10183 (N_10183,N_7345,N_6714);
nand U10184 (N_10184,N_7407,N_7820);
nor U10185 (N_10185,N_7970,N_7821);
xor U10186 (N_10186,N_8118,N_6721);
nand U10187 (N_10187,N_7968,N_6563);
nor U10188 (N_10188,N_6521,N_7286);
nor U10189 (N_10189,N_6404,N_8232);
or U10190 (N_10190,N_8130,N_8143);
and U10191 (N_10191,N_6859,N_7744);
and U10192 (N_10192,N_7505,N_6303);
nand U10193 (N_10193,N_7270,N_9079);
nand U10194 (N_10194,N_8725,N_7935);
nand U10195 (N_10195,N_9120,N_6864);
nor U10196 (N_10196,N_6338,N_7919);
nand U10197 (N_10197,N_7090,N_7595);
or U10198 (N_10198,N_6610,N_6626);
xnor U10199 (N_10199,N_8956,N_7681);
nor U10200 (N_10200,N_7993,N_6891);
nand U10201 (N_10201,N_7984,N_7227);
and U10202 (N_10202,N_9345,N_8138);
nand U10203 (N_10203,N_8563,N_8042);
nand U10204 (N_10204,N_7460,N_6930);
and U10205 (N_10205,N_8793,N_7372);
nand U10206 (N_10206,N_6504,N_7627);
xnor U10207 (N_10207,N_9064,N_9034);
or U10208 (N_10208,N_6791,N_7459);
nor U10209 (N_10209,N_7547,N_6867);
nor U10210 (N_10210,N_8548,N_8018);
nand U10211 (N_10211,N_7340,N_6280);
and U10212 (N_10212,N_9057,N_6917);
nor U10213 (N_10213,N_7202,N_7624);
xor U10214 (N_10214,N_6535,N_7873);
or U10215 (N_10215,N_9098,N_9157);
and U10216 (N_10216,N_9202,N_6296);
or U10217 (N_10217,N_6436,N_8727);
or U10218 (N_10218,N_8564,N_6866);
nand U10219 (N_10219,N_6362,N_7937);
or U10220 (N_10220,N_6417,N_8271);
nor U10221 (N_10221,N_7261,N_6276);
or U10222 (N_10222,N_6786,N_9292);
nand U10223 (N_10223,N_7422,N_9090);
xnor U10224 (N_10224,N_6839,N_8885);
nand U10225 (N_10225,N_8464,N_7731);
xor U10226 (N_10226,N_7831,N_9234);
nand U10227 (N_10227,N_9301,N_6662);
nand U10228 (N_10228,N_8882,N_7413);
nand U10229 (N_10229,N_8257,N_8559);
nor U10230 (N_10230,N_8450,N_9138);
nand U10231 (N_10231,N_8942,N_7223);
nand U10232 (N_10232,N_8546,N_8634);
or U10233 (N_10233,N_6550,N_9109);
xnor U10234 (N_10234,N_8434,N_8335);
xor U10235 (N_10235,N_8653,N_6737);
and U10236 (N_10236,N_8880,N_6530);
or U10237 (N_10237,N_9095,N_6492);
or U10238 (N_10238,N_6543,N_7558);
nor U10239 (N_10239,N_6482,N_9351);
nor U10240 (N_10240,N_6771,N_9250);
nor U10241 (N_10241,N_7190,N_6777);
xnor U10242 (N_10242,N_7443,N_7661);
or U10243 (N_10243,N_6800,N_7751);
and U10244 (N_10244,N_7075,N_8247);
xor U10245 (N_10245,N_8935,N_9083);
nand U10246 (N_10246,N_7226,N_6736);
or U10247 (N_10247,N_6268,N_6835);
or U10248 (N_10248,N_8751,N_7676);
nor U10249 (N_10249,N_6356,N_8891);
and U10250 (N_10250,N_8767,N_6684);
nand U10251 (N_10251,N_6942,N_8250);
xnor U10252 (N_10252,N_7388,N_6297);
or U10253 (N_10253,N_6837,N_8508);
and U10254 (N_10254,N_8285,N_8140);
nor U10255 (N_10255,N_6702,N_9020);
nor U10256 (N_10256,N_6478,N_8183);
and U10257 (N_10257,N_8322,N_8640);
or U10258 (N_10258,N_7618,N_7452);
or U10259 (N_10259,N_7682,N_9280);
nor U10260 (N_10260,N_6722,N_7314);
nand U10261 (N_10261,N_8648,N_8669);
and U10262 (N_10262,N_7541,N_8844);
nor U10263 (N_10263,N_7069,N_8469);
or U10264 (N_10264,N_6614,N_8852);
xor U10265 (N_10265,N_9330,N_8117);
and U10266 (N_10266,N_7662,N_6547);
and U10267 (N_10267,N_6822,N_6664);
xnor U10268 (N_10268,N_8319,N_6364);
and U10269 (N_10269,N_6766,N_7272);
or U10270 (N_10270,N_8146,N_8218);
nor U10271 (N_10271,N_9268,N_9317);
and U10272 (N_10272,N_6439,N_6371);
xnor U10273 (N_10273,N_8534,N_6566);
and U10274 (N_10274,N_7336,N_6595);
or U10275 (N_10275,N_7962,N_6650);
and U10276 (N_10276,N_7689,N_8053);
nand U10277 (N_10277,N_6938,N_6937);
and U10278 (N_10278,N_7041,N_7221);
nand U10279 (N_10279,N_8407,N_7438);
xnor U10280 (N_10280,N_8733,N_8990);
nand U10281 (N_10281,N_8204,N_9129);
nor U10282 (N_10282,N_7769,N_7903);
or U10283 (N_10283,N_6915,N_8065);
or U10284 (N_10284,N_6851,N_7680);
or U10285 (N_10285,N_8701,N_6979);
xor U10286 (N_10286,N_6432,N_7039);
nand U10287 (N_10287,N_7423,N_6512);
nand U10288 (N_10288,N_7843,N_8265);
and U10289 (N_10289,N_8461,N_8061);
nand U10290 (N_10290,N_8967,N_6860);
and U10291 (N_10291,N_8172,N_6710);
or U10292 (N_10292,N_7941,N_8312);
nor U10293 (N_10293,N_9096,N_6287);
nand U10294 (N_10294,N_6676,N_9198);
xor U10295 (N_10295,N_7125,N_6620);
and U10296 (N_10296,N_6368,N_6709);
or U10297 (N_10297,N_8877,N_8995);
xnor U10298 (N_10298,N_6264,N_6273);
nor U10299 (N_10299,N_8923,N_8983);
xnor U10300 (N_10300,N_6735,N_6435);
nand U10301 (N_10301,N_6814,N_7721);
nor U10302 (N_10302,N_6972,N_7139);
and U10303 (N_10303,N_6695,N_7081);
or U10304 (N_10304,N_8887,N_6470);
nand U10305 (N_10305,N_7670,N_7310);
xor U10306 (N_10306,N_8988,N_6681);
nor U10307 (N_10307,N_7854,N_6382);
nand U10308 (N_10308,N_6863,N_8431);
or U10309 (N_10309,N_7327,N_7537);
nand U10310 (N_10310,N_9169,N_6598);
nand U10311 (N_10311,N_8736,N_7985);
or U10312 (N_10312,N_8045,N_6677);
xnor U10313 (N_10313,N_8682,N_6536);
or U10314 (N_10314,N_7909,N_8229);
or U10315 (N_10315,N_6690,N_9299);
and U10316 (N_10316,N_8134,N_8994);
nand U10317 (N_10317,N_7648,N_6840);
and U10318 (N_10318,N_7603,N_6908);
nand U10319 (N_10319,N_8595,N_8107);
nor U10320 (N_10320,N_8422,N_8458);
nor U10321 (N_10321,N_6923,N_8325);
xnor U10322 (N_10322,N_6451,N_6699);
nor U10323 (N_10323,N_6447,N_7583);
and U10324 (N_10324,N_7358,N_6782);
or U10325 (N_10325,N_7440,N_6897);
nand U10326 (N_10326,N_6685,N_8294);
and U10327 (N_10327,N_7091,N_8040);
or U10328 (N_10328,N_7104,N_7176);
nor U10329 (N_10329,N_8907,N_8135);
nor U10330 (N_10330,N_6327,N_6920);
and U10331 (N_10331,N_7192,N_6868);
nand U10332 (N_10332,N_6358,N_8832);
and U10333 (N_10333,N_8056,N_9245);
nand U10334 (N_10334,N_8928,N_6889);
xor U10335 (N_10335,N_8547,N_7200);
or U10336 (N_10336,N_9226,N_8729);
nand U10337 (N_10337,N_8160,N_6928);
nand U10338 (N_10338,N_8525,N_7853);
xor U10339 (N_10339,N_7715,N_7412);
or U10340 (N_10340,N_8924,N_7182);
nand U10341 (N_10341,N_7895,N_7219);
and U10342 (N_10342,N_8649,N_8685);
xor U10343 (N_10343,N_7269,N_6503);
or U10344 (N_10344,N_8717,N_7415);
xnor U10345 (N_10345,N_9221,N_6970);
xor U10346 (N_10346,N_9042,N_9071);
nand U10347 (N_10347,N_8643,N_6882);
or U10348 (N_10348,N_8908,N_6959);
or U10349 (N_10349,N_7005,N_6560);
and U10350 (N_10350,N_7880,N_6873);
nand U10351 (N_10351,N_7748,N_8604);
xnor U10352 (N_10352,N_7241,N_7434);
or U10353 (N_10353,N_8925,N_6348);
or U10354 (N_10354,N_6261,N_6960);
and U10355 (N_10355,N_7385,N_8878);
xnor U10356 (N_10356,N_8141,N_6332);
nor U10357 (N_10357,N_8079,N_8976);
and U10358 (N_10358,N_7691,N_8410);
nand U10359 (N_10359,N_8472,N_8281);
and U10360 (N_10360,N_7330,N_7355);
nor U10361 (N_10361,N_7476,N_9155);
or U10362 (N_10362,N_8456,N_7693);
or U10363 (N_10363,N_8753,N_6756);
nand U10364 (N_10364,N_7535,N_6437);
nor U10365 (N_10365,N_8610,N_8625);
or U10366 (N_10366,N_6263,N_8400);
or U10367 (N_10367,N_7837,N_6418);
xor U10368 (N_10368,N_7791,N_7080);
nor U10369 (N_10369,N_7509,N_9229);
nand U10370 (N_10370,N_8601,N_6481);
and U10371 (N_10371,N_6449,N_9108);
nor U10372 (N_10372,N_7444,N_9033);
nand U10373 (N_10373,N_7087,N_8599);
xor U10374 (N_10374,N_8892,N_8528);
nand U10375 (N_10375,N_7350,N_9131);
or U10376 (N_10376,N_6340,N_6893);
nor U10377 (N_10377,N_6872,N_6555);
or U10378 (N_10378,N_7028,N_7886);
nor U10379 (N_10379,N_8764,N_7719);
or U10380 (N_10380,N_6410,N_6802);
xor U10381 (N_10381,N_6438,N_8462);
nor U10382 (N_10382,N_7463,N_8589);
xor U10383 (N_10383,N_6833,N_8081);
xor U10384 (N_10384,N_6250,N_7094);
xor U10385 (N_10385,N_8816,N_8526);
nand U10386 (N_10386,N_8697,N_8920);
nor U10387 (N_10387,N_8573,N_7654);
or U10388 (N_10388,N_7494,N_8905);
and U10389 (N_10389,N_9077,N_7747);
or U10390 (N_10390,N_7248,N_9286);
nand U10391 (N_10391,N_6318,N_7807);
xnor U10392 (N_10392,N_9215,N_8153);
and U10393 (N_10393,N_6506,N_8090);
nor U10394 (N_10394,N_7076,N_7233);
nor U10395 (N_10395,N_6957,N_6639);
nor U10396 (N_10396,N_9271,N_6719);
nand U10397 (N_10397,N_7109,N_7107);
xnor U10398 (N_10398,N_7614,N_6758);
nand U10399 (N_10399,N_8190,N_6725);
nand U10400 (N_10400,N_6671,N_7132);
xnor U10401 (N_10401,N_8977,N_6585);
nor U10402 (N_10402,N_9340,N_8943);
and U10403 (N_10403,N_6426,N_7185);
or U10404 (N_10404,N_8017,N_8026);
xor U10405 (N_10405,N_6927,N_8945);
nor U10406 (N_10406,N_7562,N_8660);
nand U10407 (N_10407,N_8747,N_8049);
or U10408 (N_10408,N_8398,N_8574);
and U10409 (N_10409,N_8647,N_9069);
nand U10410 (N_10410,N_8191,N_6583);
nor U10411 (N_10411,N_8501,N_8326);
or U10412 (N_10412,N_8480,N_7099);
nand U10413 (N_10413,N_8110,N_9316);
nor U10414 (N_10414,N_7802,N_8420);
and U10415 (N_10415,N_6277,N_8246);
and U10416 (N_10416,N_6425,N_7012);
and U10417 (N_10417,N_7017,N_9328);
xnor U10418 (N_10418,N_7761,N_8863);
and U10419 (N_10419,N_6283,N_8769);
xnor U10420 (N_10420,N_8631,N_8749);
xor U10421 (N_10421,N_8209,N_8598);
nor U10422 (N_10422,N_7533,N_7378);
nor U10423 (N_10423,N_6510,N_9349);
xnor U10424 (N_10424,N_7199,N_6934);
xnor U10425 (N_10425,N_9148,N_6850);
nor U10426 (N_10426,N_9070,N_8066);
xor U10427 (N_10427,N_8438,N_9056);
xnor U10428 (N_10428,N_8618,N_7146);
xnor U10429 (N_10429,N_8468,N_7995);
xnor U10430 (N_10430,N_9063,N_8834);
xnor U10431 (N_10431,N_8821,N_6775);
and U10432 (N_10432,N_6788,N_8098);
nor U10433 (N_10433,N_6913,N_7033);
nand U10434 (N_10434,N_8992,N_6395);
and U10435 (N_10435,N_9199,N_8944);
nor U10436 (N_10436,N_6932,N_7922);
nand U10437 (N_10437,N_7175,N_7817);
nand U10438 (N_10438,N_6384,N_7870);
nand U10439 (N_10439,N_7914,N_8455);
nand U10440 (N_10440,N_8365,N_8437);
nand U10441 (N_10441,N_7236,N_7342);
xnor U10442 (N_10442,N_9265,N_6440);
xnor U10443 (N_10443,N_8371,N_6865);
nand U10444 (N_10444,N_7262,N_7447);
and U10445 (N_10445,N_8376,N_8258);
or U10446 (N_10446,N_8370,N_7554);
and U10447 (N_10447,N_6323,N_9121);
or U10448 (N_10448,N_7130,N_8320);
and U10449 (N_10449,N_9191,N_7701);
or U10450 (N_10450,N_9254,N_8553);
nand U10451 (N_10451,N_6683,N_7568);
xnor U10452 (N_10452,N_6910,N_8357);
and U10453 (N_10453,N_7696,N_8384);
nor U10454 (N_10454,N_7514,N_8346);
xnor U10455 (N_10455,N_8982,N_7297);
nor U10456 (N_10456,N_7249,N_8214);
nor U10457 (N_10457,N_8038,N_8276);
or U10458 (N_10458,N_7410,N_7134);
and U10459 (N_10459,N_8965,N_8007);
nor U10460 (N_10460,N_7016,N_7188);
nor U10461 (N_10461,N_7281,N_6636);
nand U10462 (N_10462,N_9125,N_8321);
xnor U10463 (N_10463,N_7174,N_9336);
or U10464 (N_10464,N_7679,N_6921);
and U10465 (N_10465,N_8783,N_9105);
and U10466 (N_10466,N_8109,N_8556);
and U10467 (N_10467,N_7825,N_6301);
and U10468 (N_10468,N_6285,N_7745);
xor U10469 (N_10469,N_6391,N_8936);
and U10470 (N_10470,N_6380,N_7110);
or U10471 (N_10471,N_8862,N_6799);
and U10472 (N_10472,N_6946,N_7607);
and U10473 (N_10473,N_9279,N_8352);
nor U10474 (N_10474,N_7885,N_6849);
nor U10475 (N_10475,N_8368,N_6661);
nand U10476 (N_10476,N_6765,N_9165);
xor U10477 (N_10477,N_7173,N_7025);
or U10478 (N_10478,N_8466,N_6776);
and U10479 (N_10479,N_8961,N_7872);
nand U10480 (N_10480,N_8694,N_8290);
xor U10481 (N_10481,N_6513,N_6460);
nor U10482 (N_10482,N_7158,N_8806);
nand U10483 (N_10483,N_8158,N_8483);
nor U10484 (N_10484,N_6360,N_9231);
nor U10485 (N_10485,N_7863,N_6306);
nor U10486 (N_10486,N_6812,N_8087);
or U10487 (N_10487,N_7260,N_8331);
and U10488 (N_10488,N_7470,N_8960);
or U10489 (N_10489,N_8403,N_7808);
xnor U10490 (N_10490,N_7898,N_8768);
or U10491 (N_10491,N_7409,N_7180);
xnor U10492 (N_10492,N_9154,N_8939);
nand U10493 (N_10493,N_8672,N_6843);
xnor U10494 (N_10494,N_7115,N_7792);
or U10495 (N_10495,N_8504,N_6441);
nand U10496 (N_10496,N_6546,N_6794);
or U10497 (N_10497,N_9293,N_6706);
xor U10498 (N_10498,N_7739,N_7135);
nor U10499 (N_10499,N_7976,N_7686);
xor U10500 (N_10500,N_6663,N_6902);
nor U10501 (N_10501,N_7268,N_6514);
xor U10502 (N_10502,N_7849,N_7121);
and U10503 (N_10503,N_8731,N_6809);
and U10504 (N_10504,N_9196,N_9332);
nand U10505 (N_10505,N_8671,N_8637);
nor U10506 (N_10506,N_6445,N_7823);
xnor U10507 (N_10507,N_8949,N_8114);
xnor U10508 (N_10508,N_7635,N_9122);
xnor U10509 (N_10509,N_7394,N_7071);
nor U10510 (N_10510,N_6807,N_8256);
and U10511 (N_10511,N_6311,N_9211);
and U10512 (N_10512,N_7316,N_7114);
or U10513 (N_10513,N_6591,N_9086);
or U10514 (N_10514,N_7511,N_7072);
or U10515 (N_10515,N_9097,N_9310);
xor U10516 (N_10516,N_9135,N_6888);
nor U10517 (N_10517,N_7428,N_8219);
and U10518 (N_10518,N_6387,N_9012);
or U10519 (N_10519,N_6852,N_9307);
xor U10520 (N_10520,N_8588,N_8820);
xnor U10521 (N_10521,N_8113,N_7240);
or U10522 (N_10522,N_8329,N_6990);
xor U10523 (N_10523,N_6692,N_7794);
or U10524 (N_10524,N_6648,N_8686);
nor U10525 (N_10525,N_7455,N_9306);
nor U10526 (N_10526,N_7700,N_8819);
or U10527 (N_10527,N_9146,N_9112);
or U10528 (N_10528,N_7117,N_7545);
xnor U10529 (N_10529,N_7293,N_8524);
nand U10530 (N_10530,N_6508,N_7510);
nand U10531 (N_10531,N_9275,N_7600);
or U10532 (N_10532,N_6524,N_6294);
nand U10533 (N_10533,N_7591,N_7924);
nor U10534 (N_10534,N_6747,N_6390);
and U10535 (N_10535,N_7940,N_8463);
xor U10536 (N_10536,N_9136,N_7062);
nor U10537 (N_10537,N_8888,N_8782);
nand U10538 (N_10538,N_7239,N_6312);
or U10539 (N_10539,N_8094,N_8756);
or U10540 (N_10540,N_6686,N_9093);
or U10541 (N_10541,N_7942,N_6281);
or U10542 (N_10542,N_8606,N_7486);
and U10543 (N_10543,N_6477,N_7305);
nand U10544 (N_10544,N_8377,N_7524);
xnor U10545 (N_10545,N_8518,N_8465);
and U10546 (N_10546,N_6450,N_6540);
nor U10547 (N_10547,N_6567,N_8490);
and U10548 (N_10548,N_7949,N_7974);
xnor U10549 (N_10549,N_8185,N_7982);
xnor U10550 (N_10550,N_9298,N_8193);
or U10551 (N_10551,N_7564,N_8562);
and U10552 (N_10552,N_7499,N_8542);
and U10553 (N_10553,N_8996,N_8509);
xnor U10554 (N_10554,N_8500,N_8409);
nor U10555 (N_10555,N_8537,N_8973);
or U10556 (N_10556,N_8054,N_6275);
and U10557 (N_10557,N_6289,N_7021);
and U10558 (N_10558,N_7738,N_7998);
or U10559 (N_10559,N_7518,N_9110);
nor U10560 (N_10560,N_6308,N_8002);
nor U10561 (N_10561,N_9206,N_7833);
and U10562 (N_10562,N_7673,N_7860);
or U10563 (N_10563,N_6260,N_9088);
xnor U10564 (N_10564,N_6748,N_8351);
or U10565 (N_10565,N_7803,N_8303);
xor U10566 (N_10566,N_7382,N_7634);
nand U10567 (N_10567,N_7611,N_7196);
nor U10568 (N_10568,N_8578,N_6554);
nor U10569 (N_10569,N_8310,N_8695);
or U10570 (N_10570,N_6328,N_8347);
and U10571 (N_10571,N_7931,N_7911);
or U10572 (N_10572,N_6600,N_7437);
nand U10573 (N_10573,N_7616,N_9195);
and U10574 (N_10574,N_8856,N_7730);
and U10575 (N_10575,N_7054,N_9357);
xor U10576 (N_10576,N_9106,N_7006);
nand U10577 (N_10577,N_6707,N_6429);
nor U10578 (N_10578,N_7070,N_8077);
nor U10579 (N_10579,N_7787,N_8774);
xor U10580 (N_10580,N_7608,N_8494);
nor U10581 (N_10581,N_7126,N_8084);
nor U10582 (N_10582,N_7845,N_7613);
xnor U10583 (N_10583,N_7638,N_7275);
or U10584 (N_10584,N_8399,N_9171);
nand U10585 (N_10585,N_7343,N_6634);
nand U10586 (N_10586,N_6916,N_6764);
or U10587 (N_10587,N_8652,N_7093);
nand U10588 (N_10588,N_7512,N_6647);
nand U10589 (N_10589,N_6925,N_7009);
and U10590 (N_10590,N_6755,N_8020);
xor U10591 (N_10591,N_8841,N_7035);
or U10592 (N_10592,N_8687,N_8993);
nand U10593 (N_10593,N_8428,N_8076);
nand U10594 (N_10594,N_7065,N_9099);
or U10595 (N_10595,N_8848,N_8006);
xnor U10596 (N_10596,N_8174,N_7552);
or U10597 (N_10597,N_9010,N_6904);
xor U10598 (N_10598,N_9043,N_7398);
nor U10599 (N_10599,N_6881,N_7852);
xnor U10600 (N_10600,N_6568,N_8189);
nor U10601 (N_10601,N_7481,N_8630);
xor U10602 (N_10602,N_8491,N_8353);
or U10603 (N_10603,N_7923,N_8005);
and U10604 (N_10604,N_7897,N_8707);
nor U10605 (N_10605,N_9342,N_7023);
nand U10606 (N_10606,N_7031,N_7544);
nand U10607 (N_10607,N_8754,N_6473);
nor U10608 (N_10608,N_6751,N_8716);
and U10609 (N_10609,N_8374,N_6556);
and U10610 (N_10610,N_7593,N_8952);
xnor U10611 (N_10611,N_7980,N_6844);
and U10612 (N_10612,N_6801,N_8817);
nor U10613 (N_10613,N_8150,N_7939);
xnor U10614 (N_10614,N_8389,N_8164);
nor U10615 (N_10615,N_7456,N_7660);
nor U10616 (N_10616,N_8379,N_6511);
nand U10617 (N_10617,N_9147,N_7862);
nand U10618 (N_10618,N_6251,N_8097);
or U10619 (N_10619,N_7961,N_7877);
or U10620 (N_10620,N_7283,N_8484);
and U10621 (N_10621,N_8008,N_8938);
and U10622 (N_10622,N_7653,N_6660);
and U10623 (N_10623,N_8340,N_8843);
or U10624 (N_10624,N_8684,N_7193);
nand U10625 (N_10625,N_7380,N_6701);
xnor U10626 (N_10626,N_9177,N_8638);
or U10627 (N_10627,N_6495,N_7839);
nand U10628 (N_10628,N_9372,N_9185);
nand U10629 (N_10629,N_7688,N_7582);
or U10630 (N_10630,N_8825,N_9355);
or U10631 (N_10631,N_8662,N_6484);
nor U10632 (N_10632,N_8597,N_6836);
nand U10633 (N_10633,N_7215,N_7061);
xor U10634 (N_10634,N_6336,N_6830);
nor U10635 (N_10635,N_7112,N_8799);
xnor U10636 (N_10636,N_7373,N_6586);
xor U10637 (N_10637,N_7390,N_7913);
nand U10638 (N_10638,N_8876,N_6615);
nor U10639 (N_10639,N_7954,N_8241);
nand U10640 (N_10640,N_8950,N_6422);
nor U10641 (N_10641,N_8926,N_8108);
or U10642 (N_10642,N_6254,N_8657);
and U10643 (N_10643,N_6531,N_8436);
and U10644 (N_10644,N_9220,N_7421);
nand U10645 (N_10645,N_9039,N_7163);
or U10646 (N_10646,N_8378,N_9370);
or U10647 (N_10647,N_8289,N_8839);
nand U10648 (N_10648,N_7728,N_8275);
nor U10649 (N_10649,N_7783,N_9151);
xor U10650 (N_10650,N_8402,N_6576);
nor U10651 (N_10651,N_8367,N_7418);
or U10652 (N_10652,N_7022,N_8879);
or U10653 (N_10653,N_7529,N_8914);
xor U10654 (N_10654,N_8063,N_9248);
xor U10655 (N_10655,N_8699,N_8136);
and U10656 (N_10656,N_7349,N_7706);
xor U10657 (N_10657,N_7123,N_6516);
or U10658 (N_10658,N_9325,N_7586);
or U10659 (N_10659,N_6488,N_7029);
or U10660 (N_10660,N_7868,N_6688);
and U10661 (N_10661,N_6549,N_7684);
nor U10662 (N_10662,N_6385,N_6669);
and U10663 (N_10663,N_7912,N_7381);
nand U10664 (N_10664,N_7546,N_8609);
xor U10665 (N_10665,N_7589,N_8698);
xnor U10666 (N_10666,N_9011,N_9208);
or U10667 (N_10667,N_7282,N_8901);
nand U10668 (N_10668,N_8263,N_6603);
or U10669 (N_10669,N_6973,N_6607);
and U10670 (N_10670,N_8287,N_7387);
or U10671 (N_10671,N_8927,N_9161);
and U10672 (N_10672,N_8552,N_6672);
nor U10673 (N_10673,N_6963,N_7786);
and U10674 (N_10674,N_7755,N_7896);
and U10675 (N_10675,N_9374,N_7492);
xor U10676 (N_10676,N_8369,N_8679);
or U10677 (N_10677,N_6750,N_9137);
and U10678 (N_10678,N_8454,N_9266);
and U10679 (N_10679,N_7625,N_8594);
nand U10680 (N_10680,N_9044,N_6322);
xor U10681 (N_10681,N_6646,N_7473);
nor U10682 (N_10682,N_6944,N_8062);
nand U10683 (N_10683,N_8670,N_7720);
and U10684 (N_10684,N_8123,N_8430);
and U10685 (N_10685,N_6529,N_8449);
nor U10686 (N_10686,N_7631,N_7307);
and U10687 (N_10687,N_9001,N_7004);
xnor U10688 (N_10688,N_9052,N_8044);
and U10689 (N_10689,N_6453,N_7859);
or U10690 (N_10690,N_6587,N_9162);
or U10691 (N_10691,N_6977,N_9238);
nand U10692 (N_10692,N_7255,N_9258);
xnor U10693 (N_10693,N_6691,N_8187);
or U10694 (N_10694,N_8481,N_6298);
or U10695 (N_10695,N_6256,N_6879);
or U10696 (N_10696,N_6420,N_8165);
and U10697 (N_10697,N_8513,N_6950);
nor U10698 (N_10698,N_7707,N_7640);
xor U10699 (N_10699,N_8616,N_8315);
xnor U10700 (N_10700,N_9296,N_8811);
nand U10701 (N_10701,N_7201,N_6627);
nand U10702 (N_10702,N_7975,N_7482);
and U10703 (N_10703,N_6696,N_7687);
and U10704 (N_10704,N_8517,N_8866);
nor U10705 (N_10705,N_8612,N_7001);
nand U10706 (N_10706,N_6732,N_8283);
xor U10707 (N_10707,N_8080,N_7630);
and U10708 (N_10708,N_6496,N_7818);
and U10709 (N_10709,N_8744,N_9270);
and U10710 (N_10710,N_8800,N_8869);
or U10711 (N_10711,N_6674,N_6678);
xnor U10712 (N_10712,N_8476,N_9256);
xnor U10713 (N_10713,N_7179,N_7753);
and U10714 (N_10714,N_9014,N_8890);
nor U10715 (N_10715,N_9327,N_6502);
xor U10716 (N_10716,N_7522,N_6443);
or U10717 (N_10717,N_8567,N_7032);
and U10718 (N_10718,N_6534,N_6918);
nand U10719 (N_10719,N_8792,N_6552);
nor U10720 (N_10720,N_8680,N_8180);
or U10721 (N_10721,N_8703,N_9237);
xor U10722 (N_10722,N_6353,N_6841);
nand U10723 (N_10723,N_7869,N_9123);
or U10724 (N_10724,N_7244,N_7184);
nand U10725 (N_10725,N_7764,N_7389);
nor U10726 (N_10726,N_6670,N_9166);
nor U10727 (N_10727,N_8419,N_7726);
and U10728 (N_10728,N_7487,N_7754);
xnor U10729 (N_10729,N_6832,N_9253);
nand U10730 (N_10730,N_6901,N_6347);
or U10731 (N_10731,N_8442,N_7122);
or U10732 (N_10732,N_7578,N_7963);
nand U10733 (N_10733,N_8101,N_6465);
nor U10734 (N_10734,N_8460,N_8664);
xor U10735 (N_10735,N_6997,N_6828);
xor U10736 (N_10736,N_6980,N_8088);
or U10737 (N_10737,N_8051,N_8440);
nand U10738 (N_10738,N_8170,N_8324);
xor U10739 (N_10739,N_9322,N_7733);
and U10740 (N_10740,N_9232,N_8666);
xor U10741 (N_10741,N_8039,N_7743);
and U10742 (N_10742,N_7204,N_6472);
or U10743 (N_10743,N_9153,N_6302);
or U10744 (N_10744,N_8286,N_7242);
xnor U10745 (N_10745,N_7274,N_8313);
or U10746 (N_10746,N_8099,N_8968);
and U10747 (N_10747,N_6951,N_7892);
and U10748 (N_10748,N_8427,N_9276);
or U10749 (N_10749,N_6291,N_6675);
or U10750 (N_10750,N_8868,N_6819);
and U10751 (N_10751,N_6853,N_7992);
nor U10752 (N_10752,N_6464,N_8316);
nand U10753 (N_10753,N_8478,N_8233);
xnor U10754 (N_10754,N_8332,N_6463);
nor U10755 (N_10755,N_6265,N_7416);
nand U10756 (N_10756,N_9067,N_7053);
or U10757 (N_10757,N_8510,N_8765);
nor U10758 (N_10758,N_7584,N_6592);
nor U10759 (N_10759,N_8207,N_6763);
or U10760 (N_10760,N_7666,N_8904);
or U10761 (N_10761,N_8345,N_7057);
nand U10762 (N_10762,N_9047,N_6769);
or U10763 (N_10763,N_8284,N_8225);
nand U10764 (N_10764,N_6267,N_8913);
nor U10765 (N_10765,N_9186,N_7609);
or U10766 (N_10766,N_6914,N_7224);
nand U10767 (N_10767,N_8425,N_6366);
nor U10768 (N_10768,N_6711,N_8531);
nand U10769 (N_10769,N_7699,N_8502);
nor U10770 (N_10770,N_8805,N_7649);
xor U10771 (N_10771,N_7724,N_9193);
xor U10772 (N_10772,N_7212,N_7273);
xor U10773 (N_10773,N_6282,N_7893);
and U10774 (N_10774,N_7111,N_6886);
xor U10775 (N_10775,N_8867,N_6428);
or U10776 (N_10776,N_6738,N_6532);
nor U10777 (N_10777,N_8941,N_6813);
xor U10778 (N_10778,N_7329,N_8317);
and U10779 (N_10779,N_9118,N_7246);
and U10780 (N_10780,N_6489,N_9126);
or U10781 (N_10781,N_7278,N_6815);
nand U10782 (N_10782,N_7579,N_7516);
xnor U10783 (N_10783,N_6259,N_6787);
nand U10784 (N_10784,N_7809,N_7550);
xor U10785 (N_10785,N_8175,N_8100);
or U10786 (N_10786,N_6579,N_8132);
nand U10787 (N_10787,N_6459,N_9363);
or U10788 (N_10788,N_9007,N_6293);
or U10789 (N_10789,N_8875,N_9127);
nor U10790 (N_10790,N_7674,N_7203);
nor U10791 (N_10791,N_9172,N_8069);
xnor U10792 (N_10792,N_8655,N_6462);
nand U10793 (N_10793,N_8894,N_8238);
and U10794 (N_10794,N_8978,N_7765);
or U10795 (N_10795,N_7468,N_6383);
xnor U10796 (N_10796,N_8593,N_6403);
nand U10797 (N_10797,N_8052,N_6909);
or U10798 (N_10798,N_7318,N_8712);
xnor U10799 (N_10799,N_9367,N_7344);
nor U10800 (N_10800,N_8433,N_8718);
and U10801 (N_10801,N_6772,N_8987);
nand U10802 (N_10802,N_9068,N_6526);
or U10803 (N_10803,N_9140,N_9257);
xor U10804 (N_10804,N_7556,N_9176);
xor U10805 (N_10805,N_7592,N_7441);
xnor U10806 (N_10806,N_6703,N_6363);
and U10807 (N_10807,N_8858,N_7225);
xnor U10808 (N_10808,N_7264,N_6573);
nand U10809 (N_10809,N_6905,N_9356);
nand U10810 (N_10810,N_8809,N_7665);
or U10811 (N_10811,N_9145,N_6361);
and U10812 (N_10812,N_7581,N_7368);
xnor U10813 (N_10813,N_8198,N_6562);
xor U10814 (N_10814,N_6431,N_7491);
xor U10815 (N_10815,N_7599,N_6608);
xnor U10816 (N_10816,N_7560,N_6342);
nand U10817 (N_10817,N_8222,N_8750);
nor U10818 (N_10818,N_6890,N_8255);
and U10819 (N_10819,N_7519,N_8277);
xor U10820 (N_10820,N_8459,N_7851);
nor U10821 (N_10821,N_8139,N_8451);
nor U10822 (N_10822,N_9143,N_9040);
and U10823 (N_10823,N_9311,N_6996);
nand U10824 (N_10824,N_9004,N_6733);
nor U10825 (N_10825,N_7206,N_7465);
nand U10826 (N_10826,N_6500,N_7252);
and U10827 (N_10827,N_8182,N_8798);
or U10828 (N_10828,N_8899,N_8675);
or U10829 (N_10829,N_8530,N_7551);
and U10830 (N_10830,N_7003,N_8211);
nor U10831 (N_10831,N_8934,N_7824);
and U10832 (N_10832,N_8272,N_8851);
and U10833 (N_10833,N_8149,N_6998);
nand U10834 (N_10834,N_6616,N_9022);
xor U10835 (N_10835,N_7901,N_8112);
or U10836 (N_10836,N_7596,N_8957);
nor U10837 (N_10837,N_7669,N_8549);
xnor U10838 (N_10838,N_7301,N_7695);
xnor U10839 (N_10839,N_7768,N_8505);
nor U10840 (N_10840,N_8853,N_9080);
and U10841 (N_10841,N_8931,N_6397);
and U10842 (N_10842,N_7563,N_8497);
and U10843 (N_10843,N_8998,N_7501);
nor U10844 (N_10844,N_8511,N_8093);
nand U10845 (N_10845,N_6895,N_7905);
or U10846 (N_10846,N_8757,N_8603);
nor U10847 (N_10847,N_6310,N_9241);
nand U10848 (N_10848,N_9352,N_8708);
nand U10849 (N_10849,N_8507,N_7757);
and U10850 (N_10850,N_8642,N_8387);
nand U10851 (N_10851,N_9124,N_6968);
nand U10852 (N_10852,N_6517,N_7605);
xor U10853 (N_10853,N_8413,N_7063);
nor U10854 (N_10854,N_6295,N_6943);
nand U10855 (N_10855,N_6761,N_8473);
xnor U10856 (N_10856,N_7351,N_7641);
xnor U10857 (N_10857,N_7433,N_8299);
and U10858 (N_10858,N_7425,N_7171);
and U10859 (N_10859,N_8032,N_7448);
nand U10860 (N_10860,N_7972,N_7493);
or U10861 (N_10861,N_6638,N_7458);
or U10862 (N_10862,N_7539,N_6700);
or U10863 (N_10863,N_7637,N_8037);
or U10864 (N_10864,N_7405,N_7102);
nor U10865 (N_10865,N_6961,N_8622);
nand U10866 (N_10866,N_7376,N_8375);
or U10867 (N_10867,N_6999,N_7709);
or U10868 (N_10868,N_7643,N_7983);
xor U10869 (N_10869,N_7165,N_7313);
or U10870 (N_10870,N_9205,N_6339);
nor U10871 (N_10871,N_8551,N_6631);
nor U10872 (N_10872,N_8541,N_8188);
and U10873 (N_10873,N_8203,N_6854);
and U10874 (N_10874,N_8385,N_6789);
nor U10875 (N_10875,N_8446,N_7559);
and U10876 (N_10876,N_6544,N_9308);
nor U10877 (N_10877,N_7585,N_6415);
and U10878 (N_10878,N_7569,N_8067);
nor U10879 (N_10879,N_9320,N_7750);
nor U10880 (N_10880,N_8022,N_9082);
and U10881 (N_10881,N_8236,N_9212);
nor U10882 (N_10882,N_7656,N_8417);
nor U10883 (N_10883,N_6929,N_8495);
nor U10884 (N_10884,N_9029,N_7978);
nor U10885 (N_10885,N_6446,N_7714);
and U10886 (N_10886,N_8966,N_7642);
or U10887 (N_10887,N_7604,N_9054);
xnor U10888 (N_10888,N_6971,N_6760);
xor U10889 (N_10889,N_6964,N_7113);
or U10890 (N_10890,N_7331,N_8348);
nand U10891 (N_10891,N_7326,N_9194);
or U10892 (N_10892,N_8210,N_8406);
and U10893 (N_10893,N_8632,N_7655);
nand U10894 (N_10894,N_7084,N_6269);
nor U10895 (N_10895,N_8217,N_8693);
nand U10896 (N_10896,N_7321,N_8763);
xnor U10897 (N_10897,N_6551,N_6515);
and U10898 (N_10898,N_7194,N_7375);
xnor U10899 (N_10899,N_9141,N_6270);
or U10900 (N_10900,N_6652,N_8201);
nand U10901 (N_10901,N_8323,N_6887);
xor U10902 (N_10902,N_8048,N_6326);
nand U10903 (N_10903,N_8835,N_8027);
nand U10904 (N_10904,N_9005,N_7835);
and U10905 (N_10905,N_7209,N_6274);
and U10906 (N_10906,N_6413,N_6754);
or U10907 (N_10907,N_9026,N_8600);
nand U10908 (N_10908,N_8607,N_7332);
xnor U10909 (N_10909,N_7804,N_7472);
nand U10910 (N_10910,N_6753,N_7668);
nor U10911 (N_10911,N_8605,N_9228);
nor U10912 (N_10912,N_6430,N_7339);
or U10913 (N_10913,N_9031,N_7136);
xnor U10914 (N_10914,N_6679,N_8249);
nor U10915 (N_10915,N_6682,N_9269);
xnor U10916 (N_10916,N_7628,N_6324);
nor U10917 (N_10917,N_6656,N_7160);
or U10918 (N_10918,N_6956,N_8091);
nor U10919 (N_10919,N_6578,N_6831);
or U10920 (N_10920,N_7320,N_8177);
nor U10921 (N_10921,N_7015,N_6845);
xor U10922 (N_10922,N_6726,N_7536);
nor U10923 (N_10923,N_6538,N_6952);
nor U10924 (N_10924,N_7096,N_8746);
xnor U10925 (N_10925,N_8072,N_6594);
nand U10926 (N_10926,N_7280,N_6331);
and U10927 (N_10927,N_7296,N_8252);
nand U10928 (N_10928,N_7097,N_8168);
or U10929 (N_10929,N_7450,N_8359);
xor U10930 (N_10930,N_7644,N_7566);
nand U10931 (N_10931,N_9359,N_8974);
nor U10932 (N_10932,N_6378,N_9167);
nor U10933 (N_10933,N_8734,N_9066);
nor U10934 (N_10934,N_7276,N_8847);
or U10935 (N_10935,N_6744,N_8628);
nand U10936 (N_10936,N_6698,N_6408);
and U10937 (N_10937,N_6846,N_8142);
nand U10938 (N_10938,N_8911,N_8348);
nand U10939 (N_10939,N_7162,N_6751);
nand U10940 (N_10940,N_7098,N_7422);
nand U10941 (N_10941,N_8877,N_7761);
xnor U10942 (N_10942,N_8702,N_9280);
xnor U10943 (N_10943,N_7416,N_6657);
xor U10944 (N_10944,N_7808,N_8081);
or U10945 (N_10945,N_8464,N_8987);
nand U10946 (N_10946,N_6865,N_6930);
or U10947 (N_10947,N_8851,N_9134);
xnor U10948 (N_10948,N_8826,N_8356);
nor U10949 (N_10949,N_9044,N_6369);
nor U10950 (N_10950,N_7105,N_8911);
nand U10951 (N_10951,N_8910,N_6864);
xor U10952 (N_10952,N_8185,N_6896);
nand U10953 (N_10953,N_7199,N_8321);
xor U10954 (N_10954,N_9207,N_8687);
or U10955 (N_10955,N_7047,N_8266);
xnor U10956 (N_10956,N_8952,N_7051);
and U10957 (N_10957,N_7062,N_8282);
and U10958 (N_10958,N_8662,N_7806);
or U10959 (N_10959,N_6833,N_8061);
nor U10960 (N_10960,N_6344,N_9187);
and U10961 (N_10961,N_7291,N_7743);
nor U10962 (N_10962,N_9306,N_6397);
nor U10963 (N_10963,N_6934,N_6608);
or U10964 (N_10964,N_8513,N_6435);
nand U10965 (N_10965,N_8332,N_8393);
nand U10966 (N_10966,N_7129,N_7457);
xnor U10967 (N_10967,N_6364,N_6323);
nand U10968 (N_10968,N_6550,N_7616);
and U10969 (N_10969,N_9168,N_7593);
or U10970 (N_10970,N_7460,N_9217);
or U10971 (N_10971,N_8981,N_9180);
or U10972 (N_10972,N_9258,N_6343);
xor U10973 (N_10973,N_7613,N_6377);
or U10974 (N_10974,N_7306,N_8190);
nor U10975 (N_10975,N_6355,N_9050);
or U10976 (N_10976,N_6948,N_6283);
nand U10977 (N_10977,N_6253,N_7351);
nor U10978 (N_10978,N_8064,N_7027);
nor U10979 (N_10979,N_8210,N_6766);
or U10980 (N_10980,N_8442,N_7682);
xnor U10981 (N_10981,N_6763,N_8112);
nor U10982 (N_10982,N_8090,N_8638);
xnor U10983 (N_10983,N_6422,N_6288);
nand U10984 (N_10984,N_8947,N_7273);
and U10985 (N_10985,N_8489,N_8780);
xor U10986 (N_10986,N_6389,N_7983);
and U10987 (N_10987,N_6644,N_8979);
or U10988 (N_10988,N_8525,N_9075);
xnor U10989 (N_10989,N_9118,N_7313);
nor U10990 (N_10990,N_6871,N_6643);
nor U10991 (N_10991,N_6991,N_9038);
nor U10992 (N_10992,N_8377,N_8052);
xnor U10993 (N_10993,N_7653,N_9183);
nand U10994 (N_10994,N_7853,N_6897);
nor U10995 (N_10995,N_8085,N_7965);
and U10996 (N_10996,N_8483,N_8402);
xnor U10997 (N_10997,N_8775,N_8951);
and U10998 (N_10998,N_6747,N_8720);
nor U10999 (N_10999,N_6433,N_7022);
nand U11000 (N_11000,N_9328,N_9092);
xnor U11001 (N_11001,N_8215,N_8239);
and U11002 (N_11002,N_6825,N_8157);
xnor U11003 (N_11003,N_8988,N_6625);
xnor U11004 (N_11004,N_6574,N_6420);
or U11005 (N_11005,N_8645,N_6983);
xnor U11006 (N_11006,N_9014,N_6333);
or U11007 (N_11007,N_6395,N_9084);
nor U11008 (N_11008,N_7133,N_7252);
nand U11009 (N_11009,N_7320,N_8129);
nor U11010 (N_11010,N_7792,N_7427);
nand U11011 (N_11011,N_7819,N_8092);
nor U11012 (N_11012,N_6766,N_7431);
or U11013 (N_11013,N_6897,N_7220);
xor U11014 (N_11014,N_7787,N_6786);
or U11015 (N_11015,N_7876,N_7905);
or U11016 (N_11016,N_6872,N_8695);
and U11017 (N_11017,N_8471,N_6315);
nand U11018 (N_11018,N_8860,N_7844);
or U11019 (N_11019,N_9298,N_8025);
xnor U11020 (N_11020,N_9185,N_8762);
and U11021 (N_11021,N_6346,N_7251);
nor U11022 (N_11022,N_8328,N_6630);
nand U11023 (N_11023,N_8390,N_8797);
nor U11024 (N_11024,N_8662,N_9180);
xnor U11025 (N_11025,N_6529,N_7431);
nand U11026 (N_11026,N_8479,N_8759);
and U11027 (N_11027,N_6619,N_8258);
and U11028 (N_11028,N_8614,N_7721);
nor U11029 (N_11029,N_7700,N_6254);
nor U11030 (N_11030,N_7795,N_8571);
and U11031 (N_11031,N_8611,N_8869);
or U11032 (N_11032,N_6867,N_8912);
xor U11033 (N_11033,N_8113,N_6477);
nor U11034 (N_11034,N_7592,N_7903);
xnor U11035 (N_11035,N_8515,N_7266);
xor U11036 (N_11036,N_7167,N_9275);
and U11037 (N_11037,N_7398,N_7277);
or U11038 (N_11038,N_6893,N_8754);
nor U11039 (N_11039,N_7915,N_6987);
nand U11040 (N_11040,N_7003,N_7102);
nor U11041 (N_11041,N_6739,N_6898);
nor U11042 (N_11042,N_6253,N_7816);
xnor U11043 (N_11043,N_8661,N_8000);
or U11044 (N_11044,N_9231,N_9073);
or U11045 (N_11045,N_8104,N_8554);
xor U11046 (N_11046,N_6317,N_6657);
xor U11047 (N_11047,N_8648,N_7830);
xnor U11048 (N_11048,N_6507,N_7900);
nand U11049 (N_11049,N_9193,N_9103);
nor U11050 (N_11050,N_8111,N_8214);
nand U11051 (N_11051,N_6928,N_8275);
or U11052 (N_11052,N_6418,N_7260);
or U11053 (N_11053,N_7847,N_6526);
nand U11054 (N_11054,N_7754,N_8978);
or U11055 (N_11055,N_7963,N_8230);
and U11056 (N_11056,N_6974,N_9263);
xnor U11057 (N_11057,N_6465,N_7648);
or U11058 (N_11058,N_7915,N_9222);
nand U11059 (N_11059,N_9056,N_7735);
xnor U11060 (N_11060,N_8382,N_9278);
nand U11061 (N_11061,N_8703,N_9097);
nor U11062 (N_11062,N_8927,N_7409);
or U11063 (N_11063,N_7364,N_7785);
nor U11064 (N_11064,N_6791,N_7466);
or U11065 (N_11065,N_8750,N_9358);
and U11066 (N_11066,N_7389,N_7992);
and U11067 (N_11067,N_7544,N_8309);
xnor U11068 (N_11068,N_6815,N_9322);
nand U11069 (N_11069,N_7017,N_8728);
nand U11070 (N_11070,N_7543,N_6814);
nand U11071 (N_11071,N_7530,N_9204);
and U11072 (N_11072,N_6732,N_6761);
xnor U11073 (N_11073,N_7207,N_8443);
or U11074 (N_11074,N_8599,N_8433);
or U11075 (N_11075,N_9032,N_6597);
nand U11076 (N_11076,N_6845,N_7145);
nand U11077 (N_11077,N_8316,N_8411);
nand U11078 (N_11078,N_7722,N_8870);
and U11079 (N_11079,N_8993,N_7171);
nor U11080 (N_11080,N_6877,N_6844);
nor U11081 (N_11081,N_7963,N_7944);
xnor U11082 (N_11082,N_7246,N_8330);
nand U11083 (N_11083,N_7897,N_8608);
and U11084 (N_11084,N_7839,N_7828);
or U11085 (N_11085,N_6563,N_9355);
nor U11086 (N_11086,N_6408,N_6543);
nand U11087 (N_11087,N_8166,N_6986);
and U11088 (N_11088,N_8005,N_6662);
nand U11089 (N_11089,N_7608,N_7571);
or U11090 (N_11090,N_8001,N_7178);
and U11091 (N_11091,N_8113,N_6363);
xnor U11092 (N_11092,N_8881,N_7573);
nand U11093 (N_11093,N_7485,N_8606);
xnor U11094 (N_11094,N_8404,N_8792);
or U11095 (N_11095,N_8839,N_7641);
nand U11096 (N_11096,N_8727,N_7411);
and U11097 (N_11097,N_7404,N_8509);
nor U11098 (N_11098,N_6958,N_6570);
and U11099 (N_11099,N_8959,N_7972);
nand U11100 (N_11100,N_6750,N_6940);
nand U11101 (N_11101,N_8152,N_7757);
nor U11102 (N_11102,N_9094,N_7623);
nor U11103 (N_11103,N_6855,N_7021);
or U11104 (N_11104,N_7265,N_9248);
nor U11105 (N_11105,N_6857,N_6391);
and U11106 (N_11106,N_7057,N_8989);
nand U11107 (N_11107,N_9147,N_8136);
nand U11108 (N_11108,N_9091,N_8901);
nand U11109 (N_11109,N_6983,N_8349);
nor U11110 (N_11110,N_7336,N_8341);
or U11111 (N_11111,N_9063,N_7968);
xnor U11112 (N_11112,N_9336,N_8018);
or U11113 (N_11113,N_7090,N_7514);
xor U11114 (N_11114,N_8485,N_7616);
and U11115 (N_11115,N_9047,N_6996);
xnor U11116 (N_11116,N_8978,N_6952);
or U11117 (N_11117,N_8929,N_8979);
nand U11118 (N_11118,N_7651,N_8649);
nand U11119 (N_11119,N_7741,N_6723);
xor U11120 (N_11120,N_8716,N_8682);
nor U11121 (N_11121,N_7134,N_9266);
xnor U11122 (N_11122,N_7286,N_7784);
nor U11123 (N_11123,N_7988,N_8067);
and U11124 (N_11124,N_7220,N_8758);
or U11125 (N_11125,N_7355,N_8847);
nor U11126 (N_11126,N_8084,N_7514);
and U11127 (N_11127,N_7191,N_9119);
or U11128 (N_11128,N_8544,N_6374);
and U11129 (N_11129,N_6268,N_7627);
or U11130 (N_11130,N_7799,N_8085);
or U11131 (N_11131,N_8532,N_6991);
and U11132 (N_11132,N_8332,N_7038);
xnor U11133 (N_11133,N_9120,N_6689);
nor U11134 (N_11134,N_8933,N_8536);
or U11135 (N_11135,N_9174,N_7758);
xor U11136 (N_11136,N_9308,N_6966);
and U11137 (N_11137,N_7026,N_7877);
nand U11138 (N_11138,N_7169,N_7369);
nor U11139 (N_11139,N_8313,N_7637);
and U11140 (N_11140,N_6581,N_8203);
nand U11141 (N_11141,N_6880,N_6441);
xor U11142 (N_11142,N_6851,N_6760);
or U11143 (N_11143,N_8434,N_6885);
nor U11144 (N_11144,N_6935,N_8538);
and U11145 (N_11145,N_6255,N_8765);
nor U11146 (N_11146,N_8234,N_7692);
nand U11147 (N_11147,N_7156,N_6370);
nand U11148 (N_11148,N_8118,N_9256);
nor U11149 (N_11149,N_6468,N_7007);
nor U11150 (N_11150,N_6273,N_6948);
xnor U11151 (N_11151,N_8603,N_7951);
nand U11152 (N_11152,N_7414,N_8965);
nand U11153 (N_11153,N_8159,N_6555);
and U11154 (N_11154,N_8061,N_6933);
or U11155 (N_11155,N_7265,N_7837);
or U11156 (N_11156,N_6764,N_7950);
or U11157 (N_11157,N_7993,N_6691);
or U11158 (N_11158,N_7522,N_7376);
nand U11159 (N_11159,N_9295,N_7515);
nand U11160 (N_11160,N_7063,N_9370);
xnor U11161 (N_11161,N_8860,N_7383);
nand U11162 (N_11162,N_7316,N_6473);
nor U11163 (N_11163,N_8837,N_9321);
and U11164 (N_11164,N_6900,N_7859);
and U11165 (N_11165,N_7718,N_7662);
or U11166 (N_11166,N_6455,N_6260);
xnor U11167 (N_11167,N_7339,N_7776);
xnor U11168 (N_11168,N_6887,N_6733);
and U11169 (N_11169,N_7728,N_6501);
nor U11170 (N_11170,N_8572,N_6606);
or U11171 (N_11171,N_8374,N_8539);
xnor U11172 (N_11172,N_6704,N_8765);
nand U11173 (N_11173,N_7156,N_8770);
and U11174 (N_11174,N_7744,N_8189);
and U11175 (N_11175,N_8461,N_7791);
and U11176 (N_11176,N_7081,N_8111);
and U11177 (N_11177,N_9260,N_8874);
or U11178 (N_11178,N_8338,N_9086);
nand U11179 (N_11179,N_7262,N_9159);
nor U11180 (N_11180,N_6552,N_7119);
and U11181 (N_11181,N_7708,N_6677);
nand U11182 (N_11182,N_9256,N_8889);
and U11183 (N_11183,N_8626,N_6480);
and U11184 (N_11184,N_7589,N_6525);
or U11185 (N_11185,N_7529,N_7155);
xor U11186 (N_11186,N_7500,N_6672);
or U11187 (N_11187,N_8473,N_8572);
xor U11188 (N_11188,N_8957,N_6734);
nand U11189 (N_11189,N_9079,N_8686);
and U11190 (N_11190,N_8821,N_6653);
xnor U11191 (N_11191,N_8541,N_8917);
and U11192 (N_11192,N_8549,N_7495);
xor U11193 (N_11193,N_6820,N_8865);
xnor U11194 (N_11194,N_8421,N_8262);
nand U11195 (N_11195,N_7543,N_7831);
nand U11196 (N_11196,N_8791,N_9288);
nor U11197 (N_11197,N_8691,N_8873);
and U11198 (N_11198,N_8280,N_7043);
nor U11199 (N_11199,N_8327,N_7294);
xor U11200 (N_11200,N_8287,N_6737);
xnor U11201 (N_11201,N_6828,N_8075);
or U11202 (N_11202,N_7667,N_6352);
and U11203 (N_11203,N_6623,N_9342);
nand U11204 (N_11204,N_7566,N_8353);
and U11205 (N_11205,N_6894,N_6502);
and U11206 (N_11206,N_7717,N_6738);
or U11207 (N_11207,N_8053,N_7170);
nor U11208 (N_11208,N_6700,N_7413);
nor U11209 (N_11209,N_8971,N_6498);
and U11210 (N_11210,N_6888,N_8666);
nand U11211 (N_11211,N_8089,N_9308);
or U11212 (N_11212,N_7098,N_9082);
and U11213 (N_11213,N_7320,N_7793);
xnor U11214 (N_11214,N_7183,N_7604);
xnor U11215 (N_11215,N_7940,N_7067);
or U11216 (N_11216,N_8943,N_8317);
xor U11217 (N_11217,N_8057,N_9298);
or U11218 (N_11218,N_8018,N_7035);
xnor U11219 (N_11219,N_8395,N_8324);
nand U11220 (N_11220,N_6491,N_8605);
nor U11221 (N_11221,N_9129,N_7391);
or U11222 (N_11222,N_7841,N_8932);
nor U11223 (N_11223,N_7835,N_9053);
or U11224 (N_11224,N_7936,N_8980);
and U11225 (N_11225,N_8550,N_7946);
nor U11226 (N_11226,N_6315,N_6528);
or U11227 (N_11227,N_6773,N_9257);
or U11228 (N_11228,N_7659,N_8605);
and U11229 (N_11229,N_7716,N_8634);
nor U11230 (N_11230,N_7543,N_8968);
nor U11231 (N_11231,N_7923,N_6318);
nor U11232 (N_11232,N_6849,N_8574);
xnor U11233 (N_11233,N_9238,N_6468);
nand U11234 (N_11234,N_6459,N_8849);
and U11235 (N_11235,N_6692,N_9259);
xnor U11236 (N_11236,N_7796,N_9103);
xor U11237 (N_11237,N_7177,N_7729);
and U11238 (N_11238,N_6477,N_6560);
nand U11239 (N_11239,N_7673,N_7622);
nand U11240 (N_11240,N_6496,N_9074);
nor U11241 (N_11241,N_7667,N_9326);
nor U11242 (N_11242,N_8616,N_7700);
xor U11243 (N_11243,N_7982,N_6950);
xnor U11244 (N_11244,N_8454,N_7254);
nor U11245 (N_11245,N_8113,N_7065);
xor U11246 (N_11246,N_6523,N_6819);
or U11247 (N_11247,N_8414,N_6685);
or U11248 (N_11248,N_8350,N_8767);
xor U11249 (N_11249,N_8923,N_6411);
nor U11250 (N_11250,N_9308,N_8862);
xnor U11251 (N_11251,N_7495,N_6814);
and U11252 (N_11252,N_9249,N_7950);
or U11253 (N_11253,N_9041,N_7858);
nor U11254 (N_11254,N_7836,N_8435);
and U11255 (N_11255,N_6706,N_8673);
and U11256 (N_11256,N_9056,N_6307);
xor U11257 (N_11257,N_8725,N_6557);
nor U11258 (N_11258,N_7365,N_8896);
or U11259 (N_11259,N_6811,N_8628);
and U11260 (N_11260,N_6837,N_9350);
and U11261 (N_11261,N_8332,N_6606);
xnor U11262 (N_11262,N_8008,N_8932);
nor U11263 (N_11263,N_8093,N_9254);
or U11264 (N_11264,N_7061,N_6402);
nor U11265 (N_11265,N_7254,N_9046);
nor U11266 (N_11266,N_7513,N_6292);
xor U11267 (N_11267,N_9114,N_9310);
or U11268 (N_11268,N_9277,N_8295);
nor U11269 (N_11269,N_9048,N_8471);
nor U11270 (N_11270,N_6661,N_9122);
nor U11271 (N_11271,N_8835,N_7938);
xor U11272 (N_11272,N_7539,N_8418);
and U11273 (N_11273,N_8618,N_8965);
nor U11274 (N_11274,N_9334,N_8833);
xor U11275 (N_11275,N_9203,N_7423);
xor U11276 (N_11276,N_8853,N_7034);
nor U11277 (N_11277,N_8342,N_6537);
nor U11278 (N_11278,N_7989,N_6764);
and U11279 (N_11279,N_8171,N_9092);
nand U11280 (N_11280,N_7035,N_6646);
and U11281 (N_11281,N_6540,N_6915);
or U11282 (N_11282,N_6495,N_7421);
nor U11283 (N_11283,N_9074,N_9157);
xnor U11284 (N_11284,N_8987,N_8754);
or U11285 (N_11285,N_6633,N_8648);
or U11286 (N_11286,N_9138,N_7241);
or U11287 (N_11287,N_8182,N_8199);
nand U11288 (N_11288,N_7811,N_6784);
nand U11289 (N_11289,N_6999,N_6462);
nand U11290 (N_11290,N_7791,N_6928);
xnor U11291 (N_11291,N_9282,N_8186);
and U11292 (N_11292,N_7122,N_9259);
or U11293 (N_11293,N_7898,N_9346);
and U11294 (N_11294,N_9261,N_9314);
nand U11295 (N_11295,N_7115,N_9001);
or U11296 (N_11296,N_8725,N_7142);
or U11297 (N_11297,N_7879,N_8804);
nor U11298 (N_11298,N_8414,N_7272);
nor U11299 (N_11299,N_7533,N_8794);
or U11300 (N_11300,N_7716,N_6755);
and U11301 (N_11301,N_8157,N_7079);
nor U11302 (N_11302,N_6369,N_6884);
or U11303 (N_11303,N_6791,N_6698);
nand U11304 (N_11304,N_9113,N_8164);
nand U11305 (N_11305,N_9291,N_7472);
and U11306 (N_11306,N_8365,N_9361);
xnor U11307 (N_11307,N_8986,N_7079);
nand U11308 (N_11308,N_6645,N_8788);
and U11309 (N_11309,N_7177,N_9115);
or U11310 (N_11310,N_9232,N_7621);
and U11311 (N_11311,N_7409,N_8195);
nor U11312 (N_11312,N_8467,N_7627);
xor U11313 (N_11313,N_7370,N_9092);
and U11314 (N_11314,N_8871,N_9156);
xor U11315 (N_11315,N_8022,N_7413);
and U11316 (N_11316,N_8259,N_6943);
nor U11317 (N_11317,N_7010,N_8092);
xor U11318 (N_11318,N_8817,N_8206);
nand U11319 (N_11319,N_9175,N_7121);
nand U11320 (N_11320,N_8285,N_6746);
nor U11321 (N_11321,N_7673,N_8800);
nand U11322 (N_11322,N_7530,N_8731);
xnor U11323 (N_11323,N_8925,N_8485);
xnor U11324 (N_11324,N_8690,N_9128);
and U11325 (N_11325,N_8977,N_8882);
and U11326 (N_11326,N_7070,N_9117);
and U11327 (N_11327,N_9090,N_7683);
and U11328 (N_11328,N_8447,N_8156);
nand U11329 (N_11329,N_8814,N_7878);
and U11330 (N_11330,N_9198,N_8589);
xor U11331 (N_11331,N_7650,N_8349);
nand U11332 (N_11332,N_7206,N_7021);
nor U11333 (N_11333,N_6517,N_8837);
and U11334 (N_11334,N_6280,N_9181);
and U11335 (N_11335,N_7702,N_6337);
or U11336 (N_11336,N_6566,N_8049);
xor U11337 (N_11337,N_6470,N_8588);
xor U11338 (N_11338,N_7227,N_8572);
nand U11339 (N_11339,N_6920,N_8960);
nor U11340 (N_11340,N_7392,N_9306);
and U11341 (N_11341,N_9217,N_7626);
xor U11342 (N_11342,N_8002,N_7899);
nand U11343 (N_11343,N_9311,N_8938);
or U11344 (N_11344,N_8359,N_9284);
nand U11345 (N_11345,N_6575,N_7923);
xor U11346 (N_11346,N_7650,N_7850);
xnor U11347 (N_11347,N_8504,N_6799);
or U11348 (N_11348,N_8093,N_8139);
and U11349 (N_11349,N_9342,N_6496);
and U11350 (N_11350,N_8656,N_7402);
and U11351 (N_11351,N_6911,N_9029);
xor U11352 (N_11352,N_9184,N_6278);
xor U11353 (N_11353,N_6662,N_9192);
or U11354 (N_11354,N_6303,N_6794);
and U11355 (N_11355,N_7325,N_9286);
or U11356 (N_11356,N_7475,N_7007);
and U11357 (N_11357,N_9089,N_6734);
nor U11358 (N_11358,N_7656,N_9096);
nor U11359 (N_11359,N_9327,N_9088);
xor U11360 (N_11360,N_7122,N_8114);
nand U11361 (N_11361,N_9344,N_7128);
or U11362 (N_11362,N_7339,N_7597);
and U11363 (N_11363,N_7832,N_8783);
or U11364 (N_11364,N_6874,N_7627);
or U11365 (N_11365,N_7820,N_6377);
and U11366 (N_11366,N_9189,N_9045);
and U11367 (N_11367,N_9143,N_8762);
nand U11368 (N_11368,N_8772,N_7451);
xor U11369 (N_11369,N_8135,N_7480);
nor U11370 (N_11370,N_7097,N_8523);
and U11371 (N_11371,N_8642,N_8550);
xnor U11372 (N_11372,N_8391,N_9078);
and U11373 (N_11373,N_7993,N_9111);
nor U11374 (N_11374,N_6809,N_7067);
and U11375 (N_11375,N_9137,N_6975);
xnor U11376 (N_11376,N_8474,N_7478);
nor U11377 (N_11377,N_7010,N_8375);
or U11378 (N_11378,N_7333,N_7707);
nand U11379 (N_11379,N_6766,N_8391);
nand U11380 (N_11380,N_6783,N_7041);
or U11381 (N_11381,N_7192,N_8122);
or U11382 (N_11382,N_7030,N_8468);
or U11383 (N_11383,N_7155,N_8071);
and U11384 (N_11384,N_7206,N_6991);
nor U11385 (N_11385,N_8314,N_9102);
nor U11386 (N_11386,N_7837,N_6874);
xnor U11387 (N_11387,N_7931,N_9282);
nor U11388 (N_11388,N_8656,N_7671);
nand U11389 (N_11389,N_9218,N_8899);
xnor U11390 (N_11390,N_6257,N_8187);
and U11391 (N_11391,N_6299,N_8306);
nor U11392 (N_11392,N_7747,N_8278);
xor U11393 (N_11393,N_6612,N_7015);
and U11394 (N_11394,N_9018,N_6442);
xnor U11395 (N_11395,N_6994,N_9028);
nor U11396 (N_11396,N_8187,N_7181);
nand U11397 (N_11397,N_6933,N_7923);
nor U11398 (N_11398,N_8422,N_7800);
or U11399 (N_11399,N_7875,N_8358);
or U11400 (N_11400,N_6929,N_7002);
xnor U11401 (N_11401,N_7999,N_7788);
nor U11402 (N_11402,N_7472,N_6266);
or U11403 (N_11403,N_8293,N_6681);
nor U11404 (N_11404,N_7885,N_6714);
xor U11405 (N_11405,N_7960,N_8238);
nor U11406 (N_11406,N_9153,N_7164);
nor U11407 (N_11407,N_8055,N_8764);
xnor U11408 (N_11408,N_8836,N_6423);
and U11409 (N_11409,N_8161,N_6951);
or U11410 (N_11410,N_8305,N_8841);
nand U11411 (N_11411,N_8350,N_9268);
and U11412 (N_11412,N_7446,N_6927);
xnor U11413 (N_11413,N_7989,N_7080);
and U11414 (N_11414,N_8776,N_8398);
xor U11415 (N_11415,N_8788,N_6707);
nand U11416 (N_11416,N_7070,N_7244);
and U11417 (N_11417,N_9371,N_9196);
nand U11418 (N_11418,N_8790,N_8216);
or U11419 (N_11419,N_8211,N_7026);
and U11420 (N_11420,N_8307,N_9317);
xnor U11421 (N_11421,N_9190,N_6674);
or U11422 (N_11422,N_6916,N_7776);
and U11423 (N_11423,N_8758,N_9245);
nor U11424 (N_11424,N_8557,N_8932);
and U11425 (N_11425,N_6853,N_7870);
or U11426 (N_11426,N_9304,N_6545);
or U11427 (N_11427,N_8190,N_8273);
and U11428 (N_11428,N_8912,N_7899);
and U11429 (N_11429,N_7315,N_6814);
nor U11430 (N_11430,N_6514,N_7475);
or U11431 (N_11431,N_7087,N_7242);
xnor U11432 (N_11432,N_7137,N_7903);
and U11433 (N_11433,N_6573,N_8496);
nand U11434 (N_11434,N_7718,N_7937);
xnor U11435 (N_11435,N_8448,N_6521);
nor U11436 (N_11436,N_8449,N_6416);
nand U11437 (N_11437,N_6616,N_6397);
nand U11438 (N_11438,N_8340,N_8969);
xnor U11439 (N_11439,N_8967,N_6687);
nor U11440 (N_11440,N_6355,N_9049);
or U11441 (N_11441,N_7833,N_6553);
and U11442 (N_11442,N_7905,N_9238);
xor U11443 (N_11443,N_8608,N_7525);
or U11444 (N_11444,N_6920,N_8561);
or U11445 (N_11445,N_9256,N_9000);
xnor U11446 (N_11446,N_6596,N_7458);
and U11447 (N_11447,N_8191,N_9092);
or U11448 (N_11448,N_8651,N_7166);
nand U11449 (N_11449,N_6419,N_7487);
nor U11450 (N_11450,N_8595,N_9045);
nor U11451 (N_11451,N_7706,N_8367);
or U11452 (N_11452,N_8528,N_7007);
nor U11453 (N_11453,N_7832,N_6572);
or U11454 (N_11454,N_8771,N_8512);
nand U11455 (N_11455,N_9125,N_8177);
or U11456 (N_11456,N_6759,N_6557);
xor U11457 (N_11457,N_8268,N_8183);
nand U11458 (N_11458,N_6520,N_8030);
xor U11459 (N_11459,N_7760,N_6293);
xor U11460 (N_11460,N_8439,N_6407);
xnor U11461 (N_11461,N_7357,N_6625);
nand U11462 (N_11462,N_7432,N_8278);
and U11463 (N_11463,N_7512,N_8420);
nor U11464 (N_11464,N_6521,N_6834);
xor U11465 (N_11465,N_7632,N_7733);
nand U11466 (N_11466,N_7875,N_6491);
and U11467 (N_11467,N_8985,N_6543);
or U11468 (N_11468,N_9348,N_7559);
nor U11469 (N_11469,N_8080,N_8410);
or U11470 (N_11470,N_9206,N_7709);
xnor U11471 (N_11471,N_8612,N_9194);
xnor U11472 (N_11472,N_8579,N_9282);
nor U11473 (N_11473,N_7776,N_8574);
and U11474 (N_11474,N_9269,N_6749);
xnor U11475 (N_11475,N_7232,N_6936);
nand U11476 (N_11476,N_7856,N_8328);
nand U11477 (N_11477,N_7751,N_6340);
nor U11478 (N_11478,N_6599,N_7732);
nor U11479 (N_11479,N_8961,N_6934);
xnor U11480 (N_11480,N_7238,N_9182);
nor U11481 (N_11481,N_8303,N_7426);
nand U11482 (N_11482,N_7406,N_7056);
nor U11483 (N_11483,N_7272,N_6792);
nor U11484 (N_11484,N_8181,N_7470);
nor U11485 (N_11485,N_7740,N_7403);
or U11486 (N_11486,N_6560,N_8679);
xor U11487 (N_11487,N_6721,N_7014);
xor U11488 (N_11488,N_8412,N_6583);
and U11489 (N_11489,N_7786,N_8421);
xor U11490 (N_11490,N_8719,N_9158);
and U11491 (N_11491,N_7545,N_7127);
xor U11492 (N_11492,N_7521,N_6946);
nor U11493 (N_11493,N_6728,N_8144);
nand U11494 (N_11494,N_6796,N_7800);
nor U11495 (N_11495,N_8035,N_7636);
nand U11496 (N_11496,N_6816,N_8840);
nand U11497 (N_11497,N_6620,N_8643);
nor U11498 (N_11498,N_6363,N_7517);
nand U11499 (N_11499,N_7780,N_6469);
or U11500 (N_11500,N_8931,N_7628);
nor U11501 (N_11501,N_9298,N_8653);
nand U11502 (N_11502,N_7317,N_7670);
nand U11503 (N_11503,N_9308,N_6646);
nor U11504 (N_11504,N_8497,N_7496);
nand U11505 (N_11505,N_9257,N_6441);
xnor U11506 (N_11506,N_9165,N_7534);
nor U11507 (N_11507,N_8775,N_8229);
or U11508 (N_11508,N_7853,N_9121);
and U11509 (N_11509,N_7427,N_7451);
and U11510 (N_11510,N_6611,N_6968);
nand U11511 (N_11511,N_8821,N_6275);
and U11512 (N_11512,N_8404,N_6734);
and U11513 (N_11513,N_6267,N_9107);
nor U11514 (N_11514,N_9306,N_8147);
nand U11515 (N_11515,N_8821,N_7229);
and U11516 (N_11516,N_8498,N_7855);
nand U11517 (N_11517,N_6696,N_6710);
and U11518 (N_11518,N_7150,N_7411);
nor U11519 (N_11519,N_8142,N_9302);
and U11520 (N_11520,N_6384,N_8598);
xnor U11521 (N_11521,N_6925,N_7417);
or U11522 (N_11522,N_8038,N_8405);
nor U11523 (N_11523,N_6341,N_8569);
nand U11524 (N_11524,N_8444,N_7386);
and U11525 (N_11525,N_8413,N_7192);
nor U11526 (N_11526,N_6627,N_8348);
nand U11527 (N_11527,N_7141,N_6694);
xnor U11528 (N_11528,N_8381,N_9328);
nor U11529 (N_11529,N_6561,N_7284);
and U11530 (N_11530,N_6933,N_6752);
and U11531 (N_11531,N_7238,N_8718);
xor U11532 (N_11532,N_8013,N_6272);
nor U11533 (N_11533,N_6501,N_7748);
nor U11534 (N_11534,N_9116,N_6955);
xor U11535 (N_11535,N_7505,N_7695);
nand U11536 (N_11536,N_7189,N_8690);
and U11537 (N_11537,N_8214,N_8901);
or U11538 (N_11538,N_8976,N_8381);
xor U11539 (N_11539,N_8540,N_9145);
nand U11540 (N_11540,N_7267,N_8325);
and U11541 (N_11541,N_6900,N_7731);
nand U11542 (N_11542,N_7351,N_7585);
or U11543 (N_11543,N_6940,N_8817);
and U11544 (N_11544,N_9089,N_9213);
and U11545 (N_11545,N_7544,N_6423);
nor U11546 (N_11546,N_7195,N_8041);
and U11547 (N_11547,N_8185,N_8997);
nand U11548 (N_11548,N_7632,N_8832);
or U11549 (N_11549,N_8900,N_8769);
xnor U11550 (N_11550,N_6998,N_8971);
xor U11551 (N_11551,N_7835,N_6628);
nand U11552 (N_11552,N_7026,N_7618);
nor U11553 (N_11553,N_7388,N_6731);
nor U11554 (N_11554,N_8206,N_7518);
xnor U11555 (N_11555,N_6541,N_8688);
nor U11556 (N_11556,N_9207,N_8824);
nand U11557 (N_11557,N_6559,N_8413);
nand U11558 (N_11558,N_7548,N_8453);
and U11559 (N_11559,N_8847,N_7845);
and U11560 (N_11560,N_7905,N_7544);
and U11561 (N_11561,N_6918,N_8938);
nand U11562 (N_11562,N_7421,N_7827);
nand U11563 (N_11563,N_6541,N_8855);
and U11564 (N_11564,N_7890,N_8173);
and U11565 (N_11565,N_8187,N_9145);
xnor U11566 (N_11566,N_8398,N_6794);
xor U11567 (N_11567,N_8211,N_7558);
xor U11568 (N_11568,N_8385,N_9192);
and U11569 (N_11569,N_9146,N_8133);
xnor U11570 (N_11570,N_7453,N_8129);
xor U11571 (N_11571,N_7511,N_8124);
nand U11572 (N_11572,N_6837,N_7905);
and U11573 (N_11573,N_8186,N_9276);
and U11574 (N_11574,N_7970,N_8169);
nand U11575 (N_11575,N_9223,N_6595);
nor U11576 (N_11576,N_8461,N_8543);
or U11577 (N_11577,N_7496,N_6642);
xnor U11578 (N_11578,N_6351,N_8205);
xor U11579 (N_11579,N_8069,N_6280);
xor U11580 (N_11580,N_8415,N_8887);
xor U11581 (N_11581,N_9016,N_8471);
xor U11582 (N_11582,N_8766,N_7587);
nand U11583 (N_11583,N_7857,N_9103);
nor U11584 (N_11584,N_7771,N_6909);
xnor U11585 (N_11585,N_8807,N_6271);
or U11586 (N_11586,N_7523,N_7816);
nor U11587 (N_11587,N_6717,N_8916);
nor U11588 (N_11588,N_8228,N_6998);
and U11589 (N_11589,N_6853,N_6383);
nand U11590 (N_11590,N_8876,N_7045);
and U11591 (N_11591,N_9361,N_6622);
nor U11592 (N_11592,N_9243,N_8865);
or U11593 (N_11593,N_7113,N_6377);
and U11594 (N_11594,N_7800,N_6358);
xnor U11595 (N_11595,N_7763,N_9098);
or U11596 (N_11596,N_6586,N_7259);
nor U11597 (N_11597,N_7545,N_7936);
or U11598 (N_11598,N_8598,N_9293);
nand U11599 (N_11599,N_8874,N_6746);
nor U11600 (N_11600,N_6689,N_9182);
xor U11601 (N_11601,N_7581,N_9076);
and U11602 (N_11602,N_6974,N_8649);
or U11603 (N_11603,N_9020,N_7945);
xnor U11604 (N_11604,N_8726,N_7944);
nand U11605 (N_11605,N_7976,N_6726);
or U11606 (N_11606,N_8464,N_7085);
nor U11607 (N_11607,N_7807,N_8723);
or U11608 (N_11608,N_7790,N_6565);
nor U11609 (N_11609,N_8285,N_6859);
xor U11610 (N_11610,N_7515,N_7633);
and U11611 (N_11611,N_8543,N_6752);
nor U11612 (N_11612,N_7015,N_7892);
xor U11613 (N_11613,N_6369,N_8600);
xnor U11614 (N_11614,N_7247,N_7196);
xnor U11615 (N_11615,N_8038,N_7732);
or U11616 (N_11616,N_8513,N_7243);
xnor U11617 (N_11617,N_8211,N_9186);
nor U11618 (N_11618,N_7119,N_8137);
nor U11619 (N_11619,N_8622,N_7691);
or U11620 (N_11620,N_6894,N_8040);
nor U11621 (N_11621,N_6769,N_6511);
and U11622 (N_11622,N_8668,N_7697);
nor U11623 (N_11623,N_8545,N_6597);
or U11624 (N_11624,N_7991,N_8555);
nor U11625 (N_11625,N_8507,N_7868);
xnor U11626 (N_11626,N_6421,N_8964);
nor U11627 (N_11627,N_6561,N_7966);
nor U11628 (N_11628,N_7307,N_6403);
nor U11629 (N_11629,N_8973,N_6808);
or U11630 (N_11630,N_6668,N_9294);
and U11631 (N_11631,N_7621,N_6492);
nand U11632 (N_11632,N_7363,N_7725);
nand U11633 (N_11633,N_6940,N_7694);
nor U11634 (N_11634,N_7390,N_8487);
nor U11635 (N_11635,N_7450,N_6743);
xnor U11636 (N_11636,N_9109,N_8360);
xor U11637 (N_11637,N_7293,N_6652);
or U11638 (N_11638,N_7759,N_7029);
and U11639 (N_11639,N_6838,N_9200);
xor U11640 (N_11640,N_6330,N_6585);
xnor U11641 (N_11641,N_6334,N_7200);
nor U11642 (N_11642,N_7230,N_9047);
nand U11643 (N_11643,N_7019,N_7816);
or U11644 (N_11644,N_9319,N_6413);
and U11645 (N_11645,N_7903,N_6881);
nand U11646 (N_11646,N_7378,N_6609);
nand U11647 (N_11647,N_7921,N_8308);
nand U11648 (N_11648,N_8300,N_7866);
or U11649 (N_11649,N_8821,N_6647);
and U11650 (N_11650,N_7285,N_8673);
nand U11651 (N_11651,N_7098,N_8957);
or U11652 (N_11652,N_6908,N_7378);
xor U11653 (N_11653,N_7779,N_9205);
xnor U11654 (N_11654,N_7591,N_8713);
and U11655 (N_11655,N_9057,N_6504);
or U11656 (N_11656,N_6599,N_8224);
nor U11657 (N_11657,N_9202,N_9208);
nor U11658 (N_11658,N_6433,N_8334);
nand U11659 (N_11659,N_6648,N_6325);
nand U11660 (N_11660,N_6859,N_6549);
xnor U11661 (N_11661,N_7731,N_7534);
nand U11662 (N_11662,N_6337,N_6727);
and U11663 (N_11663,N_8305,N_7149);
xor U11664 (N_11664,N_8189,N_6474);
nand U11665 (N_11665,N_6440,N_7603);
nand U11666 (N_11666,N_6502,N_8490);
nand U11667 (N_11667,N_8082,N_8116);
nand U11668 (N_11668,N_8689,N_7959);
nor U11669 (N_11669,N_9125,N_6600);
nor U11670 (N_11670,N_8442,N_7436);
and U11671 (N_11671,N_8714,N_7559);
and U11672 (N_11672,N_8455,N_8414);
nor U11673 (N_11673,N_8152,N_8447);
and U11674 (N_11674,N_9360,N_8641);
or U11675 (N_11675,N_6758,N_6796);
xnor U11676 (N_11676,N_6306,N_7132);
and U11677 (N_11677,N_7542,N_8467);
xor U11678 (N_11678,N_6309,N_8902);
nor U11679 (N_11679,N_6748,N_6790);
and U11680 (N_11680,N_8057,N_8607);
or U11681 (N_11681,N_7345,N_6757);
and U11682 (N_11682,N_8606,N_6602);
and U11683 (N_11683,N_8339,N_8375);
and U11684 (N_11684,N_7059,N_8248);
or U11685 (N_11685,N_7869,N_9205);
or U11686 (N_11686,N_8389,N_8030);
and U11687 (N_11687,N_7232,N_8172);
xnor U11688 (N_11688,N_8516,N_9076);
nor U11689 (N_11689,N_8031,N_6385);
xor U11690 (N_11690,N_8443,N_7775);
xor U11691 (N_11691,N_8501,N_8092);
nand U11692 (N_11692,N_8459,N_9213);
and U11693 (N_11693,N_7265,N_7418);
nor U11694 (N_11694,N_9020,N_8394);
nor U11695 (N_11695,N_6412,N_8573);
or U11696 (N_11696,N_9357,N_8489);
nand U11697 (N_11697,N_6846,N_9001);
nor U11698 (N_11698,N_6259,N_8214);
nand U11699 (N_11699,N_8773,N_7147);
and U11700 (N_11700,N_6427,N_6933);
and U11701 (N_11701,N_7780,N_6572);
nor U11702 (N_11702,N_9050,N_7017);
xor U11703 (N_11703,N_7231,N_7489);
nor U11704 (N_11704,N_8951,N_8755);
nand U11705 (N_11705,N_8186,N_6965);
nor U11706 (N_11706,N_7622,N_7909);
xnor U11707 (N_11707,N_7703,N_6803);
nor U11708 (N_11708,N_7162,N_7366);
nand U11709 (N_11709,N_8640,N_8429);
xor U11710 (N_11710,N_7828,N_7831);
and U11711 (N_11711,N_9293,N_6276);
xor U11712 (N_11712,N_7043,N_9032);
nand U11713 (N_11713,N_7356,N_8470);
xor U11714 (N_11714,N_8699,N_7611);
and U11715 (N_11715,N_6321,N_7664);
and U11716 (N_11716,N_6739,N_7532);
nor U11717 (N_11717,N_7196,N_8071);
and U11718 (N_11718,N_6397,N_8197);
xor U11719 (N_11719,N_7538,N_6256);
nor U11720 (N_11720,N_7583,N_6344);
nor U11721 (N_11721,N_6271,N_9163);
and U11722 (N_11722,N_8713,N_9136);
or U11723 (N_11723,N_6987,N_6728);
nand U11724 (N_11724,N_6355,N_9330);
and U11725 (N_11725,N_7947,N_7193);
nand U11726 (N_11726,N_7172,N_9041);
or U11727 (N_11727,N_8262,N_7406);
and U11728 (N_11728,N_6834,N_8070);
xnor U11729 (N_11729,N_8834,N_6975);
xor U11730 (N_11730,N_8352,N_7923);
nor U11731 (N_11731,N_8938,N_6903);
nor U11732 (N_11732,N_8006,N_8100);
xnor U11733 (N_11733,N_9122,N_6657);
xnor U11734 (N_11734,N_8525,N_6631);
nor U11735 (N_11735,N_8436,N_8926);
nor U11736 (N_11736,N_6750,N_8279);
and U11737 (N_11737,N_6497,N_7547);
xor U11738 (N_11738,N_9301,N_9109);
or U11739 (N_11739,N_9036,N_7736);
xnor U11740 (N_11740,N_6670,N_8078);
and U11741 (N_11741,N_8121,N_8381);
or U11742 (N_11742,N_6431,N_6961);
xor U11743 (N_11743,N_7190,N_7199);
nor U11744 (N_11744,N_8840,N_6304);
nor U11745 (N_11745,N_7247,N_7306);
nor U11746 (N_11746,N_6969,N_7530);
or U11747 (N_11747,N_9343,N_8740);
and U11748 (N_11748,N_7426,N_6965);
and U11749 (N_11749,N_8842,N_8447);
nand U11750 (N_11750,N_7811,N_8336);
nor U11751 (N_11751,N_7634,N_8167);
and U11752 (N_11752,N_8507,N_8005);
nor U11753 (N_11753,N_7489,N_8756);
and U11754 (N_11754,N_8457,N_7396);
nand U11755 (N_11755,N_7718,N_8885);
nand U11756 (N_11756,N_8182,N_6905);
nand U11757 (N_11757,N_8632,N_7743);
or U11758 (N_11758,N_7050,N_7677);
or U11759 (N_11759,N_6707,N_8816);
xnor U11760 (N_11760,N_7111,N_7325);
nand U11761 (N_11761,N_7536,N_9170);
nor U11762 (N_11762,N_9027,N_6919);
xnor U11763 (N_11763,N_7987,N_6866);
nand U11764 (N_11764,N_8237,N_8944);
and U11765 (N_11765,N_8322,N_9129);
and U11766 (N_11766,N_6618,N_8629);
or U11767 (N_11767,N_8297,N_6996);
xor U11768 (N_11768,N_7425,N_9156);
xor U11769 (N_11769,N_8989,N_7434);
xor U11770 (N_11770,N_8179,N_9195);
and U11771 (N_11771,N_6927,N_6322);
nor U11772 (N_11772,N_9131,N_7316);
nand U11773 (N_11773,N_6610,N_9267);
or U11774 (N_11774,N_8808,N_7025);
or U11775 (N_11775,N_7214,N_8666);
and U11776 (N_11776,N_8529,N_8178);
xor U11777 (N_11777,N_9185,N_6488);
xnor U11778 (N_11778,N_7184,N_6525);
and U11779 (N_11779,N_9008,N_6529);
or U11780 (N_11780,N_8038,N_7501);
and U11781 (N_11781,N_7911,N_8988);
nand U11782 (N_11782,N_7612,N_8521);
nand U11783 (N_11783,N_8022,N_6274);
xnor U11784 (N_11784,N_6811,N_6964);
nand U11785 (N_11785,N_8334,N_8866);
and U11786 (N_11786,N_7509,N_6504);
xor U11787 (N_11787,N_8978,N_8958);
or U11788 (N_11788,N_6759,N_7851);
xnor U11789 (N_11789,N_7797,N_7408);
or U11790 (N_11790,N_6439,N_7082);
xor U11791 (N_11791,N_7531,N_6772);
xor U11792 (N_11792,N_6781,N_7924);
nand U11793 (N_11793,N_9193,N_8771);
and U11794 (N_11794,N_7766,N_8298);
nor U11795 (N_11795,N_8366,N_7124);
or U11796 (N_11796,N_8527,N_9318);
or U11797 (N_11797,N_6904,N_9183);
xnor U11798 (N_11798,N_7617,N_7168);
nand U11799 (N_11799,N_6356,N_7743);
nand U11800 (N_11800,N_7709,N_7301);
nor U11801 (N_11801,N_7273,N_6995);
or U11802 (N_11802,N_9065,N_7372);
xnor U11803 (N_11803,N_6482,N_8187);
and U11804 (N_11804,N_7572,N_9275);
nor U11805 (N_11805,N_6992,N_7782);
and U11806 (N_11806,N_9216,N_6730);
nand U11807 (N_11807,N_8193,N_7779);
nand U11808 (N_11808,N_7269,N_7407);
nand U11809 (N_11809,N_6993,N_7437);
and U11810 (N_11810,N_6713,N_6406);
nor U11811 (N_11811,N_8715,N_6858);
and U11812 (N_11812,N_7740,N_8970);
or U11813 (N_11813,N_8984,N_8467);
and U11814 (N_11814,N_9267,N_7164);
nor U11815 (N_11815,N_8645,N_6687);
xnor U11816 (N_11816,N_8052,N_7226);
nor U11817 (N_11817,N_8929,N_7126);
nor U11818 (N_11818,N_6690,N_8352);
and U11819 (N_11819,N_8772,N_9116);
nand U11820 (N_11820,N_7565,N_8913);
xor U11821 (N_11821,N_8466,N_8983);
nor U11822 (N_11822,N_7990,N_6913);
and U11823 (N_11823,N_7991,N_9106);
xnor U11824 (N_11824,N_6876,N_6748);
nor U11825 (N_11825,N_9078,N_7890);
and U11826 (N_11826,N_7974,N_6367);
nor U11827 (N_11827,N_6332,N_9112);
nand U11828 (N_11828,N_8750,N_7454);
and U11829 (N_11829,N_6840,N_9151);
nor U11830 (N_11830,N_8667,N_8755);
xnor U11831 (N_11831,N_8269,N_8858);
nand U11832 (N_11832,N_7791,N_9308);
and U11833 (N_11833,N_7030,N_7392);
nor U11834 (N_11834,N_8201,N_6796);
xnor U11835 (N_11835,N_8560,N_7526);
and U11836 (N_11836,N_6839,N_8437);
xor U11837 (N_11837,N_7340,N_6691);
and U11838 (N_11838,N_7404,N_7543);
xnor U11839 (N_11839,N_6761,N_9219);
and U11840 (N_11840,N_9245,N_8713);
or U11841 (N_11841,N_6502,N_7492);
and U11842 (N_11842,N_6328,N_6686);
or U11843 (N_11843,N_7190,N_8013);
nor U11844 (N_11844,N_7126,N_7272);
and U11845 (N_11845,N_9032,N_8236);
and U11846 (N_11846,N_8973,N_9256);
and U11847 (N_11847,N_9358,N_8564);
nand U11848 (N_11848,N_8573,N_9067);
nand U11849 (N_11849,N_6516,N_9370);
xnor U11850 (N_11850,N_9126,N_9292);
or U11851 (N_11851,N_7342,N_6426);
nor U11852 (N_11852,N_8883,N_6440);
nor U11853 (N_11853,N_7861,N_8788);
xnor U11854 (N_11854,N_7736,N_7882);
and U11855 (N_11855,N_6506,N_8348);
or U11856 (N_11856,N_6957,N_7471);
xor U11857 (N_11857,N_6600,N_8780);
and U11858 (N_11858,N_7581,N_8180);
nor U11859 (N_11859,N_7491,N_8589);
and U11860 (N_11860,N_6746,N_9206);
nand U11861 (N_11861,N_7386,N_8047);
and U11862 (N_11862,N_7879,N_8709);
nor U11863 (N_11863,N_7707,N_7515);
and U11864 (N_11864,N_9287,N_8012);
nand U11865 (N_11865,N_9117,N_6586);
or U11866 (N_11866,N_6408,N_8594);
and U11867 (N_11867,N_8658,N_6572);
xnor U11868 (N_11868,N_8919,N_9090);
and U11869 (N_11869,N_8011,N_8199);
xnor U11870 (N_11870,N_6253,N_8890);
xnor U11871 (N_11871,N_7880,N_8215);
xor U11872 (N_11872,N_8736,N_7143);
or U11873 (N_11873,N_8792,N_7139);
and U11874 (N_11874,N_7291,N_8476);
xor U11875 (N_11875,N_8449,N_8393);
xnor U11876 (N_11876,N_7284,N_6328);
nor U11877 (N_11877,N_6789,N_9182);
nand U11878 (N_11878,N_8797,N_8165);
xnor U11879 (N_11879,N_6950,N_8765);
xnor U11880 (N_11880,N_9101,N_6333);
nand U11881 (N_11881,N_7519,N_8955);
or U11882 (N_11882,N_8780,N_6306);
and U11883 (N_11883,N_6568,N_6698);
and U11884 (N_11884,N_8639,N_8887);
nand U11885 (N_11885,N_8155,N_6994);
xnor U11886 (N_11886,N_7758,N_9240);
nor U11887 (N_11887,N_6624,N_8451);
nand U11888 (N_11888,N_7612,N_9281);
nor U11889 (N_11889,N_8220,N_7626);
nand U11890 (N_11890,N_6311,N_8447);
and U11891 (N_11891,N_8688,N_7149);
nand U11892 (N_11892,N_6833,N_7581);
nand U11893 (N_11893,N_6652,N_7843);
xor U11894 (N_11894,N_7556,N_9364);
and U11895 (N_11895,N_8850,N_8412);
and U11896 (N_11896,N_7918,N_8364);
and U11897 (N_11897,N_8622,N_6568);
nor U11898 (N_11898,N_8384,N_8457);
nand U11899 (N_11899,N_9171,N_9317);
and U11900 (N_11900,N_9082,N_7744);
or U11901 (N_11901,N_8988,N_7831);
nor U11902 (N_11902,N_6398,N_6300);
nand U11903 (N_11903,N_8334,N_9274);
xor U11904 (N_11904,N_7016,N_6925);
nor U11905 (N_11905,N_9048,N_6388);
or U11906 (N_11906,N_6381,N_6669);
and U11907 (N_11907,N_7673,N_8072);
nor U11908 (N_11908,N_6613,N_8481);
and U11909 (N_11909,N_7785,N_7183);
xnor U11910 (N_11910,N_7957,N_9068);
xnor U11911 (N_11911,N_7834,N_7753);
nor U11912 (N_11912,N_8039,N_9146);
nand U11913 (N_11913,N_9374,N_8143);
nand U11914 (N_11914,N_6793,N_9111);
xor U11915 (N_11915,N_8159,N_6408);
nor U11916 (N_11916,N_9255,N_6817);
xor U11917 (N_11917,N_9065,N_6708);
and U11918 (N_11918,N_7039,N_6303);
nand U11919 (N_11919,N_8448,N_7203);
xnor U11920 (N_11920,N_7727,N_6401);
nand U11921 (N_11921,N_7540,N_6542);
nand U11922 (N_11922,N_7953,N_9059);
and U11923 (N_11923,N_7155,N_9225);
xor U11924 (N_11924,N_6558,N_7351);
xor U11925 (N_11925,N_6731,N_6839);
and U11926 (N_11926,N_8983,N_7676);
nor U11927 (N_11927,N_8129,N_7757);
or U11928 (N_11928,N_7372,N_8614);
nor U11929 (N_11929,N_8809,N_9331);
and U11930 (N_11930,N_9243,N_7508);
nand U11931 (N_11931,N_9308,N_6372);
and U11932 (N_11932,N_8408,N_8495);
and U11933 (N_11933,N_7693,N_8381);
nand U11934 (N_11934,N_7732,N_8821);
nor U11935 (N_11935,N_6809,N_7264);
or U11936 (N_11936,N_6631,N_8349);
nor U11937 (N_11937,N_8741,N_7475);
xnor U11938 (N_11938,N_8002,N_7126);
nand U11939 (N_11939,N_7774,N_8325);
and U11940 (N_11940,N_9222,N_6511);
nand U11941 (N_11941,N_6958,N_6972);
nor U11942 (N_11942,N_7793,N_6252);
or U11943 (N_11943,N_6566,N_7760);
xor U11944 (N_11944,N_7565,N_7038);
and U11945 (N_11945,N_9347,N_7492);
or U11946 (N_11946,N_9195,N_8311);
nand U11947 (N_11947,N_9087,N_6727);
and U11948 (N_11948,N_9263,N_9084);
or U11949 (N_11949,N_9239,N_6546);
and U11950 (N_11950,N_8248,N_8916);
xor U11951 (N_11951,N_8922,N_8626);
nor U11952 (N_11952,N_7332,N_9015);
nor U11953 (N_11953,N_9052,N_6936);
nor U11954 (N_11954,N_6385,N_7638);
and U11955 (N_11955,N_7902,N_7557);
nor U11956 (N_11956,N_7677,N_8214);
xnor U11957 (N_11957,N_8221,N_7505);
and U11958 (N_11958,N_8184,N_7300);
nand U11959 (N_11959,N_8111,N_7147);
nand U11960 (N_11960,N_9359,N_8427);
or U11961 (N_11961,N_7285,N_6654);
xor U11962 (N_11962,N_8846,N_9050);
nor U11963 (N_11963,N_7454,N_7684);
and U11964 (N_11964,N_9033,N_7816);
or U11965 (N_11965,N_6952,N_9088);
or U11966 (N_11966,N_7162,N_7838);
nand U11967 (N_11967,N_6356,N_8976);
or U11968 (N_11968,N_6974,N_8867);
nor U11969 (N_11969,N_8815,N_6775);
and U11970 (N_11970,N_6358,N_7952);
or U11971 (N_11971,N_7475,N_8360);
nor U11972 (N_11972,N_7773,N_7862);
nand U11973 (N_11973,N_7617,N_8836);
and U11974 (N_11974,N_8397,N_8388);
nand U11975 (N_11975,N_7393,N_6627);
xor U11976 (N_11976,N_8987,N_9253);
nor U11977 (N_11977,N_6270,N_8630);
or U11978 (N_11978,N_6967,N_9292);
or U11979 (N_11979,N_8749,N_6435);
or U11980 (N_11980,N_8868,N_6583);
nand U11981 (N_11981,N_9263,N_7957);
nand U11982 (N_11982,N_6387,N_6713);
nand U11983 (N_11983,N_6516,N_8044);
or U11984 (N_11984,N_8740,N_7159);
nand U11985 (N_11985,N_8229,N_6525);
nor U11986 (N_11986,N_6666,N_7447);
xor U11987 (N_11987,N_8116,N_7345);
or U11988 (N_11988,N_6271,N_9331);
and U11989 (N_11989,N_7351,N_7033);
nor U11990 (N_11990,N_6722,N_8605);
nand U11991 (N_11991,N_7398,N_8626);
or U11992 (N_11992,N_7542,N_8909);
and U11993 (N_11993,N_8446,N_9330);
nand U11994 (N_11994,N_8000,N_9010);
xnor U11995 (N_11995,N_6749,N_7051);
and U11996 (N_11996,N_7464,N_9286);
and U11997 (N_11997,N_6508,N_6372);
nor U11998 (N_11998,N_8004,N_6824);
or U11999 (N_11999,N_8723,N_7006);
nand U12000 (N_12000,N_8795,N_8976);
and U12001 (N_12001,N_8315,N_8006);
nand U12002 (N_12002,N_6559,N_7738);
or U12003 (N_12003,N_8820,N_9319);
nand U12004 (N_12004,N_7647,N_8084);
nand U12005 (N_12005,N_9122,N_8903);
nand U12006 (N_12006,N_6951,N_8844);
nor U12007 (N_12007,N_7358,N_8921);
nor U12008 (N_12008,N_9368,N_8006);
or U12009 (N_12009,N_8564,N_6880);
or U12010 (N_12010,N_6884,N_6813);
xnor U12011 (N_12011,N_6603,N_6365);
nor U12012 (N_12012,N_7172,N_8929);
or U12013 (N_12013,N_7819,N_8385);
xor U12014 (N_12014,N_6794,N_8039);
nor U12015 (N_12015,N_7279,N_6389);
or U12016 (N_12016,N_8487,N_8783);
and U12017 (N_12017,N_6969,N_9075);
xnor U12018 (N_12018,N_6707,N_6364);
nand U12019 (N_12019,N_6954,N_8179);
xnor U12020 (N_12020,N_7839,N_8802);
and U12021 (N_12021,N_8483,N_6475);
xor U12022 (N_12022,N_8995,N_7770);
xor U12023 (N_12023,N_8522,N_7043);
or U12024 (N_12024,N_8499,N_6803);
nor U12025 (N_12025,N_7775,N_6518);
and U12026 (N_12026,N_7016,N_7029);
nor U12027 (N_12027,N_7840,N_7424);
or U12028 (N_12028,N_7960,N_8656);
and U12029 (N_12029,N_8031,N_6420);
and U12030 (N_12030,N_7893,N_9334);
nand U12031 (N_12031,N_7712,N_6943);
nand U12032 (N_12032,N_8108,N_8200);
nand U12033 (N_12033,N_8740,N_6820);
nand U12034 (N_12034,N_7206,N_7326);
nor U12035 (N_12035,N_8315,N_6667);
and U12036 (N_12036,N_7925,N_8427);
nor U12037 (N_12037,N_6751,N_9203);
nand U12038 (N_12038,N_9071,N_8017);
and U12039 (N_12039,N_8356,N_8094);
and U12040 (N_12040,N_8832,N_7615);
nand U12041 (N_12041,N_7425,N_8936);
or U12042 (N_12042,N_7909,N_6451);
nand U12043 (N_12043,N_6941,N_8789);
or U12044 (N_12044,N_7584,N_9341);
or U12045 (N_12045,N_6321,N_8330);
nor U12046 (N_12046,N_8189,N_6534);
xnor U12047 (N_12047,N_8572,N_6313);
and U12048 (N_12048,N_8244,N_6583);
nand U12049 (N_12049,N_6826,N_7792);
nor U12050 (N_12050,N_7697,N_8151);
nand U12051 (N_12051,N_6921,N_6810);
and U12052 (N_12052,N_8209,N_6366);
nor U12053 (N_12053,N_7506,N_9317);
and U12054 (N_12054,N_6616,N_8738);
nand U12055 (N_12055,N_6502,N_8826);
nand U12056 (N_12056,N_8378,N_6552);
or U12057 (N_12057,N_8443,N_7443);
nand U12058 (N_12058,N_8365,N_8505);
xor U12059 (N_12059,N_6444,N_7512);
and U12060 (N_12060,N_7988,N_8187);
nand U12061 (N_12061,N_6974,N_7408);
nand U12062 (N_12062,N_6432,N_7646);
or U12063 (N_12063,N_7017,N_7507);
xor U12064 (N_12064,N_8495,N_9335);
nor U12065 (N_12065,N_8634,N_7468);
nor U12066 (N_12066,N_6528,N_9274);
or U12067 (N_12067,N_7180,N_8255);
nand U12068 (N_12068,N_8922,N_6898);
xnor U12069 (N_12069,N_9185,N_7879);
xor U12070 (N_12070,N_8160,N_8227);
nor U12071 (N_12071,N_9061,N_7193);
xnor U12072 (N_12072,N_7431,N_8683);
and U12073 (N_12073,N_7730,N_7433);
xnor U12074 (N_12074,N_6255,N_8911);
and U12075 (N_12075,N_8595,N_7221);
nor U12076 (N_12076,N_8245,N_6546);
and U12077 (N_12077,N_8137,N_7545);
or U12078 (N_12078,N_6542,N_6580);
and U12079 (N_12079,N_8259,N_8425);
or U12080 (N_12080,N_8446,N_7158);
nand U12081 (N_12081,N_6475,N_7960);
nor U12082 (N_12082,N_7952,N_7761);
and U12083 (N_12083,N_8655,N_8420);
nand U12084 (N_12084,N_6874,N_8261);
nor U12085 (N_12085,N_9198,N_7513);
xnor U12086 (N_12086,N_8306,N_6829);
or U12087 (N_12087,N_8137,N_8810);
nand U12088 (N_12088,N_8876,N_7788);
xor U12089 (N_12089,N_8668,N_8797);
and U12090 (N_12090,N_6948,N_7568);
and U12091 (N_12091,N_8789,N_7902);
nor U12092 (N_12092,N_7088,N_8617);
nor U12093 (N_12093,N_6732,N_7968);
nand U12094 (N_12094,N_7143,N_7919);
and U12095 (N_12095,N_6546,N_7643);
or U12096 (N_12096,N_9048,N_7992);
nor U12097 (N_12097,N_8276,N_7049);
or U12098 (N_12098,N_6332,N_6652);
nand U12099 (N_12099,N_7818,N_8702);
nor U12100 (N_12100,N_6341,N_7242);
nand U12101 (N_12101,N_9297,N_7457);
xnor U12102 (N_12102,N_7225,N_6508);
or U12103 (N_12103,N_9176,N_8876);
and U12104 (N_12104,N_6553,N_8729);
or U12105 (N_12105,N_9033,N_6903);
nor U12106 (N_12106,N_8425,N_6961);
nand U12107 (N_12107,N_7966,N_8070);
and U12108 (N_12108,N_9230,N_6340);
nor U12109 (N_12109,N_7624,N_7022);
xor U12110 (N_12110,N_7857,N_8553);
nand U12111 (N_12111,N_8807,N_8634);
and U12112 (N_12112,N_6981,N_7884);
nand U12113 (N_12113,N_7493,N_6519);
or U12114 (N_12114,N_6894,N_8275);
xor U12115 (N_12115,N_8794,N_8056);
or U12116 (N_12116,N_6377,N_7046);
nor U12117 (N_12117,N_6474,N_6512);
nand U12118 (N_12118,N_8805,N_8551);
xnor U12119 (N_12119,N_7714,N_7543);
xnor U12120 (N_12120,N_6721,N_9371);
and U12121 (N_12121,N_8427,N_7326);
and U12122 (N_12122,N_9194,N_7688);
nand U12123 (N_12123,N_6796,N_7631);
nor U12124 (N_12124,N_6493,N_8925);
xnor U12125 (N_12125,N_8700,N_9267);
and U12126 (N_12126,N_8592,N_7114);
xnor U12127 (N_12127,N_8826,N_7896);
nand U12128 (N_12128,N_7533,N_6775);
or U12129 (N_12129,N_6438,N_9262);
nand U12130 (N_12130,N_7008,N_8095);
nand U12131 (N_12131,N_8179,N_8462);
xnor U12132 (N_12132,N_6323,N_9041);
or U12133 (N_12133,N_7254,N_8014);
nor U12134 (N_12134,N_7233,N_6803);
and U12135 (N_12135,N_7809,N_8018);
and U12136 (N_12136,N_8538,N_8823);
nand U12137 (N_12137,N_6421,N_7128);
xnor U12138 (N_12138,N_7876,N_7359);
nor U12139 (N_12139,N_6264,N_6446);
nand U12140 (N_12140,N_8124,N_8774);
and U12141 (N_12141,N_6550,N_6974);
or U12142 (N_12142,N_9271,N_6487);
xnor U12143 (N_12143,N_7653,N_6571);
and U12144 (N_12144,N_7401,N_7880);
and U12145 (N_12145,N_8821,N_7131);
xor U12146 (N_12146,N_9279,N_8621);
and U12147 (N_12147,N_6582,N_9207);
or U12148 (N_12148,N_9262,N_9168);
and U12149 (N_12149,N_6975,N_6605);
nor U12150 (N_12150,N_6728,N_7018);
nand U12151 (N_12151,N_7960,N_6530);
nor U12152 (N_12152,N_8032,N_7425);
and U12153 (N_12153,N_8439,N_6434);
or U12154 (N_12154,N_8611,N_8786);
nand U12155 (N_12155,N_6376,N_8581);
nor U12156 (N_12156,N_6929,N_8538);
nor U12157 (N_12157,N_6509,N_6933);
nand U12158 (N_12158,N_6682,N_8416);
or U12159 (N_12159,N_7178,N_9044);
and U12160 (N_12160,N_7441,N_7523);
nand U12161 (N_12161,N_6457,N_9346);
nand U12162 (N_12162,N_7731,N_7579);
xor U12163 (N_12163,N_8971,N_7990);
and U12164 (N_12164,N_8575,N_6271);
xnor U12165 (N_12165,N_8795,N_6738);
xnor U12166 (N_12166,N_8482,N_7634);
and U12167 (N_12167,N_7020,N_7261);
and U12168 (N_12168,N_7418,N_9139);
and U12169 (N_12169,N_7414,N_9266);
or U12170 (N_12170,N_9287,N_8748);
or U12171 (N_12171,N_8045,N_6469);
and U12172 (N_12172,N_7046,N_7269);
nand U12173 (N_12173,N_8150,N_7668);
or U12174 (N_12174,N_9165,N_7280);
nor U12175 (N_12175,N_6936,N_6342);
xor U12176 (N_12176,N_9025,N_7944);
xor U12177 (N_12177,N_6733,N_9179);
and U12178 (N_12178,N_7084,N_8798);
and U12179 (N_12179,N_6563,N_6348);
nor U12180 (N_12180,N_7528,N_8929);
xor U12181 (N_12181,N_7120,N_8551);
or U12182 (N_12182,N_8462,N_7413);
nor U12183 (N_12183,N_6627,N_9001);
nor U12184 (N_12184,N_7778,N_8666);
nand U12185 (N_12185,N_9172,N_8200);
nor U12186 (N_12186,N_7894,N_6596);
nor U12187 (N_12187,N_6434,N_7142);
nor U12188 (N_12188,N_6617,N_6760);
and U12189 (N_12189,N_6732,N_9124);
nor U12190 (N_12190,N_7055,N_6253);
nor U12191 (N_12191,N_8987,N_7003);
and U12192 (N_12192,N_8845,N_6791);
and U12193 (N_12193,N_6263,N_7534);
nor U12194 (N_12194,N_8176,N_7335);
or U12195 (N_12195,N_7638,N_9093);
xor U12196 (N_12196,N_9029,N_7904);
or U12197 (N_12197,N_8499,N_9166);
and U12198 (N_12198,N_7168,N_6654);
nor U12199 (N_12199,N_7304,N_6641);
xor U12200 (N_12200,N_7310,N_6926);
nand U12201 (N_12201,N_6451,N_6658);
nand U12202 (N_12202,N_7843,N_6727);
nor U12203 (N_12203,N_7471,N_7098);
xor U12204 (N_12204,N_6844,N_6872);
xnor U12205 (N_12205,N_6396,N_7791);
or U12206 (N_12206,N_8120,N_8089);
nand U12207 (N_12207,N_8174,N_6831);
or U12208 (N_12208,N_7294,N_8457);
and U12209 (N_12209,N_8087,N_6856);
or U12210 (N_12210,N_8896,N_9281);
nand U12211 (N_12211,N_6624,N_8513);
xnor U12212 (N_12212,N_9171,N_6889);
or U12213 (N_12213,N_8022,N_7263);
nor U12214 (N_12214,N_9198,N_9254);
xnor U12215 (N_12215,N_8966,N_7368);
nand U12216 (N_12216,N_9137,N_8171);
xnor U12217 (N_12217,N_8977,N_8954);
nor U12218 (N_12218,N_8050,N_9144);
nor U12219 (N_12219,N_8480,N_7040);
and U12220 (N_12220,N_7172,N_7391);
xnor U12221 (N_12221,N_6561,N_7526);
xor U12222 (N_12222,N_7159,N_7654);
nand U12223 (N_12223,N_8356,N_6333);
and U12224 (N_12224,N_6777,N_6673);
and U12225 (N_12225,N_8891,N_8641);
nor U12226 (N_12226,N_9372,N_8722);
nand U12227 (N_12227,N_8828,N_9080);
or U12228 (N_12228,N_8252,N_8749);
or U12229 (N_12229,N_7675,N_7314);
nor U12230 (N_12230,N_6771,N_6979);
nand U12231 (N_12231,N_9212,N_8406);
and U12232 (N_12232,N_8799,N_6423);
xor U12233 (N_12233,N_9265,N_7499);
xor U12234 (N_12234,N_6252,N_7452);
nor U12235 (N_12235,N_7131,N_7936);
and U12236 (N_12236,N_7945,N_7384);
xor U12237 (N_12237,N_6839,N_8666);
nand U12238 (N_12238,N_8561,N_8819);
xnor U12239 (N_12239,N_8804,N_6738);
xor U12240 (N_12240,N_7986,N_8651);
nand U12241 (N_12241,N_6997,N_7773);
and U12242 (N_12242,N_8412,N_7946);
xor U12243 (N_12243,N_8775,N_7872);
nor U12244 (N_12244,N_8959,N_7333);
or U12245 (N_12245,N_6613,N_8545);
or U12246 (N_12246,N_9356,N_6367);
xor U12247 (N_12247,N_7582,N_6859);
nor U12248 (N_12248,N_6284,N_7975);
nor U12249 (N_12249,N_8306,N_8238);
and U12250 (N_12250,N_6893,N_7025);
or U12251 (N_12251,N_6906,N_6803);
or U12252 (N_12252,N_8650,N_8759);
or U12253 (N_12253,N_7969,N_7746);
nand U12254 (N_12254,N_8317,N_6538);
and U12255 (N_12255,N_7714,N_7444);
nor U12256 (N_12256,N_7668,N_6573);
nor U12257 (N_12257,N_6621,N_6534);
xnor U12258 (N_12258,N_6607,N_9360);
nand U12259 (N_12259,N_7845,N_7974);
nor U12260 (N_12260,N_8742,N_7134);
xnor U12261 (N_12261,N_8491,N_8356);
or U12262 (N_12262,N_9347,N_8800);
nand U12263 (N_12263,N_7548,N_6873);
xnor U12264 (N_12264,N_8975,N_6421);
xor U12265 (N_12265,N_8702,N_6608);
and U12266 (N_12266,N_8071,N_7576);
and U12267 (N_12267,N_7840,N_7954);
and U12268 (N_12268,N_8522,N_6314);
and U12269 (N_12269,N_7479,N_6987);
and U12270 (N_12270,N_7964,N_8346);
xor U12271 (N_12271,N_6854,N_6296);
nand U12272 (N_12272,N_9348,N_8139);
nor U12273 (N_12273,N_7275,N_7954);
nand U12274 (N_12274,N_6753,N_8220);
nand U12275 (N_12275,N_6463,N_9163);
nor U12276 (N_12276,N_6856,N_6978);
or U12277 (N_12277,N_7656,N_8702);
nor U12278 (N_12278,N_7939,N_7133);
xor U12279 (N_12279,N_9105,N_7797);
nand U12280 (N_12280,N_7158,N_8590);
xnor U12281 (N_12281,N_8893,N_8815);
nor U12282 (N_12282,N_8747,N_8341);
and U12283 (N_12283,N_6680,N_7131);
and U12284 (N_12284,N_9190,N_7973);
or U12285 (N_12285,N_7747,N_7679);
or U12286 (N_12286,N_6931,N_9257);
xnor U12287 (N_12287,N_8213,N_9262);
or U12288 (N_12288,N_7199,N_6628);
or U12289 (N_12289,N_6634,N_6587);
and U12290 (N_12290,N_6340,N_6267);
nor U12291 (N_12291,N_8925,N_7993);
nor U12292 (N_12292,N_6361,N_7947);
and U12293 (N_12293,N_7596,N_8207);
xnor U12294 (N_12294,N_6516,N_8531);
nor U12295 (N_12295,N_8276,N_8678);
nand U12296 (N_12296,N_6854,N_7767);
or U12297 (N_12297,N_9114,N_7182);
and U12298 (N_12298,N_9293,N_9346);
or U12299 (N_12299,N_8666,N_9298);
nand U12300 (N_12300,N_6909,N_9047);
nor U12301 (N_12301,N_7268,N_8613);
nand U12302 (N_12302,N_8697,N_7521);
xnor U12303 (N_12303,N_7967,N_8143);
nand U12304 (N_12304,N_8992,N_7900);
nand U12305 (N_12305,N_7388,N_8966);
and U12306 (N_12306,N_8672,N_6251);
nor U12307 (N_12307,N_8852,N_7805);
xor U12308 (N_12308,N_8573,N_6743);
xor U12309 (N_12309,N_9071,N_7464);
xnor U12310 (N_12310,N_6926,N_7049);
nand U12311 (N_12311,N_8285,N_8865);
nor U12312 (N_12312,N_7763,N_8892);
or U12313 (N_12313,N_7350,N_8597);
and U12314 (N_12314,N_8199,N_9300);
xor U12315 (N_12315,N_7406,N_9026);
nand U12316 (N_12316,N_6884,N_8313);
nand U12317 (N_12317,N_7930,N_7085);
nor U12318 (N_12318,N_8785,N_6649);
or U12319 (N_12319,N_8698,N_7664);
nor U12320 (N_12320,N_6870,N_7425);
or U12321 (N_12321,N_9009,N_9206);
or U12322 (N_12322,N_6623,N_6774);
or U12323 (N_12323,N_9215,N_6358);
nor U12324 (N_12324,N_7763,N_7146);
or U12325 (N_12325,N_8802,N_9268);
xor U12326 (N_12326,N_6335,N_7764);
and U12327 (N_12327,N_7742,N_9359);
xnor U12328 (N_12328,N_9335,N_6663);
or U12329 (N_12329,N_8063,N_8816);
xor U12330 (N_12330,N_6745,N_7836);
xor U12331 (N_12331,N_7708,N_7507);
nor U12332 (N_12332,N_8498,N_8905);
and U12333 (N_12333,N_8717,N_6919);
and U12334 (N_12334,N_6941,N_6863);
nor U12335 (N_12335,N_9287,N_8625);
nand U12336 (N_12336,N_8327,N_6771);
nor U12337 (N_12337,N_6261,N_8514);
nand U12338 (N_12338,N_8966,N_7087);
or U12339 (N_12339,N_6716,N_6337);
or U12340 (N_12340,N_8322,N_6461);
nand U12341 (N_12341,N_6529,N_6348);
nand U12342 (N_12342,N_8537,N_9004);
and U12343 (N_12343,N_8829,N_8621);
nor U12344 (N_12344,N_8402,N_6732);
nand U12345 (N_12345,N_9040,N_6734);
nand U12346 (N_12346,N_6801,N_8574);
and U12347 (N_12347,N_8752,N_8934);
nand U12348 (N_12348,N_8632,N_8455);
xor U12349 (N_12349,N_6820,N_9189);
nand U12350 (N_12350,N_8357,N_9300);
and U12351 (N_12351,N_6896,N_8948);
nor U12352 (N_12352,N_8073,N_7965);
xor U12353 (N_12353,N_8961,N_7954);
or U12354 (N_12354,N_9174,N_6771);
and U12355 (N_12355,N_7968,N_7541);
or U12356 (N_12356,N_8118,N_7715);
or U12357 (N_12357,N_8602,N_7837);
and U12358 (N_12358,N_6317,N_8542);
and U12359 (N_12359,N_8572,N_6253);
nand U12360 (N_12360,N_6352,N_6823);
and U12361 (N_12361,N_8705,N_7562);
and U12362 (N_12362,N_6759,N_8231);
or U12363 (N_12363,N_7335,N_8459);
and U12364 (N_12364,N_8546,N_8058);
nand U12365 (N_12365,N_8488,N_8861);
nand U12366 (N_12366,N_7641,N_8515);
and U12367 (N_12367,N_7513,N_7211);
nand U12368 (N_12368,N_6848,N_9050);
nand U12369 (N_12369,N_8183,N_6600);
and U12370 (N_12370,N_8696,N_6714);
nor U12371 (N_12371,N_8355,N_8351);
xor U12372 (N_12372,N_7914,N_8546);
nand U12373 (N_12373,N_7430,N_8157);
and U12374 (N_12374,N_8650,N_9184);
and U12375 (N_12375,N_9318,N_8209);
and U12376 (N_12376,N_7153,N_9236);
nor U12377 (N_12377,N_8912,N_8632);
and U12378 (N_12378,N_6935,N_9169);
or U12379 (N_12379,N_9095,N_8844);
xnor U12380 (N_12380,N_6535,N_8803);
nand U12381 (N_12381,N_7366,N_9305);
nor U12382 (N_12382,N_9146,N_6541);
xor U12383 (N_12383,N_6311,N_8394);
nand U12384 (N_12384,N_9248,N_8243);
and U12385 (N_12385,N_8788,N_8535);
nand U12386 (N_12386,N_7948,N_8581);
or U12387 (N_12387,N_7049,N_8166);
nor U12388 (N_12388,N_9209,N_9109);
nand U12389 (N_12389,N_6279,N_7563);
nor U12390 (N_12390,N_6724,N_8717);
and U12391 (N_12391,N_6388,N_8242);
or U12392 (N_12392,N_9048,N_8994);
xnor U12393 (N_12393,N_9282,N_8401);
nor U12394 (N_12394,N_9157,N_7705);
xnor U12395 (N_12395,N_7689,N_6746);
xor U12396 (N_12396,N_6452,N_8081);
or U12397 (N_12397,N_7723,N_8269);
xnor U12398 (N_12398,N_7141,N_8734);
or U12399 (N_12399,N_9231,N_9272);
and U12400 (N_12400,N_8983,N_8663);
or U12401 (N_12401,N_7558,N_7277);
or U12402 (N_12402,N_7733,N_6797);
xnor U12403 (N_12403,N_8329,N_7100);
nand U12404 (N_12404,N_7455,N_7370);
or U12405 (N_12405,N_8231,N_8596);
nor U12406 (N_12406,N_7540,N_7871);
nor U12407 (N_12407,N_8174,N_8529);
and U12408 (N_12408,N_8765,N_8191);
nand U12409 (N_12409,N_7057,N_9151);
and U12410 (N_12410,N_8127,N_6780);
nand U12411 (N_12411,N_8240,N_8539);
xor U12412 (N_12412,N_7972,N_8589);
and U12413 (N_12413,N_8146,N_8215);
and U12414 (N_12414,N_6300,N_9349);
xor U12415 (N_12415,N_7580,N_8838);
xnor U12416 (N_12416,N_6701,N_7534);
and U12417 (N_12417,N_7573,N_8401);
or U12418 (N_12418,N_8176,N_8928);
and U12419 (N_12419,N_6320,N_7403);
nor U12420 (N_12420,N_8604,N_7876);
and U12421 (N_12421,N_7162,N_7079);
and U12422 (N_12422,N_6432,N_7489);
and U12423 (N_12423,N_9097,N_8529);
and U12424 (N_12424,N_7553,N_8477);
nand U12425 (N_12425,N_6582,N_8822);
and U12426 (N_12426,N_9311,N_6372);
or U12427 (N_12427,N_7720,N_8738);
or U12428 (N_12428,N_7359,N_6959);
nor U12429 (N_12429,N_8382,N_6974);
xnor U12430 (N_12430,N_7248,N_7637);
xnor U12431 (N_12431,N_8384,N_9286);
and U12432 (N_12432,N_8044,N_8796);
and U12433 (N_12433,N_8319,N_6274);
xor U12434 (N_12434,N_8354,N_7626);
xnor U12435 (N_12435,N_7852,N_6742);
nor U12436 (N_12436,N_8742,N_8769);
and U12437 (N_12437,N_7415,N_6806);
nor U12438 (N_12438,N_7708,N_8268);
or U12439 (N_12439,N_6514,N_9097);
xor U12440 (N_12440,N_6832,N_7149);
xor U12441 (N_12441,N_8795,N_6876);
or U12442 (N_12442,N_8386,N_6457);
xnor U12443 (N_12443,N_7101,N_6602);
nor U12444 (N_12444,N_8948,N_8501);
xor U12445 (N_12445,N_7879,N_9000);
nand U12446 (N_12446,N_8367,N_9187);
xnor U12447 (N_12447,N_7544,N_8765);
nor U12448 (N_12448,N_6519,N_8006);
xnor U12449 (N_12449,N_7454,N_9028);
nand U12450 (N_12450,N_8735,N_6470);
nand U12451 (N_12451,N_6475,N_6596);
xnor U12452 (N_12452,N_9063,N_7915);
nand U12453 (N_12453,N_6994,N_9170);
nand U12454 (N_12454,N_6842,N_7694);
nand U12455 (N_12455,N_8156,N_6885);
nor U12456 (N_12456,N_8125,N_7022);
xor U12457 (N_12457,N_8498,N_6920);
and U12458 (N_12458,N_6491,N_8348);
or U12459 (N_12459,N_8888,N_9154);
nand U12460 (N_12460,N_8272,N_6660);
xor U12461 (N_12461,N_8205,N_8725);
nor U12462 (N_12462,N_8532,N_6343);
and U12463 (N_12463,N_8962,N_8514);
or U12464 (N_12464,N_7273,N_8800);
xor U12465 (N_12465,N_6891,N_7066);
and U12466 (N_12466,N_7600,N_8591);
nor U12467 (N_12467,N_7031,N_7051);
and U12468 (N_12468,N_7988,N_7829);
and U12469 (N_12469,N_8967,N_7790);
nand U12470 (N_12470,N_8486,N_7263);
nand U12471 (N_12471,N_9219,N_8197);
and U12472 (N_12472,N_6351,N_6440);
and U12473 (N_12473,N_6562,N_8418);
nand U12474 (N_12474,N_8463,N_8966);
xor U12475 (N_12475,N_8065,N_6475);
nor U12476 (N_12476,N_6743,N_8323);
or U12477 (N_12477,N_8935,N_6871);
xnor U12478 (N_12478,N_7274,N_7249);
nand U12479 (N_12479,N_7678,N_8408);
nor U12480 (N_12480,N_8735,N_7870);
nor U12481 (N_12481,N_8277,N_6347);
nand U12482 (N_12482,N_8106,N_6804);
or U12483 (N_12483,N_7046,N_7078);
nand U12484 (N_12484,N_7446,N_9136);
and U12485 (N_12485,N_6680,N_8102);
xnor U12486 (N_12486,N_7436,N_7139);
nor U12487 (N_12487,N_7974,N_8864);
nor U12488 (N_12488,N_9371,N_6589);
nand U12489 (N_12489,N_8118,N_8577);
xor U12490 (N_12490,N_9261,N_8903);
nand U12491 (N_12491,N_7286,N_8266);
nand U12492 (N_12492,N_9137,N_6311);
or U12493 (N_12493,N_7034,N_7621);
xor U12494 (N_12494,N_8413,N_6656);
xnor U12495 (N_12495,N_7082,N_7654);
and U12496 (N_12496,N_6998,N_6462);
nand U12497 (N_12497,N_6880,N_6741);
or U12498 (N_12498,N_7838,N_8660);
or U12499 (N_12499,N_9276,N_6565);
xnor U12500 (N_12500,N_10567,N_11478);
or U12501 (N_12501,N_11481,N_11801);
nand U12502 (N_12502,N_11748,N_9909);
or U12503 (N_12503,N_12338,N_11244);
and U12504 (N_12504,N_11012,N_10622);
nor U12505 (N_12505,N_12489,N_10082);
and U12506 (N_12506,N_11625,N_10204);
and U12507 (N_12507,N_9904,N_11807);
xnor U12508 (N_12508,N_10661,N_11149);
and U12509 (N_12509,N_9679,N_11958);
xnor U12510 (N_12510,N_11952,N_10614);
or U12511 (N_12511,N_11838,N_12498);
nand U12512 (N_12512,N_10077,N_12151);
xnor U12513 (N_12513,N_10882,N_12067);
nand U12514 (N_12514,N_11110,N_11351);
and U12515 (N_12515,N_12036,N_9652);
xor U12516 (N_12516,N_10926,N_11679);
nand U12517 (N_12517,N_11578,N_11642);
nor U12518 (N_12518,N_10382,N_9568);
or U12519 (N_12519,N_12419,N_11242);
xnor U12520 (N_12520,N_10149,N_11472);
and U12521 (N_12521,N_11218,N_10813);
nand U12522 (N_12522,N_11795,N_11320);
nand U12523 (N_12523,N_10133,N_10105);
and U12524 (N_12524,N_10880,N_10618);
nand U12525 (N_12525,N_9818,N_10623);
nand U12526 (N_12526,N_10144,N_10219);
xnor U12527 (N_12527,N_10521,N_11659);
or U12528 (N_12528,N_9874,N_10765);
or U12529 (N_12529,N_12331,N_9720);
nor U12530 (N_12530,N_12294,N_11518);
xnor U12531 (N_12531,N_12046,N_11014);
nand U12532 (N_12532,N_11825,N_11383);
nand U12533 (N_12533,N_11694,N_11687);
nand U12534 (N_12534,N_9965,N_9537);
or U12535 (N_12535,N_9545,N_9921);
or U12536 (N_12536,N_10986,N_9757);
nor U12537 (N_12537,N_11233,N_10202);
or U12538 (N_12538,N_12104,N_11224);
nor U12539 (N_12539,N_12119,N_11720);
or U12540 (N_12540,N_11048,N_9505);
nor U12541 (N_12541,N_11096,N_9748);
or U12542 (N_12542,N_9711,N_10901);
nor U12543 (N_12543,N_10557,N_11073);
nor U12544 (N_12544,N_11606,N_10635);
xnor U12545 (N_12545,N_11076,N_12187);
xnor U12546 (N_12546,N_10110,N_10467);
or U12547 (N_12547,N_9826,N_10950);
and U12548 (N_12548,N_10859,N_9459);
or U12549 (N_12549,N_10914,N_9585);
nand U12550 (N_12550,N_9954,N_10319);
nand U12551 (N_12551,N_9644,N_12199);
nor U12552 (N_12552,N_10751,N_12141);
or U12553 (N_12553,N_11199,N_12383);
or U12554 (N_12554,N_11272,N_11997);
xnor U12555 (N_12555,N_9663,N_12291);
nor U12556 (N_12556,N_11443,N_12314);
xor U12557 (N_12557,N_10108,N_11844);
xnor U12558 (N_12558,N_10266,N_10334);
nor U12559 (N_12559,N_10072,N_9469);
or U12560 (N_12560,N_11716,N_10491);
xnor U12561 (N_12561,N_11358,N_11792);
nand U12562 (N_12562,N_12364,N_11563);
nor U12563 (N_12563,N_11152,N_11975);
nand U12564 (N_12564,N_9816,N_11793);
and U12565 (N_12565,N_10695,N_10345);
and U12566 (N_12566,N_11496,N_9991);
nand U12567 (N_12567,N_12076,N_11289);
nor U12568 (N_12568,N_10747,N_10095);
nor U12569 (N_12569,N_10928,N_11401);
or U12570 (N_12570,N_9603,N_11196);
nor U12571 (N_12571,N_9792,N_11768);
nand U12572 (N_12572,N_12252,N_11163);
xnor U12573 (N_12573,N_12487,N_12296);
or U12574 (N_12574,N_9735,N_9739);
xor U12575 (N_12575,N_12081,N_12433);
or U12576 (N_12576,N_11534,N_10426);
nand U12577 (N_12577,N_11709,N_11011);
or U12578 (N_12578,N_11821,N_12039);
nor U12579 (N_12579,N_9598,N_9495);
or U12580 (N_12580,N_9432,N_10230);
nand U12581 (N_12581,N_10285,N_11460);
and U12582 (N_12582,N_10698,N_9674);
or U12583 (N_12583,N_9517,N_10865);
nor U12584 (N_12584,N_11368,N_9591);
xnor U12585 (N_12585,N_10729,N_10076);
and U12586 (N_12586,N_12392,N_9397);
nor U12587 (N_12587,N_10257,N_10134);
xor U12588 (N_12588,N_11780,N_11582);
or U12589 (N_12589,N_10418,N_12476);
xnor U12590 (N_12590,N_10783,N_10590);
nor U12591 (N_12591,N_12345,N_10093);
nand U12592 (N_12592,N_11644,N_11551);
nor U12593 (N_12593,N_10242,N_12420);
and U12594 (N_12594,N_11678,N_11256);
nand U12595 (N_12595,N_10657,N_12122);
nor U12596 (N_12596,N_10518,N_11751);
nand U12597 (N_12597,N_12227,N_10430);
or U12598 (N_12598,N_9615,N_12258);
or U12599 (N_12599,N_9628,N_11211);
or U12600 (N_12600,N_12134,N_10985);
nand U12601 (N_12601,N_10486,N_10044);
or U12602 (N_12602,N_11470,N_11866);
and U12603 (N_12603,N_9827,N_10469);
and U12604 (N_12604,N_9872,N_9718);
nand U12605 (N_12605,N_9883,N_12087);
nand U12606 (N_12606,N_9880,N_10852);
nand U12607 (N_12607,N_12232,N_11832);
xor U12608 (N_12608,N_10290,N_9836);
nand U12609 (N_12609,N_10015,N_9888);
nand U12610 (N_12610,N_9656,N_11041);
and U12611 (N_12611,N_9868,N_9911);
nor U12612 (N_12612,N_10723,N_11944);
and U12613 (N_12613,N_12013,N_10042);
xor U12614 (N_12614,N_10908,N_9492);
nor U12615 (N_12615,N_9688,N_11531);
and U12616 (N_12616,N_9813,N_9801);
nand U12617 (N_12617,N_12210,N_10707);
nor U12618 (N_12618,N_10611,N_9547);
xor U12619 (N_12619,N_9631,N_12177);
xnor U12620 (N_12620,N_9942,N_12064);
nor U12621 (N_12621,N_11493,N_9655);
nor U12622 (N_12622,N_10088,N_9572);
xor U12623 (N_12623,N_9482,N_12037);
and U12624 (N_12624,N_9392,N_11584);
or U12625 (N_12625,N_9993,N_10484);
nor U12626 (N_12626,N_10542,N_12479);
or U12627 (N_12627,N_12175,N_10966);
nand U12628 (N_12628,N_12200,N_11013);
nor U12629 (N_12629,N_11107,N_9574);
or U12630 (N_12630,N_9595,N_9564);
or U12631 (N_12631,N_10744,N_9925);
nor U12632 (N_12632,N_12299,N_11567);
xnor U12633 (N_12633,N_12322,N_11180);
or U12634 (N_12634,N_9383,N_11937);
or U12635 (N_12635,N_11423,N_11317);
xor U12636 (N_12636,N_10849,N_10700);
nand U12637 (N_12637,N_10036,N_11138);
nor U12638 (N_12638,N_11495,N_10066);
and U12639 (N_12639,N_9571,N_10330);
nand U12640 (N_12640,N_11992,N_9584);
nand U12641 (N_12641,N_9630,N_9839);
or U12642 (N_12642,N_11685,N_11396);
xor U12643 (N_12643,N_12408,N_10026);
xor U12644 (N_12644,N_9765,N_9789);
nand U12645 (N_12645,N_10048,N_11055);
nor U12646 (N_12646,N_10544,N_10029);
or U12647 (N_12647,N_10838,N_9832);
nand U12648 (N_12648,N_11938,N_11286);
xnor U12649 (N_12649,N_10957,N_10593);
and U12650 (N_12650,N_11184,N_12268);
and U12651 (N_12651,N_10224,N_9995);
and U12652 (N_12652,N_12301,N_11360);
or U12653 (N_12653,N_10617,N_10314);
xnor U12654 (N_12654,N_10085,N_11929);
nand U12655 (N_12655,N_9693,N_11161);
nand U12656 (N_12656,N_12212,N_11082);
xor U12657 (N_12657,N_9716,N_10779);
or U12658 (N_12658,N_11539,N_10647);
nand U12659 (N_12659,N_12219,N_12121);
nand U12660 (N_12660,N_12255,N_10996);
nand U12661 (N_12661,N_9471,N_10216);
and U12662 (N_12662,N_10642,N_10761);
nor U12663 (N_12663,N_10278,N_9708);
nor U12664 (N_12664,N_10458,N_11640);
and U12665 (N_12665,N_11226,N_11089);
nand U12666 (N_12666,N_12045,N_11888);
nor U12667 (N_12667,N_11239,N_11840);
and U12668 (N_12668,N_11160,N_11742);
nor U12669 (N_12669,N_10295,N_11033);
xor U12670 (N_12670,N_10293,N_10890);
and U12671 (N_12671,N_10798,N_9898);
nand U12672 (N_12672,N_11336,N_11835);
xnor U12673 (N_12673,N_10710,N_10644);
nor U12674 (N_12674,N_9980,N_9989);
nor U12675 (N_12675,N_11965,N_11817);
nor U12676 (N_12676,N_10817,N_9951);
nor U12677 (N_12677,N_11127,N_12350);
and U12678 (N_12678,N_10829,N_12478);
and U12679 (N_12679,N_10102,N_10532);
and U12680 (N_12680,N_11707,N_11141);
nand U12681 (N_12681,N_9536,N_9956);
xnor U12682 (N_12682,N_12080,N_12469);
nand U12683 (N_12683,N_11969,N_10079);
nand U12684 (N_12684,N_12482,N_11266);
nor U12685 (N_12685,N_11344,N_12155);
nor U12686 (N_12686,N_12333,N_10184);
or U12687 (N_12687,N_12140,N_10419);
nor U12688 (N_12688,N_9763,N_11072);
nand U12689 (N_12689,N_11186,N_9696);
nand U12690 (N_12690,N_11222,N_9377);
nor U12691 (N_12691,N_10280,N_10718);
nor U12692 (N_12692,N_11604,N_9913);
and U12693 (N_12693,N_9756,N_11673);
or U12694 (N_12694,N_10959,N_10704);
and U12695 (N_12695,N_11131,N_9619);
nand U12696 (N_12696,N_12162,N_11389);
nor U12697 (N_12697,N_11592,N_11400);
xnor U12698 (N_12698,N_9701,N_12198);
nor U12699 (N_12699,N_11206,N_10871);
nand U12700 (N_12700,N_10953,N_10171);
nand U12701 (N_12701,N_9480,N_9997);
nand U12702 (N_12702,N_9793,N_11208);
xnor U12703 (N_12703,N_9848,N_11977);
nand U12704 (N_12704,N_9667,N_11021);
nor U12705 (N_12705,N_11613,N_9742);
or U12706 (N_12706,N_11862,N_9819);
nand U12707 (N_12707,N_11125,N_11112);
xnor U12708 (N_12708,N_11858,N_11546);
xnor U12709 (N_12709,N_10612,N_10949);
nand U12710 (N_12710,N_10403,N_10531);
nor U12711 (N_12711,N_10193,N_10109);
xnor U12712 (N_12712,N_10436,N_9648);
and U12713 (N_12713,N_11191,N_9702);
nand U12714 (N_12714,N_11734,N_9838);
nor U12715 (N_12715,N_12384,N_12040);
and U12716 (N_12716,N_11532,N_9817);
and U12717 (N_12717,N_10059,N_11830);
and U12718 (N_12718,N_12493,N_9544);
or U12719 (N_12719,N_10627,N_11241);
nand U12720 (N_12720,N_9607,N_12370);
nor U12721 (N_12721,N_9788,N_11018);
and U12722 (N_12722,N_9446,N_9719);
nor U12723 (N_12723,N_11354,N_11232);
nand U12724 (N_12724,N_11932,N_11427);
or U12725 (N_12725,N_11797,N_9890);
nand U12726 (N_12726,N_9770,N_9875);
and U12727 (N_12727,N_10757,N_11598);
nand U12728 (N_12728,N_10666,N_10115);
xor U12729 (N_12729,N_9927,N_11798);
and U12730 (N_12730,N_10619,N_11881);
xnor U12731 (N_12731,N_12259,N_10424);
nor U12732 (N_12732,N_9439,N_11255);
and U12733 (N_12733,N_11855,N_11105);
or U12734 (N_12734,N_9475,N_10279);
and U12735 (N_12735,N_10206,N_10306);
and U12736 (N_12736,N_11966,N_11192);
nand U12737 (N_12737,N_11706,N_10487);
or U12738 (N_12738,N_11869,N_11263);
or U12739 (N_12739,N_11094,N_10652);
xnor U12740 (N_12740,N_9751,N_9772);
and U12741 (N_12741,N_9723,N_10646);
nand U12742 (N_12742,N_12109,N_12000);
xnor U12743 (N_12743,N_10307,N_10283);
xor U12744 (N_12744,N_10929,N_10506);
xnor U12745 (N_12745,N_9632,N_11507);
nand U12746 (N_12746,N_11579,N_10889);
and U12747 (N_12747,N_10743,N_10001);
nor U12748 (N_12748,N_11133,N_11210);
xor U12749 (N_12749,N_9579,N_10510);
nor U12750 (N_12750,N_10951,N_10490);
and U12751 (N_12751,N_10119,N_11137);
or U12752 (N_12752,N_11010,N_10522);
xnor U12753 (N_12753,N_9806,N_10106);
nand U12754 (N_12754,N_11346,N_9577);
nor U12755 (N_12755,N_10089,N_10651);
and U12756 (N_12756,N_9758,N_12049);
nor U12757 (N_12757,N_12465,N_10069);
nor U12758 (N_12758,N_10947,N_10005);
nand U12759 (N_12759,N_12060,N_9388);
nand U12760 (N_12760,N_10324,N_11303);
nand U12761 (N_12761,N_10804,N_11297);
xor U12762 (N_12762,N_12285,N_11409);
and U12763 (N_12763,N_11465,N_11200);
nand U12764 (N_12764,N_11819,N_10898);
nor U12765 (N_12765,N_11322,N_11547);
xor U12766 (N_12766,N_11426,N_12437);
nor U12767 (N_12767,N_11328,N_10084);
or U12768 (N_12768,N_10348,N_9949);
nand U12769 (N_12769,N_9589,N_12211);
or U12770 (N_12770,N_12218,N_10445);
xnor U12771 (N_12771,N_11848,N_9919);
xnor U12772 (N_12772,N_10988,N_9820);
nor U12773 (N_12773,N_10363,N_10113);
or U12774 (N_12774,N_12378,N_11772);
nor U12775 (N_12775,N_10591,N_9976);
nor U12776 (N_12776,N_9861,N_9881);
or U12777 (N_12777,N_11674,N_11001);
xor U12778 (N_12778,N_12048,N_10800);
and U12779 (N_12779,N_11670,N_10485);
or U12780 (N_12780,N_11924,N_11656);
nor U12781 (N_12781,N_11544,N_9664);
nand U12782 (N_12782,N_10006,N_10053);
xor U12783 (N_12783,N_9510,N_11714);
and U12784 (N_12784,N_10794,N_9532);
nor U12785 (N_12785,N_10713,N_10287);
xnor U12786 (N_12786,N_9409,N_10474);
nor U12787 (N_12787,N_9933,N_9625);
and U12788 (N_12788,N_9437,N_12074);
xor U12789 (N_12789,N_9730,N_11189);
and U12790 (N_12790,N_11281,N_10555);
xnor U12791 (N_12791,N_10196,N_9671);
nand U12792 (N_12792,N_10136,N_11851);
nor U12793 (N_12793,N_12095,N_10178);
nor U12794 (N_12794,N_11750,N_10970);
nor U12795 (N_12795,N_10357,N_10819);
nor U12796 (N_12796,N_11058,N_10263);
or U12797 (N_12797,N_9798,N_11267);
and U12798 (N_12798,N_11065,N_10158);
xor U12799 (N_12799,N_11319,N_9743);
and U12800 (N_12800,N_11139,N_11690);
and U12801 (N_12801,N_10176,N_10601);
and U12802 (N_12802,N_11875,N_11867);
nor U12803 (N_12803,N_11619,N_11775);
xnor U12804 (N_12804,N_10442,N_9922);
nor U12805 (N_12805,N_10180,N_11052);
nand U12806 (N_12806,N_11955,N_9586);
or U12807 (N_12807,N_11647,N_10459);
or U12808 (N_12808,N_10473,N_10168);
xor U12809 (N_12809,N_10905,N_9727);
or U12810 (N_12810,N_11220,N_11243);
xnor U12811 (N_12811,N_11727,N_11134);
xnor U12812 (N_12812,N_12310,N_10373);
and U12813 (N_12813,N_11559,N_12295);
nand U12814 (N_12814,N_11448,N_10845);
xnor U12815 (N_12815,N_10896,N_11412);
or U12816 (N_12816,N_12123,N_10660);
xnor U12817 (N_12817,N_12279,N_12415);
nor U12818 (N_12818,N_11996,N_10320);
and U12819 (N_12819,N_9618,N_9842);
and U12820 (N_12820,N_11904,N_9390);
xor U12821 (N_12821,N_9410,N_11658);
or U12822 (N_12822,N_10937,N_11558);
or U12823 (N_12823,N_9979,N_9613);
or U12824 (N_12824,N_10463,N_10537);
nor U12825 (N_12825,N_9415,N_11121);
or U12826 (N_12826,N_12451,N_11485);
and U12827 (N_12827,N_10528,N_12137);
and U12828 (N_12828,N_9519,N_10769);
or U12829 (N_12829,N_11590,N_12222);
or U12830 (N_12830,N_10610,N_11918);
nor U12831 (N_12831,N_12035,N_9498);
xor U12832 (N_12832,N_12307,N_10046);
nand U12833 (N_12833,N_10847,N_9414);
nand U12834 (N_12834,N_9562,N_10302);
nor U12835 (N_12835,N_9647,N_11803);
or U12836 (N_12836,N_11629,N_12239);
and U12837 (N_12837,N_12010,N_12369);
nor U12838 (N_12838,N_10840,N_10616);
or U12839 (N_12839,N_10602,N_11972);
or U12840 (N_12840,N_11649,N_9749);
nor U12841 (N_12841,N_12455,N_11390);
nor U12842 (N_12842,N_10276,N_9681);
nor U12843 (N_12843,N_12019,N_10692);
xor U12844 (N_12844,N_10270,N_11779);
or U12845 (N_12845,N_11873,N_11951);
nand U12846 (N_12846,N_11859,N_11806);
and U12847 (N_12847,N_11925,N_9810);
nand U12848 (N_12848,N_9752,N_12416);
xnor U12849 (N_12849,N_11540,N_12261);
nor U12850 (N_12850,N_9614,N_11275);
nand U12851 (N_12851,N_11111,N_10738);
nand U12852 (N_12852,N_12336,N_11070);
xnor U12853 (N_12853,N_10179,N_10497);
xnor U12854 (N_12854,N_9736,N_10766);
or U12855 (N_12855,N_10796,N_12340);
and U12856 (N_12856,N_11403,N_12143);
nor U12857 (N_12857,N_12387,N_11870);
nor U12858 (N_12858,N_12431,N_10200);
nor U12859 (N_12859,N_9401,N_10778);
and U12860 (N_12860,N_9815,N_11251);
nand U12861 (N_12861,N_9876,N_10821);
or U12862 (N_12862,N_10464,N_11307);
or U12863 (N_12863,N_10043,N_10126);
nor U12864 (N_12864,N_10254,N_9393);
nor U12865 (N_12865,N_10068,N_12447);
nand U12866 (N_12866,N_11337,N_10645);
xnor U12867 (N_12867,N_9462,N_9797);
or U12868 (N_12868,N_11549,N_9900);
or U12869 (N_12869,N_10221,N_9996);
nand U12870 (N_12870,N_11877,N_11093);
nand U12871 (N_12871,N_9986,N_9744);
or U12872 (N_12872,N_12072,N_11049);
or U12873 (N_12873,N_12099,N_12118);
or U12874 (N_12874,N_10944,N_12267);
or U12875 (N_12875,N_11476,N_9485);
nand U12876 (N_12876,N_10223,N_9703);
nor U12877 (N_12877,N_12214,N_11684);
xor U12878 (N_12878,N_10886,N_11444);
nor U12879 (N_12879,N_11339,N_11978);
or U12880 (N_12880,N_11726,N_12092);
xnor U12881 (N_12881,N_9773,N_10303);
xor U12882 (N_12882,N_9893,N_12495);
xor U12883 (N_12883,N_9382,N_10595);
nor U12884 (N_12884,N_11228,N_11363);
and U12885 (N_12885,N_11909,N_9704);
xnor U12886 (N_12886,N_11442,N_10325);
or U12887 (N_12887,N_9928,N_12246);
nand U12888 (N_12888,N_12202,N_11756);
nand U12889 (N_12889,N_9745,N_11057);
or U12890 (N_12890,N_10099,N_9522);
and U12891 (N_12891,N_9606,N_11741);
nor U12892 (N_12892,N_12225,N_12287);
xnor U12893 (N_12893,N_10620,N_10391);
nand U12894 (N_12894,N_10575,N_11466);
nor U12895 (N_12895,N_11379,N_9481);
nor U12896 (N_12896,N_9561,N_11494);
and U12897 (N_12897,N_11576,N_10316);
nor U12898 (N_12898,N_11378,N_10706);
nor U12899 (N_12899,N_10454,N_9538);
and U12900 (N_12900,N_10777,N_11535);
nor U12901 (N_12901,N_10654,N_9588);
or U12902 (N_12902,N_10569,N_11433);
nor U12903 (N_12903,N_10900,N_10140);
nor U12904 (N_12904,N_10913,N_11015);
nand U12905 (N_12905,N_10879,N_10904);
nand U12906 (N_12906,N_10406,N_11198);
or U12907 (N_12907,N_9837,N_10020);
nand U12908 (N_12908,N_11516,N_11475);
xnor U12909 (N_12909,N_12382,N_9698);
xnor U12910 (N_12910,N_12017,N_12107);
xnor U12911 (N_12911,N_10669,N_9649);
xnor U12912 (N_12912,N_9566,N_10767);
or U12913 (N_12913,N_11016,N_11829);
xor U12914 (N_12914,N_11473,N_11868);
xnor U12915 (N_12915,N_10737,N_9665);
nor U12916 (N_12916,N_11815,N_11188);
xnor U12917 (N_12917,N_11260,N_10736);
xor U12918 (N_12918,N_11813,N_12473);
and U12919 (N_12919,N_9534,N_10351);
and U12920 (N_12920,N_10417,N_10447);
and U12921 (N_12921,N_10443,N_10500);
nand U12922 (N_12922,N_10183,N_10942);
and U12923 (N_12923,N_12142,N_9957);
and U12924 (N_12924,N_9594,N_10201);
nand U12925 (N_12925,N_11405,N_10199);
nand U12926 (N_12926,N_9474,N_12311);
xnor U12927 (N_12927,N_11902,N_11294);
or U12928 (N_12928,N_10261,N_11047);
xnor U12929 (N_12929,N_10613,N_12464);
and U12930 (N_12930,N_9912,N_10259);
or U12931 (N_12931,N_11982,N_9809);
nand U12932 (N_12932,N_12161,N_9795);
nand U12933 (N_12933,N_10630,N_10498);
nor U12934 (N_12934,N_9882,N_10786);
xnor U12935 (N_12935,N_11760,N_9528);
nor U12936 (N_12936,N_11528,N_12302);
or U12937 (N_12937,N_10087,N_12423);
nand U12938 (N_12938,N_11253,N_11689);
and U12939 (N_12939,N_10980,N_9541);
nor U12940 (N_12940,N_11235,N_9405);
nand U12941 (N_12941,N_9582,N_12147);
nor U12942 (N_12942,N_12070,N_11114);
xor U12943 (N_12943,N_11890,N_11833);
nand U12944 (N_12944,N_12023,N_10922);
or U12945 (N_12945,N_10739,N_10665);
and U12946 (N_12946,N_10984,N_12317);
xor U12947 (N_12947,N_11419,N_12324);
nand U12948 (N_12948,N_10289,N_11926);
nand U12949 (N_12949,N_9943,N_11062);
or U12950 (N_12950,N_10477,N_11812);
and U12951 (N_12951,N_10993,N_10958);
xor U12952 (N_12952,N_9472,N_11668);
nor U12953 (N_12953,N_10994,N_12009);
xor U12954 (N_12954,N_10892,N_12368);
nor U12955 (N_12955,N_11878,N_10217);
or U12956 (N_12956,N_10860,N_12321);
or U12957 (N_12957,N_11754,N_11115);
and U12958 (N_12958,N_9822,N_10679);
or U12959 (N_12959,N_10407,N_9559);
xnor U12960 (N_12960,N_10038,N_10203);
and U12961 (N_12961,N_12312,N_9600);
xnor U12962 (N_12962,N_10013,N_9500);
nand U12963 (N_12963,N_11770,N_9878);
or U12964 (N_12964,N_10992,N_10598);
nor U12965 (N_12965,N_9602,N_10983);
and U12966 (N_12966,N_10205,N_11157);
nand U12967 (N_12967,N_9914,N_11602);
nor U12968 (N_12968,N_10333,N_10116);
xnor U12969 (N_12969,N_9761,N_11386);
nand U12970 (N_12970,N_9969,N_9673);
and U12971 (N_12971,N_11633,N_11037);
xnor U12972 (N_12972,N_12006,N_11749);
nand U12973 (N_12973,N_9846,N_9461);
or U12974 (N_12974,N_12127,N_12256);
and U12975 (N_12975,N_10551,N_11823);
nand U12976 (N_12976,N_12260,N_11099);
and U12977 (N_12977,N_11459,N_9952);
nand U12978 (N_12978,N_9489,N_12264);
or U12979 (N_12979,N_11343,N_12245);
nand U12980 (N_12980,N_10065,N_9635);
xnor U12981 (N_12981,N_12342,N_10097);
nand U12982 (N_12982,N_10138,N_9915);
and U12983 (N_12983,N_12289,N_10262);
xor U12984 (N_12984,N_11150,N_9948);
nand U12985 (N_12985,N_11142,N_11901);
nor U12986 (N_12986,N_9622,N_9504);
nand U12987 (N_12987,N_10060,N_10714);
nand U12988 (N_12988,N_11364,N_9569);
nor U12989 (N_12989,N_11710,N_10733);
nor U12990 (N_12990,N_11006,N_10960);
and U12991 (N_12991,N_11169,N_11652);
or U12992 (N_12992,N_10828,N_12250);
nand U12993 (N_12993,N_11743,N_12004);
and U12994 (N_12994,N_11456,N_9685);
and U12995 (N_12995,N_10034,N_9378);
nand U12996 (N_12996,N_11591,N_12435);
nand U12997 (N_12997,N_11510,N_12192);
nor U12998 (N_12998,N_10375,N_11638);
and U12999 (N_12999,N_11983,N_11923);
xor U13000 (N_13000,N_9609,N_11511);
nor U13001 (N_13001,N_9905,N_11355);
and U13002 (N_13002,N_10174,N_9887);
xnor U13003 (N_13003,N_11147,N_10425);
xnor U13004 (N_13004,N_11330,N_12458);
and U13005 (N_13005,N_11257,N_10000);
nand U13006 (N_13006,N_10527,N_10021);
nand U13007 (N_13007,N_9403,N_11555);
or U13008 (N_13008,N_10211,N_11118);
xor U13009 (N_13009,N_9764,N_10604);
or U13010 (N_13010,N_10272,N_11025);
nor U13011 (N_13011,N_11564,N_11035);
or U13012 (N_13012,N_10475,N_10160);
nand U13013 (N_13013,N_11007,N_11588);
nor U13014 (N_13014,N_11891,N_11414);
nand U13015 (N_13015,N_11653,N_9521);
xnor U13016 (N_13016,N_9916,N_9486);
or U13017 (N_13017,N_11595,N_12188);
nor U13018 (N_13018,N_10299,N_12400);
and U13019 (N_13019,N_10823,N_11661);
nand U13020 (N_13020,N_10514,N_12441);
nor U13021 (N_13021,N_11686,N_12234);
xnor U13022 (N_13022,N_10626,N_11201);
or U13023 (N_13023,N_11711,N_11836);
xor U13024 (N_13024,N_12160,N_10494);
xnor U13025 (N_13025,N_9808,N_12197);
nor U13026 (N_13026,N_10853,N_11327);
or U13027 (N_13027,N_10340,N_12226);
xnor U13028 (N_13028,N_11831,N_12283);
or U13029 (N_13029,N_10260,N_10636);
nand U13030 (N_13030,N_9964,N_9970);
nor U13031 (N_13031,N_11611,N_12244);
nor U13032 (N_13032,N_9592,N_10018);
nand U13033 (N_13033,N_11764,N_12124);
and U13034 (N_13034,N_11042,N_9851);
or U13035 (N_13035,N_12332,N_11247);
and U13036 (N_13036,N_10930,N_9766);
xor U13037 (N_13037,N_9930,N_10142);
nor U13038 (N_13038,N_12230,N_11348);
nand U13039 (N_13039,N_11101,N_11846);
nor U13040 (N_13040,N_11985,N_11722);
or U13041 (N_13041,N_12149,N_11026);
nor U13042 (N_13042,N_11318,N_11217);
nand U13043 (N_13043,N_12399,N_10120);
xor U13044 (N_13044,N_10549,N_11762);
nor U13045 (N_13045,N_12236,N_10912);
xor U13046 (N_13046,N_9807,N_9389);
nand U13047 (N_13047,N_11406,N_11769);
xnor U13048 (N_13048,N_11036,N_11863);
nor U13049 (N_13049,N_9558,N_10344);
xor U13050 (N_13050,N_10215,N_9570);
nor U13051 (N_13051,N_11240,N_12097);
nor U13052 (N_13052,N_12293,N_9885);
nand U13053 (N_13053,N_10368,N_9643);
and U13054 (N_13054,N_10231,N_9529);
or U13055 (N_13055,N_10502,N_11103);
xor U13056 (N_13056,N_9960,N_11000);
nor U13057 (N_13057,N_9857,N_11560);
and U13058 (N_13058,N_10249,N_9540);
or U13059 (N_13059,N_11704,N_10366);
or U13060 (N_13060,N_11497,N_11331);
xnor U13061 (N_13061,N_12485,N_12304);
and U13062 (N_13062,N_11372,N_11723);
xor U13063 (N_13063,N_10039,N_9852);
xor U13064 (N_13064,N_9733,N_11436);
or U13065 (N_13065,N_9940,N_11504);
nor U13066 (N_13066,N_12168,N_10481);
and U13067 (N_13067,N_10253,N_11900);
nor U13068 (N_13068,N_9934,N_10460);
and U13069 (N_13069,N_9408,N_10322);
nor U13070 (N_13070,N_9824,N_11498);
nor U13071 (N_13071,N_11527,N_9712);
or U13072 (N_13072,N_12221,N_11071);
xnor U13073 (N_13073,N_9825,N_12089);
and U13074 (N_13074,N_11135,N_11991);
nor U13075 (N_13075,N_9515,N_10394);
xnor U13076 (N_13076,N_12281,N_10526);
nand U13077 (N_13077,N_10478,N_10377);
and U13078 (N_13078,N_11648,N_9958);
nand U13079 (N_13079,N_11215,N_12051);
xnor U13080 (N_13080,N_11906,N_10818);
and U13081 (N_13081,N_10650,N_11671);
nand U13082 (N_13082,N_11092,N_11946);
and U13083 (N_13083,N_12131,N_10715);
and U13084 (N_13084,N_10288,N_11277);
and U13085 (N_13085,N_12357,N_11044);
xor U13086 (N_13086,N_10702,N_9590);
or U13087 (N_13087,N_9460,N_9513);
and U13088 (N_13088,N_11313,N_9535);
or U13089 (N_13089,N_11672,N_11799);
or U13090 (N_13090,N_10347,N_12249);
nand U13091 (N_13091,N_11090,N_12446);
xor U13092 (N_13092,N_10045,N_12330);
nor U13093 (N_13093,N_10883,N_10237);
nand U13094 (N_13094,N_9855,N_10047);
xor U13095 (N_13095,N_12410,N_10504);
nor U13096 (N_13096,N_9983,N_11411);
and U13097 (N_13097,N_10894,N_10875);
nor U13098 (N_13098,N_12203,N_12363);
nand U13099 (N_13099,N_12282,N_10573);
and U13100 (N_13100,N_10248,N_12057);
or U13101 (N_13101,N_9821,N_11271);
and U13102 (N_13102,N_10839,N_11884);
nor U13103 (N_13103,N_11538,N_10063);
or U13104 (N_13104,N_10681,N_9687);
xor U13105 (N_13105,N_10396,N_10427);
nor U13106 (N_13106,N_11980,N_10037);
or U13107 (N_13107,N_10705,N_10916);
nor U13108 (N_13108,N_9897,N_9465);
and U13109 (N_13109,N_11626,N_12186);
and U13110 (N_13110,N_9938,N_11597);
or U13111 (N_13111,N_11566,N_11854);
and U13112 (N_13112,N_9714,N_10027);
xor U13113 (N_13113,N_12117,N_12031);
or U13114 (N_13114,N_12030,N_10100);
and U13115 (N_13115,N_11765,N_12398);
nor U13116 (N_13116,N_12079,N_11523);
xor U13117 (N_13117,N_11197,N_11306);
nor U13118 (N_13118,N_11834,N_9850);
nor U13119 (N_13119,N_10155,N_12253);
nand U13120 (N_13120,N_10452,N_11586);
nor U13121 (N_13121,N_9402,N_10884);
and U13122 (N_13122,N_10235,N_11695);
nor U13123 (N_13123,N_11713,N_12024);
or U13124 (N_13124,N_12381,N_11418);
xor U13125 (N_13125,N_12001,N_12014);
or U13126 (N_13126,N_11178,N_9684);
xor U13127 (N_13127,N_10525,N_11308);
nand U13128 (N_13128,N_11826,N_10732);
nand U13129 (N_13129,N_10195,N_10264);
xor U13130 (N_13130,N_11631,N_9604);
nand U13131 (N_13131,N_10450,N_10023);
nor U13132 (N_13132,N_11064,N_10740);
xnor U13133 (N_13133,N_11600,N_11811);
nand U13134 (N_13134,N_10606,N_11931);
nand U13135 (N_13135,N_12355,N_10717);
xor U13136 (N_13136,N_11361,N_9478);
xnor U13137 (N_13137,N_11245,N_9918);
xnor U13138 (N_13138,N_10004,N_12044);
nor U13139 (N_13139,N_12078,N_10359);
nor U13140 (N_13140,N_10999,N_11957);
xor U13141 (N_13141,N_9777,N_9497);
and U13142 (N_13142,N_9463,N_10938);
or U13143 (N_13143,N_10965,N_11612);
xor U13144 (N_13144,N_12273,N_11278);
xor U13145 (N_13145,N_11259,N_11288);
nand U13146 (N_13146,N_11144,N_11919);
and U13147 (N_13147,N_11818,N_11223);
xnor U13148 (N_13148,N_10014,N_12318);
or U13149 (N_13149,N_11187,N_10343);
or U13150 (N_13150,N_10887,N_10104);
xor U13151 (N_13151,N_11369,N_11804);
or U13152 (N_13152,N_12265,N_10387);
nand U13153 (N_13153,N_10415,N_11782);
nand U13154 (N_13154,N_11948,N_10255);
and U13155 (N_13155,N_11839,N_11615);
xnor U13156 (N_13156,N_10583,N_10973);
xnor U13157 (N_13157,N_11505,N_11124);
xor U13158 (N_13158,N_11249,N_12367);
nor U13159 (N_13159,N_10429,N_11897);
nor U13160 (N_13160,N_10846,N_10592);
nand U13161 (N_13161,N_10906,N_9877);
nor U13162 (N_13162,N_9760,N_11565);
and U13163 (N_13163,N_11916,N_12323);
and U13164 (N_13164,N_11651,N_12290);
nor U13165 (N_13165,N_9710,N_10691);
or U13166 (N_13166,N_10741,N_11181);
and U13167 (N_13167,N_10139,N_12185);
nor U13168 (N_13168,N_10934,N_10600);
nand U13169 (N_13169,N_9705,N_9543);
or U13170 (N_13170,N_12271,N_11999);
xnor U13171 (N_13171,N_10421,N_11876);
nor U13172 (N_13172,N_10008,N_11349);
or U13173 (N_13173,N_10848,N_11552);
and U13174 (N_13174,N_10011,N_12278);
nand U13175 (N_13175,N_11404,N_9672);
or U13176 (N_13176,N_10788,N_10716);
and U13177 (N_13177,N_9599,N_10123);
or U13178 (N_13178,N_10917,N_10156);
and U13179 (N_13179,N_10678,N_10932);
nor U13180 (N_13180,N_11159,N_10243);
xnor U13181 (N_13181,N_12426,N_9484);
or U13182 (N_13182,N_11503,N_11524);
and U13183 (N_13183,N_11847,N_11896);
xor U13184 (N_13184,N_11699,N_11634);
or U13185 (N_13185,N_11513,N_11989);
nor U13186 (N_13186,N_10785,N_12372);
xor U13187 (N_13187,N_11156,N_9458);
and U13188 (N_13188,N_11587,N_9653);
or U13189 (N_13189,N_9884,N_10955);
or U13190 (N_13190,N_11637,N_12180);
nand U13191 (N_13191,N_10878,N_11441);
nor U13192 (N_13192,N_10812,N_12171);
nor U13193 (N_13193,N_12274,N_11574);
nor U13194 (N_13194,N_11079,N_9610);
or U13195 (N_13195,N_12216,N_10869);
xnor U13196 (N_13196,N_9971,N_10759);
and U13197 (N_13197,N_12195,N_10317);
nor U13198 (N_13198,N_12102,N_9843);
xor U13199 (N_13199,N_11117,N_9438);
nor U13200 (N_13200,N_11454,N_9468);
and U13201 (N_13201,N_10159,N_10362);
xor U13202 (N_13202,N_9988,N_10667);
or U13203 (N_13203,N_10055,N_9549);
nor U13204 (N_13204,N_10220,N_9858);
or U13205 (N_13205,N_10028,N_11915);
or U13206 (N_13206,N_11087,N_11061);
xnor U13207 (N_13207,N_9924,N_11899);
or U13208 (N_13208,N_10784,N_12213);
nor U13209 (N_13209,N_10148,N_9491);
and U13210 (N_13210,N_12490,N_10998);
nor U13211 (N_13211,N_12052,N_9732);
nand U13212 (N_13212,N_10435,N_10493);
nand U13213 (N_13213,N_10843,N_10050);
nand U13214 (N_13214,N_12360,N_10010);
and U13215 (N_13215,N_10770,N_10192);
nor U13216 (N_13216,N_12499,N_12496);
and U13217 (N_13217,N_10833,N_9962);
or U13218 (N_13218,N_10304,N_9677);
xor U13219 (N_13219,N_11802,N_9706);
or U13220 (N_13220,N_10850,N_11643);
nand U13221 (N_13221,N_11167,N_10327);
or U13222 (N_13222,N_9738,N_12033);
xor U13223 (N_13223,N_12038,N_12034);
and U13224 (N_13224,N_10685,N_11942);
or U13225 (N_13225,N_9533,N_10353);
nand U13226 (N_13226,N_11913,N_10772);
and U13227 (N_13227,N_10931,N_12073);
or U13228 (N_13228,N_10933,N_10920);
nor U13229 (N_13229,N_11575,N_11279);
and U13230 (N_13230,N_11777,N_9662);
or U13231 (N_13231,N_9923,N_10381);
nor U13232 (N_13232,N_9802,N_10194);
xor U13233 (N_13233,N_11234,N_9617);
or U13234 (N_13234,N_11113,N_11660);
and U13235 (N_13235,N_11622,N_10358);
nor U13236 (N_13236,N_10392,N_10731);
and U13237 (N_13237,N_11562,N_11976);
and U13238 (N_13238,N_9565,N_11205);
xnor U13239 (N_13239,N_11824,N_9982);
nand U13240 (N_13240,N_9512,N_10842);
and U13241 (N_13241,N_12454,N_10480);
xor U13242 (N_13242,N_11808,N_11373);
nor U13243 (N_13243,N_9400,N_9436);
or U13244 (N_13244,N_11457,N_12272);
nor U13245 (N_13245,N_10432,N_10507);
and U13246 (N_13246,N_10564,N_9697);
xor U13247 (N_13247,N_11353,N_11788);
nor U13248 (N_13248,N_12237,N_10401);
or U13249 (N_13249,N_10816,N_9961);
xnor U13250 (N_13250,N_12228,N_11543);
nor U13251 (N_13251,N_12391,N_11721);
xnor U13252 (N_13252,N_11083,N_11501);
nand U13253 (N_13253,N_10247,N_10643);
or U13254 (N_13254,N_11728,N_10125);
and U13255 (N_13255,N_9841,N_10455);
nor U13256 (N_13256,N_11347,N_9487);
and U13257 (N_13257,N_9434,N_9676);
nor U13258 (N_13258,N_12462,N_12327);
nor U13259 (N_13259,N_10807,N_12477);
and U13260 (N_13260,N_11086,N_10689);
nor U13261 (N_13261,N_9774,N_12207);
or U13262 (N_13262,N_11388,N_10165);
xnor U13263 (N_13263,N_10457,N_11274);
and U13264 (N_13264,N_11449,N_11022);
xnor U13265 (N_13265,N_10815,N_11050);
and U13266 (N_13266,N_11309,N_10400);
and U13267 (N_13267,N_12320,N_10694);
and U13268 (N_13268,N_10559,N_12166);
nor U13269 (N_13269,N_10177,N_10040);
and U13270 (N_13270,N_10052,N_12385);
xnor U13271 (N_13271,N_10378,N_11794);
and U13272 (N_13272,N_11905,N_10488);
nor U13273 (N_13273,N_11359,N_12427);
and U13274 (N_13274,N_12397,N_11295);
nand U13275 (N_13275,N_10117,N_10721);
xor U13276 (N_13276,N_11979,N_12269);
nor U13277 (N_13277,N_10893,N_10354);
and U13278 (N_13278,N_11827,N_10131);
nor U13279 (N_13279,N_9420,N_10873);
xor U13280 (N_13280,N_10789,N_12215);
nor U13281 (N_13281,N_9479,N_11735);
nor U13282 (N_13282,N_12438,N_11236);
xnor U13283 (N_13283,N_10775,N_10127);
xor U13284 (N_13284,N_11949,N_11168);
xor U13285 (N_13285,N_12414,N_9926);
nor U13286 (N_13286,N_12075,N_11039);
nand U13287 (N_13287,N_12439,N_11356);
nand U13288 (N_13288,N_12315,N_10639);
nand U13289 (N_13289,N_10599,N_10605);
nand U13290 (N_13290,N_9670,N_11805);
and U13291 (N_13291,N_9692,N_12442);
xnor U13292 (N_13292,N_9636,N_9896);
or U13293 (N_13293,N_9966,N_10758);
nor U13294 (N_13294,N_12375,N_11262);
nand U13295 (N_13295,N_10897,N_10699);
or U13296 (N_13296,N_11415,N_10153);
nor U13297 (N_13297,N_12243,N_12088);
nand U13298 (N_13298,N_11129,N_10535);
nand U13299 (N_13299,N_12128,N_11264);
and U13300 (N_13300,N_9831,N_11323);
xor U13301 (N_13301,N_11500,N_9494);
nand U13302 (N_13302,N_12157,N_11301);
or U13303 (N_13303,N_10300,N_11822);
or U13304 (N_13304,N_10874,N_10703);
nand U13305 (N_13305,N_10019,N_10782);
and U13306 (N_13306,N_9659,N_10903);
xor U13307 (N_13307,N_12116,N_10730);
or U13308 (N_13308,N_12497,N_12425);
xor U13309 (N_13309,N_10298,N_10607);
or U13310 (N_13310,N_11043,N_10675);
nor U13311 (N_13311,N_10797,N_10437);
nand U13312 (N_13312,N_12276,N_10748);
nor U13313 (N_13313,N_11889,N_10746);
or U13314 (N_13314,N_9423,N_10383);
xor U13315 (N_13315,N_12316,N_12401);
xnor U13316 (N_13316,N_10308,N_11202);
or U13317 (N_13317,N_10546,N_10462);
or U13318 (N_13318,N_9661,N_11885);
nor U13319 (N_13319,N_9412,N_10628);
xnor U13320 (N_13320,N_11871,N_10456);
or U13321 (N_13321,N_11407,N_11185);
nand U13322 (N_13322,N_10208,N_10103);
or U13323 (N_13323,N_10925,N_12093);
xnor U13324 (N_13324,N_11338,N_10318);
and U13325 (N_13325,N_9612,N_10172);
nand U13326 (N_13326,N_9803,N_11557);
nand U13327 (N_13327,N_9715,N_12041);
nor U13328 (N_13328,N_9394,N_11212);
nor U13329 (N_13329,N_9419,N_9456);
nor U13330 (N_13330,N_12460,N_11767);
and U13331 (N_13331,N_11548,N_9424);
xor U13332 (N_13332,N_10948,N_10446);
xnor U13333 (N_13333,N_12393,N_12298);
xnor U13334 (N_13334,N_12150,N_12334);
nor U13335 (N_13335,N_12174,N_12082);
and U13336 (N_13336,N_9690,N_9539);
nor U13337 (N_13337,N_9906,N_10690);
nor U13338 (N_13338,N_9786,N_11095);
nand U13339 (N_13339,N_10822,N_11607);
nand U13340 (N_13340,N_10568,N_11688);
or U13341 (N_13341,N_10609,N_11059);
xnor U13342 (N_13342,N_12020,N_11635);
and U13343 (N_13343,N_11231,N_10041);
or U13344 (N_13344,N_9941,N_10633);
nor U13345 (N_13345,N_9844,N_12405);
nor U13346 (N_13346,N_10022,N_10070);
xor U13347 (N_13347,N_11171,N_11376);
nor U13348 (N_13348,N_10680,N_12319);
or U13349 (N_13349,N_9404,N_12135);
and U13350 (N_13350,N_9721,N_12235);
or U13351 (N_13351,N_10449,N_10064);
and U13352 (N_13352,N_11691,N_9526);
nand U13353 (N_13353,N_11663,N_12450);
nor U13354 (N_13354,N_12091,N_9455);
or U13355 (N_13355,N_12471,N_10389);
or U13356 (N_13356,N_11785,N_12068);
or U13357 (N_13357,N_9645,N_10560);
xor U13358 (N_13358,N_10831,N_10438);
or U13359 (N_13359,N_10711,N_10505);
xnor U13360 (N_13360,N_11054,N_10885);
xor U13361 (N_13361,N_10753,N_12306);
nand U13362 (N_13362,N_10461,N_11326);
nor U13363 (N_13363,N_12422,N_12139);
xnor U13364 (N_13364,N_10124,N_12448);
nand U13365 (N_13365,N_11746,N_12480);
nor U13366 (N_13366,N_11479,N_10371);
nor U13367 (N_13367,N_10030,N_10540);
nand U13368 (N_13368,N_10073,N_11384);
or U13369 (N_13369,N_10529,N_11737);
or U13370 (N_13370,N_11031,N_10856);
and U13371 (N_13371,N_12103,N_12086);
nand U13372 (N_13372,N_10911,N_12388);
and U13373 (N_13373,N_12418,N_11471);
nor U13374 (N_13374,N_10524,N_10975);
and U13375 (N_13375,N_9499,N_12184);
and U13376 (N_13376,N_11455,N_11486);
and U13377 (N_13377,N_10597,N_9683);
and U13378 (N_13378,N_10096,N_11002);
or U13379 (N_13379,N_12026,N_10062);
or U13380 (N_13380,N_12483,N_12467);
xor U13381 (N_13381,N_12475,N_10146);
and U13382 (N_13382,N_11657,N_10547);
and U13383 (N_13383,N_12347,N_11312);
xor U13384 (N_13384,N_10801,N_11489);
xnor U13385 (N_13385,N_12101,N_12286);
nor U13386 (N_13386,N_12335,N_9830);
nand U13387 (N_13387,N_9974,N_11908);
or U13388 (N_13388,N_9407,N_10024);
and U13389 (N_13389,N_11282,N_9849);
nand U13390 (N_13390,N_10752,N_11842);
and U13391 (N_13391,N_10058,N_12201);
and U13392 (N_13392,N_9581,N_11719);
and U13393 (N_13393,N_10150,N_10129);
or U13394 (N_13394,N_11759,N_10367);
and U13395 (N_13395,N_10631,N_10961);
and U13396 (N_13396,N_12389,N_12193);
or U13397 (N_13397,N_10380,N_10080);
xor U13398 (N_13398,N_11800,N_11702);
and U13399 (N_13399,N_9678,N_12136);
xnor U13400 (N_13400,N_12359,N_9399);
nand U13401 (N_13401,N_11175,N_10226);
nor U13402 (N_13402,N_9731,N_11238);
nand U13403 (N_13403,N_11708,N_12432);
nand U13404 (N_13404,N_9418,N_12251);
nor U13405 (N_13405,N_11680,N_12406);
nor U13406 (N_13406,N_11213,N_11366);
or U13407 (N_13407,N_11219,N_9411);
and U13408 (N_13408,N_11393,N_11960);
or U13409 (N_13409,N_11814,N_12409);
and U13410 (N_13410,N_12066,N_10971);
and U13411 (N_13411,N_12362,N_11753);
nand U13412 (N_13412,N_10756,N_11123);
nand U13413 (N_13413,N_9507,N_10423);
xnor U13414 (N_13414,N_11614,N_9932);
and U13415 (N_13415,N_11594,N_10167);
or U13416 (N_13416,N_10579,N_11886);
nand U13417 (N_13417,N_10810,N_11261);
xor U13418 (N_13418,N_9639,N_11450);
or U13419 (N_13419,N_11796,N_10157);
nand U13420 (N_13420,N_10182,N_10907);
nor U13421 (N_13421,N_11452,N_11128);
and U13422 (N_13422,N_9994,N_10439);
and U13423 (N_13423,N_12108,N_11654);
nor U13424 (N_13424,N_10754,N_10441);
and U13425 (N_13425,N_9642,N_11964);
nand U13426 (N_13426,N_11385,N_11487);
nand U13427 (N_13427,N_9724,N_10659);
or U13428 (N_13428,N_11182,N_10346);
xnor U13429 (N_13429,N_11298,N_10697);
nor U13430 (N_13430,N_11941,N_11484);
nor U13431 (N_13431,N_10384,N_11382);
and U13432 (N_13432,N_10083,N_9759);
or U13433 (N_13433,N_9637,N_12303);
nor U13434 (N_13434,N_9554,N_10112);
nand U13435 (N_13435,N_11646,N_11116);
or U13436 (N_13436,N_11074,N_9901);
nor U13437 (N_13437,N_10232,N_10556);
xor U13438 (N_13438,N_12208,N_11968);
nand U13439 (N_13439,N_12133,N_9725);
and U13440 (N_13440,N_11910,N_12377);
nand U13441 (N_13441,N_12339,N_11367);
nand U13442 (N_13442,N_12308,N_10941);
and U13443 (N_13443,N_11571,N_10708);
or U13444 (N_13444,N_11529,N_11787);
xnor U13445 (N_13445,N_10143,N_12257);
nand U13446 (N_13446,N_10727,N_12069);
or U13447 (N_13447,N_12288,N_11067);
nand U13448 (N_13448,N_10919,N_9587);
nand U13449 (N_13449,N_10867,N_9722);
and U13450 (N_13450,N_11194,N_11287);
or U13451 (N_13451,N_11304,N_10997);
xnor U13452 (N_13452,N_11705,N_9779);
and U13453 (N_13453,N_11758,N_10049);
and U13454 (N_13454,N_10868,N_12390);
nor U13455 (N_13455,N_11335,N_11724);
xnor U13456 (N_13456,N_10025,N_11340);
nor U13457 (N_13457,N_12346,N_10749);
nand U13458 (N_13458,N_10499,N_10902);
xor U13459 (N_13459,N_11664,N_11729);
nor U13460 (N_13460,N_11314,N_11791);
or U13461 (N_13461,N_11861,N_9531);
nand U13462 (N_13462,N_9518,N_10335);
nand U13463 (N_13463,N_11046,N_9865);
nor U13464 (N_13464,N_10265,N_10668);
and U13465 (N_13465,N_11216,N_10003);
or U13466 (N_13466,N_10326,N_12050);
and U13467 (N_13467,N_9555,N_11864);
or U13468 (N_13468,N_11225,N_11252);
nor U13469 (N_13469,N_11745,N_10790);
and U13470 (N_13470,N_9823,N_10899);
nor U13471 (N_13471,N_10489,N_10188);
and U13472 (N_13472,N_10809,N_12059);
nand U13473 (N_13473,N_9641,N_9987);
or U13474 (N_13474,N_12443,N_11447);
nand U13475 (N_13475,N_10061,N_10978);
xnor U13476 (N_13476,N_9907,N_10570);
and U13477 (N_13477,N_11019,N_9814);
xor U13478 (N_13478,N_10292,N_10648);
or U13479 (N_13479,N_12220,N_11434);
and U13480 (N_13480,N_12153,N_12191);
nand U13481 (N_13481,N_10519,N_11730);
nor U13482 (N_13482,N_11943,N_10924);
and U13483 (N_13483,N_10578,N_10742);
and U13484 (N_13484,N_10057,N_10301);
and U13485 (N_13485,N_11158,N_11850);
nand U13486 (N_13486,N_10338,N_9945);
or U13487 (N_13487,N_9386,N_9552);
nand U13488 (N_13488,N_11917,N_9623);
and U13489 (N_13489,N_11945,N_11474);
xor U13490 (N_13490,N_12434,N_11075);
and U13491 (N_13491,N_10350,N_12328);
or U13492 (N_13492,N_12277,N_11939);
nand U13493 (N_13493,N_9709,N_11431);
or U13494 (N_13494,N_11258,N_11820);
xor U13495 (N_13495,N_10273,N_10275);
or U13496 (N_13496,N_11623,N_10543);
nand U13497 (N_13497,N_11581,N_12182);
xor U13498 (N_13498,N_10799,N_10586);
xor U13499 (N_13499,N_10750,N_10137);
nor U13500 (N_13500,N_10832,N_10101);
nand U13501 (N_13501,N_12115,N_11214);
or U13502 (N_13502,N_12029,N_11172);
and U13503 (N_13503,N_9785,N_12305);
or U13504 (N_13504,N_10864,N_12196);
xnor U13505 (N_13505,N_10393,N_10258);
xor U13506 (N_13506,N_12173,N_9483);
and U13507 (N_13507,N_9473,N_12247);
nor U13508 (N_13508,N_11296,N_9640);
nand U13509 (N_13509,N_12156,N_11786);
nand U13510 (N_13510,N_11933,N_11569);
and U13511 (N_13511,N_10571,N_10236);
xor U13512 (N_13512,N_11003,N_12096);
nor U13513 (N_13513,N_11573,N_12110);
nand U13514 (N_13514,N_12413,N_11421);
xnor U13515 (N_13515,N_10550,N_10877);
xnor U13516 (N_13516,N_10281,N_9429);
nand U13517 (N_13517,N_10638,N_11550);
nor U13518 (N_13518,N_12356,N_10565);
nand U13519 (N_13519,N_10416,N_10448);
or U13520 (N_13520,N_11148,N_11577);
nand U13521 (N_13521,N_10212,N_9550);
nor U13522 (N_13522,N_11589,N_10834);
nor U13523 (N_13523,N_11081,N_10927);
xnor U13524 (N_13524,N_12054,N_9937);
or U13525 (N_13525,N_11437,N_12179);
xor U13526 (N_13526,N_11530,N_10081);
xnor U13527 (N_13527,N_12254,N_12011);
nor U13528 (N_13528,N_9944,N_12456);
xnor U13529 (N_13529,N_9892,N_9445);
nor U13530 (N_13530,N_11329,N_10946);
xor U13531 (N_13531,N_11108,N_12266);
xor U13532 (N_13532,N_12229,N_9859);
xnor U13533 (N_13533,N_11482,N_11733);
or U13534 (N_13534,N_12484,N_12085);
and U13535 (N_13535,N_10972,N_11617);
or U13536 (N_13536,N_10841,N_11620);
and U13537 (N_13537,N_11974,N_9754);
xnor U13538 (N_13538,N_12452,N_10332);
nand U13539 (N_13539,N_10186,N_9769);
or U13540 (N_13540,N_10269,N_11912);
or U13541 (N_13541,N_9381,N_11395);
nand U13542 (N_13542,N_10825,N_12436);
nor U13543 (N_13543,N_10305,N_10166);
xnor U13544 (N_13544,N_12113,N_10688);
nand U13545 (N_13545,N_11357,N_10857);
or U13546 (N_13546,N_10724,N_11321);
nor U13547 (N_13547,N_9840,N_12459);
xor U13548 (N_13548,N_10655,N_9689);
xor U13549 (N_13549,N_11284,N_11140);
nand U13550 (N_13550,N_12240,N_11422);
nand U13551 (N_13551,N_12491,N_10244);
nand U13552 (N_13552,N_11068,N_9576);
xnor U13553 (N_13553,N_11852,N_10603);
xnor U13554 (N_13554,N_9380,N_11293);
xor U13555 (N_13555,N_11265,N_10701);
nor U13556 (N_13556,N_10508,N_9750);
and U13557 (N_13557,N_9454,N_10982);
nor U13558 (N_13558,N_10566,N_10637);
or U13559 (N_13559,N_10376,N_11963);
and U13560 (N_13560,N_10672,N_10981);
xnor U13561 (N_13561,N_10414,N_10175);
nand U13562 (N_13562,N_11693,N_10355);
nand U13563 (N_13563,N_11077,N_9955);
and U13564 (N_13564,N_11398,N_11603);
nand U13565 (N_13565,N_10121,N_11993);
or U13566 (N_13566,N_10238,N_11162);
nand U13567 (N_13567,N_12374,N_10090);
xnor U13568 (N_13568,N_11166,N_10145);
nor U13569 (N_13569,N_9421,N_10835);
and U13570 (N_13570,N_9866,N_11066);
nor U13571 (N_13571,N_9448,N_11956);
nor U13572 (N_13572,N_10802,N_11120);
xnor U13573 (N_13573,N_9985,N_10092);
xor U13574 (N_13574,N_9440,N_9891);
nand U13575 (N_13575,N_9496,N_12032);
nor U13576 (N_13576,N_11136,N_11725);
and U13577 (N_13577,N_11477,N_9886);
or U13578 (N_13578,N_10764,N_9936);
and U13579 (N_13579,N_9427,N_10440);
xnor U13580 (N_13580,N_11132,N_9553);
or U13581 (N_13581,N_12412,N_9889);
nor U13582 (N_13582,N_11204,N_12470);
and U13583 (N_13583,N_9686,N_12403);
or U13584 (N_13584,N_9451,N_12440);
xor U13585 (N_13585,N_10939,N_10051);
and U13586 (N_13586,N_9523,N_10855);
nand U13587 (N_13587,N_9567,N_10173);
or U13588 (N_13588,N_10130,N_12417);
or U13589 (N_13589,N_11636,N_11387);
nor U13590 (N_13590,N_12404,N_11736);
and U13591 (N_13591,N_9530,N_12300);
and U13592 (N_13592,N_10964,N_11865);
nor U13593 (N_13593,N_10311,N_10677);
nor U13594 (N_13594,N_12309,N_11731);
xnor U13595 (N_13595,N_11480,N_10954);
nand U13596 (N_13596,N_10935,N_9476);
and U13597 (N_13597,N_10408,N_10372);
and U13598 (N_13598,N_9493,N_9780);
xor U13599 (N_13599,N_9629,N_9968);
and U13600 (N_13600,N_12468,N_9675);
and U13601 (N_13601,N_11572,N_11416);
xor U13602 (N_13602,N_9782,N_12043);
xor U13603 (N_13603,N_11596,N_9833);
nand U13604 (N_13604,N_10552,N_11898);
or U13605 (N_13605,N_9746,N_10164);
nand U13606 (N_13606,N_12275,N_10858);
and U13607 (N_13607,N_11930,N_11790);
xor U13608 (N_13608,N_12007,N_11954);
xor U13609 (N_13609,N_11440,N_11051);
nor U13610 (N_13610,N_11950,N_10227);
and U13611 (N_13611,N_9734,N_10956);
xnor U13612 (N_13612,N_10197,N_10331);
nand U13613 (N_13613,N_9449,N_12280);
or U13614 (N_13614,N_10495,N_11420);
and U13615 (N_13615,N_10615,N_11874);
nor U13616 (N_13616,N_9430,N_10395);
or U13617 (N_13617,N_10154,N_9514);
nand U13618 (N_13618,N_12379,N_11230);
or U13619 (N_13619,N_12169,N_9516);
xor U13620 (N_13620,N_11292,N_9753);
and U13621 (N_13621,N_10693,N_10774);
xor U13622 (N_13622,N_9867,N_11776);
nand U13623 (N_13623,N_10563,N_10413);
nand U13624 (N_13624,N_10687,N_11894);
and U13625 (N_13625,N_10517,N_10501);
and U13626 (N_13626,N_10608,N_10674);
nand U13627 (N_13627,N_11843,N_9728);
nand U13628 (N_13628,N_9984,N_11458);
or U13629 (N_13629,N_11461,N_11375);
or U13630 (N_13630,N_12238,N_9747);
and U13631 (N_13631,N_11069,N_12486);
nor U13632 (N_13632,N_11333,N_11605);
nand U13633 (N_13633,N_10161,N_10824);
or U13634 (N_13634,N_10676,N_12430);
or U13635 (N_13635,N_11445,N_10763);
or U13636 (N_13636,N_10356,N_12021);
nand U13637 (N_13637,N_11310,N_10342);
nor U13638 (N_13638,N_10107,N_11370);
or U13639 (N_13639,N_12386,N_12354);
or U13640 (N_13640,N_11397,N_10921);
nand U13641 (N_13641,N_12284,N_11632);
and U13642 (N_13642,N_10181,N_9593);
and U13643 (N_13643,N_10323,N_11580);
nor U13644 (N_13644,N_10649,N_9560);
nor U13645 (N_13645,N_11104,N_11492);
and U13646 (N_13646,N_10539,N_9506);
and U13647 (N_13647,N_12111,N_9694);
or U13648 (N_13648,N_10315,N_11273);
and U13649 (N_13649,N_10515,N_11438);
nor U13650 (N_13650,N_10658,N_10974);
nor U13651 (N_13651,N_10032,N_12292);
nor U13652 (N_13652,N_10588,N_12005);
nand U13653 (N_13653,N_10388,N_12380);
nor U13654 (N_13654,N_10091,N_9778);
or U13655 (N_13655,N_10943,N_11841);
nand U13656 (N_13656,N_12112,N_9443);
and U13657 (N_13657,N_11509,N_10781);
and U13658 (N_13658,N_10274,N_10576);
or U13659 (N_13659,N_11020,N_11165);
and U13660 (N_13660,N_12231,N_12352);
nor U13661 (N_13661,N_10337,N_9657);
or U13662 (N_13662,N_11947,N_11300);
xor U13663 (N_13663,N_10872,N_10291);
xor U13664 (N_13664,N_12138,N_10814);
xor U13665 (N_13665,N_10963,N_10851);
nand U13666 (N_13666,N_10352,N_12376);
or U13667 (N_13667,N_12341,N_10321);
or U13668 (N_13668,N_12463,N_9527);
nor U13669 (N_13669,N_12077,N_9967);
xnor U13670 (N_13670,N_11541,N_10207);
nor U13671 (N_13671,N_11342,N_11880);
nand U13672 (N_13672,N_9804,N_10007);
xor U13673 (N_13673,N_10585,N_11463);
or U13674 (N_13674,N_11024,N_11374);
and U13675 (N_13675,N_10067,N_12297);
or U13676 (N_13676,N_10191,N_9583);
and U13677 (N_13677,N_9624,N_11971);
xor U13678 (N_13678,N_11146,N_9428);
xor U13679 (N_13679,N_9646,N_10945);
xor U13680 (N_13680,N_11446,N_12167);
nand U13681 (N_13681,N_10187,N_12042);
or U13682 (N_13682,N_12365,N_11519);
nor U13683 (N_13683,N_10811,N_11100);
nor U13684 (N_13684,N_10209,N_11627);
nor U13685 (N_13685,N_11280,N_11641);
nor U13686 (N_13686,N_11766,N_9616);
or U13687 (N_13687,N_10969,N_9834);
xnor U13688 (N_13688,N_12056,N_11774);
nor U13689 (N_13689,N_11763,N_9442);
nand U13690 (N_13690,N_11789,N_9947);
and U13691 (N_13691,N_11143,N_9796);
or U13692 (N_13692,N_10791,N_11053);
nand U13693 (N_13693,N_10952,N_11683);
and U13694 (N_13694,N_10267,N_12209);
and U13695 (N_13695,N_11645,N_10594);
or U13696 (N_13696,N_11032,N_10968);
and U13697 (N_13697,N_10035,N_9762);
nand U13698 (N_13698,N_11040,N_12361);
xor U13699 (N_13699,N_10755,N_10492);
nor U13700 (N_13700,N_11380,N_11508);
xor U13701 (N_13701,N_10365,N_11715);
and U13702 (N_13702,N_10122,N_10012);
nor U13703 (N_13703,N_9931,N_12090);
nand U13704 (N_13704,N_11872,N_11153);
xnor U13705 (N_13705,N_10141,N_11879);
or U13706 (N_13706,N_11703,N_11402);
nor U13707 (N_13707,N_10803,N_11060);
nor U13708 (N_13708,N_12351,N_9634);
xor U13709 (N_13709,N_9860,N_11514);
nand U13710 (N_13710,N_12159,N_9680);
nand U13711 (N_13711,N_12329,N_10483);
or U13712 (N_13712,N_11717,N_10296);
nand U13713 (N_13713,N_10163,N_9790);
nand U13714 (N_13714,N_11170,N_10918);
or U13715 (N_13715,N_10162,N_11593);
nor U13716 (N_13716,N_9596,N_12148);
or U13717 (N_13717,N_11250,N_9990);
or U13718 (N_13718,N_11316,N_11299);
xor U13719 (N_13719,N_10776,N_11816);
nand U13720 (N_13720,N_9768,N_9490);
xnor U13721 (N_13721,N_11752,N_11429);
nor U13722 (N_13722,N_11922,N_10625);
nor U13723 (N_13723,N_10683,N_10339);
xnor U13724 (N_13724,N_10213,N_12358);
nand U13725 (N_13725,N_9939,N_11381);
or U13726 (N_13726,N_10808,N_9737);
xnor U13727 (N_13727,N_10189,N_9376);
nand U13728 (N_13728,N_11554,N_9977);
xnor U13729 (N_13729,N_10735,N_9396);
or U13730 (N_13730,N_10398,N_11285);
or U13731 (N_13731,N_10111,N_12114);
nand U13732 (N_13732,N_12217,N_12373);
xor U13733 (N_13733,N_10596,N_9953);
nor U13734 (N_13734,N_11773,N_9398);
nor U13735 (N_13735,N_10147,N_9406);
or U13736 (N_13736,N_11556,N_11145);
or U13737 (N_13737,N_11887,N_9845);
nand U13738 (N_13738,N_9929,N_11377);
nand U13739 (N_13739,N_11882,N_10379);
xor U13740 (N_13740,N_12407,N_11853);
nor U13741 (N_13741,N_11392,N_12313);
nand U13742 (N_13742,N_11221,N_9413);
or U13743 (N_13743,N_10031,N_11681);
xor U13744 (N_13744,N_9755,N_9601);
nor U13745 (N_13745,N_10516,N_12084);
or U13746 (N_13746,N_11085,N_10132);
nor U13747 (N_13747,N_11732,N_9828);
xnor U13748 (N_13748,N_10888,N_11502);
xor U13749 (N_13749,N_10580,N_10218);
nor U13750 (N_13750,N_12242,N_11936);
and U13751 (N_13751,N_12349,N_11856);
nand U13752 (N_13752,N_11761,N_12481);
nand U13753 (N_13753,N_10277,N_9611);
xor U13754 (N_13754,N_11371,N_10472);
nor U13755 (N_13755,N_11987,N_9973);
nor U13756 (N_13756,N_11849,N_9666);
xor U13757 (N_13757,N_9435,N_11464);
nand U13758 (N_13758,N_11755,N_10135);
or U13759 (N_13759,N_12018,N_10386);
nand U13760 (N_13760,N_9902,N_10152);
and U13761 (N_13761,N_10409,N_10663);
nor U13762 (N_13762,N_12474,N_11325);
xnor U13763 (N_13763,N_9650,N_10805);
or U13764 (N_13764,N_9767,N_10151);
nor U13765 (N_13765,N_11621,N_11030);
nor U13766 (N_13766,N_12106,N_10722);
nor U13767 (N_13767,N_11453,N_10228);
or U13768 (N_13768,N_10745,N_12466);
nor U13769 (N_13769,N_11332,N_9972);
and U13770 (N_13770,N_11778,N_10793);
xnor U13771 (N_13771,N_11712,N_11362);
xor U13772 (N_13772,N_9508,N_11151);
nor U13773 (N_13773,N_10634,N_11276);
or U13774 (N_13774,N_9605,N_10895);
or U13775 (N_13775,N_11542,N_11097);
or U13776 (N_13776,N_10361,N_9488);
nand U13777 (N_13777,N_10621,N_11895);
or U13778 (N_13778,N_11738,N_11837);
and U13779 (N_13779,N_12449,N_11098);
or U13780 (N_13780,N_9864,N_12154);
and U13781 (N_13781,N_12241,N_11229);
nand U13782 (N_13782,N_11311,N_11155);
nor U13783 (N_13783,N_9869,N_9963);
nand U13784 (N_13784,N_9729,N_9805);
or U13785 (N_13785,N_10496,N_11669);
xor U13786 (N_13786,N_9935,N_10422);
or U13787 (N_13787,N_9626,N_11961);
xnor U13788 (N_13788,N_12206,N_10553);
nor U13789 (N_13789,N_10482,N_12183);
and U13790 (N_13790,N_10762,N_9717);
or U13791 (N_13791,N_10792,N_11953);
nand U13792 (N_13792,N_12194,N_9422);
nand U13793 (N_13793,N_11525,N_10476);
xor U13794 (N_13794,N_10170,N_10967);
nor U13795 (N_13795,N_10545,N_9854);
nor U13796 (N_13796,N_10520,N_9981);
nor U13797 (N_13797,N_10534,N_10225);
and U13798 (N_13798,N_10009,N_10561);
nand U13799 (N_13799,N_11334,N_11451);
nand U13800 (N_13800,N_11119,N_12326);
nand U13801 (N_13801,N_10991,N_9829);
or U13802 (N_13802,N_12453,N_11038);
nor U13803 (N_13803,N_9548,N_10511);
and U13804 (N_13804,N_12053,N_12371);
nand U13805 (N_13805,N_12158,N_11970);
nor U13806 (N_13806,N_11618,N_11269);
or U13807 (N_13807,N_10844,N_9395);
and U13808 (N_13808,N_12270,N_12025);
and U13809 (N_13809,N_11462,N_9466);
xnor U13810 (N_13810,N_10428,N_11410);
or U13811 (N_13811,N_9551,N_10836);
xor U13812 (N_13812,N_12152,N_11130);
xor U13813 (N_13813,N_10523,N_9575);
and U13814 (N_13814,N_9450,N_12457);
xor U13815 (N_13815,N_9417,N_10404);
nand U13816 (N_13816,N_11608,N_10726);
nand U13817 (N_13817,N_12396,N_11106);
nand U13818 (N_13818,N_11628,N_10827);
nor U13819 (N_13819,N_12003,N_10536);
nor U13820 (N_13820,N_11207,N_12494);
xnor U13821 (N_13821,N_11246,N_11432);
nor U13822 (N_13822,N_10370,N_9856);
or U13823 (N_13823,N_10240,N_12395);
or U13824 (N_13824,N_11771,N_11176);
nand U13825 (N_13825,N_11193,N_10470);
xnor U13826 (N_13826,N_9998,N_12083);
and U13827 (N_13827,N_9791,N_9862);
or U13828 (N_13828,N_11091,N_10870);
nor U13829 (N_13829,N_11959,N_12058);
and U13830 (N_13830,N_10820,N_10468);
nor U13831 (N_13831,N_9959,N_10094);
and U13832 (N_13832,N_10190,N_11424);
xor U13833 (N_13833,N_11570,N_9794);
and U13834 (N_13834,N_12164,N_9433);
and U13835 (N_13835,N_10312,N_10719);
xor U13836 (N_13836,N_11920,N_9425);
xor U13837 (N_13837,N_9669,N_11439);
nor U13838 (N_13838,N_12224,N_10234);
or U13839 (N_13839,N_11195,N_10405);
xnor U13840 (N_13840,N_12343,N_11352);
or U13841 (N_13841,N_10509,N_10686);
nor U13842 (N_13842,N_9391,N_11028);
and U13843 (N_13843,N_9431,N_12262);
or U13844 (N_13844,N_10664,N_12421);
nor U13845 (N_13845,N_11967,N_9895);
and U13846 (N_13846,N_12190,N_11536);
xnor U13847 (N_13847,N_12424,N_10310);
xor U13848 (N_13848,N_12223,N_12366);
nand U13849 (N_13849,N_12411,N_10962);
and U13850 (N_13850,N_10910,N_10169);
and U13851 (N_13851,N_9707,N_9899);
or U13852 (N_13852,N_11428,N_11365);
or U13853 (N_13853,N_9668,N_9658);
nor U13854 (N_13854,N_9621,N_9799);
nor U13855 (N_13855,N_9520,N_11739);
nand U13856 (N_13856,N_9578,N_9700);
nor U13857 (N_13857,N_11927,N_10399);
or U13858 (N_13858,N_12008,N_11209);
xor U13859 (N_13859,N_11177,N_11675);
nor U13860 (N_13860,N_10632,N_11757);
nor U13861 (N_13861,N_12062,N_10720);
nand U13862 (N_13862,N_9563,N_10861);
xnor U13863 (N_13863,N_9873,N_12233);
nor U13864 (N_13864,N_10466,N_9573);
xor U13865 (N_13865,N_10385,N_10245);
nand U13866 (N_13866,N_11630,N_11394);
nor U13867 (N_13867,N_11609,N_11345);
nor U13868 (N_13868,N_11718,N_11747);
xor U13869 (N_13869,N_12488,N_9908);
and U13870 (N_13870,N_10656,N_11023);
nor U13871 (N_13871,N_10684,N_10780);
xor U13872 (N_13872,N_12205,N_10431);
nand U13873 (N_13873,N_9776,N_11305);
nand U13874 (N_13874,N_10056,N_10256);
and U13875 (N_13875,N_11499,N_10734);
nor U13876 (N_13876,N_11599,N_11183);
xnor U13877 (N_13877,N_9638,N_12176);
nor U13878 (N_13878,N_11029,N_11008);
and U13879 (N_13879,N_10479,N_9379);
xor U13880 (N_13880,N_11677,N_11860);
nand U13881 (N_13881,N_10629,N_12348);
nor U13882 (N_13882,N_10471,N_11994);
nand U13883 (N_13883,N_9384,N_12248);
nor U13884 (N_13884,N_10282,N_10360);
or U13885 (N_13885,N_11034,N_9387);
nor U13886 (N_13886,N_12263,N_12325);
nor U13887 (N_13887,N_10624,N_9787);
xnor U13888 (N_13888,N_11698,N_11857);
xor U13889 (N_13889,N_11408,N_10017);
nand U13890 (N_13890,N_12047,N_10830);
and U13891 (N_13891,N_11701,N_10641);
xor U13892 (N_13892,N_11583,N_11892);
or U13893 (N_13893,N_10402,N_12015);
xnor U13894 (N_13894,N_10309,N_11893);
xnor U13895 (N_13895,N_10513,N_10584);
nor U13896 (N_13896,N_11088,N_11682);
nor U13897 (N_13897,N_9903,N_10562);
nor U13898 (N_13898,N_12146,N_10074);
and U13899 (N_13899,N_11056,N_10075);
nor U13900 (N_13900,N_9726,N_9682);
or U13901 (N_13901,N_11254,N_12170);
or U13902 (N_13902,N_9894,N_9627);
nand U13903 (N_13903,N_11676,N_11940);
xnor U13904 (N_13904,N_11302,N_10795);
nor U13905 (N_13905,N_10572,N_12165);
and U13906 (N_13906,N_12445,N_10589);
xor U13907 (N_13907,N_11483,N_12204);
nor U13908 (N_13908,N_11650,N_11102);
xor U13909 (N_13909,N_9950,N_9847);
xnor U13910 (N_13910,N_11078,N_10582);
nand U13911 (N_13911,N_11430,N_9452);
nor U13912 (N_13912,N_11810,N_10979);
nor U13913 (N_13913,N_12130,N_9385);
xnor U13914 (N_13914,N_10434,N_12125);
or U13915 (N_13915,N_11568,N_11520);
xor U13916 (N_13916,N_10239,N_10787);
nand U13917 (N_13917,N_11981,N_9740);
nand U13918 (N_13918,N_9863,N_10987);
or U13919 (N_13919,N_12126,N_10862);
nor U13920 (N_13920,N_11515,N_12022);
nand U13921 (N_13921,N_10771,N_11017);
xor U13922 (N_13922,N_10989,N_12394);
or U13923 (N_13923,N_10670,N_11467);
nor U13924 (N_13924,N_11914,N_11526);
nor U13925 (N_13925,N_10033,N_9999);
or U13926 (N_13926,N_10444,N_12172);
nand U13927 (N_13927,N_10541,N_10252);
nand U13928 (N_13928,N_10369,N_11696);
nand U13929 (N_13929,N_11935,N_9426);
and U13930 (N_13930,N_11928,N_10390);
nand U13931 (N_13931,N_12100,N_9542);
nand U13932 (N_13932,N_10574,N_12337);
nor U13933 (N_13933,N_12055,N_9917);
xnor U13934 (N_13934,N_11154,N_9447);
nor U13935 (N_13935,N_12444,N_11122);
or U13936 (N_13936,N_10229,N_12402);
or U13937 (N_13937,N_12028,N_10940);
nand U13938 (N_13938,N_11227,N_12163);
nor U13939 (N_13939,N_10530,N_9620);
nand U13940 (N_13940,N_10923,N_11655);
and U13941 (N_13941,N_10453,N_9580);
nor U13942 (N_13942,N_11203,N_10725);
xor U13943 (N_13943,N_11521,N_11934);
xnor U13944 (N_13944,N_9546,N_10533);
and U13945 (N_13945,N_11522,N_10837);
and U13946 (N_13946,N_9375,N_11553);
and U13947 (N_13947,N_10233,N_11005);
nor U13948 (N_13948,N_10451,N_11488);
and U13949 (N_13949,N_11783,N_11740);
nor U13950 (N_13950,N_9853,N_9556);
nand U13951 (N_13951,N_12144,N_12428);
nand U13952 (N_13952,N_9695,N_12145);
nor U13953 (N_13953,N_10078,N_10936);
and U13954 (N_13954,N_10587,N_11903);
or U13955 (N_13955,N_9811,N_9597);
nand U13956 (N_13956,N_9660,N_10671);
or U13957 (N_13957,N_11700,N_9835);
or U13958 (N_13958,N_10086,N_10341);
or U13959 (N_13959,N_10854,N_12061);
and U13960 (N_13960,N_11585,N_9477);
nand U13961 (N_13961,N_12016,N_10512);
xnor U13962 (N_13962,N_9783,N_10712);
xor U13963 (N_13963,N_11045,N_10410);
xnor U13964 (N_13964,N_9713,N_11164);
nor U13965 (N_13965,N_9524,N_12461);
nand U13966 (N_13966,N_10336,N_9651);
nand U13967 (N_13967,N_12132,N_9464);
nand U13968 (N_13968,N_9978,N_11545);
xnor U13969 (N_13969,N_10328,N_10538);
nor U13970 (N_13970,N_10990,N_10696);
and U13971 (N_13971,N_10760,N_11435);
nand U13972 (N_13972,N_11883,N_9654);
xnor U13973 (N_13973,N_11350,N_11665);
or U13974 (N_13974,N_10054,N_10364);
nor U13975 (N_13975,N_11911,N_12129);
xor U13976 (N_13976,N_9812,N_12472);
nand U13977 (N_13977,N_10728,N_11126);
and U13978 (N_13978,N_11268,N_11324);
xnor U13979 (N_13979,N_10002,N_11537);
and U13980 (N_13980,N_9781,N_11004);
xnor U13981 (N_13981,N_9992,N_10098);
nor U13982 (N_13982,N_10673,N_11270);
and U13983 (N_13983,N_10682,N_10214);
nor U13984 (N_13984,N_10284,N_9910);
nor U13985 (N_13985,N_12012,N_10185);
or U13986 (N_13986,N_11962,N_11027);
xnor U13987 (N_13987,N_9871,N_11512);
and U13988 (N_13988,N_11973,N_11984);
or U13989 (N_13989,N_9509,N_11988);
or U13990 (N_13990,N_10118,N_10768);
nand U13991 (N_13991,N_9920,N_9441);
or U13992 (N_13992,N_9771,N_9502);
or U13993 (N_13993,N_11315,N_11921);
and U13994 (N_13994,N_10250,N_11601);
or U13995 (N_13995,N_11697,N_9557);
or U13996 (N_13996,N_11610,N_10114);
xor U13997 (N_13997,N_11080,N_10503);
nand U13998 (N_13998,N_11109,N_10297);
and U13999 (N_13999,N_10976,N_10251);
nand U14000 (N_14000,N_11468,N_11399);
xor U14001 (N_14001,N_11341,N_10411);
nor U14002 (N_14002,N_9775,N_11283);
and U14003 (N_14003,N_9741,N_9503);
and U14004 (N_14004,N_10420,N_12189);
xnor U14005 (N_14005,N_11990,N_11413);
xnor U14006 (N_14006,N_11784,N_10915);
and U14007 (N_14007,N_11469,N_11692);
or U14008 (N_14008,N_10876,N_9879);
and U14009 (N_14009,N_10558,N_9975);
nand U14010 (N_14010,N_9784,N_11506);
or U14011 (N_14011,N_10433,N_11809);
nand U14012 (N_14012,N_12094,N_10554);
nor U14013 (N_14013,N_11009,N_10397);
and U14014 (N_14014,N_11173,N_11998);
and U14015 (N_14015,N_9457,N_11063);
xor U14016 (N_14016,N_9691,N_9444);
and U14017 (N_14017,N_11174,N_10198);
nor U14018 (N_14018,N_11667,N_11662);
xnor U14019 (N_14019,N_10548,N_10662);
and U14020 (N_14020,N_10349,N_9800);
xor U14021 (N_14021,N_10268,N_9633);
nor U14022 (N_14022,N_11666,N_10241);
or U14023 (N_14023,N_12120,N_10465);
and U14024 (N_14024,N_10653,N_11237);
nor U14025 (N_14025,N_11907,N_11291);
and U14026 (N_14026,N_10222,N_11828);
xnor U14027 (N_14027,N_11533,N_11616);
or U14028 (N_14028,N_12353,N_12344);
or U14029 (N_14029,N_10806,N_9946);
xor U14030 (N_14030,N_10286,N_9870);
and U14031 (N_14031,N_10709,N_10294);
or U14032 (N_14032,N_12002,N_12181);
xnor U14033 (N_14033,N_9470,N_11517);
or U14034 (N_14034,N_11639,N_10071);
nand U14035 (N_14035,N_12429,N_10977);
or U14036 (N_14036,N_11248,N_11781);
or U14037 (N_14037,N_9511,N_11084);
or U14038 (N_14038,N_9467,N_9699);
and U14039 (N_14039,N_10329,N_11490);
xor U14040 (N_14040,N_11744,N_11425);
nor U14041 (N_14041,N_10313,N_11624);
nor U14042 (N_14042,N_11986,N_11179);
nand U14043 (N_14043,N_9525,N_10210);
and U14044 (N_14044,N_12492,N_11845);
nand U14045 (N_14045,N_10640,N_9416);
nand U14046 (N_14046,N_10412,N_11995);
or U14047 (N_14047,N_9453,N_10866);
or U14048 (N_14048,N_12063,N_10128);
and U14049 (N_14049,N_12065,N_9501);
nand U14050 (N_14050,N_10881,N_12105);
and U14051 (N_14051,N_11561,N_11417);
nand U14052 (N_14052,N_10826,N_12178);
and U14053 (N_14053,N_11190,N_9608);
and U14054 (N_14054,N_10891,N_10863);
nand U14055 (N_14055,N_11290,N_10995);
nand U14056 (N_14056,N_10374,N_12027);
nor U14057 (N_14057,N_11391,N_10581);
nor U14058 (N_14058,N_12098,N_10016);
xnor U14059 (N_14059,N_10773,N_10909);
nor U14060 (N_14060,N_10271,N_10577);
xnor U14061 (N_14061,N_11491,N_12071);
or U14062 (N_14062,N_10246,N_10754);
nor U14063 (N_14063,N_11861,N_12289);
or U14064 (N_14064,N_10644,N_11949);
and U14065 (N_14065,N_10445,N_9437);
and U14066 (N_14066,N_12368,N_9508);
or U14067 (N_14067,N_10666,N_12139);
and U14068 (N_14068,N_10044,N_11948);
or U14069 (N_14069,N_11234,N_10711);
nor U14070 (N_14070,N_9513,N_9786);
nor U14071 (N_14071,N_10366,N_12144);
and U14072 (N_14072,N_10215,N_9870);
or U14073 (N_14073,N_12291,N_12432);
nand U14074 (N_14074,N_10708,N_9613);
nor U14075 (N_14075,N_10910,N_10188);
or U14076 (N_14076,N_12151,N_10557);
or U14077 (N_14077,N_11802,N_11886);
xnor U14078 (N_14078,N_12129,N_10574);
nand U14079 (N_14079,N_10880,N_9788);
nor U14080 (N_14080,N_12295,N_11727);
and U14081 (N_14081,N_10405,N_11958);
xnor U14082 (N_14082,N_12369,N_11376);
or U14083 (N_14083,N_9433,N_11827);
nand U14084 (N_14084,N_10768,N_12280);
nand U14085 (N_14085,N_11202,N_9811);
and U14086 (N_14086,N_12242,N_12025);
nor U14087 (N_14087,N_11894,N_10162);
nor U14088 (N_14088,N_10081,N_11888);
nor U14089 (N_14089,N_10956,N_12155);
nand U14090 (N_14090,N_12409,N_10952);
nand U14091 (N_14091,N_9854,N_10357);
or U14092 (N_14092,N_9641,N_11944);
nand U14093 (N_14093,N_9996,N_11771);
nor U14094 (N_14094,N_12418,N_10576);
xor U14095 (N_14095,N_10115,N_10151);
and U14096 (N_14096,N_10210,N_10740);
and U14097 (N_14097,N_11155,N_10377);
nand U14098 (N_14098,N_12304,N_11116);
or U14099 (N_14099,N_11806,N_12388);
and U14100 (N_14100,N_11961,N_12034);
nand U14101 (N_14101,N_11155,N_9693);
and U14102 (N_14102,N_11156,N_12421);
nand U14103 (N_14103,N_10424,N_10697);
nand U14104 (N_14104,N_12329,N_11375);
nor U14105 (N_14105,N_10353,N_10058);
nand U14106 (N_14106,N_10068,N_10157);
xnor U14107 (N_14107,N_9562,N_10803);
or U14108 (N_14108,N_11651,N_9517);
nand U14109 (N_14109,N_11696,N_9549);
nor U14110 (N_14110,N_11710,N_10291);
nand U14111 (N_14111,N_9866,N_12498);
and U14112 (N_14112,N_10418,N_11251);
xnor U14113 (N_14113,N_10897,N_12139);
or U14114 (N_14114,N_9532,N_11506);
and U14115 (N_14115,N_11665,N_9402);
or U14116 (N_14116,N_11154,N_11753);
nor U14117 (N_14117,N_10095,N_10505);
or U14118 (N_14118,N_9808,N_12241);
and U14119 (N_14119,N_11256,N_12184);
nor U14120 (N_14120,N_9718,N_9879);
nor U14121 (N_14121,N_9689,N_10495);
or U14122 (N_14122,N_9832,N_9526);
nor U14123 (N_14123,N_11017,N_10875);
xnor U14124 (N_14124,N_10962,N_11776);
nand U14125 (N_14125,N_9882,N_10529);
nand U14126 (N_14126,N_12002,N_11506);
nor U14127 (N_14127,N_10898,N_9713);
nor U14128 (N_14128,N_10358,N_9790);
or U14129 (N_14129,N_9556,N_11639);
and U14130 (N_14130,N_11500,N_9752);
and U14131 (N_14131,N_10446,N_11479);
nor U14132 (N_14132,N_11046,N_11463);
nor U14133 (N_14133,N_12287,N_12434);
xor U14134 (N_14134,N_11790,N_11435);
and U14135 (N_14135,N_11438,N_9608);
xor U14136 (N_14136,N_11810,N_11965);
or U14137 (N_14137,N_11586,N_9854);
nor U14138 (N_14138,N_12259,N_10370);
nand U14139 (N_14139,N_11324,N_10201);
and U14140 (N_14140,N_10889,N_11193);
nor U14141 (N_14141,N_10460,N_12160);
or U14142 (N_14142,N_12249,N_12074);
xor U14143 (N_14143,N_11888,N_10610);
nand U14144 (N_14144,N_11602,N_10363);
nor U14145 (N_14145,N_9427,N_10834);
nor U14146 (N_14146,N_10798,N_9924);
xnor U14147 (N_14147,N_12140,N_10895);
and U14148 (N_14148,N_10777,N_11618);
or U14149 (N_14149,N_12216,N_11999);
nand U14150 (N_14150,N_10542,N_12242);
and U14151 (N_14151,N_9448,N_9737);
nor U14152 (N_14152,N_9655,N_12052);
nor U14153 (N_14153,N_11799,N_10553);
and U14154 (N_14154,N_9937,N_9965);
and U14155 (N_14155,N_12237,N_12197);
xor U14156 (N_14156,N_11801,N_10741);
and U14157 (N_14157,N_10986,N_12137);
xor U14158 (N_14158,N_12198,N_12499);
nand U14159 (N_14159,N_11644,N_12340);
nor U14160 (N_14160,N_10413,N_10878);
and U14161 (N_14161,N_10513,N_11028);
nor U14162 (N_14162,N_11952,N_10836);
or U14163 (N_14163,N_12012,N_10339);
nand U14164 (N_14164,N_12319,N_9527);
nor U14165 (N_14165,N_11858,N_10031);
or U14166 (N_14166,N_11065,N_11050);
or U14167 (N_14167,N_9542,N_11246);
xnor U14168 (N_14168,N_10160,N_10467);
or U14169 (N_14169,N_11889,N_12136);
xor U14170 (N_14170,N_10627,N_11290);
nand U14171 (N_14171,N_11203,N_10062);
nor U14172 (N_14172,N_9528,N_12291);
and U14173 (N_14173,N_10964,N_10912);
and U14174 (N_14174,N_9381,N_10455);
or U14175 (N_14175,N_11538,N_10276);
nor U14176 (N_14176,N_11027,N_11057);
nand U14177 (N_14177,N_11747,N_10144);
xnor U14178 (N_14178,N_10370,N_9585);
or U14179 (N_14179,N_10452,N_10167);
nand U14180 (N_14180,N_9917,N_11311);
and U14181 (N_14181,N_10690,N_10267);
xnor U14182 (N_14182,N_10538,N_11247);
and U14183 (N_14183,N_9453,N_10514);
nand U14184 (N_14184,N_9499,N_10449);
or U14185 (N_14185,N_10813,N_10795);
xor U14186 (N_14186,N_11854,N_11370);
nor U14187 (N_14187,N_12285,N_12249);
nor U14188 (N_14188,N_9635,N_12479);
and U14189 (N_14189,N_10723,N_11448);
nor U14190 (N_14190,N_12244,N_11345);
nor U14191 (N_14191,N_10801,N_10555);
nor U14192 (N_14192,N_11340,N_11531);
and U14193 (N_14193,N_9451,N_10100);
and U14194 (N_14194,N_11499,N_11838);
nand U14195 (N_14195,N_11182,N_10539);
and U14196 (N_14196,N_10597,N_11264);
nor U14197 (N_14197,N_11748,N_10333);
or U14198 (N_14198,N_9863,N_10747);
or U14199 (N_14199,N_10070,N_9704);
nor U14200 (N_14200,N_11203,N_10624);
nand U14201 (N_14201,N_9426,N_9977);
nor U14202 (N_14202,N_11277,N_9776);
xor U14203 (N_14203,N_12477,N_10271);
xnor U14204 (N_14204,N_10494,N_10417);
xnor U14205 (N_14205,N_10255,N_11974);
and U14206 (N_14206,N_11783,N_10637);
or U14207 (N_14207,N_11539,N_11921);
and U14208 (N_14208,N_9771,N_10964);
nor U14209 (N_14209,N_10340,N_11019);
nor U14210 (N_14210,N_11535,N_11215);
or U14211 (N_14211,N_12105,N_9576);
and U14212 (N_14212,N_10745,N_9477);
and U14213 (N_14213,N_10333,N_12389);
nand U14214 (N_14214,N_12375,N_11629);
nor U14215 (N_14215,N_12100,N_10253);
nand U14216 (N_14216,N_10721,N_10741);
or U14217 (N_14217,N_12007,N_12184);
nor U14218 (N_14218,N_11021,N_10820);
xnor U14219 (N_14219,N_9550,N_12263);
or U14220 (N_14220,N_10908,N_11899);
nand U14221 (N_14221,N_10564,N_9736);
xnor U14222 (N_14222,N_9914,N_11262);
nor U14223 (N_14223,N_11349,N_11272);
nor U14224 (N_14224,N_11931,N_11635);
xnor U14225 (N_14225,N_11897,N_10849);
xor U14226 (N_14226,N_11319,N_9476);
nor U14227 (N_14227,N_12198,N_10295);
nor U14228 (N_14228,N_11282,N_9577);
and U14229 (N_14229,N_11622,N_9792);
nor U14230 (N_14230,N_11749,N_10515);
and U14231 (N_14231,N_10193,N_12376);
nand U14232 (N_14232,N_11761,N_12119);
and U14233 (N_14233,N_11703,N_10893);
nor U14234 (N_14234,N_11595,N_10665);
nand U14235 (N_14235,N_10967,N_11068);
nand U14236 (N_14236,N_10954,N_9449);
nor U14237 (N_14237,N_9443,N_10964);
nand U14238 (N_14238,N_10926,N_10231);
xnor U14239 (N_14239,N_12053,N_9743);
or U14240 (N_14240,N_11340,N_10937);
or U14241 (N_14241,N_9809,N_12241);
nor U14242 (N_14242,N_9964,N_11589);
and U14243 (N_14243,N_9787,N_10176);
xnor U14244 (N_14244,N_10746,N_11477);
nand U14245 (N_14245,N_10711,N_11527);
xor U14246 (N_14246,N_10157,N_12020);
nor U14247 (N_14247,N_10303,N_10957);
or U14248 (N_14248,N_12394,N_11331);
xnor U14249 (N_14249,N_12164,N_11341);
xnor U14250 (N_14250,N_11415,N_12199);
nor U14251 (N_14251,N_11469,N_11308);
nor U14252 (N_14252,N_11848,N_11282);
nand U14253 (N_14253,N_12361,N_11431);
or U14254 (N_14254,N_10294,N_10318);
xor U14255 (N_14255,N_9436,N_9926);
nand U14256 (N_14256,N_11770,N_10024);
or U14257 (N_14257,N_10128,N_9676);
nor U14258 (N_14258,N_11190,N_11182);
xnor U14259 (N_14259,N_10242,N_12295);
nand U14260 (N_14260,N_11598,N_10732);
and U14261 (N_14261,N_12089,N_11105);
and U14262 (N_14262,N_11272,N_9434);
xor U14263 (N_14263,N_11255,N_11567);
and U14264 (N_14264,N_9461,N_10188);
nand U14265 (N_14265,N_11968,N_9492);
xnor U14266 (N_14266,N_9693,N_10127);
and U14267 (N_14267,N_10752,N_11736);
or U14268 (N_14268,N_9538,N_11387);
nor U14269 (N_14269,N_11622,N_11877);
or U14270 (N_14270,N_11500,N_12111);
or U14271 (N_14271,N_11619,N_11035);
nor U14272 (N_14272,N_10132,N_10478);
and U14273 (N_14273,N_10363,N_9740);
xnor U14274 (N_14274,N_11496,N_12108);
nand U14275 (N_14275,N_10281,N_10833);
or U14276 (N_14276,N_12177,N_10278);
nor U14277 (N_14277,N_11259,N_9827);
and U14278 (N_14278,N_12462,N_11288);
and U14279 (N_14279,N_12299,N_12182);
and U14280 (N_14280,N_11092,N_9685);
or U14281 (N_14281,N_12039,N_10647);
nand U14282 (N_14282,N_12146,N_12205);
and U14283 (N_14283,N_10546,N_10990);
xor U14284 (N_14284,N_10829,N_11884);
and U14285 (N_14285,N_12323,N_9539);
nand U14286 (N_14286,N_11681,N_9990);
nand U14287 (N_14287,N_10386,N_12288);
and U14288 (N_14288,N_11036,N_11297);
nor U14289 (N_14289,N_9881,N_12309);
nand U14290 (N_14290,N_10760,N_12308);
xnor U14291 (N_14291,N_10870,N_9850);
xor U14292 (N_14292,N_11610,N_10337);
or U14293 (N_14293,N_9442,N_9867);
and U14294 (N_14294,N_9855,N_9740);
nor U14295 (N_14295,N_11158,N_11412);
or U14296 (N_14296,N_11394,N_9583);
xor U14297 (N_14297,N_9733,N_9902);
nand U14298 (N_14298,N_12154,N_10199);
or U14299 (N_14299,N_10879,N_10101);
xor U14300 (N_14300,N_9817,N_9826);
nor U14301 (N_14301,N_9696,N_11214);
and U14302 (N_14302,N_9685,N_10095);
xnor U14303 (N_14303,N_12353,N_10290);
nand U14304 (N_14304,N_11352,N_10404);
xor U14305 (N_14305,N_11198,N_12381);
nor U14306 (N_14306,N_10057,N_12287);
and U14307 (N_14307,N_9768,N_9863);
or U14308 (N_14308,N_10317,N_11096);
or U14309 (N_14309,N_12064,N_10169);
nor U14310 (N_14310,N_11670,N_11684);
nand U14311 (N_14311,N_11425,N_10065);
and U14312 (N_14312,N_11515,N_10970);
or U14313 (N_14313,N_10414,N_12089);
and U14314 (N_14314,N_10065,N_9438);
xnor U14315 (N_14315,N_12121,N_11844);
nor U14316 (N_14316,N_11325,N_9476);
and U14317 (N_14317,N_12078,N_11845);
and U14318 (N_14318,N_12029,N_11405);
nor U14319 (N_14319,N_10474,N_11443);
or U14320 (N_14320,N_9522,N_10006);
or U14321 (N_14321,N_11347,N_9567);
and U14322 (N_14322,N_9603,N_10539);
and U14323 (N_14323,N_11080,N_11886);
nand U14324 (N_14324,N_9505,N_12362);
or U14325 (N_14325,N_10023,N_12114);
or U14326 (N_14326,N_10121,N_10673);
nor U14327 (N_14327,N_10589,N_10406);
nand U14328 (N_14328,N_10211,N_12050);
xnor U14329 (N_14329,N_12398,N_11672);
xor U14330 (N_14330,N_9584,N_12431);
and U14331 (N_14331,N_11930,N_9769);
nor U14332 (N_14332,N_12490,N_9804);
xor U14333 (N_14333,N_9958,N_12433);
nor U14334 (N_14334,N_11078,N_10144);
and U14335 (N_14335,N_10087,N_12316);
xnor U14336 (N_14336,N_12065,N_12114);
nor U14337 (N_14337,N_11911,N_10737);
and U14338 (N_14338,N_9854,N_11899);
and U14339 (N_14339,N_9504,N_12018);
or U14340 (N_14340,N_11935,N_12443);
nand U14341 (N_14341,N_9750,N_11203);
xor U14342 (N_14342,N_10471,N_10535);
xor U14343 (N_14343,N_11727,N_9922);
or U14344 (N_14344,N_11909,N_9636);
nor U14345 (N_14345,N_10168,N_12299);
or U14346 (N_14346,N_12236,N_11795);
nor U14347 (N_14347,N_10045,N_11976);
or U14348 (N_14348,N_10096,N_11551);
or U14349 (N_14349,N_9612,N_9876);
or U14350 (N_14350,N_12313,N_12364);
nor U14351 (N_14351,N_9950,N_12330);
and U14352 (N_14352,N_10896,N_12241);
nand U14353 (N_14353,N_10871,N_12131);
nand U14354 (N_14354,N_11550,N_11525);
nor U14355 (N_14355,N_10824,N_11792);
or U14356 (N_14356,N_12352,N_12116);
nand U14357 (N_14357,N_11871,N_11965);
nand U14358 (N_14358,N_9408,N_12441);
and U14359 (N_14359,N_10603,N_12089);
xor U14360 (N_14360,N_10763,N_9426);
or U14361 (N_14361,N_11702,N_9572);
and U14362 (N_14362,N_10990,N_10426);
xnor U14363 (N_14363,N_10555,N_12339);
xor U14364 (N_14364,N_9907,N_11904);
nand U14365 (N_14365,N_11809,N_12195);
nand U14366 (N_14366,N_11884,N_11797);
or U14367 (N_14367,N_12059,N_12315);
xor U14368 (N_14368,N_10948,N_11676);
xor U14369 (N_14369,N_9832,N_9889);
and U14370 (N_14370,N_11106,N_11637);
nor U14371 (N_14371,N_10388,N_10613);
nand U14372 (N_14372,N_9732,N_11188);
nand U14373 (N_14373,N_10519,N_11190);
nor U14374 (N_14374,N_9873,N_11884);
or U14375 (N_14375,N_11029,N_10600);
and U14376 (N_14376,N_11487,N_11956);
xnor U14377 (N_14377,N_10477,N_10525);
xnor U14378 (N_14378,N_12497,N_10471);
or U14379 (N_14379,N_11916,N_10018);
xor U14380 (N_14380,N_11100,N_12035);
and U14381 (N_14381,N_12430,N_9378);
or U14382 (N_14382,N_10086,N_12243);
xor U14383 (N_14383,N_11326,N_11538);
nand U14384 (N_14384,N_12431,N_11919);
or U14385 (N_14385,N_11495,N_9588);
and U14386 (N_14386,N_12208,N_11648);
nand U14387 (N_14387,N_11633,N_12421);
nand U14388 (N_14388,N_9737,N_11937);
nor U14389 (N_14389,N_11016,N_10497);
and U14390 (N_14390,N_12338,N_11436);
nand U14391 (N_14391,N_12109,N_10398);
nor U14392 (N_14392,N_11416,N_10323);
and U14393 (N_14393,N_10464,N_11291);
xor U14394 (N_14394,N_11191,N_11514);
or U14395 (N_14395,N_10520,N_9835);
xor U14396 (N_14396,N_11180,N_11920);
and U14397 (N_14397,N_10550,N_11796);
or U14398 (N_14398,N_9556,N_9425);
xnor U14399 (N_14399,N_10851,N_10916);
nand U14400 (N_14400,N_11511,N_9596);
and U14401 (N_14401,N_9956,N_9629);
nand U14402 (N_14402,N_9616,N_12186);
nand U14403 (N_14403,N_10179,N_10971);
or U14404 (N_14404,N_12044,N_10868);
nand U14405 (N_14405,N_9900,N_11851);
or U14406 (N_14406,N_10359,N_12271);
xor U14407 (N_14407,N_10634,N_9674);
nand U14408 (N_14408,N_10286,N_11870);
nor U14409 (N_14409,N_9642,N_9930);
xor U14410 (N_14410,N_11317,N_10280);
nand U14411 (N_14411,N_12297,N_11646);
xor U14412 (N_14412,N_11947,N_10297);
xor U14413 (N_14413,N_11788,N_11862);
nand U14414 (N_14414,N_10571,N_9511);
or U14415 (N_14415,N_12096,N_12462);
and U14416 (N_14416,N_10606,N_10873);
nor U14417 (N_14417,N_12246,N_9982);
nor U14418 (N_14418,N_10855,N_11908);
nand U14419 (N_14419,N_12044,N_10601);
or U14420 (N_14420,N_10779,N_11257);
or U14421 (N_14421,N_9447,N_10974);
nand U14422 (N_14422,N_11564,N_11627);
and U14423 (N_14423,N_12168,N_11739);
nand U14424 (N_14424,N_11354,N_9791);
nand U14425 (N_14425,N_10671,N_12099);
xor U14426 (N_14426,N_10901,N_10903);
nand U14427 (N_14427,N_12033,N_10085);
xor U14428 (N_14428,N_9576,N_11495);
and U14429 (N_14429,N_9446,N_11254);
nor U14430 (N_14430,N_9950,N_10521);
nor U14431 (N_14431,N_10189,N_11455);
nand U14432 (N_14432,N_10359,N_11607);
nor U14433 (N_14433,N_10736,N_11483);
and U14434 (N_14434,N_11388,N_9555);
and U14435 (N_14435,N_11257,N_11026);
nand U14436 (N_14436,N_10200,N_11416);
nand U14437 (N_14437,N_9845,N_10486);
nor U14438 (N_14438,N_10752,N_10299);
and U14439 (N_14439,N_12174,N_9674);
nor U14440 (N_14440,N_9710,N_11346);
or U14441 (N_14441,N_10549,N_12099);
or U14442 (N_14442,N_9793,N_10551);
nor U14443 (N_14443,N_9706,N_12414);
or U14444 (N_14444,N_10515,N_11678);
and U14445 (N_14445,N_11429,N_10223);
nor U14446 (N_14446,N_10195,N_10741);
or U14447 (N_14447,N_12382,N_10432);
xnor U14448 (N_14448,N_10760,N_9552);
and U14449 (N_14449,N_11844,N_10496);
nand U14450 (N_14450,N_9791,N_10424);
xnor U14451 (N_14451,N_10722,N_10223);
xor U14452 (N_14452,N_10293,N_11492);
nand U14453 (N_14453,N_9874,N_11272);
xor U14454 (N_14454,N_11525,N_10704);
xnor U14455 (N_14455,N_11466,N_12448);
xnor U14456 (N_14456,N_11441,N_12221);
and U14457 (N_14457,N_10784,N_10464);
or U14458 (N_14458,N_12103,N_12318);
nand U14459 (N_14459,N_9880,N_12236);
nor U14460 (N_14460,N_11386,N_10828);
nor U14461 (N_14461,N_10903,N_11265);
xor U14462 (N_14462,N_9474,N_11952);
or U14463 (N_14463,N_12391,N_10670);
nand U14464 (N_14464,N_10472,N_9685);
nand U14465 (N_14465,N_9395,N_11292);
nand U14466 (N_14466,N_10169,N_11665);
or U14467 (N_14467,N_11379,N_9618);
nand U14468 (N_14468,N_9790,N_10824);
and U14469 (N_14469,N_9446,N_11659);
and U14470 (N_14470,N_9508,N_10674);
nand U14471 (N_14471,N_12442,N_10139);
xor U14472 (N_14472,N_10009,N_11962);
xor U14473 (N_14473,N_11707,N_9745);
and U14474 (N_14474,N_9892,N_12095);
and U14475 (N_14475,N_12254,N_12091);
nand U14476 (N_14476,N_11501,N_12031);
nand U14477 (N_14477,N_12459,N_9925);
nand U14478 (N_14478,N_11676,N_10385);
nor U14479 (N_14479,N_9448,N_11842);
or U14480 (N_14480,N_10823,N_10608);
or U14481 (N_14481,N_10741,N_10554);
nor U14482 (N_14482,N_9870,N_11608);
nand U14483 (N_14483,N_9711,N_10379);
xor U14484 (N_14484,N_10132,N_10109);
nor U14485 (N_14485,N_12023,N_10538);
xor U14486 (N_14486,N_9656,N_9579);
or U14487 (N_14487,N_11541,N_9510);
nor U14488 (N_14488,N_12025,N_10390);
xnor U14489 (N_14489,N_11919,N_11312);
nand U14490 (N_14490,N_11735,N_11797);
xnor U14491 (N_14491,N_10239,N_9403);
and U14492 (N_14492,N_12393,N_11380);
nor U14493 (N_14493,N_11941,N_9683);
and U14494 (N_14494,N_10161,N_11139);
xnor U14495 (N_14495,N_10735,N_10143);
nor U14496 (N_14496,N_10731,N_10006);
xnor U14497 (N_14497,N_11922,N_9584);
and U14498 (N_14498,N_11765,N_10204);
xnor U14499 (N_14499,N_9863,N_11909);
nor U14500 (N_14500,N_11552,N_10424);
and U14501 (N_14501,N_9944,N_11394);
nor U14502 (N_14502,N_10631,N_9490);
and U14503 (N_14503,N_12091,N_10312);
nor U14504 (N_14504,N_10954,N_11084);
nor U14505 (N_14505,N_12378,N_11054);
or U14506 (N_14506,N_11426,N_12103);
nor U14507 (N_14507,N_11843,N_11853);
and U14508 (N_14508,N_10569,N_10379);
and U14509 (N_14509,N_11949,N_11687);
nor U14510 (N_14510,N_12015,N_12390);
and U14511 (N_14511,N_9678,N_10513);
nor U14512 (N_14512,N_12269,N_10191);
nand U14513 (N_14513,N_12410,N_12114);
xnor U14514 (N_14514,N_11860,N_10616);
xnor U14515 (N_14515,N_10654,N_12285);
or U14516 (N_14516,N_12074,N_9681);
nand U14517 (N_14517,N_10473,N_11015);
xnor U14518 (N_14518,N_11602,N_10614);
xnor U14519 (N_14519,N_10035,N_12414);
or U14520 (N_14520,N_12475,N_11900);
nand U14521 (N_14521,N_9892,N_10616);
and U14522 (N_14522,N_10689,N_11685);
and U14523 (N_14523,N_10474,N_11681);
xor U14524 (N_14524,N_11973,N_10321);
xnor U14525 (N_14525,N_10620,N_12091);
nand U14526 (N_14526,N_12358,N_11817);
and U14527 (N_14527,N_12004,N_11410);
xnor U14528 (N_14528,N_10162,N_12104);
xor U14529 (N_14529,N_9739,N_10835);
or U14530 (N_14530,N_10590,N_11357);
or U14531 (N_14531,N_11676,N_9737);
xor U14532 (N_14532,N_12129,N_10894);
nand U14533 (N_14533,N_9389,N_9388);
or U14534 (N_14534,N_10982,N_10549);
and U14535 (N_14535,N_9536,N_10284);
or U14536 (N_14536,N_9528,N_9426);
nand U14537 (N_14537,N_12390,N_10398);
or U14538 (N_14538,N_9462,N_10807);
or U14539 (N_14539,N_11178,N_10382);
xnor U14540 (N_14540,N_11390,N_10062);
nand U14541 (N_14541,N_12385,N_11184);
nand U14542 (N_14542,N_12058,N_10636);
nor U14543 (N_14543,N_10316,N_9788);
xor U14544 (N_14544,N_11159,N_10279);
xnor U14545 (N_14545,N_9923,N_12349);
nand U14546 (N_14546,N_11392,N_10018);
nor U14547 (N_14547,N_10233,N_12357);
and U14548 (N_14548,N_11510,N_11134);
and U14549 (N_14549,N_12202,N_10685);
nand U14550 (N_14550,N_11561,N_12456);
nand U14551 (N_14551,N_12079,N_12299);
and U14552 (N_14552,N_11415,N_11517);
and U14553 (N_14553,N_10743,N_11810);
or U14554 (N_14554,N_9533,N_12155);
nand U14555 (N_14555,N_11505,N_10239);
nand U14556 (N_14556,N_9955,N_9845);
nand U14557 (N_14557,N_10949,N_9415);
nand U14558 (N_14558,N_10405,N_10451);
xor U14559 (N_14559,N_11273,N_12469);
or U14560 (N_14560,N_12135,N_11792);
xor U14561 (N_14561,N_9476,N_11631);
and U14562 (N_14562,N_12450,N_10867);
xnor U14563 (N_14563,N_10188,N_12272);
or U14564 (N_14564,N_10875,N_10122);
nor U14565 (N_14565,N_11686,N_11056);
xnor U14566 (N_14566,N_11086,N_12109);
xor U14567 (N_14567,N_11953,N_10594);
or U14568 (N_14568,N_10015,N_9959);
or U14569 (N_14569,N_10153,N_11867);
nand U14570 (N_14570,N_12173,N_11123);
or U14571 (N_14571,N_10729,N_10388);
and U14572 (N_14572,N_9673,N_11815);
and U14573 (N_14573,N_11357,N_10900);
nand U14574 (N_14574,N_11122,N_11764);
or U14575 (N_14575,N_11396,N_11094);
or U14576 (N_14576,N_10063,N_11776);
xnor U14577 (N_14577,N_9517,N_11921);
or U14578 (N_14578,N_11255,N_12495);
xnor U14579 (N_14579,N_11233,N_11853);
or U14580 (N_14580,N_10805,N_9970);
and U14581 (N_14581,N_11839,N_10760);
and U14582 (N_14582,N_11795,N_12109);
or U14583 (N_14583,N_9612,N_11106);
and U14584 (N_14584,N_9999,N_9865);
and U14585 (N_14585,N_12165,N_9928);
or U14586 (N_14586,N_11279,N_12219);
xor U14587 (N_14587,N_12344,N_10580);
and U14588 (N_14588,N_9968,N_12393);
nand U14589 (N_14589,N_10112,N_10176);
nor U14590 (N_14590,N_11508,N_12266);
and U14591 (N_14591,N_10519,N_10333);
nor U14592 (N_14592,N_12282,N_10738);
or U14593 (N_14593,N_11296,N_11392);
nor U14594 (N_14594,N_12186,N_10575);
xor U14595 (N_14595,N_10716,N_12380);
or U14596 (N_14596,N_11644,N_9622);
nor U14597 (N_14597,N_11666,N_11051);
or U14598 (N_14598,N_12475,N_11887);
or U14599 (N_14599,N_12314,N_11782);
nand U14600 (N_14600,N_12250,N_10485);
nand U14601 (N_14601,N_10693,N_9918);
or U14602 (N_14602,N_12186,N_11258);
xnor U14603 (N_14603,N_10636,N_9622);
nor U14604 (N_14604,N_11136,N_9689);
or U14605 (N_14605,N_10796,N_11902);
and U14606 (N_14606,N_11137,N_11047);
nor U14607 (N_14607,N_11177,N_10818);
nor U14608 (N_14608,N_10051,N_9828);
and U14609 (N_14609,N_11442,N_12385);
and U14610 (N_14610,N_10230,N_11952);
or U14611 (N_14611,N_12123,N_11657);
or U14612 (N_14612,N_12472,N_12394);
nor U14613 (N_14613,N_10298,N_11630);
nand U14614 (N_14614,N_10026,N_9823);
xor U14615 (N_14615,N_9956,N_10285);
or U14616 (N_14616,N_12350,N_10510);
or U14617 (N_14617,N_12243,N_11767);
nor U14618 (N_14618,N_11806,N_10243);
or U14619 (N_14619,N_10568,N_12469);
xor U14620 (N_14620,N_11047,N_9579);
and U14621 (N_14621,N_12279,N_11291);
and U14622 (N_14622,N_11366,N_10234);
nand U14623 (N_14623,N_9470,N_9940);
or U14624 (N_14624,N_9877,N_10644);
or U14625 (N_14625,N_9401,N_11527);
nor U14626 (N_14626,N_11414,N_12410);
and U14627 (N_14627,N_12240,N_12307);
or U14628 (N_14628,N_10361,N_9455);
nand U14629 (N_14629,N_12001,N_11079);
nand U14630 (N_14630,N_10472,N_12024);
xnor U14631 (N_14631,N_12162,N_10642);
nor U14632 (N_14632,N_10980,N_11649);
or U14633 (N_14633,N_11978,N_9481);
and U14634 (N_14634,N_11534,N_10736);
xnor U14635 (N_14635,N_10638,N_9847);
and U14636 (N_14636,N_11399,N_9711);
nand U14637 (N_14637,N_9596,N_9934);
nand U14638 (N_14638,N_9668,N_9423);
nor U14639 (N_14639,N_11723,N_11660);
or U14640 (N_14640,N_11583,N_9487);
nor U14641 (N_14641,N_11612,N_10262);
and U14642 (N_14642,N_10902,N_12179);
nor U14643 (N_14643,N_11988,N_10293);
and U14644 (N_14644,N_10529,N_9431);
and U14645 (N_14645,N_12370,N_9834);
nor U14646 (N_14646,N_10395,N_10731);
and U14647 (N_14647,N_9390,N_12481);
nand U14648 (N_14648,N_9502,N_9652);
nand U14649 (N_14649,N_9402,N_11530);
nor U14650 (N_14650,N_12409,N_10648);
or U14651 (N_14651,N_11399,N_11001);
nor U14652 (N_14652,N_12324,N_10311);
xnor U14653 (N_14653,N_11083,N_10775);
nand U14654 (N_14654,N_10826,N_10288);
nor U14655 (N_14655,N_10103,N_10297);
nand U14656 (N_14656,N_11671,N_10789);
nor U14657 (N_14657,N_10413,N_11068);
nor U14658 (N_14658,N_10277,N_11543);
xnor U14659 (N_14659,N_10350,N_12494);
or U14660 (N_14660,N_11707,N_10608);
and U14661 (N_14661,N_10913,N_12196);
xor U14662 (N_14662,N_10311,N_9645);
nand U14663 (N_14663,N_10210,N_10762);
and U14664 (N_14664,N_9501,N_10241);
xnor U14665 (N_14665,N_9434,N_10144);
and U14666 (N_14666,N_11371,N_11908);
xnor U14667 (N_14667,N_11878,N_12388);
or U14668 (N_14668,N_11357,N_9856);
and U14669 (N_14669,N_9773,N_10422);
xor U14670 (N_14670,N_11807,N_11201);
and U14671 (N_14671,N_10236,N_10218);
or U14672 (N_14672,N_10573,N_10587);
nor U14673 (N_14673,N_11631,N_10425);
or U14674 (N_14674,N_11775,N_11089);
xnor U14675 (N_14675,N_9925,N_9482);
and U14676 (N_14676,N_11804,N_9771);
or U14677 (N_14677,N_10333,N_11239);
or U14678 (N_14678,N_9505,N_10506);
xor U14679 (N_14679,N_11743,N_11234);
xnor U14680 (N_14680,N_10773,N_10431);
and U14681 (N_14681,N_10058,N_10431);
or U14682 (N_14682,N_9500,N_11522);
and U14683 (N_14683,N_11707,N_11208);
xor U14684 (N_14684,N_11173,N_12495);
or U14685 (N_14685,N_10673,N_10853);
or U14686 (N_14686,N_12153,N_12315);
xor U14687 (N_14687,N_9802,N_11293);
xor U14688 (N_14688,N_9968,N_9828);
nor U14689 (N_14689,N_10798,N_10093);
nor U14690 (N_14690,N_9776,N_10841);
xnor U14691 (N_14691,N_11421,N_10122);
nor U14692 (N_14692,N_12245,N_9614);
xor U14693 (N_14693,N_9987,N_11004);
xnor U14694 (N_14694,N_11588,N_10281);
or U14695 (N_14695,N_10804,N_12281);
xor U14696 (N_14696,N_11975,N_10180);
nand U14697 (N_14697,N_10577,N_9883);
nand U14698 (N_14698,N_10163,N_11194);
nand U14699 (N_14699,N_9561,N_9535);
or U14700 (N_14700,N_11236,N_10683);
or U14701 (N_14701,N_10780,N_11267);
nand U14702 (N_14702,N_11823,N_10022);
and U14703 (N_14703,N_11731,N_9530);
and U14704 (N_14704,N_11027,N_9971);
or U14705 (N_14705,N_12049,N_10617);
xor U14706 (N_14706,N_11049,N_11038);
and U14707 (N_14707,N_9469,N_12238);
or U14708 (N_14708,N_12297,N_12298);
nor U14709 (N_14709,N_11712,N_10721);
nand U14710 (N_14710,N_9928,N_10932);
xnor U14711 (N_14711,N_10553,N_10291);
and U14712 (N_14712,N_10946,N_10242);
xnor U14713 (N_14713,N_11212,N_11152);
xor U14714 (N_14714,N_10802,N_10857);
xor U14715 (N_14715,N_10823,N_9944);
xor U14716 (N_14716,N_9921,N_9512);
nand U14717 (N_14717,N_10991,N_11494);
nand U14718 (N_14718,N_11967,N_11461);
and U14719 (N_14719,N_9673,N_10260);
xor U14720 (N_14720,N_9598,N_11831);
nor U14721 (N_14721,N_9408,N_11947);
and U14722 (N_14722,N_11808,N_9595);
nor U14723 (N_14723,N_12095,N_10007);
or U14724 (N_14724,N_10810,N_12063);
or U14725 (N_14725,N_11575,N_10461);
nand U14726 (N_14726,N_10245,N_10938);
xor U14727 (N_14727,N_11478,N_11200);
xnor U14728 (N_14728,N_10605,N_11686);
nand U14729 (N_14729,N_10008,N_11674);
or U14730 (N_14730,N_12062,N_10936);
nor U14731 (N_14731,N_11925,N_10039);
or U14732 (N_14732,N_12219,N_10738);
nand U14733 (N_14733,N_10240,N_10162);
and U14734 (N_14734,N_10948,N_9967);
nand U14735 (N_14735,N_12314,N_9687);
xor U14736 (N_14736,N_9974,N_11135);
and U14737 (N_14737,N_10340,N_10842);
or U14738 (N_14738,N_10308,N_9621);
xor U14739 (N_14739,N_10956,N_10886);
nor U14740 (N_14740,N_11994,N_11159);
nand U14741 (N_14741,N_10384,N_10837);
and U14742 (N_14742,N_11365,N_10695);
nand U14743 (N_14743,N_11366,N_10554);
xor U14744 (N_14744,N_9662,N_12028);
xor U14745 (N_14745,N_10808,N_11266);
nor U14746 (N_14746,N_12318,N_9387);
nor U14747 (N_14747,N_9953,N_11523);
or U14748 (N_14748,N_10753,N_11910);
and U14749 (N_14749,N_9574,N_10814);
nor U14750 (N_14750,N_11085,N_9786);
and U14751 (N_14751,N_10586,N_9481);
nand U14752 (N_14752,N_10600,N_12012);
and U14753 (N_14753,N_11925,N_11620);
and U14754 (N_14754,N_9457,N_12387);
nor U14755 (N_14755,N_12324,N_9803);
xnor U14756 (N_14756,N_9741,N_9556);
and U14757 (N_14757,N_9490,N_10134);
or U14758 (N_14758,N_9675,N_10322);
and U14759 (N_14759,N_10638,N_10319);
nand U14760 (N_14760,N_12321,N_10640);
nand U14761 (N_14761,N_10844,N_10270);
nand U14762 (N_14762,N_10821,N_11762);
and U14763 (N_14763,N_9641,N_10159);
xor U14764 (N_14764,N_12439,N_10838);
nor U14765 (N_14765,N_11526,N_10166);
nand U14766 (N_14766,N_12246,N_12219);
xnor U14767 (N_14767,N_11088,N_10124);
xnor U14768 (N_14768,N_12039,N_10470);
or U14769 (N_14769,N_10581,N_11235);
nor U14770 (N_14770,N_11374,N_9650);
xnor U14771 (N_14771,N_11240,N_10984);
and U14772 (N_14772,N_10219,N_10123);
or U14773 (N_14773,N_9776,N_12316);
or U14774 (N_14774,N_11069,N_10269);
xor U14775 (N_14775,N_10326,N_10630);
or U14776 (N_14776,N_9504,N_11982);
or U14777 (N_14777,N_12359,N_10508);
and U14778 (N_14778,N_12442,N_10510);
nand U14779 (N_14779,N_9934,N_10127);
and U14780 (N_14780,N_11742,N_12276);
nor U14781 (N_14781,N_11210,N_9379);
or U14782 (N_14782,N_12007,N_11310);
xnor U14783 (N_14783,N_12227,N_12078);
nand U14784 (N_14784,N_10021,N_10128);
nand U14785 (N_14785,N_11007,N_11991);
nor U14786 (N_14786,N_9887,N_9965);
nand U14787 (N_14787,N_9952,N_11596);
nand U14788 (N_14788,N_10476,N_10969);
xor U14789 (N_14789,N_12258,N_10598);
xnor U14790 (N_14790,N_10682,N_10201);
and U14791 (N_14791,N_11164,N_10672);
nand U14792 (N_14792,N_10271,N_9748);
xor U14793 (N_14793,N_9769,N_9781);
nor U14794 (N_14794,N_10925,N_10921);
and U14795 (N_14795,N_11957,N_11926);
nor U14796 (N_14796,N_11713,N_12195);
xor U14797 (N_14797,N_12242,N_10683);
nand U14798 (N_14798,N_9472,N_12362);
xor U14799 (N_14799,N_10850,N_12203);
and U14800 (N_14800,N_11982,N_10635);
nor U14801 (N_14801,N_11148,N_9586);
and U14802 (N_14802,N_11985,N_9430);
xnor U14803 (N_14803,N_11746,N_11160);
and U14804 (N_14804,N_11383,N_10113);
or U14805 (N_14805,N_9632,N_10928);
xnor U14806 (N_14806,N_10047,N_12401);
and U14807 (N_14807,N_11080,N_11705);
and U14808 (N_14808,N_11849,N_9834);
nor U14809 (N_14809,N_12192,N_9849);
and U14810 (N_14810,N_12405,N_11250);
nand U14811 (N_14811,N_9669,N_11954);
or U14812 (N_14812,N_9521,N_10511);
nor U14813 (N_14813,N_11596,N_10410);
or U14814 (N_14814,N_11720,N_10783);
nand U14815 (N_14815,N_9446,N_9601);
and U14816 (N_14816,N_11935,N_12234);
or U14817 (N_14817,N_11925,N_9820);
xor U14818 (N_14818,N_12475,N_10273);
nor U14819 (N_14819,N_12132,N_10823);
xor U14820 (N_14820,N_10652,N_11520);
and U14821 (N_14821,N_11494,N_11291);
nand U14822 (N_14822,N_10248,N_10138);
nand U14823 (N_14823,N_11805,N_10985);
nand U14824 (N_14824,N_10978,N_12154);
nand U14825 (N_14825,N_9546,N_11786);
or U14826 (N_14826,N_9819,N_11423);
or U14827 (N_14827,N_11162,N_10529);
or U14828 (N_14828,N_12116,N_12197);
nand U14829 (N_14829,N_10913,N_10492);
xnor U14830 (N_14830,N_11023,N_10379);
or U14831 (N_14831,N_9780,N_9620);
xor U14832 (N_14832,N_11590,N_9514);
and U14833 (N_14833,N_11096,N_11454);
or U14834 (N_14834,N_11396,N_9612);
nand U14835 (N_14835,N_10046,N_11569);
or U14836 (N_14836,N_10034,N_10752);
and U14837 (N_14837,N_10126,N_10161);
and U14838 (N_14838,N_11486,N_11757);
nor U14839 (N_14839,N_9931,N_9995);
xnor U14840 (N_14840,N_9818,N_11194);
nand U14841 (N_14841,N_10269,N_12277);
or U14842 (N_14842,N_9453,N_11911);
xnor U14843 (N_14843,N_10018,N_10037);
nand U14844 (N_14844,N_12270,N_11080);
xnor U14845 (N_14845,N_9478,N_11854);
or U14846 (N_14846,N_9461,N_10648);
nand U14847 (N_14847,N_9800,N_11792);
xnor U14848 (N_14848,N_11272,N_11277);
and U14849 (N_14849,N_10634,N_10841);
nand U14850 (N_14850,N_11092,N_12165);
nor U14851 (N_14851,N_11560,N_11811);
nor U14852 (N_14852,N_11979,N_11689);
and U14853 (N_14853,N_9504,N_12492);
nand U14854 (N_14854,N_9706,N_9939);
nand U14855 (N_14855,N_10225,N_11099);
xor U14856 (N_14856,N_10435,N_11744);
nand U14857 (N_14857,N_12045,N_12356);
nand U14858 (N_14858,N_12357,N_12343);
nand U14859 (N_14859,N_9664,N_11355);
nor U14860 (N_14860,N_9996,N_9832);
and U14861 (N_14861,N_10519,N_11267);
nand U14862 (N_14862,N_10707,N_9810);
nand U14863 (N_14863,N_12316,N_11002);
nor U14864 (N_14864,N_12074,N_11505);
and U14865 (N_14865,N_9821,N_9998);
nor U14866 (N_14866,N_11246,N_12145);
nor U14867 (N_14867,N_10262,N_10806);
and U14868 (N_14868,N_10429,N_11314);
nor U14869 (N_14869,N_11563,N_9491);
and U14870 (N_14870,N_11239,N_11510);
nor U14871 (N_14871,N_12087,N_10877);
and U14872 (N_14872,N_9620,N_9579);
and U14873 (N_14873,N_9761,N_10691);
nor U14874 (N_14874,N_12411,N_12104);
or U14875 (N_14875,N_11308,N_11348);
or U14876 (N_14876,N_10331,N_12385);
and U14877 (N_14877,N_11869,N_10012);
xnor U14878 (N_14878,N_10273,N_9918);
and U14879 (N_14879,N_11588,N_10809);
nand U14880 (N_14880,N_9790,N_11018);
or U14881 (N_14881,N_9557,N_9814);
or U14882 (N_14882,N_9472,N_11341);
nand U14883 (N_14883,N_10621,N_11786);
nand U14884 (N_14884,N_11016,N_10239);
nand U14885 (N_14885,N_10838,N_12257);
nand U14886 (N_14886,N_11679,N_9581);
xor U14887 (N_14887,N_12436,N_12320);
or U14888 (N_14888,N_10579,N_11997);
nor U14889 (N_14889,N_9841,N_12396);
nor U14890 (N_14890,N_10970,N_12472);
nand U14891 (N_14891,N_9415,N_11133);
and U14892 (N_14892,N_9947,N_11070);
or U14893 (N_14893,N_12384,N_10234);
nand U14894 (N_14894,N_9639,N_12263);
xor U14895 (N_14895,N_10503,N_12168);
nand U14896 (N_14896,N_12414,N_9736);
and U14897 (N_14897,N_12122,N_9712);
nand U14898 (N_14898,N_10584,N_10237);
and U14899 (N_14899,N_11169,N_9623);
nand U14900 (N_14900,N_11166,N_11606);
nor U14901 (N_14901,N_11816,N_12083);
or U14902 (N_14902,N_11746,N_9704);
and U14903 (N_14903,N_9818,N_12256);
xnor U14904 (N_14904,N_9869,N_10321);
nor U14905 (N_14905,N_9824,N_12146);
nand U14906 (N_14906,N_12164,N_11515);
nor U14907 (N_14907,N_9847,N_10789);
or U14908 (N_14908,N_10612,N_10092);
nor U14909 (N_14909,N_9523,N_12009);
nand U14910 (N_14910,N_10177,N_11558);
or U14911 (N_14911,N_11800,N_10484);
nor U14912 (N_14912,N_10097,N_11738);
nor U14913 (N_14913,N_10332,N_10317);
and U14914 (N_14914,N_12019,N_10116);
and U14915 (N_14915,N_11263,N_12148);
and U14916 (N_14916,N_10731,N_11293);
and U14917 (N_14917,N_10716,N_12426);
nand U14918 (N_14918,N_9422,N_11420);
xor U14919 (N_14919,N_10426,N_9952);
nor U14920 (N_14920,N_12260,N_10390);
nor U14921 (N_14921,N_11414,N_12412);
nor U14922 (N_14922,N_9524,N_12081);
xnor U14923 (N_14923,N_9775,N_12343);
nor U14924 (N_14924,N_12470,N_10781);
nand U14925 (N_14925,N_9861,N_11346);
xnor U14926 (N_14926,N_12116,N_11764);
and U14927 (N_14927,N_10522,N_12136);
nor U14928 (N_14928,N_9532,N_10340);
or U14929 (N_14929,N_11100,N_9538);
xor U14930 (N_14930,N_9917,N_9915);
xnor U14931 (N_14931,N_10363,N_10626);
xnor U14932 (N_14932,N_12291,N_10810);
or U14933 (N_14933,N_11518,N_10386);
xnor U14934 (N_14934,N_10194,N_10454);
xor U14935 (N_14935,N_9763,N_11186);
nor U14936 (N_14936,N_10294,N_12206);
nand U14937 (N_14937,N_9947,N_11291);
nor U14938 (N_14938,N_12239,N_11491);
nand U14939 (N_14939,N_9473,N_10277);
xnor U14940 (N_14940,N_11065,N_9882);
nand U14941 (N_14941,N_12354,N_9911);
xnor U14942 (N_14942,N_11978,N_10985);
xnor U14943 (N_14943,N_10773,N_11621);
xor U14944 (N_14944,N_12010,N_11281);
and U14945 (N_14945,N_11056,N_12129);
and U14946 (N_14946,N_11395,N_11177);
and U14947 (N_14947,N_10094,N_10090);
and U14948 (N_14948,N_12044,N_10111);
nand U14949 (N_14949,N_11380,N_9705);
and U14950 (N_14950,N_12325,N_10136);
nand U14951 (N_14951,N_9395,N_11491);
nand U14952 (N_14952,N_12198,N_11765);
and U14953 (N_14953,N_10391,N_12296);
and U14954 (N_14954,N_11994,N_11798);
nand U14955 (N_14955,N_10620,N_9695);
and U14956 (N_14956,N_12061,N_12209);
or U14957 (N_14957,N_12091,N_11947);
and U14958 (N_14958,N_10221,N_12200);
or U14959 (N_14959,N_11103,N_9696);
xor U14960 (N_14960,N_9427,N_11361);
and U14961 (N_14961,N_12344,N_12448);
and U14962 (N_14962,N_9584,N_12498);
xnor U14963 (N_14963,N_11250,N_9852);
or U14964 (N_14964,N_10730,N_11915);
nand U14965 (N_14965,N_11981,N_9505);
and U14966 (N_14966,N_10603,N_10539);
and U14967 (N_14967,N_9895,N_10243);
xnor U14968 (N_14968,N_10769,N_9806);
nor U14969 (N_14969,N_10616,N_9649);
or U14970 (N_14970,N_11993,N_11313);
and U14971 (N_14971,N_11636,N_12304);
nor U14972 (N_14972,N_10021,N_11298);
and U14973 (N_14973,N_11955,N_10316);
or U14974 (N_14974,N_9930,N_11702);
or U14975 (N_14975,N_10900,N_9419);
and U14976 (N_14976,N_9866,N_11578);
nand U14977 (N_14977,N_10208,N_10591);
nor U14978 (N_14978,N_11127,N_11595);
and U14979 (N_14979,N_11437,N_9453);
nand U14980 (N_14980,N_12273,N_9538);
nor U14981 (N_14981,N_10583,N_10578);
xor U14982 (N_14982,N_10927,N_10232);
and U14983 (N_14983,N_11756,N_9665);
and U14984 (N_14984,N_9591,N_10787);
xnor U14985 (N_14985,N_11183,N_10538);
and U14986 (N_14986,N_11196,N_11335);
nand U14987 (N_14987,N_12210,N_11904);
xor U14988 (N_14988,N_11301,N_10880);
xor U14989 (N_14989,N_9711,N_10479);
or U14990 (N_14990,N_10045,N_10795);
xor U14991 (N_14991,N_11811,N_9577);
nand U14992 (N_14992,N_9428,N_11100);
nand U14993 (N_14993,N_10662,N_12219);
or U14994 (N_14994,N_12002,N_11295);
xor U14995 (N_14995,N_11424,N_10510);
nand U14996 (N_14996,N_12053,N_11392);
and U14997 (N_14997,N_9918,N_10039);
and U14998 (N_14998,N_12316,N_11540);
nand U14999 (N_14999,N_9965,N_9520);
nand U15000 (N_15000,N_11829,N_12019);
xnor U15001 (N_15001,N_9498,N_10989);
nand U15002 (N_15002,N_10823,N_10567);
and U15003 (N_15003,N_10649,N_10011);
xnor U15004 (N_15004,N_10520,N_10471);
and U15005 (N_15005,N_12147,N_11057);
nor U15006 (N_15006,N_12333,N_11551);
xnor U15007 (N_15007,N_10081,N_10484);
xnor U15008 (N_15008,N_11613,N_11126);
nor U15009 (N_15009,N_12175,N_10466);
and U15010 (N_15010,N_9710,N_11556);
nand U15011 (N_15011,N_9784,N_12325);
xor U15012 (N_15012,N_10610,N_12044);
or U15013 (N_15013,N_12084,N_9746);
xnor U15014 (N_15014,N_9415,N_11750);
or U15015 (N_15015,N_9547,N_9483);
and U15016 (N_15016,N_9621,N_12427);
and U15017 (N_15017,N_10121,N_11781);
xnor U15018 (N_15018,N_10941,N_11251);
nand U15019 (N_15019,N_11831,N_12025);
nor U15020 (N_15020,N_10488,N_10394);
nand U15021 (N_15021,N_11757,N_9977);
or U15022 (N_15022,N_10065,N_11793);
or U15023 (N_15023,N_11721,N_10921);
nor U15024 (N_15024,N_9773,N_10672);
nand U15025 (N_15025,N_12330,N_9678);
nor U15026 (N_15026,N_11412,N_11749);
and U15027 (N_15027,N_10765,N_10545);
or U15028 (N_15028,N_11177,N_10714);
xnor U15029 (N_15029,N_11669,N_11841);
nor U15030 (N_15030,N_9519,N_10790);
xor U15031 (N_15031,N_10800,N_11884);
or U15032 (N_15032,N_10955,N_9640);
nor U15033 (N_15033,N_9537,N_10702);
nand U15034 (N_15034,N_9543,N_10315);
and U15035 (N_15035,N_12022,N_11644);
or U15036 (N_15036,N_9575,N_10735);
nor U15037 (N_15037,N_12087,N_10873);
nand U15038 (N_15038,N_11410,N_10204);
xor U15039 (N_15039,N_10595,N_9881);
and U15040 (N_15040,N_9791,N_11537);
or U15041 (N_15041,N_10567,N_11217);
or U15042 (N_15042,N_10569,N_11308);
nand U15043 (N_15043,N_12499,N_12324);
nand U15044 (N_15044,N_9453,N_12057);
nor U15045 (N_15045,N_10198,N_11733);
nor U15046 (N_15046,N_11995,N_12078);
or U15047 (N_15047,N_12244,N_11896);
or U15048 (N_15048,N_12434,N_11412);
or U15049 (N_15049,N_11130,N_11458);
or U15050 (N_15050,N_11061,N_11920);
and U15051 (N_15051,N_10478,N_10946);
nand U15052 (N_15052,N_10907,N_11649);
or U15053 (N_15053,N_11477,N_11149);
xor U15054 (N_15054,N_10597,N_12230);
nor U15055 (N_15055,N_10000,N_10808);
nor U15056 (N_15056,N_9888,N_11790);
nand U15057 (N_15057,N_12222,N_11588);
xor U15058 (N_15058,N_9756,N_9555);
or U15059 (N_15059,N_9556,N_11424);
nor U15060 (N_15060,N_9536,N_10136);
nor U15061 (N_15061,N_11770,N_11140);
and U15062 (N_15062,N_9719,N_9756);
or U15063 (N_15063,N_10968,N_11139);
nand U15064 (N_15064,N_12036,N_11120);
or U15065 (N_15065,N_10853,N_10942);
or U15066 (N_15066,N_11103,N_11839);
or U15067 (N_15067,N_12041,N_10654);
xor U15068 (N_15068,N_11432,N_9716);
nand U15069 (N_15069,N_12279,N_12431);
nor U15070 (N_15070,N_11231,N_11437);
xor U15071 (N_15071,N_10413,N_10090);
and U15072 (N_15072,N_10485,N_11801);
and U15073 (N_15073,N_9910,N_9889);
or U15074 (N_15074,N_9584,N_12009);
nor U15075 (N_15075,N_11559,N_11141);
nor U15076 (N_15076,N_12325,N_12464);
and U15077 (N_15077,N_10482,N_11445);
or U15078 (N_15078,N_10221,N_10568);
nor U15079 (N_15079,N_9429,N_10604);
or U15080 (N_15080,N_9950,N_12256);
xor U15081 (N_15081,N_10482,N_9824);
and U15082 (N_15082,N_10351,N_11047);
or U15083 (N_15083,N_9989,N_10477);
xor U15084 (N_15084,N_11287,N_11204);
xnor U15085 (N_15085,N_10217,N_10827);
nor U15086 (N_15086,N_10437,N_11030);
nor U15087 (N_15087,N_11570,N_9440);
nand U15088 (N_15088,N_10609,N_12251);
and U15089 (N_15089,N_9694,N_11341);
or U15090 (N_15090,N_12494,N_11688);
nor U15091 (N_15091,N_10351,N_11417);
or U15092 (N_15092,N_10258,N_11375);
nand U15093 (N_15093,N_12345,N_11637);
nand U15094 (N_15094,N_11872,N_11126);
nor U15095 (N_15095,N_11467,N_9755);
or U15096 (N_15096,N_10297,N_10728);
or U15097 (N_15097,N_10844,N_12312);
or U15098 (N_15098,N_9716,N_10731);
xor U15099 (N_15099,N_11981,N_11322);
or U15100 (N_15100,N_12273,N_12070);
or U15101 (N_15101,N_11356,N_9659);
and U15102 (N_15102,N_10128,N_11854);
xnor U15103 (N_15103,N_12045,N_11217);
or U15104 (N_15104,N_11957,N_12376);
nor U15105 (N_15105,N_9728,N_10012);
or U15106 (N_15106,N_12114,N_10665);
and U15107 (N_15107,N_10832,N_9718);
or U15108 (N_15108,N_9968,N_10455);
nor U15109 (N_15109,N_11272,N_12138);
nor U15110 (N_15110,N_9898,N_11053);
nand U15111 (N_15111,N_10248,N_11094);
nand U15112 (N_15112,N_10373,N_12019);
and U15113 (N_15113,N_9563,N_10274);
nor U15114 (N_15114,N_11978,N_12214);
and U15115 (N_15115,N_12159,N_10769);
xor U15116 (N_15116,N_11678,N_12458);
xor U15117 (N_15117,N_12260,N_11113);
and U15118 (N_15118,N_11893,N_10617);
xnor U15119 (N_15119,N_11988,N_10183);
nor U15120 (N_15120,N_9967,N_12118);
nand U15121 (N_15121,N_11523,N_11791);
or U15122 (N_15122,N_10073,N_11729);
nor U15123 (N_15123,N_10829,N_11999);
or U15124 (N_15124,N_11701,N_10332);
or U15125 (N_15125,N_10483,N_10270);
nand U15126 (N_15126,N_12214,N_10358);
and U15127 (N_15127,N_12424,N_9596);
nand U15128 (N_15128,N_10506,N_10587);
nand U15129 (N_15129,N_12014,N_12280);
or U15130 (N_15130,N_11963,N_10197);
nor U15131 (N_15131,N_9904,N_10461);
nand U15132 (N_15132,N_11350,N_9897);
or U15133 (N_15133,N_10742,N_12372);
or U15134 (N_15134,N_12362,N_9813);
and U15135 (N_15135,N_9892,N_10456);
nor U15136 (N_15136,N_9662,N_9569);
or U15137 (N_15137,N_9823,N_9547);
nor U15138 (N_15138,N_9695,N_10119);
xor U15139 (N_15139,N_11734,N_10600);
xor U15140 (N_15140,N_10450,N_10924);
and U15141 (N_15141,N_9916,N_11826);
nand U15142 (N_15142,N_10646,N_11945);
xor U15143 (N_15143,N_11525,N_10222);
or U15144 (N_15144,N_10452,N_9985);
xor U15145 (N_15145,N_11290,N_10517);
xor U15146 (N_15146,N_10993,N_10322);
nor U15147 (N_15147,N_11468,N_12443);
or U15148 (N_15148,N_10660,N_12312);
xor U15149 (N_15149,N_10502,N_12381);
nand U15150 (N_15150,N_11404,N_10461);
or U15151 (N_15151,N_11702,N_12032);
xnor U15152 (N_15152,N_12141,N_10156);
and U15153 (N_15153,N_12136,N_10728);
or U15154 (N_15154,N_10414,N_9572);
xor U15155 (N_15155,N_10729,N_10620);
or U15156 (N_15156,N_11052,N_11995);
or U15157 (N_15157,N_10326,N_10440);
and U15158 (N_15158,N_11023,N_10297);
xor U15159 (N_15159,N_10466,N_9614);
xor U15160 (N_15160,N_10628,N_9879);
or U15161 (N_15161,N_10514,N_12430);
nand U15162 (N_15162,N_11502,N_11817);
xnor U15163 (N_15163,N_11762,N_10473);
nand U15164 (N_15164,N_9404,N_11816);
nand U15165 (N_15165,N_10417,N_11897);
nand U15166 (N_15166,N_11410,N_11462);
and U15167 (N_15167,N_11553,N_9989);
and U15168 (N_15168,N_11351,N_11326);
xor U15169 (N_15169,N_9555,N_11161);
and U15170 (N_15170,N_11842,N_11247);
or U15171 (N_15171,N_12055,N_12417);
nor U15172 (N_15172,N_9707,N_10441);
and U15173 (N_15173,N_10205,N_10430);
xnor U15174 (N_15174,N_12231,N_11118);
or U15175 (N_15175,N_10785,N_10381);
xor U15176 (N_15176,N_11407,N_12473);
or U15177 (N_15177,N_10454,N_10336);
xnor U15178 (N_15178,N_10580,N_11395);
or U15179 (N_15179,N_11040,N_12001);
nand U15180 (N_15180,N_11131,N_11407);
xnor U15181 (N_15181,N_12367,N_12066);
xnor U15182 (N_15182,N_11448,N_12403);
or U15183 (N_15183,N_9763,N_12232);
and U15184 (N_15184,N_12078,N_12267);
nor U15185 (N_15185,N_12170,N_10694);
xnor U15186 (N_15186,N_10028,N_12357);
or U15187 (N_15187,N_11977,N_12161);
or U15188 (N_15188,N_10897,N_10115);
nand U15189 (N_15189,N_12107,N_11445);
and U15190 (N_15190,N_10030,N_10913);
or U15191 (N_15191,N_10191,N_12183);
xnor U15192 (N_15192,N_10334,N_9694);
nor U15193 (N_15193,N_12338,N_12225);
nand U15194 (N_15194,N_9962,N_11183);
xnor U15195 (N_15195,N_10702,N_9428);
nand U15196 (N_15196,N_9946,N_11822);
nand U15197 (N_15197,N_11386,N_10605);
or U15198 (N_15198,N_9792,N_10573);
or U15199 (N_15199,N_12132,N_9704);
nor U15200 (N_15200,N_11247,N_10410);
and U15201 (N_15201,N_11054,N_10818);
and U15202 (N_15202,N_9900,N_9849);
nor U15203 (N_15203,N_11926,N_9598);
xor U15204 (N_15204,N_10492,N_11035);
xnor U15205 (N_15205,N_10964,N_12370);
and U15206 (N_15206,N_9943,N_9504);
xnor U15207 (N_15207,N_10194,N_11050);
nor U15208 (N_15208,N_11931,N_10151);
nand U15209 (N_15209,N_11395,N_10933);
and U15210 (N_15210,N_10825,N_10074);
xor U15211 (N_15211,N_9533,N_9471);
and U15212 (N_15212,N_12272,N_10757);
nor U15213 (N_15213,N_12124,N_9984);
nand U15214 (N_15214,N_11466,N_9969);
xor U15215 (N_15215,N_11935,N_12020);
nor U15216 (N_15216,N_11627,N_9731);
and U15217 (N_15217,N_12309,N_11757);
nor U15218 (N_15218,N_11308,N_12202);
nor U15219 (N_15219,N_9568,N_11694);
nor U15220 (N_15220,N_10652,N_10085);
or U15221 (N_15221,N_12404,N_12085);
xnor U15222 (N_15222,N_9964,N_11071);
nand U15223 (N_15223,N_11500,N_10860);
nand U15224 (N_15224,N_10078,N_10753);
nor U15225 (N_15225,N_10116,N_10039);
and U15226 (N_15226,N_12393,N_11565);
nor U15227 (N_15227,N_10686,N_11958);
nand U15228 (N_15228,N_10587,N_11597);
and U15229 (N_15229,N_10385,N_12065);
and U15230 (N_15230,N_11590,N_9586);
and U15231 (N_15231,N_10405,N_11565);
and U15232 (N_15232,N_11449,N_11218);
and U15233 (N_15233,N_12349,N_10974);
nor U15234 (N_15234,N_12352,N_11470);
nand U15235 (N_15235,N_12244,N_9614);
nor U15236 (N_15236,N_9680,N_11484);
and U15237 (N_15237,N_10755,N_9884);
or U15238 (N_15238,N_11455,N_10378);
nor U15239 (N_15239,N_12360,N_10343);
xor U15240 (N_15240,N_10001,N_10491);
or U15241 (N_15241,N_10001,N_10500);
xnor U15242 (N_15242,N_11628,N_11005);
nor U15243 (N_15243,N_11565,N_11279);
or U15244 (N_15244,N_12355,N_10122);
xor U15245 (N_15245,N_10800,N_11739);
nand U15246 (N_15246,N_10582,N_12125);
and U15247 (N_15247,N_9598,N_10817);
nor U15248 (N_15248,N_10923,N_10598);
xor U15249 (N_15249,N_12073,N_11175);
nor U15250 (N_15250,N_10173,N_11684);
nand U15251 (N_15251,N_12206,N_10620);
and U15252 (N_15252,N_12307,N_11441);
nor U15253 (N_15253,N_11507,N_10786);
or U15254 (N_15254,N_9995,N_12010);
nand U15255 (N_15255,N_10025,N_9968);
nand U15256 (N_15256,N_9380,N_12393);
nand U15257 (N_15257,N_9645,N_10234);
xnor U15258 (N_15258,N_11163,N_10809);
xnor U15259 (N_15259,N_11631,N_11887);
nand U15260 (N_15260,N_11321,N_9889);
or U15261 (N_15261,N_10680,N_11968);
or U15262 (N_15262,N_11888,N_11029);
and U15263 (N_15263,N_9790,N_10238);
or U15264 (N_15264,N_10427,N_10454);
nand U15265 (N_15265,N_11316,N_10764);
nor U15266 (N_15266,N_9468,N_9587);
nand U15267 (N_15267,N_12380,N_11337);
xor U15268 (N_15268,N_9920,N_11509);
or U15269 (N_15269,N_11000,N_12386);
nand U15270 (N_15270,N_12288,N_11820);
nand U15271 (N_15271,N_10547,N_10900);
or U15272 (N_15272,N_11505,N_9908);
nand U15273 (N_15273,N_9518,N_11117);
nand U15274 (N_15274,N_10399,N_11786);
or U15275 (N_15275,N_10591,N_9857);
nand U15276 (N_15276,N_10291,N_12017);
or U15277 (N_15277,N_10026,N_10243);
xnor U15278 (N_15278,N_10453,N_10415);
and U15279 (N_15279,N_11322,N_12151);
xnor U15280 (N_15280,N_9943,N_9764);
xor U15281 (N_15281,N_11147,N_9481);
nor U15282 (N_15282,N_11224,N_10715);
or U15283 (N_15283,N_11819,N_10289);
nand U15284 (N_15284,N_10740,N_11566);
nand U15285 (N_15285,N_10555,N_10253);
or U15286 (N_15286,N_10015,N_11153);
or U15287 (N_15287,N_11848,N_9903);
nand U15288 (N_15288,N_11020,N_11598);
or U15289 (N_15289,N_11835,N_10599);
or U15290 (N_15290,N_11858,N_10277);
and U15291 (N_15291,N_10934,N_11712);
nand U15292 (N_15292,N_10830,N_9848);
xnor U15293 (N_15293,N_11453,N_10746);
or U15294 (N_15294,N_10564,N_12480);
nand U15295 (N_15295,N_12473,N_11199);
nand U15296 (N_15296,N_10429,N_10717);
nor U15297 (N_15297,N_10756,N_10471);
nand U15298 (N_15298,N_12405,N_10499);
and U15299 (N_15299,N_10376,N_10987);
nand U15300 (N_15300,N_10285,N_9587);
or U15301 (N_15301,N_9731,N_11230);
nor U15302 (N_15302,N_10713,N_11373);
xnor U15303 (N_15303,N_9545,N_10700);
xor U15304 (N_15304,N_12417,N_12035);
and U15305 (N_15305,N_11325,N_12043);
xnor U15306 (N_15306,N_11064,N_11364);
nand U15307 (N_15307,N_9775,N_9474);
and U15308 (N_15308,N_12420,N_10352);
xnor U15309 (N_15309,N_10449,N_11844);
and U15310 (N_15310,N_9910,N_9776);
nand U15311 (N_15311,N_11507,N_11476);
nor U15312 (N_15312,N_10789,N_12087);
nor U15313 (N_15313,N_12134,N_9629);
nor U15314 (N_15314,N_10827,N_12355);
nand U15315 (N_15315,N_10354,N_11851);
nand U15316 (N_15316,N_10368,N_10403);
xnor U15317 (N_15317,N_12461,N_10525);
nor U15318 (N_15318,N_10238,N_9660);
and U15319 (N_15319,N_11597,N_11665);
or U15320 (N_15320,N_12386,N_9594);
nand U15321 (N_15321,N_11287,N_11277);
and U15322 (N_15322,N_11303,N_9498);
nor U15323 (N_15323,N_11041,N_10954);
nor U15324 (N_15324,N_10236,N_11106);
xnor U15325 (N_15325,N_10297,N_9654);
nand U15326 (N_15326,N_11086,N_9452);
and U15327 (N_15327,N_11354,N_12349);
or U15328 (N_15328,N_10860,N_12063);
and U15329 (N_15329,N_9577,N_9545);
nand U15330 (N_15330,N_12109,N_11640);
and U15331 (N_15331,N_10861,N_10770);
and U15332 (N_15332,N_12242,N_11538);
and U15333 (N_15333,N_10782,N_10619);
and U15334 (N_15334,N_10666,N_11068);
nand U15335 (N_15335,N_11065,N_12339);
nor U15336 (N_15336,N_11703,N_12113);
nand U15337 (N_15337,N_12328,N_11604);
and U15338 (N_15338,N_11089,N_11236);
nor U15339 (N_15339,N_11727,N_11229);
nand U15340 (N_15340,N_11657,N_10845);
nand U15341 (N_15341,N_11412,N_10244);
nor U15342 (N_15342,N_10319,N_11160);
and U15343 (N_15343,N_12016,N_11967);
and U15344 (N_15344,N_11726,N_9888);
nand U15345 (N_15345,N_11436,N_11889);
nor U15346 (N_15346,N_11166,N_11343);
xnor U15347 (N_15347,N_11941,N_11118);
and U15348 (N_15348,N_11490,N_12448);
nor U15349 (N_15349,N_11591,N_11202);
nand U15350 (N_15350,N_9389,N_11580);
and U15351 (N_15351,N_11402,N_11277);
nand U15352 (N_15352,N_10306,N_10041);
xnor U15353 (N_15353,N_10243,N_12152);
and U15354 (N_15354,N_10117,N_11509);
or U15355 (N_15355,N_10730,N_10583);
nand U15356 (N_15356,N_10717,N_12277);
nand U15357 (N_15357,N_11521,N_9568);
nand U15358 (N_15358,N_11449,N_11403);
nand U15359 (N_15359,N_12427,N_10506);
nand U15360 (N_15360,N_12411,N_12191);
xor U15361 (N_15361,N_11766,N_10929);
xor U15362 (N_15362,N_10902,N_11532);
nor U15363 (N_15363,N_9735,N_11290);
nor U15364 (N_15364,N_11170,N_11946);
xor U15365 (N_15365,N_12484,N_10740);
nor U15366 (N_15366,N_10130,N_11466);
nor U15367 (N_15367,N_10144,N_9898);
and U15368 (N_15368,N_11978,N_10858);
nor U15369 (N_15369,N_10918,N_10993);
or U15370 (N_15370,N_10772,N_10803);
nor U15371 (N_15371,N_11815,N_10276);
nand U15372 (N_15372,N_10267,N_11659);
or U15373 (N_15373,N_10391,N_10816);
or U15374 (N_15374,N_9460,N_11182);
nor U15375 (N_15375,N_9986,N_11756);
xor U15376 (N_15376,N_12355,N_11084);
and U15377 (N_15377,N_10552,N_10801);
and U15378 (N_15378,N_9388,N_11743);
nor U15379 (N_15379,N_12404,N_11157);
xnor U15380 (N_15380,N_11645,N_9835);
or U15381 (N_15381,N_10141,N_11427);
or U15382 (N_15382,N_11294,N_12258);
or U15383 (N_15383,N_11524,N_11039);
and U15384 (N_15384,N_10074,N_12194);
and U15385 (N_15385,N_10853,N_12449);
and U15386 (N_15386,N_10010,N_12309);
nand U15387 (N_15387,N_9774,N_12413);
nor U15388 (N_15388,N_11517,N_10732);
or U15389 (N_15389,N_11519,N_10983);
xor U15390 (N_15390,N_10602,N_12178);
nor U15391 (N_15391,N_11195,N_10776);
and U15392 (N_15392,N_12044,N_9822);
xnor U15393 (N_15393,N_11195,N_9572);
xor U15394 (N_15394,N_11818,N_10363);
nor U15395 (N_15395,N_12178,N_11100);
xnor U15396 (N_15396,N_9402,N_10606);
xor U15397 (N_15397,N_10193,N_11429);
and U15398 (N_15398,N_12336,N_9866);
or U15399 (N_15399,N_10816,N_11399);
nor U15400 (N_15400,N_11366,N_9659);
or U15401 (N_15401,N_10562,N_11237);
or U15402 (N_15402,N_9826,N_10513);
or U15403 (N_15403,N_12425,N_11195);
xor U15404 (N_15404,N_11942,N_11220);
nand U15405 (N_15405,N_10151,N_12420);
nand U15406 (N_15406,N_10288,N_12195);
or U15407 (N_15407,N_10263,N_10340);
or U15408 (N_15408,N_11137,N_11007);
nand U15409 (N_15409,N_11054,N_10166);
or U15410 (N_15410,N_12492,N_9639);
nor U15411 (N_15411,N_12169,N_11661);
nor U15412 (N_15412,N_10699,N_10038);
xnor U15413 (N_15413,N_10837,N_11050);
xnor U15414 (N_15414,N_11552,N_10563);
and U15415 (N_15415,N_12211,N_9773);
xnor U15416 (N_15416,N_9992,N_10509);
or U15417 (N_15417,N_10961,N_10469);
or U15418 (N_15418,N_11696,N_11748);
nor U15419 (N_15419,N_12332,N_9973);
nand U15420 (N_15420,N_9867,N_11176);
or U15421 (N_15421,N_10653,N_11303);
or U15422 (N_15422,N_11758,N_10235);
nor U15423 (N_15423,N_10783,N_12099);
nor U15424 (N_15424,N_10696,N_11521);
nand U15425 (N_15425,N_9861,N_10959);
or U15426 (N_15426,N_11835,N_12450);
or U15427 (N_15427,N_12340,N_11441);
xnor U15428 (N_15428,N_11685,N_12450);
and U15429 (N_15429,N_11489,N_11935);
nor U15430 (N_15430,N_12038,N_9718);
or U15431 (N_15431,N_11816,N_10357);
nor U15432 (N_15432,N_9821,N_9927);
and U15433 (N_15433,N_11540,N_12192);
xnor U15434 (N_15434,N_11491,N_11111);
nor U15435 (N_15435,N_12057,N_9956);
and U15436 (N_15436,N_10797,N_11169);
nand U15437 (N_15437,N_11106,N_9978);
xor U15438 (N_15438,N_11744,N_11364);
xnor U15439 (N_15439,N_11984,N_10011);
nor U15440 (N_15440,N_11019,N_10617);
nand U15441 (N_15441,N_11824,N_11944);
nand U15442 (N_15442,N_10990,N_10646);
xor U15443 (N_15443,N_12265,N_11437);
nor U15444 (N_15444,N_10580,N_10640);
and U15445 (N_15445,N_10295,N_12432);
nor U15446 (N_15446,N_10278,N_11244);
xor U15447 (N_15447,N_9405,N_12127);
nand U15448 (N_15448,N_11872,N_10483);
nor U15449 (N_15449,N_11850,N_11738);
xor U15450 (N_15450,N_11739,N_10748);
nand U15451 (N_15451,N_11988,N_11632);
or U15452 (N_15452,N_12480,N_10126);
nor U15453 (N_15453,N_10746,N_10976);
nor U15454 (N_15454,N_10864,N_11761);
or U15455 (N_15455,N_9453,N_11828);
nor U15456 (N_15456,N_11414,N_12000);
nor U15457 (N_15457,N_9455,N_11109);
nand U15458 (N_15458,N_11133,N_9941);
xnor U15459 (N_15459,N_11225,N_12285);
nand U15460 (N_15460,N_9663,N_12301);
or U15461 (N_15461,N_11150,N_9624);
nand U15462 (N_15462,N_10070,N_9764);
and U15463 (N_15463,N_11377,N_10825);
and U15464 (N_15464,N_10858,N_10889);
xnor U15465 (N_15465,N_10485,N_11704);
and U15466 (N_15466,N_10455,N_11606);
and U15467 (N_15467,N_11995,N_10662);
and U15468 (N_15468,N_9653,N_10353);
xnor U15469 (N_15469,N_9534,N_12281);
and U15470 (N_15470,N_10716,N_10838);
nor U15471 (N_15471,N_11800,N_12068);
nor U15472 (N_15472,N_10446,N_11684);
or U15473 (N_15473,N_9604,N_10349);
nand U15474 (N_15474,N_10960,N_9679);
or U15475 (N_15475,N_10982,N_12140);
xor U15476 (N_15476,N_11063,N_10069);
nand U15477 (N_15477,N_12313,N_9808);
xnor U15478 (N_15478,N_12152,N_10686);
xor U15479 (N_15479,N_11950,N_9896);
nand U15480 (N_15480,N_9425,N_11731);
nand U15481 (N_15481,N_12189,N_9492);
xnor U15482 (N_15482,N_10271,N_10744);
xnor U15483 (N_15483,N_11360,N_12093);
or U15484 (N_15484,N_11000,N_11505);
nor U15485 (N_15485,N_11672,N_12429);
nand U15486 (N_15486,N_10261,N_11615);
or U15487 (N_15487,N_11132,N_11245);
and U15488 (N_15488,N_11613,N_11087);
nor U15489 (N_15489,N_9974,N_9747);
and U15490 (N_15490,N_11420,N_9899);
or U15491 (N_15491,N_10366,N_11415);
nand U15492 (N_15492,N_12433,N_10095);
or U15493 (N_15493,N_10215,N_9709);
nand U15494 (N_15494,N_11296,N_10653);
or U15495 (N_15495,N_10266,N_12439);
xor U15496 (N_15496,N_11141,N_10932);
and U15497 (N_15497,N_10926,N_11202);
nor U15498 (N_15498,N_12135,N_10059);
or U15499 (N_15499,N_11245,N_9608);
xnor U15500 (N_15500,N_10488,N_9821);
xor U15501 (N_15501,N_10081,N_9802);
or U15502 (N_15502,N_9838,N_11564);
nor U15503 (N_15503,N_11680,N_10702);
nor U15504 (N_15504,N_10685,N_10406);
xor U15505 (N_15505,N_11605,N_11924);
xnor U15506 (N_15506,N_9399,N_10754);
and U15507 (N_15507,N_9593,N_10606);
xnor U15508 (N_15508,N_9532,N_10381);
or U15509 (N_15509,N_11764,N_10230);
nor U15510 (N_15510,N_9621,N_9916);
nor U15511 (N_15511,N_11690,N_10808);
nand U15512 (N_15512,N_11108,N_11959);
xnor U15513 (N_15513,N_10685,N_10057);
nand U15514 (N_15514,N_9694,N_9464);
nand U15515 (N_15515,N_10953,N_9712);
or U15516 (N_15516,N_11894,N_9992);
and U15517 (N_15517,N_11741,N_9970);
nand U15518 (N_15518,N_10739,N_11841);
nand U15519 (N_15519,N_10926,N_10479);
nand U15520 (N_15520,N_10053,N_11544);
xor U15521 (N_15521,N_10604,N_11799);
or U15522 (N_15522,N_9769,N_11702);
nor U15523 (N_15523,N_11425,N_11528);
nor U15524 (N_15524,N_9815,N_12242);
or U15525 (N_15525,N_10429,N_11150);
or U15526 (N_15526,N_9448,N_11427);
nor U15527 (N_15527,N_11741,N_11170);
nor U15528 (N_15528,N_11334,N_9961);
and U15529 (N_15529,N_10467,N_11907);
and U15530 (N_15530,N_11290,N_9757);
nor U15531 (N_15531,N_12429,N_12482);
nor U15532 (N_15532,N_11349,N_12316);
or U15533 (N_15533,N_11815,N_9471);
and U15534 (N_15534,N_10645,N_11802);
nor U15535 (N_15535,N_11665,N_11233);
or U15536 (N_15536,N_11059,N_10158);
and U15537 (N_15537,N_11524,N_10852);
and U15538 (N_15538,N_12396,N_11111);
nand U15539 (N_15539,N_10456,N_9937);
or U15540 (N_15540,N_11687,N_10536);
or U15541 (N_15541,N_9661,N_10869);
nor U15542 (N_15542,N_11124,N_12166);
nor U15543 (N_15543,N_9709,N_9785);
xnor U15544 (N_15544,N_11666,N_9982);
nor U15545 (N_15545,N_12451,N_11002);
and U15546 (N_15546,N_10616,N_12183);
nand U15547 (N_15547,N_10731,N_9731);
nor U15548 (N_15548,N_11209,N_12037);
nand U15549 (N_15549,N_11514,N_10391);
nand U15550 (N_15550,N_11115,N_12459);
nor U15551 (N_15551,N_11901,N_11605);
nand U15552 (N_15552,N_10330,N_11361);
and U15553 (N_15553,N_10057,N_9496);
nor U15554 (N_15554,N_10553,N_10859);
xor U15555 (N_15555,N_11826,N_10590);
nor U15556 (N_15556,N_12140,N_9717);
nor U15557 (N_15557,N_11813,N_9897);
xnor U15558 (N_15558,N_11256,N_10972);
and U15559 (N_15559,N_12071,N_11894);
and U15560 (N_15560,N_12138,N_12066);
or U15561 (N_15561,N_12305,N_10383);
nand U15562 (N_15562,N_9537,N_11706);
and U15563 (N_15563,N_9963,N_9588);
xnor U15564 (N_15564,N_10447,N_9508);
and U15565 (N_15565,N_9798,N_11082);
xnor U15566 (N_15566,N_12024,N_11838);
nor U15567 (N_15567,N_9489,N_10361);
xor U15568 (N_15568,N_11157,N_11491);
nand U15569 (N_15569,N_10054,N_11783);
nand U15570 (N_15570,N_9454,N_10070);
nor U15571 (N_15571,N_11312,N_9585);
nand U15572 (N_15572,N_11012,N_10031);
nor U15573 (N_15573,N_9980,N_10833);
or U15574 (N_15574,N_9449,N_11984);
or U15575 (N_15575,N_12148,N_11801);
nor U15576 (N_15576,N_9666,N_12388);
nor U15577 (N_15577,N_10073,N_10135);
xor U15578 (N_15578,N_10509,N_12422);
and U15579 (N_15579,N_12379,N_10402);
and U15580 (N_15580,N_11272,N_12161);
nand U15581 (N_15581,N_9755,N_9664);
or U15582 (N_15582,N_9849,N_11327);
and U15583 (N_15583,N_11427,N_10582);
xnor U15584 (N_15584,N_11122,N_10765);
nor U15585 (N_15585,N_11399,N_9815);
nand U15586 (N_15586,N_11702,N_10567);
and U15587 (N_15587,N_12112,N_9987);
or U15588 (N_15588,N_11713,N_10693);
xor U15589 (N_15589,N_9405,N_11826);
nand U15590 (N_15590,N_9679,N_9855);
nor U15591 (N_15591,N_11232,N_9419);
nor U15592 (N_15592,N_12365,N_11711);
nand U15593 (N_15593,N_10815,N_11141);
and U15594 (N_15594,N_9848,N_10902);
or U15595 (N_15595,N_10238,N_11775);
or U15596 (N_15596,N_10182,N_9886);
nor U15597 (N_15597,N_9715,N_9497);
nor U15598 (N_15598,N_10424,N_10221);
xor U15599 (N_15599,N_10053,N_11968);
or U15600 (N_15600,N_11633,N_11618);
nor U15601 (N_15601,N_10881,N_10552);
or U15602 (N_15602,N_10362,N_12369);
nand U15603 (N_15603,N_11810,N_9974);
nand U15604 (N_15604,N_10735,N_10113);
nor U15605 (N_15605,N_10273,N_10448);
nand U15606 (N_15606,N_9995,N_12127);
and U15607 (N_15607,N_10955,N_9460);
or U15608 (N_15608,N_12468,N_11743);
and U15609 (N_15609,N_12337,N_10228);
or U15610 (N_15610,N_12472,N_9604);
nand U15611 (N_15611,N_10569,N_11129);
nor U15612 (N_15612,N_10557,N_12447);
nor U15613 (N_15613,N_9927,N_11094);
or U15614 (N_15614,N_10135,N_12290);
xor U15615 (N_15615,N_11202,N_11939);
or U15616 (N_15616,N_11465,N_9843);
nor U15617 (N_15617,N_11279,N_10464);
nand U15618 (N_15618,N_10279,N_12046);
or U15619 (N_15619,N_11887,N_12118);
and U15620 (N_15620,N_11310,N_10957);
nor U15621 (N_15621,N_9760,N_10326);
and U15622 (N_15622,N_9857,N_10453);
nor U15623 (N_15623,N_9834,N_12193);
nand U15624 (N_15624,N_10290,N_11115);
and U15625 (N_15625,N_14044,N_12573);
nand U15626 (N_15626,N_13722,N_14387);
nor U15627 (N_15627,N_13031,N_13934);
xnor U15628 (N_15628,N_14606,N_15209);
xor U15629 (N_15629,N_15294,N_13056);
and U15630 (N_15630,N_14610,N_13775);
and U15631 (N_15631,N_12774,N_12500);
nand U15632 (N_15632,N_14503,N_15512);
or U15633 (N_15633,N_15271,N_15088);
xnor U15634 (N_15634,N_14195,N_13490);
xor U15635 (N_15635,N_12601,N_13165);
xnor U15636 (N_15636,N_13032,N_14285);
nand U15637 (N_15637,N_12881,N_15003);
nor U15638 (N_15638,N_15538,N_12989);
and U15639 (N_15639,N_13250,N_13900);
and U15640 (N_15640,N_15492,N_15503);
xor U15641 (N_15641,N_13871,N_15035);
and U15642 (N_15642,N_14164,N_14047);
or U15643 (N_15643,N_15004,N_13870);
or U15644 (N_15644,N_12505,N_13478);
nand U15645 (N_15645,N_13026,N_15570);
or U15646 (N_15646,N_15133,N_12713);
nand U15647 (N_15647,N_14201,N_13242);
nor U15648 (N_15648,N_12818,N_12645);
and U15649 (N_15649,N_15379,N_14672);
nor U15650 (N_15650,N_14985,N_13646);
nor U15651 (N_15651,N_15285,N_15459);
nand U15652 (N_15652,N_14323,N_12787);
or U15653 (N_15653,N_13517,N_15486);
nand U15654 (N_15654,N_15001,N_13547);
nand U15655 (N_15655,N_14141,N_15248);
and U15656 (N_15656,N_13773,N_12673);
or U15657 (N_15657,N_14296,N_15615);
or U15658 (N_15658,N_14349,N_12718);
xnor U15659 (N_15659,N_14601,N_13048);
xnor U15660 (N_15660,N_14984,N_14670);
and U15661 (N_15661,N_13066,N_12501);
nor U15662 (N_15662,N_14171,N_13702);
and U15663 (N_15663,N_15465,N_13541);
xnor U15664 (N_15664,N_14170,N_14350);
nor U15665 (N_15665,N_13125,N_13312);
xnor U15666 (N_15666,N_14098,N_14854);
and U15667 (N_15667,N_12855,N_13064);
nand U15668 (N_15668,N_13703,N_12865);
xnor U15669 (N_15669,N_12981,N_14504);
xor U15670 (N_15670,N_15147,N_15124);
xnor U15671 (N_15671,N_15603,N_13856);
and U15672 (N_15672,N_13169,N_14911);
nand U15673 (N_15673,N_14915,N_13384);
nand U15674 (N_15674,N_14219,N_15373);
nor U15675 (N_15675,N_13415,N_13206);
or U15676 (N_15676,N_13244,N_13099);
and U15677 (N_15677,N_15278,N_12803);
and U15678 (N_15678,N_12832,N_13552);
nand U15679 (N_15679,N_13075,N_15410);
and U15680 (N_15680,N_14161,N_13661);
nor U15681 (N_15681,N_14183,N_14810);
nand U15682 (N_15682,N_13698,N_14925);
or U15683 (N_15683,N_15036,N_15113);
xnor U15684 (N_15684,N_14301,N_14591);
xor U15685 (N_15685,N_14423,N_14530);
and U15686 (N_15686,N_15165,N_14172);
nor U15687 (N_15687,N_14325,N_14061);
xor U15688 (N_15688,N_14443,N_15376);
xnor U15689 (N_15689,N_15094,N_13969);
nor U15690 (N_15690,N_13989,N_13264);
xor U15691 (N_15691,N_14176,N_14033);
or U15692 (N_15692,N_12871,N_13378);
nor U15693 (N_15693,N_14807,N_14457);
nor U15694 (N_15694,N_15554,N_13493);
nand U15695 (N_15695,N_14417,N_14905);
xor U15696 (N_15696,N_15108,N_15205);
and U15697 (N_15697,N_13807,N_15276);
or U15698 (N_15698,N_13874,N_14022);
or U15699 (N_15699,N_14151,N_13053);
xor U15700 (N_15700,N_12559,N_14186);
nand U15701 (N_15701,N_12754,N_14050);
and U15702 (N_15702,N_15284,N_15065);
or U15703 (N_15703,N_13472,N_14036);
nor U15704 (N_15704,N_14346,N_13611);
xor U15705 (N_15705,N_13893,N_13291);
and U15706 (N_15706,N_13286,N_14641);
and U15707 (N_15707,N_14676,N_14834);
nand U15708 (N_15708,N_13952,N_15167);
or U15709 (N_15709,N_14785,N_13281);
and U15710 (N_15710,N_13944,N_14305);
nand U15711 (N_15711,N_14225,N_13531);
or U15712 (N_15712,N_14193,N_13802);
and U15713 (N_15713,N_15493,N_14567);
nand U15714 (N_15714,N_12536,N_13367);
nor U15715 (N_15715,N_12615,N_15595);
nand U15716 (N_15716,N_13859,N_15236);
nand U15717 (N_15717,N_15090,N_12892);
nor U15718 (N_15718,N_14966,N_15196);
and U15719 (N_15719,N_13007,N_15401);
and U15720 (N_15720,N_15234,N_13683);
nand U15721 (N_15721,N_15115,N_14689);
xor U15722 (N_15722,N_13507,N_14144);
or U15723 (N_15723,N_15238,N_12912);
xor U15724 (N_15724,N_12627,N_14125);
and U15725 (N_15725,N_13176,N_15008);
and U15726 (N_15726,N_14024,N_14425);
nor U15727 (N_15727,N_14717,N_14989);
nand U15728 (N_15728,N_14939,N_13070);
nor U15729 (N_15729,N_12745,N_13821);
nand U15730 (N_15730,N_15363,N_13835);
nand U15731 (N_15731,N_12691,N_14001);
nor U15732 (N_15732,N_13783,N_12709);
and U15733 (N_15733,N_15227,N_13498);
and U15734 (N_15734,N_15589,N_13950);
and U15735 (N_15735,N_14986,N_13617);
nand U15736 (N_15736,N_14298,N_15349);
and U15737 (N_15737,N_12917,N_14786);
nand U15738 (N_15738,N_13529,N_12593);
and U15739 (N_15739,N_13423,N_14299);
or U15740 (N_15740,N_15142,N_13596);
or U15741 (N_15741,N_13267,N_13920);
xnor U15742 (N_15742,N_13522,N_15571);
or U15743 (N_15743,N_13956,N_12863);
nor U15744 (N_15744,N_13413,N_15028);
and U15745 (N_15745,N_15219,N_15399);
nor U15746 (N_15746,N_13135,N_13542);
xnor U15747 (N_15747,N_13284,N_12888);
nand U15748 (N_15748,N_14344,N_14005);
nor U15749 (N_15749,N_14289,N_15352);
nor U15750 (N_15750,N_13028,N_15599);
nand U15751 (N_15751,N_14435,N_14572);
or U15752 (N_15752,N_14592,N_14332);
nor U15753 (N_15753,N_15509,N_15327);
or U15754 (N_15754,N_15257,N_13548);
nor U15755 (N_15755,N_12646,N_14231);
and U15756 (N_15756,N_13393,N_13084);
nand U15757 (N_15757,N_14732,N_15267);
and U15758 (N_15758,N_14877,N_13919);
xnor U15759 (N_15759,N_14103,N_12607);
nor U15760 (N_15760,N_13477,N_14267);
xor U15761 (N_15761,N_15160,N_15223);
or U15762 (N_15762,N_12983,N_12827);
xnor U15763 (N_15763,N_15273,N_14642);
nor U15764 (N_15764,N_14449,N_13023);
nand U15765 (N_15765,N_15573,N_14744);
xnor U15766 (N_15766,N_14916,N_15302);
nor U15767 (N_15767,N_12920,N_13623);
nor U15768 (N_15768,N_13037,N_13705);
xnor U15769 (N_15769,N_14228,N_13838);
and U15770 (N_15770,N_13771,N_13685);
nand U15771 (N_15771,N_15254,N_15188);
and U15772 (N_15772,N_13012,N_14018);
and U15773 (N_15773,N_14499,N_14181);
and U15774 (N_15774,N_13813,N_14278);
nor U15775 (N_15775,N_13076,N_13229);
or U15776 (N_15776,N_12711,N_14060);
nand U15777 (N_15777,N_13655,N_13690);
or U15778 (N_15778,N_14890,N_13193);
nand U15779 (N_15779,N_12659,N_14317);
or U15780 (N_15780,N_12651,N_15092);
or U15781 (N_15781,N_15555,N_14869);
or U15782 (N_15782,N_14666,N_14166);
and U15783 (N_15783,N_12597,N_15025);
nand U15784 (N_15784,N_14716,N_14462);
nor U15785 (N_15785,N_12828,N_14092);
and U15786 (N_15786,N_14746,N_13155);
nand U15787 (N_15787,N_15344,N_14356);
and U15788 (N_15788,N_14973,N_13297);
nand U15789 (N_15789,N_13659,N_15045);
and U15790 (N_15790,N_14863,N_15384);
nand U15791 (N_15791,N_14607,N_14284);
xor U15792 (N_15792,N_12668,N_13963);
nor U15793 (N_15793,N_13743,N_14002);
nand U15794 (N_15794,N_13373,N_13781);
or U15795 (N_15795,N_15048,N_14808);
and U15796 (N_15796,N_13767,N_14742);
nand U15797 (N_15797,N_15433,N_13146);
or U15798 (N_15798,N_14197,N_13330);
nor U15799 (N_15799,N_13207,N_13129);
and U15800 (N_15800,N_14494,N_14371);
nor U15801 (N_15801,N_15545,N_15063);
xnor U15802 (N_15802,N_14945,N_12901);
nor U15803 (N_15803,N_13201,N_15371);
nand U15804 (N_15804,N_15128,N_13454);
and U15805 (N_15805,N_13553,N_13689);
xor U15806 (N_15806,N_14375,N_12781);
nor U15807 (N_15807,N_12548,N_13977);
nand U15808 (N_15808,N_14380,N_15221);
xnor U15809 (N_15809,N_13846,N_13828);
xor U15810 (N_15810,N_13383,N_12882);
xnor U15811 (N_15811,N_14980,N_12686);
and U15812 (N_15812,N_12734,N_12523);
nand U15813 (N_15813,N_14010,N_14426);
nand U15814 (N_15814,N_14698,N_12879);
nand U15815 (N_15815,N_12589,N_15397);
nor U15816 (N_15816,N_13959,N_15089);
nor U15817 (N_15817,N_13170,N_12546);
nand U15818 (N_15818,N_14561,N_14922);
nand U15819 (N_15819,N_12928,N_15068);
and U15820 (N_15820,N_13868,N_13460);
nand U15821 (N_15821,N_13039,N_15579);
nor U15822 (N_15822,N_14329,N_13220);
nor U15823 (N_15823,N_15533,N_15015);
or U15824 (N_15824,N_13530,N_15307);
xor U15825 (N_15825,N_15064,N_12698);
xnor U15826 (N_15826,N_13386,N_13883);
xor U15827 (N_15827,N_13480,N_14415);
xnor U15828 (N_15828,N_15342,N_14846);
nand U15829 (N_15829,N_14832,N_14995);
xnor U15830 (N_15830,N_15134,N_15542);
nand U15831 (N_15831,N_15386,N_12595);
xnor U15832 (N_15832,N_13570,N_12579);
and U15833 (N_15833,N_12695,N_13607);
and U15834 (N_15834,N_14236,N_13216);
and U15835 (N_15835,N_14573,N_14445);
or U15836 (N_15836,N_14816,N_14118);
or U15837 (N_15837,N_15237,N_14977);
and U15838 (N_15838,N_14920,N_14781);
or U15839 (N_15839,N_13184,N_14074);
and U15840 (N_15840,N_13525,N_13610);
nand U15841 (N_15841,N_12567,N_14105);
and U15842 (N_15842,N_14145,N_14835);
and U15843 (N_15843,N_13124,N_14390);
and U15844 (N_15844,N_15481,N_14611);
nand U15845 (N_15845,N_14414,N_12996);
nand U15846 (N_15846,N_14697,N_15548);
nor U15847 (N_15847,N_13044,N_13528);
nand U15848 (N_15848,N_14958,N_13426);
or U15849 (N_15849,N_15075,N_13353);
nor U15850 (N_15850,N_12689,N_12999);
or U15851 (N_15851,N_15031,N_13234);
or U15852 (N_15852,N_14839,N_13660);
nand U15853 (N_15853,N_14514,N_15138);
or U15854 (N_15854,N_14643,N_12578);
or U15855 (N_15855,N_14680,N_13022);
or U15856 (N_15856,N_13306,N_12613);
and U15857 (N_15857,N_15345,N_13765);
nand U15858 (N_15858,N_12716,N_13167);
and U15859 (N_15859,N_12964,N_13879);
and U15860 (N_15860,N_15365,N_14130);
and U15861 (N_15861,N_13658,N_13709);
nand U15862 (N_15862,N_14042,N_13038);
nand U15863 (N_15863,N_15245,N_13348);
xnor U15864 (N_15864,N_15303,N_13142);
or U15865 (N_15865,N_14307,N_13035);
nor U15866 (N_15866,N_13591,N_13484);
and U15867 (N_15867,N_14968,N_12534);
nand U15868 (N_15868,N_15258,N_14729);
or U15869 (N_15869,N_14677,N_14538);
or U15870 (N_15870,N_13120,N_14271);
or U15871 (N_15871,N_15059,N_15498);
and U15872 (N_15872,N_12801,N_13079);
and U15873 (N_15873,N_15461,N_12785);
and U15874 (N_15874,N_15163,N_14998);
nor U15875 (N_15875,N_13109,N_14411);
nor U15876 (N_15876,N_15305,N_13412);
nor U15877 (N_15877,N_13223,N_14838);
xor U15878 (N_15878,N_15424,N_15170);
and U15879 (N_15879,N_15242,N_15558);
or U15880 (N_15880,N_15460,N_14793);
or U15881 (N_15881,N_12761,N_13582);
and U15882 (N_15882,N_13392,N_14248);
xor U15883 (N_15883,N_14454,N_13976);
and U15884 (N_15884,N_13533,N_15427);
or U15885 (N_15885,N_15593,N_14952);
and U15886 (N_15886,N_13600,N_13937);
or U15887 (N_15887,N_14882,N_13209);
and U15888 (N_15888,N_12963,N_14795);
and U15889 (N_15889,N_14027,N_13006);
xnor U15890 (N_15890,N_14324,N_15039);
xor U15891 (N_15891,N_14308,N_13344);
nand U15892 (N_15892,N_14992,N_14819);
xnor U15893 (N_15893,N_14593,N_12532);
nor U15894 (N_15894,N_15340,N_14871);
nand U15895 (N_15895,N_15056,N_14178);
and U15896 (N_15896,N_14082,N_15140);
nand U15897 (N_15897,N_14859,N_14482);
xor U15898 (N_15898,N_13416,N_15444);
or U15899 (N_15899,N_15246,N_14971);
xnor U15900 (N_15900,N_14148,N_12862);
nand U15901 (N_15901,N_15332,N_13979);
nand U15902 (N_15902,N_15588,N_14331);
nand U15903 (N_15903,N_13086,N_14306);
nor U15904 (N_15904,N_14908,N_14522);
or U15905 (N_15905,N_13875,N_14885);
nand U15906 (N_15906,N_12635,N_13073);
nor U15907 (N_15907,N_15168,N_15208);
xnor U15908 (N_15908,N_14263,N_13824);
xnor U15909 (N_15909,N_13102,N_12557);
nor U15910 (N_15910,N_14929,N_13843);
or U15911 (N_15911,N_13701,N_14318);
nor U15912 (N_15912,N_13299,N_14055);
or U15913 (N_15913,N_13823,N_14481);
xnor U15914 (N_15914,N_12634,N_13496);
and U15915 (N_15915,N_12528,N_13136);
nor U15916 (N_15916,N_14139,N_15122);
nor U15917 (N_15917,N_14759,N_13670);
nand U15918 (N_15918,N_13625,N_15544);
nor U15919 (N_15919,N_12509,N_13973);
nand U15920 (N_15920,N_12675,N_13764);
or U15921 (N_15921,N_13562,N_13957);
nand U15922 (N_15922,N_14058,N_15295);
nor U15923 (N_15923,N_15292,N_14474);
xor U15924 (N_15924,N_14628,N_15146);
xnor U15925 (N_15925,N_15348,N_15298);
or U15926 (N_15926,N_12932,N_13932);
or U15927 (N_15927,N_13931,N_14407);
or U15928 (N_15928,N_13329,N_15395);
or U15929 (N_15929,N_13827,N_15319);
xnor U15930 (N_15930,N_14924,N_15289);
or U15931 (N_15931,N_14737,N_13401);
or U15932 (N_15932,N_13631,N_13217);
or U15933 (N_15933,N_15323,N_14475);
nor U15934 (N_15934,N_14327,N_13514);
nand U15935 (N_15935,N_12592,N_14218);
or U15936 (N_15936,N_15186,N_12518);
and U15937 (N_15937,N_12919,N_13753);
xor U15938 (N_15938,N_13004,N_14498);
nand U15939 (N_15939,N_15280,N_13322);
nand U15940 (N_15940,N_13595,N_13841);
nand U15941 (N_15941,N_13104,N_14769);
nor U15942 (N_15942,N_14274,N_14903);
nor U15943 (N_15943,N_15118,N_14686);
xnor U15944 (N_15944,N_12993,N_13847);
xnor U15945 (N_15945,N_13812,N_13748);
or U15946 (N_15946,N_15421,N_12558);
nor U15947 (N_15947,N_15597,N_14003);
or U15948 (N_15948,N_14987,N_14736);
nand U15949 (N_15949,N_13839,N_14364);
xnor U15950 (N_15950,N_14800,N_14599);
nand U15951 (N_15951,N_14473,N_13368);
and U15952 (N_15952,N_15244,N_15213);
or U15953 (N_15953,N_14661,N_13901);
xnor U15954 (N_15954,N_15197,N_13198);
xor U15955 (N_15955,N_13723,N_14710);
nor U15956 (N_15956,N_15480,N_14537);
or U15957 (N_15957,N_13080,N_14917);
xor U15958 (N_15958,N_13776,N_14930);
nor U15959 (N_15959,N_12618,N_14630);
nor U15960 (N_15960,N_12563,N_15351);
nor U15961 (N_15961,N_15477,N_15220);
nor U15962 (N_15962,N_15261,N_14243);
and U15963 (N_15963,N_12840,N_12608);
nor U15964 (N_15964,N_13523,N_13059);
nor U15965 (N_15965,N_12736,N_13675);
nand U15966 (N_15966,N_13536,N_13309);
xnor U15967 (N_15967,N_15338,N_12979);
or U15968 (N_15968,N_13350,N_13226);
or U15969 (N_15969,N_14699,N_15600);
and U15970 (N_15970,N_15448,N_12520);
xnor U15971 (N_15971,N_14604,N_13430);
nand U15972 (N_15972,N_14476,N_13626);
and U15973 (N_15973,N_13147,N_13994);
xnor U15974 (N_15974,N_13001,N_13779);
xor U15975 (N_15975,N_14811,N_14725);
xor U15976 (N_15976,N_14730,N_13805);
or U15977 (N_15977,N_14406,N_12741);
nor U15978 (N_15978,N_15020,N_12904);
or U15979 (N_15979,N_14276,N_15306);
or U15980 (N_15980,N_13276,N_14856);
xnor U15981 (N_15981,N_14333,N_13270);
nand U15982 (N_15982,N_12719,N_15191);
nor U15983 (N_15983,N_12572,N_14135);
xor U15984 (N_15984,N_14765,N_13062);
xnor U15985 (N_15985,N_15489,N_15225);
nand U15986 (N_15986,N_13832,N_12867);
nand U15987 (N_15987,N_14095,N_14613);
nand U15988 (N_15988,N_13618,N_14873);
nand U15989 (N_15989,N_14054,N_13172);
or U15990 (N_15990,N_12853,N_12533);
nor U15991 (N_15991,N_12599,N_14501);
and U15992 (N_15992,N_13361,N_14366);
or U15993 (N_15993,N_14480,N_14855);
nor U15994 (N_15994,N_13050,N_14146);
nor U15995 (N_15995,N_15508,N_13587);
nand U15996 (N_15996,N_12681,N_15182);
nand U15997 (N_15997,N_13235,N_14815);
nand U15998 (N_15998,N_12927,N_15099);
and U15999 (N_15999,N_13636,N_12986);
nor U16000 (N_16000,N_12980,N_13712);
xor U16001 (N_16001,N_13461,N_15491);
or U16002 (N_16002,N_15007,N_13740);
and U16003 (N_16003,N_15497,N_14297);
nand U16004 (N_16004,N_14075,N_15178);
xnor U16005 (N_16005,N_15511,N_13688);
nor U16006 (N_16006,N_14959,N_13578);
or U16007 (N_16007,N_13614,N_14099);
nor U16008 (N_16008,N_15296,N_13787);
nand U16009 (N_16009,N_14261,N_13819);
xor U16010 (N_16010,N_13481,N_14720);
and U16011 (N_16011,N_12955,N_15083);
nor U16012 (N_16012,N_13325,N_13972);
xor U16013 (N_16013,N_14918,N_14159);
xnor U16014 (N_16014,N_15613,N_12577);
and U16015 (N_16015,N_14382,N_14957);
nand U16016 (N_16016,N_12938,N_14581);
or U16017 (N_16017,N_15443,N_13947);
nand U16018 (N_16018,N_12662,N_13594);
nand U16019 (N_16019,N_15496,N_13105);
nand U16020 (N_16020,N_14747,N_13987);
or U16021 (N_16021,N_15249,N_12540);
xnor U16022 (N_16022,N_13314,N_12729);
nor U16023 (N_16023,N_12603,N_15476);
xor U16024 (N_16024,N_14496,N_13047);
xor U16025 (N_16025,N_14771,N_14185);
and U16026 (N_16026,N_14463,N_13898);
nand U16027 (N_16027,N_12680,N_12795);
xor U16028 (N_16028,N_12583,N_15131);
nor U16029 (N_16029,N_15392,N_15451);
and U16030 (N_16030,N_14794,N_13185);
or U16031 (N_16031,N_12594,N_12949);
xnor U16032 (N_16032,N_14688,N_13777);
or U16033 (N_16033,N_13860,N_13786);
nor U16034 (N_16034,N_14809,N_14352);
xnor U16035 (N_16035,N_13680,N_14634);
and U16036 (N_16036,N_13682,N_15622);
xnor U16037 (N_16037,N_14767,N_15574);
nor U16038 (N_16038,N_13820,N_15576);
nor U16039 (N_16039,N_14638,N_15546);
and U16040 (N_16040,N_13449,N_15504);
nor U16041 (N_16041,N_12845,N_15226);
nor U16042 (N_16042,N_15315,N_15473);
xnor U16043 (N_16043,N_12682,N_14011);
nor U16044 (N_16044,N_14461,N_14889);
and U16045 (N_16045,N_13290,N_12972);
and U16046 (N_16046,N_13891,N_12749);
xnor U16047 (N_16047,N_13708,N_13140);
or U16048 (N_16048,N_14441,N_12930);
xor U16049 (N_16049,N_13720,N_13117);
and U16050 (N_16050,N_15591,N_15116);
nor U16051 (N_16051,N_12529,N_13347);
nand U16052 (N_16052,N_14951,N_13794);
and U16053 (N_16053,N_13518,N_13577);
nand U16054 (N_16054,N_14131,N_14629);
nor U16055 (N_16055,N_12580,N_12722);
nor U16056 (N_16056,N_13943,N_15057);
or U16057 (N_16057,N_12933,N_13095);
xnor U16058 (N_16058,N_15328,N_12571);
and U16059 (N_16059,N_14740,N_13981);
xor U16060 (N_16060,N_12826,N_15187);
nand U16061 (N_16061,N_13138,N_12747);
xor U16062 (N_16062,N_15228,N_13261);
and U16063 (N_16063,N_14438,N_14520);
xor U16064 (N_16064,N_14316,N_15347);
and U16065 (N_16065,N_13806,N_15470);
nor U16066 (N_16066,N_14486,N_14814);
or U16067 (N_16067,N_14883,N_15177);
xnor U16068 (N_16068,N_14207,N_15474);
or U16069 (N_16069,N_12956,N_14400);
xor U16070 (N_16070,N_13593,N_14353);
and U16071 (N_16071,N_13667,N_14374);
or U16072 (N_16072,N_14244,N_15114);
and U16073 (N_16073,N_13257,N_12706);
or U16074 (N_16074,N_13154,N_14554);
nor U16075 (N_16075,N_13153,N_15091);
and U16076 (N_16076,N_12512,N_14860);
or U16077 (N_16077,N_14468,N_14345);
or U16078 (N_16078,N_13985,N_15010);
nor U16079 (N_16079,N_14937,N_14963);
nand U16080 (N_16080,N_15535,N_12970);
and U16081 (N_16081,N_14967,N_12586);
and U16082 (N_16082,N_14682,N_14653);
xor U16083 (N_16083,N_13238,N_12946);
nor U16084 (N_16084,N_15123,N_15176);
nand U16085 (N_16085,N_15026,N_14077);
or U16086 (N_16086,N_14283,N_14953);
nor U16087 (N_16087,N_13913,N_14822);
and U16088 (N_16088,N_14427,N_15155);
and U16089 (N_16089,N_14431,N_12708);
or U16090 (N_16090,N_14852,N_13465);
nor U16091 (N_16091,N_14960,N_14745);
nand U16092 (N_16092,N_15367,N_14041);
or U16093 (N_16093,N_14096,N_13872);
nand U16094 (N_16094,N_14000,N_13017);
xnor U16095 (N_16095,N_14659,N_14657);
or U16096 (N_16096,N_15516,N_12649);
nor U16097 (N_16097,N_12982,N_12755);
or U16098 (N_16098,N_12648,N_14051);
nor U16099 (N_16099,N_15297,N_13650);
or U16100 (N_16100,N_13228,N_13321);
xor U16101 (N_16101,N_13043,N_15321);
xor U16102 (N_16102,N_13160,N_13666);
xnor U16103 (N_16103,N_14086,N_15314);
nand U16104 (N_16104,N_15500,N_14107);
nand U16105 (N_16105,N_13572,N_14862);
nand U16106 (N_16106,N_15530,N_13113);
nor U16107 (N_16107,N_12878,N_14497);
and U16108 (N_16108,N_15194,N_13569);
xnor U16109 (N_16109,N_14512,N_14751);
and U16110 (N_16110,N_13091,N_15353);
nand U16111 (N_16111,N_12638,N_13657);
nor U16112 (N_16112,N_14648,N_13686);
xnor U16113 (N_16113,N_15272,N_14637);
and U16114 (N_16114,N_13046,N_13566);
xnor U16115 (N_16115,N_14156,N_13679);
nand U16116 (N_16116,N_15370,N_15011);
or U16117 (N_16117,N_12652,N_12902);
xnor U16118 (N_16118,N_12576,N_13474);
xor U16119 (N_16119,N_12656,N_13747);
or U16120 (N_16120,N_12760,N_13240);
nor U16121 (N_16121,N_13190,N_13277);
xor U16122 (N_16122,N_14764,N_14351);
nor U16123 (N_16123,N_13958,N_14715);
or U16124 (N_16124,N_13203,N_13087);
nand U16125 (N_16125,N_13656,N_13563);
and U16126 (N_16126,N_15121,N_14339);
nor U16127 (N_16127,N_14645,N_12905);
nor U16128 (N_16128,N_14588,N_15419);
and U16129 (N_16129,N_13830,N_13940);
xnor U16130 (N_16130,N_14252,N_12666);
nor U16131 (N_16131,N_14545,N_15580);
and U16132 (N_16132,N_13211,N_13882);
nand U16133 (N_16133,N_13538,N_14803);
xor U16134 (N_16134,N_14235,N_12596);
and U16135 (N_16135,N_13333,N_13231);
xnor U16136 (N_16136,N_12690,N_13997);
nor U16137 (N_16137,N_14830,N_14045);
nand U16138 (N_16138,N_14451,N_14064);
nor U16139 (N_16139,N_15256,N_13041);
and U16140 (N_16140,N_13274,N_12775);
nor U16141 (N_16141,N_13310,N_14052);
or U16142 (N_16142,N_12759,N_13519);
nand U16143 (N_16143,N_15567,N_12590);
nor U16144 (N_16144,N_14119,N_14673);
xor U16145 (N_16145,N_14175,N_12547);
and U16146 (N_16146,N_13307,N_12684);
nand U16147 (N_16147,N_14442,N_13419);
nand U16148 (N_16148,N_12744,N_13025);
and U16149 (N_16149,N_14386,N_12786);
xor U16150 (N_16150,N_15202,N_14750);
and U16151 (N_16151,N_13254,N_14355);
nor U16152 (N_16152,N_12808,N_14290);
xnor U16153 (N_16153,N_14241,N_14829);
xor U16154 (N_16154,N_14721,N_14311);
nand U16155 (N_16155,N_14874,N_13420);
nand U16156 (N_16156,N_12812,N_14849);
nand U16157 (N_16157,N_14928,N_14965);
nor U16158 (N_16158,N_14544,N_12872);
nor U16159 (N_16159,N_15084,N_14568);
nor U16160 (N_16160,N_13557,N_14288);
or U16161 (N_16161,N_14741,N_14211);
nand U16162 (N_16162,N_14065,N_13766);
nand U16163 (N_16163,N_14626,N_14748);
or U16164 (N_16164,N_13888,N_15040);
nor U16165 (N_16165,N_14358,N_15012);
xor U16166 (N_16166,N_13908,N_14338);
or U16167 (N_16167,N_15531,N_12721);
and U16168 (N_16168,N_13571,N_12630);
and U16169 (N_16169,N_13964,N_13724);
nand U16170 (N_16170,N_12866,N_14770);
xnor U16171 (N_16171,N_13106,N_14777);
nor U16172 (N_16172,N_12822,N_14583);
xor U16173 (N_16173,N_14517,N_13030);
or U16174 (N_16174,N_15488,N_12617);
or U16175 (N_16175,N_13744,N_12790);
nor U16176 (N_16176,N_14255,N_13398);
nand U16177 (N_16177,N_15310,N_14222);
and U16178 (N_16178,N_14652,N_12626);
nand U16179 (N_16179,N_15438,N_12699);
nand U16180 (N_16180,N_12903,N_13822);
nor U16181 (N_16181,N_13866,N_12765);
nor U16182 (N_16182,N_13400,N_13033);
and U16183 (N_16183,N_12778,N_15215);
nor U16184 (N_16184,N_12602,N_14505);
and U16185 (N_16185,N_14214,N_13691);
xnor U16186 (N_16186,N_14247,N_14878);
xor U16187 (N_16187,N_15522,N_14194);
nor U16188 (N_16188,N_12816,N_14787);
or U16189 (N_16189,N_12647,N_13447);
xnor U16190 (N_16190,N_13852,N_14017);
xnor U16191 (N_16191,N_14357,N_13145);
or U16192 (N_16192,N_14681,N_13337);
or U16193 (N_16193,N_14596,N_13164);
or U16194 (N_16194,N_13520,N_14253);
or U16195 (N_16195,N_14238,N_14436);
nand U16196 (N_16196,N_12895,N_15283);
nand U16197 (N_16197,N_13424,N_14469);
or U16198 (N_16198,N_13818,N_14887);
and U16199 (N_16199,N_13369,N_13341);
xor U16200 (N_16200,N_13372,N_13249);
and U16201 (N_16201,N_13791,N_13564);
or U16202 (N_16202,N_14016,N_13283);
nand U16203 (N_16203,N_15098,N_14397);
nand U16204 (N_16204,N_13521,N_12884);
nand U16205 (N_16205,N_14365,N_14614);
nor U16206 (N_16206,N_12710,N_14724);
and U16207 (N_16207,N_14633,N_13717);
nor U16208 (N_16208,N_15184,N_15466);
or U16209 (N_16209,N_13986,N_14948);
and U16210 (N_16210,N_13619,N_13082);
xnor U16211 (N_16211,N_14927,N_14162);
and U16212 (N_16212,N_12942,N_13093);
and U16213 (N_16213,N_15117,N_12995);
nor U16214 (N_16214,N_14179,N_15224);
or U16215 (N_16215,N_14651,N_13735);
or U16216 (N_16216,N_14420,N_13808);
nor U16217 (N_16217,N_14384,N_12733);
xnor U16218 (N_16218,N_15357,N_14116);
nor U16219 (N_16219,N_13601,N_14752);
nor U16220 (N_16220,N_12819,N_13354);
and U16221 (N_16221,N_12960,N_15577);
and U16222 (N_16222,N_13725,N_13230);
and U16223 (N_16223,N_13945,N_14618);
nor U16224 (N_16224,N_14379,N_13224);
and U16225 (N_16225,N_12654,N_14076);
nor U16226 (N_16226,N_13980,N_12931);
nand U16227 (N_16227,N_12504,N_14021);
nand U16228 (N_16228,N_13936,N_14089);
xor U16229 (N_16229,N_14007,N_15044);
xor U16230 (N_16230,N_14768,N_15425);
nand U16231 (N_16231,N_15078,N_12731);
or U16232 (N_16232,N_14706,N_15190);
or U16233 (N_16233,N_12772,N_15050);
and U16234 (N_16234,N_15534,N_14602);
nand U16235 (N_16235,N_12606,N_15612);
nand U16236 (N_16236,N_14578,N_14361);
and U16237 (N_16237,N_14556,N_15259);
or U16238 (N_16238,N_13641,N_14704);
or U16239 (N_16239,N_13928,N_13191);
or U16240 (N_16240,N_13359,N_14539);
or U16241 (N_16241,N_12985,N_12544);
nor U16242 (N_16242,N_13598,N_13550);
xor U16243 (N_16243,N_13624,N_14687);
and U16244 (N_16244,N_15107,N_15200);
xor U16245 (N_16245,N_12870,N_13559);
nor U16246 (N_16246,N_14574,N_15525);
nor U16247 (N_16247,N_15594,N_14693);
or U16248 (N_16248,N_14932,N_15437);
nand U16249 (N_16249,N_14217,N_14806);
nand U16250 (N_16250,N_13444,N_14779);
xor U16251 (N_16251,N_14650,N_15192);
and U16252 (N_16252,N_13482,N_14152);
nor U16253 (N_16253,N_14026,N_13532);
nand U16254 (N_16254,N_12517,N_15037);
and U16255 (N_16255,N_15616,N_13946);
or U16256 (N_16256,N_15447,N_14395);
xnor U16257 (N_16257,N_15210,N_13721);
nand U16258 (N_16258,N_15543,N_14956);
or U16259 (N_16259,N_13402,N_15181);
or U16260 (N_16260,N_15405,N_13237);
nand U16261 (N_16261,N_13829,N_13436);
or U16262 (N_16262,N_13464,N_13929);
nor U16263 (N_16263,N_15563,N_13364);
nor U16264 (N_16264,N_13479,N_12890);
nor U16265 (N_16265,N_13092,N_14079);
nor U16266 (N_16266,N_12735,N_15189);
nor U16267 (N_16267,N_14109,N_14341);
and U16268 (N_16268,N_14674,N_15453);
or U16269 (N_16269,N_15456,N_13923);
nor U16270 (N_16270,N_13456,N_15312);
and U16271 (N_16271,N_12730,N_13966);
xor U16272 (N_16272,N_13739,N_12727);
and U16273 (N_16273,N_12624,N_14902);
nand U16274 (N_16274,N_13726,N_12555);
or U16275 (N_16275,N_14595,N_12537);
or U16276 (N_16276,N_13560,N_13751);
xor U16277 (N_16277,N_13885,N_15266);
xor U16278 (N_16278,N_12636,N_14898);
nor U16279 (N_16279,N_14388,N_12857);
and U16280 (N_16280,N_13516,N_13094);
and U16281 (N_16281,N_13907,N_14550);
xor U16282 (N_16282,N_13652,N_15510);
nor U16283 (N_16283,N_13716,N_14378);
nand U16284 (N_16284,N_15100,N_13371);
nand U16285 (N_16285,N_14553,N_14413);
and U16286 (N_16286,N_15301,N_13455);
nor U16287 (N_16287,N_15120,N_15212);
and U16288 (N_16288,N_13534,N_15617);
nand U16289 (N_16289,N_13027,N_14424);
xnor U16290 (N_16290,N_12850,N_13115);
or U16291 (N_16291,N_13366,N_15552);
nor U16292 (N_16292,N_12791,N_13788);
nand U16293 (N_16293,N_15093,N_14090);
or U16294 (N_16294,N_14063,N_14376);
nand U16295 (N_16295,N_13074,N_13640);
xor U16296 (N_16296,N_12678,N_15462);
nand U16297 (N_16297,N_15339,N_14876);
or U16298 (N_16298,N_14962,N_13055);
or U16299 (N_16299,N_13475,N_12915);
nor U16300 (N_16300,N_13639,N_14408);
xnor U16301 (N_16301,N_13857,N_15478);
and U16302 (N_16302,N_13175,N_13834);
xor U16303 (N_16303,N_12798,N_13158);
nor U16304 (N_16304,N_12825,N_12876);
nand U16305 (N_16305,N_15368,N_13067);
xnor U16306 (N_16306,N_15449,N_13849);
nor U16307 (N_16307,N_14073,N_14813);
nand U16308 (N_16308,N_15429,N_14587);
and U16309 (N_16309,N_15198,N_12898);
or U16310 (N_16310,N_14487,N_13642);
xnor U16311 (N_16311,N_13263,N_14230);
xnor U16312 (N_16312,N_13797,N_14342);
xnor U16313 (N_16313,N_14049,N_13643);
nand U16314 (N_16314,N_14133,N_14826);
xor U16315 (N_16315,N_14735,N_13647);
nand U16316 (N_16316,N_14205,N_13362);
xnor U16317 (N_16317,N_13210,N_13311);
or U16318 (N_16318,N_12951,N_13406);
xor U16319 (N_16319,N_13509,N_13328);
nor U16320 (N_16320,N_14362,N_14210);
xor U16321 (N_16321,N_15326,N_15529);
or U16322 (N_16322,N_12502,N_13500);
nor U16323 (N_16323,N_14190,N_14892);
nor U16324 (N_16324,N_14761,N_13243);
nand U16325 (N_16325,N_14600,N_13749);
xor U16326 (N_16326,N_14609,N_14734);
nand U16327 (N_16327,N_14203,N_15564);
and U16328 (N_16328,N_13495,N_15293);
and U16329 (N_16329,N_12820,N_13285);
nor U16330 (N_16330,N_13305,N_15061);
or U16331 (N_16331,N_13065,N_15551);
and U16332 (N_16332,N_14667,N_13902);
or U16333 (N_16333,N_15164,N_15407);
xnor U16334 (N_16334,N_15144,N_12789);
nor U16335 (N_16335,N_14733,N_13645);
and U16336 (N_16336,N_13139,N_14066);
nand U16337 (N_16337,N_14774,N_14836);
and U16338 (N_16338,N_14531,N_13878);
and U16339 (N_16339,N_14032,N_14996);
xor U16340 (N_16340,N_15559,N_12792);
or U16341 (N_16341,N_13417,N_13195);
or U16342 (N_16342,N_13774,N_14723);
nor U16343 (N_16343,N_13034,N_13837);
xnor U16344 (N_16344,N_14312,N_14282);
and U16345 (N_16345,N_14558,N_13382);
xnor U16346 (N_16346,N_15260,N_12692);
xor U16347 (N_16347,N_13971,N_13324);
and U16348 (N_16348,N_13590,N_13941);
xnor U16349 (N_16349,N_14383,N_13540);
or U16350 (N_16350,N_12625,N_14206);
nand U16351 (N_16351,N_14121,N_15033);
and U16352 (N_16352,N_14784,N_13403);
or U16353 (N_16353,N_15358,N_13280);
and U16354 (N_16354,N_14631,N_14535);
xor U16355 (N_16355,N_13673,N_14646);
or U16356 (N_16356,N_13543,N_12641);
xor U16357 (N_16357,N_12683,N_15105);
or U16358 (N_16358,N_14907,N_12839);
or U16359 (N_16359,N_14961,N_13227);
nand U16360 (N_16360,N_13083,N_15507);
xnor U16361 (N_16361,N_13815,N_13317);
xor U16362 (N_16362,N_13298,N_15262);
nand U16363 (N_16363,N_15290,N_12861);
nor U16364 (N_16364,N_13895,N_12856);
xor U16365 (N_16365,N_12950,N_14373);
or U16366 (N_16366,N_12793,N_15027);
nand U16367 (N_16367,N_13678,N_13360);
xor U16368 (N_16368,N_14009,N_14880);
and U16369 (N_16369,N_13487,N_14934);
nor U16370 (N_16370,N_15207,N_13103);
xor U16371 (N_16371,N_15060,N_15051);
and U16372 (N_16372,N_12965,N_14272);
and U16373 (N_16373,N_13020,N_12834);
or U16374 (N_16374,N_13483,N_13151);
xor U16375 (N_16375,N_13301,N_12854);
nor U16376 (N_16376,N_12570,N_13905);
xnor U16377 (N_16377,N_15584,N_13011);
or U16378 (N_16378,N_15375,N_12587);
nand U16379 (N_16379,N_14547,N_13457);
and U16380 (N_16380,N_15414,N_13912);
or U16381 (N_16381,N_15103,N_12978);
nor U16382 (N_16382,N_13873,N_12851);
xnor U16383 (N_16383,N_12899,N_13674);
nand U16384 (N_16384,N_15204,N_14310);
nor U16385 (N_16385,N_15043,N_13880);
nand U16386 (N_16386,N_14555,N_15049);
nor U16387 (N_16387,N_13476,N_14616);
xor U16388 (N_16388,N_14070,N_15607);
nor U16389 (N_16389,N_14493,N_13130);
nor U16390 (N_16390,N_12810,N_15505);
nand U16391 (N_16391,N_12957,N_13575);
nand U16392 (N_16392,N_14220,N_14264);
xnor U16393 (N_16393,N_13991,N_13377);
nand U16394 (N_16394,N_14403,N_14412);
or U16395 (N_16395,N_14091,N_13029);
nor U16396 (N_16396,N_14502,N_14756);
nand U16397 (N_16397,N_13664,N_13225);
or U16398 (N_16398,N_15175,N_14844);
nand U16399 (N_16399,N_15334,N_14279);
or U16400 (N_16400,N_12542,N_14192);
nor U16401 (N_16401,N_13016,N_14824);
and U16402 (N_16402,N_12535,N_13921);
xnor U16403 (N_16403,N_14084,N_15452);
xnor U16404 (N_16404,N_13289,N_14025);
nand U16405 (N_16405,N_13974,N_14208);
and U16406 (N_16406,N_13396,N_14897);
nand U16407 (N_16407,N_13613,N_15066);
nor U16408 (N_16408,N_15263,N_15286);
and U16409 (N_16409,N_14845,N_15233);
and U16410 (N_16410,N_13999,N_13300);
xor U16411 (N_16411,N_15519,N_14866);
xnor U16412 (N_16412,N_14444,N_15152);
or U16413 (N_16413,N_12947,N_15016);
nand U16414 (N_16414,N_15528,N_15320);
nor U16415 (N_16415,N_15171,N_13732);
nor U16416 (N_16416,N_15377,N_12860);
and U16417 (N_16417,N_14043,N_13427);
and U16418 (N_16418,N_13345,N_14150);
xnor U16419 (N_16419,N_12574,N_12653);
nor U16420 (N_16420,N_14484,N_15605);
and U16421 (N_16421,N_15536,N_12622);
and U16422 (N_16422,N_14589,N_12846);
nor U16423 (N_16423,N_13869,N_12660);
and U16424 (N_16424,N_15413,N_15046);
and U16425 (N_16425,N_13545,N_14979);
nor U16426 (N_16426,N_13551,N_13303);
and U16427 (N_16427,N_13338,N_14048);
and U16428 (N_16428,N_15609,N_13850);
and U16429 (N_16429,N_13288,N_13616);
and U16430 (N_16430,N_14543,N_14295);
xor U16431 (N_16431,N_14817,N_14978);
and U16432 (N_16432,N_14335,N_13515);
or U16433 (N_16433,N_13128,N_15445);
nor U16434 (N_16434,N_13097,N_12550);
xnor U16435 (N_16435,N_13669,N_13390);
and U16436 (N_16436,N_12707,N_14046);
nor U16437 (N_16437,N_12700,N_13439);
and U16438 (N_16438,N_15111,N_14639);
nor U16439 (N_16439,N_14936,N_15148);
nand U16440 (N_16440,N_13466,N_14842);
nand U16441 (N_16441,N_13316,N_13446);
or U16442 (N_16442,N_14363,N_13924);
and U16443 (N_16443,N_15232,N_13052);
xnor U16444 (N_16444,N_13181,N_15408);
and U16445 (N_16445,N_12788,N_12629);
nor U16446 (N_16446,N_13554,N_15274);
nand U16447 (N_16447,N_14577,N_14701);
nor U16448 (N_16448,N_14196,N_15277);
nor U16449 (N_16449,N_15382,N_13876);
xor U16450 (N_16450,N_14722,N_14256);
or U16451 (N_16451,N_13114,N_15592);
and U16452 (N_16452,N_13699,N_14300);
nor U16453 (N_16453,N_15325,N_15402);
or U16454 (N_16454,N_13308,N_13537);
nand U16455 (N_16455,N_14100,N_12541);
and U16456 (N_16456,N_13218,N_13734);
nand U16457 (N_16457,N_14711,N_15130);
xor U16458 (N_16458,N_15082,N_12837);
nor U16459 (N_16459,N_13719,N_13894);
nand U16460 (N_16460,N_13770,N_15282);
xor U16461 (N_16461,N_13741,N_14488);
or U16462 (N_16462,N_13486,N_13696);
or U16463 (N_16463,N_13862,N_13763);
nor U16464 (N_16464,N_14755,N_15154);
nor U16465 (N_16465,N_12813,N_15426);
xnor U16466 (N_16466,N_15471,N_15052);
nand U16467 (N_16467,N_14399,N_13428);
xnor U16468 (N_16468,N_13918,N_15136);
nor U16469 (N_16469,N_12916,N_15125);
nand U16470 (N_16470,N_15313,N_12925);
and U16471 (N_16471,N_13555,N_14564);
nand U16472 (N_16472,N_15537,N_15411);
nand U16473 (N_16473,N_12859,N_14586);
and U16474 (N_16474,N_13318,N_13653);
nor U16475 (N_16475,N_14801,N_14526);
and U16476 (N_16476,N_14158,N_14069);
nor U16477 (N_16477,N_14921,N_14919);
nor U16478 (N_16478,N_14775,N_15404);
xor U16479 (N_16479,N_13793,N_14656);
nor U16480 (N_16480,N_15141,N_13326);
nor U16481 (N_16481,N_12969,N_14981);
or U16482 (N_16482,N_14763,N_15062);
and U16483 (N_16483,N_14277,N_15578);
nand U16484 (N_16484,N_14062,N_15479);
nor U16485 (N_16485,N_14251,N_13634);
nand U16486 (N_16486,N_14990,N_15513);
xnor U16487 (N_16487,N_14792,N_15406);
nand U16488 (N_16488,N_13178,N_15374);
or U16489 (N_16489,N_14865,N_12771);
nand U16490 (N_16490,N_12843,N_14030);
and U16491 (N_16491,N_15112,N_13809);
xnor U16492 (N_16492,N_14847,N_12714);
nand U16493 (N_16493,N_13488,N_14056);
xnor U16494 (N_16494,N_13222,N_13246);
xnor U16495 (N_16495,N_14293,N_12545);
nor U16496 (N_16496,N_14422,N_13177);
xnor U16497 (N_16497,N_13255,N_15430);
xnor U16498 (N_16498,N_12748,N_15350);
or U16499 (N_16499,N_14891,N_12516);
nor U16500 (N_16500,N_15316,N_14394);
xor U16501 (N_16501,N_14460,N_13759);
nand U16502 (N_16502,N_13836,N_15250);
nand U16503 (N_16503,N_14612,N_13864);
and U16504 (N_16504,N_13205,N_13355);
and U16505 (N_16505,N_12934,N_12514);
nand U16506 (N_16506,N_15054,N_15434);
or U16507 (N_16507,N_12796,N_13897);
or U16508 (N_16508,N_14738,N_14249);
nand U16509 (N_16509,N_13271,N_14585);
and U16510 (N_16510,N_14623,N_13995);
or U16511 (N_16511,N_13000,N_14142);
or U16512 (N_16512,N_14226,N_12696);
xnor U16513 (N_16513,N_14184,N_15166);
nor U16514 (N_16514,N_15341,N_12685);
or U16515 (N_16515,N_15527,N_14541);
or U16516 (N_16516,N_13024,N_12780);
or U16517 (N_16517,N_15308,N_12835);
xnor U16518 (N_16518,N_14040,N_14012);
xnor U16519 (N_16519,N_12661,N_13295);
or U16520 (N_16520,N_12891,N_13253);
or U16521 (N_16521,N_14097,N_14088);
or U16522 (N_16522,N_12943,N_13458);
nor U16523 (N_16523,N_13851,N_12869);
nand U16524 (N_16524,N_13526,N_13710);
nor U16525 (N_16525,N_13409,N_14129);
nand U16526 (N_16526,N_15024,N_12794);
or U16527 (N_16527,N_14695,N_13605);
nand U16528 (N_16528,N_15299,N_13968);
xnor U16529 (N_16529,N_14120,N_14309);
nor U16530 (N_16530,N_12975,N_13009);
nor U16531 (N_16531,N_14843,N_14974);
nand U16532 (N_16532,N_12936,N_14136);
nor U16533 (N_16533,N_15441,N_12672);
nor U16534 (N_16534,N_13018,N_14067);
or U16535 (N_16535,N_13302,N_13760);
and U16536 (N_16536,N_12677,N_14215);
nand U16537 (N_16537,N_14381,N_13877);
nor U16538 (N_16538,N_13118,N_15520);
or U16539 (N_16539,N_12746,N_15569);
xor U16540 (N_16540,N_14521,N_13335);
xor U16541 (N_16541,N_12575,N_12561);
and U16542 (N_16542,N_14796,N_14432);
and U16543 (N_16543,N_13539,N_13199);
nor U16544 (N_16544,N_15304,N_12962);
nor U16545 (N_16545,N_15038,N_15361);
nor U16546 (N_16546,N_13861,N_13405);
and U16547 (N_16547,N_15018,N_12974);
nand U16548 (N_16548,N_12511,N_14947);
xor U16549 (N_16549,N_13269,N_14354);
or U16550 (N_16550,N_14286,N_13845);
or U16551 (N_16551,N_14246,N_14134);
nor U16552 (N_16552,N_13214,N_12720);
and U16553 (N_16553,N_14421,N_14579);
xor U16554 (N_16554,N_14821,N_13896);
xnor U16555 (N_16555,N_13599,N_12883);
xor U16556 (N_16556,N_14685,N_14780);
or U16557 (N_16557,N_14896,N_13955);
nor U16558 (N_16558,N_13068,N_13245);
or U16559 (N_16559,N_13914,N_14013);
xnor U16560 (N_16560,N_13817,N_15582);
xor U16561 (N_16561,N_14692,N_15174);
xnor U16562 (N_16562,N_14875,N_14605);
and U16563 (N_16563,N_13331,N_14524);
and U16564 (N_16564,N_12954,N_12873);
nor U16565 (N_16565,N_14518,N_14464);
xor U16566 (N_16566,N_14994,N_15364);
xor U16567 (N_16567,N_15396,N_14202);
xnor U16568 (N_16568,N_13425,N_13970);
xnor U16569 (N_16569,N_15022,N_13633);
nand U16570 (N_16570,N_14712,N_14812);
nor U16571 (N_16571,N_15017,N_13241);
xor U16572 (N_16572,N_15230,N_12565);
xor U16573 (N_16573,N_13268,N_13471);
xnor U16574 (N_16574,N_13292,N_15309);
xnor U16575 (N_16575,N_13854,N_15506);
nand U16576 (N_16576,N_13884,N_13592);
nor U16577 (N_16577,N_15359,N_12921);
xnor U16578 (N_16578,N_13906,N_15080);
nor U16579 (N_16579,N_15523,N_14410);
xor U16580 (N_16580,N_12598,N_14177);
nand U16581 (N_16581,N_14273,N_13143);
or U16582 (N_16582,N_14124,N_15586);
and U16583 (N_16583,N_12701,N_15069);
and U16584 (N_16584,N_15317,N_12724);
xnor U16585 (N_16585,N_15587,N_13694);
xnor U16586 (N_16586,N_13704,N_14182);
nand U16587 (N_16587,N_14944,N_14392);
nand U16588 (N_16588,N_13746,N_15029);
and U16589 (N_16589,N_13993,N_13013);
or U16590 (N_16590,N_12961,N_13282);
xnor U16591 (N_16591,N_13327,N_14627);
xnor U16592 (N_16592,N_14258,N_14534);
nor U16593 (N_16593,N_14527,N_13998);
nand U16594 (N_16594,N_15560,N_14169);
xor U16595 (N_16595,N_12640,N_12526);
xnor U16596 (N_16596,N_14008,N_13903);
or U16597 (N_16597,N_13443,N_13568);
nand U16598 (N_16598,N_14204,N_12552);
and U16599 (N_16599,N_14857,N_13262);
and U16600 (N_16600,N_13189,N_13435);
and U16601 (N_16601,N_14110,N_14625);
nor U16602 (N_16602,N_13790,N_14085);
nor U16603 (N_16603,N_15268,N_12732);
and U16604 (N_16604,N_13266,N_13433);
and U16605 (N_16605,N_14168,N_14731);
nor U16606 (N_16606,N_15081,N_14014);
nand U16607 (N_16607,N_14198,N_13489);
xor U16608 (N_16608,N_14840,N_15585);
nand U16609 (N_16609,N_13462,N_15070);
or U16610 (N_16610,N_12605,N_15173);
nand U16611 (N_16611,N_15549,N_15279);
xnor U16612 (N_16612,N_15021,N_13501);
or U16613 (N_16613,N_15265,N_15097);
nor U16614 (N_16614,N_15072,N_15389);
nor U16615 (N_16615,N_13411,N_13171);
or U16616 (N_16616,N_13942,N_12769);
or U16617 (N_16617,N_14360,N_13695);
or U16618 (N_16618,N_13983,N_12833);
nor U16619 (N_16619,N_12663,N_14754);
nand U16620 (N_16620,N_13058,N_13780);
nand U16621 (N_16621,N_13953,N_15079);
nor U16622 (N_16622,N_14709,N_15568);
nand U16623 (N_16623,N_14268,N_13407);
and U16624 (N_16624,N_14690,N_14034);
nor U16625 (N_16625,N_13693,N_14370);
xor U16626 (N_16626,N_14385,N_14292);
and U16627 (N_16627,N_14827,N_15482);
nor U16628 (N_16628,N_13320,N_13126);
xnor U16629 (N_16629,N_15240,N_14313);
nand U16630 (N_16630,N_12604,N_13840);
and U16631 (N_16631,N_14180,N_15398);
nor U16632 (N_16632,N_15539,N_12620);
nand U16633 (N_16633,N_14536,N_13323);
or U16634 (N_16634,N_14209,N_13910);
nand U16635 (N_16635,N_15110,N_15566);
nand U16636 (N_16636,N_13194,N_15620);
xor U16637 (N_16637,N_15442,N_13442);
or U16638 (N_16638,N_14991,N_14714);
or U16639 (N_16639,N_12510,N_14848);
or U16640 (N_16640,N_14879,N_13408);
nor U16641 (N_16641,N_14935,N_12937);
xor U16642 (N_16642,N_13168,N_12519);
and U16643 (N_16643,N_12738,N_12918);
or U16644 (N_16644,N_14233,N_13085);
or U16645 (N_16645,N_15495,N_14389);
nand U16646 (N_16646,N_15085,N_12582);
and U16647 (N_16647,N_14678,N_13252);
nand U16648 (N_16648,N_13975,N_15403);
nand U16649 (N_16649,N_13711,N_14684);
and U16650 (N_16650,N_13399,N_12619);
and U16651 (N_16651,N_13287,N_14456);
or U16652 (N_16652,N_12522,N_14515);
nor U16653 (N_16653,N_15180,N_15013);
and U16654 (N_16654,N_13395,N_13684);
and U16655 (N_16655,N_15387,N_13576);
or U16656 (N_16656,N_15515,N_14707);
and U16657 (N_16657,N_14696,N_14111);
nor U16658 (N_16658,N_14322,N_14997);
nor U16659 (N_16659,N_12935,N_13917);
nand U16660 (N_16660,N_14428,N_14805);
or U16661 (N_16661,N_13731,N_13831);
nand U16662 (N_16662,N_15621,N_14260);
and U16663 (N_16663,N_15158,N_13663);
and U16664 (N_16664,N_15216,N_14719);
nand U16665 (N_16665,N_14450,N_13506);
and U16666 (N_16666,N_14402,N_14655);
or U16667 (N_16667,N_13909,N_15532);
xor U16668 (N_16668,N_13798,N_12959);
nor U16669 (N_16669,N_14072,N_14466);
nor U16670 (N_16670,N_15436,N_12926);
and U16671 (N_16671,N_13304,N_12667);
nor U16672 (N_16672,N_14240,N_15596);
nand U16673 (N_16673,N_13622,N_15311);
nor U16674 (N_16674,N_15322,N_13567);
and U16675 (N_16675,N_15446,N_14820);
nand U16676 (N_16676,N_12907,N_15330);
and U16677 (N_16677,N_15378,N_13259);
nand U16678 (N_16678,N_14881,N_13293);
nor U16679 (N_16679,N_13714,N_15251);
nand U16680 (N_16680,N_15484,N_12655);
nor U16681 (N_16681,N_15422,N_12782);
nor U16682 (N_16682,N_15455,N_13935);
nor U16683 (N_16683,N_13278,N_14229);
xor U16684 (N_16684,N_14478,N_14160);
nor U16685 (N_16685,N_15391,N_13200);
xor U16686 (N_16686,N_13922,N_13247);
and U16687 (N_16687,N_13021,N_14485);
nand U16688 (N_16688,N_14546,N_14405);
xor U16689 (N_16689,N_14287,N_13697);
xor U16690 (N_16690,N_14157,N_13204);
or U16691 (N_16691,N_12952,N_13612);
nor U16692 (N_16692,N_14128,N_13467);
or U16693 (N_16693,N_14580,N_12836);
nor U16694 (N_16694,N_14223,N_15483);
nand U16695 (N_16695,N_15157,N_13119);
nand U16696 (N_16696,N_12911,N_14946);
xor U16697 (N_16697,N_15218,N_13296);
nand U16698 (N_16698,N_15199,N_14472);
nand U16699 (N_16699,N_14340,N_14635);
nor U16700 (N_16700,N_14529,N_13081);
xor U16701 (N_16701,N_12991,N_15235);
nor U16702 (N_16702,N_14941,N_14559);
or U16703 (N_16703,N_12823,N_15499);
nand U16704 (N_16704,N_12530,N_15417);
nor U16705 (N_16705,N_14019,N_14727);
or U16706 (N_16706,N_15550,N_13108);
and U16707 (N_16707,N_13132,N_12948);
nor U16708 (N_16708,N_15087,N_13911);
nand U16709 (N_16709,N_13040,N_12984);
nand U16710 (N_16710,N_12844,N_15463);
and U16711 (N_16711,N_12784,N_15324);
or U16712 (N_16712,N_12824,N_12990);
nor U16713 (N_16713,N_15231,N_13351);
or U16714 (N_16714,N_14094,N_13580);
nand U16715 (N_16715,N_14455,N_13459);
nor U16716 (N_16716,N_14265,N_14837);
nand U16717 (N_16717,N_15109,N_12809);
nand U16718 (N_16718,N_13982,N_12703);
xnor U16719 (N_16719,N_13549,N_15169);
nand U16720 (N_16720,N_12889,N_14654);
nand U16721 (N_16721,N_13632,N_13144);
nand U16722 (N_16722,N_12694,N_13221);
nor U16723 (N_16723,N_13422,N_15602);
nor U16724 (N_16724,N_12609,N_13313);
and U16725 (N_16725,N_15400,N_13996);
xnor U16726 (N_16726,N_15624,N_15337);
nand U16727 (N_16727,N_15409,N_15547);
nand U16728 (N_16728,N_13833,N_12503);
nand U16729 (N_16729,N_13448,N_13609);
or U16730 (N_16730,N_14647,N_15195);
nor U16731 (N_16731,N_13644,N_13502);
nand U16732 (N_16732,N_13814,N_15346);
nand U16733 (N_16733,N_15360,N_13434);
xor U16734 (N_16734,N_13131,N_14540);
nor U16735 (N_16735,N_15106,N_12539);
and U16736 (N_16736,N_12549,N_14068);
xor U16737 (N_16737,N_14254,N_13858);
and U16738 (N_16738,N_13608,N_13397);
nand U16739 (N_16739,N_13379,N_13629);
nor U16740 (N_16740,N_14886,N_13855);
or U16741 (N_16741,N_13556,N_15336);
and U16742 (N_16742,N_13676,N_15435);
xnor U16743 (N_16743,N_13008,N_12768);
nor U16744 (N_16744,N_13107,N_13100);
nand U16745 (N_16745,N_15185,N_13978);
or U16746 (N_16746,N_13340,N_14433);
nor U16747 (N_16747,N_13588,N_15514);
nor U16748 (N_16748,N_15390,N_14035);
xor U16749 (N_16749,N_14224,N_12777);
or U16750 (N_16750,N_13069,N_12756);
nand U16751 (N_16751,N_12723,N_14683);
nor U16752 (N_16752,N_12642,N_14108);
nor U16753 (N_16753,N_14500,N_13792);
or U16754 (N_16754,N_14525,N_13452);
nand U16755 (N_16755,N_14492,N_15132);
and U16756 (N_16756,N_14250,N_14749);
nor U16757 (N_16757,N_12665,N_12562);
nor U16758 (N_16758,N_12909,N_13188);
or U16759 (N_16759,N_14189,N_15318);
or U16760 (N_16760,N_13801,N_15067);
nor U16761 (N_16761,N_14314,N_13414);
nor U16762 (N_16762,N_14575,N_12908);
nand U16763 (N_16763,N_12966,N_13088);
or U16764 (N_16764,N_12621,N_13150);
nor U16765 (N_16765,N_14636,N_12740);
nor U16766 (N_16766,N_14083,N_13157);
nor U16767 (N_16767,N_12702,N_14900);
nand U16768 (N_16768,N_15139,N_13930);
nor U16769 (N_16769,N_13899,N_12506);
or U16770 (N_16770,N_14954,N_13163);
xor U16771 (N_16771,N_12527,N_13183);
or U16772 (N_16772,N_14242,N_14590);
and U16773 (N_16773,N_14582,N_14416);
and U16774 (N_16774,N_13491,N_15193);
xor U16775 (N_16775,N_12997,N_14336);
nand U16776 (N_16776,N_13573,N_13294);
and U16777 (N_16777,N_14964,N_13078);
nand U16778 (N_16778,N_13597,N_12584);
xor U16779 (N_16779,N_14347,N_14776);
and U16780 (N_16780,N_14037,N_14038);
nor U16781 (N_16781,N_13867,N_13497);
xnor U16782 (N_16782,N_14562,N_14841);
xnor U16783 (N_16783,N_13904,N_13825);
or U16784 (N_16784,N_15487,N_13418);
or U16785 (N_16785,N_13527,N_14906);
and U16786 (N_16786,N_14372,N_15331);
nand U16787 (N_16787,N_13202,N_13057);
and U16788 (N_16788,N_14671,N_13810);
nand U16789 (N_16789,N_12988,N_13123);
and U16790 (N_16790,N_13485,N_15475);
nand U16791 (N_16791,N_12628,N_13621);
nand U16792 (N_16792,N_12631,N_14147);
or U16793 (N_16793,N_13339,N_14679);
or U16794 (N_16794,N_13638,N_14057);
or U16795 (N_16795,N_12751,N_14199);
xor U16796 (N_16796,N_14938,N_12581);
and U16797 (N_16797,N_13651,N_15101);
and U16798 (N_16798,N_14798,N_14409);
nor U16799 (N_16799,N_14823,N_14140);
and U16800 (N_16800,N_14955,N_13071);
nand U16801 (N_16801,N_12877,N_14275);
or U16802 (N_16802,N_12847,N_15241);
nor U16803 (N_16803,N_14106,N_15102);
or U16804 (N_16804,N_13336,N_13156);
or U16805 (N_16805,N_14122,N_14901);
xor U16806 (N_16806,N_15418,N_13799);
or U16807 (N_16807,N_14893,N_14471);
or U16808 (N_16808,N_12543,N_13440);
nor U16809 (N_16809,N_15575,N_12894);
nor U16810 (N_16810,N_15222,N_13450);
nor U16811 (N_16811,N_13803,N_14328);
xnor U16812 (N_16812,N_14087,N_13503);
nand U16813 (N_16813,N_13005,N_14483);
or U16814 (N_16814,N_14081,N_15354);
and U16815 (N_16815,N_13811,N_13692);
nand U16816 (N_16816,N_14429,N_14491);
or U16817 (N_16817,N_14926,N_14603);
xor U16818 (N_16818,N_15454,N_14982);
nor U16819 (N_16819,N_13662,N_13045);
or U16820 (N_16820,N_15524,N_13887);
xor U16821 (N_16821,N_15394,N_14668);
xor U16822 (N_16822,N_12637,N_12643);
xnor U16823 (N_16823,N_12697,N_13429);
nor U16824 (N_16824,N_13951,N_14858);
xnor U16825 (N_16825,N_13387,N_12762);
and U16826 (N_16826,N_13090,N_15619);
nand U16827 (N_16827,N_13453,N_14078);
nand U16828 (N_16828,N_15172,N_13926);
nor U16829 (N_16829,N_12800,N_13003);
or U16830 (N_16830,N_14804,N_12657);
and U16831 (N_16831,N_15608,N_14155);
or U16832 (N_16832,N_14112,N_14080);
and U16833 (N_16833,N_12524,N_13729);
or U16834 (N_16834,N_14799,N_14269);
nor U16835 (N_16835,N_12679,N_12923);
and U16836 (N_16836,N_14418,N_13960);
and U16837 (N_16837,N_15159,N_13002);
or U16838 (N_16838,N_15183,N_15053);
and U16839 (N_16839,N_13750,N_13358);
xor U16840 (N_16840,N_12568,N_14923);
xor U16841 (N_16841,N_15428,N_14020);
and U16842 (N_16842,N_14702,N_13391);
and U16843 (N_16843,N_14833,N_15042);
nor U16844 (N_16844,N_15467,N_15032);
nand U16845 (N_16845,N_13174,N_14703);
nand U16846 (N_16846,N_13604,N_15485);
xnor U16847 (N_16847,N_15472,N_14868);
xnor U16848 (N_16848,N_13745,N_13890);
nor U16849 (N_16849,N_15557,N_13558);
and U16850 (N_16850,N_14788,N_15565);
xor U16851 (N_16851,N_14367,N_15517);
or U16852 (N_16852,N_12739,N_15119);
nor U16853 (N_16853,N_15287,N_13654);
or U16854 (N_16854,N_15153,N_13182);
nand U16855 (N_16855,N_12600,N_13795);
and U16856 (N_16856,N_12797,N_13933);
nor U16857 (N_16857,N_13627,N_15556);
nor U16858 (N_16858,N_14101,N_13248);
nor U16859 (N_16859,N_14302,N_15077);
or U16860 (N_16860,N_15415,N_13394);
nor U16861 (N_16861,N_15611,N_15030);
nor U16862 (N_16862,N_12814,N_15239);
nor U16863 (N_16863,N_14570,N_13180);
nand U16864 (N_16864,N_12633,N_14495);
xor U16865 (N_16865,N_13927,N_15269);
nor U16866 (N_16866,N_13187,N_15129);
or U16867 (N_16867,N_13049,N_14114);
xnor U16868 (N_16868,N_14213,N_14864);
nand U16869 (N_16869,N_13778,N_13758);
nor U16870 (N_16870,N_14154,N_13173);
xor U16871 (N_16871,N_13374,N_12752);
xor U16872 (N_16872,N_13603,N_13356);
xor U16873 (N_16873,N_13737,N_14675);
and U16874 (N_16874,N_15009,N_15058);
nor U16875 (N_16875,N_15366,N_13742);
and U16876 (N_16876,N_13589,N_13121);
or U16877 (N_16877,N_13233,N_13346);
nand U16878 (N_16878,N_12821,N_14975);
nor U16879 (N_16879,N_14943,N_13375);
nand U16880 (N_16880,N_14713,N_13015);
and U16881 (N_16881,N_14280,N_13583);
and U16882 (N_16882,N_14391,N_15458);
or U16883 (N_16883,N_13256,N_14245);
or U16884 (N_16884,N_13315,N_14319);
nor U16885 (N_16885,N_14691,N_14718);
xnor U16886 (N_16886,N_13468,N_12971);
xor U16887 (N_16887,N_14551,N_13615);
or U16888 (N_16888,N_12910,N_13886);
or U16889 (N_16889,N_13804,N_14434);
nor U16890 (N_16890,N_13042,N_13738);
nand U16891 (N_16891,N_12758,N_12508);
nand U16892 (N_16892,N_13665,N_12676);
xor U16893 (N_16893,N_13060,N_14728);
nand U16894 (N_16894,N_12553,N_14970);
nand U16895 (N_16895,N_12556,N_13162);
or U16896 (N_16896,N_15071,N_12776);
nand U16897 (N_16897,N_14173,N_14910);
nand U16898 (N_16898,N_15161,N_13186);
or U16899 (N_16899,N_14598,N_13889);
xor U16900 (N_16900,N_14113,N_15468);
nand U16901 (N_16901,N_12841,N_14563);
xnor U16902 (N_16902,N_14532,N_15149);
and U16903 (N_16903,N_12848,N_14700);
or U16904 (N_16904,N_15457,N_12614);
nor U16905 (N_16905,N_12531,N_13649);
or U16906 (N_16906,N_13385,N_14789);
and U16907 (N_16907,N_13511,N_13881);
nand U16908 (N_16908,N_12693,N_15562);
and U16909 (N_16909,N_12941,N_13648);
or U16910 (N_16910,N_13984,N_14153);
xor U16911 (N_16911,N_13961,N_14490);
nor U16912 (N_16912,N_14753,N_15135);
and U16913 (N_16913,N_14867,N_12886);
xnor U16914 (N_16914,N_15610,N_14872);
nand U16915 (N_16915,N_13736,N_12829);
xnor U16916 (N_16916,N_15450,N_14950);
nand U16917 (N_16917,N_13826,N_14348);
and U16918 (N_16918,N_14569,N_13275);
nor U16919 (N_16919,N_13463,N_14743);
nor U16920 (N_16920,N_13370,N_13404);
xor U16921 (N_16921,N_15381,N_15583);
nor U16922 (N_16922,N_15162,N_15490);
and U16923 (N_16923,N_14227,N_13535);
or U16924 (N_16924,N_14446,N_12842);
xnor U16925 (N_16925,N_14093,N_15150);
xor U16926 (N_16926,N_13431,N_13581);
and U16927 (N_16927,N_14138,N_14257);
nor U16928 (N_16928,N_13579,N_12838);
xnor U16929 (N_16929,N_14621,N_12849);
and U16930 (N_16930,N_13785,N_15047);
or U16931 (N_16931,N_15553,N_12807);
or U16932 (N_16932,N_15614,N_13148);
nand U16933 (N_16933,N_14132,N_12753);
xnor U16934 (N_16934,N_14262,N_14359);
and U16935 (N_16935,N_12551,N_12924);
or U16936 (N_16936,N_13134,N_13179);
or U16937 (N_16937,N_13754,N_12670);
and U16938 (N_16938,N_14115,N_13343);
nand U16939 (N_16939,N_12987,N_14187);
nand U16940 (N_16940,N_14617,N_13388);
nor U16941 (N_16941,N_15253,N_13376);
xor U16942 (N_16942,N_13706,N_12914);
or U16943 (N_16943,N_15247,N_13718);
and U16944 (N_16944,N_12564,N_14739);
xor U16945 (N_16945,N_12585,N_13036);
xor U16946 (N_16946,N_14576,N_14513);
xnor U16947 (N_16947,N_13272,N_13389);
nand U16948 (N_16948,N_13584,N_14028);
and U16949 (N_16949,N_14023,N_13441);
nand U16950 (N_16950,N_13089,N_15281);
nand U16951 (N_16951,N_12639,N_15014);
xnor U16952 (N_16952,N_14694,N_14239);
xnor U16953 (N_16953,N_13939,N_14511);
or U16954 (N_16954,N_13752,N_12687);
and U16955 (N_16955,N_14663,N_15383);
nor U16956 (N_16956,N_12852,N_15086);
nand U16957 (N_16957,N_13437,N_12893);
or U16958 (N_16958,N_13504,N_14216);
or U16959 (N_16959,N_13865,N_13844);
or U16960 (N_16960,N_14584,N_13965);
or U16961 (N_16961,N_14393,N_15601);
nand U16962 (N_16962,N_15074,N_13602);
xor U16963 (N_16963,N_12664,N_14790);
xnor U16964 (N_16964,N_14163,N_12632);
xor U16965 (N_16965,N_14452,N_12705);
and U16966 (N_16966,N_12817,N_14662);
and U16967 (N_16967,N_13260,N_14221);
or U16968 (N_16968,N_13561,N_13762);
xor U16969 (N_16969,N_13761,N_15151);
nand U16970 (N_16970,N_14467,N_14783);
and U16971 (N_16971,N_13279,N_14059);
and U16972 (N_16972,N_12616,N_14828);
nand U16973 (N_16973,N_14516,N_13524);
nand U16974 (N_16974,N_15076,N_13410);
and U16975 (N_16975,N_13677,N_13668);
and U16976 (N_16976,N_14039,N_13251);
xor U16977 (N_16977,N_12779,N_12802);
or U16978 (N_16978,N_13630,N_12944);
or U16979 (N_16979,N_12704,N_13782);
xnor U16980 (N_16980,N_13586,N_13273);
xor U16981 (N_16981,N_15431,N_13954);
nor U16982 (N_16982,N_15252,N_13505);
nand U16983 (N_16983,N_15355,N_14888);
nand U16984 (N_16984,N_14940,N_12750);
nand U16985 (N_16985,N_15275,N_13166);
xnor U16986 (N_16986,N_12897,N_14437);
and U16987 (N_16987,N_14377,N_13730);
xor U16988 (N_16988,N_14519,N_15380);
nor U16989 (N_16989,N_14949,N_13700);
or U16990 (N_16990,N_15362,N_12953);
xor U16991 (N_16991,N_14831,N_14972);
xnor U16992 (N_16992,N_13816,N_15372);
xnor U16993 (N_16993,N_14510,N_14404);
and U16994 (N_16994,N_15388,N_14477);
nor U16995 (N_16995,N_14942,N_13494);
nor U16996 (N_16996,N_12958,N_14104);
or U16997 (N_16997,N_15203,N_13967);
nand U16998 (N_16998,N_14708,N_13236);
or U16999 (N_16999,N_14766,N_12566);
nand U17000 (N_17000,N_15217,N_13510);
nand U17001 (N_17001,N_15540,N_13159);
or U17002 (N_17002,N_14999,N_13432);
nor U17003 (N_17003,N_13077,N_14006);
nand U17004 (N_17004,N_12728,N_13014);
and U17005 (N_17005,N_13789,N_13111);
or U17006 (N_17006,N_15335,N_14281);
xor U17007 (N_17007,N_13342,N_15623);
and U17008 (N_17008,N_14620,N_15288);
xor U17009 (N_17009,N_12994,N_13352);
and U17010 (N_17010,N_13681,N_12805);
or U17011 (N_17011,N_13492,N_13101);
nor U17012 (N_17012,N_14660,N_14931);
nor U17013 (N_17013,N_13707,N_12806);
and U17014 (N_17014,N_15618,N_12742);
xor U17015 (N_17015,N_13733,N_15179);
and U17016 (N_17016,N_12515,N_12588);
nand U17017 (N_17017,N_13212,N_14597);
and U17018 (N_17018,N_15502,N_14401);
or U17019 (N_17019,N_14127,N_12799);
xnor U17020 (N_17020,N_15291,N_14549);
or U17021 (N_17021,N_13365,N_14594);
or U17022 (N_17022,N_12939,N_15420);
xor U17023 (N_17023,N_13990,N_12976);
nand U17024 (N_17024,N_13768,N_15264);
and U17025 (N_17025,N_14458,N_14419);
nand U17026 (N_17026,N_13149,N_14664);
xnor U17027 (N_17027,N_14448,N_12896);
xor U17028 (N_17028,N_12610,N_12770);
or U17029 (N_17029,N_15412,N_13544);
nand U17030 (N_17030,N_15005,N_15581);
or U17031 (N_17031,N_14850,N_13949);
nor U17032 (N_17032,N_14632,N_13469);
and U17033 (N_17033,N_13756,N_13451);
and U17034 (N_17034,N_14004,N_13842);
xor U17035 (N_17035,N_14398,N_15055);
xor U17036 (N_17036,N_13925,N_13892);
and U17037 (N_17037,N_13192,N_12913);
nor U17038 (N_17038,N_14320,N_13098);
or U17039 (N_17039,N_14523,N_13152);
nand U17040 (N_17040,N_12725,N_13606);
and U17041 (N_17041,N_14528,N_15385);
and U17042 (N_17042,N_14303,N_14622);
and U17043 (N_17043,N_14608,N_15333);
or U17044 (N_17044,N_12766,N_14465);
nor U17045 (N_17045,N_12757,N_15300);
xor U17046 (N_17046,N_15369,N_13122);
nand U17047 (N_17047,N_15041,N_12538);
or U17048 (N_17048,N_14913,N_13438);
nand U17049 (N_17049,N_15590,N_14137);
and U17050 (N_17050,N_12831,N_14029);
nand U17051 (N_17051,N_15440,N_12804);
or U17052 (N_17052,N_12623,N_13473);
or U17053 (N_17053,N_12726,N_14149);
xor U17054 (N_17054,N_14914,N_13916);
nor U17055 (N_17055,N_12658,N_12887);
xor U17056 (N_17056,N_14851,N_14976);
xnor U17057 (N_17057,N_14234,N_14870);
nor U17058 (N_17058,N_13948,N_14270);
or U17059 (N_17059,N_14479,N_12743);
nor U17060 (N_17060,N_15270,N_12525);
nand U17061 (N_17061,N_14232,N_14343);
nand U17062 (N_17062,N_12875,N_13728);
xor U17063 (N_17063,N_14757,N_12998);
nor U17064 (N_17064,N_12712,N_14884);
or U17065 (N_17065,N_13988,N_13713);
and U17066 (N_17066,N_15464,N_14772);
and U17067 (N_17067,N_14565,N_14895);
and U17068 (N_17068,N_12967,N_13380);
or U17069 (N_17069,N_13213,N_14758);
or U17070 (N_17070,N_14053,N_14315);
nand U17071 (N_17071,N_14983,N_14294);
nand U17072 (N_17072,N_14304,N_14188);
nor U17073 (N_17073,N_15521,N_13672);
nand U17074 (N_17074,N_12922,N_15526);
xor U17075 (N_17075,N_14861,N_13258);
or U17076 (N_17076,N_13546,N_14508);
nand U17077 (N_17077,N_15572,N_14489);
nand U17078 (N_17078,N_14143,N_13332);
nand U17079 (N_17079,N_14615,N_15201);
xnor U17080 (N_17080,N_15006,N_13357);
and U17081 (N_17081,N_14212,N_15096);
and U17082 (N_17082,N_14552,N_14507);
nand U17083 (N_17083,N_15329,N_12830);
or U17084 (N_17084,N_13215,N_13470);
nand U17085 (N_17085,N_14440,N_15126);
and U17086 (N_17086,N_14797,N_15019);
and U17087 (N_17087,N_13992,N_14102);
xnor U17088 (N_17088,N_15423,N_13232);
and U17089 (N_17089,N_14533,N_14658);
or U17090 (N_17090,N_13208,N_14904);
and U17091 (N_17091,N_15439,N_15356);
and U17092 (N_17092,N_13319,N_14782);
or U17093 (N_17093,N_12868,N_14969);
nand U17094 (N_17094,N_13137,N_12764);
nor U17095 (N_17095,N_14649,N_13755);
nor U17096 (N_17096,N_15393,N_12929);
and U17097 (N_17097,N_15211,N_14368);
nor U17098 (N_17098,N_12715,N_15494);
nor U17099 (N_17099,N_15541,N_12717);
nand U17100 (N_17100,N_14760,N_13161);
xnor U17101 (N_17101,N_12507,N_13381);
xor U17102 (N_17102,N_13628,N_14542);
and U17103 (N_17103,N_14853,N_13110);
and U17104 (N_17104,N_13116,N_12885);
nor U17105 (N_17105,N_14988,N_12650);
nor U17106 (N_17106,N_14818,N_14509);
or U17107 (N_17107,N_13796,N_13962);
nand U17108 (N_17108,N_13265,N_12612);
nor U17109 (N_17109,N_14031,N_13019);
nor U17110 (N_17110,N_14557,N_15432);
or U17111 (N_17111,N_14619,N_15002);
xor U17112 (N_17112,N_14396,N_15343);
xnor U17113 (N_17113,N_14669,N_13421);
or U17114 (N_17114,N_14117,N_14899);
xnor U17115 (N_17115,N_14993,N_13096);
and U17116 (N_17116,N_12560,N_15034);
xnor U17117 (N_17117,N_12977,N_13784);
or U17118 (N_17118,N_15604,N_13010);
or U17119 (N_17119,N_15229,N_13051);
xnor U17120 (N_17120,N_12815,N_15561);
nor U17121 (N_17121,N_13915,N_14167);
and U17122 (N_17122,N_13574,N_14762);
xnor U17123 (N_17123,N_15156,N_12973);
nand U17124 (N_17124,N_15243,N_14644);
and U17125 (N_17125,N_13637,N_12737);
or U17126 (N_17126,N_13141,N_13061);
nor U17127 (N_17127,N_14571,N_14123);
nor U17128 (N_17128,N_12783,N_14334);
or U17129 (N_17129,N_15127,N_12669);
xnor U17130 (N_17130,N_12644,N_13054);
nor U17131 (N_17131,N_14369,N_14337);
nand U17132 (N_17132,N_13769,N_13197);
nand U17133 (N_17133,N_15137,N_14773);
or U17134 (N_17134,N_12906,N_14191);
and U17135 (N_17135,N_14200,N_12900);
nand U17136 (N_17136,N_15518,N_13938);
and U17137 (N_17137,N_13112,N_15104);
or U17138 (N_17138,N_14726,N_14330);
xnor U17139 (N_17139,N_15095,N_13334);
nand U17140 (N_17140,N_12763,N_12858);
xnor U17141 (N_17141,N_14909,N_15143);
xor U17142 (N_17142,N_14566,N_12940);
nand U17143 (N_17143,N_13671,N_14802);
and U17144 (N_17144,N_14548,N_14506);
and U17145 (N_17145,N_13772,N_14778);
or U17146 (N_17146,N_14933,N_14640);
and U17147 (N_17147,N_14470,N_14447);
xor U17148 (N_17148,N_13063,N_13565);
and U17149 (N_17149,N_13127,N_14165);
and U17150 (N_17150,N_14912,N_14174);
xor U17151 (N_17151,N_14453,N_14459);
or U17152 (N_17152,N_12591,N_15214);
nor U17153 (N_17153,N_15416,N_15206);
and U17154 (N_17154,N_14624,N_13687);
nor U17155 (N_17155,N_14321,N_14291);
xor U17156 (N_17156,N_12992,N_13635);
xnor U17157 (N_17157,N_15606,N_14259);
nand U17158 (N_17158,N_12611,N_15073);
and U17159 (N_17159,N_12554,N_12874);
and U17160 (N_17160,N_13757,N_13800);
xor U17161 (N_17161,N_15469,N_12521);
xor U17162 (N_17162,N_13133,N_14894);
xor U17163 (N_17163,N_15000,N_14430);
or U17164 (N_17164,N_15501,N_14015);
or U17165 (N_17165,N_12688,N_14237);
nand U17166 (N_17166,N_13853,N_13349);
xor U17167 (N_17167,N_12513,N_13219);
or U17168 (N_17168,N_12968,N_13508);
xnor U17169 (N_17169,N_13715,N_14326);
nor U17170 (N_17170,N_15145,N_13363);
nor U17171 (N_17171,N_13863,N_14071);
nor U17172 (N_17172,N_13499,N_14665);
and U17173 (N_17173,N_13445,N_12864);
or U17174 (N_17174,N_15255,N_14791);
and U17175 (N_17175,N_12569,N_14439);
xnor U17176 (N_17176,N_13512,N_12671);
nand U17177 (N_17177,N_14560,N_13513);
and U17178 (N_17178,N_15023,N_13239);
xnor U17179 (N_17179,N_14705,N_12945);
and U17180 (N_17180,N_13620,N_12767);
nand U17181 (N_17181,N_14126,N_12880);
or U17182 (N_17182,N_12773,N_13585);
or U17183 (N_17183,N_13196,N_14266);
or U17184 (N_17184,N_15598,N_12811);
nor U17185 (N_17185,N_14825,N_13848);
or U17186 (N_17186,N_13727,N_13072);
xnor U17187 (N_17187,N_12674,N_15387);
nand U17188 (N_17188,N_12892,N_13052);
and U17189 (N_17189,N_12831,N_13527);
xnor U17190 (N_17190,N_13408,N_14050);
nand U17191 (N_17191,N_13282,N_14682);
nor U17192 (N_17192,N_13497,N_14485);
and U17193 (N_17193,N_14780,N_14615);
and U17194 (N_17194,N_12867,N_15500);
or U17195 (N_17195,N_14259,N_13388);
nor U17196 (N_17196,N_13318,N_12514);
nand U17197 (N_17197,N_13906,N_14170);
nand U17198 (N_17198,N_13347,N_12994);
and U17199 (N_17199,N_14109,N_13463);
and U17200 (N_17200,N_14324,N_13843);
and U17201 (N_17201,N_13424,N_14626);
or U17202 (N_17202,N_13649,N_15344);
and U17203 (N_17203,N_13335,N_14775);
nor U17204 (N_17204,N_12941,N_13483);
nor U17205 (N_17205,N_13098,N_12801);
nand U17206 (N_17206,N_14777,N_15593);
nor U17207 (N_17207,N_15178,N_14213);
nand U17208 (N_17208,N_13562,N_13782);
nor U17209 (N_17209,N_12515,N_13581);
xnor U17210 (N_17210,N_14010,N_15396);
and U17211 (N_17211,N_13171,N_13242);
and U17212 (N_17212,N_14575,N_13515);
xnor U17213 (N_17213,N_13916,N_13426);
and U17214 (N_17214,N_13489,N_14378);
or U17215 (N_17215,N_14406,N_12799);
nand U17216 (N_17216,N_15269,N_14262);
nor U17217 (N_17217,N_12602,N_12920);
nor U17218 (N_17218,N_13142,N_14060);
nand U17219 (N_17219,N_12994,N_14654);
xor U17220 (N_17220,N_13827,N_13894);
nand U17221 (N_17221,N_14872,N_14459);
nand U17222 (N_17222,N_12580,N_13398);
and U17223 (N_17223,N_15228,N_12810);
and U17224 (N_17224,N_13085,N_12918);
or U17225 (N_17225,N_12636,N_14275);
or U17226 (N_17226,N_15063,N_15204);
or U17227 (N_17227,N_15380,N_14055);
nor U17228 (N_17228,N_13294,N_12975);
nand U17229 (N_17229,N_14805,N_15206);
nand U17230 (N_17230,N_15398,N_15540);
nand U17231 (N_17231,N_15312,N_12678);
and U17232 (N_17232,N_15096,N_14466);
or U17233 (N_17233,N_13664,N_13779);
nand U17234 (N_17234,N_15496,N_13487);
and U17235 (N_17235,N_13874,N_14229);
or U17236 (N_17236,N_15448,N_13547);
xor U17237 (N_17237,N_13786,N_14747);
or U17238 (N_17238,N_12650,N_12625);
or U17239 (N_17239,N_13524,N_13999);
xor U17240 (N_17240,N_13133,N_13630);
and U17241 (N_17241,N_14186,N_14817);
nand U17242 (N_17242,N_15374,N_15185);
and U17243 (N_17243,N_15226,N_14659);
and U17244 (N_17244,N_15568,N_13229);
nand U17245 (N_17245,N_15436,N_13382);
or U17246 (N_17246,N_13102,N_15258);
xor U17247 (N_17247,N_12695,N_15510);
and U17248 (N_17248,N_15091,N_12668);
or U17249 (N_17249,N_14243,N_13545);
nor U17250 (N_17250,N_13900,N_15604);
nor U17251 (N_17251,N_13038,N_13851);
or U17252 (N_17252,N_13533,N_13803);
or U17253 (N_17253,N_12559,N_15307);
nand U17254 (N_17254,N_12623,N_12949);
nor U17255 (N_17255,N_14722,N_13203);
nor U17256 (N_17256,N_13135,N_12699);
nor U17257 (N_17257,N_15095,N_15123);
or U17258 (N_17258,N_15396,N_15609);
nor U17259 (N_17259,N_15347,N_14074);
nand U17260 (N_17260,N_14837,N_12775);
xor U17261 (N_17261,N_15209,N_15395);
nor U17262 (N_17262,N_12624,N_13591);
xnor U17263 (N_17263,N_13560,N_13719);
xor U17264 (N_17264,N_13660,N_12516);
xnor U17265 (N_17265,N_14044,N_13239);
or U17266 (N_17266,N_14453,N_15349);
and U17267 (N_17267,N_14043,N_12773);
or U17268 (N_17268,N_14082,N_12968);
and U17269 (N_17269,N_14314,N_13086);
nor U17270 (N_17270,N_13861,N_12600);
nor U17271 (N_17271,N_14664,N_14047);
nor U17272 (N_17272,N_12857,N_12891);
xnor U17273 (N_17273,N_15146,N_14116);
nor U17274 (N_17274,N_14850,N_13428);
xnor U17275 (N_17275,N_15060,N_14293);
or U17276 (N_17276,N_12531,N_13659);
nand U17277 (N_17277,N_13984,N_15498);
nor U17278 (N_17278,N_13104,N_12721);
nor U17279 (N_17279,N_14454,N_13425);
and U17280 (N_17280,N_13523,N_12615);
xor U17281 (N_17281,N_13924,N_14664);
xnor U17282 (N_17282,N_14536,N_14718);
or U17283 (N_17283,N_14653,N_13276);
xor U17284 (N_17284,N_14949,N_14349);
or U17285 (N_17285,N_15469,N_14659);
nor U17286 (N_17286,N_15361,N_13091);
nand U17287 (N_17287,N_13567,N_14092);
nand U17288 (N_17288,N_14918,N_14716);
xor U17289 (N_17289,N_14573,N_13882);
or U17290 (N_17290,N_13324,N_14494);
or U17291 (N_17291,N_13318,N_12526);
and U17292 (N_17292,N_15129,N_15288);
and U17293 (N_17293,N_12961,N_13496);
and U17294 (N_17294,N_13704,N_14113);
or U17295 (N_17295,N_12839,N_12528);
nor U17296 (N_17296,N_12903,N_14488);
or U17297 (N_17297,N_12990,N_13450);
or U17298 (N_17298,N_13311,N_14086);
nand U17299 (N_17299,N_14606,N_14160);
nor U17300 (N_17300,N_14018,N_15123);
and U17301 (N_17301,N_14774,N_12721);
nor U17302 (N_17302,N_13282,N_14259);
and U17303 (N_17303,N_14428,N_14416);
or U17304 (N_17304,N_13704,N_13062);
and U17305 (N_17305,N_13941,N_15177);
or U17306 (N_17306,N_14319,N_14497);
nand U17307 (N_17307,N_14397,N_13775);
xor U17308 (N_17308,N_13551,N_12957);
xor U17309 (N_17309,N_15217,N_13080);
and U17310 (N_17310,N_14101,N_13828);
nor U17311 (N_17311,N_14338,N_14456);
xor U17312 (N_17312,N_15195,N_15050);
xnor U17313 (N_17313,N_13156,N_13899);
nor U17314 (N_17314,N_15350,N_14049);
nand U17315 (N_17315,N_14203,N_14971);
and U17316 (N_17316,N_12647,N_14492);
nand U17317 (N_17317,N_13650,N_14292);
and U17318 (N_17318,N_14935,N_14296);
xor U17319 (N_17319,N_14504,N_13622);
and U17320 (N_17320,N_13979,N_15512);
xor U17321 (N_17321,N_13785,N_14209);
nor U17322 (N_17322,N_13632,N_13998);
xnor U17323 (N_17323,N_13694,N_12735);
or U17324 (N_17324,N_13097,N_14971);
nor U17325 (N_17325,N_14819,N_14716);
or U17326 (N_17326,N_15009,N_13001);
or U17327 (N_17327,N_13390,N_14078);
nand U17328 (N_17328,N_13007,N_13082);
and U17329 (N_17329,N_14090,N_14714);
nor U17330 (N_17330,N_14304,N_14539);
nand U17331 (N_17331,N_14875,N_14546);
xnor U17332 (N_17332,N_15258,N_13207);
nand U17333 (N_17333,N_13448,N_15110);
nand U17334 (N_17334,N_14795,N_13423);
xor U17335 (N_17335,N_14779,N_15271);
xor U17336 (N_17336,N_13948,N_15083);
nand U17337 (N_17337,N_14227,N_14445);
xnor U17338 (N_17338,N_15160,N_15365);
or U17339 (N_17339,N_14031,N_13215);
nand U17340 (N_17340,N_15013,N_12571);
and U17341 (N_17341,N_14035,N_13201);
xnor U17342 (N_17342,N_13719,N_14776);
or U17343 (N_17343,N_12506,N_12925);
nand U17344 (N_17344,N_14790,N_14808);
nor U17345 (N_17345,N_14525,N_12771);
xnor U17346 (N_17346,N_14275,N_15333);
and U17347 (N_17347,N_14161,N_12654);
or U17348 (N_17348,N_13296,N_13640);
and U17349 (N_17349,N_15013,N_13952);
and U17350 (N_17350,N_14620,N_15266);
or U17351 (N_17351,N_14477,N_14437);
or U17352 (N_17352,N_14707,N_13039);
xor U17353 (N_17353,N_15033,N_13859);
or U17354 (N_17354,N_13330,N_12592);
or U17355 (N_17355,N_13794,N_12878);
and U17356 (N_17356,N_13704,N_14129);
or U17357 (N_17357,N_14048,N_15451);
and U17358 (N_17358,N_14103,N_14205);
or U17359 (N_17359,N_12727,N_12716);
or U17360 (N_17360,N_14319,N_14404);
xnor U17361 (N_17361,N_15390,N_14168);
nor U17362 (N_17362,N_14556,N_14250);
xnor U17363 (N_17363,N_12970,N_14370);
nor U17364 (N_17364,N_13121,N_13995);
and U17365 (N_17365,N_13889,N_12998);
nor U17366 (N_17366,N_15350,N_14936);
nor U17367 (N_17367,N_13892,N_14122);
and U17368 (N_17368,N_14834,N_15454);
xnor U17369 (N_17369,N_13662,N_13227);
or U17370 (N_17370,N_13628,N_14126);
or U17371 (N_17371,N_12722,N_14600);
or U17372 (N_17372,N_13257,N_14147);
and U17373 (N_17373,N_13632,N_13762);
or U17374 (N_17374,N_12762,N_15156);
nand U17375 (N_17375,N_15592,N_13024);
and U17376 (N_17376,N_13845,N_12782);
nor U17377 (N_17377,N_12540,N_14749);
and U17378 (N_17378,N_15034,N_14694);
or U17379 (N_17379,N_14939,N_14831);
xor U17380 (N_17380,N_15218,N_13153);
nor U17381 (N_17381,N_13031,N_12980);
nor U17382 (N_17382,N_15069,N_14618);
nor U17383 (N_17383,N_15483,N_12655);
and U17384 (N_17384,N_14521,N_14136);
and U17385 (N_17385,N_14731,N_13333);
or U17386 (N_17386,N_12901,N_12890);
nor U17387 (N_17387,N_13349,N_14451);
nand U17388 (N_17388,N_13982,N_14874);
or U17389 (N_17389,N_14445,N_12637);
nand U17390 (N_17390,N_13708,N_14935);
xor U17391 (N_17391,N_13362,N_14124);
nand U17392 (N_17392,N_12592,N_13618);
xnor U17393 (N_17393,N_14436,N_13738);
nor U17394 (N_17394,N_14111,N_14846);
or U17395 (N_17395,N_13216,N_13227);
nor U17396 (N_17396,N_12899,N_13149);
and U17397 (N_17397,N_14132,N_12890);
and U17398 (N_17398,N_14374,N_13675);
or U17399 (N_17399,N_13410,N_14327);
or U17400 (N_17400,N_15501,N_15403);
xor U17401 (N_17401,N_15069,N_15239);
nand U17402 (N_17402,N_15113,N_14035);
and U17403 (N_17403,N_12698,N_13484);
nand U17404 (N_17404,N_14770,N_14117);
nand U17405 (N_17405,N_12641,N_14571);
xnor U17406 (N_17406,N_12852,N_12908);
and U17407 (N_17407,N_14228,N_13823);
nor U17408 (N_17408,N_13624,N_15370);
and U17409 (N_17409,N_14765,N_15428);
or U17410 (N_17410,N_13921,N_12785);
xor U17411 (N_17411,N_14145,N_12977);
xor U17412 (N_17412,N_13111,N_13152);
xnor U17413 (N_17413,N_15362,N_12541);
nor U17414 (N_17414,N_14512,N_14056);
nor U17415 (N_17415,N_13322,N_13516);
nand U17416 (N_17416,N_13107,N_14411);
nor U17417 (N_17417,N_13183,N_14872);
nand U17418 (N_17418,N_13903,N_14489);
nand U17419 (N_17419,N_14410,N_14295);
and U17420 (N_17420,N_14961,N_13062);
and U17421 (N_17421,N_13701,N_14036);
nand U17422 (N_17422,N_14735,N_13162);
or U17423 (N_17423,N_14464,N_13082);
nor U17424 (N_17424,N_13003,N_15137);
and U17425 (N_17425,N_14800,N_12963);
nand U17426 (N_17426,N_14291,N_15114);
and U17427 (N_17427,N_13821,N_14744);
xnor U17428 (N_17428,N_13645,N_13045);
nand U17429 (N_17429,N_14306,N_15235);
nor U17430 (N_17430,N_12591,N_13584);
nand U17431 (N_17431,N_13071,N_12825);
nand U17432 (N_17432,N_13491,N_15058);
and U17433 (N_17433,N_15383,N_15515);
nand U17434 (N_17434,N_12545,N_13951);
or U17435 (N_17435,N_12711,N_14428);
nor U17436 (N_17436,N_14479,N_13106);
and U17437 (N_17437,N_15114,N_15103);
or U17438 (N_17438,N_13670,N_15049);
nor U17439 (N_17439,N_13339,N_15483);
and U17440 (N_17440,N_14246,N_13291);
or U17441 (N_17441,N_14177,N_13376);
or U17442 (N_17442,N_13659,N_13058);
nand U17443 (N_17443,N_14955,N_12700);
nand U17444 (N_17444,N_14418,N_14743);
xor U17445 (N_17445,N_14017,N_12950);
xor U17446 (N_17446,N_13212,N_13846);
nand U17447 (N_17447,N_14444,N_13143);
nand U17448 (N_17448,N_13494,N_14835);
xnor U17449 (N_17449,N_14828,N_15343);
or U17450 (N_17450,N_13475,N_13039);
nor U17451 (N_17451,N_13480,N_15112);
nor U17452 (N_17452,N_15195,N_15548);
or U17453 (N_17453,N_14540,N_15341);
nand U17454 (N_17454,N_13603,N_14577);
or U17455 (N_17455,N_15369,N_13619);
nand U17456 (N_17456,N_14913,N_12958);
or U17457 (N_17457,N_15124,N_12686);
xor U17458 (N_17458,N_12904,N_14869);
xnor U17459 (N_17459,N_13924,N_14785);
or U17460 (N_17460,N_13000,N_15058);
xor U17461 (N_17461,N_12533,N_14436);
nand U17462 (N_17462,N_13295,N_14195);
xor U17463 (N_17463,N_13856,N_12862);
xor U17464 (N_17464,N_15094,N_14236);
nand U17465 (N_17465,N_13447,N_14984);
xnor U17466 (N_17466,N_13158,N_13659);
or U17467 (N_17467,N_13355,N_12618);
nand U17468 (N_17468,N_15329,N_14708);
xor U17469 (N_17469,N_14526,N_14629);
xnor U17470 (N_17470,N_13395,N_13507);
and U17471 (N_17471,N_13459,N_13356);
nor U17472 (N_17472,N_13044,N_13731);
nor U17473 (N_17473,N_12757,N_15041);
and U17474 (N_17474,N_15141,N_15087);
and U17475 (N_17475,N_12737,N_12882);
xor U17476 (N_17476,N_14448,N_13871);
nor U17477 (N_17477,N_13642,N_12513);
or U17478 (N_17478,N_12606,N_13316);
and U17479 (N_17479,N_14719,N_14472);
or U17480 (N_17480,N_15269,N_12831);
or U17481 (N_17481,N_15165,N_13292);
xor U17482 (N_17482,N_15558,N_13904);
or U17483 (N_17483,N_13732,N_14808);
and U17484 (N_17484,N_12844,N_12876);
or U17485 (N_17485,N_15064,N_15162);
nand U17486 (N_17486,N_13378,N_12524);
nand U17487 (N_17487,N_15254,N_13837);
xnor U17488 (N_17488,N_14823,N_14188);
xor U17489 (N_17489,N_13094,N_14873);
xor U17490 (N_17490,N_13737,N_13543);
nor U17491 (N_17491,N_14692,N_15530);
xor U17492 (N_17492,N_14667,N_14956);
or U17493 (N_17493,N_13781,N_13495);
and U17494 (N_17494,N_15294,N_13554);
nor U17495 (N_17495,N_14259,N_14805);
or U17496 (N_17496,N_15065,N_13836);
and U17497 (N_17497,N_12588,N_12737);
nor U17498 (N_17498,N_14657,N_13560);
nor U17499 (N_17499,N_13776,N_14120);
or U17500 (N_17500,N_13673,N_14908);
and U17501 (N_17501,N_13382,N_13435);
or U17502 (N_17502,N_13621,N_14283);
or U17503 (N_17503,N_13318,N_13929);
or U17504 (N_17504,N_15306,N_14840);
nand U17505 (N_17505,N_14115,N_14338);
or U17506 (N_17506,N_13849,N_13883);
or U17507 (N_17507,N_13343,N_15355);
nand U17508 (N_17508,N_14468,N_14418);
and U17509 (N_17509,N_12835,N_13892);
nor U17510 (N_17510,N_13283,N_14637);
xor U17511 (N_17511,N_15473,N_14734);
nand U17512 (N_17512,N_12857,N_15006);
nor U17513 (N_17513,N_14683,N_14532);
nor U17514 (N_17514,N_13816,N_15589);
nor U17515 (N_17515,N_13164,N_12740);
xnor U17516 (N_17516,N_12882,N_14675);
and U17517 (N_17517,N_15148,N_13453);
and U17518 (N_17518,N_15205,N_13554);
xor U17519 (N_17519,N_15123,N_15073);
and U17520 (N_17520,N_12829,N_15021);
and U17521 (N_17521,N_14940,N_13345);
nand U17522 (N_17522,N_14721,N_13054);
nor U17523 (N_17523,N_14554,N_13713);
xnor U17524 (N_17524,N_14785,N_12677);
nor U17525 (N_17525,N_14973,N_14577);
xor U17526 (N_17526,N_12861,N_12881);
nor U17527 (N_17527,N_13612,N_14455);
and U17528 (N_17528,N_14021,N_13688);
or U17529 (N_17529,N_14322,N_13480);
xnor U17530 (N_17530,N_12621,N_13874);
and U17531 (N_17531,N_13935,N_14283);
nor U17532 (N_17532,N_15161,N_14663);
or U17533 (N_17533,N_14631,N_14603);
or U17534 (N_17534,N_14649,N_14944);
nand U17535 (N_17535,N_15222,N_13964);
or U17536 (N_17536,N_12860,N_15153);
and U17537 (N_17537,N_14665,N_14604);
or U17538 (N_17538,N_12638,N_13256);
and U17539 (N_17539,N_15140,N_15494);
and U17540 (N_17540,N_13251,N_14440);
or U17541 (N_17541,N_14245,N_13800);
nand U17542 (N_17542,N_14434,N_15114);
nand U17543 (N_17543,N_14189,N_14585);
nand U17544 (N_17544,N_13897,N_13294);
or U17545 (N_17545,N_13564,N_12956);
nor U17546 (N_17546,N_14996,N_13163);
xnor U17547 (N_17547,N_14324,N_14848);
nand U17548 (N_17548,N_14204,N_12984);
or U17549 (N_17549,N_12599,N_13873);
or U17550 (N_17550,N_12878,N_13160);
xor U17551 (N_17551,N_15530,N_15358);
and U17552 (N_17552,N_12634,N_13812);
or U17553 (N_17553,N_12771,N_12638);
nand U17554 (N_17554,N_13101,N_12894);
nand U17555 (N_17555,N_13028,N_13674);
and U17556 (N_17556,N_14538,N_15615);
nand U17557 (N_17557,N_13304,N_15360);
xnor U17558 (N_17558,N_15590,N_14311);
and U17559 (N_17559,N_15595,N_13431);
or U17560 (N_17560,N_12937,N_15254);
or U17561 (N_17561,N_13766,N_14664);
or U17562 (N_17562,N_12976,N_14044);
or U17563 (N_17563,N_14808,N_15071);
nand U17564 (N_17564,N_15229,N_14795);
nand U17565 (N_17565,N_15532,N_14763);
nor U17566 (N_17566,N_14031,N_14141);
or U17567 (N_17567,N_12668,N_13272);
nand U17568 (N_17568,N_14838,N_14928);
nor U17569 (N_17569,N_12554,N_12952);
xnor U17570 (N_17570,N_13636,N_12792);
nand U17571 (N_17571,N_14946,N_12992);
and U17572 (N_17572,N_14592,N_15194);
and U17573 (N_17573,N_12717,N_13215);
xor U17574 (N_17574,N_12816,N_15235);
xor U17575 (N_17575,N_14251,N_15287);
nor U17576 (N_17576,N_14140,N_15395);
xnor U17577 (N_17577,N_14392,N_12785);
xnor U17578 (N_17578,N_14259,N_13736);
nor U17579 (N_17579,N_14441,N_14846);
and U17580 (N_17580,N_14011,N_14519);
and U17581 (N_17581,N_13092,N_15149);
xor U17582 (N_17582,N_14077,N_14016);
nor U17583 (N_17583,N_14959,N_15041);
nor U17584 (N_17584,N_14575,N_12802);
or U17585 (N_17585,N_13139,N_15144);
nand U17586 (N_17586,N_15304,N_14028);
nor U17587 (N_17587,N_13697,N_14267);
or U17588 (N_17588,N_13139,N_15154);
nand U17589 (N_17589,N_14677,N_12705);
or U17590 (N_17590,N_12849,N_15214);
or U17591 (N_17591,N_15536,N_15425);
xor U17592 (N_17592,N_13470,N_13776);
xor U17593 (N_17593,N_12576,N_13489);
nor U17594 (N_17594,N_15108,N_13548);
xnor U17595 (N_17595,N_13863,N_14408);
nand U17596 (N_17596,N_14292,N_14674);
xnor U17597 (N_17597,N_13839,N_13981);
nand U17598 (N_17598,N_14505,N_14227);
xnor U17599 (N_17599,N_13735,N_12670);
nor U17600 (N_17600,N_14415,N_13883);
and U17601 (N_17601,N_14620,N_12814);
nand U17602 (N_17602,N_15611,N_14931);
and U17603 (N_17603,N_14688,N_14331);
xor U17604 (N_17604,N_14819,N_12911);
or U17605 (N_17605,N_14467,N_12841);
and U17606 (N_17606,N_12810,N_15068);
and U17607 (N_17607,N_13988,N_14171);
and U17608 (N_17608,N_13710,N_14426);
nor U17609 (N_17609,N_14967,N_13096);
xor U17610 (N_17610,N_14070,N_13955);
xor U17611 (N_17611,N_13791,N_15093);
xor U17612 (N_17612,N_12629,N_12508);
and U17613 (N_17613,N_12576,N_13337);
nand U17614 (N_17614,N_14308,N_15256);
nand U17615 (N_17615,N_12505,N_12969);
xnor U17616 (N_17616,N_15614,N_12761);
or U17617 (N_17617,N_13136,N_13067);
and U17618 (N_17618,N_13460,N_14776);
nor U17619 (N_17619,N_14304,N_13241);
xnor U17620 (N_17620,N_13862,N_12969);
and U17621 (N_17621,N_13204,N_13259);
or U17622 (N_17622,N_13226,N_13519);
xnor U17623 (N_17623,N_14568,N_12884);
xor U17624 (N_17624,N_12594,N_14993);
nand U17625 (N_17625,N_14690,N_12607);
and U17626 (N_17626,N_15402,N_13937);
xor U17627 (N_17627,N_12974,N_13749);
and U17628 (N_17628,N_13978,N_13025);
xor U17629 (N_17629,N_15008,N_15016);
nand U17630 (N_17630,N_14010,N_12722);
and U17631 (N_17631,N_13472,N_13841);
nor U17632 (N_17632,N_12952,N_14444);
or U17633 (N_17633,N_14360,N_14755);
xor U17634 (N_17634,N_14488,N_14055);
or U17635 (N_17635,N_14568,N_15614);
or U17636 (N_17636,N_14162,N_15318);
or U17637 (N_17637,N_13469,N_14910);
and U17638 (N_17638,N_14661,N_13793);
nor U17639 (N_17639,N_13604,N_13942);
nand U17640 (N_17640,N_13726,N_14593);
nand U17641 (N_17641,N_13728,N_14140);
nand U17642 (N_17642,N_12655,N_12642);
nand U17643 (N_17643,N_13180,N_13124);
xor U17644 (N_17644,N_13710,N_13619);
or U17645 (N_17645,N_13657,N_13662);
nand U17646 (N_17646,N_15224,N_15077);
or U17647 (N_17647,N_14070,N_15237);
nor U17648 (N_17648,N_14701,N_13622);
and U17649 (N_17649,N_13587,N_13511);
nor U17650 (N_17650,N_14010,N_12842);
xnor U17651 (N_17651,N_14883,N_15004);
nor U17652 (N_17652,N_12760,N_12701);
or U17653 (N_17653,N_12609,N_15454);
nand U17654 (N_17654,N_13222,N_15001);
nand U17655 (N_17655,N_15540,N_13760);
and U17656 (N_17656,N_13232,N_14662);
nor U17657 (N_17657,N_14144,N_12701);
nand U17658 (N_17658,N_13928,N_14271);
and U17659 (N_17659,N_13420,N_14970);
nor U17660 (N_17660,N_13492,N_14956);
and U17661 (N_17661,N_12987,N_14343);
nand U17662 (N_17662,N_14009,N_13340);
nand U17663 (N_17663,N_13655,N_14802);
and U17664 (N_17664,N_12762,N_14594);
nand U17665 (N_17665,N_13611,N_13519);
xor U17666 (N_17666,N_15476,N_15242);
nor U17667 (N_17667,N_15443,N_13123);
nand U17668 (N_17668,N_13035,N_15107);
xor U17669 (N_17669,N_13623,N_13330);
or U17670 (N_17670,N_14595,N_14636);
and U17671 (N_17671,N_15564,N_13863);
nand U17672 (N_17672,N_15598,N_15550);
nand U17673 (N_17673,N_15409,N_14469);
or U17674 (N_17674,N_12826,N_12646);
xnor U17675 (N_17675,N_12771,N_12949);
nand U17676 (N_17676,N_13343,N_13809);
xnor U17677 (N_17677,N_14603,N_12779);
xnor U17678 (N_17678,N_14050,N_15006);
nand U17679 (N_17679,N_14033,N_13911);
nor U17680 (N_17680,N_13806,N_15399);
and U17681 (N_17681,N_13789,N_13004);
nand U17682 (N_17682,N_14408,N_15385);
and U17683 (N_17683,N_13815,N_14361);
nand U17684 (N_17684,N_14169,N_12639);
nand U17685 (N_17685,N_15600,N_15128);
and U17686 (N_17686,N_12634,N_15037);
nor U17687 (N_17687,N_12614,N_15588);
xnor U17688 (N_17688,N_15066,N_13397);
nor U17689 (N_17689,N_12848,N_12706);
xnor U17690 (N_17690,N_13042,N_14806);
nand U17691 (N_17691,N_14163,N_13380);
nand U17692 (N_17692,N_14415,N_13097);
nor U17693 (N_17693,N_15041,N_13409);
and U17694 (N_17694,N_12652,N_13802);
and U17695 (N_17695,N_15443,N_15098);
or U17696 (N_17696,N_13587,N_13392);
or U17697 (N_17697,N_14656,N_14341);
xnor U17698 (N_17698,N_13167,N_14809);
xnor U17699 (N_17699,N_12674,N_13080);
xnor U17700 (N_17700,N_13103,N_13949);
xnor U17701 (N_17701,N_14255,N_15282);
nand U17702 (N_17702,N_14558,N_15219);
nor U17703 (N_17703,N_15538,N_15356);
or U17704 (N_17704,N_13054,N_15484);
nor U17705 (N_17705,N_15361,N_13683);
nor U17706 (N_17706,N_13374,N_15013);
nand U17707 (N_17707,N_14177,N_13529);
nand U17708 (N_17708,N_13637,N_14658);
and U17709 (N_17709,N_15474,N_14647);
nor U17710 (N_17710,N_14591,N_15237);
nand U17711 (N_17711,N_13805,N_13382);
and U17712 (N_17712,N_13300,N_15395);
and U17713 (N_17713,N_14798,N_15544);
nor U17714 (N_17714,N_14582,N_14112);
nor U17715 (N_17715,N_15257,N_14197);
nand U17716 (N_17716,N_14185,N_14488);
nand U17717 (N_17717,N_14317,N_12502);
nand U17718 (N_17718,N_12533,N_13405);
and U17719 (N_17719,N_13817,N_13161);
or U17720 (N_17720,N_15107,N_12796);
or U17721 (N_17721,N_12975,N_15484);
and U17722 (N_17722,N_14601,N_15214);
nand U17723 (N_17723,N_13528,N_15622);
and U17724 (N_17724,N_13220,N_13560);
or U17725 (N_17725,N_12703,N_14822);
xor U17726 (N_17726,N_15433,N_14651);
and U17727 (N_17727,N_14278,N_13328);
and U17728 (N_17728,N_14934,N_15520);
nand U17729 (N_17729,N_14983,N_12604);
nor U17730 (N_17730,N_14188,N_12602);
xnor U17731 (N_17731,N_15541,N_14844);
or U17732 (N_17732,N_13493,N_14907);
and U17733 (N_17733,N_12956,N_13169);
nand U17734 (N_17734,N_14362,N_14821);
xor U17735 (N_17735,N_12552,N_13190);
or U17736 (N_17736,N_13654,N_14585);
and U17737 (N_17737,N_13821,N_14915);
or U17738 (N_17738,N_15596,N_12518);
nor U17739 (N_17739,N_13324,N_13634);
or U17740 (N_17740,N_14885,N_13845);
and U17741 (N_17741,N_13182,N_13993);
xor U17742 (N_17742,N_12900,N_12667);
and U17743 (N_17743,N_13484,N_14104);
and U17744 (N_17744,N_12908,N_12674);
nor U17745 (N_17745,N_13996,N_13849);
xor U17746 (N_17746,N_14930,N_12915);
and U17747 (N_17747,N_15450,N_14935);
nor U17748 (N_17748,N_15583,N_14717);
nor U17749 (N_17749,N_13811,N_13324);
nor U17750 (N_17750,N_14620,N_14184);
xnor U17751 (N_17751,N_15005,N_15231);
nor U17752 (N_17752,N_14926,N_13903);
xor U17753 (N_17753,N_14909,N_13618);
and U17754 (N_17754,N_14301,N_13527);
nand U17755 (N_17755,N_12991,N_12627);
and U17756 (N_17756,N_13338,N_13918);
xnor U17757 (N_17757,N_13278,N_14253);
nand U17758 (N_17758,N_14721,N_12702);
nand U17759 (N_17759,N_12638,N_14938);
nor U17760 (N_17760,N_12577,N_13092);
xor U17761 (N_17761,N_14382,N_12953);
and U17762 (N_17762,N_13278,N_13130);
nand U17763 (N_17763,N_15209,N_14101);
nand U17764 (N_17764,N_12589,N_14535);
and U17765 (N_17765,N_14134,N_15163);
or U17766 (N_17766,N_13430,N_12539);
xor U17767 (N_17767,N_14956,N_14344);
nand U17768 (N_17768,N_12570,N_15340);
xor U17769 (N_17769,N_14019,N_15185);
nand U17770 (N_17770,N_13592,N_15374);
xnor U17771 (N_17771,N_14225,N_14426);
or U17772 (N_17772,N_12889,N_13842);
and U17773 (N_17773,N_15505,N_15160);
nand U17774 (N_17774,N_15201,N_14862);
or U17775 (N_17775,N_15276,N_13000);
nor U17776 (N_17776,N_13166,N_13836);
or U17777 (N_17777,N_13097,N_14981);
nor U17778 (N_17778,N_14108,N_15185);
nand U17779 (N_17779,N_14627,N_13292);
or U17780 (N_17780,N_14895,N_13335);
or U17781 (N_17781,N_15566,N_13939);
nand U17782 (N_17782,N_14939,N_15392);
nand U17783 (N_17783,N_13177,N_15073);
nor U17784 (N_17784,N_15483,N_14493);
nor U17785 (N_17785,N_14743,N_12752);
nor U17786 (N_17786,N_13209,N_14254);
nor U17787 (N_17787,N_15591,N_13986);
nand U17788 (N_17788,N_13279,N_13979);
nor U17789 (N_17789,N_14380,N_13898);
nor U17790 (N_17790,N_14404,N_14987);
and U17791 (N_17791,N_12634,N_13696);
nand U17792 (N_17792,N_14031,N_14602);
nand U17793 (N_17793,N_14559,N_12924);
nor U17794 (N_17794,N_15097,N_13050);
and U17795 (N_17795,N_13096,N_15041);
nor U17796 (N_17796,N_14435,N_14860);
nor U17797 (N_17797,N_15406,N_12603);
and U17798 (N_17798,N_12780,N_13181);
nand U17799 (N_17799,N_13769,N_15171);
nor U17800 (N_17800,N_14221,N_14696);
and U17801 (N_17801,N_14989,N_14304);
xnor U17802 (N_17802,N_12948,N_13442);
and U17803 (N_17803,N_13517,N_14496);
nand U17804 (N_17804,N_13474,N_15439);
xor U17805 (N_17805,N_12829,N_13511);
and U17806 (N_17806,N_13232,N_15280);
and U17807 (N_17807,N_14620,N_14199);
xor U17808 (N_17808,N_14045,N_14873);
or U17809 (N_17809,N_13035,N_13592);
nand U17810 (N_17810,N_15513,N_13817);
xor U17811 (N_17811,N_13237,N_12620);
nand U17812 (N_17812,N_14162,N_14057);
or U17813 (N_17813,N_14468,N_14705);
or U17814 (N_17814,N_14004,N_14143);
nor U17815 (N_17815,N_14751,N_13822);
or U17816 (N_17816,N_13950,N_13976);
nand U17817 (N_17817,N_14841,N_13428);
xnor U17818 (N_17818,N_13675,N_15278);
or U17819 (N_17819,N_13418,N_15075);
nand U17820 (N_17820,N_14097,N_14509);
nand U17821 (N_17821,N_12692,N_13256);
nor U17822 (N_17822,N_15068,N_15035);
or U17823 (N_17823,N_14872,N_13894);
nor U17824 (N_17824,N_13677,N_14161);
and U17825 (N_17825,N_15542,N_13660);
or U17826 (N_17826,N_15521,N_14357);
nor U17827 (N_17827,N_13769,N_14905);
nand U17828 (N_17828,N_14325,N_13881);
and U17829 (N_17829,N_13333,N_12604);
nand U17830 (N_17830,N_14591,N_13498);
nand U17831 (N_17831,N_15243,N_12667);
nor U17832 (N_17832,N_13031,N_15411);
xnor U17833 (N_17833,N_15468,N_15031);
or U17834 (N_17834,N_15306,N_14225);
xnor U17835 (N_17835,N_12829,N_13732);
nor U17836 (N_17836,N_15344,N_13774);
nor U17837 (N_17837,N_13955,N_14502);
nand U17838 (N_17838,N_15125,N_12698);
and U17839 (N_17839,N_13962,N_13156);
or U17840 (N_17840,N_14138,N_12511);
and U17841 (N_17841,N_13117,N_14318);
or U17842 (N_17842,N_15432,N_12705);
or U17843 (N_17843,N_13503,N_13234);
nand U17844 (N_17844,N_14754,N_15555);
nor U17845 (N_17845,N_14086,N_13746);
nor U17846 (N_17846,N_15466,N_14786);
nand U17847 (N_17847,N_15001,N_12804);
and U17848 (N_17848,N_15599,N_15541);
nor U17849 (N_17849,N_15193,N_13338);
nand U17850 (N_17850,N_12896,N_12736);
nor U17851 (N_17851,N_13399,N_15217);
nand U17852 (N_17852,N_13362,N_15346);
xnor U17853 (N_17853,N_14599,N_14603);
nand U17854 (N_17854,N_13151,N_13756);
or U17855 (N_17855,N_14632,N_13384);
xor U17856 (N_17856,N_12526,N_14380);
and U17857 (N_17857,N_12951,N_13654);
nor U17858 (N_17858,N_15550,N_12662);
or U17859 (N_17859,N_14921,N_15548);
nor U17860 (N_17860,N_12695,N_12779);
nor U17861 (N_17861,N_13929,N_15330);
nor U17862 (N_17862,N_15068,N_15554);
nor U17863 (N_17863,N_14311,N_15079);
nand U17864 (N_17864,N_13625,N_13924);
xnor U17865 (N_17865,N_13594,N_12953);
xor U17866 (N_17866,N_13716,N_13314);
or U17867 (N_17867,N_14423,N_15366);
xor U17868 (N_17868,N_14646,N_14403);
xnor U17869 (N_17869,N_12624,N_13788);
or U17870 (N_17870,N_13045,N_15157);
or U17871 (N_17871,N_15307,N_15568);
nor U17872 (N_17872,N_13642,N_13208);
nand U17873 (N_17873,N_14054,N_15579);
nand U17874 (N_17874,N_13212,N_12696);
and U17875 (N_17875,N_14424,N_15176);
or U17876 (N_17876,N_13682,N_12634);
nand U17877 (N_17877,N_13518,N_14723);
and U17878 (N_17878,N_13254,N_15044);
nor U17879 (N_17879,N_13594,N_14352);
or U17880 (N_17880,N_14858,N_14587);
and U17881 (N_17881,N_14090,N_13765);
xor U17882 (N_17882,N_14101,N_13167);
or U17883 (N_17883,N_13665,N_15464);
nand U17884 (N_17884,N_14720,N_14222);
nand U17885 (N_17885,N_12881,N_12772);
xnor U17886 (N_17886,N_15415,N_12507);
or U17887 (N_17887,N_14194,N_13748);
or U17888 (N_17888,N_15505,N_14704);
xnor U17889 (N_17889,N_13426,N_13466);
nand U17890 (N_17890,N_15026,N_12608);
nand U17891 (N_17891,N_15449,N_13434);
and U17892 (N_17892,N_13276,N_15351);
or U17893 (N_17893,N_13971,N_14495);
or U17894 (N_17894,N_12856,N_12933);
nor U17895 (N_17895,N_14808,N_15434);
xnor U17896 (N_17896,N_13802,N_14049);
nor U17897 (N_17897,N_14860,N_12549);
nand U17898 (N_17898,N_14523,N_13189);
xnor U17899 (N_17899,N_12648,N_15508);
nor U17900 (N_17900,N_14816,N_15445);
nand U17901 (N_17901,N_15578,N_13931);
xor U17902 (N_17902,N_13767,N_14101);
or U17903 (N_17903,N_15404,N_13180);
or U17904 (N_17904,N_13926,N_14870);
nand U17905 (N_17905,N_12738,N_13588);
and U17906 (N_17906,N_14178,N_13119);
or U17907 (N_17907,N_15488,N_15540);
nor U17908 (N_17908,N_14504,N_13981);
and U17909 (N_17909,N_14525,N_14211);
or U17910 (N_17910,N_14971,N_13952);
nand U17911 (N_17911,N_13578,N_15034);
xnor U17912 (N_17912,N_14285,N_12726);
xnor U17913 (N_17913,N_15208,N_13786);
nor U17914 (N_17914,N_14799,N_13513);
xor U17915 (N_17915,N_14026,N_13239);
nor U17916 (N_17916,N_15616,N_13287);
xor U17917 (N_17917,N_13736,N_14062);
nor U17918 (N_17918,N_15607,N_15573);
and U17919 (N_17919,N_15048,N_13999);
nor U17920 (N_17920,N_14453,N_14877);
xor U17921 (N_17921,N_12899,N_14167);
nor U17922 (N_17922,N_14508,N_15332);
or U17923 (N_17923,N_14445,N_14562);
and U17924 (N_17924,N_14967,N_15295);
and U17925 (N_17925,N_12954,N_14861);
nand U17926 (N_17926,N_14930,N_13079);
or U17927 (N_17927,N_13178,N_13466);
nor U17928 (N_17928,N_14208,N_14748);
xnor U17929 (N_17929,N_15543,N_13128);
nor U17930 (N_17930,N_14028,N_14247);
xnor U17931 (N_17931,N_13814,N_13185);
xor U17932 (N_17932,N_13486,N_14040);
xnor U17933 (N_17933,N_13433,N_13857);
xor U17934 (N_17934,N_13318,N_14241);
nand U17935 (N_17935,N_13855,N_15446);
nand U17936 (N_17936,N_12655,N_12771);
nand U17937 (N_17937,N_14783,N_14162);
and U17938 (N_17938,N_14635,N_13684);
nor U17939 (N_17939,N_14108,N_14812);
and U17940 (N_17940,N_14235,N_13242);
nand U17941 (N_17941,N_14131,N_13046);
nor U17942 (N_17942,N_13313,N_14697);
nor U17943 (N_17943,N_14262,N_15222);
or U17944 (N_17944,N_13639,N_14269);
and U17945 (N_17945,N_15287,N_14989);
or U17946 (N_17946,N_13382,N_13368);
or U17947 (N_17947,N_12556,N_12650);
xor U17948 (N_17948,N_15155,N_14395);
nor U17949 (N_17949,N_15256,N_13851);
nand U17950 (N_17950,N_13733,N_14805);
and U17951 (N_17951,N_15159,N_14851);
nor U17952 (N_17952,N_14603,N_13636);
and U17953 (N_17953,N_13310,N_13108);
nor U17954 (N_17954,N_13732,N_13106);
and U17955 (N_17955,N_14743,N_14974);
nor U17956 (N_17956,N_14598,N_15199);
nor U17957 (N_17957,N_14001,N_12829);
xor U17958 (N_17958,N_14821,N_15013);
nor U17959 (N_17959,N_12956,N_13693);
and U17960 (N_17960,N_12662,N_14482);
xnor U17961 (N_17961,N_13147,N_12948);
or U17962 (N_17962,N_15319,N_13955);
xnor U17963 (N_17963,N_14421,N_13400);
nor U17964 (N_17964,N_15343,N_12571);
and U17965 (N_17965,N_12730,N_13597);
or U17966 (N_17966,N_15312,N_15272);
xor U17967 (N_17967,N_15063,N_15453);
nor U17968 (N_17968,N_15089,N_14755);
nor U17969 (N_17969,N_12779,N_13900);
nor U17970 (N_17970,N_12851,N_15134);
or U17971 (N_17971,N_14990,N_14738);
or U17972 (N_17972,N_13742,N_15621);
xor U17973 (N_17973,N_12917,N_15282);
or U17974 (N_17974,N_12839,N_12746);
nand U17975 (N_17975,N_14832,N_14868);
or U17976 (N_17976,N_12588,N_13401);
nor U17977 (N_17977,N_14590,N_15476);
nor U17978 (N_17978,N_15201,N_13834);
or U17979 (N_17979,N_13091,N_13205);
xnor U17980 (N_17980,N_13726,N_13967);
xor U17981 (N_17981,N_14574,N_14493);
xor U17982 (N_17982,N_14427,N_13428);
and U17983 (N_17983,N_15326,N_15435);
xor U17984 (N_17984,N_13694,N_13099);
and U17985 (N_17985,N_12853,N_12773);
nand U17986 (N_17986,N_13280,N_14499);
nor U17987 (N_17987,N_14231,N_12704);
xnor U17988 (N_17988,N_15205,N_13400);
and U17989 (N_17989,N_12855,N_13322);
nor U17990 (N_17990,N_12940,N_15455);
and U17991 (N_17991,N_15222,N_13417);
xor U17992 (N_17992,N_12955,N_13797);
nand U17993 (N_17993,N_12965,N_14841);
xor U17994 (N_17994,N_14934,N_14575);
or U17995 (N_17995,N_12633,N_14843);
nand U17996 (N_17996,N_13792,N_14331);
nor U17997 (N_17997,N_14449,N_14729);
nor U17998 (N_17998,N_12924,N_14718);
nand U17999 (N_17999,N_13445,N_15346);
nor U18000 (N_18000,N_12760,N_13284);
or U18001 (N_18001,N_13956,N_14110);
xor U18002 (N_18002,N_14858,N_14063);
and U18003 (N_18003,N_14795,N_14688);
xor U18004 (N_18004,N_14363,N_15617);
or U18005 (N_18005,N_13998,N_13723);
nor U18006 (N_18006,N_13801,N_14698);
nor U18007 (N_18007,N_13295,N_12653);
or U18008 (N_18008,N_13233,N_13966);
nor U18009 (N_18009,N_12658,N_13222);
xor U18010 (N_18010,N_14180,N_14251);
and U18011 (N_18011,N_15137,N_12849);
xnor U18012 (N_18012,N_13350,N_14676);
and U18013 (N_18013,N_12617,N_15623);
nand U18014 (N_18014,N_15159,N_13540);
nand U18015 (N_18015,N_15262,N_13381);
and U18016 (N_18016,N_15588,N_13931);
nor U18017 (N_18017,N_14671,N_14794);
or U18018 (N_18018,N_13336,N_15474);
and U18019 (N_18019,N_12534,N_15029);
or U18020 (N_18020,N_13823,N_13827);
nand U18021 (N_18021,N_13028,N_13560);
xor U18022 (N_18022,N_15607,N_14065);
and U18023 (N_18023,N_12739,N_15120);
nand U18024 (N_18024,N_15216,N_12720);
nand U18025 (N_18025,N_12867,N_13015);
nand U18026 (N_18026,N_13983,N_15114);
or U18027 (N_18027,N_15156,N_14253);
nor U18028 (N_18028,N_13647,N_15001);
and U18029 (N_18029,N_12884,N_13881);
or U18030 (N_18030,N_13718,N_13117);
nor U18031 (N_18031,N_13163,N_14345);
and U18032 (N_18032,N_12890,N_13806);
nand U18033 (N_18033,N_13602,N_13673);
xor U18034 (N_18034,N_13044,N_12899);
or U18035 (N_18035,N_13277,N_13324);
or U18036 (N_18036,N_13525,N_13618);
xor U18037 (N_18037,N_13238,N_12721);
nor U18038 (N_18038,N_15356,N_14250);
nor U18039 (N_18039,N_12814,N_14965);
nand U18040 (N_18040,N_13918,N_13572);
xnor U18041 (N_18041,N_13193,N_13678);
xnor U18042 (N_18042,N_15488,N_14446);
and U18043 (N_18043,N_15033,N_15570);
xor U18044 (N_18044,N_12564,N_13639);
nand U18045 (N_18045,N_15554,N_15155);
or U18046 (N_18046,N_14830,N_14288);
nor U18047 (N_18047,N_13455,N_13166);
and U18048 (N_18048,N_15197,N_13108);
nor U18049 (N_18049,N_15220,N_15127);
nor U18050 (N_18050,N_15068,N_13252);
nor U18051 (N_18051,N_13370,N_14064);
xor U18052 (N_18052,N_14761,N_12868);
xor U18053 (N_18053,N_14755,N_14026);
xnor U18054 (N_18054,N_13303,N_14021);
and U18055 (N_18055,N_15141,N_14326);
nand U18056 (N_18056,N_15092,N_14591);
nand U18057 (N_18057,N_12732,N_12690);
nor U18058 (N_18058,N_12946,N_14177);
xor U18059 (N_18059,N_15209,N_13750);
xnor U18060 (N_18060,N_14764,N_14951);
xor U18061 (N_18061,N_12509,N_12991);
nand U18062 (N_18062,N_12994,N_14628);
or U18063 (N_18063,N_13221,N_12877);
nand U18064 (N_18064,N_14601,N_14817);
and U18065 (N_18065,N_14066,N_13380);
xor U18066 (N_18066,N_15469,N_12988);
and U18067 (N_18067,N_14181,N_14880);
nand U18068 (N_18068,N_13703,N_13668);
or U18069 (N_18069,N_15423,N_13451);
or U18070 (N_18070,N_13032,N_13651);
nand U18071 (N_18071,N_13598,N_13325);
xnor U18072 (N_18072,N_12851,N_15354);
and U18073 (N_18073,N_14597,N_14510);
xor U18074 (N_18074,N_15214,N_13763);
xor U18075 (N_18075,N_14268,N_13615);
and U18076 (N_18076,N_13775,N_15101);
or U18077 (N_18077,N_14317,N_15005);
xnor U18078 (N_18078,N_13983,N_12865);
or U18079 (N_18079,N_13423,N_13345);
xnor U18080 (N_18080,N_14362,N_14988);
or U18081 (N_18081,N_14790,N_13183);
or U18082 (N_18082,N_12667,N_14513);
nand U18083 (N_18083,N_12941,N_12555);
xnor U18084 (N_18084,N_14039,N_13643);
nor U18085 (N_18085,N_15056,N_12784);
xnor U18086 (N_18086,N_14559,N_13970);
xor U18087 (N_18087,N_13291,N_13403);
and U18088 (N_18088,N_15463,N_15336);
nor U18089 (N_18089,N_15530,N_15398);
or U18090 (N_18090,N_13766,N_13725);
and U18091 (N_18091,N_14493,N_13837);
xor U18092 (N_18092,N_14068,N_14126);
nand U18093 (N_18093,N_15197,N_13732);
or U18094 (N_18094,N_14363,N_13579);
or U18095 (N_18095,N_13309,N_14531);
and U18096 (N_18096,N_12685,N_14996);
or U18097 (N_18097,N_14525,N_15535);
and U18098 (N_18098,N_15151,N_14877);
xnor U18099 (N_18099,N_14445,N_15292);
xor U18100 (N_18100,N_14311,N_15320);
nor U18101 (N_18101,N_14070,N_12660);
nor U18102 (N_18102,N_14152,N_13351);
or U18103 (N_18103,N_12736,N_12766);
or U18104 (N_18104,N_13019,N_13971);
or U18105 (N_18105,N_15335,N_13739);
nor U18106 (N_18106,N_12721,N_14928);
nand U18107 (N_18107,N_14489,N_13803);
or U18108 (N_18108,N_15478,N_14321);
nor U18109 (N_18109,N_14352,N_13522);
and U18110 (N_18110,N_14334,N_13762);
nor U18111 (N_18111,N_14057,N_14158);
xnor U18112 (N_18112,N_13837,N_15349);
nand U18113 (N_18113,N_15594,N_14285);
nand U18114 (N_18114,N_14081,N_14604);
nand U18115 (N_18115,N_13964,N_14571);
nor U18116 (N_18116,N_12913,N_13590);
nor U18117 (N_18117,N_13015,N_14230);
nor U18118 (N_18118,N_13968,N_12580);
nor U18119 (N_18119,N_14167,N_14874);
nand U18120 (N_18120,N_14484,N_12872);
nand U18121 (N_18121,N_15569,N_15127);
nor U18122 (N_18122,N_15115,N_12903);
nor U18123 (N_18123,N_13076,N_13477);
or U18124 (N_18124,N_12914,N_14114);
or U18125 (N_18125,N_14631,N_13277);
or U18126 (N_18126,N_13002,N_14257);
and U18127 (N_18127,N_14010,N_15588);
nand U18128 (N_18128,N_13776,N_14876);
xor U18129 (N_18129,N_12933,N_15120);
xor U18130 (N_18130,N_12915,N_13035);
and U18131 (N_18131,N_14391,N_13416);
and U18132 (N_18132,N_13463,N_15578);
or U18133 (N_18133,N_14233,N_14424);
and U18134 (N_18134,N_12790,N_13463);
and U18135 (N_18135,N_12537,N_14546);
nand U18136 (N_18136,N_14258,N_14423);
and U18137 (N_18137,N_14588,N_14260);
and U18138 (N_18138,N_14996,N_13249);
nor U18139 (N_18139,N_12957,N_14058);
or U18140 (N_18140,N_12704,N_15512);
xnor U18141 (N_18141,N_15229,N_14568);
nand U18142 (N_18142,N_15192,N_15145);
or U18143 (N_18143,N_13712,N_12896);
or U18144 (N_18144,N_12564,N_12578);
xnor U18145 (N_18145,N_13390,N_14630);
nor U18146 (N_18146,N_13494,N_13902);
nor U18147 (N_18147,N_12800,N_12804);
nor U18148 (N_18148,N_14391,N_13019);
or U18149 (N_18149,N_13195,N_15473);
nand U18150 (N_18150,N_13018,N_15615);
nor U18151 (N_18151,N_12595,N_14882);
nor U18152 (N_18152,N_14046,N_15294);
xnor U18153 (N_18153,N_13913,N_13492);
nand U18154 (N_18154,N_15153,N_15456);
nand U18155 (N_18155,N_14509,N_14471);
or U18156 (N_18156,N_14025,N_12790);
nand U18157 (N_18157,N_13177,N_14159);
xnor U18158 (N_18158,N_13917,N_13433);
nand U18159 (N_18159,N_13596,N_14997);
and U18160 (N_18160,N_13761,N_15010);
nor U18161 (N_18161,N_13392,N_15251);
nor U18162 (N_18162,N_15215,N_12686);
and U18163 (N_18163,N_12667,N_14212);
xnor U18164 (N_18164,N_12606,N_13821);
xor U18165 (N_18165,N_13645,N_14108);
and U18166 (N_18166,N_14317,N_12583);
or U18167 (N_18167,N_12736,N_15335);
and U18168 (N_18168,N_15120,N_14138);
nor U18169 (N_18169,N_15507,N_12542);
nand U18170 (N_18170,N_14634,N_13112);
nand U18171 (N_18171,N_13240,N_14373);
nand U18172 (N_18172,N_13592,N_15512);
xnor U18173 (N_18173,N_14271,N_13515);
nor U18174 (N_18174,N_13769,N_14928);
nand U18175 (N_18175,N_14264,N_13844);
xor U18176 (N_18176,N_12911,N_14832);
xnor U18177 (N_18177,N_13764,N_12635);
or U18178 (N_18178,N_14767,N_12927);
nand U18179 (N_18179,N_15274,N_12746);
and U18180 (N_18180,N_12595,N_14389);
and U18181 (N_18181,N_14465,N_13247);
nand U18182 (N_18182,N_13647,N_15333);
nand U18183 (N_18183,N_13534,N_13783);
or U18184 (N_18184,N_12555,N_13997);
and U18185 (N_18185,N_13076,N_13767);
nand U18186 (N_18186,N_15462,N_15119);
and U18187 (N_18187,N_13906,N_12987);
xor U18188 (N_18188,N_14164,N_13209);
nand U18189 (N_18189,N_15563,N_13187);
or U18190 (N_18190,N_15144,N_14731);
or U18191 (N_18191,N_15547,N_14329);
and U18192 (N_18192,N_14161,N_14704);
or U18193 (N_18193,N_12707,N_14932);
nor U18194 (N_18194,N_13142,N_14395);
and U18195 (N_18195,N_14840,N_12691);
nor U18196 (N_18196,N_14749,N_14436);
or U18197 (N_18197,N_12739,N_14158);
and U18198 (N_18198,N_14876,N_14450);
xnor U18199 (N_18199,N_13131,N_15244);
nor U18200 (N_18200,N_13781,N_12705);
nor U18201 (N_18201,N_15375,N_14459);
nand U18202 (N_18202,N_14435,N_13256);
or U18203 (N_18203,N_14603,N_14704);
nor U18204 (N_18204,N_13347,N_15556);
nor U18205 (N_18205,N_13690,N_12917);
xor U18206 (N_18206,N_12593,N_14186);
nor U18207 (N_18207,N_13470,N_14220);
nor U18208 (N_18208,N_14048,N_14844);
xor U18209 (N_18209,N_12685,N_15445);
or U18210 (N_18210,N_12911,N_14687);
nor U18211 (N_18211,N_15451,N_13895);
nor U18212 (N_18212,N_13110,N_12915);
and U18213 (N_18213,N_14767,N_12595);
and U18214 (N_18214,N_12747,N_15400);
xor U18215 (N_18215,N_13337,N_14854);
or U18216 (N_18216,N_12698,N_13146);
xor U18217 (N_18217,N_14611,N_15010);
xor U18218 (N_18218,N_12877,N_14388);
nand U18219 (N_18219,N_13648,N_13045);
nand U18220 (N_18220,N_13038,N_15289);
and U18221 (N_18221,N_13446,N_15240);
and U18222 (N_18222,N_13770,N_12853);
and U18223 (N_18223,N_12561,N_13829);
nor U18224 (N_18224,N_14370,N_14926);
nand U18225 (N_18225,N_13384,N_13120);
nand U18226 (N_18226,N_13682,N_15065);
xor U18227 (N_18227,N_12970,N_14215);
xor U18228 (N_18228,N_12616,N_15237);
or U18229 (N_18229,N_13136,N_15325);
nand U18230 (N_18230,N_12780,N_13828);
or U18231 (N_18231,N_15615,N_15324);
and U18232 (N_18232,N_12649,N_12902);
nor U18233 (N_18233,N_15250,N_14583);
or U18234 (N_18234,N_14408,N_14314);
xor U18235 (N_18235,N_14962,N_13658);
or U18236 (N_18236,N_13112,N_15467);
xor U18237 (N_18237,N_13406,N_13941);
xnor U18238 (N_18238,N_12663,N_13546);
nand U18239 (N_18239,N_12736,N_15000);
nand U18240 (N_18240,N_13699,N_14545);
and U18241 (N_18241,N_13752,N_13422);
and U18242 (N_18242,N_14730,N_15004);
or U18243 (N_18243,N_14065,N_14690);
nor U18244 (N_18244,N_15196,N_15092);
nor U18245 (N_18245,N_12583,N_14374);
nand U18246 (N_18246,N_13319,N_14156);
xor U18247 (N_18247,N_12917,N_15173);
nand U18248 (N_18248,N_13479,N_13645);
nand U18249 (N_18249,N_14392,N_13704);
nand U18250 (N_18250,N_14965,N_14907);
and U18251 (N_18251,N_14224,N_15340);
xnor U18252 (N_18252,N_13950,N_14097);
and U18253 (N_18253,N_14223,N_15247);
nand U18254 (N_18254,N_13094,N_13446);
xnor U18255 (N_18255,N_12861,N_12846);
nor U18256 (N_18256,N_13612,N_13754);
xnor U18257 (N_18257,N_13160,N_14404);
and U18258 (N_18258,N_15014,N_14641);
nand U18259 (N_18259,N_13811,N_15402);
or U18260 (N_18260,N_14721,N_14583);
or U18261 (N_18261,N_14532,N_14358);
or U18262 (N_18262,N_12864,N_13603);
and U18263 (N_18263,N_13266,N_13228);
nand U18264 (N_18264,N_12947,N_14881);
or U18265 (N_18265,N_13514,N_14625);
or U18266 (N_18266,N_14510,N_15357);
xnor U18267 (N_18267,N_14850,N_13872);
xnor U18268 (N_18268,N_15520,N_12761);
nand U18269 (N_18269,N_15068,N_14747);
nor U18270 (N_18270,N_15029,N_13150);
or U18271 (N_18271,N_15436,N_12859);
and U18272 (N_18272,N_14106,N_13081);
xor U18273 (N_18273,N_15462,N_15581);
or U18274 (N_18274,N_13934,N_14925);
nor U18275 (N_18275,N_13422,N_13664);
nand U18276 (N_18276,N_12644,N_15060);
or U18277 (N_18277,N_12787,N_13332);
nor U18278 (N_18278,N_13596,N_15412);
xor U18279 (N_18279,N_13940,N_14845);
and U18280 (N_18280,N_14467,N_15109);
nand U18281 (N_18281,N_14832,N_14843);
or U18282 (N_18282,N_14813,N_14784);
and U18283 (N_18283,N_14102,N_13784);
nor U18284 (N_18284,N_15617,N_14290);
nand U18285 (N_18285,N_13577,N_13166);
nand U18286 (N_18286,N_12938,N_15379);
nand U18287 (N_18287,N_12878,N_15025);
and U18288 (N_18288,N_13409,N_12655);
nor U18289 (N_18289,N_14381,N_14345);
nand U18290 (N_18290,N_13099,N_13236);
and U18291 (N_18291,N_15435,N_13133);
xnor U18292 (N_18292,N_15290,N_14140);
nand U18293 (N_18293,N_12946,N_14564);
nand U18294 (N_18294,N_13233,N_14353);
nor U18295 (N_18295,N_14095,N_13360);
xnor U18296 (N_18296,N_14130,N_13961);
and U18297 (N_18297,N_13854,N_13115);
nand U18298 (N_18298,N_12926,N_15261);
xor U18299 (N_18299,N_14194,N_14197);
or U18300 (N_18300,N_14280,N_14666);
xor U18301 (N_18301,N_14922,N_14020);
nor U18302 (N_18302,N_12795,N_15542);
nor U18303 (N_18303,N_13335,N_15243);
and U18304 (N_18304,N_14537,N_12638);
and U18305 (N_18305,N_14512,N_14761);
xor U18306 (N_18306,N_14553,N_12892);
nand U18307 (N_18307,N_13118,N_12855);
nor U18308 (N_18308,N_12925,N_14164);
and U18309 (N_18309,N_15142,N_12502);
or U18310 (N_18310,N_14931,N_13809);
and U18311 (N_18311,N_13826,N_12860);
and U18312 (N_18312,N_13017,N_12927);
or U18313 (N_18313,N_14074,N_14293);
or U18314 (N_18314,N_14302,N_13515);
or U18315 (N_18315,N_12940,N_13147);
xor U18316 (N_18316,N_15512,N_12697);
or U18317 (N_18317,N_13658,N_13001);
or U18318 (N_18318,N_15359,N_13469);
or U18319 (N_18319,N_12554,N_14795);
xor U18320 (N_18320,N_13599,N_14809);
and U18321 (N_18321,N_15455,N_14474);
xor U18322 (N_18322,N_14523,N_14589);
nor U18323 (N_18323,N_13734,N_14125);
and U18324 (N_18324,N_15090,N_13570);
nand U18325 (N_18325,N_13887,N_13297);
or U18326 (N_18326,N_13271,N_12680);
and U18327 (N_18327,N_13460,N_14144);
nand U18328 (N_18328,N_13947,N_13855);
or U18329 (N_18329,N_15368,N_13991);
nand U18330 (N_18330,N_13930,N_14279);
xor U18331 (N_18331,N_13716,N_13201);
nand U18332 (N_18332,N_13498,N_13981);
nand U18333 (N_18333,N_13691,N_15138);
and U18334 (N_18334,N_15308,N_12608);
nor U18335 (N_18335,N_13653,N_14888);
xnor U18336 (N_18336,N_14789,N_13573);
and U18337 (N_18337,N_12857,N_15244);
and U18338 (N_18338,N_15509,N_12577);
or U18339 (N_18339,N_13433,N_14597);
or U18340 (N_18340,N_13130,N_14056);
nor U18341 (N_18341,N_12622,N_14097);
nor U18342 (N_18342,N_14000,N_15316);
and U18343 (N_18343,N_12899,N_14204);
xor U18344 (N_18344,N_12964,N_14617);
or U18345 (N_18345,N_14599,N_14967);
xnor U18346 (N_18346,N_15017,N_13983);
xnor U18347 (N_18347,N_15616,N_14042);
or U18348 (N_18348,N_13487,N_14238);
nor U18349 (N_18349,N_15618,N_12522);
or U18350 (N_18350,N_13205,N_12771);
or U18351 (N_18351,N_15287,N_13528);
xnor U18352 (N_18352,N_12835,N_15448);
and U18353 (N_18353,N_15604,N_12630);
and U18354 (N_18354,N_13275,N_13544);
and U18355 (N_18355,N_13408,N_12506);
nand U18356 (N_18356,N_14129,N_14782);
xnor U18357 (N_18357,N_15602,N_15185);
or U18358 (N_18358,N_15099,N_15330);
nor U18359 (N_18359,N_12798,N_15303);
or U18360 (N_18360,N_14456,N_15288);
nand U18361 (N_18361,N_15159,N_13822);
and U18362 (N_18362,N_13906,N_14671);
xnor U18363 (N_18363,N_13687,N_14372);
xnor U18364 (N_18364,N_13670,N_14984);
and U18365 (N_18365,N_14087,N_14665);
or U18366 (N_18366,N_14583,N_14710);
or U18367 (N_18367,N_13971,N_13065);
or U18368 (N_18368,N_12956,N_14378);
xnor U18369 (N_18369,N_13417,N_13312);
nor U18370 (N_18370,N_13160,N_14224);
nor U18371 (N_18371,N_14314,N_13493);
xnor U18372 (N_18372,N_14427,N_14638);
or U18373 (N_18373,N_14903,N_14216);
xnor U18374 (N_18374,N_14323,N_12607);
xor U18375 (N_18375,N_12638,N_14314);
nand U18376 (N_18376,N_14972,N_12752);
nand U18377 (N_18377,N_15096,N_15570);
and U18378 (N_18378,N_12900,N_15420);
or U18379 (N_18379,N_15334,N_15560);
and U18380 (N_18380,N_12509,N_15455);
nand U18381 (N_18381,N_12500,N_13644);
nand U18382 (N_18382,N_12529,N_12941);
xnor U18383 (N_18383,N_14655,N_13455);
nand U18384 (N_18384,N_15186,N_14970);
xnor U18385 (N_18385,N_13061,N_13950);
or U18386 (N_18386,N_15495,N_14409);
xnor U18387 (N_18387,N_13704,N_14099);
or U18388 (N_18388,N_14952,N_14148);
nor U18389 (N_18389,N_13224,N_13421);
nand U18390 (N_18390,N_14301,N_14135);
nor U18391 (N_18391,N_13365,N_12567);
xor U18392 (N_18392,N_14528,N_14334);
xnor U18393 (N_18393,N_12536,N_12628);
nand U18394 (N_18394,N_12796,N_14558);
xor U18395 (N_18395,N_14671,N_13134);
nand U18396 (N_18396,N_12940,N_14750);
nand U18397 (N_18397,N_13179,N_13339);
nor U18398 (N_18398,N_13953,N_14865);
and U18399 (N_18399,N_13660,N_15197);
xnor U18400 (N_18400,N_14162,N_12584);
and U18401 (N_18401,N_12855,N_15568);
nand U18402 (N_18402,N_14737,N_12846);
nand U18403 (N_18403,N_14823,N_12897);
nor U18404 (N_18404,N_15263,N_15291);
and U18405 (N_18405,N_15336,N_14967);
and U18406 (N_18406,N_13815,N_15079);
xor U18407 (N_18407,N_12639,N_12899);
nand U18408 (N_18408,N_13979,N_13225);
nand U18409 (N_18409,N_14614,N_15443);
nor U18410 (N_18410,N_14448,N_15465);
and U18411 (N_18411,N_14417,N_14284);
and U18412 (N_18412,N_14133,N_14021);
nand U18413 (N_18413,N_15197,N_13776);
nor U18414 (N_18414,N_14197,N_15272);
and U18415 (N_18415,N_12772,N_12756);
or U18416 (N_18416,N_14412,N_12983);
xnor U18417 (N_18417,N_15334,N_13557);
nand U18418 (N_18418,N_13457,N_15272);
and U18419 (N_18419,N_14392,N_13194);
xnor U18420 (N_18420,N_14919,N_14470);
xnor U18421 (N_18421,N_14148,N_14857);
nand U18422 (N_18422,N_12916,N_13824);
nor U18423 (N_18423,N_13435,N_14815);
nand U18424 (N_18424,N_12899,N_13114);
or U18425 (N_18425,N_14303,N_14518);
nand U18426 (N_18426,N_14475,N_15234);
xnor U18427 (N_18427,N_14947,N_12600);
nand U18428 (N_18428,N_14488,N_12942);
or U18429 (N_18429,N_14057,N_14959);
or U18430 (N_18430,N_13648,N_14408);
nor U18431 (N_18431,N_13896,N_14395);
nand U18432 (N_18432,N_14706,N_13770);
or U18433 (N_18433,N_14000,N_14181);
nor U18434 (N_18434,N_12941,N_13869);
nor U18435 (N_18435,N_14086,N_15533);
nand U18436 (N_18436,N_14035,N_13774);
xor U18437 (N_18437,N_13780,N_15182);
or U18438 (N_18438,N_14686,N_12805);
and U18439 (N_18439,N_12718,N_12816);
and U18440 (N_18440,N_12891,N_12544);
nor U18441 (N_18441,N_14170,N_13353);
nor U18442 (N_18442,N_12940,N_13948);
xor U18443 (N_18443,N_13096,N_13514);
and U18444 (N_18444,N_12796,N_12958);
xnor U18445 (N_18445,N_14095,N_15257);
and U18446 (N_18446,N_13586,N_14838);
or U18447 (N_18447,N_12730,N_13895);
or U18448 (N_18448,N_12987,N_12832);
and U18449 (N_18449,N_13913,N_15278);
or U18450 (N_18450,N_12811,N_15454);
nor U18451 (N_18451,N_13570,N_13723);
nor U18452 (N_18452,N_14205,N_14593);
nor U18453 (N_18453,N_12769,N_15268);
nand U18454 (N_18454,N_14038,N_13004);
and U18455 (N_18455,N_14894,N_14189);
nor U18456 (N_18456,N_15085,N_14801);
xor U18457 (N_18457,N_13934,N_14066);
nand U18458 (N_18458,N_14925,N_14300);
or U18459 (N_18459,N_12631,N_15350);
or U18460 (N_18460,N_14409,N_15446);
nand U18461 (N_18461,N_14913,N_15201);
nand U18462 (N_18462,N_15143,N_15127);
nor U18463 (N_18463,N_12634,N_15190);
nor U18464 (N_18464,N_14819,N_14656);
and U18465 (N_18465,N_15434,N_12708);
nand U18466 (N_18466,N_14352,N_12827);
or U18467 (N_18467,N_15010,N_13184);
xnor U18468 (N_18468,N_14295,N_14148);
or U18469 (N_18469,N_12716,N_14928);
nand U18470 (N_18470,N_12685,N_12865);
xnor U18471 (N_18471,N_13489,N_14058);
nand U18472 (N_18472,N_13606,N_13117);
xnor U18473 (N_18473,N_14842,N_14412);
nand U18474 (N_18474,N_12564,N_12876);
xnor U18475 (N_18475,N_13926,N_15444);
nor U18476 (N_18476,N_12571,N_14757);
nor U18477 (N_18477,N_13850,N_14245);
xor U18478 (N_18478,N_15306,N_13902);
xnor U18479 (N_18479,N_12816,N_14616);
and U18480 (N_18480,N_14044,N_14892);
nand U18481 (N_18481,N_14125,N_14126);
or U18482 (N_18482,N_12745,N_14611);
and U18483 (N_18483,N_13373,N_15352);
or U18484 (N_18484,N_12982,N_13758);
and U18485 (N_18485,N_12683,N_14670);
or U18486 (N_18486,N_13508,N_14820);
and U18487 (N_18487,N_13780,N_14154);
or U18488 (N_18488,N_13267,N_14753);
nor U18489 (N_18489,N_15144,N_13261);
nand U18490 (N_18490,N_13646,N_14771);
and U18491 (N_18491,N_13767,N_12517);
or U18492 (N_18492,N_14804,N_13958);
nand U18493 (N_18493,N_13632,N_13339);
and U18494 (N_18494,N_12675,N_13641);
xor U18495 (N_18495,N_13385,N_13839);
nand U18496 (N_18496,N_15094,N_13392);
and U18497 (N_18497,N_14965,N_14732);
nor U18498 (N_18498,N_13345,N_13013);
or U18499 (N_18499,N_12819,N_12885);
or U18500 (N_18500,N_13613,N_15364);
nor U18501 (N_18501,N_14423,N_15393);
xnor U18502 (N_18502,N_15266,N_15254);
xnor U18503 (N_18503,N_15412,N_13921);
xor U18504 (N_18504,N_15125,N_14140);
xnor U18505 (N_18505,N_12550,N_14135);
and U18506 (N_18506,N_12968,N_12845);
nand U18507 (N_18507,N_13609,N_14915);
or U18508 (N_18508,N_13883,N_12913);
nand U18509 (N_18509,N_15178,N_15332);
nor U18510 (N_18510,N_13163,N_13810);
xnor U18511 (N_18511,N_15216,N_14273);
xnor U18512 (N_18512,N_15111,N_15580);
nor U18513 (N_18513,N_14047,N_15039);
or U18514 (N_18514,N_12511,N_14607);
nand U18515 (N_18515,N_13307,N_14523);
or U18516 (N_18516,N_14045,N_15476);
and U18517 (N_18517,N_13591,N_14937);
or U18518 (N_18518,N_14230,N_13408);
nor U18519 (N_18519,N_14400,N_13079);
and U18520 (N_18520,N_12695,N_13007);
or U18521 (N_18521,N_14107,N_14058);
xor U18522 (N_18522,N_13223,N_12933);
nor U18523 (N_18523,N_14147,N_14625);
and U18524 (N_18524,N_12718,N_15288);
or U18525 (N_18525,N_14093,N_14341);
nand U18526 (N_18526,N_15388,N_14600);
nand U18527 (N_18527,N_14625,N_15086);
xor U18528 (N_18528,N_14887,N_13417);
nand U18529 (N_18529,N_13379,N_13211);
xnor U18530 (N_18530,N_13272,N_12733);
nand U18531 (N_18531,N_12936,N_14911);
nand U18532 (N_18532,N_13887,N_12601);
xnor U18533 (N_18533,N_13125,N_12782);
nand U18534 (N_18534,N_12831,N_13750);
nand U18535 (N_18535,N_14458,N_15087);
and U18536 (N_18536,N_14197,N_13549);
xnor U18537 (N_18537,N_13256,N_15016);
nor U18538 (N_18538,N_12893,N_15079);
or U18539 (N_18539,N_14375,N_15597);
nor U18540 (N_18540,N_14884,N_12751);
and U18541 (N_18541,N_12568,N_14537);
nand U18542 (N_18542,N_12947,N_13355);
nand U18543 (N_18543,N_14477,N_14897);
or U18544 (N_18544,N_13541,N_15559);
and U18545 (N_18545,N_14748,N_14696);
and U18546 (N_18546,N_13424,N_14914);
nor U18547 (N_18547,N_14834,N_14293);
nor U18548 (N_18548,N_14398,N_13778);
or U18549 (N_18549,N_12797,N_13980);
nor U18550 (N_18550,N_15410,N_15353);
and U18551 (N_18551,N_13752,N_14000);
xor U18552 (N_18552,N_12935,N_15467);
nand U18553 (N_18553,N_13668,N_14357);
or U18554 (N_18554,N_14361,N_15002);
xor U18555 (N_18555,N_13175,N_13311);
and U18556 (N_18556,N_14315,N_15321);
nand U18557 (N_18557,N_14305,N_14132);
and U18558 (N_18558,N_14657,N_12809);
xnor U18559 (N_18559,N_14747,N_13191);
and U18560 (N_18560,N_15222,N_15139);
xnor U18561 (N_18561,N_15335,N_13615);
nand U18562 (N_18562,N_13236,N_14553);
or U18563 (N_18563,N_14059,N_14402);
nor U18564 (N_18564,N_14111,N_14372);
nand U18565 (N_18565,N_15176,N_12709);
or U18566 (N_18566,N_12865,N_12816);
nor U18567 (N_18567,N_14903,N_15529);
and U18568 (N_18568,N_12736,N_13632);
or U18569 (N_18569,N_13712,N_13158);
and U18570 (N_18570,N_13785,N_15580);
or U18571 (N_18571,N_13736,N_15179);
and U18572 (N_18572,N_13363,N_14180);
nand U18573 (N_18573,N_13524,N_15530);
xor U18574 (N_18574,N_13579,N_13954);
or U18575 (N_18575,N_15427,N_12940);
xor U18576 (N_18576,N_15156,N_13357);
nand U18577 (N_18577,N_12508,N_13272);
nand U18578 (N_18578,N_12969,N_12898);
or U18579 (N_18579,N_13381,N_13811);
xnor U18580 (N_18580,N_14145,N_15362);
nor U18581 (N_18581,N_15349,N_13459);
nand U18582 (N_18582,N_15220,N_15079);
nor U18583 (N_18583,N_14468,N_13013);
or U18584 (N_18584,N_14580,N_13612);
or U18585 (N_18585,N_14553,N_14824);
and U18586 (N_18586,N_13464,N_14153);
nor U18587 (N_18587,N_12566,N_13763);
and U18588 (N_18588,N_13815,N_13727);
nand U18589 (N_18589,N_14964,N_14218);
nand U18590 (N_18590,N_13003,N_13956);
nor U18591 (N_18591,N_14478,N_14214);
nand U18592 (N_18592,N_15266,N_13006);
or U18593 (N_18593,N_15044,N_14008);
and U18594 (N_18594,N_13792,N_15236);
and U18595 (N_18595,N_14265,N_12823);
xor U18596 (N_18596,N_13027,N_14113);
or U18597 (N_18597,N_12631,N_12585);
nand U18598 (N_18598,N_13787,N_15096);
nor U18599 (N_18599,N_14551,N_13458);
or U18600 (N_18600,N_12904,N_14432);
nor U18601 (N_18601,N_13508,N_14012);
and U18602 (N_18602,N_14022,N_14609);
or U18603 (N_18603,N_13859,N_14163);
nand U18604 (N_18604,N_13539,N_14406);
nor U18605 (N_18605,N_14136,N_13965);
nor U18606 (N_18606,N_14352,N_14366);
and U18607 (N_18607,N_14451,N_14882);
nor U18608 (N_18608,N_14924,N_15106);
or U18609 (N_18609,N_15143,N_15149);
nor U18610 (N_18610,N_13732,N_15593);
or U18611 (N_18611,N_14650,N_12638);
or U18612 (N_18612,N_13201,N_15163);
nand U18613 (N_18613,N_15169,N_14984);
xnor U18614 (N_18614,N_14136,N_15192);
nand U18615 (N_18615,N_13162,N_15291);
nor U18616 (N_18616,N_15042,N_14216);
nand U18617 (N_18617,N_15583,N_13649);
and U18618 (N_18618,N_13423,N_14796);
xor U18619 (N_18619,N_14224,N_14803);
xnor U18620 (N_18620,N_13092,N_15509);
xnor U18621 (N_18621,N_13627,N_14421);
or U18622 (N_18622,N_14645,N_14594);
and U18623 (N_18623,N_13573,N_15072);
and U18624 (N_18624,N_12814,N_14860);
and U18625 (N_18625,N_14131,N_12594);
and U18626 (N_18626,N_14692,N_15356);
and U18627 (N_18627,N_14710,N_14959);
nor U18628 (N_18628,N_12801,N_12839);
nor U18629 (N_18629,N_14654,N_13823);
and U18630 (N_18630,N_15361,N_15171);
nand U18631 (N_18631,N_13759,N_12605);
or U18632 (N_18632,N_13643,N_13911);
nand U18633 (N_18633,N_15087,N_14876);
or U18634 (N_18634,N_13920,N_14464);
nand U18635 (N_18635,N_14754,N_13229);
and U18636 (N_18636,N_14533,N_13255);
xnor U18637 (N_18637,N_13295,N_12533);
nor U18638 (N_18638,N_14383,N_14713);
nand U18639 (N_18639,N_12904,N_15616);
or U18640 (N_18640,N_13338,N_15382);
and U18641 (N_18641,N_13374,N_15552);
nand U18642 (N_18642,N_13253,N_15506);
and U18643 (N_18643,N_13487,N_14564);
nand U18644 (N_18644,N_15550,N_13371);
nor U18645 (N_18645,N_14289,N_12955);
nor U18646 (N_18646,N_13818,N_12698);
or U18647 (N_18647,N_13832,N_14038);
nand U18648 (N_18648,N_14196,N_12870);
and U18649 (N_18649,N_13369,N_13073);
and U18650 (N_18650,N_14956,N_12942);
nand U18651 (N_18651,N_15180,N_15148);
nand U18652 (N_18652,N_14831,N_14572);
and U18653 (N_18653,N_13433,N_13587);
nand U18654 (N_18654,N_13247,N_14469);
xnor U18655 (N_18655,N_13278,N_14538);
nor U18656 (N_18656,N_14867,N_14672);
nor U18657 (N_18657,N_13138,N_14507);
xor U18658 (N_18658,N_13648,N_14481);
and U18659 (N_18659,N_12848,N_14610);
and U18660 (N_18660,N_15612,N_13347);
nor U18661 (N_18661,N_12634,N_13913);
and U18662 (N_18662,N_12516,N_14253);
xnor U18663 (N_18663,N_14843,N_13507);
nand U18664 (N_18664,N_13791,N_13214);
or U18665 (N_18665,N_12825,N_13771);
or U18666 (N_18666,N_13282,N_14971);
nor U18667 (N_18667,N_15199,N_14891);
nor U18668 (N_18668,N_13105,N_14227);
and U18669 (N_18669,N_14497,N_14511);
or U18670 (N_18670,N_14034,N_15006);
and U18671 (N_18671,N_14891,N_15520);
and U18672 (N_18672,N_14242,N_14717);
xnor U18673 (N_18673,N_13364,N_15448);
and U18674 (N_18674,N_14341,N_13052);
nand U18675 (N_18675,N_14728,N_15223);
xor U18676 (N_18676,N_13567,N_15021);
nand U18677 (N_18677,N_14224,N_13013);
and U18678 (N_18678,N_14553,N_13843);
nand U18679 (N_18679,N_14448,N_15460);
nor U18680 (N_18680,N_13375,N_14780);
and U18681 (N_18681,N_15273,N_13552);
xnor U18682 (N_18682,N_14162,N_14920);
and U18683 (N_18683,N_14031,N_15227);
nor U18684 (N_18684,N_13434,N_13301);
and U18685 (N_18685,N_12804,N_13614);
and U18686 (N_18686,N_15169,N_15535);
and U18687 (N_18687,N_13963,N_14473);
nand U18688 (N_18688,N_13557,N_12833);
or U18689 (N_18689,N_13886,N_13682);
xor U18690 (N_18690,N_14677,N_14407);
xnor U18691 (N_18691,N_14154,N_15080);
and U18692 (N_18692,N_13951,N_14713);
nor U18693 (N_18693,N_13070,N_14886);
nand U18694 (N_18694,N_15122,N_15084);
nand U18695 (N_18695,N_13761,N_12505);
xnor U18696 (N_18696,N_13534,N_14126);
and U18697 (N_18697,N_13653,N_13871);
or U18698 (N_18698,N_15013,N_14378);
and U18699 (N_18699,N_12848,N_14362);
nor U18700 (N_18700,N_15609,N_13561);
nor U18701 (N_18701,N_13594,N_12847);
or U18702 (N_18702,N_14428,N_12706);
nand U18703 (N_18703,N_15018,N_14546);
xor U18704 (N_18704,N_12629,N_15342);
and U18705 (N_18705,N_13735,N_14766);
nor U18706 (N_18706,N_14064,N_13684);
or U18707 (N_18707,N_14064,N_14074);
or U18708 (N_18708,N_13296,N_14169);
xor U18709 (N_18709,N_14817,N_13677);
xor U18710 (N_18710,N_15394,N_12557);
nand U18711 (N_18711,N_15099,N_12793);
or U18712 (N_18712,N_13976,N_13569);
or U18713 (N_18713,N_13203,N_12815);
nand U18714 (N_18714,N_13814,N_15164);
or U18715 (N_18715,N_13106,N_13053);
and U18716 (N_18716,N_14864,N_13298);
nor U18717 (N_18717,N_13970,N_13173);
xnor U18718 (N_18718,N_13241,N_15595);
and U18719 (N_18719,N_15580,N_12848);
or U18720 (N_18720,N_13606,N_14335);
nand U18721 (N_18721,N_14910,N_14907);
or U18722 (N_18722,N_13829,N_14515);
nand U18723 (N_18723,N_14710,N_13809);
or U18724 (N_18724,N_12718,N_14765);
xnor U18725 (N_18725,N_12519,N_13885);
xnor U18726 (N_18726,N_15557,N_13881);
nand U18727 (N_18727,N_12883,N_14295);
nor U18728 (N_18728,N_15613,N_13832);
xnor U18729 (N_18729,N_12663,N_13462);
xnor U18730 (N_18730,N_13106,N_14598);
xnor U18731 (N_18731,N_13271,N_14910);
nor U18732 (N_18732,N_14555,N_13909);
nor U18733 (N_18733,N_12630,N_14053);
and U18734 (N_18734,N_14123,N_15351);
xor U18735 (N_18735,N_13199,N_13670);
nand U18736 (N_18736,N_13436,N_14358);
xor U18737 (N_18737,N_12703,N_13085);
and U18738 (N_18738,N_13794,N_14876);
nor U18739 (N_18739,N_13584,N_12783);
nor U18740 (N_18740,N_13106,N_14654);
or U18741 (N_18741,N_14394,N_13065);
nor U18742 (N_18742,N_14558,N_14737);
nand U18743 (N_18743,N_14422,N_13891);
nand U18744 (N_18744,N_14567,N_13690);
and U18745 (N_18745,N_14788,N_13090);
nor U18746 (N_18746,N_15281,N_12603);
nor U18747 (N_18747,N_14877,N_12693);
and U18748 (N_18748,N_14904,N_15230);
or U18749 (N_18749,N_15379,N_12795);
nor U18750 (N_18750,N_17334,N_16817);
or U18751 (N_18751,N_17706,N_15955);
nor U18752 (N_18752,N_16400,N_15768);
nor U18753 (N_18753,N_16434,N_17109);
xor U18754 (N_18754,N_17506,N_18110);
xor U18755 (N_18755,N_17142,N_17918);
xor U18756 (N_18756,N_15647,N_17790);
or U18757 (N_18757,N_15762,N_18303);
nand U18758 (N_18758,N_17499,N_15975);
nand U18759 (N_18759,N_16268,N_18468);
and U18760 (N_18760,N_16372,N_18215);
xor U18761 (N_18761,N_18599,N_16438);
and U18762 (N_18762,N_17247,N_16304);
and U18763 (N_18763,N_17006,N_17822);
nand U18764 (N_18764,N_18305,N_16704);
xor U18765 (N_18765,N_16148,N_16053);
and U18766 (N_18766,N_15731,N_16516);
or U18767 (N_18767,N_16139,N_16935);
nor U18768 (N_18768,N_17675,N_16557);
and U18769 (N_18769,N_18180,N_18315);
nand U18770 (N_18770,N_17877,N_17814);
xnor U18771 (N_18771,N_18157,N_17632);
and U18772 (N_18772,N_16582,N_18564);
nand U18773 (N_18773,N_17562,N_16506);
and U18774 (N_18774,N_16157,N_16484);
nor U18775 (N_18775,N_15856,N_18246);
xor U18776 (N_18776,N_17543,N_18448);
nor U18777 (N_18777,N_16262,N_16041);
and U18778 (N_18778,N_18071,N_16292);
nand U18779 (N_18779,N_17697,N_16101);
nand U18780 (N_18780,N_18511,N_15643);
and U18781 (N_18781,N_16260,N_18690);
xnor U18782 (N_18782,N_16699,N_18452);
xor U18783 (N_18783,N_17252,N_17497);
or U18784 (N_18784,N_17883,N_18548);
and U18785 (N_18785,N_18674,N_17507);
nand U18786 (N_18786,N_17825,N_17719);
nor U18787 (N_18787,N_17279,N_17625);
xnor U18788 (N_18788,N_16963,N_17937);
nand U18789 (N_18789,N_16684,N_17585);
or U18790 (N_18790,N_17452,N_17687);
and U18791 (N_18791,N_16369,N_16532);
and U18792 (N_18792,N_17523,N_15864);
nand U18793 (N_18793,N_17828,N_15688);
nor U18794 (N_18794,N_17531,N_18447);
or U18795 (N_18795,N_16601,N_16514);
nand U18796 (N_18796,N_15741,N_16063);
nor U18797 (N_18797,N_16667,N_18334);
nor U18798 (N_18798,N_18076,N_16643);
nand U18799 (N_18799,N_17626,N_17462);
nand U18800 (N_18800,N_16005,N_16952);
or U18801 (N_18801,N_15928,N_16927);
and U18802 (N_18802,N_17301,N_16217);
xor U18803 (N_18803,N_16492,N_17821);
xor U18804 (N_18804,N_16705,N_15716);
nand U18805 (N_18805,N_18039,N_17286);
xnor U18806 (N_18806,N_17668,N_15759);
nor U18807 (N_18807,N_18089,N_17480);
nand U18808 (N_18808,N_16026,N_16814);
or U18809 (N_18809,N_17624,N_18026);
nor U18810 (N_18810,N_16614,N_17358);
nor U18811 (N_18811,N_17032,N_18285);
nand U18812 (N_18812,N_17979,N_18450);
nor U18813 (N_18813,N_17983,N_18366);
xnor U18814 (N_18814,N_18086,N_16512);
xnor U18815 (N_18815,N_18224,N_18238);
and U18816 (N_18816,N_15721,N_17193);
nand U18817 (N_18817,N_15627,N_18604);
nand U18818 (N_18818,N_18239,N_16067);
nor U18819 (N_18819,N_17038,N_17800);
xnor U18820 (N_18820,N_18014,N_16622);
nor U18821 (N_18821,N_16336,N_18547);
nor U18822 (N_18822,N_17617,N_18236);
and U18823 (N_18823,N_18104,N_17492);
and U18824 (N_18824,N_16723,N_17303);
xor U18825 (N_18825,N_17984,N_16736);
or U18826 (N_18826,N_16273,N_15652);
and U18827 (N_18827,N_18118,N_17349);
xnor U18828 (N_18828,N_17691,N_16447);
or U18829 (N_18829,N_17775,N_18418);
nor U18830 (N_18830,N_17879,N_18323);
nor U18831 (N_18831,N_16591,N_16066);
or U18832 (N_18832,N_16778,N_15964);
and U18833 (N_18833,N_15654,N_18029);
and U18834 (N_18834,N_18376,N_18154);
nor U18835 (N_18835,N_18423,N_18383);
nor U18836 (N_18836,N_18333,N_15971);
nand U18837 (N_18837,N_16445,N_15668);
nand U18838 (N_18838,N_15789,N_16465);
xor U18839 (N_18839,N_17659,N_18731);
nor U18840 (N_18840,N_18730,N_18225);
and U18841 (N_18841,N_18216,N_16930);
nand U18842 (N_18842,N_17986,N_17282);
or U18843 (N_18843,N_15715,N_17759);
nor U18844 (N_18844,N_16297,N_16692);
nand U18845 (N_18845,N_18654,N_17402);
xnor U18846 (N_18846,N_16224,N_16872);
and U18847 (N_18847,N_16923,N_17258);
nand U18848 (N_18848,N_18403,N_18072);
nor U18849 (N_18849,N_15909,N_17850);
or U18850 (N_18850,N_17200,N_17586);
or U18851 (N_18851,N_17926,N_16842);
or U18852 (N_18852,N_16290,N_16884);
nor U18853 (N_18853,N_17036,N_17249);
nand U18854 (N_18854,N_16785,N_16362);
or U18855 (N_18855,N_18529,N_18313);
and U18856 (N_18856,N_18196,N_16654);
nand U18857 (N_18857,N_16974,N_17673);
and U18858 (N_18858,N_18397,N_18142);
and U18859 (N_18859,N_17166,N_15807);
and U18860 (N_18860,N_18633,N_17327);
and U18861 (N_18861,N_17149,N_16034);
or U18862 (N_18862,N_17220,N_16385);
xor U18863 (N_18863,N_16665,N_17265);
nand U18864 (N_18864,N_17540,N_18257);
and U18865 (N_18865,N_16620,N_16382);
nand U18866 (N_18866,N_16676,N_16401);
or U18867 (N_18867,N_15932,N_17328);
or U18868 (N_18868,N_16395,N_18724);
nor U18869 (N_18869,N_15933,N_16464);
and U18870 (N_18870,N_17155,N_17250);
nand U18871 (N_18871,N_16964,N_18369);
or U18872 (N_18872,N_18412,N_16856);
xnor U18873 (N_18873,N_16386,N_15782);
or U18874 (N_18874,N_17664,N_18056);
or U18875 (N_18875,N_17027,N_17544);
xnor U18876 (N_18876,N_17805,N_16639);
nor U18877 (N_18877,N_18617,N_17439);
nand U18878 (N_18878,N_18600,N_17855);
xnor U18879 (N_18879,N_17113,N_17550);
nand U18880 (N_18880,N_16973,N_16587);
nor U18881 (N_18881,N_18302,N_18358);
xnor U18882 (N_18882,N_17779,N_18677);
and U18883 (N_18883,N_18706,N_16957);
and U18884 (N_18884,N_18141,N_17799);
and U18885 (N_18885,N_18166,N_18590);
xnor U18886 (N_18886,N_15858,N_17718);
and U18887 (N_18887,N_16370,N_16602);
or U18888 (N_18888,N_17931,N_17630);
and U18889 (N_18889,N_16649,N_16215);
nor U18890 (N_18890,N_17844,N_16777);
and U18891 (N_18891,N_16206,N_18531);
xnor U18892 (N_18892,N_16106,N_16278);
xnor U18893 (N_18893,N_16827,N_17558);
xor U18894 (N_18894,N_18497,N_18569);
or U18895 (N_18895,N_18459,N_17880);
or U18896 (N_18896,N_17486,N_18640);
xnor U18897 (N_18897,N_16311,N_16112);
and U18898 (N_18898,N_16211,N_17614);
or U18899 (N_18899,N_17138,N_16795);
xnor U18900 (N_18900,N_16521,N_16167);
nor U18901 (N_18901,N_18061,N_17817);
and U18902 (N_18902,N_18133,N_16460);
xor U18903 (N_18903,N_16284,N_17432);
and U18904 (N_18904,N_15816,N_15703);
xnor U18905 (N_18905,N_17660,N_17577);
nand U18906 (N_18906,N_16763,N_17270);
or U18907 (N_18907,N_18126,N_18115);
nor U18908 (N_18908,N_17627,N_18117);
nand U18909 (N_18909,N_16774,N_16909);
and U18910 (N_18910,N_15693,N_18454);
nand U18911 (N_18911,N_17517,N_17228);
nor U18912 (N_18912,N_18184,N_17902);
and U18913 (N_18913,N_17703,N_18370);
nand U18914 (N_18914,N_18003,N_17663);
nor U18915 (N_18915,N_18554,N_16715);
and U18916 (N_18916,N_16307,N_16073);
nor U18917 (N_18917,N_18637,N_17953);
nor U18918 (N_18918,N_18553,N_18000);
or U18919 (N_18919,N_16749,N_16926);
nand U18920 (N_18920,N_18693,N_15787);
and U18921 (N_18921,N_16531,N_15718);
or U18922 (N_18922,N_16046,N_17650);
or U18923 (N_18923,N_17119,N_17067);
or U18924 (N_18924,N_17016,N_16200);
xnor U18925 (N_18925,N_17580,N_17542);
or U18926 (N_18926,N_17564,N_16503);
nand U18927 (N_18927,N_17310,N_18328);
xor U18928 (N_18928,N_17620,N_16976);
or U18929 (N_18929,N_17893,N_15879);
nor U18930 (N_18930,N_16631,N_16078);
nor U18931 (N_18931,N_16708,N_17251);
nand U18932 (N_18932,N_16186,N_16308);
and U18933 (N_18933,N_16703,N_17741);
nand U18934 (N_18934,N_17406,N_16394);
and U18935 (N_18935,N_15779,N_17366);
nand U18936 (N_18936,N_17904,N_16943);
xor U18937 (N_18937,N_18145,N_18433);
and U18938 (N_18938,N_16127,N_16992);
or U18939 (N_18939,N_18623,N_16012);
or U18940 (N_18940,N_16373,N_17864);
nand U18941 (N_18941,N_17901,N_17921);
nor U18942 (N_18942,N_15870,N_16613);
or U18943 (N_18943,N_15685,N_16580);
and U18944 (N_18944,N_17304,N_16184);
nand U18945 (N_18945,N_18012,N_18296);
nand U18946 (N_18946,N_18507,N_15899);
or U18947 (N_18947,N_16068,N_18259);
xor U18948 (N_18948,N_16096,N_18669);
and U18949 (N_18949,N_17876,N_16743);
and U18950 (N_18950,N_18463,N_18361);
nand U18951 (N_18951,N_17407,N_17804);
nor U18952 (N_18952,N_18137,N_16932);
nor U18953 (N_18953,N_16192,N_16389);
nand U18954 (N_18954,N_15637,N_17377);
xnor U18955 (N_18955,N_16657,N_17306);
nor U18956 (N_18956,N_16618,N_17831);
and U18957 (N_18957,N_17040,N_16809);
xor U18958 (N_18958,N_16753,N_16775);
nor U18959 (N_18959,N_18228,N_17281);
xor U18960 (N_18960,N_16874,N_18001);
and U18961 (N_18961,N_18703,N_17399);
or U18962 (N_18962,N_18588,N_17750);
or U18963 (N_18963,N_17778,N_15752);
nor U18964 (N_18964,N_18011,N_16728);
or U18965 (N_18965,N_18127,N_17280);
nand U18966 (N_18966,N_15941,N_17992);
or U18967 (N_18967,N_18040,N_16534);
and U18968 (N_18968,N_15904,N_17842);
xnor U18969 (N_18969,N_18211,N_17557);
and U18970 (N_18970,N_17830,N_17030);
nand U18971 (N_18971,N_17218,N_17034);
xor U18972 (N_18972,N_16845,N_16549);
xnor U18973 (N_18973,N_18414,N_17299);
xor U18974 (N_18974,N_16493,N_17444);
nor U18975 (N_18975,N_17742,N_16494);
xnor U18976 (N_18976,N_18518,N_16018);
xnor U18977 (N_18977,N_17665,N_16244);
and U18978 (N_18978,N_17049,N_17256);
xor U18979 (N_18979,N_18720,N_18645);
nor U18980 (N_18980,N_17043,N_17930);
or U18981 (N_18981,N_16746,N_17647);
nor U18982 (N_18982,N_17035,N_16387);
and U18983 (N_18983,N_16410,N_17309);
nand U18984 (N_18984,N_16031,N_17803);
nor U18985 (N_18985,N_16553,N_16942);
and U18986 (N_18986,N_17686,N_17246);
nand U18987 (N_18987,N_18292,N_16677);
xnor U18988 (N_18988,N_16419,N_16655);
nand U18989 (N_18989,N_16700,N_17526);
and U18990 (N_18990,N_18605,N_17928);
and U18991 (N_18991,N_18657,N_17257);
and U18992 (N_18992,N_17160,N_17423);
or U18993 (N_18993,N_15963,N_18695);
or U18994 (N_18994,N_18424,N_18644);
xor U18995 (N_18995,N_17722,N_17774);
xnor U18996 (N_18996,N_16301,N_16662);
or U18997 (N_18997,N_18140,N_17989);
or U18998 (N_18998,N_17757,N_18055);
or U18999 (N_18999,N_16427,N_16265);
or U19000 (N_19000,N_16478,N_16044);
and U19001 (N_19001,N_17987,N_17797);
xor U19002 (N_19002,N_18460,N_17955);
or U19003 (N_19003,N_15672,N_18359);
and U19004 (N_19004,N_17766,N_16183);
nand U19005 (N_19005,N_18010,N_15838);
and U19006 (N_19006,N_17416,N_16858);
and U19007 (N_19007,N_18129,N_18562);
nand U19008 (N_19008,N_16489,N_18063);
nand U19009 (N_19009,N_16145,N_18200);
nor U19010 (N_19010,N_16533,N_15810);
or U19011 (N_19011,N_15737,N_16016);
and U19012 (N_19012,N_17115,N_16697);
nor U19013 (N_19013,N_17853,N_16783);
and U19014 (N_19014,N_18636,N_16691);
nand U19015 (N_19015,N_16014,N_16366);
nand U19016 (N_19016,N_18610,N_18496);
nor U19017 (N_19017,N_17430,N_17938);
xor U19018 (N_19018,N_18429,N_16568);
and U19019 (N_19019,N_17044,N_17175);
nor U19020 (N_19020,N_18603,N_16756);
nand U19021 (N_19021,N_15937,N_16844);
nand U19022 (N_19022,N_17451,N_15891);
nand U19023 (N_19023,N_18567,N_16017);
nand U19024 (N_19024,N_15645,N_15842);
nor U19025 (N_19025,N_16983,N_18593);
and U19026 (N_19026,N_16590,N_17765);
nor U19027 (N_19027,N_17272,N_17939);
nor U19028 (N_19028,N_16737,N_18156);
and U19029 (N_19029,N_17317,N_17212);
nor U19030 (N_19030,N_17888,N_16539);
nor U19031 (N_19031,N_16421,N_16230);
xor U19032 (N_19032,N_16559,N_17436);
nand U19033 (N_19033,N_15832,N_17022);
or U19034 (N_19034,N_15653,N_15991);
nor U19035 (N_19035,N_18167,N_17581);
and U19036 (N_19036,N_17005,N_17404);
nand U19037 (N_19037,N_18365,N_17391);
and U19038 (N_19038,N_18719,N_16889);
nor U19039 (N_19039,N_16837,N_17133);
or U19040 (N_19040,N_17078,N_18467);
and U19041 (N_19041,N_17141,N_15750);
xnor U19042 (N_19042,N_17111,N_17368);
and U19043 (N_19043,N_17371,N_17125);
nor U19044 (N_19044,N_18676,N_16047);
nand U19045 (N_19045,N_15689,N_18023);
nor U19046 (N_19046,N_15747,N_17187);
and U19047 (N_19047,N_15720,N_18632);
xnor U19048 (N_19048,N_18464,N_18143);
and U19049 (N_19049,N_18155,N_18389);
and U19050 (N_19050,N_18715,N_17999);
and U19051 (N_19051,N_16325,N_15809);
xnor U19052 (N_19052,N_17575,N_17372);
xor U19053 (N_19053,N_15986,N_16270);
xnor U19054 (N_19054,N_17375,N_17001);
or U19055 (N_19055,N_17426,N_18712);
or U19056 (N_19056,N_17000,N_16042);
or U19057 (N_19057,N_18421,N_16686);
or U19058 (N_19058,N_16589,N_17041);
and U19059 (N_19059,N_16538,N_17355);
or U19060 (N_19060,N_17527,N_17116);
nand U19061 (N_19061,N_16470,N_16334);
nor U19062 (N_19062,N_16713,N_16733);
and U19063 (N_19063,N_17730,N_15895);
nor U19064 (N_19064,N_16712,N_18324);
and U19065 (N_19065,N_17818,N_16725);
nor U19066 (N_19066,N_17165,N_17677);
nand U19067 (N_19067,N_18408,N_16196);
xor U19068 (N_19068,N_16288,N_17071);
nand U19069 (N_19069,N_17300,N_18121);
and U19070 (N_19070,N_15996,N_17923);
nand U19071 (N_19071,N_17052,N_16058);
or U19072 (N_19072,N_16501,N_15918);
xor U19073 (N_19073,N_16579,N_16679);
nor U19074 (N_19074,N_18349,N_17737);
xnor U19075 (N_19075,N_16852,N_16787);
nor U19076 (N_19076,N_15764,N_16586);
xor U19077 (N_19077,N_15755,N_16352);
and U19078 (N_19078,N_17701,N_18019);
xnor U19079 (N_19079,N_17960,N_16111);
or U19080 (N_19080,N_15985,N_16381);
or U19081 (N_19081,N_18209,N_17454);
or U19082 (N_19082,N_17743,N_16804);
or U19083 (N_19083,N_17520,N_16955);
or U19084 (N_19084,N_16571,N_17393);
and U19085 (N_19085,N_15657,N_18540);
nand U19086 (N_19086,N_17106,N_16626);
and U19087 (N_19087,N_18269,N_16335);
nor U19088 (N_19088,N_17360,N_16767);
nand U19089 (N_19089,N_18387,N_18456);
nand U19090 (N_19090,N_17117,N_18083);
nor U19091 (N_19091,N_17661,N_17491);
nand U19092 (N_19092,N_16818,N_18405);
or U19093 (N_19093,N_15894,N_17356);
nand U19094 (N_19094,N_17796,N_16082);
xor U19095 (N_19095,N_17636,N_16898);
xor U19096 (N_19096,N_17079,N_16209);
nor U19097 (N_19097,N_18013,N_16102);
and U19098 (N_19098,N_16529,N_16981);
and U19099 (N_19099,N_17498,N_17561);
or U19100 (N_19100,N_18021,N_17178);
nor U19101 (N_19101,N_18560,N_18346);
nand U19102 (N_19102,N_18700,N_18252);
or U19103 (N_19103,N_17185,N_18686);
and U19104 (N_19104,N_18671,N_17235);
nor U19105 (N_19105,N_15871,N_17466);
xnor U19106 (N_19106,N_16754,N_18608);
nand U19107 (N_19107,N_18481,N_15679);
nor U19108 (N_19108,N_15992,N_16772);
or U19109 (N_19109,N_18404,N_17209);
and U19110 (N_19110,N_15698,N_17020);
nand U19111 (N_19111,N_17188,N_16323);
xnor U19112 (N_19112,N_18661,N_16103);
or U19113 (N_19113,N_16758,N_16543);
or U19114 (N_19114,N_16796,N_16770);
and U19115 (N_19115,N_18530,N_17483);
nand U19116 (N_19116,N_16822,N_16393);
nand U19117 (N_19117,N_16136,N_15994);
or U19118 (N_19118,N_16537,N_17887);
or U19119 (N_19119,N_15709,N_16024);
nand U19120 (N_19120,N_18559,N_17489);
nand U19121 (N_19121,N_16418,N_18298);
or U19122 (N_19122,N_18667,N_17101);
nor U19123 (N_19123,N_16940,N_18173);
nand U19124 (N_19124,N_17764,N_16583);
nand U19125 (N_19125,N_18572,N_16566);
xnor U19126 (N_19126,N_16698,N_18525);
and U19127 (N_19127,N_16322,N_18628);
nand U19128 (N_19128,N_18697,N_16162);
nor U19129 (N_19129,N_18339,N_15893);
or U19130 (N_19130,N_17823,N_16810);
or U19131 (N_19131,N_16987,N_16309);
xor U19132 (N_19132,N_16247,N_18622);
nand U19133 (N_19133,N_16187,N_18325);
or U19134 (N_19134,N_17386,N_16956);
or U19135 (N_19135,N_16371,N_17934);
nand U19136 (N_19136,N_16864,N_16415);
nor U19137 (N_19137,N_16263,N_17680);
nor U19138 (N_19138,N_17087,N_18015);
xor U19139 (N_19139,N_18374,N_17996);
xor U19140 (N_19140,N_18379,N_16638);
nand U19141 (N_19141,N_16922,N_18054);
nor U19142 (N_19142,N_15770,N_17551);
xnor U19143 (N_19143,N_17990,N_17223);
and U19144 (N_19144,N_17157,N_16104);
nand U19145 (N_19145,N_18746,N_18392);
nor U19146 (N_19146,N_15837,N_16132);
nor U19147 (N_19147,N_18192,N_15930);
or U19148 (N_19148,N_15820,N_16074);
xor U19149 (N_19149,N_15812,N_18396);
or U19150 (N_19150,N_17214,N_16199);
and U19151 (N_19151,N_18718,N_16599);
nor U19152 (N_19152,N_18487,N_18739);
xor U19153 (N_19153,N_18186,N_16218);
nor U19154 (N_19154,N_16165,N_18563);
xnor U19155 (N_19155,N_17758,N_17882);
nand U19156 (N_19156,N_17894,N_18742);
nand U19157 (N_19157,N_18197,N_16632);
nand U19158 (N_19158,N_17461,N_16857);
and U19159 (N_19159,N_16422,N_18651);
xnor U19160 (N_19160,N_18291,N_17457);
or U19161 (N_19161,N_17903,N_16895);
xor U19162 (N_19162,N_15890,N_18509);
xnor U19163 (N_19163,N_17954,N_18624);
and U19164 (N_19164,N_16870,N_17198);
or U19165 (N_19165,N_17819,N_16281);
or U19166 (N_19166,N_18230,N_15630);
and U19167 (N_19167,N_17453,N_18362);
or U19168 (N_19168,N_17177,N_17392);
nor U19169 (N_19169,N_17786,N_18635);
nor U19170 (N_19170,N_16469,N_16236);
xor U19171 (N_19171,N_18357,N_18368);
xnor U19172 (N_19172,N_18103,N_16688);
xnor U19173 (N_19173,N_17860,N_18229);
nor U19174 (N_19174,N_17050,N_17202);
xnor U19175 (N_19175,N_16285,N_17136);
or U19176 (N_19176,N_16741,N_18082);
or U19177 (N_19177,N_16023,N_17023);
or U19178 (N_19178,N_16189,N_17025);
xor U19179 (N_19179,N_15961,N_16330);
nor U19180 (N_19180,N_16908,N_15699);
nand U19181 (N_19181,N_17288,N_17770);
and U19182 (N_19182,N_18130,N_17781);
xor U19183 (N_19183,N_17835,N_18288);
or U19184 (N_19184,N_17290,N_17857);
nand U19185 (N_19185,N_17717,N_18504);
nand U19186 (N_19186,N_17287,N_18411);
nor U19187 (N_19187,N_17525,N_17126);
xnor U19188 (N_19188,N_18297,N_15924);
nand U19189 (N_19189,N_17827,N_17653);
xnor U19190 (N_19190,N_16841,N_16672);
and U19191 (N_19191,N_17144,N_17112);
or U19192 (N_19192,N_16780,N_16666);
or U19193 (N_19193,N_18726,N_15999);
and U19194 (N_19194,N_17007,N_17973);
nor U19195 (N_19195,N_16015,N_18025);
nand U19196 (N_19196,N_15970,N_15775);
nand U19197 (N_19197,N_16091,N_16541);
nand U19198 (N_19198,N_15665,N_18522);
nand U19199 (N_19199,N_17982,N_18377);
nor U19200 (N_19200,N_16246,N_17514);
and U19201 (N_19201,N_15944,N_16072);
or U19202 (N_19202,N_17225,N_15841);
xnor U19203 (N_19203,N_16762,N_18213);
xor U19204 (N_19204,N_16659,N_16353);
nor U19205 (N_19205,N_16994,N_17843);
nor U19206 (N_19206,N_16122,N_16037);
or U19207 (N_19207,N_17980,N_18568);
nor U19208 (N_19208,N_17807,N_16630);
nor U19209 (N_19209,N_16612,N_16750);
xnor U19210 (N_19210,N_17897,N_17541);
or U19211 (N_19211,N_16181,N_16197);
or U19212 (N_19212,N_18735,N_17216);
nor U19213 (N_19213,N_16522,N_15885);
nor U19214 (N_19214,N_18242,N_16714);
nor U19215 (N_19215,N_18049,N_15777);
nand U19216 (N_19216,N_17529,N_17608);
or U19217 (N_19217,N_16569,N_16163);
nor U19218 (N_19218,N_17376,N_18652);
nand U19219 (N_19219,N_18432,N_15868);
xnor U19220 (N_19220,N_18535,N_17201);
and U19221 (N_19221,N_18091,N_15998);
nand U19222 (N_19222,N_18098,N_15936);
nor U19223 (N_19223,N_15650,N_17648);
nand U19224 (N_19224,N_16635,N_18364);
and U19225 (N_19225,N_17508,N_17456);
or U19226 (N_19226,N_17325,N_17048);
or U19227 (N_19227,N_16359,N_17271);
xnor U19228 (N_19228,N_18314,N_16761);
nand U19229 (N_19229,N_16257,N_18048);
nand U19230 (N_19230,N_18017,N_16020);
nor U19231 (N_19231,N_17278,N_16830);
nand U19232 (N_19232,N_17276,N_17365);
nor U19233 (N_19233,N_16114,N_16039);
and U19234 (N_19234,N_16921,N_16116);
nor U19235 (N_19235,N_15923,N_16242);
or U19236 (N_19236,N_16479,N_15704);
and U19237 (N_19237,N_15902,N_17840);
nand U19238 (N_19238,N_17726,N_15960);
and U19239 (N_19239,N_15995,N_16152);
nand U19240 (N_19240,N_15788,N_16097);
nand U19241 (N_19241,N_18596,N_16071);
and U19242 (N_19242,N_18282,N_17801);
xnor U19243 (N_19243,N_18308,N_17751);
or U19244 (N_19244,N_17236,N_17080);
nand U19245 (N_19245,N_16887,N_16156);
xnor U19246 (N_19246,N_18451,N_17054);
nor U19247 (N_19247,N_16982,N_17802);
nand U19248 (N_19248,N_18702,N_16180);
xnor U19249 (N_19249,N_16918,N_15743);
nand U19250 (N_19250,N_18526,N_17316);
xnor U19251 (N_19251,N_17073,N_18638);
xnor U19252 (N_19252,N_18233,N_16911);
nor U19253 (N_19253,N_18639,N_18193);
xnor U19254 (N_19254,N_17846,N_16355);
xnor U19255 (N_19255,N_17100,N_16882);
xnor U19256 (N_19256,N_15676,N_17951);
nand U19257 (N_19257,N_18337,N_17875);
nor U19258 (N_19258,N_17587,N_16271);
or U19259 (N_19259,N_17074,N_18018);
xor U19260 (N_19260,N_17560,N_16941);
or U19261 (N_19261,N_18330,N_17907);
nand U19262 (N_19262,N_17832,N_17629);
or U19263 (N_19263,N_16511,N_15742);
nand U19264 (N_19264,N_16624,N_15667);
nor U19265 (N_19265,N_16815,N_17611);
nor U19266 (N_19266,N_15953,N_18745);
nor U19267 (N_19267,N_16576,N_17192);
and U19268 (N_19268,N_16191,N_18457);
or U19269 (N_19269,N_15833,N_18744);
nand U19270 (N_19270,N_16129,N_18177);
nor U19271 (N_19271,N_17072,N_16623);
nor U19272 (N_19272,N_18717,N_17064);
xor U19273 (N_19273,N_17705,N_16350);
nor U19274 (N_19274,N_17771,N_17578);
or U19275 (N_19275,N_17215,N_17602);
or U19276 (N_19276,N_17333,N_15910);
or U19277 (N_19277,N_17095,N_18251);
nor U19278 (N_19278,N_16435,N_16821);
nor U19279 (N_19279,N_15734,N_16695);
or U19280 (N_19280,N_15951,N_16825);
nand U19281 (N_19281,N_16650,N_18538);
nand U19282 (N_19282,N_17400,N_17754);
nor U19283 (N_19283,N_16651,N_16969);
xor U19284 (N_19284,N_15857,N_15927);
nor U19285 (N_19285,N_16258,N_17021);
nor U19286 (N_19286,N_16899,N_17045);
nand U19287 (N_19287,N_18256,N_16076);
and U19288 (N_19288,N_18629,N_17961);
or U19289 (N_19289,N_16117,N_16070);
nor U19290 (N_19290,N_15666,N_18470);
and U19291 (N_19291,N_18271,N_15957);
nand U19292 (N_19292,N_17345,N_18147);
xnor U19293 (N_19293,N_17570,N_17572);
and U19294 (N_19294,N_16443,N_18514);
nor U19295 (N_19295,N_16253,N_17692);
and U19296 (N_19296,N_17566,N_18112);
or U19297 (N_19297,N_18664,N_16064);
xor U19298 (N_19298,N_16995,N_16879);
nor U19299 (N_19299,N_18503,N_18248);
nand U19300 (N_19300,N_17576,N_16838);
xnor U19301 (N_19301,N_16680,N_18268);
nor U19302 (N_19302,N_18144,N_18434);
nor U19303 (N_19303,N_16061,N_17735);
nor U19304 (N_19304,N_18153,N_17003);
nor U19305 (N_19305,N_16604,N_18449);
xor U19306 (N_19306,N_17197,N_17469);
xor U19307 (N_19307,N_15738,N_18453);
nand U19308 (N_19308,N_18249,N_17128);
and U19309 (N_19309,N_17084,N_16384);
or U19310 (N_19310,N_16719,N_18428);
or U19311 (N_19311,N_17976,N_18609);
nand U19312 (N_19312,N_17046,N_16458);
or U19313 (N_19313,N_18595,N_17884);
and U19314 (N_19314,N_16890,N_17411);
nand U19315 (N_19315,N_17676,N_17331);
nor U19316 (N_19316,N_17208,N_17862);
xor U19317 (N_19317,N_18692,N_17662);
nand U19318 (N_19318,N_16151,N_18301);
nor U19319 (N_19319,N_16043,N_17847);
xnor U19320 (N_19320,N_16220,N_15943);
or U19321 (N_19321,N_18465,N_16900);
and U19322 (N_19322,N_16453,N_15935);
xnor U19323 (N_19323,N_16634,N_16933);
nor U19324 (N_19324,N_17156,N_17460);
nand U19325 (N_19325,N_17622,N_16967);
and U19326 (N_19326,N_16439,N_16222);
and U19327 (N_19327,N_17307,N_16945);
nor U19328 (N_19328,N_16998,N_17417);
xor U19329 (N_19329,N_16993,N_16077);
and U19330 (N_19330,N_16906,N_17645);
and U19331 (N_19331,N_17104,N_18489);
or U19332 (N_19332,N_16836,N_18024);
xor U19333 (N_19333,N_16305,N_18343);
and U19334 (N_19334,N_17793,N_16588);
nor U19335 (N_19335,N_16153,N_17174);
or U19336 (N_19336,N_17545,N_17350);
xor U19337 (N_19337,N_18169,N_16938);
nor U19338 (N_19338,N_16594,N_18163);
or U19339 (N_19339,N_16975,N_17274);
and U19340 (N_19340,N_17899,N_15922);
nand U19341 (N_19341,N_16351,N_17302);
nand U19342 (N_19342,N_18698,N_16931);
nand U19343 (N_19343,N_17769,N_16146);
nor U19344 (N_19344,N_17806,N_17912);
nor U19345 (N_19345,N_17914,N_16644);
nor U19346 (N_19346,N_17579,N_16202);
and U19347 (N_19347,N_16223,N_16851);
or U19348 (N_19348,N_15724,N_16764);
nand U19349 (N_19349,N_17180,N_18232);
nor U19350 (N_19350,N_17619,N_18747);
or U19351 (N_19351,N_17612,N_18131);
and U19352 (N_19352,N_16021,N_16515);
xnor U19353 (N_19353,N_16429,N_16978);
and U19354 (N_19354,N_16251,N_17448);
nor U19355 (N_19355,N_18513,N_18655);
nand U19356 (N_19356,N_18394,N_16452);
and U19357 (N_19357,N_16170,N_17684);
or U19358 (N_19358,N_18139,N_18185);
nand U19359 (N_19359,N_16628,N_18534);
nor U19360 (N_19360,N_17556,N_17656);
and U19361 (N_19361,N_17695,N_15980);
xnor U19362 (N_19362,N_16524,N_17727);
and U19363 (N_19363,N_16954,N_16883);
xnor U19364 (N_19364,N_17908,N_15695);
xnor U19365 (N_19365,N_16451,N_17829);
nand U19366 (N_19366,N_18659,N_16147);
nand U19367 (N_19367,N_15914,N_17638);
and U19368 (N_19368,N_17413,N_17204);
nand U19369 (N_19369,N_17988,N_18352);
nor U19370 (N_19370,N_15648,N_17496);
or U19371 (N_19371,N_17711,N_16653);
nor U19372 (N_19372,N_15908,N_18069);
nand U19373 (N_19373,N_18512,N_18202);
nor U19374 (N_19374,N_18729,N_15877);
or U19375 (N_19375,N_17870,N_18340);
and U19376 (N_19376,N_17978,N_16341);
or U19377 (N_19377,N_17037,N_18594);
nand U19378 (N_19378,N_16233,N_18519);
nor U19379 (N_19379,N_18311,N_18276);
and U19380 (N_19380,N_17515,N_17925);
and U19381 (N_19381,N_17026,N_17420);
or U19382 (N_19382,N_17553,N_15800);
nand U19383 (N_19383,N_15897,N_17061);
nand U19384 (N_19384,N_15780,N_17582);
or U19385 (N_19385,N_18626,N_16939);
and U19386 (N_19386,N_17213,N_18066);
xor U19387 (N_19387,N_16806,N_15797);
or U19388 (N_19388,N_17528,N_16637);
nand U19389 (N_19389,N_15806,N_16925);
and U19390 (N_19390,N_18164,N_15956);
xor U19391 (N_19391,N_16446,N_16660);
xnor U19392 (N_19392,N_17445,N_18508);
nor U19393 (N_19393,N_16221,N_17651);
xnor U19394 (N_19394,N_17364,N_16648);
nor U19395 (N_19395,N_18727,N_16913);
or U19396 (N_19396,N_16302,N_17667);
nor U19397 (N_19397,N_17519,N_16585);
or U19398 (N_19398,N_17066,N_17158);
xor U19399 (N_19399,N_18279,N_18101);
nand U19400 (N_19400,N_16876,N_17296);
nor U19401 (N_19401,N_18042,N_17964);
xnor U19402 (N_19402,N_18036,N_17872);
nand U19403 (N_19403,N_15678,N_17941);
nand U19404 (N_19404,N_16138,N_16702);
nand U19405 (N_19405,N_15646,N_17164);
nor U19406 (N_19406,N_16166,N_17412);
or U19407 (N_19407,N_16597,N_16463);
and U19408 (N_19408,N_18341,N_16142);
nand U19409 (N_19409,N_17443,N_18065);
nor U19410 (N_19410,N_17091,N_18310);
nor U19411 (N_19411,N_17267,N_16792);
nor U19412 (N_19412,N_16252,N_18583);
nand U19413 (N_19413,N_16573,N_17315);
nor U19414 (N_19414,N_18107,N_17977);
nand U19415 (N_19415,N_17163,N_16853);
and U19416 (N_19416,N_17446,N_15733);
and U19417 (N_19417,N_17172,N_17378);
or U19418 (N_19418,N_18443,N_16903);
nand U19419 (N_19419,N_15796,N_18435);
nand U19420 (N_19420,N_17985,N_17082);
xor U19421 (N_19421,N_16732,N_17707);
xor U19422 (N_19422,N_17284,N_16765);
or U19423 (N_19423,N_18516,N_18125);
and U19424 (N_19424,N_16875,N_17437);
xor U19425 (N_19425,N_17255,N_18052);
nor U19426 (N_19426,N_16361,N_18650);
and U19427 (N_19427,N_16317,N_17487);
or U19428 (N_19428,N_17184,N_16488);
nand U19429 (N_19429,N_15711,N_17194);
and U19430 (N_19430,N_15834,N_16124);
nor U19431 (N_19431,N_18060,N_17203);
xnor U19432 (N_19432,N_17183,N_17425);
and U19433 (N_19433,N_17681,N_17485);
nor U19434 (N_19434,N_17024,N_15847);
xnor U19435 (N_19435,N_18390,N_17539);
nand U19436 (N_19436,N_18565,N_16798);
nor U19437 (N_19437,N_18338,N_16348);
xnor U19438 (N_19438,N_18344,N_17513);
and U19439 (N_19439,N_18354,N_18031);
or U19440 (N_19440,N_18461,N_17308);
nor U19441 (N_19441,N_16605,N_17981);
nand U19442 (N_19442,N_18416,N_16726);
nor U19443 (N_19443,N_16950,N_17671);
or U19444 (N_19444,N_16542,N_16050);
nor U19445 (N_19445,N_15825,N_16407);
xnor U19446 (N_19446,N_16340,N_17971);
nor U19447 (N_19447,N_16990,N_16420);
and U19448 (N_19448,N_16669,N_18493);
nand U19449 (N_19449,N_17099,N_18351);
or U19450 (N_19450,N_15748,N_16840);
nand U19451 (N_19451,N_18375,N_17736);
xor U19452 (N_19452,N_16079,N_18350);
and U19453 (N_19453,N_18046,N_16641);
xnor U19454 (N_19454,N_15694,N_17913);
or U19455 (N_19455,N_15968,N_18273);
nor U19456 (N_19456,N_18492,N_16345);
nor U19457 (N_19457,N_17708,N_16300);
or U19458 (N_19458,N_18067,N_18087);
nand U19459 (N_19459,N_18290,N_15817);
nand U19460 (N_19460,N_15954,N_16368);
or U19461 (N_19461,N_17081,N_17217);
and U19462 (N_19462,N_18217,N_17114);
xnor U19463 (N_19463,N_16828,N_17810);
or U19464 (N_19464,N_16929,N_16490);
xnor U19465 (N_19465,N_18475,N_18212);
nand U19466 (N_19466,N_16962,N_17776);
nor U19467 (N_19467,N_17699,N_17051);
nor U19468 (N_19468,N_16045,N_17505);
nor U19469 (N_19469,N_16204,N_15815);
xor U19470 (N_19470,N_17493,N_16897);
nand U19471 (N_19471,N_17920,N_18662);
nand U19472 (N_19472,N_16476,N_17297);
nor U19473 (N_19473,N_16551,N_18485);
nor U19474 (N_19474,N_17326,N_18445);
or U19475 (N_19475,N_15859,N_16971);
nand U19476 (N_19476,N_16486,N_16555);
nand U19477 (N_19477,N_16473,N_16598);
and U19478 (N_19478,N_16567,N_16256);
xor U19479 (N_19479,N_16358,N_16740);
and U19480 (N_19480,N_16693,N_16919);
nor U19481 (N_19481,N_18293,N_17590);
or U19482 (N_19482,N_16141,N_16149);
nor U19483 (N_19483,N_16109,N_18627);
nand U19484 (N_19484,N_17077,N_16527);
or U19485 (N_19485,N_17533,N_18116);
xnor U19486 (N_19486,N_18149,N_16760);
xor U19487 (N_19487,N_18722,N_16805);
and U19488 (N_19488,N_17968,N_16724);
nand U19489 (N_19489,N_18181,N_16694);
or U19490 (N_19490,N_18007,N_16519);
nor U19491 (N_19491,N_18683,N_17820);
nand U19492 (N_19492,N_16459,N_17569);
xnor U19493 (N_19493,N_17841,N_16800);
or U19494 (N_19494,N_18119,N_17382);
xor U19495 (N_19495,N_18584,N_16269);
xnor U19496 (N_19496,N_17945,N_17615);
xnor U19497 (N_19497,N_16701,N_17243);
or U19498 (N_19498,N_16808,N_18549);
or U19499 (N_19499,N_17919,N_17748);
xor U19500 (N_19500,N_15692,N_17530);
nor U19501 (N_19501,N_16862,N_17784);
nor U19502 (N_19502,N_15687,N_17500);
nor U19503 (N_19503,N_18472,N_16412);
and U19504 (N_19504,N_17521,N_18734);
xnor U19505 (N_19505,N_16087,N_17524);
nand U19506 (N_19506,N_16140,N_17105);
nand U19507 (N_19507,N_17599,N_18168);
and U19508 (N_19508,N_16028,N_18591);
nand U19509 (N_19509,N_15946,N_16988);
xor U19510 (N_19510,N_15826,N_16564);
nor U19511 (N_19511,N_16896,N_16985);
xor U19512 (N_19512,N_16188,N_18419);
nand U19513 (N_19513,N_15706,N_18307);
or U19514 (N_19514,N_18444,N_16854);
or U19515 (N_19515,N_15690,N_16751);
xnor U19516 (N_19516,N_16617,N_18395);
nor U19517 (N_19517,N_18566,N_17063);
xor U19518 (N_19518,N_16134,N_16055);
nor U19519 (N_19519,N_15739,N_18597);
and U19520 (N_19520,N_17859,N_16303);
or U19521 (N_19521,N_16801,N_17442);
nand U19522 (N_19522,N_17042,N_15855);
and U19523 (N_19523,N_18732,N_17729);
nor U19524 (N_19524,N_18619,N_16869);
or U19525 (N_19525,N_16496,N_15712);
or U19526 (N_19526,N_18064,N_18436);
nor U19527 (N_19527,N_16243,N_17689);
or U19528 (N_19528,N_17892,N_16721);
and U19529 (N_19529,N_18312,N_18221);
nand U19530 (N_19530,N_17683,N_16462);
nand U19531 (N_19531,N_16859,N_15990);
and U19532 (N_19532,N_15640,N_17324);
nor U19533 (N_19533,N_18716,N_16548);
xnor U19534 (N_19534,N_16917,N_16060);
and U19535 (N_19535,N_16275,N_18684);
nand U19536 (N_19536,N_16294,N_18663);
and U19537 (N_19537,N_15873,N_17195);
nor U19538 (N_19538,N_18265,N_18648);
or U19539 (N_19539,N_16615,N_16027);
and U19540 (N_19540,N_18078,N_15916);
or U19541 (N_19541,N_18124,N_18439);
and U19542 (N_19542,N_16980,N_16722);
and U19543 (N_19543,N_16901,N_15979);
or U19544 (N_19544,N_17649,N_17475);
nor U19545 (N_19545,N_18322,N_17482);
and U19546 (N_19546,N_18701,N_15628);
and U19547 (N_19547,N_16173,N_16377);
xnor U19548 (N_19548,N_18080,N_16216);
nand U19549 (N_19549,N_16049,N_18401);
and U19550 (N_19550,N_15824,N_16121);
nor U19551 (N_19551,N_16466,N_17169);
nor U19552 (N_19552,N_18032,N_16327);
or U19553 (N_19553,N_16779,N_16086);
and U19554 (N_19554,N_18474,N_18425);
or U19555 (N_19555,N_15852,N_17268);
nand U19556 (N_19556,N_15860,N_18455);
and U19557 (N_19557,N_16467,N_16850);
xor U19558 (N_19558,N_16572,N_18205);
or U19559 (N_19559,N_17885,N_15631);
nor U19560 (N_19560,N_15636,N_15633);
or U19561 (N_19561,N_17019,N_16457);
or U19562 (N_19562,N_18483,N_17359);
xnor U19563 (N_19563,N_16888,N_16409);
xor U19564 (N_19564,N_17410,N_16380);
or U19565 (N_19565,N_17869,N_18309);
nor U19566 (N_19566,N_18151,N_17792);
xor U19567 (N_19567,N_17467,N_16241);
nor U19568 (N_19568,N_15940,N_17518);
and U19569 (N_19569,N_17396,N_15680);
and U19570 (N_19570,N_18289,N_18266);
and U19571 (N_19571,N_16629,N_17479);
or U19572 (N_19572,N_16907,N_17056);
nand U19573 (N_19573,N_17749,N_17009);
xor U19574 (N_19574,N_15728,N_18008);
nand U19575 (N_19575,N_17601,N_16391);
xor U19576 (N_19576,N_15677,N_16450);
nor U19577 (N_19577,N_16480,N_18585);
or U19578 (N_19578,N_16291,N_17890);
nor U19579 (N_19579,N_15882,N_16848);
nor U19580 (N_19580,N_17320,N_16812);
nor U19581 (N_19581,N_16324,N_16010);
nand U19582 (N_19582,N_18582,N_16449);
xnor U19583 (N_19583,N_16936,N_16826);
xor U19584 (N_19584,N_17096,N_15969);
xnor U19585 (N_19585,N_18191,N_17589);
nand U19586 (N_19586,N_17851,N_16248);
and U19587 (N_19587,N_16239,N_18391);
nor U19588 (N_19588,N_16402,N_15794);
and U19589 (N_19589,N_18625,N_16731);
xor U19590 (N_19590,N_18318,N_16773);
or U19591 (N_19591,N_17004,N_18551);
or U19592 (N_19592,N_17055,N_16108);
nor U19593 (N_19593,N_18316,N_18533);
or U19594 (N_19594,N_15656,N_16120);
or U19595 (N_19595,N_16871,N_16675);
xnor U19596 (N_19596,N_17495,N_17658);
or U19597 (N_19597,N_18575,N_16396);
xor U19598 (N_19598,N_16711,N_16225);
nand U19599 (N_19599,N_15735,N_18294);
or U19600 (N_19600,N_17596,N_16966);
nor U19601 (N_19601,N_17949,N_15749);
xor U19602 (N_19602,N_17440,N_17415);
and U19603 (N_19603,N_16279,N_17549);
nor U19604 (N_19604,N_16332,N_16755);
or U19605 (N_19605,N_16803,N_16855);
or U19606 (N_19606,N_17678,N_17623);
and U19607 (N_19607,N_15710,N_16378);
and U19608 (N_19608,N_17470,N_18345);
nor U19609 (N_19609,N_15670,N_18206);
xnor U19610 (N_19610,N_16509,N_17568);
xnor U19611 (N_19611,N_16658,N_18705);
or U19612 (N_19612,N_17374,N_18275);
and U19613 (N_19613,N_16289,N_16337);
and U19614 (N_19614,N_16578,N_18606);
or U19615 (N_19615,N_18203,N_15854);
and U19616 (N_19616,N_17121,N_17917);
or U19617 (N_19617,N_16160,N_18355);
and U19618 (N_19618,N_16690,N_18317);
and U19619 (N_19619,N_17924,N_16276);
nor U19620 (N_19620,N_18653,N_18673);
nand U19621 (N_19621,N_15972,N_18607);
or U19622 (N_19622,N_16006,N_15888);
nand U19623 (N_19623,N_15911,N_16234);
nand U19624 (N_19624,N_16878,N_16948);
and U19625 (N_19625,N_16240,N_16329);
or U19626 (N_19626,N_17168,N_16894);
nand U19627 (N_19627,N_18162,N_17186);
and U19628 (N_19628,N_15836,N_16912);
nand U19629 (N_19629,N_17403,N_15931);
and U19630 (N_19630,N_17867,N_17791);
or U19631 (N_19631,N_18523,N_18602);
nand U19632 (N_19632,N_15921,N_16363);
xnor U19633 (N_19633,N_17767,N_16219);
nor U19634 (N_19634,N_18499,N_15912);
and U19635 (N_19635,N_17090,N_17639);
and U19636 (N_19636,N_16172,N_17339);
or U19637 (N_19637,N_15708,N_17273);
and U19638 (N_19638,N_16593,N_17455);
and U19639 (N_19639,N_17322,N_17747);
nand U19640 (N_19640,N_16036,N_18372);
xnor U19641 (N_19641,N_17777,N_15808);
xor U19642 (N_19642,N_17836,N_17329);
and U19643 (N_19643,N_17600,N_17260);
or U19644 (N_19644,N_16552,N_17785);
nor U19645 (N_19645,N_17261,N_15804);
nand U19646 (N_19646,N_18410,N_17474);
nand U19647 (N_19647,N_16430,N_17631);
xor U19648 (N_19648,N_16349,N_18556);
nor U19649 (N_19649,N_17787,N_16970);
and U19650 (N_19650,N_15831,N_18708);
or U19651 (N_19651,N_17812,N_17245);
xor U19652 (N_19652,N_16379,N_17389);
and U19653 (N_19653,N_16295,N_16717);
nor U19654 (N_19654,N_16277,N_17755);
nand U19655 (N_19655,N_16161,N_16080);
and U19656 (N_19656,N_17598,N_17849);
nor U19657 (N_19657,N_16991,N_17935);
nor U19658 (N_19658,N_17353,N_17838);
and U19659 (N_19659,N_16207,N_16185);
or U19660 (N_19660,N_15811,N_15634);
nand U19661 (N_19661,N_18044,N_17768);
nor U19662 (N_19662,N_16306,N_16647);
nor U19663 (N_19663,N_16143,N_16267);
xnor U19664 (N_19664,N_17434,N_18539);
xnor U19665 (N_19665,N_17633,N_17944);
nor U19666 (N_19666,N_17464,N_16392);
or U19667 (N_19667,N_17146,N_17672);
nor U19668 (N_19668,N_18045,N_15781);
or U19669 (N_19669,N_18120,N_16802);
nand U19670 (N_19670,N_16004,N_17896);
or U19671 (N_19671,N_17574,N_16428);
nor U19672 (N_19672,N_17909,N_18532);
or U19673 (N_19673,N_18441,N_15915);
or U19674 (N_19674,N_15863,N_17230);
and U19675 (N_19675,N_15754,N_15950);
nor U19676 (N_19676,N_16782,N_17811);
xor U19677 (N_19677,N_17405,N_17148);
xor U19678 (N_19678,N_17642,N_17429);
xor U19679 (N_19679,N_18495,N_16475);
and U19680 (N_19680,N_17795,N_18247);
or U19681 (N_19681,N_18694,N_16417);
or U19682 (N_19682,N_17013,N_16646);
and U19683 (N_19683,N_16454,N_17607);
or U19684 (N_19684,N_17900,N_15929);
nand U19685 (N_19685,N_17343,N_17874);
xnor U19686 (N_19686,N_17210,N_15845);
and U19687 (N_19687,N_18009,N_17266);
xnor U19688 (N_19688,N_17745,N_17794);
and U19689 (N_19689,N_16829,N_17277);
and U19690 (N_19690,N_15840,N_17932);
and U19691 (N_19691,N_15883,N_17809);
nand U19692 (N_19692,N_18544,N_18255);
and U19693 (N_19693,N_17394,N_18427);
xor U19694 (N_19694,N_18555,N_16867);
and U19695 (N_19695,N_17537,N_18002);
nor U19696 (N_19696,N_16574,N_15795);
xnor U19697 (N_19697,N_17710,N_18473);
and U19698 (N_19698,N_18020,N_17962);
or U19699 (N_19699,N_17291,N_16550);
xor U19700 (N_19700,N_16052,N_17094);
nand U19701 (N_19701,N_17414,N_17011);
xnor U19702 (N_19702,N_17583,N_16595);
xor U19703 (N_19703,N_15886,N_16190);
or U19704 (N_19704,N_17380,N_16621);
xnor U19705 (N_19705,N_17012,N_16914);
nand U19706 (N_19706,N_18174,N_17127);
and U19707 (N_19707,N_16357,N_17118);
xor U19708 (N_19708,N_16177,N_16229);
nor U19709 (N_19709,N_18577,N_15763);
xor U19710 (N_19710,N_16937,N_18327);
and U19711 (N_19711,N_17408,N_17337);
and U19712 (N_19712,N_16797,N_16863);
nor U19713 (N_19713,N_17057,N_16397);
xor U19714 (N_19714,N_18413,N_16860);
or U19715 (N_19715,N_18096,N_16296);
or U19716 (N_19716,N_17788,N_16416);
nand U19717 (N_19717,N_18380,N_17123);
nand U19718 (N_19718,N_16861,N_17244);
and U19719 (N_19719,N_16663,N_17696);
nand U19720 (N_19720,N_18621,N_16611);
nor U19721 (N_19721,N_16338,N_16642);
nand U19722 (N_19722,N_17232,N_15827);
and U19723 (N_19723,N_15632,N_17383);
xnor U19724 (N_19724,N_17167,N_18571);
xnor U19725 (N_19725,N_16603,N_16110);
or U19726 (N_19726,N_17298,N_18198);
nor U19727 (N_19727,N_15730,N_17690);
nand U19728 (N_19728,N_16769,N_17646);
and U19729 (N_19729,N_16789,N_15821);
or U19730 (N_19730,N_15976,N_16333);
nor U19731 (N_19731,N_15938,N_17637);
or U19732 (N_19732,N_16811,N_18725);
and U19733 (N_19733,N_16893,N_16007);
and U19734 (N_19734,N_16316,N_16816);
nand U19735 (N_19735,N_16905,N_17031);
nor U19736 (N_19736,N_16502,N_16193);
and U19737 (N_19737,N_18360,N_18736);
nor U19738 (N_19738,N_17447,N_16094);
nor U19739 (N_19739,N_18264,N_18458);
xor U19740 (N_19740,N_17390,N_15862);
or U19741 (N_19741,N_18160,N_18135);
or U19742 (N_19742,N_16833,N_17367);
nor U19743 (N_19743,N_15850,N_18620);
and U19744 (N_19744,N_17346,N_18398);
nor U19745 (N_19745,N_17047,N_18402);
nor U19746 (N_19746,N_18172,N_17889);
xnor U19747 (N_19747,N_16344,N_17654);
and U19748 (N_19748,N_18570,N_16510);
or U19749 (N_19749,N_18749,N_16877);
nor U19750 (N_19750,N_18558,N_18043);
or U19751 (N_19751,N_15675,N_18385);
nor U19752 (N_19752,N_18332,N_18670);
nand U19753 (N_19753,N_17813,N_17886);
nand U19754 (N_19754,N_17856,N_16168);
nor U19755 (N_19755,N_17227,N_16771);
and U19756 (N_19756,N_18171,N_18201);
nor U19757 (N_19757,N_17336,N_18182);
nand U19758 (N_19758,N_18161,N_17263);
nand U19759 (N_19759,N_16089,N_18490);
nand U19760 (N_19760,N_17975,N_15844);
nand U19761 (N_19761,N_16383,N_16471);
nand U19762 (N_19762,N_18016,N_18240);
nand U19763 (N_19763,N_16057,N_15949);
and U19764 (N_19764,N_16846,N_17154);
and U19765 (N_19765,N_18528,N_16610);
and U19766 (N_19766,N_16790,N_17606);
nor U19767 (N_19767,N_15671,N_16786);
or U19768 (N_19768,N_17915,N_16517);
xnor U19769 (N_19769,N_17780,N_18476);
nor U19770 (N_19770,N_17970,N_18260);
xnor U19771 (N_19771,N_18237,N_17958);
and U19772 (N_19772,N_17592,N_15942);
nand U19773 (N_19773,N_18254,N_16011);
and U19774 (N_19774,N_17547,N_17181);
and U19775 (N_19775,N_17756,N_16339);
and U19776 (N_19776,N_18111,N_16742);
or U19777 (N_19777,N_15978,N_16009);
xor U19778 (N_19778,N_17147,N_17340);
xor U19779 (N_19779,N_17963,N_16886);
nor U19780 (N_19780,N_15853,N_18100);
nand U19781 (N_19781,N_15849,N_17254);
xor U19782 (N_19782,N_16274,N_17609);
nand U19783 (N_19783,N_18261,N_18241);
nand U19784 (N_19784,N_15813,N_16504);
and U19785 (N_19785,N_16326,N_15988);
xor U19786 (N_19786,N_17357,N_15659);
nor U19787 (N_19787,N_15867,N_18477);
or U19788 (N_19788,N_16468,N_18073);
nor U19789 (N_19789,N_17994,N_17594);
xor U19790 (N_19790,N_16685,N_17222);
and U19791 (N_19791,N_16739,N_17744);
xnor U19792 (N_19792,N_16709,N_15835);
nor U19793 (N_19793,N_17132,N_16228);
nand U19794 (N_19794,N_16250,N_16508);
and U19795 (N_19795,N_17362,N_17852);
and U19796 (N_19796,N_15892,N_17728);
xor U19797 (N_19797,N_16164,N_15757);
nand U19798 (N_19798,N_18188,N_16310);
nand U19799 (N_19799,N_17153,N_18178);
or U19800 (N_19800,N_16431,N_17905);
or U19801 (N_19801,N_15798,N_17891);
and U19802 (N_19802,N_18146,N_16892);
xnor U19803 (N_19803,N_17933,N_17418);
or U19804 (N_19804,N_15761,N_17002);
or U19805 (N_19805,N_17871,N_16823);
and U19806 (N_19806,N_17341,N_17732);
or U19807 (N_19807,N_16640,N_16347);
nand U19808 (N_19808,N_15638,N_16674);
and U19809 (N_19809,N_16425,N_17484);
nor U19810 (N_19810,N_16972,N_16885);
nor U19811 (N_19811,N_17398,N_18034);
nand U19812 (N_19812,N_16095,N_16123);
and U19813 (N_19813,N_16706,N_16398);
nand U19814 (N_19814,N_17536,N_16526);
xnor U19815 (N_19815,N_16374,N_15965);
xor U19816 (N_19816,N_18227,N_15736);
xor U19817 (N_19817,N_17773,N_16213);
xor U19818 (N_19818,N_17387,N_18542);
nand U19819 (N_19819,N_16194,N_16839);
nor U19820 (N_19820,N_17704,N_17863);
xnor U19821 (N_19821,N_16520,N_15625);
or U19822 (N_19822,N_17219,N_16544);
or U19823 (N_19823,N_16904,N_16033);
nand U19824 (N_19824,N_17173,N_16540);
or U19825 (N_19825,N_15848,N_17929);
and U19826 (N_19826,N_18552,N_17435);
nand U19827 (N_19827,N_15767,N_18253);
or U19828 (N_19828,N_18004,N_17370);
nand U19829 (N_19829,N_18342,N_17170);
nand U19830 (N_19830,N_18381,N_16423);
or U19831 (N_19831,N_17753,N_17140);
or U19832 (N_19832,N_16996,N_17458);
or U19833 (N_19833,N_17010,N_17477);
nor U19834 (N_19834,N_17338,N_16563);
nor U19835 (N_19835,N_17868,N_16226);
xor U19836 (N_19836,N_18728,N_18680);
or U19837 (N_19837,N_18170,N_16609);
xor U19838 (N_19838,N_18231,N_15658);
and U19839 (N_19839,N_17014,N_17103);
nand U19840 (N_19840,N_17221,N_16054);
and U19841 (N_19841,N_17069,N_18738);
nand U19842 (N_19842,N_16002,N_18660);
and U19843 (N_19843,N_18326,N_16280);
nor U19844 (N_19844,N_16999,N_18306);
xnor U19845 (N_19845,N_18498,N_16364);
xor U19846 (N_19846,N_17789,N_17264);
nor U19847 (N_19847,N_16832,N_18295);
nor U19848 (N_19848,N_17685,N_18109);
or U19849 (N_19849,N_18068,N_16671);
nor U19850 (N_19850,N_17940,N_16203);
nand U19851 (N_19851,N_17431,N_15982);
xor U19852 (N_19852,N_16100,N_18278);
and U19853 (N_19853,N_18721,N_16411);
nand U19854 (N_19854,N_16038,N_17231);
or U19855 (N_19855,N_18723,N_17731);
nor U19856 (N_19856,N_17397,N_18704);
xnor U19857 (N_19857,N_17740,N_16208);
and U19858 (N_19858,N_16154,N_15784);
nand U19859 (N_19859,N_16499,N_18696);
nor U19860 (N_19860,N_16312,N_17947);
or U19861 (N_19861,N_17028,N_18263);
nand U19862 (N_19862,N_15745,N_17957);
xnor U19863 (N_19863,N_18527,N_18243);
xor U19864 (N_19864,N_17866,N_17969);
and U19865 (N_19865,N_17563,N_17655);
nand U19866 (N_19866,N_17129,N_17993);
and U19867 (N_19867,N_17229,N_18737);
nor U19868 (N_19868,N_16254,N_16781);
or U19869 (N_19869,N_17956,N_17571);
or U19870 (N_19870,N_16195,N_16433);
and U19871 (N_19871,N_18122,N_18272);
or U19872 (N_19872,N_16040,N_16865);
nand U19873 (N_19873,N_15966,N_17734);
and U19874 (N_19874,N_17108,N_17384);
nand U19875 (N_19875,N_17965,N_17488);
or U19876 (N_19876,N_16318,N_15726);
or U19877 (N_19877,N_17516,N_16924);
nor U19878 (N_19878,N_16513,N_16968);
nor U19879 (N_19879,N_18517,N_17826);
or U19880 (N_19880,N_17351,N_17293);
or U19881 (N_19881,N_18642,N_17865);
nand U19882 (N_19882,N_17233,N_17712);
xnor U19883 (N_19883,N_18194,N_16032);
nor U19884 (N_19884,N_18541,N_15758);
and U19885 (N_19885,N_16873,N_17700);
nand U19886 (N_19886,N_17363,N_16791);
xnor U19887 (N_19887,N_16375,N_16824);
nand U19888 (N_19888,N_17369,N_17465);
nor U19889 (N_19889,N_16003,N_18687);
and U19890 (N_19890,N_15691,N_16596);
xnor U19891 (N_19891,N_18022,N_16556);
and U19892 (N_19892,N_17422,N_18050);
and U19893 (N_19893,N_18176,N_18226);
or U19894 (N_19894,N_15830,N_17294);
nand U19895 (N_19895,N_15962,N_18488);
xor U19896 (N_19896,N_18543,N_18576);
nand U19897 (N_19897,N_17305,N_15865);
nor U19898 (N_19898,N_16619,N_16673);
nand U19899 (N_19899,N_16633,N_16313);
xnor U19900 (N_19900,N_16716,N_16404);
and U19901 (N_19901,N_18152,N_17352);
or U19902 (N_19902,N_15802,N_17725);
nor U19903 (N_19903,N_16788,N_17643);
nand U19904 (N_19904,N_17546,N_18187);
or U19905 (N_19905,N_18378,N_15783);
nand U19906 (N_19906,N_18041,N_17824);
and U19907 (N_19907,N_18128,N_17347);
or U19908 (N_19908,N_16315,N_16118);
nor U19909 (N_19909,N_16342,N_17783);
or U19910 (N_19910,N_15803,N_15655);
xor U19911 (N_19911,N_17224,N_17124);
nor U19912 (N_19912,N_16505,N_16158);
nand U19913 (N_19913,N_16947,N_16682);
nand U19914 (N_19914,N_17714,N_17059);
or U19915 (N_19915,N_17952,N_17122);
and U19916 (N_19916,N_18081,N_18280);
xnor U19917 (N_19917,N_17421,N_17379);
or U19918 (N_19918,N_17861,N_17772);
xor U19919 (N_19919,N_18613,N_15701);
nor U19920 (N_19920,N_16681,N_15948);
xnor U19921 (N_19921,N_18006,N_18214);
nor U19922 (N_19922,N_17463,N_17565);
or U19923 (N_19923,N_15717,N_18592);
or U19924 (N_19924,N_16997,N_17927);
and U19925 (N_19925,N_17752,N_16444);
nand U19926 (N_19926,N_15661,N_17135);
xnor U19927 (N_19927,N_16656,N_16616);
nor U19928 (N_19928,N_18105,N_15905);
nor U19929 (N_19929,N_16442,N_16266);
xor U19930 (N_19930,N_17211,N_16210);
and U19931 (N_19931,N_18748,N_17873);
nand U19932 (N_19932,N_18095,N_15799);
and U19933 (N_19933,N_18179,N_15700);
and U19934 (N_19934,N_16198,N_18093);
or U19935 (N_19935,N_17239,N_16099);
and U19936 (N_19936,N_17644,N_18113);
and U19937 (N_19937,N_17834,N_18356);
or U19938 (N_19938,N_17076,N_15793);
nand U19939 (N_19939,N_16085,N_15729);
xnor U19940 (N_19940,N_16961,N_18707);
nand U19941 (N_19941,N_17995,N_18220);
xnor U19942 (N_19942,N_18479,N_17060);
nor U19943 (N_19943,N_18612,N_18175);
xor U19944 (N_19944,N_17319,N_18579);
nand U19945 (N_19945,N_18666,N_15644);
or U19946 (N_19946,N_16916,N_16729);
or U19947 (N_19947,N_17538,N_17029);
and U19948 (N_19948,N_16949,N_16868);
nand U19949 (N_19949,N_16399,N_15866);
or U19950 (N_19950,N_16965,N_17248);
xnor U19951 (N_19951,N_18329,N_16231);
nand U19952 (N_19952,N_17275,N_15993);
or U19953 (N_19953,N_18085,N_16979);
nor U19954 (N_19954,N_18320,N_17641);
and U19955 (N_19955,N_18641,N_17145);
nor U19956 (N_19956,N_17966,N_15828);
and U19957 (N_19957,N_17196,N_17502);
nor U19958 (N_19958,N_16607,N_15987);
nor U19959 (N_19959,N_17015,N_16664);
xor U19960 (N_19960,N_15814,N_17226);
nand U19961 (N_19961,N_18510,N_16115);
xor U19962 (N_19962,N_15727,N_16668);
nor U19963 (N_19963,N_18084,N_17698);
xor U19964 (N_19964,N_15626,N_17640);
or U19965 (N_19965,N_17151,N_18733);
xnor U19966 (N_19966,N_17062,N_17381);
and U19967 (N_19967,N_16035,N_17318);
or U19968 (N_19968,N_16437,N_16214);
or U19969 (N_19969,N_15989,N_15887);
and U19970 (N_19970,N_15686,N_18234);
xnor U19971 (N_19971,N_17159,N_17259);
nand U19972 (N_19972,N_18484,N_15925);
or U19973 (N_19973,N_15973,N_17427);
nand U19974 (N_19974,N_16600,N_17635);
nand U19975 (N_19975,N_17895,N_17241);
and U19976 (N_19976,N_15926,N_17762);
nor U19977 (N_19977,N_15958,N_16915);
and U19978 (N_19978,N_15919,N_16944);
nand U19979 (N_19979,N_16636,N_16528);
or U19980 (N_19980,N_15660,N_16441);
nor U19981 (N_19981,N_17097,N_18348);
nor U19982 (N_19982,N_15769,N_16577);
and U19983 (N_19983,N_17401,N_16354);
nand U19984 (N_19984,N_18422,N_17335);
nor U19985 (N_19985,N_16436,N_17373);
nand U19986 (N_19986,N_16205,N_16238);
or U19987 (N_19987,N_16029,N_17567);
nand U19988 (N_19988,N_18299,N_17130);
nor U19989 (N_19989,N_16175,N_16670);
or U19990 (N_19990,N_15740,N_18114);
nor U19991 (N_19991,N_18123,N_18070);
xor U19992 (N_19992,N_18494,N_18587);
xnor U19993 (N_19993,N_18300,N_17494);
nand U19994 (N_19994,N_16495,N_16390);
nand U19995 (N_19995,N_18195,N_18331);
nor U19996 (N_19996,N_17881,N_18537);
or U19997 (N_19997,N_17237,N_18075);
or U19998 (N_19998,N_18150,N_16535);
and U19999 (N_19999,N_15901,N_16813);
nor U20000 (N_20000,N_18466,N_18373);
nand U20001 (N_20001,N_15900,N_16689);
nor U20002 (N_20002,N_15662,N_16314);
and U20003 (N_20003,N_16730,N_16546);
or U20004 (N_20004,N_17503,N_18675);
or U20005 (N_20005,N_16013,N_18030);
or U20006 (N_20006,N_17242,N_17845);
nor U20007 (N_20007,N_17313,N_18630);
xor U20008 (N_20008,N_18321,N_17152);
nand U20009 (N_20009,N_16951,N_15880);
or U20010 (N_20010,N_15682,N_18482);
and U20011 (N_20011,N_17143,N_15719);
nand U20012 (N_20012,N_15696,N_15673);
nand U20013 (N_20013,N_16182,N_16727);
or U20014 (N_20014,N_17991,N_16536);
or U20015 (N_20015,N_17723,N_17089);
and U20016 (N_20016,N_16891,N_18611);
nand U20017 (N_20017,N_16554,N_15684);
or U20018 (N_20018,N_17314,N_17911);
nor U20019 (N_20019,N_16986,N_18367);
and U20020 (N_20020,N_16799,N_18681);
nor U20021 (N_20021,N_16367,N_17068);
and U20022 (N_20022,N_16581,N_16093);
nor U20023 (N_20023,N_16376,N_16558);
or U20024 (N_20024,N_17837,N_18614);
nor U20025 (N_20025,N_18283,N_18258);
nor U20026 (N_20026,N_16748,N_18647);
nand U20027 (N_20027,N_17075,N_17597);
and U20028 (N_20028,N_18284,N_17262);
nor U20029 (N_20029,N_18656,N_15766);
nor U20030 (N_20030,N_17535,N_17361);
or U20031 (N_20031,N_16820,N_18274);
nand U20032 (N_20032,N_16365,N_16113);
xnor U20033 (N_20033,N_16720,N_15681);
nor U20034 (N_20034,N_17283,N_17833);
and U20035 (N_20035,N_16174,N_17922);
or U20036 (N_20036,N_18051,N_16227);
xor U20037 (N_20037,N_18037,N_17910);
nor U20038 (N_20038,N_18088,N_15898);
nor U20039 (N_20039,N_16133,N_15974);
nor U20040 (N_20040,N_17522,N_18685);
and U20041 (N_20041,N_18393,N_17760);
nand U20042 (N_20042,N_17323,N_16472);
or U20043 (N_20043,N_18406,N_17974);
xnor U20044 (N_20044,N_16056,N_16481);
and U20045 (N_20045,N_16562,N_18058);
or U20046 (N_20046,N_15725,N_17657);
xor U20047 (N_20047,N_18210,N_17504);
and U20048 (N_20048,N_16343,N_18035);
or U20049 (N_20049,N_17110,N_16831);
and U20050 (N_20050,N_15843,N_17449);
nand U20051 (N_20051,N_18678,N_18270);
or U20052 (N_20052,N_17131,N_16155);
nor U20053 (N_20053,N_16030,N_18668);
and U20054 (N_20054,N_17510,N_18646);
nor U20055 (N_20055,N_15642,N_16977);
nor U20056 (N_20056,N_16298,N_16282);
and U20057 (N_20057,N_15702,N_16652);
or U20058 (N_20058,N_16752,N_15977);
xor U20059 (N_20059,N_17058,N_18047);
and U20060 (N_20060,N_18148,N_17534);
xnor U20061 (N_20061,N_18616,N_15786);
or U20062 (N_20062,N_17906,N_16405);
nand U20063 (N_20063,N_18094,N_15981);
and U20064 (N_20064,N_18442,N_15744);
or U20065 (N_20065,N_17595,N_18711);
or U20066 (N_20066,N_17409,N_18462);
or U20067 (N_20067,N_16059,N_18138);
nor U20068 (N_20068,N_15997,N_18208);
nand U20069 (N_20069,N_18382,N_18545);
and U20070 (N_20070,N_16119,N_16331);
nand U20071 (N_20071,N_18471,N_16171);
xor U20072 (N_20072,N_18057,N_17674);
nand U20073 (N_20073,N_18190,N_17573);
or U20074 (N_20074,N_16176,N_15822);
and U20075 (N_20075,N_18709,N_18437);
nor U20076 (N_20076,N_17782,N_17816);
xnor U20077 (N_20077,N_18689,N_17997);
nand U20078 (N_20078,N_17344,N_16683);
nand U20079 (N_20079,N_17878,N_16849);
nand U20080 (N_20080,N_17613,N_18743);
nand U20081 (N_20081,N_16346,N_18245);
xnor U20082 (N_20082,N_17950,N_18165);
and U20083 (N_20083,N_18415,N_16518);
or U20084 (N_20084,N_15669,N_16019);
nor U20085 (N_20085,N_16560,N_16048);
nor U20086 (N_20086,N_17354,N_17120);
nor U20087 (N_20087,N_18589,N_15705);
nor U20088 (N_20088,N_18218,N_16584);
and U20089 (N_20089,N_16910,N_16461);
nor U20090 (N_20090,N_17070,N_16001);
or U20091 (N_20091,N_16249,N_16051);
nor U20092 (N_20092,N_17916,N_15913);
and U20093 (N_20093,N_17972,N_17688);
nand U20094 (N_20094,N_16128,N_17682);
nor U20095 (N_20095,N_18092,N_16360);
xor U20096 (N_20096,N_17584,N_18561);
xnor U20097 (N_20097,N_15907,N_16498);
or U20098 (N_20098,N_16958,N_16547);
and U20099 (N_20099,N_17295,N_15649);
xnor U20100 (N_20100,N_17559,N_17808);
nor U20101 (N_20101,N_16661,N_16098);
nor U20102 (N_20102,N_16237,N_18615);
nand U20103 (N_20103,N_16232,N_16482);
nand U20104 (N_20104,N_18108,N_16455);
nor U20105 (N_20105,N_16687,N_17205);
nand U20106 (N_20106,N_16090,N_17385);
nor U20107 (N_20107,N_17321,N_17715);
or U20108 (N_20108,N_17669,N_16259);
and U20109 (N_20109,N_15878,N_16286);
xnor U20110 (N_20110,N_16819,N_17898);
nor U20111 (N_20111,N_16953,N_18520);
and U20112 (N_20112,N_15906,N_17428);
xor U20113 (N_20113,N_16606,N_15753);
nand U20114 (N_20114,N_17179,N_16523);
nor U20115 (N_20115,N_17238,N_17694);
and U20116 (N_20116,N_17348,N_18478);
xnor U20117 (N_20117,N_15641,N_18438);
xor U20118 (N_20118,N_18581,N_18665);
xor U20119 (N_20119,N_16283,N_18699);
nand U20120 (N_20120,N_15778,N_18420);
and U20121 (N_20121,N_17388,N_15651);
and U20122 (N_20122,N_18574,N_18550);
nor U20123 (N_20123,N_17433,N_16920);
or U20124 (N_20124,N_18235,N_18062);
and U20125 (N_20125,N_15917,N_15945);
or U20126 (N_20126,N_17666,N_17738);
nand U20127 (N_20127,N_15774,N_16793);
or U20128 (N_20128,N_16025,N_18400);
and U20129 (N_20129,N_16989,N_17652);
or U20130 (N_20130,N_16738,N_17332);
or U20131 (N_20131,N_18159,N_16261);
nand U20132 (N_20132,N_17967,N_15984);
xor U20133 (N_20133,N_17511,N_17424);
nor U20134 (N_20134,N_15903,N_17588);
xor U20135 (N_20135,N_16062,N_17199);
xor U20136 (N_20136,N_16734,N_16179);
nor U20137 (N_20137,N_17191,N_16545);
and U20138 (N_20138,N_17509,N_18336);
and U20139 (N_20139,N_15674,N_17190);
or U20140 (N_20140,N_17161,N_17253);
nor U20141 (N_20141,N_16413,N_17450);
or U20142 (N_20142,N_18505,N_17936);
and U20143 (N_20143,N_17269,N_15818);
or U20144 (N_20144,N_15629,N_16406);
and U20145 (N_20145,N_18353,N_17471);
nor U20146 (N_20146,N_15707,N_18262);
and U20147 (N_20147,N_16137,N_16745);
xnor U20148 (N_20148,N_15664,N_15697);
nand U20149 (N_20149,N_17441,N_18386);
and U20150 (N_20150,N_17468,N_16356);
nand U20151 (N_20151,N_17206,N_16946);
xor U20152 (N_20152,N_18586,N_16144);
xor U20153 (N_20153,N_16483,N_16608);
xnor U20154 (N_20154,N_17107,N_16388);
nand U20155 (N_20155,N_18027,N_16866);
nor U20156 (N_20156,N_18207,N_16834);
or U20157 (N_20157,N_15663,N_15746);
or U20158 (N_20158,N_17548,N_18005);
and U20159 (N_20159,N_16744,N_16299);
xnor U20160 (N_20160,N_17098,N_16092);
xor U20161 (N_20161,N_18399,N_17093);
and U20162 (N_20162,N_15765,N_18250);
nor U20163 (N_20163,N_18740,N_17713);
or U20164 (N_20164,N_18741,N_17033);
xor U20165 (N_20165,N_18033,N_18536);
nor U20166 (N_20166,N_16000,N_16759);
nand U20167 (N_20167,N_17634,N_18649);
nor U20168 (N_20168,N_18501,N_16928);
xnor U20169 (N_20169,N_17171,N_15875);
or U20170 (N_20170,N_18134,N_16424);
xnor U20171 (N_20171,N_18222,N_15756);
nor U20172 (N_20172,N_18053,N_17139);
nand U20173 (N_20173,N_16592,N_18500);
nand U20174 (N_20174,N_17137,N_16081);
nor U20175 (N_20175,N_18480,N_18281);
or U20176 (N_20176,N_16245,N_16525);
and U20177 (N_20177,N_15872,N_18183);
xnor U20178 (N_20178,N_15639,N_18431);
nor U20179 (N_20179,N_18189,N_16432);
nand U20180 (N_20180,N_18524,N_15967);
nor U20181 (N_20181,N_18546,N_16293);
or U20182 (N_20182,N_18714,N_17234);
nand U20183 (N_20183,N_18363,N_15959);
and U20184 (N_20184,N_17670,N_15773);
nor U20185 (N_20185,N_16131,N_16507);
xnor U20186 (N_20186,N_16625,N_17419);
nand U20187 (N_20187,N_15889,N_16959);
nand U20188 (N_20188,N_15776,N_16485);
or U20189 (N_20189,N_18059,N_17604);
or U20190 (N_20190,N_16934,N_16075);
nand U20191 (N_20191,N_17946,N_15771);
and U20192 (N_20192,N_16264,N_17085);
nor U20193 (N_20193,N_18038,N_18219);
nor U20194 (N_20194,N_18407,N_18132);
nor U20195 (N_20195,N_17998,N_17621);
or U20196 (N_20196,N_15839,N_16069);
or U20197 (N_20197,N_17815,N_15851);
nand U20198 (N_20198,N_16150,N_18580);
and U20199 (N_20199,N_16880,N_17438);
xnor U20200 (N_20200,N_18643,N_17240);
xor U20201 (N_20201,N_17854,N_16159);
nand U20202 (N_20202,N_15791,N_16065);
or U20203 (N_20203,N_16530,N_18440);
and U20204 (N_20204,N_17763,N_16757);
or U20205 (N_20205,N_17628,N_15952);
and U20206 (N_20206,N_17616,N_16440);
nand U20207 (N_20207,N_17942,N_15983);
xnor U20208 (N_20208,N_17724,N_15732);
or U20209 (N_20209,N_16022,N_17746);
xor U20210 (N_20210,N_16255,N_18515);
nand U20211 (N_20211,N_17008,N_16902);
and U20212 (N_20212,N_17490,N_17839);
nor U20213 (N_20213,N_18491,N_18521);
or U20214 (N_20214,N_18598,N_17017);
and U20215 (N_20215,N_17679,N_18557);
and U20216 (N_20216,N_16776,N_18469);
or U20217 (N_20217,N_15722,N_15790);
xnor U20218 (N_20218,N_17459,N_16645);
nand U20219 (N_20219,N_15934,N_16487);
nor U20220 (N_20220,N_18417,N_17086);
nor U20221 (N_20221,N_15751,N_15861);
nor U20222 (N_20222,N_18672,N_17959);
nor U20223 (N_20223,N_16212,N_16477);
and U20224 (N_20224,N_17292,N_16130);
xnor U20225 (N_20225,N_18106,N_17554);
nor U20226 (N_20226,N_18158,N_16784);
or U20227 (N_20227,N_16169,N_17532);
nand U20228 (N_20228,N_16448,N_17720);
or U20229 (N_20229,N_16710,N_15939);
xnor U20230 (N_20230,N_17702,N_17716);
and U20231 (N_20231,N_18426,N_17948);
xor U20232 (N_20232,N_16678,N_18136);
nand U20233 (N_20233,N_18658,N_17848);
or U20234 (N_20234,N_18371,N_16491);
xnor U20235 (N_20235,N_17207,N_17312);
xnor U20236 (N_20236,N_17189,N_18199);
nand U20237 (N_20237,N_18486,N_16235);
nand U20238 (N_20238,N_15896,N_17618);
or U20239 (N_20239,N_15819,N_15829);
or U20240 (N_20240,N_18578,N_15846);
nor U20241 (N_20241,N_16201,N_15823);
nor U20242 (N_20242,N_16561,N_17761);
or U20243 (N_20243,N_17342,N_15713);
nor U20244 (N_20244,N_16474,N_15723);
or U20245 (N_20245,N_18102,N_18090);
nor U20246 (N_20246,N_17311,N_15881);
nor U20247 (N_20247,N_18502,N_18077);
nor U20248 (N_20248,N_18618,N_18335);
xnor U20249 (N_20249,N_18304,N_16627);
and U20250 (N_20250,N_16707,N_17733);
nand U20251 (N_20251,N_18573,N_17092);
nand U20252 (N_20252,N_18286,N_15683);
and U20253 (N_20253,N_16272,N_18277);
nand U20254 (N_20254,N_15792,N_15947);
xnor U20255 (N_20255,N_17472,N_18682);
or U20256 (N_20256,N_18601,N_15635);
xnor U20257 (N_20257,N_18384,N_16107);
nor U20258 (N_20258,N_17289,N_16835);
nand U20259 (N_20259,N_17593,N_17552);
xnor U20260 (N_20260,N_16735,N_16426);
or U20261 (N_20261,N_17478,N_17721);
xnor U20262 (N_20262,N_17476,N_17473);
nand U20263 (N_20263,N_15920,N_16843);
nor U20264 (N_20264,N_16768,N_18244);
nand U20265 (N_20265,N_18287,N_18347);
and U20266 (N_20266,N_17395,N_18710);
xor U20267 (N_20267,N_16328,N_17134);
xnor U20268 (N_20268,N_18223,N_16497);
nor U20269 (N_20269,N_17176,N_17591);
and U20270 (N_20270,N_17330,N_15869);
nand U20271 (N_20271,N_16570,N_18028);
xor U20272 (N_20272,N_17605,N_17858);
xor U20273 (N_20273,N_17943,N_16575);
xnor U20274 (N_20274,N_16135,N_17481);
nor U20275 (N_20275,N_16696,N_15874);
xor U20276 (N_20276,N_16408,N_18713);
and U20277 (N_20277,N_17285,N_16126);
and U20278 (N_20278,N_16565,N_16984);
nor U20279 (N_20279,N_18634,N_16807);
or U20280 (N_20280,N_18430,N_18446);
xnor U20281 (N_20281,N_16794,N_18074);
or U20282 (N_20282,N_16125,N_16414);
nor U20283 (N_20283,N_18506,N_17102);
nor U20284 (N_20284,N_18204,N_15760);
xor U20285 (N_20285,N_17065,N_17610);
nand U20286 (N_20286,N_17501,N_18631);
and U20287 (N_20287,N_17150,N_16320);
or U20288 (N_20288,N_18097,N_18688);
nand U20289 (N_20289,N_17603,N_15714);
xor U20290 (N_20290,N_18079,N_17798);
or U20291 (N_20291,N_16960,N_16178);
and U20292 (N_20292,N_16403,N_16456);
and U20293 (N_20293,N_16083,N_17088);
and U20294 (N_20294,N_15801,N_16319);
xnor U20295 (N_20295,N_18099,N_18409);
xor U20296 (N_20296,N_16321,N_17693);
nor U20297 (N_20297,N_17083,N_16847);
and U20298 (N_20298,N_18267,N_16008);
xor U20299 (N_20299,N_16105,N_16088);
xor U20300 (N_20300,N_18691,N_15805);
nand U20301 (N_20301,N_15876,N_17162);
nor U20302 (N_20302,N_17709,N_15785);
nor U20303 (N_20303,N_16881,N_18319);
nand U20304 (N_20304,N_16766,N_15884);
nor U20305 (N_20305,N_17053,N_17555);
or U20306 (N_20306,N_16084,N_17039);
nor U20307 (N_20307,N_18679,N_17512);
or U20308 (N_20308,N_18388,N_15772);
nor U20309 (N_20309,N_16747,N_16500);
xor U20310 (N_20310,N_17018,N_17182);
nor U20311 (N_20311,N_17739,N_16718);
nor U20312 (N_20312,N_16287,N_15760);
xor U20313 (N_20313,N_16960,N_15734);
xor U20314 (N_20314,N_17036,N_17447);
nor U20315 (N_20315,N_16983,N_17412);
nand U20316 (N_20316,N_18423,N_18739);
nor U20317 (N_20317,N_16199,N_18019);
or U20318 (N_20318,N_16997,N_18678);
nand U20319 (N_20319,N_18150,N_18720);
and U20320 (N_20320,N_18053,N_18339);
nor U20321 (N_20321,N_15991,N_16431);
and U20322 (N_20322,N_17390,N_18142);
nor U20323 (N_20323,N_17155,N_16630);
and U20324 (N_20324,N_15995,N_17174);
nor U20325 (N_20325,N_17054,N_18288);
nor U20326 (N_20326,N_18487,N_16936);
or U20327 (N_20327,N_15994,N_18212);
and U20328 (N_20328,N_18056,N_16437);
nand U20329 (N_20329,N_17691,N_15946);
nor U20330 (N_20330,N_18359,N_16916);
nor U20331 (N_20331,N_16045,N_15747);
and U20332 (N_20332,N_17014,N_17425);
and U20333 (N_20333,N_18656,N_16008);
and U20334 (N_20334,N_17068,N_18408);
and U20335 (N_20335,N_15891,N_16090);
nor U20336 (N_20336,N_16727,N_18249);
nor U20337 (N_20337,N_17700,N_16595);
nand U20338 (N_20338,N_15934,N_15799);
nor U20339 (N_20339,N_17650,N_15736);
nor U20340 (N_20340,N_16816,N_18278);
and U20341 (N_20341,N_18354,N_16748);
and U20342 (N_20342,N_17843,N_16238);
xnor U20343 (N_20343,N_16898,N_16547);
nand U20344 (N_20344,N_17688,N_18110);
and U20345 (N_20345,N_17840,N_16384);
or U20346 (N_20346,N_18137,N_17761);
nand U20347 (N_20347,N_17410,N_16076);
xnor U20348 (N_20348,N_18733,N_16257);
or U20349 (N_20349,N_16123,N_18314);
and U20350 (N_20350,N_18078,N_15895);
nor U20351 (N_20351,N_17369,N_17381);
nand U20352 (N_20352,N_17634,N_17759);
or U20353 (N_20353,N_15954,N_18734);
and U20354 (N_20354,N_16155,N_16758);
and U20355 (N_20355,N_17038,N_18205);
xnor U20356 (N_20356,N_17367,N_17747);
nor U20357 (N_20357,N_16264,N_18561);
xnor U20358 (N_20358,N_18113,N_17530);
nand U20359 (N_20359,N_17063,N_18228);
nand U20360 (N_20360,N_17735,N_16154);
nor U20361 (N_20361,N_17527,N_17747);
or U20362 (N_20362,N_17145,N_17806);
nand U20363 (N_20363,N_18363,N_16737);
nand U20364 (N_20364,N_17788,N_17152);
and U20365 (N_20365,N_17704,N_17956);
nor U20366 (N_20366,N_16897,N_18030);
and U20367 (N_20367,N_16637,N_17102);
and U20368 (N_20368,N_16881,N_16777);
xor U20369 (N_20369,N_16099,N_17747);
xor U20370 (N_20370,N_17728,N_17874);
or U20371 (N_20371,N_17307,N_17411);
nand U20372 (N_20372,N_15952,N_15666);
nor U20373 (N_20373,N_17073,N_16932);
xnor U20374 (N_20374,N_18306,N_17058);
and U20375 (N_20375,N_17460,N_16976);
or U20376 (N_20376,N_18734,N_18351);
nand U20377 (N_20377,N_17569,N_16686);
xnor U20378 (N_20378,N_16636,N_16527);
or U20379 (N_20379,N_16343,N_16900);
or U20380 (N_20380,N_18451,N_18657);
or U20381 (N_20381,N_16258,N_18027);
nor U20382 (N_20382,N_15737,N_16570);
xnor U20383 (N_20383,N_17146,N_16519);
nand U20384 (N_20384,N_15659,N_16090);
nand U20385 (N_20385,N_16977,N_17092);
nor U20386 (N_20386,N_16058,N_18021);
xor U20387 (N_20387,N_17584,N_17618);
nand U20388 (N_20388,N_15805,N_17678);
xor U20389 (N_20389,N_16767,N_16108);
nand U20390 (N_20390,N_16431,N_17967);
or U20391 (N_20391,N_18054,N_15669);
and U20392 (N_20392,N_17202,N_17162);
and U20393 (N_20393,N_17507,N_18697);
or U20394 (N_20394,N_16142,N_17038);
xnor U20395 (N_20395,N_15657,N_15683);
or U20396 (N_20396,N_15667,N_16162);
xor U20397 (N_20397,N_15677,N_17146);
or U20398 (N_20398,N_17286,N_18099);
or U20399 (N_20399,N_16312,N_16672);
nand U20400 (N_20400,N_15903,N_16249);
xor U20401 (N_20401,N_18618,N_16329);
nor U20402 (N_20402,N_17667,N_18558);
nor U20403 (N_20403,N_15790,N_16179);
and U20404 (N_20404,N_18193,N_18662);
nor U20405 (N_20405,N_16268,N_16823);
or U20406 (N_20406,N_17604,N_18649);
nand U20407 (N_20407,N_17892,N_17088);
nor U20408 (N_20408,N_15810,N_17241);
or U20409 (N_20409,N_17011,N_16625);
nand U20410 (N_20410,N_17165,N_15725);
nand U20411 (N_20411,N_18309,N_17629);
or U20412 (N_20412,N_18697,N_17133);
xnor U20413 (N_20413,N_17747,N_18513);
xnor U20414 (N_20414,N_15804,N_16397);
or U20415 (N_20415,N_17705,N_18251);
xor U20416 (N_20416,N_16123,N_17172);
xor U20417 (N_20417,N_16110,N_18472);
and U20418 (N_20418,N_16326,N_15896);
and U20419 (N_20419,N_15787,N_16089);
nand U20420 (N_20420,N_17665,N_18580);
xnor U20421 (N_20421,N_17498,N_17083);
nand U20422 (N_20422,N_17683,N_18233);
xor U20423 (N_20423,N_18551,N_16389);
and U20424 (N_20424,N_18252,N_18376);
nor U20425 (N_20425,N_17462,N_16424);
or U20426 (N_20426,N_18264,N_16989);
or U20427 (N_20427,N_18107,N_15810);
xnor U20428 (N_20428,N_17673,N_17135);
and U20429 (N_20429,N_17384,N_18137);
or U20430 (N_20430,N_17485,N_16910);
nand U20431 (N_20431,N_16379,N_16678);
or U20432 (N_20432,N_18666,N_16132);
xnor U20433 (N_20433,N_18503,N_15870);
and U20434 (N_20434,N_18312,N_18433);
nand U20435 (N_20435,N_17262,N_16916);
nand U20436 (N_20436,N_18710,N_16817);
or U20437 (N_20437,N_16877,N_17508);
nand U20438 (N_20438,N_17619,N_16599);
xor U20439 (N_20439,N_18137,N_17231);
and U20440 (N_20440,N_18615,N_16224);
and U20441 (N_20441,N_16462,N_16803);
nand U20442 (N_20442,N_18412,N_16953);
xnor U20443 (N_20443,N_15925,N_16345);
xnor U20444 (N_20444,N_16102,N_16344);
nand U20445 (N_20445,N_16217,N_18337);
xnor U20446 (N_20446,N_16427,N_17760);
nor U20447 (N_20447,N_15958,N_16760);
nor U20448 (N_20448,N_16149,N_17039);
nand U20449 (N_20449,N_18712,N_18387);
or U20450 (N_20450,N_18505,N_16575);
or U20451 (N_20451,N_17273,N_17648);
xnor U20452 (N_20452,N_16522,N_16124);
and U20453 (N_20453,N_18562,N_17992);
and U20454 (N_20454,N_17118,N_18573);
xnor U20455 (N_20455,N_17428,N_18637);
nor U20456 (N_20456,N_18373,N_16959);
xnor U20457 (N_20457,N_16861,N_16591);
nand U20458 (N_20458,N_16067,N_18514);
and U20459 (N_20459,N_15802,N_16414);
nor U20460 (N_20460,N_16048,N_15702);
nand U20461 (N_20461,N_17189,N_18416);
nand U20462 (N_20462,N_18090,N_18046);
and U20463 (N_20463,N_17041,N_18155);
xor U20464 (N_20464,N_18670,N_18699);
nand U20465 (N_20465,N_17855,N_17631);
xor U20466 (N_20466,N_17590,N_16369);
or U20467 (N_20467,N_18349,N_16319);
nor U20468 (N_20468,N_18146,N_16933);
xor U20469 (N_20469,N_17966,N_17863);
or U20470 (N_20470,N_16860,N_18319);
nand U20471 (N_20471,N_17975,N_17364);
nand U20472 (N_20472,N_18112,N_17060);
or U20473 (N_20473,N_18512,N_17910);
or U20474 (N_20474,N_17641,N_16902);
and U20475 (N_20475,N_18728,N_17586);
and U20476 (N_20476,N_16135,N_18380);
nand U20477 (N_20477,N_16308,N_18535);
nand U20478 (N_20478,N_16500,N_16021);
nand U20479 (N_20479,N_17415,N_17290);
and U20480 (N_20480,N_18661,N_16743);
and U20481 (N_20481,N_17485,N_16864);
nand U20482 (N_20482,N_18229,N_18508);
xnor U20483 (N_20483,N_16145,N_17573);
and U20484 (N_20484,N_17866,N_16741);
nor U20485 (N_20485,N_17291,N_15939);
nand U20486 (N_20486,N_17145,N_16655);
xor U20487 (N_20487,N_18110,N_15956);
xor U20488 (N_20488,N_17697,N_17780);
nor U20489 (N_20489,N_17981,N_18636);
and U20490 (N_20490,N_17697,N_16549);
or U20491 (N_20491,N_16955,N_18106);
or U20492 (N_20492,N_17594,N_15850);
xor U20493 (N_20493,N_16355,N_18266);
xnor U20494 (N_20494,N_16267,N_16638);
nor U20495 (N_20495,N_18119,N_18461);
nand U20496 (N_20496,N_18214,N_16428);
nand U20497 (N_20497,N_15709,N_18325);
xor U20498 (N_20498,N_16972,N_16108);
and U20499 (N_20499,N_18260,N_17591);
xnor U20500 (N_20500,N_16007,N_18630);
xnor U20501 (N_20501,N_18185,N_16181);
nand U20502 (N_20502,N_16370,N_18409);
xor U20503 (N_20503,N_18390,N_17295);
nor U20504 (N_20504,N_15642,N_17082);
or U20505 (N_20505,N_18713,N_17329);
nand U20506 (N_20506,N_16754,N_16700);
xor U20507 (N_20507,N_15932,N_18714);
nor U20508 (N_20508,N_18538,N_16168);
nand U20509 (N_20509,N_16705,N_17402);
nor U20510 (N_20510,N_16833,N_18225);
xor U20511 (N_20511,N_17393,N_16059);
xnor U20512 (N_20512,N_18368,N_16177);
nor U20513 (N_20513,N_18372,N_16881);
nor U20514 (N_20514,N_18121,N_17575);
xnor U20515 (N_20515,N_16742,N_18038);
nand U20516 (N_20516,N_16139,N_15722);
or U20517 (N_20517,N_18709,N_17712);
nand U20518 (N_20518,N_17146,N_18467);
or U20519 (N_20519,N_18674,N_15725);
nand U20520 (N_20520,N_17083,N_17589);
xnor U20521 (N_20521,N_16298,N_16353);
xor U20522 (N_20522,N_17014,N_18556);
nand U20523 (N_20523,N_16984,N_16685);
and U20524 (N_20524,N_16668,N_18099);
nand U20525 (N_20525,N_18691,N_18328);
and U20526 (N_20526,N_17085,N_18595);
xor U20527 (N_20527,N_18690,N_18153);
xnor U20528 (N_20528,N_16172,N_16349);
and U20529 (N_20529,N_16484,N_18282);
nand U20530 (N_20530,N_16499,N_17390);
xnor U20531 (N_20531,N_18357,N_17051);
and U20532 (N_20532,N_16314,N_18335);
or U20533 (N_20533,N_17285,N_16415);
xor U20534 (N_20534,N_17295,N_17929);
nand U20535 (N_20535,N_17190,N_16542);
or U20536 (N_20536,N_16192,N_17820);
nand U20537 (N_20537,N_15736,N_18697);
xnor U20538 (N_20538,N_17460,N_16680);
and U20539 (N_20539,N_16417,N_17831);
or U20540 (N_20540,N_16010,N_18094);
and U20541 (N_20541,N_18649,N_16362);
nor U20542 (N_20542,N_15649,N_17724);
or U20543 (N_20543,N_16905,N_15645);
and U20544 (N_20544,N_16812,N_18492);
xor U20545 (N_20545,N_18742,N_17715);
xor U20546 (N_20546,N_16803,N_15950);
and U20547 (N_20547,N_17393,N_17991);
and U20548 (N_20548,N_17246,N_15747);
nor U20549 (N_20549,N_15998,N_17981);
nor U20550 (N_20550,N_16095,N_15846);
nor U20551 (N_20551,N_18153,N_15912);
xor U20552 (N_20552,N_16829,N_16485);
xor U20553 (N_20553,N_17516,N_16181);
or U20554 (N_20554,N_16701,N_16496);
nor U20555 (N_20555,N_16137,N_15875);
and U20556 (N_20556,N_18448,N_17359);
nor U20557 (N_20557,N_18737,N_17153);
or U20558 (N_20558,N_15866,N_15983);
or U20559 (N_20559,N_17997,N_18198);
nand U20560 (N_20560,N_17064,N_16551);
and U20561 (N_20561,N_15750,N_16802);
or U20562 (N_20562,N_16811,N_15685);
xnor U20563 (N_20563,N_16497,N_18513);
xnor U20564 (N_20564,N_17580,N_16968);
or U20565 (N_20565,N_17622,N_15984);
and U20566 (N_20566,N_16937,N_16957);
nand U20567 (N_20567,N_16428,N_18304);
or U20568 (N_20568,N_17494,N_18362);
or U20569 (N_20569,N_16274,N_18614);
xnor U20570 (N_20570,N_16673,N_18637);
or U20571 (N_20571,N_17541,N_18283);
nor U20572 (N_20572,N_17560,N_17383);
and U20573 (N_20573,N_18626,N_16071);
and U20574 (N_20574,N_17042,N_15952);
nand U20575 (N_20575,N_17251,N_18193);
nor U20576 (N_20576,N_16512,N_17217);
nand U20577 (N_20577,N_15793,N_17195);
xor U20578 (N_20578,N_17128,N_16799);
nand U20579 (N_20579,N_18192,N_18098);
and U20580 (N_20580,N_18054,N_18177);
nand U20581 (N_20581,N_18221,N_18512);
xnor U20582 (N_20582,N_18277,N_17429);
or U20583 (N_20583,N_16364,N_18559);
or U20584 (N_20584,N_16504,N_17839);
nand U20585 (N_20585,N_15851,N_16500);
or U20586 (N_20586,N_15926,N_17618);
nand U20587 (N_20587,N_16322,N_18280);
nor U20588 (N_20588,N_17850,N_16471);
nand U20589 (N_20589,N_15995,N_16892);
nor U20590 (N_20590,N_16152,N_17791);
nor U20591 (N_20591,N_16569,N_18620);
and U20592 (N_20592,N_17229,N_16659);
nor U20593 (N_20593,N_16287,N_16245);
nor U20594 (N_20594,N_17037,N_18431);
or U20595 (N_20595,N_18220,N_18740);
nor U20596 (N_20596,N_18639,N_18625);
xnor U20597 (N_20597,N_17056,N_18498);
and U20598 (N_20598,N_16803,N_16351);
nand U20599 (N_20599,N_17554,N_16176);
and U20600 (N_20600,N_16757,N_18087);
and U20601 (N_20601,N_18557,N_18208);
and U20602 (N_20602,N_16853,N_15822);
nor U20603 (N_20603,N_17026,N_18438);
xor U20604 (N_20604,N_16381,N_16735);
nor U20605 (N_20605,N_18109,N_17009);
nand U20606 (N_20606,N_17125,N_17895);
or U20607 (N_20607,N_17993,N_16953);
or U20608 (N_20608,N_18070,N_16746);
xor U20609 (N_20609,N_16742,N_17866);
or U20610 (N_20610,N_18749,N_17159);
nor U20611 (N_20611,N_16468,N_18267);
xnor U20612 (N_20612,N_16651,N_16102);
xor U20613 (N_20613,N_16475,N_16566);
nand U20614 (N_20614,N_16996,N_17324);
and U20615 (N_20615,N_17349,N_17829);
nand U20616 (N_20616,N_16083,N_16495);
nand U20617 (N_20617,N_17489,N_16920);
nand U20618 (N_20618,N_15691,N_16602);
nor U20619 (N_20619,N_17291,N_16471);
or U20620 (N_20620,N_16505,N_16659);
or U20621 (N_20621,N_17841,N_18398);
nor U20622 (N_20622,N_17806,N_16039);
nor U20623 (N_20623,N_18307,N_17634);
or U20624 (N_20624,N_18390,N_17299);
and U20625 (N_20625,N_16831,N_16027);
nand U20626 (N_20626,N_15803,N_18714);
or U20627 (N_20627,N_16699,N_17166);
xor U20628 (N_20628,N_17716,N_15960);
and U20629 (N_20629,N_16608,N_16546);
xnor U20630 (N_20630,N_15760,N_18683);
and U20631 (N_20631,N_17543,N_16909);
or U20632 (N_20632,N_17339,N_16939);
nand U20633 (N_20633,N_17201,N_17159);
xor U20634 (N_20634,N_16486,N_16271);
nor U20635 (N_20635,N_16334,N_18021);
nor U20636 (N_20636,N_17498,N_17622);
nor U20637 (N_20637,N_17301,N_17045);
nand U20638 (N_20638,N_16465,N_18179);
or U20639 (N_20639,N_16195,N_17313);
and U20640 (N_20640,N_15768,N_18222);
nand U20641 (N_20641,N_18735,N_16036);
nor U20642 (N_20642,N_16138,N_17697);
or U20643 (N_20643,N_17426,N_18388);
and U20644 (N_20644,N_16675,N_17162);
xnor U20645 (N_20645,N_16944,N_18616);
nor U20646 (N_20646,N_15881,N_16860);
and U20647 (N_20647,N_16299,N_16453);
nand U20648 (N_20648,N_15662,N_15671);
nand U20649 (N_20649,N_16456,N_17236);
nand U20650 (N_20650,N_18407,N_15862);
xnor U20651 (N_20651,N_18497,N_16536);
xor U20652 (N_20652,N_18036,N_17577);
xnor U20653 (N_20653,N_17034,N_17288);
nand U20654 (N_20654,N_16081,N_17407);
xnor U20655 (N_20655,N_16862,N_17609);
nand U20656 (N_20656,N_17363,N_16665);
nand U20657 (N_20657,N_17472,N_16055);
nor U20658 (N_20658,N_17043,N_16465);
nor U20659 (N_20659,N_18416,N_17605);
nor U20660 (N_20660,N_16408,N_16291);
nand U20661 (N_20661,N_15846,N_18671);
xor U20662 (N_20662,N_18191,N_17839);
nand U20663 (N_20663,N_15660,N_17365);
xnor U20664 (N_20664,N_18710,N_18522);
and U20665 (N_20665,N_18144,N_17411);
nor U20666 (N_20666,N_18704,N_16838);
and U20667 (N_20667,N_15709,N_18126);
nand U20668 (N_20668,N_15808,N_18313);
nand U20669 (N_20669,N_17096,N_17106);
or U20670 (N_20670,N_17270,N_18148);
and U20671 (N_20671,N_16790,N_17978);
xnor U20672 (N_20672,N_16296,N_17397);
nor U20673 (N_20673,N_18432,N_17137);
or U20674 (N_20674,N_17450,N_16166);
xor U20675 (N_20675,N_16368,N_15945);
nand U20676 (N_20676,N_16903,N_16120);
and U20677 (N_20677,N_16530,N_16014);
or U20678 (N_20678,N_18274,N_17294);
nand U20679 (N_20679,N_17856,N_17734);
and U20680 (N_20680,N_15686,N_17644);
xor U20681 (N_20681,N_18344,N_16170);
xnor U20682 (N_20682,N_15730,N_16909);
xor U20683 (N_20683,N_16823,N_17404);
nor U20684 (N_20684,N_16071,N_16302);
or U20685 (N_20685,N_18702,N_16154);
xor U20686 (N_20686,N_16246,N_17078);
nand U20687 (N_20687,N_18729,N_16700);
xnor U20688 (N_20688,N_15955,N_16544);
or U20689 (N_20689,N_16861,N_18464);
xnor U20690 (N_20690,N_15926,N_18629);
xor U20691 (N_20691,N_16708,N_15954);
nor U20692 (N_20692,N_16987,N_17950);
nand U20693 (N_20693,N_18687,N_18335);
xnor U20694 (N_20694,N_15652,N_18128);
and U20695 (N_20695,N_16267,N_16163);
nand U20696 (N_20696,N_17942,N_15763);
nor U20697 (N_20697,N_16237,N_16976);
nor U20698 (N_20698,N_15915,N_16735);
and U20699 (N_20699,N_18427,N_18033);
nor U20700 (N_20700,N_18515,N_15841);
and U20701 (N_20701,N_17990,N_16968);
and U20702 (N_20702,N_17190,N_17554);
and U20703 (N_20703,N_15810,N_18452);
xor U20704 (N_20704,N_17385,N_18331);
nor U20705 (N_20705,N_17401,N_17151);
nand U20706 (N_20706,N_17702,N_17393);
xnor U20707 (N_20707,N_18206,N_17656);
xor U20708 (N_20708,N_16633,N_17014);
xnor U20709 (N_20709,N_16747,N_16297);
nor U20710 (N_20710,N_18176,N_17907);
nor U20711 (N_20711,N_16328,N_18685);
xnor U20712 (N_20712,N_17681,N_15653);
nor U20713 (N_20713,N_16278,N_17778);
nand U20714 (N_20714,N_16341,N_17932);
nor U20715 (N_20715,N_16847,N_16139);
or U20716 (N_20716,N_17866,N_16539);
xor U20717 (N_20717,N_17894,N_17351);
xnor U20718 (N_20718,N_16650,N_18401);
nor U20719 (N_20719,N_17835,N_17471);
or U20720 (N_20720,N_16534,N_16250);
and U20721 (N_20721,N_18155,N_15828);
and U20722 (N_20722,N_16881,N_17676);
or U20723 (N_20723,N_17584,N_17489);
nand U20724 (N_20724,N_18197,N_16962);
and U20725 (N_20725,N_16773,N_16368);
nand U20726 (N_20726,N_15634,N_18144);
or U20727 (N_20727,N_16591,N_17276);
xnor U20728 (N_20728,N_17245,N_17259);
nor U20729 (N_20729,N_18068,N_17736);
or U20730 (N_20730,N_16298,N_17935);
or U20731 (N_20731,N_17506,N_17313);
and U20732 (N_20732,N_16310,N_18529);
nor U20733 (N_20733,N_15987,N_16845);
nor U20734 (N_20734,N_17260,N_17273);
nor U20735 (N_20735,N_18691,N_18212);
xor U20736 (N_20736,N_15833,N_16088);
nor U20737 (N_20737,N_17815,N_17648);
or U20738 (N_20738,N_16146,N_17286);
or U20739 (N_20739,N_15782,N_17275);
and U20740 (N_20740,N_16720,N_16705);
and U20741 (N_20741,N_16337,N_15675);
nand U20742 (N_20742,N_16227,N_16092);
xnor U20743 (N_20743,N_18534,N_17655);
and U20744 (N_20744,N_16264,N_17481);
or U20745 (N_20745,N_18267,N_16646);
xnor U20746 (N_20746,N_17147,N_15852);
nor U20747 (N_20747,N_17446,N_17274);
or U20748 (N_20748,N_17502,N_18275);
and U20749 (N_20749,N_15986,N_16834);
or U20750 (N_20750,N_16895,N_16367);
and U20751 (N_20751,N_16157,N_17014);
and U20752 (N_20752,N_17412,N_17370);
nand U20753 (N_20753,N_16978,N_18649);
or U20754 (N_20754,N_17873,N_15862);
or U20755 (N_20755,N_18517,N_15907);
or U20756 (N_20756,N_17540,N_16453);
and U20757 (N_20757,N_17275,N_17135);
xnor U20758 (N_20758,N_18615,N_16840);
or U20759 (N_20759,N_16906,N_17660);
or U20760 (N_20760,N_18678,N_16403);
nand U20761 (N_20761,N_18009,N_18408);
or U20762 (N_20762,N_18385,N_17495);
nand U20763 (N_20763,N_17849,N_16054);
or U20764 (N_20764,N_16876,N_16124);
and U20765 (N_20765,N_18675,N_16849);
nand U20766 (N_20766,N_18513,N_17654);
xor U20767 (N_20767,N_17391,N_15676);
xor U20768 (N_20768,N_17796,N_17131);
or U20769 (N_20769,N_16189,N_17109);
nand U20770 (N_20770,N_18536,N_18475);
nand U20771 (N_20771,N_16175,N_18000);
xnor U20772 (N_20772,N_16325,N_18366);
xor U20773 (N_20773,N_17351,N_18147);
nor U20774 (N_20774,N_16526,N_18338);
xor U20775 (N_20775,N_17044,N_17082);
xor U20776 (N_20776,N_17077,N_17199);
or U20777 (N_20777,N_18546,N_17266);
nor U20778 (N_20778,N_18195,N_18438);
nor U20779 (N_20779,N_17205,N_16324);
xnor U20780 (N_20780,N_16993,N_16288);
or U20781 (N_20781,N_17042,N_16549);
nor U20782 (N_20782,N_16772,N_16556);
xor U20783 (N_20783,N_16181,N_15629);
nand U20784 (N_20784,N_16389,N_17901);
and U20785 (N_20785,N_18169,N_16980);
nor U20786 (N_20786,N_18325,N_17160);
or U20787 (N_20787,N_15981,N_17510);
xor U20788 (N_20788,N_18020,N_15838);
and U20789 (N_20789,N_18587,N_18398);
xor U20790 (N_20790,N_18128,N_17120);
and U20791 (N_20791,N_16099,N_17379);
and U20792 (N_20792,N_16231,N_15943);
nor U20793 (N_20793,N_18513,N_18682);
and U20794 (N_20794,N_17069,N_18249);
nand U20795 (N_20795,N_17883,N_16263);
xnor U20796 (N_20796,N_18578,N_15794);
and U20797 (N_20797,N_15692,N_16824);
nand U20798 (N_20798,N_16282,N_17042);
xnor U20799 (N_20799,N_16011,N_18011);
xnor U20800 (N_20800,N_16357,N_17787);
and U20801 (N_20801,N_18372,N_15785);
and U20802 (N_20802,N_16644,N_18405);
nor U20803 (N_20803,N_18408,N_17728);
nand U20804 (N_20804,N_18519,N_16034);
xnor U20805 (N_20805,N_16243,N_17892);
xor U20806 (N_20806,N_18341,N_17274);
and U20807 (N_20807,N_16419,N_17735);
and U20808 (N_20808,N_15826,N_17140);
or U20809 (N_20809,N_18355,N_16029);
nand U20810 (N_20810,N_18376,N_15876);
nand U20811 (N_20811,N_15991,N_16947);
and U20812 (N_20812,N_18565,N_17864);
or U20813 (N_20813,N_15730,N_16201);
nor U20814 (N_20814,N_18013,N_16269);
nor U20815 (N_20815,N_16465,N_16187);
or U20816 (N_20816,N_15738,N_18207);
nor U20817 (N_20817,N_17111,N_17524);
xor U20818 (N_20818,N_18002,N_17175);
nand U20819 (N_20819,N_16778,N_17012);
nor U20820 (N_20820,N_17472,N_16963);
xnor U20821 (N_20821,N_18229,N_18368);
xor U20822 (N_20822,N_17626,N_16153);
xor U20823 (N_20823,N_16768,N_15814);
or U20824 (N_20824,N_17405,N_16228);
nor U20825 (N_20825,N_17948,N_16797);
xnor U20826 (N_20826,N_17366,N_17581);
xnor U20827 (N_20827,N_18047,N_17964);
nand U20828 (N_20828,N_16162,N_18615);
nor U20829 (N_20829,N_18687,N_18428);
and U20830 (N_20830,N_18187,N_16015);
and U20831 (N_20831,N_17032,N_16559);
nand U20832 (N_20832,N_17641,N_17256);
and U20833 (N_20833,N_17149,N_18502);
nor U20834 (N_20834,N_18065,N_17467);
xnor U20835 (N_20835,N_16079,N_16874);
xor U20836 (N_20836,N_18700,N_18102);
xnor U20837 (N_20837,N_18594,N_16225);
nor U20838 (N_20838,N_18551,N_17234);
and U20839 (N_20839,N_17857,N_16666);
and U20840 (N_20840,N_18413,N_16735);
nor U20841 (N_20841,N_17153,N_18236);
nor U20842 (N_20842,N_16060,N_18318);
or U20843 (N_20843,N_16817,N_17758);
or U20844 (N_20844,N_16980,N_18241);
nand U20845 (N_20845,N_17916,N_17600);
nor U20846 (N_20846,N_18116,N_18669);
or U20847 (N_20847,N_15798,N_16332);
or U20848 (N_20848,N_15809,N_16580);
xnor U20849 (N_20849,N_17872,N_15963);
nand U20850 (N_20850,N_16279,N_16154);
xnor U20851 (N_20851,N_17457,N_16810);
nor U20852 (N_20852,N_17609,N_17441);
nor U20853 (N_20853,N_17501,N_18509);
nand U20854 (N_20854,N_17247,N_16714);
and U20855 (N_20855,N_16117,N_18575);
or U20856 (N_20856,N_17760,N_15770);
nor U20857 (N_20857,N_17872,N_15915);
nor U20858 (N_20858,N_15754,N_17669);
nand U20859 (N_20859,N_16883,N_17604);
xor U20860 (N_20860,N_18337,N_15809);
nor U20861 (N_20861,N_18533,N_16875);
or U20862 (N_20862,N_18077,N_16023);
nand U20863 (N_20863,N_18291,N_16361);
xor U20864 (N_20864,N_16409,N_18281);
nor U20865 (N_20865,N_16034,N_16758);
or U20866 (N_20866,N_18717,N_18657);
nor U20867 (N_20867,N_15766,N_16034);
or U20868 (N_20868,N_15770,N_17225);
xnor U20869 (N_20869,N_16472,N_18339);
nand U20870 (N_20870,N_15669,N_16778);
or U20871 (N_20871,N_17420,N_17501);
nand U20872 (N_20872,N_17153,N_17189);
nor U20873 (N_20873,N_16673,N_18222);
xnor U20874 (N_20874,N_18675,N_17294);
and U20875 (N_20875,N_17978,N_17187);
xor U20876 (N_20876,N_18529,N_17027);
xor U20877 (N_20877,N_17216,N_16031);
and U20878 (N_20878,N_17551,N_18041);
nand U20879 (N_20879,N_17184,N_17711);
and U20880 (N_20880,N_17026,N_16164);
nor U20881 (N_20881,N_18037,N_18266);
nor U20882 (N_20882,N_16738,N_16631);
and U20883 (N_20883,N_16443,N_16552);
xnor U20884 (N_20884,N_17432,N_16132);
xnor U20885 (N_20885,N_17294,N_17292);
nand U20886 (N_20886,N_17483,N_18299);
and U20887 (N_20887,N_16534,N_18091);
and U20888 (N_20888,N_17635,N_16869);
xor U20889 (N_20889,N_15681,N_16455);
or U20890 (N_20890,N_17419,N_16120);
nand U20891 (N_20891,N_17909,N_18476);
nor U20892 (N_20892,N_15799,N_15664);
and U20893 (N_20893,N_17725,N_18211);
xnor U20894 (N_20894,N_17135,N_17103);
or U20895 (N_20895,N_17040,N_18282);
xor U20896 (N_20896,N_16802,N_16799);
xor U20897 (N_20897,N_16700,N_16846);
xor U20898 (N_20898,N_18328,N_17811);
xnor U20899 (N_20899,N_16009,N_16486);
and U20900 (N_20900,N_16660,N_18381);
nor U20901 (N_20901,N_16737,N_16906);
nor U20902 (N_20902,N_17577,N_16537);
and U20903 (N_20903,N_16291,N_15805);
or U20904 (N_20904,N_17134,N_18717);
nor U20905 (N_20905,N_15982,N_15768);
xor U20906 (N_20906,N_15770,N_16545);
or U20907 (N_20907,N_16327,N_15939);
nor U20908 (N_20908,N_18417,N_16738);
xnor U20909 (N_20909,N_16230,N_16277);
nor U20910 (N_20910,N_17959,N_15628);
nand U20911 (N_20911,N_17980,N_18148);
or U20912 (N_20912,N_18652,N_16616);
and U20913 (N_20913,N_15921,N_17989);
xnor U20914 (N_20914,N_17901,N_15662);
nand U20915 (N_20915,N_17470,N_17252);
nand U20916 (N_20916,N_15899,N_18130);
nand U20917 (N_20917,N_15633,N_18103);
xnor U20918 (N_20918,N_16236,N_18419);
xor U20919 (N_20919,N_15992,N_16843);
xor U20920 (N_20920,N_17101,N_18287);
and U20921 (N_20921,N_18422,N_16370);
nor U20922 (N_20922,N_16506,N_15896);
and U20923 (N_20923,N_16024,N_15717);
nor U20924 (N_20924,N_15822,N_16459);
and U20925 (N_20925,N_17554,N_18712);
or U20926 (N_20926,N_18571,N_18154);
nand U20927 (N_20927,N_17051,N_17296);
or U20928 (N_20928,N_17479,N_18102);
xnor U20929 (N_20929,N_16070,N_17884);
xnor U20930 (N_20930,N_16381,N_16501);
or U20931 (N_20931,N_16798,N_17768);
nor U20932 (N_20932,N_18021,N_17284);
nand U20933 (N_20933,N_17991,N_17377);
and U20934 (N_20934,N_17448,N_18216);
xor U20935 (N_20935,N_16551,N_15840);
and U20936 (N_20936,N_18409,N_16386);
xnor U20937 (N_20937,N_16369,N_16313);
nor U20938 (N_20938,N_17266,N_15827);
nand U20939 (N_20939,N_16459,N_16641);
or U20940 (N_20940,N_18185,N_16941);
xor U20941 (N_20941,N_15648,N_16260);
nor U20942 (N_20942,N_17247,N_17003);
and U20943 (N_20943,N_17650,N_17656);
or U20944 (N_20944,N_17313,N_17254);
nor U20945 (N_20945,N_17616,N_17565);
nor U20946 (N_20946,N_15918,N_17207);
nand U20947 (N_20947,N_17542,N_16936);
xnor U20948 (N_20948,N_17313,N_16574);
and U20949 (N_20949,N_16119,N_18572);
or U20950 (N_20950,N_16899,N_18612);
xnor U20951 (N_20951,N_18067,N_15769);
and U20952 (N_20952,N_17365,N_17987);
or U20953 (N_20953,N_16783,N_16240);
nand U20954 (N_20954,N_18366,N_17044);
xnor U20955 (N_20955,N_18194,N_18340);
xnor U20956 (N_20956,N_17417,N_16965);
or U20957 (N_20957,N_17327,N_16394);
xnor U20958 (N_20958,N_18348,N_17417);
nor U20959 (N_20959,N_18183,N_16561);
nand U20960 (N_20960,N_16056,N_17212);
or U20961 (N_20961,N_18329,N_18474);
nand U20962 (N_20962,N_15863,N_18695);
nor U20963 (N_20963,N_16799,N_16807);
nor U20964 (N_20964,N_17895,N_18169);
and U20965 (N_20965,N_17890,N_18651);
or U20966 (N_20966,N_18324,N_16345);
and U20967 (N_20967,N_17044,N_17214);
or U20968 (N_20968,N_17300,N_18528);
xor U20969 (N_20969,N_16128,N_17147);
xnor U20970 (N_20970,N_16890,N_16852);
xor U20971 (N_20971,N_17029,N_16603);
nor U20972 (N_20972,N_18381,N_17482);
xor U20973 (N_20973,N_17699,N_17732);
or U20974 (N_20974,N_16061,N_17772);
and U20975 (N_20975,N_16655,N_17858);
and U20976 (N_20976,N_18082,N_18710);
nor U20977 (N_20977,N_18647,N_17966);
or U20978 (N_20978,N_18249,N_18088);
and U20979 (N_20979,N_16461,N_16604);
xor U20980 (N_20980,N_18168,N_15992);
and U20981 (N_20981,N_18254,N_17777);
or U20982 (N_20982,N_17269,N_15632);
xnor U20983 (N_20983,N_18342,N_17558);
nand U20984 (N_20984,N_18294,N_15836);
xor U20985 (N_20985,N_18440,N_18618);
or U20986 (N_20986,N_17414,N_18011);
and U20987 (N_20987,N_17452,N_18397);
nand U20988 (N_20988,N_17152,N_17826);
xnor U20989 (N_20989,N_16179,N_18737);
or U20990 (N_20990,N_17577,N_15880);
or U20991 (N_20991,N_17104,N_18708);
or U20992 (N_20992,N_16449,N_17011);
xnor U20993 (N_20993,N_16467,N_18363);
xnor U20994 (N_20994,N_16964,N_15824);
xnor U20995 (N_20995,N_16332,N_15857);
and U20996 (N_20996,N_16667,N_18666);
or U20997 (N_20997,N_18102,N_16284);
nand U20998 (N_20998,N_16187,N_18393);
nor U20999 (N_20999,N_18642,N_17117);
nand U21000 (N_21000,N_17262,N_16541);
and U21001 (N_21001,N_16550,N_18415);
and U21002 (N_21002,N_17838,N_15637);
nand U21003 (N_21003,N_16675,N_16570);
nand U21004 (N_21004,N_16479,N_16207);
nand U21005 (N_21005,N_16554,N_17452);
nor U21006 (N_21006,N_15814,N_17340);
nand U21007 (N_21007,N_17733,N_16160);
nand U21008 (N_21008,N_18434,N_17553);
or U21009 (N_21009,N_17454,N_17933);
and U21010 (N_21010,N_17619,N_17335);
nor U21011 (N_21011,N_17599,N_16959);
nand U21012 (N_21012,N_15788,N_18141);
nand U21013 (N_21013,N_17268,N_17528);
or U21014 (N_21014,N_18564,N_17893);
nand U21015 (N_21015,N_16971,N_15771);
and U21016 (N_21016,N_15838,N_17478);
or U21017 (N_21017,N_17471,N_18175);
nor U21018 (N_21018,N_15815,N_17112);
xnor U21019 (N_21019,N_17638,N_16691);
nor U21020 (N_21020,N_18610,N_17462);
nor U21021 (N_21021,N_16810,N_15925);
or U21022 (N_21022,N_16194,N_17861);
and U21023 (N_21023,N_16385,N_17042);
nand U21024 (N_21024,N_17278,N_18133);
xnor U21025 (N_21025,N_18650,N_16764);
and U21026 (N_21026,N_16203,N_17129);
xnor U21027 (N_21027,N_15754,N_15900);
and U21028 (N_21028,N_17855,N_16781);
nand U21029 (N_21029,N_16784,N_17434);
nor U21030 (N_21030,N_16453,N_16918);
nor U21031 (N_21031,N_18485,N_16805);
xor U21032 (N_21032,N_17082,N_16599);
and U21033 (N_21033,N_18556,N_17492);
or U21034 (N_21034,N_17987,N_18358);
nand U21035 (N_21035,N_18745,N_17427);
or U21036 (N_21036,N_17675,N_16091);
xnor U21037 (N_21037,N_15924,N_17729);
nor U21038 (N_21038,N_17274,N_18073);
nor U21039 (N_21039,N_17919,N_18632);
xor U21040 (N_21040,N_15971,N_18020);
nor U21041 (N_21041,N_18387,N_18699);
nor U21042 (N_21042,N_16950,N_17510);
or U21043 (N_21043,N_17202,N_17654);
nand U21044 (N_21044,N_15707,N_18089);
nand U21045 (N_21045,N_17964,N_16214);
or U21046 (N_21046,N_18613,N_16550);
nand U21047 (N_21047,N_17387,N_15715);
or U21048 (N_21048,N_15814,N_15675);
nor U21049 (N_21049,N_18180,N_18490);
xnor U21050 (N_21050,N_16915,N_17687);
xor U21051 (N_21051,N_16263,N_18533);
xor U21052 (N_21052,N_16642,N_16521);
nor U21053 (N_21053,N_18189,N_17602);
or U21054 (N_21054,N_17304,N_16829);
xor U21055 (N_21055,N_16342,N_18038);
or U21056 (N_21056,N_18331,N_16669);
or U21057 (N_21057,N_17959,N_15855);
nor U21058 (N_21058,N_16410,N_18018);
nor U21059 (N_21059,N_16152,N_18342);
or U21060 (N_21060,N_15896,N_18276);
nand U21061 (N_21061,N_17357,N_18404);
nor U21062 (N_21062,N_16544,N_16676);
or U21063 (N_21063,N_15852,N_18322);
nor U21064 (N_21064,N_17194,N_18033);
xnor U21065 (N_21065,N_17507,N_16888);
nand U21066 (N_21066,N_16296,N_17948);
nand U21067 (N_21067,N_16389,N_17919);
and U21068 (N_21068,N_18580,N_17284);
xnor U21069 (N_21069,N_16171,N_15904);
nand U21070 (N_21070,N_17538,N_15722);
and U21071 (N_21071,N_15678,N_17981);
xnor U21072 (N_21072,N_17336,N_16336);
nand U21073 (N_21073,N_15988,N_17259);
or U21074 (N_21074,N_17916,N_16256);
xor U21075 (N_21075,N_17804,N_16597);
or U21076 (N_21076,N_16336,N_18301);
and U21077 (N_21077,N_15927,N_17203);
nor U21078 (N_21078,N_18498,N_17289);
and U21079 (N_21079,N_17738,N_18424);
or U21080 (N_21080,N_16130,N_17860);
nand U21081 (N_21081,N_16197,N_17371);
or U21082 (N_21082,N_16205,N_16649);
xnor U21083 (N_21083,N_18642,N_17716);
nand U21084 (N_21084,N_16755,N_16866);
xor U21085 (N_21085,N_18646,N_18606);
nand U21086 (N_21086,N_16710,N_15912);
nand U21087 (N_21087,N_17070,N_18139);
nand U21088 (N_21088,N_18183,N_15847);
xor U21089 (N_21089,N_17298,N_18310);
and U21090 (N_21090,N_16560,N_17149);
or U21091 (N_21091,N_16143,N_17322);
or U21092 (N_21092,N_15942,N_18293);
nor U21093 (N_21093,N_15880,N_15911);
or U21094 (N_21094,N_15959,N_17818);
or U21095 (N_21095,N_15813,N_17959);
nand U21096 (N_21096,N_16472,N_16626);
xnor U21097 (N_21097,N_17641,N_17303);
nand U21098 (N_21098,N_16748,N_17189);
nand U21099 (N_21099,N_16397,N_17584);
and U21100 (N_21100,N_16284,N_18127);
and U21101 (N_21101,N_16356,N_16435);
xor U21102 (N_21102,N_16629,N_18066);
nand U21103 (N_21103,N_16970,N_17791);
xor U21104 (N_21104,N_16653,N_16860);
and U21105 (N_21105,N_18597,N_15662);
nor U21106 (N_21106,N_17112,N_18399);
and U21107 (N_21107,N_16719,N_17344);
nand U21108 (N_21108,N_15852,N_17418);
nor U21109 (N_21109,N_17098,N_16079);
and U21110 (N_21110,N_16119,N_18067);
nand U21111 (N_21111,N_17187,N_18484);
nor U21112 (N_21112,N_16957,N_16996);
xor U21113 (N_21113,N_17847,N_18242);
or U21114 (N_21114,N_16920,N_17220);
or U21115 (N_21115,N_18087,N_16688);
and U21116 (N_21116,N_16674,N_16375);
nor U21117 (N_21117,N_18104,N_17137);
xor U21118 (N_21118,N_16025,N_18134);
xor U21119 (N_21119,N_16883,N_18612);
or U21120 (N_21120,N_15857,N_18459);
nor U21121 (N_21121,N_17023,N_18739);
xor U21122 (N_21122,N_18536,N_15692);
or U21123 (N_21123,N_18336,N_18098);
nor U21124 (N_21124,N_18165,N_18724);
nand U21125 (N_21125,N_17580,N_17422);
nand U21126 (N_21126,N_16017,N_16424);
nand U21127 (N_21127,N_18319,N_18551);
nor U21128 (N_21128,N_17341,N_17953);
or U21129 (N_21129,N_18120,N_15830);
or U21130 (N_21130,N_17392,N_17143);
or U21131 (N_21131,N_18066,N_17146);
xor U21132 (N_21132,N_18564,N_17402);
nand U21133 (N_21133,N_17498,N_18518);
nor U21134 (N_21134,N_18389,N_17926);
or U21135 (N_21135,N_16872,N_16896);
and U21136 (N_21136,N_17556,N_17932);
nand U21137 (N_21137,N_17528,N_16538);
nand U21138 (N_21138,N_18509,N_17814);
nor U21139 (N_21139,N_17971,N_17948);
or U21140 (N_21140,N_16058,N_16926);
and U21141 (N_21141,N_16029,N_17093);
nand U21142 (N_21142,N_16760,N_17165);
nand U21143 (N_21143,N_16952,N_17004);
and U21144 (N_21144,N_18603,N_18697);
and U21145 (N_21145,N_15852,N_15654);
nor U21146 (N_21146,N_18088,N_18182);
nor U21147 (N_21147,N_18321,N_17009);
or U21148 (N_21148,N_16309,N_17198);
xnor U21149 (N_21149,N_18004,N_16779);
nor U21150 (N_21150,N_16086,N_17810);
or U21151 (N_21151,N_16884,N_16336);
nand U21152 (N_21152,N_17593,N_16919);
xor U21153 (N_21153,N_16695,N_18437);
and U21154 (N_21154,N_16638,N_15685);
nand U21155 (N_21155,N_18305,N_15705);
xnor U21156 (N_21156,N_16424,N_18322);
nand U21157 (N_21157,N_17856,N_16785);
nor U21158 (N_21158,N_17627,N_17986);
nor U21159 (N_21159,N_16867,N_16879);
nor U21160 (N_21160,N_16325,N_17988);
or U21161 (N_21161,N_16706,N_17409);
xnor U21162 (N_21162,N_15862,N_18509);
and U21163 (N_21163,N_16082,N_15671);
and U21164 (N_21164,N_18583,N_16023);
and U21165 (N_21165,N_16175,N_16387);
and U21166 (N_21166,N_17474,N_16071);
xnor U21167 (N_21167,N_17885,N_18676);
nor U21168 (N_21168,N_16327,N_17112);
nor U21169 (N_21169,N_18027,N_16253);
and U21170 (N_21170,N_17574,N_15756);
and U21171 (N_21171,N_17892,N_16089);
nor U21172 (N_21172,N_18000,N_16453);
or U21173 (N_21173,N_17893,N_18204);
and U21174 (N_21174,N_17087,N_17478);
xnor U21175 (N_21175,N_17195,N_15875);
and U21176 (N_21176,N_17955,N_16828);
xor U21177 (N_21177,N_18539,N_17092);
and U21178 (N_21178,N_17750,N_16069);
nor U21179 (N_21179,N_16358,N_15755);
xnor U21180 (N_21180,N_17916,N_16473);
and U21181 (N_21181,N_16475,N_16570);
nand U21182 (N_21182,N_16265,N_16874);
nand U21183 (N_21183,N_17829,N_16782);
nand U21184 (N_21184,N_16016,N_18087);
xnor U21185 (N_21185,N_16937,N_16789);
xor U21186 (N_21186,N_15848,N_18076);
or U21187 (N_21187,N_16458,N_18616);
nand U21188 (N_21188,N_16947,N_17672);
nor U21189 (N_21189,N_17354,N_15669);
and U21190 (N_21190,N_16345,N_17714);
and U21191 (N_21191,N_18409,N_17235);
xnor U21192 (N_21192,N_17208,N_16820);
nor U21193 (N_21193,N_16722,N_16653);
xor U21194 (N_21194,N_16295,N_16383);
nor U21195 (N_21195,N_17971,N_16916);
or U21196 (N_21196,N_18409,N_16238);
nand U21197 (N_21197,N_15826,N_15825);
and U21198 (N_21198,N_16515,N_16220);
xnor U21199 (N_21199,N_16335,N_17011);
nor U21200 (N_21200,N_18362,N_15796);
and U21201 (N_21201,N_17334,N_17397);
and U21202 (N_21202,N_16155,N_17759);
and U21203 (N_21203,N_17617,N_18512);
or U21204 (N_21204,N_16769,N_16121);
nor U21205 (N_21205,N_17901,N_18000);
or U21206 (N_21206,N_18538,N_16040);
nand U21207 (N_21207,N_17940,N_16840);
or U21208 (N_21208,N_16778,N_17162);
nand U21209 (N_21209,N_18230,N_18516);
nor U21210 (N_21210,N_18609,N_18226);
or U21211 (N_21211,N_18658,N_18724);
nor U21212 (N_21212,N_16108,N_18100);
nand U21213 (N_21213,N_15957,N_16103);
nand U21214 (N_21214,N_16370,N_17173);
and U21215 (N_21215,N_18077,N_17234);
and U21216 (N_21216,N_17558,N_17351);
nand U21217 (N_21217,N_18621,N_17432);
nor U21218 (N_21218,N_18468,N_17123);
and U21219 (N_21219,N_18297,N_16707);
and U21220 (N_21220,N_18350,N_18103);
xor U21221 (N_21221,N_17810,N_18354);
and U21222 (N_21222,N_16379,N_17908);
nor U21223 (N_21223,N_16973,N_17349);
or U21224 (N_21224,N_16674,N_17501);
xnor U21225 (N_21225,N_17937,N_16519);
and U21226 (N_21226,N_17765,N_16503);
nand U21227 (N_21227,N_18373,N_18037);
xor U21228 (N_21228,N_16003,N_17562);
xnor U21229 (N_21229,N_18327,N_16770);
nor U21230 (N_21230,N_15729,N_17919);
and U21231 (N_21231,N_17542,N_15865);
and U21232 (N_21232,N_16583,N_15773);
and U21233 (N_21233,N_16973,N_15705);
or U21234 (N_21234,N_16538,N_18010);
xor U21235 (N_21235,N_15977,N_18325);
xor U21236 (N_21236,N_17136,N_17003);
nor U21237 (N_21237,N_17211,N_16877);
nand U21238 (N_21238,N_16709,N_17744);
nand U21239 (N_21239,N_18194,N_16757);
and U21240 (N_21240,N_16043,N_18461);
nand U21241 (N_21241,N_18187,N_18253);
and U21242 (N_21242,N_15885,N_17064);
nor U21243 (N_21243,N_16649,N_18057);
nor U21244 (N_21244,N_15936,N_16074);
nor U21245 (N_21245,N_16753,N_17014);
nand U21246 (N_21246,N_18065,N_16766);
nor U21247 (N_21247,N_17667,N_17930);
and U21248 (N_21248,N_18642,N_17112);
nor U21249 (N_21249,N_18414,N_15664);
and U21250 (N_21250,N_15998,N_16337);
nor U21251 (N_21251,N_16813,N_16335);
or U21252 (N_21252,N_15746,N_18014);
xnor U21253 (N_21253,N_18674,N_16812);
and U21254 (N_21254,N_17874,N_18663);
nor U21255 (N_21255,N_18174,N_15719);
nor U21256 (N_21256,N_18291,N_16106);
nand U21257 (N_21257,N_16364,N_18269);
nand U21258 (N_21258,N_17252,N_16866);
and U21259 (N_21259,N_15960,N_17818);
nand U21260 (N_21260,N_18363,N_16969);
nand U21261 (N_21261,N_18084,N_15897);
and U21262 (N_21262,N_17682,N_18521);
nor U21263 (N_21263,N_16307,N_17323);
xnor U21264 (N_21264,N_16793,N_17799);
and U21265 (N_21265,N_16185,N_17060);
and U21266 (N_21266,N_18696,N_16816);
and U21267 (N_21267,N_15869,N_15876);
and U21268 (N_21268,N_15874,N_17499);
nor U21269 (N_21269,N_15795,N_17642);
nor U21270 (N_21270,N_16850,N_17242);
or U21271 (N_21271,N_16758,N_15870);
xor U21272 (N_21272,N_16896,N_17318);
or U21273 (N_21273,N_16637,N_17675);
nand U21274 (N_21274,N_16858,N_17933);
and U21275 (N_21275,N_17154,N_15906);
nand U21276 (N_21276,N_18557,N_17450);
nand U21277 (N_21277,N_16854,N_18586);
or U21278 (N_21278,N_16763,N_16224);
and U21279 (N_21279,N_18168,N_16949);
nand U21280 (N_21280,N_16776,N_18680);
and U21281 (N_21281,N_15746,N_15713);
xnor U21282 (N_21282,N_16666,N_15818);
xnor U21283 (N_21283,N_17833,N_16599);
nand U21284 (N_21284,N_18330,N_17382);
xor U21285 (N_21285,N_17231,N_18705);
or U21286 (N_21286,N_18426,N_17853);
xor U21287 (N_21287,N_16840,N_18220);
xnor U21288 (N_21288,N_16569,N_15697);
and U21289 (N_21289,N_16105,N_18497);
and U21290 (N_21290,N_18175,N_18314);
xnor U21291 (N_21291,N_17770,N_15742);
xnor U21292 (N_21292,N_17165,N_16577);
and U21293 (N_21293,N_18583,N_15775);
or U21294 (N_21294,N_16347,N_16005);
nand U21295 (N_21295,N_18193,N_16147);
xnor U21296 (N_21296,N_17010,N_18570);
or U21297 (N_21297,N_18476,N_16966);
nand U21298 (N_21298,N_17322,N_17304);
xnor U21299 (N_21299,N_16506,N_16067);
or U21300 (N_21300,N_18595,N_16436);
nor U21301 (N_21301,N_16332,N_17415);
nor U21302 (N_21302,N_17940,N_15729);
nand U21303 (N_21303,N_16919,N_16141);
or U21304 (N_21304,N_16498,N_15650);
and U21305 (N_21305,N_18051,N_18100);
nor U21306 (N_21306,N_17022,N_18176);
or U21307 (N_21307,N_18422,N_17233);
xnor U21308 (N_21308,N_16735,N_17098);
and U21309 (N_21309,N_16690,N_17267);
xor U21310 (N_21310,N_17906,N_18306);
or U21311 (N_21311,N_16337,N_16250);
and U21312 (N_21312,N_15863,N_18047);
and U21313 (N_21313,N_17715,N_18569);
or U21314 (N_21314,N_16602,N_17309);
xor U21315 (N_21315,N_18495,N_17665);
nand U21316 (N_21316,N_17970,N_15829);
and U21317 (N_21317,N_17983,N_16310);
nand U21318 (N_21318,N_17606,N_16752);
nor U21319 (N_21319,N_15864,N_17944);
nand U21320 (N_21320,N_17263,N_17500);
or U21321 (N_21321,N_18171,N_15685);
and U21322 (N_21322,N_17500,N_17444);
nand U21323 (N_21323,N_18098,N_16312);
xnor U21324 (N_21324,N_18021,N_15796);
nand U21325 (N_21325,N_18683,N_18290);
nand U21326 (N_21326,N_16973,N_16739);
or U21327 (N_21327,N_17652,N_15907);
or U21328 (N_21328,N_17773,N_16043);
nor U21329 (N_21329,N_18288,N_16293);
xor U21330 (N_21330,N_17354,N_18585);
nand U21331 (N_21331,N_17072,N_16311);
or U21332 (N_21332,N_17672,N_17041);
or U21333 (N_21333,N_17898,N_16346);
or U21334 (N_21334,N_17117,N_15788);
nor U21335 (N_21335,N_15897,N_17807);
nor U21336 (N_21336,N_17578,N_17985);
nand U21337 (N_21337,N_17449,N_16008);
and U21338 (N_21338,N_18066,N_18085);
or U21339 (N_21339,N_15925,N_16183);
or U21340 (N_21340,N_17690,N_18028);
nor U21341 (N_21341,N_16599,N_18501);
or U21342 (N_21342,N_18138,N_16823);
xor U21343 (N_21343,N_15719,N_18383);
or U21344 (N_21344,N_18007,N_17267);
nand U21345 (N_21345,N_15817,N_17248);
xnor U21346 (N_21346,N_15765,N_18029);
nor U21347 (N_21347,N_18222,N_15823);
nand U21348 (N_21348,N_18493,N_17799);
xnor U21349 (N_21349,N_17895,N_16166);
xnor U21350 (N_21350,N_15733,N_16991);
and U21351 (N_21351,N_17354,N_16111);
xor U21352 (N_21352,N_16602,N_16562);
nor U21353 (N_21353,N_18560,N_16290);
xor U21354 (N_21354,N_16321,N_16772);
and U21355 (N_21355,N_17986,N_17577);
or U21356 (N_21356,N_17012,N_17398);
xor U21357 (N_21357,N_15842,N_17924);
nand U21358 (N_21358,N_16390,N_17409);
and U21359 (N_21359,N_17107,N_15725);
nor U21360 (N_21360,N_17854,N_18094);
nor U21361 (N_21361,N_15869,N_17460);
and U21362 (N_21362,N_17956,N_16205);
and U21363 (N_21363,N_16281,N_18660);
xor U21364 (N_21364,N_17056,N_17547);
or U21365 (N_21365,N_18331,N_18358);
xor U21366 (N_21366,N_18681,N_18712);
or U21367 (N_21367,N_17595,N_18470);
nor U21368 (N_21368,N_16890,N_16506);
xor U21369 (N_21369,N_15726,N_18488);
xnor U21370 (N_21370,N_15721,N_15993);
nand U21371 (N_21371,N_16242,N_17295);
nand U21372 (N_21372,N_18328,N_17427);
nand U21373 (N_21373,N_16182,N_16363);
xnor U21374 (N_21374,N_17364,N_18248);
and U21375 (N_21375,N_18048,N_16480);
or U21376 (N_21376,N_18039,N_17554);
or U21377 (N_21377,N_17324,N_18647);
and U21378 (N_21378,N_15794,N_18394);
and U21379 (N_21379,N_18289,N_17102);
xor U21380 (N_21380,N_16454,N_17434);
xor U21381 (N_21381,N_17075,N_16650);
and U21382 (N_21382,N_17420,N_16488);
nand U21383 (N_21383,N_17224,N_16344);
xnor U21384 (N_21384,N_15690,N_18012);
nor U21385 (N_21385,N_15886,N_16687);
xnor U21386 (N_21386,N_15661,N_15864);
and U21387 (N_21387,N_18647,N_16836);
nor U21388 (N_21388,N_18707,N_15841);
and U21389 (N_21389,N_17290,N_18692);
or U21390 (N_21390,N_16540,N_16389);
xnor U21391 (N_21391,N_16495,N_16934);
nor U21392 (N_21392,N_18641,N_16258);
nand U21393 (N_21393,N_17478,N_18125);
and U21394 (N_21394,N_17003,N_16900);
or U21395 (N_21395,N_15739,N_15846);
xnor U21396 (N_21396,N_16802,N_18043);
nand U21397 (N_21397,N_16300,N_17805);
or U21398 (N_21398,N_15804,N_16206);
nand U21399 (N_21399,N_17976,N_18019);
xnor U21400 (N_21400,N_17574,N_18521);
or U21401 (N_21401,N_17410,N_15639);
nor U21402 (N_21402,N_18606,N_18686);
nor U21403 (N_21403,N_17726,N_15821);
or U21404 (N_21404,N_16624,N_16117);
nor U21405 (N_21405,N_16682,N_17770);
nand U21406 (N_21406,N_17530,N_16889);
nor U21407 (N_21407,N_18217,N_18694);
and U21408 (N_21408,N_18001,N_16476);
or U21409 (N_21409,N_18737,N_16536);
or U21410 (N_21410,N_17874,N_15915);
or U21411 (N_21411,N_17542,N_16897);
and U21412 (N_21412,N_16119,N_18440);
xnor U21413 (N_21413,N_16659,N_17984);
or U21414 (N_21414,N_17782,N_15767);
or U21415 (N_21415,N_17763,N_15982);
nand U21416 (N_21416,N_18557,N_17687);
nand U21417 (N_21417,N_17675,N_17920);
or U21418 (N_21418,N_16209,N_16275);
and U21419 (N_21419,N_18467,N_16752);
xnor U21420 (N_21420,N_15778,N_17425);
and U21421 (N_21421,N_15909,N_17666);
nor U21422 (N_21422,N_17119,N_17098);
xnor U21423 (N_21423,N_18113,N_15743);
nor U21424 (N_21424,N_15758,N_18649);
nor U21425 (N_21425,N_15633,N_18641);
and U21426 (N_21426,N_18040,N_16440);
and U21427 (N_21427,N_16827,N_17554);
or U21428 (N_21428,N_15759,N_16946);
xor U21429 (N_21429,N_16813,N_18236);
nand U21430 (N_21430,N_18017,N_16197);
nor U21431 (N_21431,N_16749,N_15834);
nor U21432 (N_21432,N_18276,N_16121);
nor U21433 (N_21433,N_18571,N_16517);
nand U21434 (N_21434,N_16284,N_18244);
nor U21435 (N_21435,N_17701,N_17640);
nand U21436 (N_21436,N_17241,N_15851);
and U21437 (N_21437,N_18358,N_16643);
xor U21438 (N_21438,N_17197,N_16234);
or U21439 (N_21439,N_17873,N_17204);
or U21440 (N_21440,N_16930,N_17181);
nand U21441 (N_21441,N_18117,N_16658);
nor U21442 (N_21442,N_15652,N_17649);
nor U21443 (N_21443,N_17673,N_16881);
nand U21444 (N_21444,N_16307,N_15761);
and U21445 (N_21445,N_16249,N_16687);
or U21446 (N_21446,N_18693,N_17727);
xor U21447 (N_21447,N_17263,N_15811);
xor U21448 (N_21448,N_15684,N_16822);
nand U21449 (N_21449,N_16501,N_18123);
and U21450 (N_21450,N_17576,N_15714);
nand U21451 (N_21451,N_18708,N_17647);
xnor U21452 (N_21452,N_16284,N_18661);
or U21453 (N_21453,N_16640,N_16115);
or U21454 (N_21454,N_17254,N_16297);
nor U21455 (N_21455,N_18125,N_17577);
nor U21456 (N_21456,N_18294,N_16757);
nand U21457 (N_21457,N_17828,N_15854);
or U21458 (N_21458,N_16186,N_16336);
xnor U21459 (N_21459,N_17469,N_16027);
and U21460 (N_21460,N_17096,N_16044);
and U21461 (N_21461,N_18217,N_17164);
xnor U21462 (N_21462,N_15951,N_18555);
and U21463 (N_21463,N_17074,N_16550);
xor U21464 (N_21464,N_18466,N_17845);
and U21465 (N_21465,N_16395,N_15665);
nand U21466 (N_21466,N_15637,N_16922);
nor U21467 (N_21467,N_16782,N_16136);
nand U21468 (N_21468,N_16776,N_16843);
nand U21469 (N_21469,N_18235,N_16780);
xor U21470 (N_21470,N_18318,N_16943);
or U21471 (N_21471,N_16370,N_18632);
nand U21472 (N_21472,N_18339,N_18446);
xor U21473 (N_21473,N_17494,N_17101);
xnor U21474 (N_21474,N_16546,N_17318);
nand U21475 (N_21475,N_18553,N_17197);
nor U21476 (N_21476,N_16773,N_18126);
nor U21477 (N_21477,N_18488,N_18084);
nor U21478 (N_21478,N_17869,N_16311);
nand U21479 (N_21479,N_18490,N_18014);
nand U21480 (N_21480,N_17852,N_18461);
xnor U21481 (N_21481,N_17794,N_17155);
xnor U21482 (N_21482,N_15631,N_18598);
and U21483 (N_21483,N_17180,N_18011);
or U21484 (N_21484,N_17334,N_17497);
nor U21485 (N_21485,N_15746,N_16257);
or U21486 (N_21486,N_16835,N_16451);
xnor U21487 (N_21487,N_18415,N_17480);
xnor U21488 (N_21488,N_15922,N_17699);
nor U21489 (N_21489,N_16926,N_18032);
and U21490 (N_21490,N_16777,N_17216);
and U21491 (N_21491,N_16519,N_16068);
nand U21492 (N_21492,N_18707,N_17397);
and U21493 (N_21493,N_17631,N_16231);
nor U21494 (N_21494,N_16610,N_18075);
nor U21495 (N_21495,N_17347,N_16251);
xor U21496 (N_21496,N_17025,N_16760);
xor U21497 (N_21497,N_16683,N_15762);
nor U21498 (N_21498,N_16066,N_18225);
or U21499 (N_21499,N_16898,N_17309);
and U21500 (N_21500,N_16227,N_16253);
or U21501 (N_21501,N_18621,N_18525);
and U21502 (N_21502,N_15971,N_15798);
and U21503 (N_21503,N_16627,N_16967);
nand U21504 (N_21504,N_18578,N_16795);
nor U21505 (N_21505,N_16063,N_18529);
nand U21506 (N_21506,N_16539,N_15718);
xnor U21507 (N_21507,N_18187,N_17945);
nand U21508 (N_21508,N_16201,N_17085);
nor U21509 (N_21509,N_16981,N_16422);
and U21510 (N_21510,N_18637,N_18020);
and U21511 (N_21511,N_18170,N_16627);
xor U21512 (N_21512,N_17637,N_16840);
xor U21513 (N_21513,N_17113,N_17220);
nand U21514 (N_21514,N_18243,N_16296);
nor U21515 (N_21515,N_17991,N_17586);
nand U21516 (N_21516,N_16213,N_17839);
nor U21517 (N_21517,N_17523,N_17119);
and U21518 (N_21518,N_16720,N_18532);
nor U21519 (N_21519,N_17214,N_17642);
and U21520 (N_21520,N_18731,N_17194);
nand U21521 (N_21521,N_16217,N_16283);
or U21522 (N_21522,N_18571,N_17554);
nor U21523 (N_21523,N_18246,N_18348);
or U21524 (N_21524,N_18729,N_18204);
nor U21525 (N_21525,N_17404,N_17653);
nor U21526 (N_21526,N_18396,N_16921);
nor U21527 (N_21527,N_16043,N_15736);
nor U21528 (N_21528,N_17832,N_15880);
nand U21529 (N_21529,N_16163,N_16792);
nand U21530 (N_21530,N_16286,N_18427);
nor U21531 (N_21531,N_16339,N_17809);
or U21532 (N_21532,N_17517,N_16253);
and U21533 (N_21533,N_15867,N_17791);
and U21534 (N_21534,N_18111,N_16176);
or U21535 (N_21535,N_17290,N_17301);
nor U21536 (N_21536,N_18042,N_18187);
and U21537 (N_21537,N_18373,N_16682);
nor U21538 (N_21538,N_15685,N_16602);
and U21539 (N_21539,N_17582,N_18504);
nor U21540 (N_21540,N_17300,N_15809);
or U21541 (N_21541,N_17611,N_17876);
xnor U21542 (N_21542,N_18711,N_15702);
nand U21543 (N_21543,N_16744,N_18333);
nor U21544 (N_21544,N_17254,N_16474);
nand U21545 (N_21545,N_17898,N_18676);
and U21546 (N_21546,N_18657,N_15905);
xnor U21547 (N_21547,N_17353,N_15977);
nor U21548 (N_21548,N_17860,N_15969);
nor U21549 (N_21549,N_16550,N_18437);
and U21550 (N_21550,N_16763,N_16504);
nand U21551 (N_21551,N_18026,N_17840);
and U21552 (N_21552,N_17708,N_15902);
and U21553 (N_21553,N_16689,N_18745);
or U21554 (N_21554,N_17459,N_16035);
nand U21555 (N_21555,N_17568,N_18447);
or U21556 (N_21556,N_17771,N_16165);
and U21557 (N_21557,N_17769,N_18328);
and U21558 (N_21558,N_17999,N_16988);
and U21559 (N_21559,N_17394,N_16253);
nand U21560 (N_21560,N_18185,N_18108);
xor U21561 (N_21561,N_18399,N_16070);
xnor U21562 (N_21562,N_17313,N_16916);
or U21563 (N_21563,N_17098,N_15827);
nand U21564 (N_21564,N_17923,N_17271);
xor U21565 (N_21565,N_16094,N_17443);
nor U21566 (N_21566,N_16418,N_18405);
nor U21567 (N_21567,N_16388,N_16458);
xor U21568 (N_21568,N_17646,N_15784);
and U21569 (N_21569,N_18146,N_17645);
xor U21570 (N_21570,N_17775,N_18242);
nand U21571 (N_21571,N_18458,N_15898);
and U21572 (N_21572,N_16973,N_17340);
nor U21573 (N_21573,N_16964,N_17993);
nand U21574 (N_21574,N_16005,N_18551);
nand U21575 (N_21575,N_16450,N_18434);
xor U21576 (N_21576,N_17302,N_17218);
and U21577 (N_21577,N_17613,N_17387);
nor U21578 (N_21578,N_17936,N_17813);
or U21579 (N_21579,N_17804,N_18468);
nor U21580 (N_21580,N_17920,N_18307);
xnor U21581 (N_21581,N_15627,N_17298);
nor U21582 (N_21582,N_18367,N_18251);
nor U21583 (N_21583,N_16994,N_16948);
xnor U21584 (N_21584,N_18715,N_17270);
or U21585 (N_21585,N_18681,N_16148);
and U21586 (N_21586,N_16148,N_17239);
and U21587 (N_21587,N_17060,N_16794);
nand U21588 (N_21588,N_17674,N_17662);
and U21589 (N_21589,N_16360,N_17441);
nor U21590 (N_21590,N_18174,N_17275);
and U21591 (N_21591,N_18061,N_15827);
xnor U21592 (N_21592,N_18567,N_18568);
nand U21593 (N_21593,N_16188,N_17258);
nand U21594 (N_21594,N_18478,N_18382);
and U21595 (N_21595,N_16014,N_16532);
and U21596 (N_21596,N_18555,N_16548);
or U21597 (N_21597,N_18176,N_17522);
nor U21598 (N_21598,N_16648,N_17844);
or U21599 (N_21599,N_16951,N_15996);
nor U21600 (N_21600,N_17055,N_16558);
and U21601 (N_21601,N_17359,N_17672);
or U21602 (N_21602,N_16848,N_16307);
xor U21603 (N_21603,N_16887,N_17922);
xor U21604 (N_21604,N_15886,N_17515);
nor U21605 (N_21605,N_16557,N_17188);
xor U21606 (N_21606,N_15736,N_17512);
nand U21607 (N_21607,N_17569,N_17833);
nor U21608 (N_21608,N_18384,N_16566);
xnor U21609 (N_21609,N_16203,N_16427);
and U21610 (N_21610,N_15764,N_15938);
xor U21611 (N_21611,N_18544,N_15677);
xnor U21612 (N_21612,N_16450,N_15915);
nand U21613 (N_21613,N_18048,N_17431);
or U21614 (N_21614,N_16907,N_16858);
nor U21615 (N_21615,N_16791,N_16166);
and U21616 (N_21616,N_16530,N_17335);
and U21617 (N_21617,N_17273,N_18269);
nor U21618 (N_21618,N_16251,N_17068);
and U21619 (N_21619,N_17182,N_16452);
and U21620 (N_21620,N_16607,N_17773);
nand U21621 (N_21621,N_17201,N_16020);
nor U21622 (N_21622,N_16192,N_18098);
xnor U21623 (N_21623,N_17483,N_17670);
nor U21624 (N_21624,N_17199,N_16930);
or U21625 (N_21625,N_17570,N_18140);
nor U21626 (N_21626,N_17746,N_17026);
nand U21627 (N_21627,N_17770,N_18414);
and U21628 (N_21628,N_16367,N_16840);
and U21629 (N_21629,N_18604,N_16002);
nor U21630 (N_21630,N_17242,N_16751);
nand U21631 (N_21631,N_17483,N_18037);
or U21632 (N_21632,N_16518,N_18204);
and U21633 (N_21633,N_16424,N_17696);
or U21634 (N_21634,N_15807,N_17690);
and U21635 (N_21635,N_16988,N_16521);
or U21636 (N_21636,N_18396,N_18512);
nand U21637 (N_21637,N_16687,N_18421);
nor U21638 (N_21638,N_18498,N_16985);
or U21639 (N_21639,N_17893,N_18406);
and U21640 (N_21640,N_18088,N_18053);
and U21641 (N_21641,N_16650,N_18377);
and U21642 (N_21642,N_18498,N_15849);
nor U21643 (N_21643,N_18622,N_17336);
nand U21644 (N_21644,N_17068,N_15834);
or U21645 (N_21645,N_18075,N_16663);
xor U21646 (N_21646,N_18268,N_16433);
nor U21647 (N_21647,N_17081,N_18594);
nand U21648 (N_21648,N_15936,N_15682);
or U21649 (N_21649,N_18553,N_18635);
xnor U21650 (N_21650,N_16481,N_18120);
nand U21651 (N_21651,N_17631,N_18079);
xnor U21652 (N_21652,N_16874,N_16728);
nand U21653 (N_21653,N_18666,N_17332);
nand U21654 (N_21654,N_17002,N_16174);
nor U21655 (N_21655,N_18483,N_16084);
and U21656 (N_21656,N_16374,N_16737);
xnor U21657 (N_21657,N_17783,N_16049);
nor U21658 (N_21658,N_17175,N_17656);
nand U21659 (N_21659,N_17897,N_16718);
nand U21660 (N_21660,N_16743,N_17941);
and U21661 (N_21661,N_15893,N_17105);
or U21662 (N_21662,N_15794,N_17498);
and U21663 (N_21663,N_16340,N_16720);
nand U21664 (N_21664,N_17794,N_16783);
xor U21665 (N_21665,N_16614,N_18727);
or U21666 (N_21666,N_18166,N_18462);
nor U21667 (N_21667,N_16320,N_18220);
nor U21668 (N_21668,N_17845,N_16643);
nand U21669 (N_21669,N_17616,N_16642);
and U21670 (N_21670,N_17903,N_16015);
and U21671 (N_21671,N_15731,N_17442);
and U21672 (N_21672,N_16999,N_17847);
or U21673 (N_21673,N_16164,N_16822);
nand U21674 (N_21674,N_18296,N_16244);
and U21675 (N_21675,N_18730,N_17855);
or U21676 (N_21676,N_16510,N_18086);
xnor U21677 (N_21677,N_16671,N_17227);
or U21678 (N_21678,N_17029,N_17555);
nand U21679 (N_21679,N_18199,N_18087);
or U21680 (N_21680,N_16098,N_17962);
nor U21681 (N_21681,N_15973,N_16936);
nand U21682 (N_21682,N_17255,N_18206);
nand U21683 (N_21683,N_17529,N_15912);
nor U21684 (N_21684,N_17447,N_18595);
xnor U21685 (N_21685,N_16591,N_16846);
nor U21686 (N_21686,N_16101,N_16698);
nor U21687 (N_21687,N_16691,N_16004);
or U21688 (N_21688,N_16849,N_17951);
xor U21689 (N_21689,N_17946,N_18221);
and U21690 (N_21690,N_17502,N_17937);
and U21691 (N_21691,N_18241,N_17842);
nand U21692 (N_21692,N_16287,N_17710);
and U21693 (N_21693,N_17900,N_17516);
xor U21694 (N_21694,N_15650,N_16606);
or U21695 (N_21695,N_16835,N_18432);
nor U21696 (N_21696,N_17911,N_18061);
nand U21697 (N_21697,N_16951,N_15839);
nor U21698 (N_21698,N_18653,N_16143);
nand U21699 (N_21699,N_18487,N_18216);
and U21700 (N_21700,N_18228,N_17413);
or U21701 (N_21701,N_18671,N_16765);
or U21702 (N_21702,N_18349,N_17943);
nor U21703 (N_21703,N_16554,N_18633);
or U21704 (N_21704,N_17200,N_16408);
xor U21705 (N_21705,N_18018,N_16421);
nand U21706 (N_21706,N_16770,N_18612);
and U21707 (N_21707,N_16611,N_17335);
nand U21708 (N_21708,N_17447,N_18367);
or U21709 (N_21709,N_18485,N_17618);
or U21710 (N_21710,N_18366,N_17800);
and U21711 (N_21711,N_17450,N_15695);
xor U21712 (N_21712,N_17641,N_16468);
or U21713 (N_21713,N_18388,N_17296);
and U21714 (N_21714,N_17220,N_18204);
nand U21715 (N_21715,N_17332,N_16702);
xnor U21716 (N_21716,N_16355,N_16032);
or U21717 (N_21717,N_16658,N_16560);
and U21718 (N_21718,N_15917,N_18712);
xor U21719 (N_21719,N_17375,N_16615);
nor U21720 (N_21720,N_18155,N_16791);
nand U21721 (N_21721,N_17655,N_17429);
nor U21722 (N_21722,N_17250,N_17749);
xor U21723 (N_21723,N_16316,N_16167);
nor U21724 (N_21724,N_15770,N_16359);
or U21725 (N_21725,N_15653,N_17416);
or U21726 (N_21726,N_15861,N_18353);
and U21727 (N_21727,N_18379,N_17869);
or U21728 (N_21728,N_16159,N_16555);
xnor U21729 (N_21729,N_17395,N_17437);
nand U21730 (N_21730,N_17786,N_16906);
nor U21731 (N_21731,N_16682,N_16536);
or U21732 (N_21732,N_16391,N_17403);
xnor U21733 (N_21733,N_15727,N_17962);
and U21734 (N_21734,N_17948,N_17001);
nand U21735 (N_21735,N_18446,N_17356);
and U21736 (N_21736,N_17942,N_18148);
nand U21737 (N_21737,N_17814,N_15788);
xor U21738 (N_21738,N_16286,N_17193);
nand U21739 (N_21739,N_18427,N_18707);
and U21740 (N_21740,N_16509,N_18508);
xnor U21741 (N_21741,N_15757,N_16639);
and U21742 (N_21742,N_17562,N_18391);
or U21743 (N_21743,N_16644,N_18077);
or U21744 (N_21744,N_18491,N_16767);
nand U21745 (N_21745,N_15647,N_16798);
or U21746 (N_21746,N_17985,N_17419);
nor U21747 (N_21747,N_17355,N_17648);
or U21748 (N_21748,N_18316,N_17362);
xor U21749 (N_21749,N_17488,N_15644);
xnor U21750 (N_21750,N_16314,N_17406);
and U21751 (N_21751,N_16648,N_16234);
nand U21752 (N_21752,N_18287,N_17642);
nor U21753 (N_21753,N_18486,N_18262);
and U21754 (N_21754,N_16049,N_18529);
nor U21755 (N_21755,N_15641,N_17254);
nor U21756 (N_21756,N_16504,N_18363);
and U21757 (N_21757,N_16907,N_15980);
xnor U21758 (N_21758,N_15856,N_17294);
and U21759 (N_21759,N_16312,N_16332);
or U21760 (N_21760,N_16242,N_18046);
and U21761 (N_21761,N_17785,N_16021);
nand U21762 (N_21762,N_15813,N_16581);
and U21763 (N_21763,N_16934,N_16285);
nor U21764 (N_21764,N_15962,N_17851);
xor U21765 (N_21765,N_18669,N_17949);
and U21766 (N_21766,N_17951,N_18332);
nor U21767 (N_21767,N_16311,N_18613);
nor U21768 (N_21768,N_16155,N_17764);
nor U21769 (N_21769,N_17930,N_18063);
or U21770 (N_21770,N_16914,N_15953);
and U21771 (N_21771,N_17722,N_17869);
nand U21772 (N_21772,N_15975,N_16979);
or U21773 (N_21773,N_17228,N_16072);
and U21774 (N_21774,N_17119,N_17935);
nor U21775 (N_21775,N_18334,N_18611);
xnor U21776 (N_21776,N_18286,N_17482);
xnor U21777 (N_21777,N_18098,N_16111);
nand U21778 (N_21778,N_16565,N_16350);
xnor U21779 (N_21779,N_17133,N_18052);
nor U21780 (N_21780,N_17476,N_18265);
nor U21781 (N_21781,N_18354,N_16290);
nor U21782 (N_21782,N_16398,N_17989);
nand U21783 (N_21783,N_17622,N_17438);
or U21784 (N_21784,N_17622,N_17040);
nand U21785 (N_21785,N_18267,N_16038);
or U21786 (N_21786,N_17028,N_16274);
xnor U21787 (N_21787,N_17177,N_17987);
nand U21788 (N_21788,N_17051,N_15922);
nand U21789 (N_21789,N_16533,N_18062);
nand U21790 (N_21790,N_17265,N_17492);
and U21791 (N_21791,N_18526,N_18218);
nand U21792 (N_21792,N_18239,N_15699);
or U21793 (N_21793,N_17674,N_15647);
and U21794 (N_21794,N_17411,N_17761);
nand U21795 (N_21795,N_18348,N_15873);
nand U21796 (N_21796,N_16707,N_17742);
nor U21797 (N_21797,N_16820,N_15877);
nand U21798 (N_21798,N_17017,N_18484);
or U21799 (N_21799,N_17238,N_18052);
xnor U21800 (N_21800,N_16463,N_18518);
xor U21801 (N_21801,N_17040,N_15645);
nor U21802 (N_21802,N_16738,N_18227);
xor U21803 (N_21803,N_17884,N_18587);
xnor U21804 (N_21804,N_17018,N_16829);
nor U21805 (N_21805,N_18458,N_17064);
nand U21806 (N_21806,N_16654,N_17549);
nand U21807 (N_21807,N_18401,N_18307);
nor U21808 (N_21808,N_18004,N_16894);
xor U21809 (N_21809,N_18004,N_18694);
nor U21810 (N_21810,N_17826,N_18580);
xnor U21811 (N_21811,N_18085,N_17243);
nor U21812 (N_21812,N_17323,N_18539);
xor U21813 (N_21813,N_17546,N_15668);
xor U21814 (N_21814,N_15892,N_18042);
nor U21815 (N_21815,N_16223,N_16326);
and U21816 (N_21816,N_18489,N_17172);
xnor U21817 (N_21817,N_16640,N_16771);
nand U21818 (N_21818,N_15697,N_15847);
xor U21819 (N_21819,N_16137,N_15714);
and U21820 (N_21820,N_17963,N_16455);
xor U21821 (N_21821,N_15704,N_18277);
or U21822 (N_21822,N_16596,N_17541);
nand U21823 (N_21823,N_17602,N_18052);
nand U21824 (N_21824,N_17492,N_15876);
and U21825 (N_21825,N_17523,N_16865);
xor U21826 (N_21826,N_17002,N_18474);
nor U21827 (N_21827,N_16863,N_18725);
xor U21828 (N_21828,N_18040,N_16903);
and U21829 (N_21829,N_18192,N_18567);
or U21830 (N_21830,N_17687,N_16819);
nor U21831 (N_21831,N_16860,N_16426);
xor U21832 (N_21832,N_16563,N_17508);
or U21833 (N_21833,N_18550,N_18505);
nor U21834 (N_21834,N_17351,N_17154);
and U21835 (N_21835,N_16901,N_18612);
xnor U21836 (N_21836,N_18373,N_18475);
or U21837 (N_21837,N_16866,N_16856);
and U21838 (N_21838,N_16001,N_17351);
and U21839 (N_21839,N_18281,N_17499);
nor U21840 (N_21840,N_17363,N_17339);
nand U21841 (N_21841,N_16995,N_18240);
xor U21842 (N_21842,N_17641,N_18190);
and U21843 (N_21843,N_16474,N_16862);
or U21844 (N_21844,N_18057,N_17387);
and U21845 (N_21845,N_16808,N_15947);
xnor U21846 (N_21846,N_17461,N_17049);
nand U21847 (N_21847,N_16908,N_16299);
xnor U21848 (N_21848,N_15938,N_17883);
nor U21849 (N_21849,N_17744,N_15899);
nor U21850 (N_21850,N_15954,N_15848);
nor U21851 (N_21851,N_18133,N_16237);
nand U21852 (N_21852,N_16180,N_17214);
or U21853 (N_21853,N_18126,N_18450);
nand U21854 (N_21854,N_15823,N_18422);
nand U21855 (N_21855,N_17728,N_18090);
and U21856 (N_21856,N_15867,N_17162);
or U21857 (N_21857,N_15891,N_18056);
nor U21858 (N_21858,N_18661,N_18282);
and U21859 (N_21859,N_15651,N_18274);
or U21860 (N_21860,N_17843,N_16686);
and U21861 (N_21861,N_18247,N_15743);
or U21862 (N_21862,N_16562,N_18589);
nand U21863 (N_21863,N_16671,N_17827);
and U21864 (N_21864,N_17548,N_16956);
and U21865 (N_21865,N_16152,N_15775);
xnor U21866 (N_21866,N_18138,N_18134);
or U21867 (N_21867,N_18626,N_15790);
or U21868 (N_21868,N_16348,N_18062);
and U21869 (N_21869,N_15898,N_15730);
nor U21870 (N_21870,N_17963,N_16909);
nor U21871 (N_21871,N_16834,N_17196);
or U21872 (N_21872,N_17855,N_15628);
and U21873 (N_21873,N_17586,N_16985);
nor U21874 (N_21874,N_16376,N_17057);
nand U21875 (N_21875,N_18802,N_21621);
or U21876 (N_21876,N_19255,N_20076);
nand U21877 (N_21877,N_20959,N_21619);
nand U21878 (N_21878,N_20659,N_19478);
and U21879 (N_21879,N_20316,N_21831);
and U21880 (N_21880,N_19900,N_19110);
or U21881 (N_21881,N_20674,N_19233);
and U21882 (N_21882,N_20779,N_21008);
nand U21883 (N_21883,N_19827,N_19027);
xnor U21884 (N_21884,N_21862,N_21517);
nand U21885 (N_21885,N_18835,N_19712);
nand U21886 (N_21886,N_20236,N_19582);
and U21887 (N_21887,N_20960,N_21686);
nor U21888 (N_21888,N_19783,N_20664);
xor U21889 (N_21889,N_20486,N_19336);
xor U21890 (N_21890,N_21440,N_20349);
xnor U21891 (N_21891,N_21286,N_21179);
or U21892 (N_21892,N_21501,N_20689);
nand U21893 (N_21893,N_19050,N_18768);
and U21894 (N_21894,N_19412,N_19379);
nand U21895 (N_21895,N_21403,N_19766);
xor U21896 (N_21896,N_18757,N_19654);
nor U21897 (N_21897,N_19554,N_21860);
xor U21898 (N_21898,N_20625,N_19703);
and U21899 (N_21899,N_18910,N_20690);
nand U21900 (N_21900,N_21184,N_20116);
and U21901 (N_21901,N_18939,N_20729);
and U21902 (N_21902,N_19548,N_18997);
and U21903 (N_21903,N_19729,N_19293);
nand U21904 (N_21904,N_19687,N_19552);
and U21905 (N_21905,N_20113,N_19365);
and U21906 (N_21906,N_21176,N_21005);
xnor U21907 (N_21907,N_20547,N_19203);
xor U21908 (N_21908,N_19580,N_20623);
nor U21909 (N_21909,N_21788,N_19467);
xnor U21910 (N_21910,N_21525,N_21052);
or U21911 (N_21911,N_20152,N_19061);
and U21912 (N_21912,N_20816,N_19571);
nand U21913 (N_21913,N_21426,N_19794);
or U21914 (N_21914,N_20418,N_19830);
nand U21915 (N_21915,N_20315,N_18914);
nor U21916 (N_21916,N_20091,N_19640);
nor U21917 (N_21917,N_21596,N_20396);
xnor U21918 (N_21918,N_19182,N_20600);
nor U21919 (N_21919,N_18862,N_19925);
or U21920 (N_21920,N_21233,N_20943);
or U21921 (N_21921,N_21528,N_20063);
xor U21922 (N_21922,N_19612,N_21143);
xnor U21923 (N_21923,N_20071,N_20042);
and U21924 (N_21924,N_18787,N_18796);
nor U21925 (N_21925,N_20074,N_20484);
xnor U21926 (N_21926,N_20402,N_19496);
nand U21927 (N_21927,N_18853,N_21503);
nand U21928 (N_21928,N_21427,N_19284);
nand U21929 (N_21929,N_21420,N_19948);
nand U21930 (N_21930,N_19859,N_20187);
and U21931 (N_21931,N_19710,N_21119);
xor U21932 (N_21932,N_21785,N_21077);
and U21933 (N_21933,N_20324,N_21446);
or U21934 (N_21934,N_21188,N_19808);
xnor U21935 (N_21935,N_21631,N_20475);
or U21936 (N_21936,N_19502,N_21173);
and U21937 (N_21937,N_18903,N_19305);
nor U21938 (N_21938,N_20066,N_21057);
nor U21939 (N_21939,N_18842,N_20836);
and U21940 (N_21940,N_20250,N_19306);
nor U21941 (N_21941,N_19286,N_20967);
xor U21942 (N_21942,N_21402,N_18826);
nor U21943 (N_21943,N_19706,N_19234);
nor U21944 (N_21944,N_21358,N_21062);
nand U21945 (N_21945,N_19810,N_21130);
nand U21946 (N_21946,N_19367,N_20764);
and U21947 (N_21947,N_21813,N_20183);
or U21948 (N_21948,N_18893,N_21527);
or U21949 (N_21949,N_20523,N_20920);
xor U21950 (N_21950,N_19457,N_21676);
xor U21951 (N_21951,N_20902,N_20753);
and U21952 (N_21952,N_19121,N_21393);
and U21953 (N_21953,N_19297,N_19184);
nand U21954 (N_21954,N_20509,N_20574);
nand U21955 (N_21955,N_21304,N_20782);
nand U21956 (N_21956,N_19299,N_20085);
xnor U21957 (N_21957,N_21565,N_19991);
xor U21958 (N_21958,N_19949,N_19543);
xnor U21959 (N_21959,N_19635,N_19483);
and U21960 (N_21960,N_20134,N_19103);
or U21961 (N_21961,N_19285,N_20846);
or U21962 (N_21962,N_20772,N_21209);
nand U21963 (N_21963,N_20388,N_19556);
or U21964 (N_21964,N_19106,N_21362);
xnor U21965 (N_21965,N_21083,N_21064);
xnor U21966 (N_21966,N_19875,N_21482);
nand U21967 (N_21967,N_21486,N_18815);
and U21968 (N_21968,N_19417,N_21659);
nand U21969 (N_21969,N_19340,N_21193);
or U21970 (N_21970,N_21037,N_18917);
nor U21971 (N_21971,N_20064,N_21855);
xnor U21972 (N_21972,N_19484,N_21392);
and U21973 (N_21973,N_19490,N_19091);
nand U21974 (N_21974,N_20551,N_19388);
nand U21975 (N_21975,N_20898,N_19998);
and U21976 (N_21976,N_20459,N_21727);
nor U21977 (N_21977,N_21725,N_19081);
or U21978 (N_21978,N_19385,N_20221);
nand U21979 (N_21979,N_19972,N_21397);
nand U21980 (N_21980,N_21866,N_19252);
xor U21981 (N_21981,N_21016,N_21459);
xnor U21982 (N_21982,N_20518,N_20696);
and U21983 (N_21983,N_19598,N_19207);
nor U21984 (N_21984,N_21322,N_21371);
xnor U21985 (N_21985,N_20421,N_21776);
and U21986 (N_21986,N_19476,N_19149);
and U21987 (N_21987,N_19592,N_19477);
nand U21988 (N_21988,N_19220,N_19368);
and U21989 (N_21989,N_19696,N_20254);
or U21990 (N_21990,N_20088,N_21638);
or U21991 (N_21991,N_19115,N_19173);
xnor U21992 (N_21992,N_20617,N_19782);
or U21993 (N_21993,N_21819,N_20011);
xnor U21994 (N_21994,N_20525,N_21049);
nor U21995 (N_21995,N_19382,N_20142);
nor U21996 (N_21996,N_19452,N_19242);
and U21997 (N_21997,N_20800,N_20302);
or U21998 (N_21998,N_21718,N_20885);
or U21999 (N_21999,N_21555,N_20997);
xnor U22000 (N_22000,N_20756,N_19716);
xnor U22001 (N_22001,N_19017,N_21107);
or U22002 (N_22002,N_19694,N_21025);
xnor U22003 (N_22003,N_20268,N_20407);
or U22004 (N_22004,N_19812,N_19596);
nor U22005 (N_22005,N_19021,N_20876);
and U22006 (N_22006,N_19239,N_20942);
and U22007 (N_22007,N_21096,N_19553);
and U22008 (N_22008,N_21734,N_20680);
nor U22009 (N_22009,N_19053,N_20133);
and U22010 (N_22010,N_21045,N_20629);
or U22011 (N_22011,N_19228,N_20605);
and U22012 (N_22012,N_21637,N_20383);
and U22013 (N_22013,N_21783,N_21000);
nand U22014 (N_22014,N_19399,N_20734);
nor U22015 (N_22015,N_21236,N_18790);
and U22016 (N_22016,N_20192,N_20539);
nor U22017 (N_22017,N_21810,N_19271);
xor U22018 (N_22018,N_21138,N_19424);
nand U22019 (N_22019,N_21593,N_21758);
nor U22020 (N_22020,N_19265,N_21273);
xnor U22021 (N_22021,N_20544,N_19408);
or U22022 (N_22022,N_21227,N_18913);
nor U22023 (N_22023,N_19260,N_19682);
and U22024 (N_22024,N_20498,N_19042);
nand U22025 (N_22025,N_20098,N_21518);
xor U22026 (N_22026,N_21566,N_18872);
nand U22027 (N_22027,N_19311,N_21690);
or U22028 (N_22028,N_21381,N_19443);
and U22029 (N_22029,N_20904,N_18904);
nand U22030 (N_22030,N_19451,N_19908);
nor U22031 (N_22031,N_20058,N_20826);
or U22032 (N_22032,N_21089,N_19083);
or U22033 (N_22033,N_19626,N_20233);
or U22034 (N_22034,N_19796,N_21048);
and U22035 (N_22035,N_20333,N_21443);
nand U22036 (N_22036,N_20665,N_21042);
nand U22037 (N_22037,N_19076,N_20430);
and U22038 (N_22038,N_18991,N_20285);
or U22039 (N_22039,N_19790,N_20075);
or U22040 (N_22040,N_20080,N_21159);
and U22041 (N_22041,N_20062,N_19613);
nand U22042 (N_22042,N_18763,N_19851);
nand U22043 (N_22043,N_19179,N_20578);
nand U22044 (N_22044,N_18854,N_19301);
xor U22045 (N_22045,N_19079,N_19878);
or U22046 (N_22046,N_21623,N_20613);
or U22047 (N_22047,N_20334,N_19604);
nand U22048 (N_22048,N_20561,N_21705);
and U22049 (N_22049,N_20542,N_21870);
nor U22050 (N_22050,N_19890,N_20855);
nand U22051 (N_22051,N_19289,N_18797);
and U22052 (N_22052,N_18990,N_20745);
xor U22053 (N_22053,N_21390,N_20595);
nand U22054 (N_22054,N_19531,N_21334);
or U22055 (N_22055,N_19806,N_20274);
and U22056 (N_22056,N_21697,N_19307);
and U22057 (N_22057,N_21850,N_21241);
nor U22058 (N_22058,N_19269,N_18901);
xnor U22059 (N_22059,N_19150,N_18843);
and U22060 (N_22060,N_19309,N_21075);
nand U22061 (N_22061,N_19397,N_20568);
nor U22062 (N_22062,N_20679,N_20419);
and U22063 (N_22063,N_21421,N_21435);
nor U22064 (N_22064,N_19735,N_21071);
or U22065 (N_22065,N_19159,N_20773);
xor U22066 (N_22066,N_20082,N_21191);
nand U22067 (N_22067,N_20003,N_19282);
or U22068 (N_22068,N_20394,N_18935);
nor U22069 (N_22069,N_19358,N_21803);
nand U22070 (N_22070,N_20515,N_19049);
nand U22071 (N_22071,N_18943,N_20079);
or U22072 (N_22072,N_21352,N_19300);
nand U22073 (N_22073,N_21768,N_20345);
nand U22074 (N_22074,N_20797,N_20768);
or U22075 (N_22075,N_19009,N_19739);
nor U22076 (N_22076,N_21259,N_18760);
xor U22077 (N_22077,N_21551,N_21532);
and U22078 (N_22078,N_19322,N_21576);
nor U22079 (N_22079,N_18955,N_19855);
xor U22080 (N_22080,N_20446,N_19482);
nor U22081 (N_22081,N_21124,N_19670);
or U22082 (N_22082,N_19429,N_20541);
or U22083 (N_22083,N_19369,N_20491);
or U22084 (N_22084,N_20359,N_20443);
and U22085 (N_22085,N_20757,N_20497);
nand U22086 (N_22086,N_19883,N_21232);
nor U22087 (N_22087,N_21800,N_21234);
nor U22088 (N_22088,N_21467,N_20969);
xnor U22089 (N_22089,N_19579,N_21268);
and U22090 (N_22090,N_20645,N_20417);
nand U22091 (N_22091,N_21260,N_19718);
nand U22092 (N_22092,N_19702,N_20266);
or U22093 (N_22093,N_19352,N_18941);
or U22094 (N_22094,N_20951,N_21756);
xnor U22095 (N_22095,N_21290,N_21363);
or U22096 (N_22096,N_19950,N_19688);
nand U22097 (N_22097,N_19987,N_21592);
nand U22098 (N_22098,N_20611,N_20461);
nand U22099 (N_22099,N_21340,N_20211);
xnor U22100 (N_22100,N_18944,N_21308);
nor U22101 (N_22101,N_20607,N_20338);
and U22102 (N_22102,N_21847,N_19409);
and U22103 (N_22103,N_19200,N_20146);
xor U22104 (N_22104,N_19118,N_18861);
xnor U22105 (N_22105,N_19188,N_20464);
or U22106 (N_22106,N_19161,N_21269);
or U22107 (N_22107,N_18771,N_20812);
xnor U22108 (N_22108,N_19815,N_21198);
nor U22109 (N_22109,N_20207,N_20549);
nand U22110 (N_22110,N_19054,N_21226);
nand U22111 (N_22111,N_21452,N_18887);
xnor U22112 (N_22112,N_21732,N_21121);
or U22113 (N_22113,N_20478,N_19785);
or U22114 (N_22114,N_20787,N_19099);
xor U22115 (N_22115,N_19226,N_21744);
xnor U22116 (N_22116,N_20169,N_20462);
nor U22117 (N_22117,N_21055,N_21513);
nand U22118 (N_22118,N_20286,N_19519);
xor U22119 (N_22119,N_20685,N_21182);
or U22120 (N_22120,N_21787,N_20103);
nor U22121 (N_22121,N_20013,N_21349);
and U22122 (N_22122,N_19243,N_20114);
and U22123 (N_22123,N_18954,N_18924);
xnor U22124 (N_22124,N_20073,N_18858);
nor U22125 (N_22125,N_18986,N_19669);
nand U22126 (N_22126,N_20119,N_19655);
nor U22127 (N_22127,N_20526,N_19120);
nor U22128 (N_22128,N_20360,N_21816);
and U22129 (N_22129,N_20310,N_18844);
or U22130 (N_22130,N_18918,N_20155);
or U22131 (N_22131,N_18801,N_20317);
nand U22132 (N_22132,N_21481,N_20938);
nor U22133 (N_22133,N_19676,N_19555);
nor U22134 (N_22134,N_20930,N_19296);
and U22135 (N_22135,N_19538,N_20229);
nand U22136 (N_22136,N_18788,N_20703);
xor U22137 (N_22137,N_20223,N_20164);
or U22138 (N_22138,N_19075,N_19642);
or U22139 (N_22139,N_20238,N_20809);
or U22140 (N_22140,N_21140,N_18995);
nor U22141 (N_22141,N_20552,N_21713);
and U22142 (N_22142,N_18810,N_21073);
nand U22143 (N_22143,N_20190,N_21624);
nand U22144 (N_22144,N_21583,N_21058);
nand U22145 (N_22145,N_20594,N_19673);
or U22146 (N_22146,N_21320,N_19277);
nor U22147 (N_22147,N_21142,N_20852);
or U22148 (N_22148,N_19880,N_20260);
xor U22149 (N_22149,N_21200,N_20993);
nand U22150 (N_22150,N_20457,N_19160);
and U22151 (N_22151,N_20487,N_19861);
or U22152 (N_22152,N_19512,N_20982);
or U22153 (N_22153,N_20751,N_20014);
nor U22154 (N_22154,N_19737,N_18833);
nor U22155 (N_22155,N_18850,N_19990);
and U22156 (N_22156,N_21346,N_18908);
nand U22157 (N_22157,N_18951,N_21171);
xor U22158 (N_22158,N_21401,N_18965);
nand U22159 (N_22159,N_21004,N_20635);
and U22160 (N_22160,N_21097,N_20466);
and U22161 (N_22161,N_20044,N_21802);
nor U22162 (N_22162,N_21586,N_18895);
and U22163 (N_22163,N_20506,N_21139);
or U22164 (N_22164,N_19614,N_21125);
or U22165 (N_22165,N_21265,N_19196);
or U22166 (N_22166,N_19711,N_20378);
xor U22167 (N_22167,N_20206,N_21298);
or U22168 (N_22168,N_20510,N_19544);
and U22169 (N_22169,N_21656,N_20814);
xnor U22170 (N_22170,N_21693,N_19937);
and U22171 (N_22171,N_20507,N_20175);
and U22172 (N_22172,N_21854,N_20234);
nand U22173 (N_22173,N_19947,N_19479);
nor U22174 (N_22174,N_20513,N_19852);
and U22175 (N_22175,N_21509,N_21837);
or U22176 (N_22176,N_20556,N_19195);
nand U22177 (N_22177,N_19036,N_21332);
or U22178 (N_22178,N_20222,N_21526);
nand U22179 (N_22179,N_20592,N_19974);
or U22180 (N_22180,N_21495,N_21047);
and U22181 (N_22181,N_19574,N_21530);
or U22182 (N_22182,N_21344,N_19862);
and U22183 (N_22183,N_21264,N_19371);
xnor U22184 (N_22184,N_21228,N_19051);
xnor U22185 (N_22185,N_19982,N_19455);
nor U22186 (N_22186,N_20865,N_21741);
xnor U22187 (N_22187,N_18814,N_19924);
xnor U22188 (N_22188,N_21533,N_20534);
nand U22189 (N_22189,N_20061,N_20186);
and U22190 (N_22190,N_19456,N_19645);
xor U22191 (N_22191,N_20973,N_19419);
xnor U22192 (N_22192,N_21502,N_21582);
nor U22193 (N_22193,N_21326,N_19641);
or U22194 (N_22194,N_21164,N_19074);
nand U22195 (N_22195,N_20707,N_20356);
xor U22196 (N_22196,N_20301,N_19540);
xor U22197 (N_22197,N_20963,N_21506);
nor U22198 (N_22198,N_20130,N_20488);
and U22199 (N_22199,N_21563,N_21464);
nor U22200 (N_22200,N_19686,N_19679);
and U22201 (N_22201,N_21794,N_21155);
xor U22202 (N_22202,N_18994,N_20131);
nor U22203 (N_22203,N_19910,N_19324);
or U22204 (N_22204,N_20649,N_20143);
xor U22205 (N_22205,N_19444,N_21126);
or U22206 (N_22206,N_19868,N_21818);
and U22207 (N_22207,N_19332,N_21861);
nor U22208 (N_22208,N_20666,N_20099);
nand U22209 (N_22209,N_20343,N_19691);
nor U22210 (N_22210,N_20639,N_21400);
nand U22211 (N_22211,N_21508,N_20330);
nor U22212 (N_22212,N_18829,N_20616);
nor U22213 (N_22213,N_19524,N_20282);
nand U22214 (N_22214,N_21106,N_21812);
nand U22215 (N_22215,N_20598,N_21535);
and U22216 (N_22216,N_20124,N_21383);
xnor U22217 (N_22217,N_19903,N_18778);
or U22218 (N_22218,N_19077,N_19295);
nor U22219 (N_22219,N_19917,N_20147);
nor U22220 (N_22220,N_20397,N_20636);
and U22221 (N_22221,N_19393,N_19646);
nor U22222 (N_22222,N_19130,N_21257);
xor U22223 (N_22223,N_20725,N_21858);
or U22224 (N_22224,N_18774,N_19404);
nor U22225 (N_22225,N_21019,N_19142);
xnor U22226 (N_22226,N_19189,N_20035);
or U22227 (N_22227,N_20804,N_21289);
nor U22228 (N_22228,N_19559,N_19517);
xnor U22229 (N_22229,N_20029,N_20803);
nand U22230 (N_22230,N_19698,N_21463);
and U22231 (N_22231,N_21645,N_19122);
and U22232 (N_22232,N_20723,N_19867);
xnor U22233 (N_22233,N_19532,N_21069);
nor U22234 (N_22234,N_19270,N_21374);
or U22235 (N_22235,N_19597,N_21183);
or U22236 (N_22236,N_20253,N_19897);
xor U22237 (N_22237,N_18899,N_21492);
or U22238 (N_22238,N_20882,N_19759);
xnor U22239 (N_22239,N_20365,N_19979);
or U22240 (N_22240,N_21274,N_21429);
nor U22241 (N_22241,N_19733,N_18823);
or U22242 (N_22242,N_20886,N_21333);
nand U22243 (N_22243,N_21167,N_19378);
or U22244 (N_22244,N_19885,N_21627);
and U22245 (N_22245,N_21166,N_21605);
and U22246 (N_22246,N_21448,N_18948);
xor U22247 (N_22247,N_20583,N_21033);
and U22248 (N_22248,N_21649,N_21419);
xnor U22249 (N_22249,N_21574,N_20141);
nand U22250 (N_22250,N_20467,N_21197);
and U22251 (N_22251,N_20593,N_19097);
nand U22252 (N_22252,N_20034,N_19899);
and U22253 (N_22253,N_19221,N_19176);
xnor U22254 (N_22254,N_20239,N_21225);
nor U22255 (N_22255,N_19557,N_19153);
xnor U22256 (N_22256,N_18759,N_21086);
nand U22257 (N_22257,N_21512,N_19758);
and U22258 (N_22258,N_20247,N_19154);
nand U22259 (N_22259,N_20601,N_19458);
nor U22260 (N_22260,N_19701,N_19127);
xor U22261 (N_22261,N_21302,N_19063);
nor U22262 (N_22262,N_21564,N_19112);
and U22263 (N_22263,N_18865,N_19978);
nor U22264 (N_22264,N_18945,N_20992);
and U22265 (N_22265,N_21079,N_19390);
nand U22266 (N_22266,N_19955,N_19647);
nor U22267 (N_22267,N_20995,N_18772);
or U22268 (N_22268,N_20572,N_20564);
xor U22269 (N_22269,N_21378,N_20971);
nand U22270 (N_22270,N_20395,N_21472);
and U22271 (N_22271,N_20628,N_19752);
and U22272 (N_22272,N_19506,N_20671);
and U22273 (N_22273,N_18751,N_19466);
nand U22274 (N_22274,N_19750,N_20741);
xnor U22275 (N_22275,N_20217,N_19789);
xnor U22276 (N_22276,N_20300,N_20001);
xor U22277 (N_22277,N_20245,N_21524);
xnor U22278 (N_22278,N_19414,N_21123);
xnor U22279 (N_22279,N_21132,N_21808);
or U22280 (N_22280,N_20382,N_19817);
and U22281 (N_22281,N_20620,N_21796);
nor U22282 (N_22282,N_19108,N_19846);
nor U22283 (N_22283,N_18920,N_21648);
nand U22284 (N_22284,N_19454,N_20670);
and U22285 (N_22285,N_20983,N_19858);
and U22286 (N_22286,N_21723,N_21814);
xnor U22287 (N_22287,N_20482,N_21820);
and U22288 (N_22288,N_20984,N_19799);
xor U22289 (N_22289,N_21061,N_21462);
xnor U22290 (N_22290,N_19771,N_20259);
and U22291 (N_22291,N_19346,N_21505);
nor U22292 (N_22292,N_21380,N_19914);
xor U22293 (N_22293,N_18855,N_19632);
or U22294 (N_22294,N_21792,N_21757);
nor U22295 (N_22295,N_21296,N_19534);
and U22296 (N_22296,N_18938,N_19814);
or U22297 (N_22297,N_21804,N_20759);
nand U22298 (N_22298,N_19029,N_19438);
xor U22299 (N_22299,N_21007,N_21604);
nand U22300 (N_22300,N_21293,N_21835);
nand U22301 (N_22301,N_21375,N_20808);
or U22302 (N_22302,N_19413,N_20137);
or U22303 (N_22303,N_19262,N_21663);
and U22304 (N_22304,N_18874,N_21541);
xor U22305 (N_22305,N_21108,N_20681);
or U22306 (N_22306,N_19767,N_20879);
or U22307 (N_22307,N_20070,N_20232);
xnor U22308 (N_22308,N_21266,N_20615);
or U22309 (N_22309,N_21091,N_21560);
and U22310 (N_22310,N_19832,N_19792);
and U22311 (N_22311,N_20609,N_21147);
xor U22312 (N_22312,N_21626,N_18780);
xnor U22313 (N_22313,N_20604,N_21104);
nand U22314 (N_22314,N_20610,N_18859);
or U22315 (N_22315,N_19335,N_20918);
or U22316 (N_22316,N_19876,N_19705);
nor U22317 (N_22317,N_21010,N_20897);
nor U22318 (N_22318,N_21279,N_21405);
and U22319 (N_22319,N_18761,N_19102);
or U22320 (N_22320,N_21101,N_21367);
or U22321 (N_22321,N_18931,N_21773);
nor U22322 (N_22322,N_20148,N_20145);
and U22323 (N_22323,N_21009,N_19152);
nand U22324 (N_22324,N_21588,N_19866);
or U22325 (N_22325,N_20677,N_19935);
xor U22326 (N_22326,N_21568,N_20658);
or U22327 (N_22327,N_21689,N_20728);
or U22328 (N_22328,N_20543,N_20307);
and U22329 (N_22329,N_21325,N_21616);
and U22330 (N_22330,N_18819,N_21600);
and U22331 (N_22331,N_21186,N_20017);
and U22332 (N_22332,N_21082,N_19728);
xor U22333 (N_22333,N_20669,N_20176);
nor U22334 (N_22334,N_19084,N_21129);
xnor U22335 (N_22335,N_20065,N_20084);
xor U22336 (N_22336,N_19940,N_19700);
nand U22337 (N_22337,N_20810,N_21660);
nand U22338 (N_22338,N_20648,N_21275);
and U22339 (N_22339,N_20706,N_19257);
xnor U22340 (N_22340,N_20807,N_20271);
xnor U22341 (N_22341,N_19965,N_19151);
xnor U22342 (N_22342,N_19717,N_19963);
nor U22343 (N_22343,N_20163,N_21222);
or U22344 (N_22344,N_19630,N_19088);
nand U22345 (N_22345,N_19464,N_21706);
and U22346 (N_22346,N_19396,N_21469);
and U22347 (N_22347,N_20479,N_20566);
nor U22348 (N_22348,N_19845,N_19171);
nor U22349 (N_22349,N_20914,N_18834);
or U22350 (N_22350,N_21211,N_21865);
or U22351 (N_22351,N_20980,N_20101);
xor U22352 (N_22352,N_19653,N_20844);
nor U22353 (N_22353,N_20444,N_21163);
and U22354 (N_22354,N_20102,N_18916);
or U22355 (N_22355,N_19004,N_20866);
nand U22356 (N_22356,N_19601,N_21251);
nand U22357 (N_22357,N_20196,N_21625);
and U22358 (N_22358,N_19374,N_19643);
nor U22359 (N_22359,N_21001,N_19167);
nor U22360 (N_22360,N_20505,N_21500);
or U22361 (N_22361,N_19608,N_21214);
or U22362 (N_22362,N_18851,N_19631);
nor U22363 (N_22363,N_20576,N_20758);
nor U22364 (N_22364,N_19770,N_19680);
and U22365 (N_22365,N_19005,N_21652);
or U22366 (N_22366,N_19319,N_20806);
xnor U22367 (N_22367,N_21704,N_19620);
and U22368 (N_22368,N_19567,N_21746);
and U22369 (N_22369,N_21195,N_19593);
and U22370 (N_22370,N_19435,N_21473);
nand U22371 (N_22371,N_19253,N_21743);
xor U22372 (N_22372,N_18782,N_20893);
or U22373 (N_22373,N_20783,N_20977);
and U22374 (N_22374,N_20744,N_21187);
and U22375 (N_22375,N_18791,N_19287);
nor U22376 (N_22376,N_20536,N_20288);
or U22377 (N_22377,N_20827,N_20654);
xnor U22378 (N_22378,N_21786,N_20754);
and U22379 (N_22379,N_20926,N_21577);
xor U22380 (N_22380,N_20933,N_20153);
nor U22381 (N_22381,N_19078,N_21729);
nor U22382 (N_22382,N_20954,N_21328);
nor U22383 (N_22383,N_20833,N_20752);
or U22384 (N_22384,N_20283,N_21546);
and U22385 (N_22385,N_21379,N_19663);
nand U22386 (N_22386,N_20128,N_18831);
or U22387 (N_22387,N_18839,N_21012);
nor U22388 (N_22388,N_21708,N_19545);
nor U22389 (N_22389,N_20557,N_21190);
nand U22390 (N_22390,N_20406,N_20219);
or U22391 (N_22391,N_20923,N_19241);
and U22392 (N_22392,N_19882,N_21039);
and U22393 (N_22393,N_21053,N_19321);
xor U22394 (N_22394,N_20246,N_21277);
and U22395 (N_22395,N_20244,N_20957);
nor U22396 (N_22396,N_20272,N_21702);
xor U22397 (N_22397,N_21828,N_20517);
nand U22398 (N_22398,N_18781,N_20730);
or U22399 (N_22399,N_20007,N_18973);
nand U22400 (N_22400,N_19850,N_20256);
xor U22401 (N_22401,N_20894,N_20278);
nand U22402 (N_22402,N_20854,N_18846);
nor U22403 (N_22403,N_21872,N_21115);
nand U22404 (N_22404,N_19465,N_19786);
or U22405 (N_22405,N_19304,N_19281);
or U22406 (N_22406,N_21441,N_21011);
xnor U22407 (N_22407,N_21458,N_20050);
xnor U22408 (N_22408,N_19034,N_18964);
or U22409 (N_22409,N_20676,N_20631);
or U22410 (N_22410,N_19373,N_21790);
or U22411 (N_22411,N_19504,N_19334);
or U22412 (N_22412,N_19267,N_21470);
xnor U22413 (N_22413,N_18849,N_19327);
and U22414 (N_22414,N_19090,N_20656);
nor U22415 (N_22415,N_21285,N_21315);
xnor U22416 (N_22416,N_21131,N_21679);
nand U22417 (N_22417,N_21805,N_21498);
xor U22418 (N_22418,N_19600,N_19588);
or U22419 (N_22419,N_19672,N_21242);
and U22420 (N_22420,N_21647,N_21666);
nand U22421 (N_22421,N_19828,N_19043);
nand U22422 (N_22422,N_20821,N_19162);
nor U22423 (N_22423,N_19030,N_19804);
nor U22424 (N_22424,N_21570,N_18750);
xor U22425 (N_22425,N_19372,N_21128);
xor U22426 (N_22426,N_19570,N_18809);
nor U22427 (N_22427,N_21278,N_21074);
nor U22428 (N_22428,N_20643,N_19529);
xor U22429 (N_22429,N_20599,N_20531);
and U22430 (N_22430,N_18940,N_21809);
nand U22431 (N_22431,N_19113,N_19395);
nor U22432 (N_22432,N_18966,N_20425);
nand U22433 (N_22433,N_20732,N_18902);
nor U22434 (N_22434,N_19279,N_20662);
and U22435 (N_22435,N_21372,N_21477);
nand U22436 (N_22436,N_19605,N_18767);
nor U22437 (N_22437,N_21377,N_20447);
xor U22438 (N_22438,N_21471,N_19480);
xor U22439 (N_22439,N_21747,N_19266);
nor U22440 (N_22440,N_21018,N_20401);
xor U22441 (N_22441,N_21873,N_19201);
xor U22442 (N_22442,N_21726,N_20650);
or U22443 (N_22443,N_19781,N_21050);
nand U22444 (N_22444,N_21013,N_19312);
xnor U22445 (N_22445,N_19416,N_21842);
nor U22446 (N_22446,N_20626,N_21438);
xnor U22447 (N_22447,N_21149,N_21146);
nor U22448 (N_22448,N_19264,N_20817);
nor U22449 (N_22449,N_19357,N_20093);
or U22450 (N_22450,N_21688,N_20432);
xor U22451 (N_22451,N_19576,N_21449);
and U22452 (N_22452,N_20548,N_19006);
nor U22453 (N_22453,N_19618,N_19581);
or U22454 (N_22454,N_21207,N_18907);
nor U22455 (N_22455,N_20796,N_20440);
nor U22456 (N_22456,N_21314,N_18783);
nand U22457 (N_22457,N_18892,N_19349);
nand U22458 (N_22458,N_21620,N_19183);
and U22459 (N_22459,N_20736,N_19690);
nor U22460 (N_22460,N_21384,N_19064);
xnor U22461 (N_22461,N_21357,N_20974);
or U22462 (N_22462,N_20877,N_19898);
and U22463 (N_22463,N_20589,N_19813);
or U22464 (N_22464,N_21634,N_20608);
and U22465 (N_22465,N_19460,N_19411);
nor U22466 (N_22466,N_21615,N_20916);
nor U22467 (N_22467,N_20135,N_21478);
or U22468 (N_22468,N_21365,N_19474);
or U22469 (N_22469,N_21331,N_21606);
or U22470 (N_22470,N_21622,N_19033);
and U22471 (N_22471,N_18769,N_21736);
or U22472 (N_22472,N_20040,N_19008);
nand U22473 (N_22473,N_20638,N_21673);
xor U22474 (N_22474,N_20657,N_19341);
and U22475 (N_22475,N_21738,N_21299);
xor U22476 (N_22476,N_21387,N_20262);
xor U22477 (N_22477,N_19722,N_20710);
or U22478 (N_22478,N_21617,N_21041);
xnor U22479 (N_22479,N_21554,N_20890);
nand U22480 (N_22480,N_18896,N_20937);
nor U22481 (N_22481,N_20798,N_19035);
nor U22482 (N_22482,N_21151,N_18982);
xnor U22483 (N_22483,N_19139,N_21680);
and U22484 (N_22484,N_20766,N_20896);
xnor U22485 (N_22485,N_20675,N_18981);
nor U22486 (N_22486,N_20700,N_20030);
and U22487 (N_22487,N_19218,N_21569);
nor U22488 (N_22488,N_21051,N_19709);
nand U22489 (N_22489,N_21301,N_20277);
nand U22490 (N_22490,N_18817,N_21043);
xnor U22491 (N_22491,N_20026,N_20195);
and U22492 (N_22492,N_21681,N_18922);
or U22493 (N_22493,N_19648,N_21815);
nor U22494 (N_22494,N_21695,N_20306);
xor U22495 (N_22495,N_20455,N_19764);
or U22496 (N_22496,N_21038,N_20718);
nand U22497 (N_22497,N_21210,N_19462);
nor U22498 (N_22498,N_19351,N_21060);
and U22499 (N_22499,N_20371,N_18946);
nand U22500 (N_22500,N_20978,N_20799);
nand U22501 (N_22501,N_19976,N_19802);
and U22502 (N_22502,N_20903,N_20872);
xnor U22503 (N_22503,N_20831,N_20255);
nand U22504 (N_22504,N_19740,N_19661);
nand U22505 (N_22505,N_19869,N_21817);
xor U22506 (N_22506,N_20504,N_20393);
xor U22507 (N_22507,N_18984,N_20321);
nand U22508 (N_22508,N_20911,N_19541);
nand U22509 (N_22509,N_21771,N_20750);
nor U22510 (N_22510,N_20492,N_20500);
or U22511 (N_22511,N_21567,N_20178);
nor U22512 (N_22512,N_19066,N_18934);
nor U22513 (N_22513,N_21204,N_21389);
xnor U22514 (N_22514,N_18878,N_21433);
nor U22515 (N_22515,N_20563,N_21671);
xnor U22516 (N_22516,N_19912,N_21386);
nand U22517 (N_22517,N_19048,N_19283);
nand U22518 (N_22518,N_19356,N_21580);
nor U22519 (N_22519,N_19453,N_19310);
nand U22520 (N_22520,N_18888,N_21841);
and U22521 (N_22521,N_20125,N_19909);
nor U22522 (N_22522,N_20015,N_20140);
nor U22523 (N_22523,N_21795,N_19566);
xor U22524 (N_22524,N_21116,N_20767);
nand U22525 (N_22525,N_20545,N_18976);
and U22526 (N_22526,N_21552,N_20363);
or U22527 (N_22527,N_19805,N_18897);
xor U22528 (N_22528,N_21120,N_20327);
nand U22529 (N_22529,N_19447,N_19059);
nand U22530 (N_22530,N_20473,N_20095);
nand U22531 (N_22531,N_20972,N_19494);
nor U22532 (N_22532,N_19755,N_20567);
nor U22533 (N_22533,N_20979,N_20909);
xnor U22534 (N_22534,N_19744,N_20721);
xor U22535 (N_22535,N_19499,N_21764);
xor U22536 (N_22536,N_21255,N_20588);
nor U22537 (N_22537,N_21603,N_19714);
xor U22538 (N_22538,N_20822,N_18800);
xor U22539 (N_22539,N_20642,N_20025);
nor U22540 (N_22540,N_19093,N_19587);
xor U22541 (N_22541,N_19798,N_20538);
and U22542 (N_22542,N_21066,N_20975);
or U22543 (N_22543,N_18886,N_19784);
nor U22544 (N_22544,N_21781,N_20172);
xnor U22545 (N_22545,N_20158,N_19069);
xor U22546 (N_22546,N_21499,N_19236);
and U22547 (N_22547,N_19787,N_21761);
and U22548 (N_22548,N_19359,N_18953);
and U22549 (N_22549,N_18766,N_20032);
nor U22550 (N_22550,N_20742,N_19057);
xor U22551 (N_22551,N_20090,N_20913);
nor U22552 (N_22552,N_20825,N_18930);
nor U22553 (N_22553,N_21112,N_20924);
nand U22554 (N_22554,N_21670,N_20416);
or U22555 (N_22555,N_19214,N_20049);
or U22556 (N_22556,N_21716,N_19314);
or U22557 (N_22557,N_20494,N_19564);
nand U22558 (N_22558,N_21002,N_20714);
xnor U22559 (N_22559,N_20489,N_21669);
xnor U22560 (N_22560,N_20762,N_20335);
nor U22561 (N_22561,N_21523,N_19263);
and U22562 (N_22562,N_21653,N_19268);
and U22563 (N_22563,N_19772,N_20976);
and U22564 (N_22564,N_19929,N_19222);
nand U22565 (N_22565,N_21859,N_21189);
or U22566 (N_22566,N_18890,N_20468);
or U22567 (N_22567,N_21416,N_19067);
nor U22568 (N_22568,N_20420,N_21437);
nor U22569 (N_22569,N_19278,N_19811);
and U22570 (N_22570,N_21537,N_19629);
nor U22571 (N_22571,N_19013,N_21339);
or U22572 (N_22572,N_21229,N_19999);
or U22573 (N_22573,N_20856,N_18866);
and U22574 (N_22574,N_20052,N_20313);
nand U22575 (N_22575,N_19224,N_19433);
xnor U22576 (N_22576,N_18841,N_19518);
and U22577 (N_22577,N_21407,N_19191);
nand U22578 (N_22578,N_19675,N_19488);
nor U22579 (N_22579,N_21162,N_21760);
and U22580 (N_22580,N_20204,N_21662);
nand U22581 (N_22581,N_21607,N_19854);
or U22582 (N_22582,N_20990,N_19366);
nand U22583 (N_22583,N_21319,N_19434);
or U22584 (N_22584,N_19132,N_21590);
xor U22585 (N_22585,N_20216,N_19326);
xor U22586 (N_22586,N_21461,N_18962);
or U22587 (N_22587,N_19445,N_21348);
nand U22588 (N_22588,N_19486,N_21701);
nor U22589 (N_22589,N_19240,N_21770);
and U22590 (N_22590,N_19961,N_21650);
xnor U22591 (N_22591,N_18915,N_21823);
nor U22592 (N_22592,N_19993,N_20122);
xnor U22593 (N_22593,N_21026,N_20481);
or U22594 (N_22594,N_21636,N_19932);
or U22595 (N_22595,N_21519,N_20367);
or U22596 (N_22596,N_19338,N_20558);
nand U22597 (N_22597,N_18978,N_20887);
and U22598 (N_22598,N_20828,N_19471);
nor U22599 (N_22599,N_21451,N_21347);
or U22600 (N_22600,N_19026,N_19638);
and U22601 (N_22601,N_21782,N_21633);
and U22602 (N_22602,N_21417,N_20514);
xor U22603 (N_22603,N_21807,N_20704);
and U22604 (N_22604,N_19801,N_20981);
or U22605 (N_22605,N_21798,N_19446);
and U22606 (N_22606,N_20086,N_20847);
nand U22607 (N_22607,N_21739,N_20587);
xnor U22608 (N_22608,N_18794,N_20399);
nand U22609 (N_22609,N_18884,N_19062);
and U22610 (N_22610,N_21874,N_20051);
nand U22611 (N_22611,N_21295,N_18960);
and U22612 (N_22612,N_18845,N_20372);
and U22613 (N_22613,N_18753,N_20830);
nor U22614 (N_22614,N_20715,N_20235);
nor U22615 (N_22615,N_21307,N_20795);
or U22616 (N_22616,N_19290,N_20127);
and U22617 (N_22617,N_20054,N_18807);
and U22618 (N_22618,N_20129,N_20719);
and U22619 (N_22619,N_21312,N_20597);
xnor U22620 (N_22620,N_20170,N_20451);
xor U22621 (N_22621,N_20320,N_21313);
xnor U22622 (N_22622,N_19928,N_21237);
and U22623 (N_22623,N_19902,N_20740);
and U22624 (N_22624,N_18906,N_21247);
xor U22625 (N_22625,N_20835,N_21578);
xor U22626 (N_22626,N_20991,N_19219);
nand U22627 (N_22627,N_19561,N_21224);
nor U22628 (N_22628,N_21245,N_21720);
nand U22629 (N_22629,N_21395,N_20527);
nor U22630 (N_22630,N_19313,N_19650);
nor U22631 (N_22631,N_19621,N_21468);
xnor U22632 (N_22632,N_19185,N_19501);
xnor U22633 (N_22633,N_19762,N_21177);
or U22634 (N_22634,N_20120,N_21692);
nand U22635 (N_22635,N_20834,N_19128);
nand U22636 (N_22636,N_20660,N_20932);
and U22637 (N_22637,N_20646,N_20512);
nand U22638 (N_22638,N_20585,N_20691);
nand U22639 (N_22639,N_19215,N_19020);
and U22640 (N_22640,N_20304,N_20763);
and U22641 (N_22641,N_18828,N_20709);
nand U22642 (N_22642,N_21272,N_19952);
xnor U22643 (N_22643,N_21483,N_18777);
and U22644 (N_22644,N_20094,N_20737);
nand U22645 (N_22645,N_21196,N_20329);
nand U22646 (N_22646,N_19164,N_19849);
nand U22647 (N_22647,N_19693,N_21643);
nand U22648 (N_22648,N_21418,N_19715);
nand U22649 (N_22649,N_20820,N_19459);
or U22650 (N_22650,N_20149,N_21856);
nand U22651 (N_22651,N_19768,N_20651);
and U22652 (N_22652,N_20503,N_21484);
nand U22653 (N_22653,N_21664,N_19526);
nor U22654 (N_22654,N_19521,N_20701);
xor U22655 (N_22655,N_18926,N_20717);
nor U22656 (N_22656,N_20373,N_19135);
and U22657 (N_22657,N_19187,N_19864);
or U22658 (N_22658,N_21399,N_21015);
nor U22659 (N_22659,N_19945,N_21127);
nand U22660 (N_22660,N_21557,N_21133);
and U22661 (N_22661,N_21324,N_21150);
or U22662 (N_22662,N_20619,N_21054);
nor U22663 (N_22663,N_20565,N_21691);
nor U22664 (N_22664,N_18816,N_20769);
or U22665 (N_22665,N_20874,N_20502);
xor U22666 (N_22666,N_19025,N_19904);
nand U22667 (N_22667,N_20860,N_19376);
nand U22668 (N_22668,N_21014,N_20749);
and U22669 (N_22669,N_20922,N_21413);
xnor U22670 (N_22670,N_20947,N_20540);
and U22671 (N_22671,N_19930,N_18912);
and U22672 (N_22672,N_20340,N_20682);
nor U22673 (N_22673,N_21728,N_20409);
xnor U22674 (N_22674,N_20888,N_19037);
nor U22675 (N_22675,N_19133,N_19428);
nand U22676 (N_22676,N_19157,N_20036);
or U22677 (N_22677,N_20354,N_19245);
xnor U22678 (N_22678,N_19803,N_18773);
nand U22679 (N_22679,N_20511,N_21540);
nor U22680 (N_22680,N_20469,N_19440);
or U22681 (N_22681,N_20209,N_20297);
nand U22682 (N_22682,N_19014,N_20863);
and U22683 (N_22683,N_19775,N_21317);
nor U22684 (N_22684,N_21084,N_21829);
nand U22685 (N_22685,N_20144,N_19980);
nand U22686 (N_22686,N_18885,N_19052);
and U22687 (N_22687,N_21030,N_21235);
nand U22688 (N_22688,N_21857,N_20057);
xnor U22689 (N_22689,N_20276,N_19298);
nand U22690 (N_22690,N_20325,N_20448);
nand U22691 (N_22691,N_21436,N_19844);
xor U22692 (N_22692,N_19137,N_21521);
nor U22693 (N_22693,N_20672,N_18975);
or U22694 (N_22694,N_19046,N_21547);
xor U22695 (N_22695,N_19823,N_19747);
nor U22696 (N_22696,N_21137,N_19594);
or U22697 (N_22697,N_21169,N_19777);
xnor U22698 (N_22698,N_20005,N_19586);
xnor U22699 (N_22699,N_19168,N_21102);
nand U22700 (N_22700,N_21250,N_19437);
xor U22701 (N_22701,N_18980,N_21456);
and U22702 (N_22702,N_21731,N_20053);
xor U22703 (N_22703,N_21496,N_21457);
xnor U22704 (N_22704,N_19578,N_21028);
nand U22705 (N_22705,N_20994,N_19007);
xor U22706 (N_22706,N_19087,N_20781);
xnor U22707 (N_22707,N_21871,N_19745);
and U22708 (N_22708,N_20945,N_20837);
xnor U22709 (N_22709,N_19355,N_19250);
nor U22710 (N_22710,N_21444,N_21100);
xnor U22711 (N_22711,N_20390,N_20731);
or U22712 (N_22712,N_19028,N_18792);
and U22713 (N_22713,N_18779,N_19839);
or U22714 (N_22714,N_19011,N_21310);
xnor U22715 (N_22715,N_21733,N_18812);
xnor U22716 (N_22716,N_20602,N_19819);
xor U22717 (N_22717,N_21056,N_18947);
nor U22718 (N_22718,N_20251,N_18889);
and U22719 (N_22719,N_21423,N_20892);
nor U22720 (N_22720,N_21838,N_20477);
nand U22721 (N_22721,N_20805,N_18820);
nand U22722 (N_22722,N_20220,N_21292);
or U22723 (N_22723,N_20948,N_18921);
nor U22724 (N_22724,N_20437,N_21485);
nor U22725 (N_22725,N_21544,N_21667);
nor U22726 (N_22726,N_19563,N_21715);
xor U22727 (N_22727,N_19889,N_21534);
or U22728 (N_22728,N_20434,N_21434);
xnor U22729 (N_22729,N_20068,N_20177);
and U22730 (N_22730,N_18928,N_20392);
xnor U22731 (N_22731,N_19197,N_19863);
xnor U22732 (N_22732,N_19107,N_19933);
nor U22733 (N_22733,N_20811,N_21263);
nand U22734 (N_22734,N_19760,N_20357);
xnor U22735 (N_22735,N_20339,N_19708);
nand U22736 (N_22736,N_18879,N_20632);
and U22737 (N_22737,N_21543,N_20157);
xnor U22738 (N_22738,N_21754,N_18996);
xnor U22739 (N_22739,N_21411,N_18818);
nor U22740 (N_22740,N_21572,N_20711);
nor U22741 (N_22741,N_21722,N_19975);
xor U22742 (N_22742,N_18832,N_20452);
nor U22743 (N_22743,N_21023,N_21683);
nor U22744 (N_22744,N_19757,N_19619);
or U22745 (N_22745,N_21284,N_20319);
or U22746 (N_22746,N_21267,N_19016);
or U22747 (N_22747,N_19193,N_19186);
and U22748 (N_22748,N_19237,N_21168);
nand U22749 (N_22749,N_21748,N_20279);
nand U22750 (N_22750,N_20449,N_19874);
nand U22751 (N_22751,N_20941,N_20739);
nor U22752 (N_22752,N_21424,N_20046);
and U22753 (N_22753,N_19217,N_19539);
and U22754 (N_22754,N_19109,N_20400);
or U22755 (N_22755,N_19956,N_21361);
or U22756 (N_22756,N_21678,N_20472);
or U22757 (N_22757,N_21529,N_21206);
xnor U22758 (N_22758,N_19276,N_20289);
xor U22759 (N_22759,N_20695,N_19206);
nand U22760 (N_22760,N_20765,N_21370);
or U22761 (N_22761,N_20761,N_21305);
xor U22762 (N_22762,N_19337,N_20653);
xnor U22763 (N_22763,N_20944,N_19086);
or U22764 (N_22764,N_20136,N_21465);
nor U22765 (N_22765,N_21271,N_20560);
or U22766 (N_22766,N_21822,N_19442);
nor U22767 (N_22767,N_20853,N_21613);
xor U22768 (N_22768,N_21231,N_20755);
or U22769 (N_22769,N_19865,N_20351);
nand U22770 (N_22770,N_21072,N_19165);
nor U22771 (N_22771,N_20735,N_19178);
nand U22772 (N_22772,N_20987,N_21360);
or U22773 (N_22773,N_19449,N_18942);
and U22774 (N_22774,N_20047,N_19957);
and U22775 (N_22775,N_19822,N_21215);
nand U22776 (N_22776,N_20189,N_21674);
or U22777 (N_22777,N_21801,N_19381);
nand U22778 (N_22778,N_20138,N_20683);
and U22779 (N_22779,N_20012,N_19225);
nand U22780 (N_22780,N_18754,N_19418);
and U22781 (N_22781,N_21337,N_20346);
nor U22782 (N_22782,N_19166,N_20884);
or U22783 (N_22783,N_20499,N_18827);
or U22784 (N_22784,N_19894,N_19223);
xor U22785 (N_22785,N_20883,N_18882);
nand U22786 (N_22786,N_21351,N_20341);
and U22787 (N_22787,N_20185,N_19104);
and U22788 (N_22788,N_21118,N_21221);
or U22789 (N_22789,N_21410,N_20159);
nand U22790 (N_22790,N_21153,N_21109);
xnor U22791 (N_22791,N_21584,N_21641);
nor U22792 (N_22792,N_21515,N_21460);
nand U22793 (N_22793,N_21165,N_19572);
xnor U22794 (N_22794,N_18933,N_21717);
xor U22795 (N_22795,N_19169,N_20439);
or U22796 (N_22796,N_19765,N_19422);
nand U22797 (N_22797,N_19971,N_20200);
and U22798 (N_22798,N_21612,N_19589);
and U22799 (N_22799,N_21618,N_19426);
and U22800 (N_22800,N_20655,N_19664);
nand U22801 (N_22801,N_19500,N_19926);
nand U22802 (N_22802,N_19525,N_18830);
xor U22803 (N_22803,N_19915,N_21230);
or U22804 (N_22804,N_20697,N_19942);
xnor U22805 (N_22805,N_19431,N_21254);
nor U22806 (N_22806,N_19348,N_20006);
nand U22807 (N_22807,N_19487,N_20314);
xor U22808 (N_22808,N_20027,N_20956);
xnor U22809 (N_22809,N_21094,N_20550);
and U22810 (N_22810,N_20379,N_21700);
and U22811 (N_22811,N_20493,N_21356);
xnor U22812 (N_22812,N_19848,N_20305);
or U22813 (N_22813,N_20712,N_20342);
nand U22814 (N_22814,N_20460,N_20733);
xor U22815 (N_22815,N_20713,N_21750);
xnor U22816 (N_22816,N_20880,N_21658);
and U22817 (N_22817,N_19973,N_20308);
or U22818 (N_22818,N_18877,N_20174);
xnor U22819 (N_22819,N_19361,N_18822);
nor U22820 (N_22820,N_18798,N_18909);
nand U22821 (N_22821,N_20059,N_21711);
or U22822 (N_22822,N_20858,N_20640);
and U22823 (N_22823,N_21765,N_21152);
and U22824 (N_22824,N_20398,N_19773);
nor U22825 (N_22825,N_18919,N_21753);
nand U22826 (N_22826,N_18838,N_19410);
and U22827 (N_22827,N_18883,N_20901);
and U22828 (N_22828,N_21113,N_19391);
or U22829 (N_22829,N_21318,N_19092);
nand U22830 (N_22830,N_18756,N_18968);
nand U22831 (N_22831,N_20871,N_19683);
or U22832 (N_22832,N_20428,N_20429);
and U22833 (N_22833,N_21821,N_18813);
or U22834 (N_22834,N_20555,N_19089);
and U22835 (N_22835,N_19659,N_21769);
or U22836 (N_22836,N_19274,N_21599);
nor U22837 (N_22837,N_20332,N_20166);
or U22838 (N_22838,N_21522,N_19788);
or U22839 (N_22839,N_18764,N_21511);
nor U22840 (N_22840,N_19584,N_20442);
nand U22841 (N_22841,N_20573,N_20815);
and U22842 (N_22842,N_19927,N_19116);
nor U22843 (N_22843,N_19343,N_20580);
and U22844 (N_22844,N_21369,N_20862);
or U22845 (N_22845,N_19860,N_21035);
nor U22846 (N_22846,N_19045,N_20205);
and U22847 (N_22847,N_20160,N_19401);
xnor U22848 (N_22848,N_19238,N_20191);
xnor U22849 (N_22849,N_20832,N_19041);
nand U22850 (N_22850,N_20859,N_19194);
and U22851 (N_22851,N_19681,N_19138);
and U22852 (N_22852,N_20087,N_20839);
nor U22853 (N_22853,N_21345,N_19551);
nor U22854 (N_22854,N_19002,N_20899);
xnor U22855 (N_22855,N_21343,N_20060);
nand U22856 (N_22856,N_21762,N_21217);
nor U22857 (N_22857,N_20529,N_19136);
nor U22858 (N_22858,N_20988,N_19721);
and U22859 (N_22859,N_19610,N_21174);
nand U22860 (N_22860,N_21090,N_21027);
and U22861 (N_22861,N_21202,N_21869);
nand U22862 (N_22862,N_21791,N_20150);
or U22863 (N_22863,N_20303,N_20081);
xnor U22864 (N_22864,N_19330,N_20964);
and U22865 (N_22865,N_19657,N_20318);
xnor U22866 (N_22866,N_20554,N_20441);
nand U22867 (N_22867,N_20154,N_19495);
nor U22868 (N_22868,N_21046,N_21657);
nor U22869 (N_22869,N_18799,N_19922);
nand U22870 (N_22870,N_18911,N_19211);
or U22871 (N_22871,N_20161,N_18863);
nor U22872 (N_22872,N_21258,N_20261);
xor U22873 (N_22873,N_20915,N_21826);
and U22874 (N_22874,N_20039,N_19939);
or U22875 (N_22875,N_21212,N_19622);
and U22876 (N_22876,N_20431,N_21550);
and U22877 (N_22877,N_20298,N_20179);
nor U22878 (N_22878,N_19461,N_19533);
nand U22879 (N_22879,N_19095,N_19511);
nand U22880 (N_22880,N_21767,N_20873);
nor U22881 (N_22881,N_19363,N_20702);
and U22882 (N_22882,N_20231,N_19302);
xor U22883 (N_22883,N_19344,N_19394);
nand U22884 (N_22884,N_20520,N_20115);
xor U22885 (N_22885,N_20569,N_20263);
nor U22886 (N_22886,N_21644,N_19994);
xor U22887 (N_22887,N_19144,N_20423);
or U22888 (N_22888,N_20743,N_21099);
xnor U22889 (N_22889,N_19231,N_21694);
nor U22890 (N_22890,N_21507,N_21261);
nor U22891 (N_22891,N_20112,N_21282);
nor U22892 (N_22892,N_21549,N_19436);
nand U22893 (N_22893,N_18929,N_20295);
xnor U22894 (N_22894,N_20869,N_21342);
or U22895 (N_22895,N_21665,N_21677);
or U22896 (N_22896,N_21699,N_19342);
xnor U22897 (N_22897,N_20591,N_18891);
and U22898 (N_22898,N_21175,N_21306);
or U22899 (N_22899,N_21774,N_19317);
xnor U22900 (N_22900,N_19210,N_19280);
and U22901 (N_22901,N_21561,N_21080);
or U22902 (N_22902,N_19905,N_20197);
or U22903 (N_22903,N_20939,N_18758);
nand U22904 (N_22904,N_20476,N_18864);
xnor U22905 (N_22905,N_19272,N_21684);
nand U22906 (N_22906,N_21453,N_21327);
or U22907 (N_22907,N_20072,N_19134);
nand U22908 (N_22908,N_19402,N_21201);
or U22909 (N_22909,N_19514,N_20110);
nand U22910 (N_22910,N_20198,N_19537);
or U22911 (N_22911,N_20422,N_20215);
nor U22912 (N_22912,N_20243,N_18806);
nand U22913 (N_22913,N_21480,N_19256);
nand U22914 (N_22914,N_21021,N_20720);
xor U22915 (N_22915,N_21276,N_19024);
nand U22916 (N_22916,N_19550,N_19887);
nor U22917 (N_22917,N_18770,N_19964);
nand U22918 (N_22918,N_19060,N_19800);
nor U22919 (N_22919,N_20033,N_21428);
nor U22920 (N_22920,N_19339,N_21070);
nor U22921 (N_22921,N_20323,N_20612);
and U22922 (N_22922,N_18979,N_20966);
nand U22923 (N_22923,N_19156,N_20848);
nor U22924 (N_22924,N_20907,N_21628);
nand U22925 (N_22925,N_21353,N_21476);
xor U22926 (N_22926,N_21450,N_21559);
xor U22927 (N_22927,N_20348,N_20958);
and U22928 (N_22928,N_20326,N_21594);
xor U22929 (N_22929,N_20227,N_19938);
or U22930 (N_22930,N_18821,N_21672);
xor U22931 (N_22931,N_21087,N_18932);
nand U22932 (N_22932,N_19080,N_21608);
xnor U22933 (N_22933,N_20934,N_19018);
and U22934 (N_22934,N_19634,N_20867);
nand U22935 (N_22935,N_19022,N_21778);
nor U22936 (N_22936,N_19734,N_19923);
nand U22937 (N_22937,N_20726,N_20630);
xor U22938 (N_22938,N_18963,N_21024);
nand U22939 (N_22939,N_21655,N_20331);
nor U22940 (N_22940,N_21172,N_19098);
xor U22941 (N_22941,N_21294,N_19741);
or U22942 (N_22942,N_19331,N_19603);
and U22943 (N_22943,N_19258,N_19216);
xor U22944 (N_22944,N_21542,N_21867);
nor U22945 (N_22945,N_20290,N_21059);
and U22946 (N_22946,N_20067,N_19386);
nor U22947 (N_22947,N_19988,N_20722);
xor U22948 (N_22948,N_20111,N_20870);
xnor U22949 (N_22949,N_20793,N_21514);
nand U22950 (N_22950,N_18755,N_19145);
xnor U22951 (N_22951,N_21040,N_21415);
nor U22952 (N_22952,N_20106,N_19094);
or U22953 (N_22953,N_19625,N_21598);
or U22954 (N_22954,N_19209,N_19731);
xnor U22955 (N_22955,N_21827,N_19345);
or U22956 (N_22956,N_20562,N_20673);
or U22957 (N_22957,N_21836,N_20337);
and U22958 (N_22958,N_18811,N_19856);
xor U22959 (N_22959,N_19776,N_20849);
xor U22960 (N_22960,N_21682,N_18837);
or U22961 (N_22961,N_21581,N_19901);
nand U22962 (N_22962,N_20776,N_20224);
or U22963 (N_22963,N_21712,N_20738);
nor U22964 (N_22964,N_19895,N_19375);
nor U22965 (N_22965,N_20264,N_19637);
nand U22966 (N_22966,N_20023,N_19071);
nor U22967 (N_22967,N_20577,N_19888);
and U22968 (N_22968,N_21032,N_21685);
nand U22969 (N_22969,N_19793,N_20435);
nor U22970 (N_22970,N_20570,N_21300);
and U22971 (N_22971,N_19199,N_19674);
xor U22972 (N_22972,N_19481,N_21614);
nor U22973 (N_22973,N_20627,N_19516);
nand U22974 (N_22974,N_20366,N_18957);
xnor U22975 (N_22975,N_19143,N_21316);
or U22976 (N_22976,N_19364,N_18871);
nor U22977 (N_22977,N_20201,N_20024);
nand U22978 (N_22978,N_20182,N_20985);
or U22979 (N_22979,N_21246,N_21730);
or U22980 (N_22980,N_19989,N_19261);
nor U22981 (N_22981,N_20900,N_20043);
nand U22982 (N_22982,N_20171,N_20038);
xor U22983 (N_22983,N_20850,N_20287);
nand U22984 (N_22984,N_21068,N_19884);
nor U22985 (N_22985,N_21354,N_19198);
or U22986 (N_22986,N_21775,N_19692);
and U22987 (N_22987,N_19119,N_19177);
xnor U22988 (N_22988,N_19662,N_18803);
nor U22989 (N_22989,N_20508,N_21755);
or U22990 (N_22990,N_21868,N_21103);
nand U22991 (N_22991,N_19825,N_19181);
and U22992 (N_22992,N_21154,N_21573);
xor U22993 (N_22993,N_21243,N_20242);
or U22994 (N_22994,N_18970,N_21844);
or U22995 (N_22995,N_21157,N_20433);
nor U22996 (N_22996,N_19678,N_19354);
xor U22997 (N_22997,N_19562,N_21863);
xnor U22998 (N_22998,N_19774,N_19615);
xnor U22999 (N_22999,N_20952,N_19958);
or U23000 (N_23000,N_20490,N_18937);
or U23001 (N_23001,N_21185,N_19249);
nand U23002 (N_23002,N_20532,N_19328);
xor U23003 (N_23003,N_20851,N_18824);
and U23004 (N_23004,N_20857,N_20165);
xor U23005 (N_23005,N_20188,N_21454);
or U23006 (N_23006,N_19872,N_20237);
nor U23007 (N_23007,N_21076,N_19472);
nand U23008 (N_23008,N_19510,N_20056);
nand U23009 (N_23009,N_18993,N_19689);
or U23010 (N_23010,N_18804,N_20644);
xor U23011 (N_23011,N_19816,N_20989);
nand U23012 (N_23012,N_19470,N_20584);
nand U23013 (N_23013,N_19542,N_21036);
nand U23014 (N_23014,N_20895,N_21752);
nor U23015 (N_23015,N_18847,N_20019);
and U23016 (N_23016,N_19623,N_21742);
nor U23017 (N_23017,N_20167,N_19491);
xnor U23018 (N_23018,N_19148,N_21122);
and U23019 (N_23019,N_21591,N_19100);
and U23020 (N_23020,N_20230,N_20391);
and U23021 (N_23021,N_19163,N_20045);
xnor U23022 (N_23022,N_20016,N_21497);
or U23023 (N_23023,N_20018,N_19724);
nor U23024 (N_23024,N_21601,N_18952);
nor U23025 (N_23025,N_19742,N_20352);
xor U23026 (N_23026,N_19585,N_21020);
and U23027 (N_23027,N_21065,N_18969);
and U23028 (N_23028,N_20840,N_19649);
nand U23029 (N_23029,N_20311,N_20104);
and U23030 (N_23030,N_20693,N_20668);
nor U23031 (N_23031,N_21531,N_21134);
nand U23032 (N_23032,N_19489,N_20785);
or U23033 (N_23033,N_19966,N_20083);
or U23034 (N_23034,N_19246,N_20280);
xnor U23035 (N_23035,N_19001,N_19797);
xnor U23036 (N_23036,N_20438,N_21439);
nand U23037 (N_23037,N_19085,N_20377);
and U23038 (N_23038,N_20212,N_20970);
and U23039 (N_23039,N_20575,N_19485);
or U23040 (N_23040,N_21575,N_19809);
and U23041 (N_23041,N_21253,N_21780);
xor U23042 (N_23042,N_21556,N_20322);
nand U23043 (N_23043,N_19962,N_20364);
xor U23044 (N_23044,N_19360,N_19333);
nand U23045 (N_23045,N_19441,N_21466);
nor U23046 (N_23046,N_19527,N_19273);
xnor U23047 (N_23047,N_21687,N_20841);
and U23048 (N_23048,N_20919,N_21238);
nand U23049 (N_23049,N_18950,N_19992);
nor U23050 (N_23050,N_21719,N_19227);
xor U23051 (N_23051,N_21489,N_21843);
xnor U23052 (N_23052,N_19038,N_21281);
nand U23053 (N_23053,N_20465,N_20353);
xnor U23054 (N_23054,N_20663,N_20998);
and U23055 (N_23055,N_19611,N_19155);
or U23056 (N_23056,N_20961,N_19967);
nor U23057 (N_23057,N_19607,N_19751);
or U23058 (N_23058,N_21430,N_19959);
nor U23059 (N_23059,N_19523,N_20020);
or U23060 (N_23060,N_18972,N_21661);
xor U23061 (N_23061,N_18867,N_21864);
nand U23062 (N_23062,N_19920,N_20089);
nor U23063 (N_23063,N_19170,N_18971);
nor U23064 (N_23064,N_21751,N_18992);
nand U23065 (N_23065,N_19513,N_19732);
xnor U23066 (N_23066,N_20203,N_20621);
nand U23067 (N_23067,N_19254,N_19995);
nor U23068 (N_23068,N_21793,N_20962);
and U23069 (N_23069,N_19896,N_21111);
nand U23070 (N_23070,N_18974,N_20257);
or U23071 (N_23071,N_19834,N_20784);
or U23072 (N_23072,N_20603,N_19105);
xnor U23073 (N_23073,N_20935,N_20519);
xor U23074 (N_23074,N_21368,N_19627);
or U23075 (N_23075,N_18786,N_20528);
nand U23076 (N_23076,N_20424,N_19383);
and U23077 (N_23077,N_19954,N_21442);
nor U23078 (N_23078,N_20661,N_20241);
nor U23079 (N_23079,N_20965,N_19748);
nor U23080 (N_23080,N_21364,N_21063);
or U23081 (N_23081,N_19509,N_20925);
nand U23082 (N_23082,N_20022,N_20596);
nor U23083 (N_23083,N_21330,N_19730);
nor U23084 (N_23084,N_19870,N_19906);
nand U23085 (N_23085,N_21406,N_21148);
and U23086 (N_23086,N_19590,N_19398);
xnor U23087 (N_23087,N_19229,N_20845);
nor U23088 (N_23088,N_19997,N_21409);
nand U23089 (N_23089,N_21520,N_19946);
and U23090 (N_23090,N_21646,N_20126);
or U23091 (N_23091,N_20891,N_19147);
xor U23092 (N_23092,N_21698,N_21602);
or U23093 (N_23093,N_19936,N_19140);
xor U23094 (N_23094,N_21034,N_19536);
xnor U23095 (N_23095,N_20686,N_19780);
and U23096 (N_23096,N_21160,N_19323);
xnor U23097 (N_23097,N_21853,N_21639);
or U23098 (N_23098,N_20375,N_21239);
and U23099 (N_23099,N_18881,N_21587);
nand U23100 (N_23100,N_20996,N_19660);
or U23101 (N_23101,N_20410,N_21244);
nand U23102 (N_23102,N_20427,N_19824);
nand U23103 (N_23103,N_19918,N_20698);
xnor U23104 (N_23104,N_21806,N_20881);
nand U23105 (N_23105,N_19350,N_21081);
nor U23106 (N_23106,N_20474,N_20641);
nand U23107 (N_23107,N_19294,N_19275);
xnor U23108 (N_23108,N_20096,N_21303);
or U23109 (N_23109,N_21117,N_19370);
nand U23110 (N_23110,N_19569,N_19907);
or U23111 (N_23111,N_20463,N_20921);
nand U23112 (N_23112,N_21414,N_19292);
and U23113 (N_23113,N_19247,N_19012);
nand U23114 (N_23114,N_20940,N_20917);
xnor U23115 (N_23115,N_20912,N_19886);
nand U23116 (N_23116,N_20999,N_19439);
or U23117 (N_23117,N_19248,N_21248);
nand U23118 (N_23118,N_21218,N_19892);
or U23119 (N_23119,N_19983,N_18923);
nor U23120 (N_23120,N_19853,N_21635);
nand U23121 (N_23121,N_18860,N_19023);
xnor U23122 (N_23122,N_19547,N_19841);
nor U23123 (N_23123,N_20100,N_21249);
and U23124 (N_23124,N_18775,N_19913);
nor U23125 (N_23125,N_19969,N_21558);
nor U23126 (N_23126,N_19303,N_20010);
xor U23127 (N_23127,N_21789,N_20296);
or U23128 (N_23128,N_18905,N_21192);
nor U23129 (N_23129,N_19652,N_19190);
nor U23130 (N_23130,N_21408,N_19668);
nor U23131 (N_23131,N_20404,N_19503);
nand U23132 (N_23132,N_19916,N_21763);
nand U23133 (N_23133,N_21270,N_20008);
xor U23134 (N_23134,N_20480,N_19175);
nand U23135 (N_23135,N_19230,N_20184);
and U23136 (N_23136,N_21321,N_20688);
xor U23137 (N_23137,N_21629,N_21180);
xor U23138 (N_23138,N_21373,N_21851);
and U23139 (N_23139,N_20522,N_20387);
nor U23140 (N_23140,N_20368,N_20208);
nor U23141 (N_23141,N_18998,N_20240);
nand U23142 (N_23142,N_20678,N_20267);
xor U23143 (N_23143,N_21707,N_20384);
and U23144 (N_23144,N_19639,N_20760);
xor U23145 (N_23145,N_20173,N_21849);
or U23146 (N_23146,N_19725,N_20770);
nor U23147 (N_23147,N_21609,N_19953);
nand U23148 (N_23148,N_21740,N_19497);
nand U23149 (N_23149,N_20777,N_19560);
and U23150 (N_23150,N_20031,N_21088);
nor U23151 (N_23151,N_20708,N_20535);
or U23152 (N_23152,N_18987,N_20647);
xnor U23153 (N_23153,N_18869,N_21710);
and U23154 (N_23154,N_21735,N_19753);
or U23155 (N_23155,N_20955,N_18977);
or U23156 (N_23156,N_21840,N_19778);
nor U23157 (N_23157,N_20413,N_21105);
nor U23158 (N_23158,N_20986,N_19756);
nand U23159 (N_23159,N_20385,N_20403);
xnor U23160 (N_23160,N_20292,N_19602);
nor U23161 (N_23161,N_21156,N_18793);
xnor U23162 (N_23162,N_21425,N_20344);
and U23163 (N_23163,N_21493,N_21199);
or U23164 (N_23164,N_20727,N_21022);
xnor U23165 (N_23165,N_20376,N_19308);
nor U23166 (N_23166,N_19931,N_21445);
and U23167 (N_23167,N_21548,N_19530);
xor U23168 (N_23168,N_20405,N_18805);
and U23169 (N_23169,N_19984,N_19677);
xor U23170 (N_23170,N_21848,N_18784);
nand U23171 (N_23171,N_19968,N_20109);
nand U23172 (N_23172,N_19667,N_19738);
nor U23173 (N_23173,N_20107,N_21338);
nor U23174 (N_23174,N_20624,N_19911);
or U23175 (N_23175,N_19838,N_21562);
nor U23176 (N_23176,N_20347,N_19212);
nor U23177 (N_23177,N_21388,N_18988);
or U23178 (N_23178,N_21309,N_20823);
or U23179 (N_23179,N_19493,N_20041);
nand U23180 (N_23180,N_20281,N_19697);
or U23181 (N_23181,N_19746,N_21145);
and U23182 (N_23182,N_19857,N_19821);
and U23183 (N_23183,N_18840,N_19599);
and U23184 (N_23184,N_21759,N_21797);
nor U23185 (N_23185,N_20362,N_19609);
nand U23186 (N_23186,N_21779,N_21219);
nor U23187 (N_23187,N_19840,N_19101);
nand U23188 (N_23188,N_20537,N_19726);
and U23189 (N_23189,N_20747,N_19318);
or U23190 (N_23190,N_19213,N_18999);
xnor U23191 (N_23191,N_21135,N_19921);
nor U23192 (N_23192,N_20637,N_21311);
xor U23193 (N_23193,N_20309,N_21336);
nor U23194 (N_23194,N_21825,N_20350);
nand U23195 (N_23195,N_19208,N_20618);
or U23196 (N_23196,N_21262,N_19684);
and U23197 (N_23197,N_21585,N_20312);
nor U23198 (N_23198,N_20746,N_20936);
and U23199 (N_23199,N_21178,N_19568);
xnor U23200 (N_23200,N_19111,N_19387);
nor U23201 (N_23201,N_21668,N_21291);
or U23202 (N_23202,N_20792,N_20829);
or U23203 (N_23203,N_20249,N_21092);
or U23204 (N_23204,N_21579,N_21382);
xor U23205 (N_23205,N_21640,N_19406);
xnor U23206 (N_23206,N_20546,N_20374);
nor U23207 (N_23207,N_20791,N_20864);
nor U23208 (N_23208,N_21830,N_19377);
and U23209 (N_23209,N_20097,N_19320);
nand U23210 (N_23210,N_21832,N_20579);
and U23211 (N_23211,N_19405,N_21538);
xor U23212 (N_23212,N_21216,N_21220);
xnor U23213 (N_23213,N_21845,N_20037);
or U23214 (N_23214,N_19727,N_19893);
nand U23215 (N_23215,N_18868,N_19704);
and U23216 (N_23216,N_20946,N_20450);
xnor U23217 (N_23217,N_20168,N_21784);
nand U23218 (N_23218,N_20516,N_19656);
xor U23219 (N_23219,N_21341,N_21846);
or U23220 (N_23220,N_21136,N_18898);
nand U23221 (N_23221,N_20790,N_20092);
or U23222 (N_23222,N_19591,N_19073);
or U23223 (N_23223,N_19019,N_21474);
or U23224 (N_23224,N_19068,N_19047);
nand U23225 (N_23225,N_20077,N_19970);
xnor U23226 (N_23226,N_20408,N_21067);
nand U23227 (N_23227,N_20533,N_18848);
or U23228 (N_23228,N_19977,N_20336);
nor U23229 (N_23229,N_20293,N_21703);
and U23230 (N_23230,N_20905,N_19871);
or U23231 (N_23231,N_20928,N_18927);
nand U23232 (N_23232,N_19031,N_19820);
or U23233 (N_23233,N_20426,N_21085);
nand U23234 (N_23234,N_21721,N_21283);
nand U23235 (N_23235,N_19056,N_21654);
nand U23236 (N_23236,N_21170,N_20248);
or U23237 (N_23237,N_21824,N_19515);
and U23238 (N_23238,N_20724,N_20838);
nor U23239 (N_23239,N_19546,N_19347);
xnor U23240 (N_23240,N_19943,N_20586);
and U23241 (N_23241,N_21431,N_19407);
nand U23242 (N_23242,N_21834,N_20381);
nor U23243 (N_23243,N_20380,N_20412);
xor U23244 (N_23244,N_21714,N_21144);
or U23245 (N_23245,N_18967,N_19583);
and U23246 (N_23246,N_19288,N_20889);
and U23247 (N_23247,N_20786,N_21510);
and U23248 (N_23248,N_19055,N_18870);
nand U23249 (N_23249,N_21479,N_19573);
nor U23250 (N_23250,N_20156,N_19829);
nand U23251 (N_23251,N_20181,N_20953);
xor U23252 (N_23252,N_18856,N_19015);
nand U23253 (N_23253,N_20456,N_20861);
or U23254 (N_23254,N_19082,N_20415);
or U23255 (N_23255,N_20000,N_21536);
and U23256 (N_23256,N_21651,N_19981);
nand U23257 (N_23257,N_21696,N_21031);
xor U23258 (N_23258,N_21288,N_19671);
nor U23259 (N_23259,N_19996,N_21611);
and U23260 (N_23260,N_21488,N_19713);
nor U23261 (N_23261,N_19468,N_20622);
xnor U23262 (N_23262,N_20929,N_20495);
xnor U23263 (N_23263,N_19172,N_18875);
nor U23264 (N_23264,N_20369,N_20358);
and U23265 (N_23265,N_18925,N_21194);
or U23266 (N_23266,N_20813,N_19492);
xnor U23267 (N_23267,N_19123,N_19624);
nor U23268 (N_23268,N_20908,N_19628);
and U23269 (N_23269,N_20078,N_21098);
nor U23270 (N_23270,N_19392,N_19522);
nor U23271 (N_23271,N_20225,N_21078);
nor U23272 (N_23272,N_20705,N_19114);
or U23273 (N_23273,N_19353,N_20294);
and U23274 (N_23274,N_21811,N_20411);
or U23275 (N_23275,N_21553,N_19699);
nand U23276 (N_23276,N_20151,N_20788);
or U23277 (N_23277,N_18985,N_20004);
xor U23278 (N_23278,N_19779,N_19763);
nor U23279 (N_23279,N_20496,N_20258);
and U23280 (N_23280,N_20454,N_19843);
nor U23281 (N_23281,N_19291,N_19420);
nand U23282 (N_23282,N_19117,N_19985);
nor U23283 (N_23283,N_20633,N_19891);
xor U23284 (N_23284,N_20606,N_19425);
xnor U23285 (N_23285,N_19919,N_19039);
nand U23286 (N_23286,N_19072,N_19010);
and U23287 (N_23287,N_19389,N_20483);
nor U23288 (N_23288,N_18989,N_19325);
or U23289 (N_23289,N_19316,N_20634);
nor U23290 (N_23290,N_20021,N_19707);
nor U23291 (N_23291,N_20530,N_21110);
nor U23292 (N_23292,N_20582,N_18789);
xnor U23293 (N_23293,N_20471,N_21610);
and U23294 (N_23294,N_19040,N_20716);
and U23295 (N_23295,N_20370,N_21571);
nor U23296 (N_23296,N_20202,N_20118);
nor U23297 (N_23297,N_20968,N_21044);
xnor U23298 (N_23298,N_20210,N_20771);
and U23299 (N_23299,N_21799,N_19065);
or U23300 (N_23300,N_21394,N_21029);
nor U23301 (N_23301,N_19450,N_20284);
or U23302 (N_23302,N_20218,N_21208);
nand U23303 (N_23303,N_18900,N_19565);
xor U23304 (N_23304,N_21093,N_19432);
and U23305 (N_23305,N_19807,N_21223);
nor U23306 (N_23306,N_19761,N_19944);
or U23307 (N_23307,N_20501,N_21213);
and U23308 (N_23308,N_20028,N_21252);
nand U23309 (N_23309,N_20002,N_20910);
nand U23310 (N_23310,N_20355,N_21141);
xnor U23311 (N_23311,N_19575,N_18776);
nand U23312 (N_23312,N_20180,N_20774);
and U23313 (N_23313,N_19877,N_20386);
nand U23314 (N_23314,N_20775,N_18880);
nor U23315 (N_23315,N_19743,N_21355);
nor U23316 (N_23316,N_19463,N_19000);
xnor U23317 (N_23317,N_18983,N_20117);
or U23318 (N_23318,N_19131,N_20614);
nand U23319 (N_23319,N_20778,N_18958);
xor U23320 (N_23320,N_21376,N_20868);
nor U23321 (N_23321,N_19473,N_21632);
xnor U23322 (N_23322,N_19380,N_19329);
xor U23323 (N_23323,N_18857,N_20048);
or U23324 (N_23324,N_21391,N_21205);
nand U23325 (N_23325,N_20270,N_18894);
or U23326 (N_23326,N_19644,N_19125);
or U23327 (N_23327,N_19833,N_19606);
or U23328 (N_23328,N_21749,N_20213);
or U23329 (N_23329,N_21724,N_19448);
and U23330 (N_23330,N_19244,N_21833);
nand U23331 (N_23331,N_18752,N_19126);
nor U23332 (N_23332,N_20801,N_20214);
and U23333 (N_23333,N_19769,N_20470);
nand U23334 (N_23334,N_20571,N_19549);
or U23335 (N_23335,N_19754,N_21630);
or U23336 (N_23336,N_21545,N_21432);
nor U23337 (N_23337,N_20132,N_20694);
and U23338 (N_23338,N_19421,N_18936);
xor U23339 (N_23339,N_21240,N_20521);
nand U23340 (N_23340,N_21396,N_19251);
nand U23341 (N_23341,N_19204,N_20105);
or U23342 (N_23342,N_19558,N_20559);
xor U23343 (N_23343,N_18949,N_19520);
and U23344 (N_23344,N_20299,N_20684);
xnor U23345 (N_23345,N_21366,N_19415);
or U23346 (N_23346,N_20414,N_20328);
nor U23347 (N_23347,N_20199,N_21422);
xnor U23348 (N_23348,N_20667,N_20252);
xor U23349 (N_23349,N_19535,N_19941);
and U23350 (N_23350,N_19032,N_20949);
nand U23351 (N_23351,N_21709,N_19873);
nand U23352 (N_23352,N_19695,N_19475);
and U23353 (N_23353,N_19129,N_21766);
or U23354 (N_23354,N_19818,N_19508);
nand U23355 (N_23355,N_21359,N_20878);
nor U23356 (N_23356,N_19986,N_21597);
or U23357 (N_23357,N_19146,N_20906);
or U23358 (N_23358,N_19791,N_21504);
xnor U23359 (N_23359,N_19837,N_18765);
nand U23360 (N_23360,N_19505,N_19384);
nor U23361 (N_23361,N_21490,N_19362);
xnor U23362 (N_23362,N_20055,N_21335);
xnor U23363 (N_23363,N_18785,N_20269);
xor U23364 (N_23364,N_19633,N_20692);
nand U23365 (N_23365,N_19400,N_19577);
and U23366 (N_23366,N_20139,N_20875);
xor U23367 (N_23367,N_21487,N_21475);
xor U23368 (N_23368,N_19847,N_19595);
nor U23369 (N_23369,N_19423,N_21455);
or U23370 (N_23370,N_21385,N_21595);
nand U23371 (N_23371,N_19826,N_18808);
nand U23372 (N_23372,N_19469,N_18762);
xnor U23373 (N_23373,N_20794,N_18825);
xor U23374 (N_23374,N_20069,N_20485);
and U23375 (N_23375,N_20553,N_19960);
nand U23376 (N_23376,N_20458,N_20819);
or U23377 (N_23377,N_20273,N_18873);
nand U23378 (N_23378,N_20291,N_19736);
or U23379 (N_23379,N_20789,N_21491);
or U23380 (N_23380,N_19192,N_20389);
nor U23381 (N_23381,N_19666,N_18956);
nor U23382 (N_23382,N_21675,N_19934);
xor U23383 (N_23383,N_20123,N_21017);
nand U23384 (N_23384,N_20780,N_20194);
nor U23385 (N_23385,N_20453,N_19259);
and U23386 (N_23386,N_20275,N_19180);
xor U23387 (N_23387,N_19842,N_20824);
and U23388 (N_23388,N_19665,N_19141);
or U23389 (N_23389,N_21161,N_21772);
nor U23390 (N_23390,N_19749,N_19158);
nand U23391 (N_23391,N_20445,N_20927);
or U23392 (N_23392,N_21839,N_18795);
and U23393 (N_23393,N_19430,N_21398);
nor U23394 (N_23394,N_20226,N_20193);
or U23395 (N_23395,N_19651,N_19205);
or U23396 (N_23396,N_21114,N_21297);
and U23397 (N_23397,N_19403,N_21745);
and U23398 (N_23398,N_21539,N_20818);
nor U23399 (N_23399,N_21516,N_21737);
nor U23400 (N_23400,N_21494,N_21329);
nor U23401 (N_23401,N_19658,N_21777);
nand U23402 (N_23402,N_21642,N_20748);
xor U23403 (N_23403,N_19202,N_19951);
xnor U23404 (N_23404,N_18961,N_19003);
xnor U23405 (N_23405,N_21158,N_21589);
xor U23406 (N_23406,N_19498,N_19879);
and U23407 (N_23407,N_18836,N_19617);
nand U23408 (N_23408,N_19720,N_20699);
nand U23409 (N_23409,N_19836,N_18876);
xor U23410 (N_23410,N_21412,N_19096);
xnor U23411 (N_23411,N_21287,N_19719);
and U23412 (N_23412,N_20361,N_20009);
and U23413 (N_23413,N_19795,N_20652);
nor U23414 (N_23414,N_19427,N_20687);
xor U23415 (N_23415,N_21003,N_21095);
or U23416 (N_23416,N_19831,N_19058);
or U23417 (N_23417,N_21280,N_20590);
nor U23418 (N_23418,N_20121,N_20524);
nand U23419 (N_23419,N_19044,N_18852);
xnor U23420 (N_23420,N_19507,N_19685);
or U23421 (N_23421,N_21006,N_20228);
and U23422 (N_23422,N_20950,N_19174);
and U23423 (N_23423,N_21323,N_19315);
nand U23424 (N_23424,N_19232,N_21181);
and U23425 (N_23425,N_20842,N_19835);
nand U23426 (N_23426,N_19636,N_20581);
nand U23427 (N_23427,N_20265,N_21256);
xor U23428 (N_23428,N_18959,N_19616);
xor U23429 (N_23429,N_19723,N_20802);
and U23430 (N_23430,N_21203,N_21350);
nand U23431 (N_23431,N_21852,N_20931);
and U23432 (N_23432,N_21404,N_19881);
or U23433 (N_23433,N_20108,N_20436);
nor U23434 (N_23434,N_19235,N_19070);
xnor U23435 (N_23435,N_19124,N_21447);
xnor U23436 (N_23436,N_19528,N_20843);
or U23437 (N_23437,N_20162,N_19779);
nand U23438 (N_23438,N_20299,N_19170);
nor U23439 (N_23439,N_21060,N_21673);
nand U23440 (N_23440,N_20182,N_20097);
or U23441 (N_23441,N_21650,N_21475);
xor U23442 (N_23442,N_18857,N_19355);
and U23443 (N_23443,N_19048,N_21202);
and U23444 (N_23444,N_21662,N_19653);
and U23445 (N_23445,N_21547,N_20890);
nand U23446 (N_23446,N_19422,N_21478);
or U23447 (N_23447,N_20004,N_21553);
and U23448 (N_23448,N_20984,N_21738);
or U23449 (N_23449,N_21549,N_20520);
xnor U23450 (N_23450,N_21191,N_19724);
nor U23451 (N_23451,N_20369,N_18842);
nand U23452 (N_23452,N_20394,N_20681);
or U23453 (N_23453,N_21018,N_21658);
or U23454 (N_23454,N_19935,N_21388);
nand U23455 (N_23455,N_21419,N_21235);
nor U23456 (N_23456,N_21390,N_19098);
or U23457 (N_23457,N_18866,N_21851);
and U23458 (N_23458,N_21775,N_19294);
and U23459 (N_23459,N_21574,N_20513);
nor U23460 (N_23460,N_18826,N_20178);
or U23461 (N_23461,N_21115,N_19649);
or U23462 (N_23462,N_21448,N_20914);
nand U23463 (N_23463,N_19314,N_18875);
or U23464 (N_23464,N_18942,N_18902);
and U23465 (N_23465,N_21831,N_20848);
nand U23466 (N_23466,N_20992,N_21356);
nor U23467 (N_23467,N_20368,N_20293);
xnor U23468 (N_23468,N_19481,N_20871);
and U23469 (N_23469,N_20323,N_18982);
nand U23470 (N_23470,N_21026,N_21774);
nor U23471 (N_23471,N_20827,N_18965);
or U23472 (N_23472,N_18925,N_21386);
nor U23473 (N_23473,N_19050,N_20658);
or U23474 (N_23474,N_21431,N_18972);
and U23475 (N_23475,N_19574,N_20389);
xor U23476 (N_23476,N_21771,N_19499);
or U23477 (N_23477,N_21440,N_21230);
nor U23478 (N_23478,N_19575,N_20290);
xnor U23479 (N_23479,N_20328,N_20111);
nor U23480 (N_23480,N_20570,N_19013);
nand U23481 (N_23481,N_18784,N_19427);
nor U23482 (N_23482,N_19281,N_20736);
or U23483 (N_23483,N_20848,N_21421);
nand U23484 (N_23484,N_20169,N_19959);
nand U23485 (N_23485,N_21644,N_20466);
and U23486 (N_23486,N_20886,N_21281);
nand U23487 (N_23487,N_20140,N_21367);
xor U23488 (N_23488,N_19723,N_21460);
nor U23489 (N_23489,N_20410,N_21530);
xor U23490 (N_23490,N_20683,N_19738);
and U23491 (N_23491,N_21503,N_21257);
or U23492 (N_23492,N_19063,N_19300);
nor U23493 (N_23493,N_21378,N_20359);
nor U23494 (N_23494,N_20053,N_21039);
nor U23495 (N_23495,N_21497,N_18822);
xnor U23496 (N_23496,N_19555,N_21420);
xor U23497 (N_23497,N_19358,N_21147);
and U23498 (N_23498,N_19359,N_21041);
xnor U23499 (N_23499,N_18863,N_20165);
and U23500 (N_23500,N_21259,N_21060);
and U23501 (N_23501,N_21800,N_20938);
nand U23502 (N_23502,N_19323,N_20160);
xor U23503 (N_23503,N_19410,N_21384);
nor U23504 (N_23504,N_20610,N_19887);
nor U23505 (N_23505,N_19761,N_19213);
xnor U23506 (N_23506,N_18890,N_19821);
xor U23507 (N_23507,N_18842,N_21326);
or U23508 (N_23508,N_18952,N_20344);
and U23509 (N_23509,N_21848,N_21614);
or U23510 (N_23510,N_18893,N_21617);
or U23511 (N_23511,N_21585,N_19617);
and U23512 (N_23512,N_18862,N_20058);
xnor U23513 (N_23513,N_19156,N_19257);
nor U23514 (N_23514,N_21222,N_21674);
nor U23515 (N_23515,N_20648,N_19965);
or U23516 (N_23516,N_19300,N_19741);
or U23517 (N_23517,N_21051,N_18937);
xnor U23518 (N_23518,N_20726,N_20842);
nand U23519 (N_23519,N_21540,N_20481);
and U23520 (N_23520,N_18990,N_19038);
nand U23521 (N_23521,N_18950,N_19315);
nor U23522 (N_23522,N_19144,N_20137);
or U23523 (N_23523,N_21291,N_21678);
or U23524 (N_23524,N_20325,N_19067);
or U23525 (N_23525,N_20305,N_21010);
and U23526 (N_23526,N_20962,N_19232);
xnor U23527 (N_23527,N_21754,N_21675);
nand U23528 (N_23528,N_20494,N_21136);
nor U23529 (N_23529,N_20891,N_19092);
and U23530 (N_23530,N_21572,N_19273);
and U23531 (N_23531,N_20027,N_19109);
nand U23532 (N_23532,N_20965,N_21038);
nor U23533 (N_23533,N_20505,N_19384);
nand U23534 (N_23534,N_19525,N_19238);
xor U23535 (N_23535,N_21546,N_18830);
nand U23536 (N_23536,N_20254,N_19710);
nand U23537 (N_23537,N_20394,N_18868);
nand U23538 (N_23538,N_19002,N_20014);
nand U23539 (N_23539,N_19169,N_20566);
nand U23540 (N_23540,N_21180,N_21211);
and U23541 (N_23541,N_20032,N_21557);
or U23542 (N_23542,N_21548,N_21622);
nor U23543 (N_23543,N_21873,N_20280);
xor U23544 (N_23544,N_20655,N_19144);
or U23545 (N_23545,N_20597,N_21762);
and U23546 (N_23546,N_21125,N_19021);
xor U23547 (N_23547,N_20577,N_21109);
and U23548 (N_23548,N_20600,N_19160);
nand U23549 (N_23549,N_20350,N_20640);
or U23550 (N_23550,N_19231,N_21210);
or U23551 (N_23551,N_19154,N_20704);
nor U23552 (N_23552,N_21841,N_18927);
xnor U23553 (N_23553,N_21059,N_20600);
and U23554 (N_23554,N_21304,N_20631);
nand U23555 (N_23555,N_20446,N_21451);
nor U23556 (N_23556,N_20375,N_19868);
or U23557 (N_23557,N_21091,N_19317);
nor U23558 (N_23558,N_20193,N_20286);
and U23559 (N_23559,N_20343,N_19483);
nand U23560 (N_23560,N_19708,N_19088);
nor U23561 (N_23561,N_19477,N_20970);
and U23562 (N_23562,N_20347,N_21417);
or U23563 (N_23563,N_21139,N_19327);
nand U23564 (N_23564,N_20384,N_21599);
xnor U23565 (N_23565,N_18906,N_18872);
or U23566 (N_23566,N_19949,N_21596);
nand U23567 (N_23567,N_19288,N_19996);
or U23568 (N_23568,N_21168,N_19327);
nor U23569 (N_23569,N_20940,N_20678);
nand U23570 (N_23570,N_21517,N_19750);
nor U23571 (N_23571,N_21038,N_18764);
and U23572 (N_23572,N_18782,N_19266);
and U23573 (N_23573,N_20271,N_21128);
xor U23574 (N_23574,N_19244,N_19270);
nor U23575 (N_23575,N_21209,N_19551);
nor U23576 (N_23576,N_19335,N_20890);
nor U23577 (N_23577,N_20354,N_20006);
and U23578 (N_23578,N_20808,N_19292);
nand U23579 (N_23579,N_19097,N_20262);
and U23580 (N_23580,N_19953,N_21095);
xnor U23581 (N_23581,N_21191,N_21359);
or U23582 (N_23582,N_19768,N_21293);
nand U23583 (N_23583,N_20397,N_20671);
nor U23584 (N_23584,N_20113,N_21707);
nand U23585 (N_23585,N_19222,N_19528);
and U23586 (N_23586,N_20504,N_19396);
nand U23587 (N_23587,N_20704,N_19817);
or U23588 (N_23588,N_20709,N_21247);
nand U23589 (N_23589,N_19116,N_19759);
nor U23590 (N_23590,N_19539,N_19552);
nor U23591 (N_23591,N_18930,N_21690);
or U23592 (N_23592,N_19765,N_21701);
xnor U23593 (N_23593,N_20764,N_20550);
xnor U23594 (N_23594,N_18791,N_21627);
xor U23595 (N_23595,N_20446,N_18891);
or U23596 (N_23596,N_18774,N_19558);
nor U23597 (N_23597,N_20631,N_20014);
or U23598 (N_23598,N_19503,N_21707);
and U23599 (N_23599,N_20276,N_19832);
nand U23600 (N_23600,N_19100,N_21620);
and U23601 (N_23601,N_21036,N_19845);
or U23602 (N_23602,N_20794,N_19218);
nand U23603 (N_23603,N_19343,N_21357);
nand U23604 (N_23604,N_21374,N_20363);
nand U23605 (N_23605,N_21126,N_21836);
xor U23606 (N_23606,N_20240,N_19667);
nand U23607 (N_23607,N_20970,N_20016);
nor U23608 (N_23608,N_19373,N_20638);
and U23609 (N_23609,N_19091,N_21698);
nand U23610 (N_23610,N_19505,N_20260);
xor U23611 (N_23611,N_20810,N_20351);
nor U23612 (N_23612,N_21873,N_19518);
nand U23613 (N_23613,N_21132,N_20459);
nor U23614 (N_23614,N_20742,N_21498);
nand U23615 (N_23615,N_20099,N_19125);
nand U23616 (N_23616,N_18886,N_19813);
or U23617 (N_23617,N_20315,N_19817);
nand U23618 (N_23618,N_19580,N_19421);
nor U23619 (N_23619,N_21190,N_20041);
and U23620 (N_23620,N_20630,N_19440);
xor U23621 (N_23621,N_21399,N_19953);
nor U23622 (N_23622,N_21834,N_21827);
nand U23623 (N_23623,N_21127,N_19272);
or U23624 (N_23624,N_20566,N_20012);
xnor U23625 (N_23625,N_19501,N_20757);
xor U23626 (N_23626,N_19110,N_21084);
and U23627 (N_23627,N_20974,N_20264);
nor U23628 (N_23628,N_18888,N_20259);
xnor U23629 (N_23629,N_18932,N_18947);
or U23630 (N_23630,N_21567,N_20332);
nand U23631 (N_23631,N_20191,N_19938);
xnor U23632 (N_23632,N_18865,N_20559);
or U23633 (N_23633,N_19396,N_21175);
xor U23634 (N_23634,N_19411,N_19732);
nand U23635 (N_23635,N_21484,N_19319);
nand U23636 (N_23636,N_19950,N_19561);
or U23637 (N_23637,N_19540,N_21327);
and U23638 (N_23638,N_20003,N_20485);
nand U23639 (N_23639,N_19555,N_18923);
nor U23640 (N_23640,N_20394,N_19979);
and U23641 (N_23641,N_20699,N_21155);
nand U23642 (N_23642,N_20878,N_21619);
nor U23643 (N_23643,N_21810,N_19198);
xnor U23644 (N_23644,N_20118,N_20493);
or U23645 (N_23645,N_20807,N_21160);
or U23646 (N_23646,N_19321,N_20073);
or U23647 (N_23647,N_19691,N_21728);
and U23648 (N_23648,N_18995,N_19851);
and U23649 (N_23649,N_20510,N_19028);
xor U23650 (N_23650,N_20262,N_18987);
xnor U23651 (N_23651,N_20803,N_20169);
nand U23652 (N_23652,N_19840,N_19637);
and U23653 (N_23653,N_20430,N_19459);
or U23654 (N_23654,N_21158,N_20183);
nand U23655 (N_23655,N_20172,N_18991);
or U23656 (N_23656,N_19933,N_21540);
xor U23657 (N_23657,N_19119,N_19896);
and U23658 (N_23658,N_21086,N_19777);
or U23659 (N_23659,N_19027,N_19612);
nand U23660 (N_23660,N_20417,N_19976);
xnor U23661 (N_23661,N_21610,N_19217);
xor U23662 (N_23662,N_21721,N_20715);
nor U23663 (N_23663,N_19221,N_21159);
nand U23664 (N_23664,N_20148,N_21160);
nand U23665 (N_23665,N_20583,N_20301);
nor U23666 (N_23666,N_19189,N_19992);
nor U23667 (N_23667,N_21336,N_21811);
nor U23668 (N_23668,N_21067,N_20447);
xor U23669 (N_23669,N_20277,N_19966);
nor U23670 (N_23670,N_19117,N_19828);
nand U23671 (N_23671,N_18984,N_19398);
and U23672 (N_23672,N_21125,N_21095);
or U23673 (N_23673,N_19934,N_19667);
and U23674 (N_23674,N_19081,N_19334);
and U23675 (N_23675,N_19603,N_20843);
nand U23676 (N_23676,N_21724,N_20060);
nand U23677 (N_23677,N_20306,N_20651);
or U23678 (N_23678,N_18951,N_19703);
xor U23679 (N_23679,N_19343,N_19649);
nor U23680 (N_23680,N_21843,N_18995);
and U23681 (N_23681,N_18959,N_19326);
nor U23682 (N_23682,N_19520,N_18830);
and U23683 (N_23683,N_19269,N_20780);
or U23684 (N_23684,N_20514,N_19075);
or U23685 (N_23685,N_18755,N_18959);
xnor U23686 (N_23686,N_19665,N_21055);
nand U23687 (N_23687,N_21059,N_21866);
xnor U23688 (N_23688,N_21077,N_20205);
and U23689 (N_23689,N_20798,N_20407);
nand U23690 (N_23690,N_19932,N_19200);
xor U23691 (N_23691,N_21728,N_21614);
or U23692 (N_23692,N_19641,N_19786);
or U23693 (N_23693,N_19327,N_21682);
nor U23694 (N_23694,N_21199,N_21392);
nand U23695 (N_23695,N_19433,N_19125);
and U23696 (N_23696,N_21686,N_19560);
nor U23697 (N_23697,N_18945,N_20861);
nor U23698 (N_23698,N_21672,N_21650);
xnor U23699 (N_23699,N_19167,N_21095);
or U23700 (N_23700,N_21226,N_19274);
or U23701 (N_23701,N_19292,N_20331);
xor U23702 (N_23702,N_20663,N_19786);
or U23703 (N_23703,N_20236,N_18856);
or U23704 (N_23704,N_20420,N_21693);
nor U23705 (N_23705,N_20848,N_18820);
or U23706 (N_23706,N_21385,N_20585);
xor U23707 (N_23707,N_20187,N_19817);
nor U23708 (N_23708,N_20100,N_20832);
xnor U23709 (N_23709,N_19077,N_20947);
or U23710 (N_23710,N_19934,N_19575);
nand U23711 (N_23711,N_19418,N_19302);
nand U23712 (N_23712,N_21471,N_21704);
or U23713 (N_23713,N_19226,N_19043);
nand U23714 (N_23714,N_21203,N_21728);
xnor U23715 (N_23715,N_20020,N_21241);
xnor U23716 (N_23716,N_20697,N_20608);
or U23717 (N_23717,N_18832,N_20140);
and U23718 (N_23718,N_19202,N_20476);
or U23719 (N_23719,N_21165,N_20209);
xor U23720 (N_23720,N_21421,N_19662);
or U23721 (N_23721,N_18932,N_18892);
xnor U23722 (N_23722,N_20173,N_18797);
or U23723 (N_23723,N_20965,N_20663);
nand U23724 (N_23724,N_20876,N_21590);
and U23725 (N_23725,N_19859,N_20459);
and U23726 (N_23726,N_19770,N_21839);
nor U23727 (N_23727,N_19489,N_21261);
xnor U23728 (N_23728,N_18788,N_19424);
nand U23729 (N_23729,N_19821,N_21851);
and U23730 (N_23730,N_19720,N_21161);
or U23731 (N_23731,N_21624,N_20829);
and U23732 (N_23732,N_19139,N_21473);
and U23733 (N_23733,N_19383,N_21728);
xor U23734 (N_23734,N_19199,N_21460);
and U23735 (N_23735,N_21189,N_20783);
and U23736 (N_23736,N_19617,N_20918);
nor U23737 (N_23737,N_19789,N_21771);
xor U23738 (N_23738,N_21703,N_18800);
or U23739 (N_23739,N_19936,N_20085);
xnor U23740 (N_23740,N_18990,N_21666);
or U23741 (N_23741,N_20463,N_20813);
nand U23742 (N_23742,N_20558,N_20086);
and U23743 (N_23743,N_19787,N_20747);
nand U23744 (N_23744,N_21416,N_21290);
nand U23745 (N_23745,N_21145,N_19790);
or U23746 (N_23746,N_20841,N_21454);
nor U23747 (N_23747,N_21173,N_19613);
or U23748 (N_23748,N_20804,N_21753);
nand U23749 (N_23749,N_21114,N_18908);
or U23750 (N_23750,N_20918,N_20723);
or U23751 (N_23751,N_19209,N_21569);
and U23752 (N_23752,N_20440,N_19553);
xnor U23753 (N_23753,N_19269,N_20137);
xnor U23754 (N_23754,N_20864,N_20889);
nor U23755 (N_23755,N_19620,N_20784);
and U23756 (N_23756,N_20015,N_21520);
nand U23757 (N_23757,N_19141,N_18790);
or U23758 (N_23758,N_21171,N_21673);
or U23759 (N_23759,N_21544,N_20029);
nor U23760 (N_23760,N_21692,N_18985);
xor U23761 (N_23761,N_20323,N_19659);
and U23762 (N_23762,N_19815,N_21312);
nor U23763 (N_23763,N_21595,N_20570);
or U23764 (N_23764,N_20941,N_20108);
nand U23765 (N_23765,N_19827,N_20823);
nor U23766 (N_23766,N_21347,N_21061);
and U23767 (N_23767,N_20143,N_19966);
or U23768 (N_23768,N_18926,N_19759);
nor U23769 (N_23769,N_21444,N_21824);
and U23770 (N_23770,N_19872,N_19531);
and U23771 (N_23771,N_19657,N_19155);
or U23772 (N_23772,N_20190,N_19791);
nor U23773 (N_23773,N_19520,N_19415);
nor U23774 (N_23774,N_18774,N_19956);
nand U23775 (N_23775,N_19329,N_21335);
nor U23776 (N_23776,N_20948,N_19056);
nand U23777 (N_23777,N_21560,N_19645);
nand U23778 (N_23778,N_19124,N_20520);
nand U23779 (N_23779,N_21581,N_21818);
nor U23780 (N_23780,N_20477,N_20049);
xor U23781 (N_23781,N_20698,N_20619);
nand U23782 (N_23782,N_20596,N_19979);
or U23783 (N_23783,N_20511,N_19842);
xor U23784 (N_23784,N_20361,N_19263);
nand U23785 (N_23785,N_20105,N_21459);
or U23786 (N_23786,N_20911,N_19869);
and U23787 (N_23787,N_19683,N_19463);
nand U23788 (N_23788,N_19091,N_20089);
and U23789 (N_23789,N_20400,N_20426);
xor U23790 (N_23790,N_19340,N_19715);
and U23791 (N_23791,N_21080,N_18915);
nor U23792 (N_23792,N_18880,N_20786);
or U23793 (N_23793,N_21083,N_21528);
nand U23794 (N_23794,N_18804,N_19126);
or U23795 (N_23795,N_20851,N_19466);
nand U23796 (N_23796,N_20465,N_19432);
and U23797 (N_23797,N_20576,N_19263);
or U23798 (N_23798,N_19812,N_21817);
or U23799 (N_23799,N_20224,N_20709);
nand U23800 (N_23800,N_19379,N_20274);
xnor U23801 (N_23801,N_19853,N_21412);
nor U23802 (N_23802,N_21235,N_19145);
or U23803 (N_23803,N_19021,N_21549);
nor U23804 (N_23804,N_18964,N_20970);
and U23805 (N_23805,N_21531,N_19785);
xnor U23806 (N_23806,N_21194,N_21583);
nand U23807 (N_23807,N_19148,N_20435);
nand U23808 (N_23808,N_19923,N_20277);
xnor U23809 (N_23809,N_19600,N_21167);
and U23810 (N_23810,N_20302,N_21380);
nand U23811 (N_23811,N_19510,N_20386);
nor U23812 (N_23812,N_19507,N_19123);
xnor U23813 (N_23813,N_18940,N_20207);
and U23814 (N_23814,N_19804,N_21627);
nand U23815 (N_23815,N_19642,N_20689);
nor U23816 (N_23816,N_21229,N_19528);
or U23817 (N_23817,N_19336,N_20718);
and U23818 (N_23818,N_21468,N_19236);
nor U23819 (N_23819,N_21164,N_18955);
nand U23820 (N_23820,N_20783,N_19838);
or U23821 (N_23821,N_19741,N_20209);
xnor U23822 (N_23822,N_20674,N_20264);
nor U23823 (N_23823,N_21270,N_20390);
and U23824 (N_23824,N_18944,N_20103);
or U23825 (N_23825,N_21324,N_19139);
and U23826 (N_23826,N_21366,N_19080);
nand U23827 (N_23827,N_21379,N_19290);
or U23828 (N_23828,N_21146,N_20954);
and U23829 (N_23829,N_21045,N_19262);
or U23830 (N_23830,N_20135,N_19025);
or U23831 (N_23831,N_19246,N_21674);
xnor U23832 (N_23832,N_21355,N_20510);
xor U23833 (N_23833,N_19474,N_19511);
xnor U23834 (N_23834,N_19916,N_21274);
nand U23835 (N_23835,N_19001,N_21202);
and U23836 (N_23836,N_19925,N_21381);
nor U23837 (N_23837,N_20147,N_20911);
nor U23838 (N_23838,N_21652,N_19153);
and U23839 (N_23839,N_20274,N_20668);
nor U23840 (N_23840,N_19015,N_21147);
and U23841 (N_23841,N_21634,N_21031);
nand U23842 (N_23842,N_21729,N_20502);
nor U23843 (N_23843,N_20624,N_18893);
xnor U23844 (N_23844,N_19609,N_19997);
nand U23845 (N_23845,N_21815,N_21665);
nand U23846 (N_23846,N_19128,N_18898);
nand U23847 (N_23847,N_20048,N_20682);
xor U23848 (N_23848,N_20940,N_19495);
nor U23849 (N_23849,N_20236,N_21392);
or U23850 (N_23850,N_21107,N_20002);
nand U23851 (N_23851,N_19333,N_20827);
and U23852 (N_23852,N_20528,N_19929);
nor U23853 (N_23853,N_20683,N_20920);
xor U23854 (N_23854,N_19630,N_19508);
and U23855 (N_23855,N_20735,N_20346);
nand U23856 (N_23856,N_19515,N_21751);
xnor U23857 (N_23857,N_19993,N_21850);
nor U23858 (N_23858,N_21182,N_19095);
and U23859 (N_23859,N_19808,N_20890);
or U23860 (N_23860,N_19189,N_18809);
nand U23861 (N_23861,N_19412,N_21742);
xor U23862 (N_23862,N_20039,N_20107);
or U23863 (N_23863,N_19156,N_19816);
nand U23864 (N_23864,N_20278,N_19035);
nand U23865 (N_23865,N_19794,N_20874);
nand U23866 (N_23866,N_21025,N_21324);
and U23867 (N_23867,N_20573,N_18863);
and U23868 (N_23868,N_19166,N_21614);
nand U23869 (N_23869,N_21160,N_21010);
xor U23870 (N_23870,N_21535,N_20685);
xor U23871 (N_23871,N_18833,N_20729);
nand U23872 (N_23872,N_20104,N_21703);
xor U23873 (N_23873,N_20902,N_19158);
nor U23874 (N_23874,N_20223,N_19102);
nand U23875 (N_23875,N_21538,N_19952);
and U23876 (N_23876,N_19814,N_21046);
nor U23877 (N_23877,N_20752,N_20248);
nand U23878 (N_23878,N_21836,N_21033);
nor U23879 (N_23879,N_21072,N_20058);
or U23880 (N_23880,N_20934,N_21692);
xnor U23881 (N_23881,N_21486,N_21514);
nand U23882 (N_23882,N_19626,N_19323);
nor U23883 (N_23883,N_20363,N_19429);
nor U23884 (N_23884,N_21381,N_21769);
nand U23885 (N_23885,N_21566,N_18802);
and U23886 (N_23886,N_19132,N_21798);
xor U23887 (N_23887,N_19820,N_19261);
nor U23888 (N_23888,N_20455,N_20397);
xnor U23889 (N_23889,N_19317,N_21793);
nand U23890 (N_23890,N_21465,N_18845);
nor U23891 (N_23891,N_19313,N_21082);
and U23892 (N_23892,N_20515,N_20617);
nor U23893 (N_23893,N_21465,N_19143);
nor U23894 (N_23894,N_19095,N_21670);
xnor U23895 (N_23895,N_21221,N_19730);
or U23896 (N_23896,N_19258,N_19438);
xor U23897 (N_23897,N_19675,N_21182);
or U23898 (N_23898,N_21190,N_20653);
xnor U23899 (N_23899,N_20396,N_18920);
and U23900 (N_23900,N_20929,N_18871);
or U23901 (N_23901,N_21873,N_18777);
or U23902 (N_23902,N_19335,N_20350);
nor U23903 (N_23903,N_20974,N_21026);
or U23904 (N_23904,N_20085,N_19873);
xnor U23905 (N_23905,N_21327,N_20276);
nor U23906 (N_23906,N_21698,N_21862);
or U23907 (N_23907,N_19285,N_21666);
nand U23908 (N_23908,N_19105,N_21257);
nor U23909 (N_23909,N_18811,N_20367);
xor U23910 (N_23910,N_20022,N_18799);
nor U23911 (N_23911,N_21586,N_19148);
and U23912 (N_23912,N_20039,N_19072);
nand U23913 (N_23913,N_21742,N_19136);
or U23914 (N_23914,N_20064,N_21751);
xnor U23915 (N_23915,N_19256,N_18816);
nand U23916 (N_23916,N_19469,N_19332);
and U23917 (N_23917,N_21812,N_19475);
or U23918 (N_23918,N_19390,N_20866);
and U23919 (N_23919,N_21736,N_19523);
nor U23920 (N_23920,N_20881,N_20348);
nand U23921 (N_23921,N_20944,N_21689);
nor U23922 (N_23922,N_20666,N_21674);
nor U23923 (N_23923,N_21201,N_19916);
xnor U23924 (N_23924,N_19716,N_20607);
nor U23925 (N_23925,N_21859,N_19159);
nor U23926 (N_23926,N_21721,N_19123);
or U23927 (N_23927,N_20110,N_18949);
and U23928 (N_23928,N_21498,N_21509);
or U23929 (N_23929,N_21736,N_20451);
or U23930 (N_23930,N_20670,N_20407);
nor U23931 (N_23931,N_21054,N_19193);
nor U23932 (N_23932,N_18911,N_21604);
and U23933 (N_23933,N_20142,N_19323);
and U23934 (N_23934,N_21688,N_20785);
nor U23935 (N_23935,N_18872,N_19819);
and U23936 (N_23936,N_21164,N_19247);
and U23937 (N_23937,N_20651,N_19295);
or U23938 (N_23938,N_20818,N_19844);
nor U23939 (N_23939,N_21253,N_19843);
nor U23940 (N_23940,N_21542,N_20307);
xor U23941 (N_23941,N_19632,N_21220);
and U23942 (N_23942,N_20793,N_19233);
or U23943 (N_23943,N_20435,N_19490);
or U23944 (N_23944,N_19291,N_19968);
and U23945 (N_23945,N_21485,N_21399);
or U23946 (N_23946,N_19549,N_19340);
nor U23947 (N_23947,N_20555,N_19644);
nand U23948 (N_23948,N_21288,N_20482);
or U23949 (N_23949,N_21094,N_21420);
or U23950 (N_23950,N_21081,N_21858);
xnor U23951 (N_23951,N_21551,N_20996);
nand U23952 (N_23952,N_19384,N_20261);
nand U23953 (N_23953,N_19722,N_18758);
or U23954 (N_23954,N_20554,N_21073);
and U23955 (N_23955,N_18816,N_21770);
nand U23956 (N_23956,N_21380,N_21144);
nand U23957 (N_23957,N_19727,N_20579);
nor U23958 (N_23958,N_19407,N_20927);
nor U23959 (N_23959,N_19213,N_21074);
nand U23960 (N_23960,N_21072,N_21378);
nor U23961 (N_23961,N_20964,N_19524);
xnor U23962 (N_23962,N_21540,N_21827);
xor U23963 (N_23963,N_21642,N_21770);
or U23964 (N_23964,N_19088,N_18972);
xor U23965 (N_23965,N_19097,N_21420);
xnor U23966 (N_23966,N_19244,N_19176);
or U23967 (N_23967,N_19006,N_21287);
or U23968 (N_23968,N_19110,N_19503);
nand U23969 (N_23969,N_20509,N_19191);
xor U23970 (N_23970,N_20110,N_20408);
and U23971 (N_23971,N_21147,N_21496);
and U23972 (N_23972,N_20655,N_19434);
xnor U23973 (N_23973,N_21072,N_19300);
and U23974 (N_23974,N_21170,N_21597);
and U23975 (N_23975,N_19233,N_21447);
nand U23976 (N_23976,N_20818,N_21764);
nor U23977 (N_23977,N_20504,N_18911);
nor U23978 (N_23978,N_21746,N_21232);
xor U23979 (N_23979,N_19422,N_21539);
nand U23980 (N_23980,N_19186,N_21866);
nand U23981 (N_23981,N_18773,N_21026);
and U23982 (N_23982,N_20842,N_19032);
and U23983 (N_23983,N_19876,N_19600);
xor U23984 (N_23984,N_19654,N_19397);
or U23985 (N_23985,N_19083,N_19458);
xor U23986 (N_23986,N_19995,N_19024);
and U23987 (N_23987,N_19782,N_19084);
nor U23988 (N_23988,N_19552,N_19119);
or U23989 (N_23989,N_21713,N_20713);
nor U23990 (N_23990,N_20458,N_21462);
nand U23991 (N_23991,N_21504,N_20919);
and U23992 (N_23992,N_21426,N_20635);
or U23993 (N_23993,N_20686,N_21781);
xnor U23994 (N_23994,N_19322,N_21638);
nor U23995 (N_23995,N_19058,N_19865);
nor U23996 (N_23996,N_21805,N_21355);
or U23997 (N_23997,N_19477,N_21766);
or U23998 (N_23998,N_20099,N_19012);
nand U23999 (N_23999,N_21015,N_20305);
xor U24000 (N_24000,N_21065,N_19558);
and U24001 (N_24001,N_20688,N_18886);
nand U24002 (N_24002,N_18770,N_18924);
nor U24003 (N_24003,N_20011,N_20714);
or U24004 (N_24004,N_18949,N_21489);
nor U24005 (N_24005,N_20536,N_19480);
nand U24006 (N_24006,N_18949,N_21417);
nor U24007 (N_24007,N_20179,N_21792);
or U24008 (N_24008,N_18944,N_18824);
nor U24009 (N_24009,N_19623,N_20737);
xnor U24010 (N_24010,N_20612,N_21729);
xor U24011 (N_24011,N_20484,N_21215);
nand U24012 (N_24012,N_21867,N_20201);
nand U24013 (N_24013,N_20738,N_21063);
and U24014 (N_24014,N_21081,N_20264);
xor U24015 (N_24015,N_20433,N_19451);
nand U24016 (N_24016,N_19270,N_20381);
and U24017 (N_24017,N_18946,N_21207);
or U24018 (N_24018,N_21324,N_20752);
or U24019 (N_24019,N_21511,N_21293);
xor U24020 (N_24020,N_21448,N_21407);
nor U24021 (N_24021,N_21410,N_19939);
nand U24022 (N_24022,N_21270,N_19908);
nor U24023 (N_24023,N_18935,N_21329);
nand U24024 (N_24024,N_21162,N_20229);
or U24025 (N_24025,N_20931,N_20325);
nand U24026 (N_24026,N_21648,N_21631);
or U24027 (N_24027,N_18910,N_20315);
nor U24028 (N_24028,N_19746,N_19528);
or U24029 (N_24029,N_18797,N_20191);
or U24030 (N_24030,N_20836,N_20200);
xnor U24031 (N_24031,N_21415,N_19953);
nor U24032 (N_24032,N_20135,N_19197);
nor U24033 (N_24033,N_19982,N_19087);
nand U24034 (N_24034,N_20113,N_21284);
nor U24035 (N_24035,N_19481,N_20129);
nand U24036 (N_24036,N_20907,N_20615);
and U24037 (N_24037,N_19726,N_20727);
and U24038 (N_24038,N_21813,N_20005);
nand U24039 (N_24039,N_20517,N_21707);
xnor U24040 (N_24040,N_19836,N_20949);
nand U24041 (N_24041,N_21361,N_18788);
or U24042 (N_24042,N_21546,N_19290);
or U24043 (N_24043,N_19090,N_18989);
xor U24044 (N_24044,N_19977,N_19365);
nor U24045 (N_24045,N_19188,N_21693);
xor U24046 (N_24046,N_19051,N_19039);
and U24047 (N_24047,N_19635,N_20082);
and U24048 (N_24048,N_19828,N_21707);
nor U24049 (N_24049,N_21303,N_20637);
nor U24050 (N_24050,N_20926,N_19534);
or U24051 (N_24051,N_21035,N_21810);
and U24052 (N_24052,N_19492,N_20867);
and U24053 (N_24053,N_19488,N_19526);
and U24054 (N_24054,N_20773,N_19055);
or U24055 (N_24055,N_19302,N_20275);
xor U24056 (N_24056,N_21134,N_20121);
and U24057 (N_24057,N_19396,N_20263);
nand U24058 (N_24058,N_19595,N_19707);
or U24059 (N_24059,N_20499,N_21187);
xor U24060 (N_24060,N_19958,N_21586);
or U24061 (N_24061,N_18865,N_21408);
xnor U24062 (N_24062,N_20988,N_20398);
xnor U24063 (N_24063,N_19470,N_21867);
and U24064 (N_24064,N_20422,N_21207);
nand U24065 (N_24065,N_18972,N_19053);
or U24066 (N_24066,N_20186,N_19867);
nor U24067 (N_24067,N_19019,N_20263);
xor U24068 (N_24068,N_20405,N_20378);
xnor U24069 (N_24069,N_21663,N_21826);
nor U24070 (N_24070,N_19841,N_20464);
nand U24071 (N_24071,N_20855,N_19977);
nor U24072 (N_24072,N_20208,N_20758);
and U24073 (N_24073,N_20682,N_19499);
or U24074 (N_24074,N_20212,N_21281);
nor U24075 (N_24075,N_21167,N_20102);
and U24076 (N_24076,N_20445,N_21277);
nor U24077 (N_24077,N_19467,N_21364);
and U24078 (N_24078,N_19634,N_19658);
nand U24079 (N_24079,N_20015,N_19395);
and U24080 (N_24080,N_19142,N_20608);
nand U24081 (N_24081,N_21194,N_21788);
xor U24082 (N_24082,N_20789,N_19250);
or U24083 (N_24083,N_21219,N_19764);
and U24084 (N_24084,N_21277,N_18964);
nor U24085 (N_24085,N_21746,N_21388);
nand U24086 (N_24086,N_21265,N_19088);
nor U24087 (N_24087,N_19299,N_19524);
or U24088 (N_24088,N_19906,N_19381);
nor U24089 (N_24089,N_20876,N_19995);
xor U24090 (N_24090,N_20460,N_20849);
xnor U24091 (N_24091,N_19129,N_20102);
and U24092 (N_24092,N_20545,N_21062);
or U24093 (N_24093,N_21790,N_21698);
or U24094 (N_24094,N_20322,N_21211);
and U24095 (N_24095,N_19382,N_20716);
or U24096 (N_24096,N_19255,N_20007);
nand U24097 (N_24097,N_19903,N_19960);
nand U24098 (N_24098,N_19583,N_20226);
xor U24099 (N_24099,N_18995,N_19183);
nand U24100 (N_24100,N_19644,N_18988);
or U24101 (N_24101,N_21526,N_19135);
and U24102 (N_24102,N_20464,N_21227);
xnor U24103 (N_24103,N_21034,N_19085);
nor U24104 (N_24104,N_21567,N_21491);
xnor U24105 (N_24105,N_20086,N_21001);
or U24106 (N_24106,N_20326,N_19811);
and U24107 (N_24107,N_20227,N_18875);
nand U24108 (N_24108,N_21449,N_21668);
nor U24109 (N_24109,N_20935,N_21829);
and U24110 (N_24110,N_21127,N_21406);
nor U24111 (N_24111,N_20867,N_20524);
xnor U24112 (N_24112,N_19147,N_21815);
xnor U24113 (N_24113,N_20339,N_19269);
nor U24114 (N_24114,N_21384,N_21523);
and U24115 (N_24115,N_20720,N_19025);
xnor U24116 (N_24116,N_20962,N_19100);
or U24117 (N_24117,N_20262,N_18770);
or U24118 (N_24118,N_20651,N_19586);
nor U24119 (N_24119,N_21264,N_20541);
and U24120 (N_24120,N_19491,N_19271);
and U24121 (N_24121,N_20409,N_21236);
and U24122 (N_24122,N_21772,N_21025);
or U24123 (N_24123,N_19085,N_19840);
or U24124 (N_24124,N_20023,N_19637);
nand U24125 (N_24125,N_19996,N_19095);
nor U24126 (N_24126,N_19260,N_19436);
and U24127 (N_24127,N_19445,N_20395);
or U24128 (N_24128,N_20475,N_19708);
nor U24129 (N_24129,N_19626,N_19966);
or U24130 (N_24130,N_20771,N_21066);
nand U24131 (N_24131,N_19327,N_20606);
nor U24132 (N_24132,N_20057,N_20145);
nor U24133 (N_24133,N_21420,N_21066);
nor U24134 (N_24134,N_20144,N_21155);
and U24135 (N_24135,N_20780,N_19319);
or U24136 (N_24136,N_20493,N_18880);
nand U24137 (N_24137,N_20001,N_19976);
nand U24138 (N_24138,N_20866,N_21310);
or U24139 (N_24139,N_19280,N_19491);
and U24140 (N_24140,N_19289,N_18882);
and U24141 (N_24141,N_19831,N_19660);
xor U24142 (N_24142,N_20379,N_21372);
xor U24143 (N_24143,N_19887,N_20945);
nand U24144 (N_24144,N_19738,N_20054);
nor U24145 (N_24145,N_20517,N_19960);
and U24146 (N_24146,N_21406,N_19050);
or U24147 (N_24147,N_21430,N_19975);
or U24148 (N_24148,N_19710,N_19216);
or U24149 (N_24149,N_19495,N_19436);
and U24150 (N_24150,N_19165,N_19555);
and U24151 (N_24151,N_18876,N_20470);
xor U24152 (N_24152,N_21694,N_20548);
or U24153 (N_24153,N_19750,N_19097);
nand U24154 (N_24154,N_20655,N_21633);
nor U24155 (N_24155,N_18896,N_21798);
xor U24156 (N_24156,N_18906,N_20140);
or U24157 (N_24157,N_21782,N_19240);
xor U24158 (N_24158,N_20685,N_19226);
nor U24159 (N_24159,N_18875,N_20880);
nor U24160 (N_24160,N_20993,N_19475);
nor U24161 (N_24161,N_19278,N_19994);
xnor U24162 (N_24162,N_20103,N_19278);
xnor U24163 (N_24163,N_20010,N_20222);
nand U24164 (N_24164,N_18913,N_21865);
or U24165 (N_24165,N_19219,N_21669);
xor U24166 (N_24166,N_19555,N_18835);
and U24167 (N_24167,N_18752,N_20670);
nor U24168 (N_24168,N_19005,N_21593);
and U24169 (N_24169,N_19143,N_20017);
nand U24170 (N_24170,N_18824,N_19331);
xor U24171 (N_24171,N_18849,N_21256);
nor U24172 (N_24172,N_21533,N_20209);
xnor U24173 (N_24173,N_21198,N_20441);
nor U24174 (N_24174,N_21615,N_21802);
nand U24175 (N_24175,N_20101,N_20005);
and U24176 (N_24176,N_18826,N_20602);
nand U24177 (N_24177,N_19216,N_21291);
or U24178 (N_24178,N_21630,N_19565);
or U24179 (N_24179,N_20544,N_21686);
nor U24180 (N_24180,N_20146,N_19769);
and U24181 (N_24181,N_18915,N_18762);
or U24182 (N_24182,N_21466,N_21229);
nand U24183 (N_24183,N_21265,N_21648);
nor U24184 (N_24184,N_18839,N_19469);
and U24185 (N_24185,N_19402,N_20512);
or U24186 (N_24186,N_20524,N_20109);
nand U24187 (N_24187,N_20480,N_19566);
and U24188 (N_24188,N_20029,N_20283);
nand U24189 (N_24189,N_19187,N_21674);
nand U24190 (N_24190,N_19089,N_19583);
xor U24191 (N_24191,N_19333,N_20084);
nor U24192 (N_24192,N_19143,N_21651);
or U24193 (N_24193,N_19260,N_21536);
xor U24194 (N_24194,N_20226,N_19941);
and U24195 (N_24195,N_20549,N_20749);
nand U24196 (N_24196,N_20716,N_19339);
or U24197 (N_24197,N_19509,N_19504);
nor U24198 (N_24198,N_18773,N_20328);
or U24199 (N_24199,N_20148,N_21507);
and U24200 (N_24200,N_20049,N_19707);
and U24201 (N_24201,N_20376,N_21317);
or U24202 (N_24202,N_21123,N_20878);
or U24203 (N_24203,N_21183,N_18981);
nor U24204 (N_24204,N_21543,N_19147);
xor U24205 (N_24205,N_21049,N_20506);
and U24206 (N_24206,N_18900,N_21664);
nand U24207 (N_24207,N_21164,N_21820);
nor U24208 (N_24208,N_20376,N_20130);
nand U24209 (N_24209,N_20181,N_18826);
xnor U24210 (N_24210,N_21419,N_19754);
nand U24211 (N_24211,N_21062,N_21852);
nand U24212 (N_24212,N_21229,N_19479);
xnor U24213 (N_24213,N_19269,N_20277);
and U24214 (N_24214,N_20160,N_18752);
and U24215 (N_24215,N_19635,N_21227);
and U24216 (N_24216,N_20607,N_19287);
or U24217 (N_24217,N_21191,N_20414);
or U24218 (N_24218,N_19700,N_20545);
or U24219 (N_24219,N_19448,N_19151);
nor U24220 (N_24220,N_19478,N_20253);
or U24221 (N_24221,N_20740,N_20677);
xnor U24222 (N_24222,N_19704,N_20752);
or U24223 (N_24223,N_19255,N_19870);
xor U24224 (N_24224,N_19232,N_18861);
or U24225 (N_24225,N_20225,N_19222);
nor U24226 (N_24226,N_21614,N_20987);
and U24227 (N_24227,N_21160,N_19430);
and U24228 (N_24228,N_18859,N_20085);
nor U24229 (N_24229,N_21438,N_21451);
xor U24230 (N_24230,N_19700,N_21054);
xnor U24231 (N_24231,N_21146,N_20221);
and U24232 (N_24232,N_20595,N_19650);
and U24233 (N_24233,N_21494,N_19182);
nand U24234 (N_24234,N_19745,N_18821);
nand U24235 (N_24235,N_21814,N_18750);
nor U24236 (N_24236,N_21749,N_19865);
or U24237 (N_24237,N_19785,N_19798);
xor U24238 (N_24238,N_19668,N_19651);
or U24239 (N_24239,N_20587,N_20719);
nand U24240 (N_24240,N_20556,N_20287);
xor U24241 (N_24241,N_20779,N_20053);
nand U24242 (N_24242,N_20032,N_20386);
or U24243 (N_24243,N_21307,N_18810);
and U24244 (N_24244,N_21167,N_19478);
or U24245 (N_24245,N_21666,N_18914);
or U24246 (N_24246,N_20209,N_21703);
or U24247 (N_24247,N_21508,N_20914);
xor U24248 (N_24248,N_20964,N_21691);
nor U24249 (N_24249,N_21179,N_21113);
nand U24250 (N_24250,N_20147,N_19960);
nor U24251 (N_24251,N_19389,N_20331);
and U24252 (N_24252,N_19190,N_21450);
and U24253 (N_24253,N_21762,N_19876);
or U24254 (N_24254,N_20704,N_20874);
nand U24255 (N_24255,N_18887,N_20803);
or U24256 (N_24256,N_20706,N_19453);
and U24257 (N_24257,N_21574,N_19293);
xnor U24258 (N_24258,N_21669,N_20472);
xnor U24259 (N_24259,N_21564,N_19804);
or U24260 (N_24260,N_18897,N_20623);
nor U24261 (N_24261,N_21218,N_21081);
or U24262 (N_24262,N_20041,N_19096);
xor U24263 (N_24263,N_18839,N_20612);
nand U24264 (N_24264,N_21243,N_21659);
nor U24265 (N_24265,N_19009,N_21357);
nand U24266 (N_24266,N_19603,N_21247);
xor U24267 (N_24267,N_20011,N_19703);
nor U24268 (N_24268,N_19292,N_21159);
nand U24269 (N_24269,N_19616,N_19019);
or U24270 (N_24270,N_20956,N_20256);
or U24271 (N_24271,N_21513,N_19208);
nand U24272 (N_24272,N_19259,N_21528);
or U24273 (N_24273,N_19614,N_20889);
xnor U24274 (N_24274,N_18884,N_19918);
nand U24275 (N_24275,N_19871,N_21028);
nor U24276 (N_24276,N_19579,N_20495);
nand U24277 (N_24277,N_21626,N_20218);
and U24278 (N_24278,N_20147,N_21532);
and U24279 (N_24279,N_21746,N_20669);
nand U24280 (N_24280,N_20831,N_20995);
and U24281 (N_24281,N_20022,N_19608);
nor U24282 (N_24282,N_19284,N_20493);
and U24283 (N_24283,N_20405,N_19378);
nand U24284 (N_24284,N_20990,N_20692);
or U24285 (N_24285,N_21787,N_20336);
and U24286 (N_24286,N_19635,N_20335);
nor U24287 (N_24287,N_20678,N_20941);
or U24288 (N_24288,N_19540,N_20974);
nand U24289 (N_24289,N_19824,N_21749);
xnor U24290 (N_24290,N_20225,N_19306);
and U24291 (N_24291,N_21869,N_18989);
nand U24292 (N_24292,N_21596,N_21059);
nor U24293 (N_24293,N_20588,N_21667);
or U24294 (N_24294,N_20782,N_19201);
nand U24295 (N_24295,N_20145,N_21269);
and U24296 (N_24296,N_20748,N_20276);
nor U24297 (N_24297,N_19628,N_20921);
and U24298 (N_24298,N_18987,N_20531);
nor U24299 (N_24299,N_19230,N_21770);
and U24300 (N_24300,N_20541,N_20225);
or U24301 (N_24301,N_21193,N_20011);
and U24302 (N_24302,N_20662,N_19034);
nor U24303 (N_24303,N_21414,N_20337);
and U24304 (N_24304,N_19780,N_19160);
xor U24305 (N_24305,N_20375,N_19030);
or U24306 (N_24306,N_19103,N_21663);
nor U24307 (N_24307,N_18875,N_19156);
xor U24308 (N_24308,N_19810,N_20491);
nand U24309 (N_24309,N_20650,N_20207);
nor U24310 (N_24310,N_21574,N_19397);
nor U24311 (N_24311,N_21748,N_20700);
or U24312 (N_24312,N_20109,N_20451);
and U24313 (N_24313,N_21699,N_21590);
or U24314 (N_24314,N_21006,N_19139);
or U24315 (N_24315,N_19395,N_21874);
or U24316 (N_24316,N_19297,N_21467);
nand U24317 (N_24317,N_20537,N_21116);
xnor U24318 (N_24318,N_20155,N_20800);
or U24319 (N_24319,N_20915,N_21159);
nor U24320 (N_24320,N_20143,N_21292);
and U24321 (N_24321,N_20644,N_19520);
and U24322 (N_24322,N_19096,N_20305);
nand U24323 (N_24323,N_18770,N_21196);
nand U24324 (N_24324,N_19116,N_20567);
nand U24325 (N_24325,N_20058,N_20783);
nor U24326 (N_24326,N_18854,N_21321);
nand U24327 (N_24327,N_20098,N_19592);
and U24328 (N_24328,N_18986,N_18935);
nand U24329 (N_24329,N_21719,N_19180);
or U24330 (N_24330,N_19485,N_21012);
nand U24331 (N_24331,N_20693,N_20968);
nand U24332 (N_24332,N_20497,N_20823);
xnor U24333 (N_24333,N_21685,N_18922);
nand U24334 (N_24334,N_21508,N_20696);
nand U24335 (N_24335,N_20094,N_20710);
or U24336 (N_24336,N_21822,N_20278);
nand U24337 (N_24337,N_18799,N_21061);
nor U24338 (N_24338,N_18751,N_21047);
or U24339 (N_24339,N_21759,N_20662);
or U24340 (N_24340,N_20913,N_21837);
nand U24341 (N_24341,N_19444,N_21707);
xnor U24342 (N_24342,N_19345,N_20278);
nand U24343 (N_24343,N_19404,N_19992);
or U24344 (N_24344,N_21175,N_19655);
xor U24345 (N_24345,N_20483,N_19653);
xnor U24346 (N_24346,N_21545,N_20257);
and U24347 (N_24347,N_19473,N_21855);
or U24348 (N_24348,N_21687,N_19219);
and U24349 (N_24349,N_19018,N_20670);
xnor U24350 (N_24350,N_20666,N_21857);
or U24351 (N_24351,N_20068,N_19291);
nand U24352 (N_24352,N_19741,N_20951);
nor U24353 (N_24353,N_20153,N_21396);
and U24354 (N_24354,N_21533,N_19475);
or U24355 (N_24355,N_19363,N_20633);
xor U24356 (N_24356,N_19753,N_20961);
or U24357 (N_24357,N_21225,N_20987);
nand U24358 (N_24358,N_21673,N_21242);
xor U24359 (N_24359,N_21855,N_20380);
nor U24360 (N_24360,N_19899,N_18852);
xnor U24361 (N_24361,N_21491,N_20676);
nand U24362 (N_24362,N_19339,N_20039);
nor U24363 (N_24363,N_21397,N_18833);
and U24364 (N_24364,N_21261,N_20318);
nor U24365 (N_24365,N_20794,N_20778);
and U24366 (N_24366,N_19730,N_20834);
nand U24367 (N_24367,N_21004,N_18926);
nand U24368 (N_24368,N_18884,N_20119);
nor U24369 (N_24369,N_21266,N_19229);
nand U24370 (N_24370,N_20985,N_18764);
nor U24371 (N_24371,N_18890,N_20793);
nor U24372 (N_24372,N_19579,N_20788);
and U24373 (N_24373,N_19279,N_19741);
nor U24374 (N_24374,N_19989,N_20928);
and U24375 (N_24375,N_20206,N_20842);
or U24376 (N_24376,N_19915,N_19892);
nand U24377 (N_24377,N_19842,N_19985);
or U24378 (N_24378,N_19801,N_19183);
xnor U24379 (N_24379,N_18987,N_20896);
or U24380 (N_24380,N_21681,N_19502);
and U24381 (N_24381,N_21162,N_18750);
nand U24382 (N_24382,N_19736,N_19503);
and U24383 (N_24383,N_20269,N_20809);
nand U24384 (N_24384,N_21609,N_19137);
xor U24385 (N_24385,N_18927,N_18961);
and U24386 (N_24386,N_21687,N_20199);
xor U24387 (N_24387,N_20523,N_20584);
xor U24388 (N_24388,N_21722,N_21461);
and U24389 (N_24389,N_20464,N_21531);
xnor U24390 (N_24390,N_19189,N_20515);
or U24391 (N_24391,N_20176,N_19272);
and U24392 (N_24392,N_18882,N_20543);
or U24393 (N_24393,N_21424,N_20311);
nand U24394 (N_24394,N_20169,N_21649);
or U24395 (N_24395,N_19850,N_20071);
or U24396 (N_24396,N_20933,N_20150);
or U24397 (N_24397,N_21373,N_18976);
nand U24398 (N_24398,N_19661,N_20729);
nor U24399 (N_24399,N_21643,N_19115);
nand U24400 (N_24400,N_21547,N_20627);
xnor U24401 (N_24401,N_20593,N_21077);
and U24402 (N_24402,N_20964,N_18924);
nand U24403 (N_24403,N_20638,N_20021);
nand U24404 (N_24404,N_20413,N_19159);
nor U24405 (N_24405,N_19929,N_20653);
xor U24406 (N_24406,N_19468,N_20962);
xor U24407 (N_24407,N_21505,N_19027);
nand U24408 (N_24408,N_21816,N_21662);
and U24409 (N_24409,N_21631,N_19558);
or U24410 (N_24410,N_20940,N_19255);
and U24411 (N_24411,N_19148,N_19379);
or U24412 (N_24412,N_18812,N_21505);
nor U24413 (N_24413,N_18826,N_18863);
nand U24414 (N_24414,N_20501,N_20178);
xor U24415 (N_24415,N_19113,N_20967);
and U24416 (N_24416,N_19156,N_21292);
or U24417 (N_24417,N_20964,N_21138);
and U24418 (N_24418,N_19217,N_19204);
or U24419 (N_24419,N_19510,N_19737);
or U24420 (N_24420,N_20994,N_19941);
nor U24421 (N_24421,N_19246,N_21826);
xnor U24422 (N_24422,N_19957,N_19365);
or U24423 (N_24423,N_19623,N_21531);
and U24424 (N_24424,N_19633,N_20687);
or U24425 (N_24425,N_20113,N_20510);
nand U24426 (N_24426,N_20101,N_20927);
or U24427 (N_24427,N_21605,N_20540);
nand U24428 (N_24428,N_21570,N_18774);
xor U24429 (N_24429,N_20799,N_20237);
and U24430 (N_24430,N_21160,N_20592);
xnor U24431 (N_24431,N_19125,N_19035);
nor U24432 (N_24432,N_20541,N_19311);
nor U24433 (N_24433,N_19830,N_21791);
xor U24434 (N_24434,N_19922,N_21251);
nor U24435 (N_24435,N_20001,N_21776);
nor U24436 (N_24436,N_20282,N_21157);
nor U24437 (N_24437,N_21544,N_21466);
xnor U24438 (N_24438,N_20697,N_19809);
xnor U24439 (N_24439,N_21092,N_20555);
nor U24440 (N_24440,N_19326,N_20404);
nor U24441 (N_24441,N_21318,N_20320);
and U24442 (N_24442,N_21292,N_18990);
nor U24443 (N_24443,N_19308,N_19658);
xor U24444 (N_24444,N_18936,N_19383);
nor U24445 (N_24445,N_20595,N_20090);
xor U24446 (N_24446,N_19528,N_20023);
nor U24447 (N_24447,N_20741,N_20187);
and U24448 (N_24448,N_18804,N_20467);
or U24449 (N_24449,N_19542,N_20857);
and U24450 (N_24450,N_20620,N_21363);
or U24451 (N_24451,N_19950,N_20114);
nand U24452 (N_24452,N_21396,N_19782);
nor U24453 (N_24453,N_19815,N_19139);
xnor U24454 (N_24454,N_19887,N_20914);
nand U24455 (N_24455,N_21698,N_20634);
and U24456 (N_24456,N_19841,N_18941);
nand U24457 (N_24457,N_19334,N_20803);
nand U24458 (N_24458,N_21068,N_21077);
xor U24459 (N_24459,N_21123,N_21116);
nor U24460 (N_24460,N_19281,N_21461);
xnor U24461 (N_24461,N_20443,N_19777);
xnor U24462 (N_24462,N_21761,N_21107);
nor U24463 (N_24463,N_21336,N_19770);
or U24464 (N_24464,N_21632,N_19102);
and U24465 (N_24465,N_21161,N_20576);
nor U24466 (N_24466,N_20803,N_20365);
nor U24467 (N_24467,N_19338,N_21621);
nor U24468 (N_24468,N_21699,N_18816);
or U24469 (N_24469,N_21627,N_20394);
and U24470 (N_24470,N_20656,N_19886);
nor U24471 (N_24471,N_19633,N_19723);
and U24472 (N_24472,N_21734,N_20523);
xor U24473 (N_24473,N_21143,N_19728);
xor U24474 (N_24474,N_21713,N_21262);
and U24475 (N_24475,N_19187,N_19452);
xnor U24476 (N_24476,N_20743,N_20480);
xnor U24477 (N_24477,N_20310,N_18893);
and U24478 (N_24478,N_21293,N_19350);
nand U24479 (N_24479,N_21007,N_20071);
or U24480 (N_24480,N_19556,N_19264);
and U24481 (N_24481,N_20080,N_21316);
xnor U24482 (N_24482,N_21242,N_21352);
or U24483 (N_24483,N_20670,N_21210);
nor U24484 (N_24484,N_20279,N_21379);
or U24485 (N_24485,N_19129,N_21507);
and U24486 (N_24486,N_18983,N_18768);
or U24487 (N_24487,N_21058,N_19551);
nand U24488 (N_24488,N_21584,N_20238);
nor U24489 (N_24489,N_18994,N_20394);
and U24490 (N_24490,N_20796,N_18923);
and U24491 (N_24491,N_18951,N_20011);
xnor U24492 (N_24492,N_21297,N_21295);
or U24493 (N_24493,N_21165,N_21725);
nor U24494 (N_24494,N_20201,N_18804);
nor U24495 (N_24495,N_18869,N_21401);
nand U24496 (N_24496,N_20897,N_21764);
nor U24497 (N_24497,N_19842,N_20072);
nand U24498 (N_24498,N_20903,N_21809);
nor U24499 (N_24499,N_19136,N_20939);
nor U24500 (N_24500,N_21743,N_20589);
nor U24501 (N_24501,N_18945,N_21600);
or U24502 (N_24502,N_18867,N_21727);
and U24503 (N_24503,N_21595,N_21290);
xor U24504 (N_24504,N_20232,N_20847);
xor U24505 (N_24505,N_19039,N_19266);
nor U24506 (N_24506,N_21458,N_21572);
or U24507 (N_24507,N_21109,N_18954);
nor U24508 (N_24508,N_19613,N_21762);
nor U24509 (N_24509,N_21178,N_20436);
nand U24510 (N_24510,N_21601,N_20120);
or U24511 (N_24511,N_21734,N_20348);
xnor U24512 (N_24512,N_19740,N_21421);
or U24513 (N_24513,N_20275,N_19598);
or U24514 (N_24514,N_21327,N_19538);
xor U24515 (N_24515,N_20048,N_20012);
nor U24516 (N_24516,N_19669,N_20016);
nor U24517 (N_24517,N_21625,N_20862);
or U24518 (N_24518,N_20790,N_21513);
nand U24519 (N_24519,N_19227,N_20238);
nor U24520 (N_24520,N_20777,N_19079);
xor U24521 (N_24521,N_21017,N_19567);
nand U24522 (N_24522,N_21333,N_19820);
xnor U24523 (N_24523,N_20538,N_20027);
or U24524 (N_24524,N_20956,N_18954);
and U24525 (N_24525,N_20133,N_19206);
nand U24526 (N_24526,N_18906,N_21873);
xnor U24527 (N_24527,N_19070,N_20044);
xnor U24528 (N_24528,N_21634,N_21020);
nor U24529 (N_24529,N_18780,N_20347);
and U24530 (N_24530,N_18849,N_19774);
and U24531 (N_24531,N_20443,N_20907);
xor U24532 (N_24532,N_19934,N_21439);
and U24533 (N_24533,N_19015,N_19727);
nor U24534 (N_24534,N_21429,N_21329);
nor U24535 (N_24535,N_20397,N_18944);
or U24536 (N_24536,N_19183,N_19616);
xor U24537 (N_24537,N_18840,N_18955);
and U24538 (N_24538,N_21467,N_21077);
or U24539 (N_24539,N_19437,N_19188);
or U24540 (N_24540,N_20661,N_19925);
or U24541 (N_24541,N_21506,N_19745);
and U24542 (N_24542,N_20973,N_19839);
nand U24543 (N_24543,N_19179,N_20022);
xor U24544 (N_24544,N_20782,N_21653);
xnor U24545 (N_24545,N_19124,N_20285);
nand U24546 (N_24546,N_19894,N_19387);
nor U24547 (N_24547,N_20390,N_20339);
xnor U24548 (N_24548,N_19797,N_20924);
and U24549 (N_24549,N_19631,N_18883);
xor U24550 (N_24550,N_19436,N_19075);
nand U24551 (N_24551,N_19804,N_18875);
nor U24552 (N_24552,N_19504,N_19616);
nor U24553 (N_24553,N_21423,N_19824);
xnor U24554 (N_24554,N_19300,N_19924);
xnor U24555 (N_24555,N_19067,N_19811);
nand U24556 (N_24556,N_19497,N_19796);
nor U24557 (N_24557,N_21835,N_21495);
and U24558 (N_24558,N_19306,N_21230);
and U24559 (N_24559,N_21829,N_19451);
and U24560 (N_24560,N_21440,N_19435);
and U24561 (N_24561,N_19080,N_18879);
xor U24562 (N_24562,N_20121,N_20037);
and U24563 (N_24563,N_20550,N_19627);
and U24564 (N_24564,N_19624,N_18843);
or U24565 (N_24565,N_19187,N_21559);
nand U24566 (N_24566,N_19108,N_21028);
xnor U24567 (N_24567,N_19073,N_21644);
or U24568 (N_24568,N_21668,N_21085);
and U24569 (N_24569,N_20106,N_21355);
nand U24570 (N_24570,N_21355,N_19611);
nand U24571 (N_24571,N_18957,N_20988);
xor U24572 (N_24572,N_19914,N_19449);
and U24573 (N_24573,N_19545,N_18959);
or U24574 (N_24574,N_18782,N_18988);
or U24575 (N_24575,N_20625,N_20899);
nor U24576 (N_24576,N_21037,N_20673);
nor U24577 (N_24577,N_20682,N_20113);
xor U24578 (N_24578,N_20048,N_20142);
or U24579 (N_24579,N_20929,N_18999);
xnor U24580 (N_24580,N_20602,N_18769);
xor U24581 (N_24581,N_19935,N_19305);
nand U24582 (N_24582,N_19257,N_21063);
and U24583 (N_24583,N_19145,N_20349);
xor U24584 (N_24584,N_18874,N_19623);
or U24585 (N_24585,N_19921,N_19273);
xor U24586 (N_24586,N_19998,N_21005);
xnor U24587 (N_24587,N_20574,N_19265);
nand U24588 (N_24588,N_21865,N_19096);
or U24589 (N_24589,N_19831,N_20711);
nand U24590 (N_24590,N_21738,N_19764);
or U24591 (N_24591,N_20355,N_19017);
or U24592 (N_24592,N_20782,N_20425);
and U24593 (N_24593,N_20344,N_19575);
nand U24594 (N_24594,N_18972,N_19688);
xor U24595 (N_24595,N_19922,N_19420);
and U24596 (N_24596,N_18878,N_21323);
xor U24597 (N_24597,N_19786,N_21255);
xnor U24598 (N_24598,N_20332,N_18856);
or U24599 (N_24599,N_19988,N_20691);
or U24600 (N_24600,N_21049,N_19292);
or U24601 (N_24601,N_20499,N_20767);
or U24602 (N_24602,N_20498,N_19991);
nand U24603 (N_24603,N_20415,N_19229);
and U24604 (N_24604,N_19833,N_20020);
nand U24605 (N_24605,N_19664,N_19595);
and U24606 (N_24606,N_18897,N_21050);
nand U24607 (N_24607,N_20361,N_19798);
nor U24608 (N_24608,N_20287,N_21673);
nor U24609 (N_24609,N_21659,N_21442);
or U24610 (N_24610,N_21685,N_19914);
nor U24611 (N_24611,N_18761,N_21816);
or U24612 (N_24612,N_19261,N_19644);
nand U24613 (N_24613,N_19166,N_21160);
and U24614 (N_24614,N_20737,N_20174);
xnor U24615 (N_24615,N_21069,N_18894);
nand U24616 (N_24616,N_21428,N_21305);
nor U24617 (N_24617,N_21141,N_19665);
and U24618 (N_24618,N_20156,N_19951);
xor U24619 (N_24619,N_21741,N_21114);
or U24620 (N_24620,N_21318,N_20393);
nor U24621 (N_24621,N_19360,N_19814);
nor U24622 (N_24622,N_20391,N_20540);
and U24623 (N_24623,N_19717,N_20567);
or U24624 (N_24624,N_21805,N_20226);
nor U24625 (N_24625,N_19648,N_20339);
xnor U24626 (N_24626,N_19123,N_21059);
and U24627 (N_24627,N_19639,N_18854);
or U24628 (N_24628,N_21818,N_20115);
or U24629 (N_24629,N_20274,N_21287);
and U24630 (N_24630,N_20489,N_21334);
nand U24631 (N_24631,N_21528,N_21308);
xor U24632 (N_24632,N_20878,N_21402);
nand U24633 (N_24633,N_20789,N_21823);
nand U24634 (N_24634,N_19834,N_19383);
or U24635 (N_24635,N_21804,N_20391);
or U24636 (N_24636,N_19644,N_18880);
nor U24637 (N_24637,N_20578,N_18991);
nand U24638 (N_24638,N_19515,N_19130);
nor U24639 (N_24639,N_20806,N_21580);
nand U24640 (N_24640,N_19730,N_20600);
and U24641 (N_24641,N_19665,N_20632);
or U24642 (N_24642,N_21314,N_20534);
and U24643 (N_24643,N_20128,N_18850);
or U24644 (N_24644,N_20458,N_21182);
xor U24645 (N_24645,N_21415,N_20391);
nand U24646 (N_24646,N_19397,N_19729);
nand U24647 (N_24647,N_19401,N_20348);
nand U24648 (N_24648,N_21571,N_20530);
or U24649 (N_24649,N_21174,N_19672);
and U24650 (N_24650,N_20390,N_20420);
or U24651 (N_24651,N_21202,N_19545);
nor U24652 (N_24652,N_21305,N_21010);
xnor U24653 (N_24653,N_18770,N_20070);
nand U24654 (N_24654,N_21711,N_19823);
nand U24655 (N_24655,N_18989,N_20262);
nand U24656 (N_24656,N_21782,N_19216);
and U24657 (N_24657,N_20439,N_20410);
or U24658 (N_24658,N_21353,N_21575);
nor U24659 (N_24659,N_19617,N_19024);
and U24660 (N_24660,N_21868,N_19189);
xor U24661 (N_24661,N_20269,N_20490);
and U24662 (N_24662,N_19038,N_19549);
and U24663 (N_24663,N_20163,N_19938);
and U24664 (N_24664,N_20178,N_19983);
or U24665 (N_24665,N_21257,N_19484);
xor U24666 (N_24666,N_20021,N_20892);
or U24667 (N_24667,N_19994,N_19557);
and U24668 (N_24668,N_21196,N_21688);
and U24669 (N_24669,N_20226,N_19766);
nor U24670 (N_24670,N_21401,N_20245);
and U24671 (N_24671,N_19940,N_20691);
xor U24672 (N_24672,N_21749,N_21781);
xor U24673 (N_24673,N_20726,N_20653);
nand U24674 (N_24674,N_19860,N_21647);
xor U24675 (N_24675,N_20498,N_21116);
nand U24676 (N_24676,N_21107,N_18926);
or U24677 (N_24677,N_19476,N_21289);
or U24678 (N_24678,N_18757,N_20717);
and U24679 (N_24679,N_18944,N_19278);
nor U24680 (N_24680,N_20018,N_18763);
nand U24681 (N_24681,N_21464,N_21805);
nor U24682 (N_24682,N_20934,N_20506);
or U24683 (N_24683,N_20350,N_21673);
nor U24684 (N_24684,N_19516,N_18829);
nor U24685 (N_24685,N_21157,N_21084);
or U24686 (N_24686,N_19549,N_21760);
xor U24687 (N_24687,N_19773,N_20484);
and U24688 (N_24688,N_19956,N_19989);
xor U24689 (N_24689,N_21636,N_20915);
xnor U24690 (N_24690,N_20130,N_19747);
nand U24691 (N_24691,N_19443,N_21636);
and U24692 (N_24692,N_20644,N_20283);
and U24693 (N_24693,N_20118,N_20854);
and U24694 (N_24694,N_20690,N_20165);
and U24695 (N_24695,N_19844,N_21280);
or U24696 (N_24696,N_20988,N_20192);
xor U24697 (N_24697,N_21721,N_20397);
and U24698 (N_24698,N_20335,N_19174);
or U24699 (N_24699,N_20631,N_19319);
and U24700 (N_24700,N_19081,N_19853);
and U24701 (N_24701,N_21870,N_19334);
nor U24702 (N_24702,N_21349,N_20583);
or U24703 (N_24703,N_21738,N_20767);
and U24704 (N_24704,N_21620,N_19462);
nand U24705 (N_24705,N_19573,N_21861);
or U24706 (N_24706,N_20251,N_19753);
or U24707 (N_24707,N_20643,N_18795);
xor U24708 (N_24708,N_21316,N_21737);
and U24709 (N_24709,N_20949,N_19971);
nand U24710 (N_24710,N_21363,N_20462);
nand U24711 (N_24711,N_21668,N_21830);
or U24712 (N_24712,N_20233,N_21499);
nor U24713 (N_24713,N_20938,N_19384);
nand U24714 (N_24714,N_19960,N_21106);
nor U24715 (N_24715,N_21471,N_21552);
or U24716 (N_24716,N_18756,N_20708);
nand U24717 (N_24717,N_21863,N_21765);
and U24718 (N_24718,N_20210,N_20098);
nand U24719 (N_24719,N_21575,N_20604);
nand U24720 (N_24720,N_19019,N_20194);
or U24721 (N_24721,N_19802,N_20301);
nand U24722 (N_24722,N_19931,N_21648);
nor U24723 (N_24723,N_18781,N_20185);
or U24724 (N_24724,N_20704,N_19400);
and U24725 (N_24725,N_21357,N_20156);
and U24726 (N_24726,N_20247,N_21342);
and U24727 (N_24727,N_19691,N_20651);
xnor U24728 (N_24728,N_20007,N_19283);
nand U24729 (N_24729,N_19454,N_21118);
or U24730 (N_24730,N_21626,N_19174);
nor U24731 (N_24731,N_21228,N_21254);
nand U24732 (N_24732,N_19980,N_20620);
or U24733 (N_24733,N_19889,N_20503);
nor U24734 (N_24734,N_20186,N_19955);
and U24735 (N_24735,N_19597,N_20452);
or U24736 (N_24736,N_20884,N_19851);
or U24737 (N_24737,N_19359,N_19976);
xor U24738 (N_24738,N_20105,N_21332);
nor U24739 (N_24739,N_21206,N_19546);
and U24740 (N_24740,N_21330,N_18986);
and U24741 (N_24741,N_20892,N_19466);
nand U24742 (N_24742,N_20561,N_20329);
nand U24743 (N_24743,N_19249,N_21426);
xnor U24744 (N_24744,N_20566,N_20309);
and U24745 (N_24745,N_18996,N_21643);
or U24746 (N_24746,N_21533,N_19267);
nor U24747 (N_24747,N_20307,N_20433);
nand U24748 (N_24748,N_20834,N_19839);
xor U24749 (N_24749,N_21517,N_20230);
or U24750 (N_24750,N_20419,N_19213);
and U24751 (N_24751,N_21295,N_20636);
and U24752 (N_24752,N_19773,N_19522);
and U24753 (N_24753,N_19690,N_20835);
nor U24754 (N_24754,N_21820,N_19868);
nand U24755 (N_24755,N_19884,N_19376);
and U24756 (N_24756,N_19502,N_19886);
or U24757 (N_24757,N_21463,N_20638);
and U24758 (N_24758,N_21272,N_20984);
or U24759 (N_24759,N_18870,N_19118);
or U24760 (N_24760,N_20931,N_19898);
or U24761 (N_24761,N_18775,N_20197);
nor U24762 (N_24762,N_20445,N_18903);
nand U24763 (N_24763,N_19012,N_20543);
nand U24764 (N_24764,N_21257,N_19917);
xor U24765 (N_24765,N_21433,N_21140);
and U24766 (N_24766,N_19379,N_20808);
xor U24767 (N_24767,N_21523,N_20282);
nand U24768 (N_24768,N_20511,N_21201);
or U24769 (N_24769,N_21752,N_21807);
or U24770 (N_24770,N_21788,N_20989);
nand U24771 (N_24771,N_20889,N_20329);
nand U24772 (N_24772,N_20440,N_21572);
nor U24773 (N_24773,N_20822,N_19079);
xor U24774 (N_24774,N_21772,N_21239);
nand U24775 (N_24775,N_19552,N_18788);
nor U24776 (N_24776,N_18752,N_20347);
nor U24777 (N_24777,N_21319,N_19693);
nand U24778 (N_24778,N_19214,N_21014);
xor U24779 (N_24779,N_21568,N_21121);
nand U24780 (N_24780,N_19966,N_19763);
and U24781 (N_24781,N_20050,N_21821);
or U24782 (N_24782,N_21320,N_21772);
xnor U24783 (N_24783,N_20409,N_19152);
xnor U24784 (N_24784,N_21542,N_21454);
xnor U24785 (N_24785,N_19100,N_20928);
or U24786 (N_24786,N_20543,N_19311);
nand U24787 (N_24787,N_21320,N_21303);
nor U24788 (N_24788,N_20588,N_19222);
or U24789 (N_24789,N_20216,N_19523);
or U24790 (N_24790,N_20642,N_18851);
nand U24791 (N_24791,N_21817,N_20905);
nor U24792 (N_24792,N_19949,N_21569);
nor U24793 (N_24793,N_18955,N_20817);
and U24794 (N_24794,N_21638,N_21478);
nor U24795 (N_24795,N_19663,N_20355);
or U24796 (N_24796,N_20841,N_20142);
xnor U24797 (N_24797,N_21644,N_19579);
and U24798 (N_24798,N_20836,N_19514);
or U24799 (N_24799,N_21073,N_19709);
xnor U24800 (N_24800,N_21776,N_20538);
xor U24801 (N_24801,N_21749,N_21823);
nand U24802 (N_24802,N_20552,N_18964);
nand U24803 (N_24803,N_21845,N_20178);
xnor U24804 (N_24804,N_19355,N_19230);
nand U24805 (N_24805,N_20394,N_20996);
xnor U24806 (N_24806,N_20004,N_21829);
nand U24807 (N_24807,N_19473,N_19974);
xnor U24808 (N_24808,N_20241,N_18751);
and U24809 (N_24809,N_21144,N_19175);
nor U24810 (N_24810,N_20006,N_19756);
nand U24811 (N_24811,N_20956,N_21690);
nor U24812 (N_24812,N_20340,N_19546);
nand U24813 (N_24813,N_19096,N_21829);
and U24814 (N_24814,N_21572,N_21132);
nand U24815 (N_24815,N_20785,N_18960);
and U24816 (N_24816,N_19527,N_21772);
nor U24817 (N_24817,N_20206,N_20064);
and U24818 (N_24818,N_19030,N_18931);
xor U24819 (N_24819,N_20519,N_20779);
nor U24820 (N_24820,N_19729,N_19147);
xor U24821 (N_24821,N_18753,N_20855);
nand U24822 (N_24822,N_20764,N_21203);
nor U24823 (N_24823,N_20235,N_21461);
and U24824 (N_24824,N_21297,N_20626);
nor U24825 (N_24825,N_21722,N_21333);
or U24826 (N_24826,N_20664,N_18810);
nand U24827 (N_24827,N_20091,N_21253);
nor U24828 (N_24828,N_19046,N_20724);
xor U24829 (N_24829,N_20766,N_19239);
xor U24830 (N_24830,N_20318,N_19854);
and U24831 (N_24831,N_19927,N_19515);
or U24832 (N_24832,N_21468,N_18826);
nand U24833 (N_24833,N_20690,N_19474);
or U24834 (N_24834,N_20674,N_21823);
or U24835 (N_24835,N_18787,N_21199);
or U24836 (N_24836,N_19397,N_20345);
and U24837 (N_24837,N_19836,N_21320);
and U24838 (N_24838,N_20481,N_19312);
or U24839 (N_24839,N_19826,N_19328);
nand U24840 (N_24840,N_20398,N_19246);
xor U24841 (N_24841,N_19383,N_21150);
or U24842 (N_24842,N_20410,N_18953);
nor U24843 (N_24843,N_20269,N_21781);
and U24844 (N_24844,N_20596,N_20152);
xnor U24845 (N_24845,N_19617,N_19498);
nand U24846 (N_24846,N_21607,N_19454);
nand U24847 (N_24847,N_20568,N_19676);
xor U24848 (N_24848,N_18932,N_18993);
nand U24849 (N_24849,N_21817,N_20999);
and U24850 (N_24850,N_19854,N_19484);
nand U24851 (N_24851,N_19200,N_20856);
xor U24852 (N_24852,N_20460,N_19987);
nand U24853 (N_24853,N_18944,N_19693);
nand U24854 (N_24854,N_19072,N_21658);
and U24855 (N_24855,N_19062,N_19747);
nand U24856 (N_24856,N_20561,N_19525);
and U24857 (N_24857,N_19374,N_19341);
and U24858 (N_24858,N_20821,N_20399);
nand U24859 (N_24859,N_21358,N_21667);
nor U24860 (N_24860,N_20289,N_19329);
nor U24861 (N_24861,N_20551,N_20376);
or U24862 (N_24862,N_19002,N_20472);
or U24863 (N_24863,N_20636,N_18885);
and U24864 (N_24864,N_21222,N_19989);
and U24865 (N_24865,N_20012,N_20270);
and U24866 (N_24866,N_20321,N_19256);
nor U24867 (N_24867,N_18922,N_20158);
xnor U24868 (N_24868,N_18967,N_20214);
nand U24869 (N_24869,N_20972,N_19931);
xor U24870 (N_24870,N_19737,N_21462);
xor U24871 (N_24871,N_19218,N_20311);
and U24872 (N_24872,N_18955,N_21238);
nand U24873 (N_24873,N_19288,N_20587);
xnor U24874 (N_24874,N_19364,N_19008);
and U24875 (N_24875,N_20148,N_21061);
and U24876 (N_24876,N_19229,N_21292);
xnor U24877 (N_24877,N_19104,N_19988);
and U24878 (N_24878,N_21367,N_18997);
and U24879 (N_24879,N_19910,N_21109);
nor U24880 (N_24880,N_20740,N_21734);
and U24881 (N_24881,N_19510,N_21801);
nor U24882 (N_24882,N_19105,N_20185);
nand U24883 (N_24883,N_19258,N_19416);
xnor U24884 (N_24884,N_18832,N_19033);
nand U24885 (N_24885,N_19183,N_20006);
nand U24886 (N_24886,N_20064,N_19287);
nor U24887 (N_24887,N_19220,N_21623);
and U24888 (N_24888,N_20826,N_18858);
nand U24889 (N_24889,N_19582,N_19732);
and U24890 (N_24890,N_19717,N_21868);
or U24891 (N_24891,N_20671,N_19533);
and U24892 (N_24892,N_20197,N_20543);
xnor U24893 (N_24893,N_20112,N_21362);
and U24894 (N_24894,N_20221,N_21817);
and U24895 (N_24895,N_19884,N_18880);
or U24896 (N_24896,N_21008,N_20219);
nor U24897 (N_24897,N_20062,N_20619);
nand U24898 (N_24898,N_19552,N_19443);
nor U24899 (N_24899,N_19050,N_21116);
nor U24900 (N_24900,N_20989,N_20688);
and U24901 (N_24901,N_19948,N_20057);
or U24902 (N_24902,N_21755,N_21036);
nor U24903 (N_24903,N_21865,N_21292);
nor U24904 (N_24904,N_20379,N_19948);
nor U24905 (N_24905,N_21757,N_20111);
xnor U24906 (N_24906,N_21431,N_19179);
nor U24907 (N_24907,N_19481,N_18889);
xor U24908 (N_24908,N_19146,N_19857);
xor U24909 (N_24909,N_20157,N_20311);
and U24910 (N_24910,N_21523,N_20910);
or U24911 (N_24911,N_20288,N_20845);
nor U24912 (N_24912,N_19507,N_19866);
and U24913 (N_24913,N_19376,N_18997);
nand U24914 (N_24914,N_19379,N_21010);
and U24915 (N_24915,N_21231,N_21793);
xor U24916 (N_24916,N_19104,N_21422);
and U24917 (N_24917,N_19576,N_20427);
nand U24918 (N_24918,N_19808,N_20070);
or U24919 (N_24919,N_21519,N_20518);
nand U24920 (N_24920,N_19054,N_19016);
and U24921 (N_24921,N_20660,N_20597);
nand U24922 (N_24922,N_18764,N_20108);
and U24923 (N_24923,N_20948,N_21787);
or U24924 (N_24924,N_20578,N_20955);
nor U24925 (N_24925,N_20384,N_21340);
or U24926 (N_24926,N_19195,N_19237);
nand U24927 (N_24927,N_19205,N_19215);
nor U24928 (N_24928,N_20635,N_20681);
nand U24929 (N_24929,N_21483,N_21394);
or U24930 (N_24930,N_20466,N_21390);
and U24931 (N_24931,N_21191,N_19318);
or U24932 (N_24932,N_21867,N_19476);
nand U24933 (N_24933,N_20211,N_19122);
nand U24934 (N_24934,N_19468,N_19724);
nand U24935 (N_24935,N_20463,N_19450);
or U24936 (N_24936,N_21118,N_20356);
nor U24937 (N_24937,N_19162,N_20396);
xnor U24938 (N_24938,N_20916,N_19097);
or U24939 (N_24939,N_19686,N_19891);
nand U24940 (N_24940,N_21603,N_19737);
and U24941 (N_24941,N_21480,N_21643);
nand U24942 (N_24942,N_19071,N_19890);
or U24943 (N_24943,N_20671,N_20419);
nor U24944 (N_24944,N_18798,N_20352);
and U24945 (N_24945,N_21260,N_19346);
xnor U24946 (N_24946,N_19424,N_20211);
and U24947 (N_24947,N_19194,N_21207);
nor U24948 (N_24948,N_19582,N_20893);
or U24949 (N_24949,N_19544,N_20540);
xnor U24950 (N_24950,N_21171,N_19854);
and U24951 (N_24951,N_21769,N_18880);
nor U24952 (N_24952,N_21264,N_19957);
nand U24953 (N_24953,N_19843,N_19694);
and U24954 (N_24954,N_18996,N_20728);
nand U24955 (N_24955,N_21214,N_19293);
nor U24956 (N_24956,N_19666,N_20456);
and U24957 (N_24957,N_19262,N_19788);
xnor U24958 (N_24958,N_19467,N_21440);
and U24959 (N_24959,N_20702,N_19552);
and U24960 (N_24960,N_21321,N_21036);
or U24961 (N_24961,N_19696,N_21284);
and U24962 (N_24962,N_19350,N_20019);
nor U24963 (N_24963,N_19351,N_20405);
nor U24964 (N_24964,N_19460,N_18782);
nor U24965 (N_24965,N_20928,N_20613);
or U24966 (N_24966,N_20261,N_20566);
nand U24967 (N_24967,N_21349,N_20301);
and U24968 (N_24968,N_20963,N_20323);
nor U24969 (N_24969,N_21185,N_20298);
and U24970 (N_24970,N_19474,N_20820);
or U24971 (N_24971,N_20361,N_20979);
or U24972 (N_24972,N_21792,N_19265);
or U24973 (N_24973,N_20405,N_21479);
and U24974 (N_24974,N_21206,N_18767);
nor U24975 (N_24975,N_18786,N_21048);
nor U24976 (N_24976,N_21242,N_20872);
nor U24977 (N_24977,N_20563,N_21568);
or U24978 (N_24978,N_21227,N_20455);
nor U24979 (N_24979,N_21825,N_19201);
or U24980 (N_24980,N_20115,N_19857);
nand U24981 (N_24981,N_19445,N_18960);
xor U24982 (N_24982,N_19395,N_20807);
and U24983 (N_24983,N_20812,N_19659);
nor U24984 (N_24984,N_18819,N_19896);
nand U24985 (N_24985,N_21242,N_21396);
nand U24986 (N_24986,N_20847,N_20420);
or U24987 (N_24987,N_20755,N_19230);
and U24988 (N_24988,N_19520,N_19548);
or U24989 (N_24989,N_21636,N_20657);
nand U24990 (N_24990,N_20482,N_20843);
xnor U24991 (N_24991,N_19899,N_19626);
nand U24992 (N_24992,N_21676,N_19395);
xnor U24993 (N_24993,N_19556,N_19688);
nor U24994 (N_24994,N_21788,N_20141);
xnor U24995 (N_24995,N_20174,N_19509);
nand U24996 (N_24996,N_20119,N_20688);
xor U24997 (N_24997,N_19567,N_20020);
nand U24998 (N_24998,N_20055,N_19354);
xnor U24999 (N_24999,N_18898,N_19720);
nand UO_0 (O_0,N_23898,N_22869);
nand UO_1 (O_1,N_23748,N_24288);
and UO_2 (O_2,N_24869,N_22411);
nand UO_3 (O_3,N_24104,N_22276);
nand UO_4 (O_4,N_24418,N_22206);
and UO_5 (O_5,N_24181,N_21918);
nor UO_6 (O_6,N_24233,N_24195);
or UO_7 (O_7,N_22234,N_23751);
or UO_8 (O_8,N_21876,N_23510);
nor UO_9 (O_9,N_22488,N_22487);
and UO_10 (O_10,N_23798,N_23616);
and UO_11 (O_11,N_22371,N_24782);
and UO_12 (O_12,N_23978,N_22256);
xor UO_13 (O_13,N_23319,N_23962);
nor UO_14 (O_14,N_23244,N_24067);
xor UO_15 (O_15,N_23205,N_24729);
nand UO_16 (O_16,N_23097,N_21941);
nor UO_17 (O_17,N_23493,N_24367);
or UO_18 (O_18,N_23200,N_22294);
nand UO_19 (O_19,N_23960,N_24182);
nor UO_20 (O_20,N_24454,N_22625);
and UO_21 (O_21,N_23331,N_23656);
xor UO_22 (O_22,N_21883,N_24972);
nand UO_23 (O_23,N_23637,N_23008);
xnor UO_24 (O_24,N_23268,N_22194);
nor UO_25 (O_25,N_23341,N_23462);
nor UO_26 (O_26,N_22014,N_23077);
and UO_27 (O_27,N_22860,N_23576);
xor UO_28 (O_28,N_23923,N_22938);
xnor UO_29 (O_29,N_22355,N_24394);
nand UO_30 (O_30,N_24515,N_23223);
nor UO_31 (O_31,N_23850,N_24201);
nand UO_32 (O_32,N_24508,N_24088);
xnor UO_33 (O_33,N_22956,N_22597);
nor UO_34 (O_34,N_24061,N_22244);
nand UO_35 (O_35,N_24493,N_23742);
and UO_36 (O_36,N_24518,N_24828);
and UO_37 (O_37,N_24700,N_23056);
xor UO_38 (O_38,N_23568,N_24805);
or UO_39 (O_39,N_23090,N_24446);
or UO_40 (O_40,N_24795,N_22476);
xnor UO_41 (O_41,N_23142,N_22694);
or UO_42 (O_42,N_22535,N_24392);
and UO_43 (O_43,N_24256,N_23020);
xor UO_44 (O_44,N_22501,N_23424);
nor UO_45 (O_45,N_24040,N_23972);
nand UO_46 (O_46,N_22910,N_22418);
xor UO_47 (O_47,N_23498,N_23677);
xnor UO_48 (O_48,N_23700,N_24161);
xor UO_49 (O_49,N_24970,N_23120);
nor UO_50 (O_50,N_23057,N_24160);
nand UO_51 (O_51,N_23584,N_24534);
or UO_52 (O_52,N_24262,N_23605);
xor UO_53 (O_53,N_24625,N_24445);
nand UO_54 (O_54,N_22266,N_23601);
or UO_55 (O_55,N_23704,N_22830);
and UO_56 (O_56,N_24504,N_22165);
and UO_57 (O_57,N_22275,N_23212);
xnor UO_58 (O_58,N_23563,N_23877);
nor UO_59 (O_59,N_22848,N_23418);
or UO_60 (O_60,N_24412,N_24378);
nor UO_61 (O_61,N_22708,N_22084);
and UO_62 (O_62,N_24707,N_23187);
or UO_63 (O_63,N_23685,N_23956);
and UO_64 (O_64,N_22183,N_24565);
nor UO_65 (O_65,N_22453,N_24967);
nor UO_66 (O_66,N_24029,N_24748);
or UO_67 (O_67,N_24552,N_23232);
or UO_68 (O_68,N_21959,N_23283);
and UO_69 (O_69,N_23351,N_23194);
nand UO_70 (O_70,N_22664,N_22796);
nor UO_71 (O_71,N_24985,N_23976);
nand UO_72 (O_72,N_24092,N_22849);
xnor UO_73 (O_73,N_22451,N_23373);
and UO_74 (O_74,N_23288,N_24557);
xor UO_75 (O_75,N_24395,N_22691);
and UO_76 (O_76,N_23375,N_23808);
and UO_77 (O_77,N_23535,N_22430);
and UO_78 (O_78,N_23835,N_22736);
nand UO_79 (O_79,N_22614,N_22310);
and UO_80 (O_80,N_23069,N_22247);
and UO_81 (O_81,N_23280,N_24963);
and UO_82 (O_82,N_23545,N_24488);
nand UO_83 (O_83,N_24207,N_24882);
nor UO_84 (O_84,N_23233,N_24637);
nor UO_85 (O_85,N_23740,N_22903);
nand UO_86 (O_86,N_23388,N_24750);
nor UO_87 (O_87,N_22224,N_22246);
or UO_88 (O_88,N_23345,N_24720);
nand UO_89 (O_89,N_22981,N_21892);
and UO_90 (O_90,N_22385,N_22945);
or UO_91 (O_91,N_22679,N_24325);
nand UO_92 (O_92,N_23447,N_24487);
nand UO_93 (O_93,N_23186,N_23015);
and UO_94 (O_94,N_24958,N_23692);
nand UO_95 (O_95,N_24562,N_22776);
nand UO_96 (O_96,N_23480,N_22684);
nand UO_97 (O_97,N_23661,N_22346);
xnor UO_98 (O_98,N_23362,N_24172);
nor UO_99 (O_99,N_22146,N_23285);
nor UO_100 (O_100,N_23532,N_23824);
or UO_101 (O_101,N_24678,N_21998);
nand UO_102 (O_102,N_22606,N_23075);
nand UO_103 (O_103,N_22861,N_24796);
and UO_104 (O_104,N_22201,N_22571);
and UO_105 (O_105,N_24472,N_22699);
or UO_106 (O_106,N_22949,N_24352);
nand UO_107 (O_107,N_22635,N_22342);
nor UO_108 (O_108,N_23429,N_23471);
nor UO_109 (O_109,N_24715,N_23529);
and UO_110 (O_110,N_24708,N_24587);
xnor UO_111 (O_111,N_23073,N_22857);
and UO_112 (O_112,N_22370,N_24991);
nor UO_113 (O_113,N_22583,N_22118);
nor UO_114 (O_114,N_22502,N_22397);
or UO_115 (O_115,N_23756,N_23894);
xnor UO_116 (O_116,N_22748,N_23992);
nor UO_117 (O_117,N_22965,N_23941);
and UO_118 (O_118,N_22547,N_22517);
xnor UO_119 (O_119,N_22880,N_24374);
and UO_120 (O_120,N_23414,N_24768);
nand UO_121 (O_121,N_24115,N_24163);
xnor UO_122 (O_122,N_24415,N_22454);
or UO_123 (O_123,N_24086,N_23503);
and UO_124 (O_124,N_24410,N_22859);
nor UO_125 (O_125,N_23182,N_23654);
or UO_126 (O_126,N_24408,N_24316);
xnor UO_127 (O_127,N_22053,N_22213);
and UO_128 (O_128,N_24690,N_22145);
xor UO_129 (O_129,N_22604,N_22494);
nor UO_130 (O_130,N_24491,N_21890);
or UO_131 (O_131,N_24008,N_22549);
or UO_132 (O_132,N_24691,N_23303);
xnor UO_133 (O_133,N_22124,N_23876);
nand UO_134 (O_134,N_23101,N_23128);
nor UO_135 (O_135,N_24610,N_22602);
nor UO_136 (O_136,N_21896,N_22772);
nor UO_137 (O_137,N_23509,N_24854);
nand UO_138 (O_138,N_24373,N_23027);
xor UO_139 (O_139,N_23951,N_23889);
nor UO_140 (O_140,N_24779,N_23118);
xor UO_141 (O_141,N_22022,N_24721);
nand UO_142 (O_142,N_24114,N_22700);
nand UO_143 (O_143,N_24210,N_23557);
nand UO_144 (O_144,N_22661,N_24820);
xnor UO_145 (O_145,N_24949,N_24604);
or UO_146 (O_146,N_23491,N_24226);
and UO_147 (O_147,N_22832,N_24601);
or UO_148 (O_148,N_21939,N_22396);
xnor UO_149 (O_149,N_22435,N_24851);
xor UO_150 (O_150,N_24457,N_23881);
or UO_151 (O_151,N_24248,N_24401);
and UO_152 (O_152,N_24475,N_23279);
xor UO_153 (O_153,N_23433,N_23352);
or UO_154 (O_154,N_22401,N_21935);
or UO_155 (O_155,N_22050,N_21965);
xor UO_156 (O_156,N_21977,N_23010);
xor UO_157 (O_157,N_24862,N_22218);
nand UO_158 (O_158,N_24495,N_24527);
nor UO_159 (O_159,N_22963,N_23486);
and UO_160 (O_160,N_23971,N_22185);
nand UO_161 (O_161,N_23441,N_24289);
or UO_162 (O_162,N_23914,N_24787);
or UO_163 (O_163,N_23423,N_22192);
or UO_164 (O_164,N_23011,N_24931);
and UO_165 (O_165,N_23378,N_24100);
and UO_166 (O_166,N_21968,N_24155);
and UO_167 (O_167,N_24359,N_24965);
and UO_168 (O_168,N_23045,N_23838);
nand UO_169 (O_169,N_23003,N_24536);
nor UO_170 (O_170,N_24784,N_24372);
and UO_171 (O_171,N_23794,N_22734);
or UO_172 (O_172,N_24636,N_22354);
xor UO_173 (O_173,N_24083,N_22461);
and UO_174 (O_174,N_22788,N_24821);
and UO_175 (O_175,N_22566,N_24522);
xor UO_176 (O_176,N_22127,N_21966);
and UO_177 (O_177,N_23959,N_22233);
nor UO_178 (O_178,N_22463,N_24688);
xor UO_179 (O_179,N_23591,N_22674);
nor UO_180 (O_180,N_22248,N_24878);
and UO_181 (O_181,N_23365,N_24102);
xor UO_182 (O_182,N_23500,N_24190);
or UO_183 (O_183,N_22554,N_22864);
nand UO_184 (O_184,N_22912,N_22775);
or UO_185 (O_185,N_23322,N_22977);
xnor UO_186 (O_186,N_24049,N_22836);
nand UO_187 (O_187,N_22626,N_22415);
or UO_188 (O_188,N_24089,N_23620);
nand UO_189 (O_189,N_24986,N_24643);
xor UO_190 (O_190,N_24036,N_23579);
nor UO_191 (O_191,N_22685,N_24987);
and UO_192 (O_192,N_23708,N_22120);
nor UO_193 (O_193,N_24667,N_23961);
nor UO_194 (O_194,N_24911,N_22272);
xor UO_195 (O_195,N_22364,N_23145);
xnor UO_196 (O_196,N_23136,N_24634);
nor UO_197 (O_197,N_23347,N_23445);
or UO_198 (O_198,N_24344,N_23631);
nor UO_199 (O_199,N_24922,N_22991);
xor UO_200 (O_200,N_24143,N_24663);
or UO_201 (O_201,N_22989,N_23397);
and UO_202 (O_202,N_21906,N_22045);
nor UO_203 (O_203,N_24662,N_22667);
or UO_204 (O_204,N_21911,N_22512);
nand UO_205 (O_205,N_23410,N_23088);
xnor UO_206 (O_206,N_23391,N_23337);
or UO_207 (O_207,N_22779,N_22777);
nand UO_208 (O_208,N_24261,N_24221);
nor UO_209 (O_209,N_22652,N_23848);
and UO_210 (O_210,N_21917,N_21954);
xnor UO_211 (O_211,N_22967,N_22374);
nor UO_212 (O_212,N_23925,N_22305);
nand UO_213 (O_213,N_24656,N_24430);
or UO_214 (O_214,N_22373,N_23272);
nand UO_215 (O_215,N_24753,N_22469);
nand UO_216 (O_216,N_23757,N_23866);
and UO_217 (O_217,N_21886,N_24122);
nor UO_218 (O_218,N_24918,N_24975);
xor UO_219 (O_219,N_24760,N_23609);
and UO_220 (O_220,N_23763,N_23475);
xor UO_221 (O_221,N_22363,N_23313);
or UO_222 (O_222,N_22892,N_23589);
or UO_223 (O_223,N_21936,N_23257);
or UO_224 (O_224,N_22390,N_24479);
nand UO_225 (O_225,N_23667,N_22601);
nor UO_226 (O_226,N_23921,N_24990);
nor UO_227 (O_227,N_24481,N_23977);
or UO_228 (O_228,N_23370,N_23549);
xnor UO_229 (O_229,N_22319,N_22280);
or UO_230 (O_230,N_22432,N_23728);
xnor UO_231 (O_231,N_23823,N_22387);
xnor UO_232 (O_232,N_24630,N_23098);
nand UO_233 (O_233,N_23733,N_24942);
or UO_234 (O_234,N_23376,N_24244);
xnor UO_235 (O_235,N_23566,N_22878);
or UO_236 (O_236,N_23443,N_23421);
or UO_237 (O_237,N_22842,N_24057);
and UO_238 (O_238,N_24137,N_23300);
xor UO_239 (O_239,N_21880,N_24499);
nor UO_240 (O_240,N_24300,N_22722);
xnor UO_241 (O_241,N_23317,N_24129);
xnor UO_242 (O_242,N_23301,N_23980);
nor UO_243 (O_243,N_22621,N_23691);
xnor UO_244 (O_244,N_22671,N_22564);
and UO_245 (O_245,N_21947,N_24901);
xor UO_246 (O_246,N_23093,N_24365);
xnor UO_247 (O_247,N_24361,N_24406);
or UO_248 (O_248,N_24448,N_23765);
xnor UO_249 (O_249,N_24568,N_24648);
nand UO_250 (O_250,N_23269,N_23729);
or UO_251 (O_251,N_24076,N_24347);
and UO_252 (O_252,N_24533,N_24863);
or UO_253 (O_253,N_24659,N_24896);
and UO_254 (O_254,N_24154,N_24212);
nand UO_255 (O_255,N_24250,N_23104);
xnor UO_256 (O_256,N_24801,N_22153);
nand UO_257 (O_257,N_23109,N_23786);
nor UO_258 (O_258,N_22990,N_22330);
xnor UO_259 (O_259,N_22181,N_22062);
or UO_260 (O_260,N_23001,N_22619);
and UO_261 (O_261,N_24291,N_24732);
xnor UO_262 (O_262,N_22026,N_24323);
xor UO_263 (O_263,N_22605,N_23036);
and UO_264 (O_264,N_23795,N_22980);
xnor UO_265 (O_265,N_22716,N_22530);
or UO_266 (O_266,N_24124,N_24617);
and UO_267 (O_267,N_22085,N_22816);
nand UO_268 (O_268,N_23577,N_23260);
nand UO_269 (O_269,N_24413,N_22377);
xnor UO_270 (O_270,N_23744,N_23891);
or UO_271 (O_271,N_23581,N_22267);
and UO_272 (O_272,N_23061,N_24741);
nand UO_273 (O_273,N_24169,N_22543);
or UO_274 (O_274,N_22702,N_22651);
and UO_275 (O_275,N_23647,N_23964);
xor UO_276 (O_276,N_23701,N_23641);
nor UO_277 (O_277,N_23864,N_23476);
nand UO_278 (O_278,N_21981,N_23507);
or UO_279 (O_279,N_23776,N_21976);
and UO_280 (O_280,N_22523,N_22303);
xnor UO_281 (O_281,N_23295,N_23861);
xnor UO_282 (O_282,N_24280,N_23344);
nor UO_283 (O_283,N_21999,N_24010);
nor UO_284 (O_284,N_24242,N_24332);
nand UO_285 (O_285,N_23315,N_24554);
xor UO_286 (O_286,N_23927,N_24510);
and UO_287 (O_287,N_23267,N_24001);
xnor UO_288 (O_288,N_21932,N_23856);
or UO_289 (O_289,N_23506,N_23687);
nor UO_290 (O_290,N_24393,N_22909);
nand UO_291 (O_291,N_24600,N_22255);
or UO_292 (O_292,N_22637,N_23931);
nand UO_293 (O_293,N_24765,N_23095);
and UO_294 (O_294,N_23693,N_24489);
xnor UO_295 (O_295,N_24693,N_23564);
nor UO_296 (O_296,N_24145,N_24632);
xnor UO_297 (O_297,N_24260,N_24506);
xor UO_298 (O_298,N_23502,N_22157);
xor UO_299 (O_299,N_24728,N_21912);
nor UO_300 (O_300,N_24094,N_24476);
and UO_301 (O_301,N_22129,N_22365);
and UO_302 (O_302,N_21894,N_24171);
xnor UO_303 (O_303,N_24016,N_23556);
nand UO_304 (O_304,N_24063,N_24671);
nand UO_305 (O_305,N_22791,N_23668);
nand UO_306 (O_306,N_24236,N_22813);
nor UO_307 (O_307,N_23780,N_23916);
nand UO_308 (O_308,N_24304,N_24885);
or UO_309 (O_309,N_23890,N_22103);
xnor UO_310 (O_310,N_22822,N_24184);
nand UO_311 (O_311,N_22636,N_23711);
and UO_312 (O_312,N_22988,N_24898);
or UO_313 (O_313,N_23671,N_22843);
nand UO_314 (O_314,N_24699,N_24019);
nor UO_315 (O_315,N_22942,N_23530);
nor UO_316 (O_316,N_24711,N_24031);
nand UO_317 (O_317,N_24494,N_22018);
xor UO_318 (O_318,N_22091,N_22260);
and UO_319 (O_319,N_22992,N_23067);
nor UO_320 (O_320,N_24563,N_24640);
or UO_321 (O_321,N_23330,N_22525);
nor UO_322 (O_322,N_24904,N_22874);
nand UO_323 (O_323,N_23967,N_23394);
and UO_324 (O_324,N_22057,N_24468);
nor UO_325 (O_325,N_23353,N_23108);
nor UO_326 (O_326,N_23760,N_23826);
nor UO_327 (O_327,N_22477,N_23430);
nand UO_328 (O_328,N_24984,N_23039);
and UO_329 (O_329,N_22666,N_23802);
nor UO_330 (O_330,N_24649,N_22863);
xor UO_331 (O_331,N_22111,N_24995);
and UO_332 (O_332,N_24302,N_22445);
nand UO_333 (O_333,N_24402,N_23783);
and UO_334 (O_334,N_22516,N_23173);
and UO_335 (O_335,N_24611,N_22895);
and UO_336 (O_336,N_24564,N_23516);
xnor UO_337 (O_337,N_22316,N_22376);
nand UO_338 (O_338,N_22426,N_22862);
nor UO_339 (O_339,N_23932,N_22866);
xnor UO_340 (O_340,N_23350,N_24389);
or UO_341 (O_341,N_23562,N_22296);
and UO_342 (O_342,N_22208,N_22329);
or UO_343 (O_343,N_23255,N_24382);
xor UO_344 (O_344,N_22040,N_24126);
or UO_345 (O_345,N_22473,N_22920);
or UO_346 (O_346,N_21994,N_24186);
or UO_347 (O_347,N_23640,N_22238);
xor UO_348 (O_348,N_23974,N_24022);
xnor UO_349 (O_349,N_22160,N_22505);
nor UO_350 (O_350,N_22351,N_23761);
xor UO_351 (O_351,N_24309,N_23539);
xnor UO_352 (O_352,N_21914,N_24103);
nor UO_353 (O_353,N_24698,N_22675);
and UO_354 (O_354,N_22203,N_24993);
nor UO_355 (O_355,N_24629,N_24553);
nor UO_356 (O_356,N_23467,N_23803);
nand UO_357 (O_357,N_23274,N_23906);
and UO_358 (O_358,N_22555,N_24689);
nor UO_359 (O_359,N_23335,N_23032);
nor UO_360 (O_360,N_22077,N_24523);
nand UO_361 (O_361,N_24004,N_22918);
xor UO_362 (O_362,N_23814,N_22792);
or UO_363 (O_363,N_24381,N_24832);
nor UO_364 (O_364,N_24093,N_24085);
and UO_365 (O_365,N_23204,N_22444);
xnor UO_366 (O_366,N_22802,N_24358);
or UO_367 (O_367,N_24482,N_23796);
or UO_368 (O_368,N_24191,N_22324);
nand UO_369 (O_369,N_23401,N_24015);
xor UO_370 (O_370,N_22639,N_23174);
xor UO_371 (O_371,N_23117,N_24179);
nand UO_372 (O_372,N_24722,N_24830);
and UO_373 (O_373,N_24881,N_23134);
and UO_374 (O_374,N_23707,N_23800);
xnor UO_375 (O_375,N_22035,N_22897);
nor UO_376 (O_376,N_22350,N_24345);
or UO_377 (O_377,N_24183,N_23540);
xor UO_378 (O_378,N_22184,N_24439);
and UO_379 (O_379,N_23007,N_21927);
nand UO_380 (O_380,N_24007,N_24437);
or UO_381 (O_381,N_22594,N_24380);
xnor UO_382 (O_382,N_22392,N_24694);
or UO_383 (O_383,N_24474,N_23215);
and UO_384 (O_384,N_22713,N_24567);
or UO_385 (O_385,N_24060,N_22873);
xor UO_386 (O_386,N_24798,N_24148);
and UO_387 (O_387,N_22766,N_22553);
nand UO_388 (O_388,N_23725,N_24059);
xnor UO_389 (O_389,N_22220,N_24342);
and UO_390 (O_390,N_22312,N_22946);
xnor UO_391 (O_391,N_24839,N_23788);
and UO_392 (O_392,N_22440,N_24905);
and UO_393 (O_393,N_21963,N_23377);
nor UO_394 (O_394,N_22030,N_24872);
nor UO_395 (O_395,N_23291,N_22693);
xor UO_396 (O_396,N_24274,N_21877);
xor UO_397 (O_397,N_22656,N_24000);
nor UO_398 (O_398,N_23218,N_24511);
and UO_399 (O_399,N_22982,N_24946);
or UO_400 (O_400,N_23793,N_24298);
and UO_401 (O_401,N_24793,N_23307);
xor UO_402 (O_402,N_24051,N_24313);
nand UO_403 (O_403,N_23195,N_24895);
or UO_404 (O_404,N_24902,N_23630);
nor UO_405 (O_405,N_24193,N_23806);
nand UO_406 (O_406,N_23087,N_24147);
xor UO_407 (O_407,N_24384,N_24025);
nand UO_408 (O_408,N_24594,N_23271);
xor UO_409 (O_409,N_23743,N_23459);
xnor UO_410 (O_410,N_22643,N_24285);
nand UO_411 (O_411,N_22737,N_23565);
or UO_412 (O_412,N_23821,N_23356);
and UO_413 (O_413,N_22121,N_22761);
nand UO_414 (O_414,N_23137,N_22966);
and UO_415 (O_415,N_22534,N_22793);
xnor UO_416 (O_416,N_24469,N_22572);
and UO_417 (O_417,N_23935,N_23593);
xor UO_418 (O_418,N_24937,N_22600);
or UO_419 (O_419,N_23102,N_23273);
or UO_420 (O_420,N_24919,N_23917);
or UO_421 (O_421,N_23696,N_22041);
nand UO_422 (O_422,N_22474,N_22723);
or UO_423 (O_423,N_24253,N_24329);
nor UO_424 (O_424,N_24661,N_24716);
or UO_425 (O_425,N_22872,N_22347);
nand UO_426 (O_426,N_22493,N_22361);
or UO_427 (O_427,N_23942,N_23703);
nand UO_428 (O_428,N_23496,N_22607);
xor UO_429 (O_429,N_23302,N_22406);
nor UO_430 (O_430,N_23304,N_23842);
nor UO_431 (O_431,N_22313,N_24013);
nand UO_432 (O_432,N_24296,N_24731);
or UO_433 (O_433,N_24270,N_23883);
or UO_434 (O_434,N_24203,N_24556);
xor UO_435 (O_435,N_23643,N_24002);
xnor UO_436 (O_436,N_22514,N_22235);
nand UO_437 (O_437,N_24319,N_23250);
or UO_438 (O_438,N_24945,N_21925);
nor UO_439 (O_439,N_22188,N_23550);
nor UO_440 (O_440,N_22226,N_23025);
nor UO_441 (O_441,N_24194,N_22712);
xnor UO_442 (O_442,N_24915,N_22409);
nor UO_443 (O_443,N_24762,N_24903);
or UO_444 (O_444,N_22638,N_24615);
nand UO_445 (O_445,N_22941,N_22940);
nor UO_446 (O_446,N_22780,N_22907);
or UO_447 (O_447,N_22817,N_23127);
nand UO_448 (O_448,N_23888,N_24467);
or UO_449 (O_449,N_23085,N_22252);
or UO_450 (O_450,N_24224,N_24635);
or UO_451 (O_451,N_22086,N_23446);
or UO_452 (O_452,N_23574,N_22076);
xnor UO_453 (O_453,N_22567,N_24346);
and UO_454 (O_454,N_22038,N_23277);
xnor UO_455 (O_455,N_22054,N_24547);
nor UO_456 (O_456,N_23874,N_23034);
xor UO_457 (O_457,N_22595,N_23044);
nor UO_458 (O_458,N_22341,N_24790);
nand UO_459 (O_459,N_22386,N_23764);
nand UO_460 (O_460,N_22056,N_23284);
and UO_461 (O_461,N_24497,N_24657);
nor UO_462 (O_462,N_24774,N_23266);
nor UO_463 (O_463,N_24357,N_23311);
and UO_464 (O_464,N_24355,N_23227);
and UO_465 (O_465,N_24619,N_21946);
nor UO_466 (O_466,N_23412,N_22999);
xnor UO_467 (O_467,N_24940,N_24733);
or UO_468 (O_468,N_22790,N_22998);
nand UO_469 (O_469,N_22921,N_24807);
nor UO_470 (O_470,N_22378,N_22389);
and UO_471 (O_471,N_24107,N_24151);
or UO_472 (O_472,N_24792,N_23159);
or UO_473 (O_473,N_24664,N_22152);
and UO_474 (O_474,N_22798,N_21920);
xnor UO_475 (O_475,N_23913,N_24106);
nor UO_476 (O_476,N_24530,N_23275);
and UO_477 (O_477,N_23122,N_22835);
xor UO_478 (O_478,N_24388,N_22692);
or UO_479 (O_479,N_22925,N_22245);
and UO_480 (O_480,N_24621,N_23658);
or UO_481 (O_481,N_23755,N_22804);
or UO_482 (O_482,N_24818,N_24071);
and UO_483 (O_483,N_22338,N_22789);
nor UO_484 (O_484,N_22007,N_23047);
xor UO_485 (O_485,N_21888,N_23702);
xnor UO_486 (O_486,N_23072,N_23078);
nand UO_487 (O_487,N_22683,N_23018);
xor UO_488 (O_488,N_22357,N_23997);
nand UO_489 (O_489,N_24641,N_24473);
or UO_490 (O_490,N_24880,N_24177);
and UO_491 (O_491,N_24532,N_24813);
and UO_492 (O_492,N_23332,N_24577);
or UO_493 (O_493,N_24046,N_22610);
nand UO_494 (O_494,N_24939,N_24237);
xor UO_495 (O_495,N_23939,N_24150);
nor UO_496 (O_496,N_22968,N_23621);
and UO_497 (O_497,N_23399,N_24650);
and UO_498 (O_498,N_22771,N_24804);
or UO_499 (O_499,N_24360,N_23343);
nor UO_500 (O_500,N_22508,N_22042);
and UO_501 (O_501,N_23222,N_21937);
and UO_502 (O_502,N_23296,N_21938);
xnor UO_503 (O_503,N_24566,N_24794);
or UO_504 (O_504,N_24623,N_22905);
xor UO_505 (O_505,N_24238,N_22647);
nand UO_506 (O_506,N_23096,N_23183);
or UO_507 (O_507,N_22230,N_22522);
nor UO_508 (O_508,N_23023,N_22154);
or UO_509 (O_509,N_23214,N_21929);
and UO_510 (O_510,N_22617,N_24585);
or UO_511 (O_511,N_23651,N_23680);
nand UO_512 (O_512,N_22178,N_24118);
nand UO_513 (O_513,N_24337,N_23569);
nor UO_514 (O_514,N_23149,N_24845);
xnor UO_515 (O_515,N_23022,N_23256);
xor UO_516 (O_516,N_23940,N_22900);
and UO_517 (O_517,N_24770,N_23827);
and UO_518 (O_518,N_22891,N_24426);
and UO_519 (O_519,N_23054,N_24101);
nor UO_520 (O_520,N_23650,N_24197);
nand UO_521 (O_521,N_21931,N_24537);
or UO_522 (O_522,N_22886,N_22101);
or UO_523 (O_523,N_22241,N_21875);
nand UO_524 (O_524,N_22955,N_22958);
and UO_525 (O_525,N_24159,N_23804);
and UO_526 (O_526,N_23138,N_21986);
nand UO_527 (O_527,N_24616,N_23986);
and UO_528 (O_528,N_23179,N_24219);
or UO_529 (O_529,N_22109,N_23140);
nor UO_530 (O_530,N_22531,N_22393);
xor UO_531 (O_531,N_24058,N_22011);
or UO_532 (O_532,N_22932,N_24591);
xor UO_533 (O_533,N_22130,N_23937);
or UO_534 (O_534,N_24875,N_22196);
xnor UO_535 (O_535,N_22254,N_22677);
nand UO_536 (O_536,N_23930,N_22824);
or UO_537 (O_537,N_22933,N_24470);
nor UO_538 (O_538,N_23281,N_23282);
xnor UO_539 (O_539,N_24879,N_23481);
or UO_540 (O_540,N_21960,N_23732);
or UO_541 (O_541,N_24123,N_24047);
nand UO_542 (O_542,N_24944,N_23403);
nor UO_543 (O_543,N_24864,N_22491);
nand UO_544 (O_544,N_22616,N_22036);
nor UO_545 (O_545,N_24157,N_23933);
nand UO_546 (O_546,N_24156,N_22507);
and UO_547 (O_547,N_24174,N_22485);
and UO_548 (O_548,N_23684,N_24502);
or UO_549 (O_549,N_24806,N_24275);
xnor UO_550 (O_550,N_23000,N_24865);
or UO_551 (O_551,N_23346,N_22953);
xnor UO_552 (O_552,N_24239,N_22964);
xor UO_553 (O_553,N_24167,N_22399);
nand UO_554 (O_554,N_22648,N_24379);
nand UO_555 (O_555,N_22452,N_23892);
or UO_556 (O_556,N_21923,N_23298);
or UO_557 (O_557,N_23797,N_24268);
nor UO_558 (O_558,N_21974,N_23172);
nand UO_559 (O_559,N_21972,N_23184);
xor UO_560 (O_560,N_24639,N_24670);
or UO_561 (O_561,N_24421,N_23606);
and UO_562 (O_562,N_23175,N_23193);
nand UO_563 (O_563,N_23457,N_24303);
xor UO_564 (O_564,N_24097,N_23849);
xnor UO_565 (O_565,N_23396,N_23489);
and UO_566 (O_566,N_22177,N_24999);
xor UO_567 (O_567,N_23664,N_22285);
nand UO_568 (O_568,N_23766,N_24950);
and UO_569 (O_569,N_23106,N_23949);
xor UO_570 (O_570,N_24041,N_23522);
nand UO_571 (O_571,N_24981,N_23536);
nand UO_572 (O_572,N_24840,N_21907);
xnor UO_573 (O_573,N_23816,N_21881);
xnor UO_574 (O_574,N_23151,N_24362);
xnor UO_575 (O_575,N_23306,N_22384);
xnor UO_576 (O_576,N_22805,N_24442);
xnor UO_577 (O_577,N_23813,N_23099);
xor UO_578 (O_578,N_23759,N_23709);
or UO_579 (O_579,N_23334,N_22459);
nor UO_580 (O_580,N_23596,N_22483);
xor UO_581 (O_581,N_22883,N_24673);
nor UO_582 (O_582,N_24458,N_24178);
or UO_583 (O_583,N_24139,N_24297);
nor UO_584 (O_584,N_24841,N_24718);
or UO_585 (O_585,N_24746,N_22634);
nor UO_586 (O_586,N_22009,N_24168);
nand UO_587 (O_587,N_23546,N_24520);
or UO_588 (O_588,N_24633,N_22801);
or UO_589 (O_589,N_24225,N_23604);
and UO_590 (O_590,N_24876,N_23004);
and UO_591 (O_591,N_22425,N_24397);
or UO_592 (O_592,N_23103,N_23320);
nand UO_593 (O_593,N_23610,N_22663);
xor UO_594 (O_594,N_23390,N_23846);
and UO_595 (O_595,N_22288,N_22043);
nor UO_596 (O_596,N_22122,N_23613);
xnor UO_597 (O_597,N_22322,N_24273);
and UO_598 (O_598,N_24091,N_21953);
and UO_599 (O_599,N_22975,N_24254);
and UO_600 (O_600,N_23675,N_24466);
or UO_601 (O_601,N_23870,N_23248);
nand UO_602 (O_602,N_24812,N_23470);
nand UO_603 (O_603,N_23996,N_23199);
xor UO_604 (O_604,N_22436,N_22937);
or UO_605 (O_605,N_23177,N_24582);
and UO_606 (O_606,N_23695,N_23855);
and UO_607 (O_607,N_24434,N_24899);
nor UO_608 (O_608,N_24651,N_22751);
and UO_609 (O_609,N_24558,N_23790);
nand UO_610 (O_610,N_24294,N_24377);
and UO_611 (O_611,N_23024,N_22733);
and UO_612 (O_612,N_24292,N_23338);
and UO_613 (O_613,N_21926,N_24205);
or UO_614 (O_614,N_24953,N_22471);
or UO_615 (O_615,N_22765,N_23957);
nor UO_616 (O_616,N_22405,N_23287);
nor UO_617 (O_617,N_23029,N_23561);
xnor UO_618 (O_618,N_23171,N_22741);
nor UO_619 (O_619,N_23926,N_23316);
nand UO_620 (O_620,N_24529,N_24279);
nand UO_621 (O_621,N_23595,N_23904);
and UO_622 (O_622,N_22269,N_23030);
nor UO_623 (O_623,N_24082,N_22499);
xnor UO_624 (O_624,N_22447,N_23782);
nor UO_625 (O_625,N_24333,N_24121);
nor UO_626 (O_626,N_24961,N_24120);
nand UO_627 (O_627,N_22837,N_24816);
nor UO_628 (O_628,N_24460,N_22497);
or UO_629 (O_629,N_22333,N_23290);
nand UO_630 (O_630,N_22974,N_24290);
xnor UO_631 (O_631,N_24858,N_22498);
or UO_632 (O_632,N_24714,N_24701);
xor UO_633 (O_633,N_23455,N_23224);
nand UO_634 (O_634,N_24544,N_23002);
or UO_635 (O_635,N_22264,N_22850);
or UO_636 (O_636,N_23435,N_24980);
xor UO_637 (O_637,N_24593,N_23474);
and UO_638 (O_638,N_22623,N_23213);
nor UO_639 (O_639,N_24276,N_22081);
nor UO_640 (O_640,N_24692,N_24978);
and UO_641 (O_641,N_24827,N_23652);
nand UO_642 (O_642,N_24817,N_22984);
xor UO_643 (O_643,N_24767,N_23525);
nor UO_644 (O_644,N_24012,N_22318);
and UO_645 (O_645,N_22413,N_22190);
xor UO_646 (O_646,N_22740,N_22456);
nand UO_647 (O_647,N_21885,N_22890);
nand UO_648 (O_648,N_23936,N_24606);
and UO_649 (O_649,N_24668,N_23526);
or UO_650 (O_650,N_22422,N_23543);
xor UO_651 (O_651,N_23386,N_21933);
nor UO_652 (O_652,N_24924,N_24066);
and UO_653 (O_653,N_24386,N_24561);
and UO_654 (O_654,N_22151,N_23750);
nand UO_655 (O_655,N_24087,N_24889);
nand UO_656 (O_656,N_21922,N_24459);
or UO_657 (O_657,N_24095,N_22879);
nor UO_658 (O_658,N_23712,N_22759);
nand UO_659 (O_659,N_23857,N_24829);
xnor UO_660 (O_660,N_23792,N_22845);
xor UO_661 (O_661,N_24907,N_23739);
xnor UO_662 (O_662,N_23258,N_24614);
or UO_663 (O_663,N_23357,N_22884);
xnor UO_664 (O_664,N_24815,N_24775);
or UO_665 (O_665,N_24541,N_24706);
xor UO_666 (O_666,N_24810,N_22174);
and UO_667 (O_667,N_23820,N_24441);
or UO_668 (O_668,N_22214,N_23990);
xor UO_669 (O_669,N_22381,N_23625);
nand UO_670 (O_670,N_24065,N_22348);
and UO_671 (O_671,N_24144,N_24175);
and UO_672 (O_672,N_22345,N_22079);
or UO_673 (O_673,N_22724,N_24166);
nand UO_674 (O_674,N_23392,N_24234);
xnor UO_675 (O_675,N_23147,N_23843);
xor UO_676 (O_676,N_22019,N_24020);
or UO_677 (O_677,N_22315,N_23487);
nor UO_678 (O_678,N_24119,N_23713);
xnor UO_679 (O_679,N_24890,N_24436);
nor UO_680 (O_680,N_22125,N_22380);
nand UO_681 (O_681,N_22526,N_22797);
nor UO_682 (O_682,N_24836,N_23062);
or UO_683 (O_683,N_23859,N_23166);
nand UO_684 (O_684,N_24245,N_23155);
nand UO_685 (O_685,N_24938,N_22356);
nand UO_686 (O_686,N_23135,N_24165);
nand UO_687 (O_687,N_22211,N_22673);
nand UO_688 (O_688,N_22149,N_24605);
or UO_689 (O_689,N_22136,N_24724);
and UO_690 (O_690,N_23360,N_22829);
xnor UO_691 (O_691,N_24416,N_22618);
and UO_692 (O_692,N_23772,N_23710);
xnor UO_693 (O_693,N_24744,N_24884);
or UO_694 (O_694,N_24009,N_22750);
and UO_695 (O_695,N_22686,N_24422);
xnor UO_696 (O_696,N_22987,N_22270);
and UO_697 (O_697,N_24512,N_22304);
or UO_698 (O_698,N_22585,N_24464);
xor UO_699 (O_699,N_23611,N_22037);
nand UO_700 (O_700,N_21934,N_22015);
nor UO_701 (O_701,N_24222,N_24951);
and UO_702 (O_702,N_22769,N_22856);
and UO_703 (O_703,N_23089,N_22362);
nor UO_704 (O_704,N_23981,N_22369);
or UO_705 (O_705,N_23374,N_23063);
and UO_706 (O_706,N_23091,N_23382);
nand UO_707 (O_707,N_24048,N_22279);
or UO_708 (O_708,N_22899,N_24590);
nand UO_709 (O_709,N_24079,N_23832);
xnor UO_710 (O_710,N_22858,N_22368);
and UO_711 (O_711,N_23727,N_24540);
nor UO_712 (O_712,N_23310,N_23779);
nor UO_713 (O_713,N_22913,N_22375);
or UO_714 (O_714,N_22917,N_22743);
or UO_715 (O_715,N_22462,N_23985);
nor UO_716 (O_716,N_23599,N_22576);
or UO_717 (O_717,N_21930,N_23124);
and UO_718 (O_718,N_23229,N_22970);
nor UO_719 (O_719,N_24324,N_22847);
and UO_720 (O_720,N_24069,N_24339);
nand UO_721 (O_721,N_23998,N_22110);
nand UO_722 (O_722,N_24505,N_22755);
xnor UO_723 (O_723,N_23681,N_24973);
nand UO_724 (O_724,N_22358,N_24391);
and UO_725 (O_725,N_21900,N_22821);
or UO_726 (O_726,N_24368,N_23948);
or UO_727 (O_727,N_24035,N_23895);
and UO_728 (O_728,N_23129,N_23867);
nand UO_729 (O_729,N_23406,N_22412);
and UO_730 (O_730,N_23081,N_22005);
nor UO_731 (O_731,N_24149,N_24135);
xnor UO_732 (O_732,N_22359,N_24450);
nor UO_733 (O_733,N_23381,N_23226);
or UO_734 (O_734,N_23686,N_22317);
nand UO_735 (O_735,N_24727,N_23551);
and UO_736 (O_736,N_23982,N_22825);
nor UO_737 (O_737,N_22550,N_23648);
nor UO_738 (O_738,N_22710,N_22670);
and UO_739 (O_739,N_22481,N_23600);
xor UO_740 (O_740,N_23523,N_22870);
and UO_741 (O_741,N_24132,N_24618);
and UO_742 (O_742,N_22711,N_23329);
or UO_743 (O_743,N_24586,N_22746);
nand UO_744 (O_744,N_23006,N_22479);
or UO_745 (O_745,N_24808,N_22803);
or UO_746 (O_746,N_24030,N_24516);
nor UO_747 (O_747,N_22237,N_22672);
xnor UO_748 (O_748,N_24954,N_23349);
xnor UO_749 (O_749,N_22575,N_21997);
nand UO_750 (O_750,N_22764,N_21969);
and UO_751 (O_751,N_24626,N_23170);
and UO_752 (O_752,N_22059,N_22820);
and UO_753 (O_753,N_23230,N_23771);
nor UO_754 (O_754,N_22428,N_24255);
and UO_755 (O_755,N_23466,N_22721);
or UO_756 (O_756,N_24928,N_22003);
nor UO_757 (O_757,N_24734,N_22680);
nor UO_758 (O_758,N_23513,N_22349);
xnor UO_759 (O_759,N_23178,N_23624);
or UO_760 (O_760,N_23465,N_22628);
and UO_761 (O_761,N_23520,N_24490);
nand UO_762 (O_762,N_22394,N_22046);
or UO_763 (O_763,N_22423,N_22326);
xnor UO_764 (O_764,N_24571,N_23646);
and UO_765 (O_765,N_22158,N_24870);
nand UO_766 (O_766,N_23934,N_23863);
xnor UO_767 (O_767,N_24595,N_24726);
xor UO_768 (O_768,N_22001,N_23785);
or UO_769 (O_769,N_22565,N_23408);
xnor UO_770 (O_770,N_22714,N_23425);
nor UO_771 (O_771,N_22705,N_24501);
xnor UO_772 (O_772,N_22144,N_22563);
nand UO_773 (O_773,N_21909,N_23206);
nor UO_774 (O_774,N_23146,N_23560);
nor UO_775 (O_775,N_23618,N_23494);
nand UO_776 (O_776,N_24241,N_22117);
or UO_777 (O_777,N_24471,N_23947);
nor UO_778 (O_778,N_24216,N_22106);
nand UO_779 (O_779,N_24866,N_22687);
or UO_780 (O_780,N_24886,N_24916);
nor UO_781 (O_781,N_24350,N_23905);
xor UO_782 (O_782,N_22800,N_23235);
nor UO_783 (O_783,N_23021,N_22016);
nand UO_784 (O_784,N_24349,N_22753);
nor UO_785 (O_785,N_23767,N_23236);
or UO_786 (O_786,N_24583,N_22784);
nand UO_787 (O_787,N_23969,N_23716);
xnor UO_788 (O_788,N_24281,N_24011);
nor UO_789 (O_789,N_22414,N_23309);
xor UO_790 (O_790,N_24315,N_23458);
nand UO_791 (O_791,N_23395,N_24038);
nor UO_792 (O_792,N_22088,N_22819);
and UO_793 (O_793,N_22928,N_24705);
nor UO_794 (O_794,N_24215,N_22882);
and UO_795 (O_795,N_22155,N_23839);
nand UO_796 (O_796,N_24252,N_21990);
nor UO_797 (O_797,N_24743,N_24628);
or UO_798 (O_798,N_22758,N_22996);
xnor UO_799 (O_799,N_24982,N_23860);
nand UO_800 (O_800,N_24723,N_22551);
nand UO_801 (O_801,N_23815,N_22002);
nand UO_802 (O_802,N_23544,N_24405);
and UO_803 (O_803,N_23689,N_24042);
nor UO_804 (O_804,N_23537,N_21901);
nand UO_805 (O_805,N_22199,N_22927);
nand UO_806 (O_806,N_23679,N_22725);
nand UO_807 (O_807,N_22496,N_24039);
xnor UO_808 (O_808,N_23263,N_23035);
and UO_809 (O_809,N_22660,N_24189);
and UO_810 (O_810,N_24853,N_24644);
nand UO_811 (O_811,N_22204,N_22500);
and UO_812 (O_812,N_24213,N_23369);
nand UO_813 (O_813,N_23717,N_23952);
nand UO_814 (O_814,N_23538,N_23490);
xor UO_815 (O_815,N_24783,N_24580);
and UO_816 (O_816,N_24328,N_22727);
and UO_817 (O_817,N_22277,N_22286);
xor UO_818 (O_818,N_23852,N_23644);
and UO_819 (O_819,N_23524,N_22028);
nand UO_820 (O_820,N_24761,N_24525);
nor UO_821 (O_821,N_24575,N_22559);
nor UO_822 (O_822,N_24077,N_22325);
or UO_823 (O_823,N_22838,N_22099);
xor UO_824 (O_824,N_23383,N_24271);
nor UO_825 (O_825,N_23634,N_22176);
nand UO_826 (O_826,N_22058,N_22592);
or UO_827 (O_827,N_22115,N_23293);
or UO_828 (O_828,N_23385,N_22630);
nor UO_829 (O_829,N_22402,N_22229);
nor UO_830 (O_830,N_22867,N_24396);
xor UO_831 (O_831,N_22962,N_22069);
and UO_832 (O_832,N_23775,N_23627);
or UO_833 (O_833,N_24598,N_23946);
nand UO_834 (O_834,N_24871,N_23042);
and UO_835 (O_835,N_24293,N_23837);
xnor UO_836 (O_836,N_22078,N_24134);
or UO_837 (O_837,N_23731,N_23809);
xnor UO_838 (O_838,N_23305,N_24539);
and UO_839 (O_839,N_22391,N_24068);
nand UO_840 (O_840,N_22061,N_23119);
nor UO_841 (O_841,N_22560,N_22398);
or UO_842 (O_842,N_23754,N_24752);
nor UO_843 (O_843,N_22760,N_22768);
nand UO_844 (O_844,N_23811,N_23801);
nor UO_845 (O_845,N_23639,N_22839);
nor UO_846 (O_846,N_23207,N_24314);
nor UO_847 (O_847,N_21985,N_23017);
nand UO_848 (O_848,N_24513,N_24017);
nand UO_849 (O_849,N_23588,N_23665);
and UO_850 (O_850,N_23201,N_22306);
nor UO_851 (O_851,N_23348,N_22806);
or UO_852 (O_852,N_23019,N_24759);
and UO_853 (O_853,N_24943,N_24218);
or UO_854 (O_854,N_22140,N_23294);
xnor UO_855 (O_855,N_22944,N_23202);
xnor UO_856 (O_856,N_23749,N_22271);
and UO_857 (O_857,N_22754,N_22031);
nor UO_858 (O_858,N_23583,N_22889);
or UO_859 (O_859,N_23110,N_23203);
or UO_860 (O_860,N_22645,N_24420);
and UO_861 (O_861,N_22844,N_22265);
nor UO_862 (O_862,N_24589,N_24883);
and UO_863 (O_863,N_24847,N_24906);
or UO_864 (O_864,N_22170,N_23570);
nand UO_865 (O_865,N_23666,N_22676);
nand UO_866 (O_866,N_22006,N_24131);
xor UO_867 (O_867,N_22809,N_22441);
nand UO_868 (O_868,N_22786,N_23737);
or UO_869 (O_869,N_23049,N_23989);
and UO_870 (O_870,N_23169,N_24414);
and UO_871 (O_871,N_23841,N_23107);
nor UO_872 (O_872,N_24428,N_23264);
xnor UO_873 (O_873,N_23909,N_23428);
xnor UO_874 (O_874,N_24702,N_24211);
nor UO_875 (O_875,N_23005,N_22609);
or UO_876 (O_876,N_23379,N_23597);
xnor UO_877 (O_877,N_22353,N_22442);
nand UO_878 (O_878,N_23571,N_22732);
nor UO_879 (O_879,N_23014,N_21908);
nor UO_880 (O_880,N_24326,N_22307);
or UO_881 (O_881,N_23037,N_23645);
xnor UO_882 (O_882,N_22506,N_23612);
nor UO_883 (O_883,N_24548,N_23575);
xor UO_884 (O_884,N_23176,N_22162);
nand UO_885 (O_885,N_22171,N_22653);
nor UO_886 (O_886,N_23879,N_24887);
or UO_887 (O_887,N_22403,N_24153);
nor UO_888 (O_888,N_22404,N_22986);
nand UO_889 (O_889,N_22281,N_22570);
xor UO_890 (O_890,N_24665,N_22887);
xnor UO_891 (O_891,N_22627,N_24375);
or UO_892 (O_892,N_23555,N_24703);
nand UO_893 (O_893,N_22102,N_24837);
nor UO_894 (O_894,N_23083,N_22128);
nand UO_895 (O_895,N_24427,N_24572);
nand UO_896 (O_896,N_22039,N_24573);
nor UO_897 (O_897,N_22876,N_22302);
xor UO_898 (O_898,N_24485,N_24037);
nor UO_899 (O_899,N_24596,N_24800);
xor UO_900 (O_900,N_22137,N_24697);
nand UO_901 (O_901,N_24599,N_23983);
xor UO_902 (O_902,N_24912,N_24613);
xnor UO_903 (O_903,N_24725,N_23825);
or UO_904 (O_904,N_21956,N_23910);
xnor UO_905 (O_905,N_23812,N_23799);
and UO_906 (O_906,N_22787,N_22446);
or UO_907 (O_907,N_22400,N_22416);
nor UO_908 (O_908,N_23963,N_22092);
nand UO_909 (O_909,N_24538,N_22536);
and UO_910 (O_910,N_23143,N_22282);
and UO_911 (O_911,N_23893,N_24192);
nor UO_912 (O_912,N_22135,N_22216);
or UO_913 (O_913,N_24142,N_22558);
nor UO_914 (O_914,N_22540,N_21962);
nor UO_915 (O_915,N_22421,N_24517);
nand UO_916 (O_916,N_22633,N_23773);
or UO_917 (O_917,N_23238,N_22301);
nor UO_918 (O_918,N_22207,N_21902);
nor UO_919 (O_919,N_22662,N_24240);
xnor UO_920 (O_920,N_24913,N_24612);
nor UO_921 (O_921,N_24751,N_23678);
or UO_922 (O_922,N_23882,N_23130);
or UO_923 (O_923,N_24908,N_21882);
xnor UO_924 (O_924,N_23907,N_22742);
or UO_925 (O_925,N_24892,N_24096);
nand UO_926 (O_926,N_24456,N_23060);
nand UO_927 (O_927,N_23619,N_23628);
nor UO_928 (O_928,N_24034,N_24023);
nand UO_929 (O_929,N_24180,N_22443);
nor UO_930 (O_930,N_22757,N_24844);
xnor UO_931 (O_931,N_23662,N_24797);
nand UO_932 (O_932,N_23164,N_23342);
and UO_933 (O_933,N_24974,N_24935);
nand UO_934 (O_934,N_21970,N_23592);
and UO_935 (O_935,N_21949,N_23100);
or UO_936 (O_936,N_23286,N_24531);
or UO_937 (O_937,N_23371,N_24856);
nand UO_938 (O_938,N_24251,N_24785);
xnor UO_939 (O_939,N_23533,N_22587);
and UO_940 (O_940,N_22828,N_23499);
or UO_941 (O_941,N_21984,N_22875);
or UO_942 (O_942,N_22620,N_22131);
and UO_943 (O_943,N_22846,N_24675);
or UO_944 (O_944,N_21957,N_22424);
or UO_945 (O_945,N_24660,N_23688);
nor UO_946 (O_946,N_23836,N_22641);
and UO_947 (O_947,N_24330,N_21992);
and UO_948 (O_948,N_22922,N_24998);
and UO_949 (O_949,N_23966,N_23887);
nor UO_950 (O_950,N_23308,N_23505);
or UO_951 (O_951,N_22865,N_24620);
or UO_952 (O_952,N_23191,N_22478);
xnor UO_953 (O_953,N_24679,N_22065);
or UO_954 (O_954,N_23092,N_22202);
xnor UO_955 (O_955,N_22826,N_24960);
xor UO_956 (O_956,N_24997,N_22200);
or UO_957 (O_957,N_24266,N_24078);
nand UO_958 (O_958,N_22284,N_23924);
or UO_959 (O_959,N_22642,N_21944);
xnor UO_960 (O_960,N_23573,N_23420);
xnor UO_961 (O_961,N_22898,N_22212);
or UO_962 (O_962,N_23847,N_23324);
or UO_963 (O_963,N_24480,N_23515);
and UO_964 (O_964,N_23209,N_23995);
and UO_965 (O_965,N_23511,N_24005);
or UO_966 (O_966,N_23718,N_22706);
nor UO_967 (O_967,N_23501,N_22851);
and UO_968 (O_968,N_24826,N_22320);
and UO_969 (O_969,N_22027,N_24888);
nor UO_970 (O_970,N_23831,N_23153);
xor UO_971 (O_971,N_22298,N_23440);
nand UO_972 (O_972,N_23259,N_22323);
nand UO_973 (O_973,N_21987,N_24199);
or UO_974 (O_974,N_22752,N_22449);
and UO_975 (O_975,N_24054,N_22119);
xor UO_976 (O_976,N_22116,N_23419);
and UO_977 (O_977,N_23979,N_23768);
and UO_978 (O_978,N_24478,N_22068);
xor UO_979 (O_979,N_24064,N_23869);
nand UO_980 (O_980,N_22644,N_24267);
or UO_981 (O_981,N_22089,N_22767);
or UO_982 (O_982,N_23157,N_22240);
and UO_983 (O_983,N_22709,N_24312);
xor UO_984 (O_984,N_23339,N_22704);
or UO_985 (O_985,N_24141,N_23132);
or UO_986 (O_986,N_22242,N_22021);
and UO_987 (O_987,N_23188,N_22072);
xnor UO_988 (O_988,N_23361,N_22681);
nor UO_989 (O_989,N_24500,N_22217);
and UO_990 (O_990,N_23747,N_22024);
nand UO_991 (O_991,N_21964,N_21967);
and UO_992 (O_992,N_24259,N_22906);
nor UO_993 (O_993,N_21951,N_24400);
and UO_994 (O_994,N_24799,N_23657);
nand UO_995 (O_995,N_24021,N_23774);
xnor UO_996 (O_996,N_22073,N_22868);
and UO_997 (O_997,N_23473,N_24453);
xor UO_998 (O_998,N_22090,N_22541);
xor UO_999 (O_999,N_22300,N_24230);
and UO_1000 (O_1000,N_22095,N_23994);
and UO_1001 (O_1001,N_23400,N_23694);
nor UO_1002 (O_1002,N_24338,N_22163);
or UO_1003 (O_1003,N_22261,N_24755);
and UO_1004 (O_1004,N_23585,N_24423);
nand UO_1005 (O_1005,N_23208,N_24764);
and UO_1006 (O_1006,N_23479,N_23884);
nor UO_1007 (O_1007,N_22420,N_24152);
xnor UO_1008 (O_1008,N_22715,N_23834);
xor UO_1009 (O_1009,N_24652,N_22504);
nor UO_1010 (O_1010,N_22569,N_24417);
and UO_1011 (O_1011,N_24909,N_22696);
nor UO_1012 (O_1012,N_22770,N_24383);
nand UO_1013 (O_1013,N_23252,N_23697);
or UO_1014 (O_1014,N_21995,N_24299);
or UO_1015 (O_1015,N_21996,N_22464);
nand UO_1016 (O_1016,N_22070,N_23472);
and UO_1017 (O_1017,N_22916,N_24696);
nand UO_1018 (O_1018,N_24914,N_23553);
and UO_1019 (O_1019,N_24994,N_22290);
or UO_1020 (O_1020,N_23603,N_22590);
and UO_1021 (O_1021,N_22480,N_23094);
nor UO_1022 (O_1022,N_22105,N_23854);
and UO_1023 (O_1023,N_22209,N_22197);
xor UO_1024 (O_1024,N_22934,N_21980);
nor UO_1025 (O_1025,N_24814,N_22960);
and UO_1026 (O_1026,N_22902,N_23340);
xnor UO_1027 (O_1027,N_23261,N_22719);
xor UO_1028 (O_1028,N_23231,N_23126);
xnor UO_1029 (O_1029,N_21889,N_24894);
or UO_1030 (O_1030,N_24786,N_24229);
nor UO_1031 (O_1031,N_22383,N_23150);
xor UO_1032 (O_1032,N_23066,N_23185);
and UO_1033 (O_1033,N_22186,N_23278);
or UO_1034 (O_1034,N_23817,N_22658);
nor UO_1035 (O_1035,N_24717,N_24492);
nor UO_1036 (O_1036,N_21971,N_24545);
and UO_1037 (O_1037,N_22438,N_24209);
or UO_1038 (O_1038,N_22509,N_23777);
nand UO_1039 (O_1039,N_22588,N_23908);
xnor UO_1040 (O_1040,N_24483,N_22482);
nand UO_1041 (O_1041,N_24900,N_22268);
or UO_1042 (O_1042,N_23013,N_22466);
and UO_1043 (O_1043,N_24404,N_24803);
and UO_1044 (O_1044,N_24070,N_23722);
nand UO_1045 (O_1045,N_22799,N_23051);
nand UO_1046 (O_1046,N_22274,N_23221);
or UO_1047 (O_1047,N_23328,N_22142);
nand UO_1048 (O_1048,N_23528,N_23918);
nor UO_1049 (O_1049,N_24535,N_22904);
xnor UO_1050 (O_1050,N_23911,N_22327);
xnor UO_1051 (O_1051,N_21919,N_24578);
nor UO_1052 (O_1052,N_23594,N_21988);
nand UO_1053 (O_1053,N_24027,N_22429);
or UO_1054 (O_1054,N_24006,N_22259);
and UO_1055 (O_1055,N_22717,N_22823);
or UO_1056 (O_1056,N_22147,N_24112);
nor UO_1057 (O_1057,N_22343,N_23240);
and UO_1058 (O_1058,N_24438,N_24235);
and UO_1059 (O_1059,N_22948,N_23405);
or UO_1060 (O_1060,N_22580,N_23297);
nor UO_1061 (O_1061,N_22896,N_24739);
nor UO_1062 (O_1062,N_22344,N_24848);
xnor UO_1063 (O_1063,N_24208,N_24683);
and UO_1064 (O_1064,N_24976,N_23950);
nand UO_1065 (O_1065,N_23086,N_23211);
and UO_1066 (O_1066,N_24966,N_23970);
nor UO_1067 (O_1067,N_22107,N_24327);
nor UO_1068 (O_1068,N_22336,N_23426);
nor UO_1069 (O_1069,N_24331,N_23954);
nand UO_1070 (O_1070,N_23497,N_23875);
or UO_1071 (O_1071,N_24874,N_24930);
nand UO_1072 (O_1072,N_23653,N_24932);
and UO_1073 (O_1073,N_22195,N_23026);
nor UO_1074 (O_1074,N_22689,N_24433);
nor UO_1075 (O_1075,N_24125,N_21924);
and UO_1076 (O_1076,N_22164,N_24407);
nor UO_1077 (O_1077,N_23262,N_23028);
or UO_1078 (O_1078,N_21945,N_23698);
nand UO_1079 (O_1079,N_24957,N_24857);
nand UO_1080 (O_1080,N_23818,N_23483);
xnor UO_1081 (O_1081,N_24477,N_24555);
nor UO_1082 (O_1082,N_23163,N_23038);
or UO_1083 (O_1083,N_22020,N_23398);
or UO_1084 (O_1084,N_24936,N_22337);
nor UO_1085 (O_1085,N_23393,N_21910);
xnor UO_1086 (O_1086,N_24045,N_23354);
or UO_1087 (O_1087,N_23050,N_22289);
or UO_1088 (O_1088,N_22738,N_24322);
or UO_1089 (O_1089,N_24646,N_24642);
xor UO_1090 (O_1090,N_24923,N_22004);
or UO_1091 (O_1091,N_24409,N_22707);
xnor UO_1092 (O_1092,N_24669,N_24719);
xnor UO_1093 (O_1093,N_23508,N_23862);
nor UO_1094 (O_1094,N_21943,N_24850);
and UO_1095 (O_1095,N_24246,N_22756);
and UO_1096 (O_1096,N_22539,N_24130);
xor UO_1097 (O_1097,N_21879,N_24353);
nand UO_1098 (O_1098,N_22807,N_24831);
nor UO_1099 (O_1099,N_22961,N_22083);
or UO_1100 (O_1100,N_23495,N_22132);
nand UO_1101 (O_1101,N_24363,N_22419);
xnor UO_1102 (O_1102,N_22655,N_24278);
nand UO_1103 (O_1103,N_23168,N_24033);
nor UO_1104 (O_1104,N_24948,N_24341);
nor UO_1105 (O_1105,N_23189,N_22774);
nand UO_1106 (O_1106,N_23778,N_22104);
nand UO_1107 (O_1107,N_23141,N_22589);
or UO_1108 (O_1108,N_24072,N_24672);
or UO_1109 (O_1109,N_24766,N_23853);
nand UO_1110 (O_1110,N_22908,N_24507);
or UO_1111 (O_1111,N_23958,N_24735);
or UO_1112 (O_1112,N_23387,N_24140);
nor UO_1113 (O_1113,N_23438,N_22262);
nor UO_1114 (O_1114,N_23789,N_23431);
or UO_1115 (O_1115,N_23672,N_22794);
nor UO_1116 (O_1116,N_24173,N_24977);
nand UO_1117 (O_1117,N_23514,N_22063);
nand UO_1118 (O_1118,N_23384,N_24834);
nand UO_1119 (O_1119,N_22448,N_24802);
nor UO_1120 (O_1120,N_22976,N_23635);
xnor UO_1121 (O_1121,N_22098,N_24917);
nand UO_1122 (O_1122,N_24306,N_22697);
nor UO_1123 (O_1123,N_22278,N_23706);
nor UO_1124 (O_1124,N_24496,N_24846);
and UO_1125 (O_1125,N_24366,N_24788);
or UO_1126 (O_1126,N_23674,N_23364);
nor UO_1127 (O_1127,N_23719,N_23076);
nor UO_1128 (O_1128,N_24399,N_21973);
xnor UO_1129 (O_1129,N_22339,N_24989);
xnor UO_1130 (O_1130,N_22071,N_23217);
nor UO_1131 (O_1131,N_22060,N_22744);
and UO_1132 (O_1132,N_22852,N_24983);
nand UO_1133 (O_1133,N_22994,N_23243);
nor UO_1134 (O_1134,N_23844,N_24431);
and UO_1135 (O_1135,N_23052,N_21921);
or UO_1136 (O_1136,N_22854,N_24429);
nor UO_1137 (O_1137,N_23531,N_23469);
nor UO_1138 (O_1138,N_24204,N_23068);
and UO_1139 (O_1139,N_23673,N_22985);
nor UO_1140 (O_1140,N_22603,N_24674);
nor UO_1141 (O_1141,N_22795,N_22257);
nor UO_1142 (O_1142,N_23456,N_22971);
nor UO_1143 (O_1143,N_22952,N_24354);
or UO_1144 (O_1144,N_24443,N_22979);
nor UO_1145 (O_1145,N_22379,N_24247);
xnor UO_1146 (O_1146,N_23900,N_22808);
nand UO_1147 (O_1147,N_23265,N_24926);
nand UO_1148 (O_1148,N_24075,N_23559);
xnor UO_1149 (O_1149,N_23048,N_23512);
nand UO_1150 (O_1150,N_23123,N_21942);
nor UO_1151 (O_1151,N_22995,N_24073);
and UO_1152 (O_1152,N_24317,N_24138);
xor UO_1153 (O_1153,N_23915,N_24243);
nand UO_1154 (O_1154,N_22785,N_24318);
nor UO_1155 (O_1155,N_24920,N_22548);
xor UO_1156 (O_1156,N_22596,N_23548);
and UO_1157 (O_1157,N_23181,N_22690);
nand UO_1158 (O_1158,N_24952,N_22537);
nor UO_1159 (O_1159,N_24370,N_22219);
nor UO_1160 (O_1160,N_23886,N_24758);
nor UO_1161 (O_1161,N_24655,N_22388);
xor UO_1162 (O_1162,N_24771,N_21884);
nor UO_1163 (O_1163,N_23442,N_22834);
xor UO_1164 (O_1164,N_23542,N_22044);
nand UO_1165 (O_1165,N_22297,N_23973);
nand UO_1166 (O_1166,N_22556,N_22141);
nand UO_1167 (O_1167,N_22033,N_22778);
and UO_1168 (O_1168,N_23987,N_23239);
nand UO_1169 (O_1169,N_24461,N_22465);
xnor UO_1170 (O_1170,N_23922,N_23016);
nand UO_1171 (O_1171,N_23041,N_24220);
xor UO_1172 (O_1172,N_23590,N_24780);
or UO_1173 (O_1173,N_24891,N_22064);
xor UO_1174 (O_1174,N_24647,N_24056);
nand UO_1175 (O_1175,N_22901,N_23247);
nor UO_1176 (O_1176,N_23372,N_24927);
or UO_1177 (O_1177,N_24849,N_23868);
nand UO_1178 (O_1178,N_24044,N_24968);
or UO_1179 (O_1179,N_23810,N_22840);
and UO_1180 (O_1180,N_24449,N_22518);
and UO_1181 (O_1181,N_22167,N_23158);
or UO_1182 (O_1182,N_24108,N_23920);
nand UO_1183 (O_1183,N_23241,N_21898);
and UO_1184 (O_1184,N_24645,N_24432);
xnor UO_1185 (O_1185,N_22287,N_22926);
nand UO_1186 (O_1186,N_23807,N_23578);
or UO_1187 (O_1187,N_22314,N_22973);
nand UO_1188 (O_1188,N_23452,N_24282);
and UO_1189 (O_1189,N_23070,N_22811);
nor UO_1190 (O_1190,N_23033,N_22735);
nor UO_1191 (O_1191,N_22168,N_22258);
xor UO_1192 (O_1192,N_23485,N_24897);
or UO_1193 (O_1193,N_24925,N_23402);
nand UO_1194 (O_1194,N_22295,N_23752);
or UO_1195 (O_1195,N_21948,N_24773);
nand UO_1196 (O_1196,N_22515,N_22228);
nor UO_1197 (O_1197,N_23955,N_24320);
nor UO_1198 (O_1198,N_24519,N_23121);
xor UO_1199 (O_1199,N_22250,N_22100);
and UO_1200 (O_1200,N_23629,N_24343);
xor UO_1201 (O_1201,N_24934,N_23878);
and UO_1202 (O_1202,N_24133,N_23938);
and UO_1203 (O_1203,N_23554,N_22993);
xnor UO_1204 (O_1204,N_22407,N_22292);
and UO_1205 (O_1205,N_24754,N_22205);
nor UO_1206 (O_1206,N_23461,N_23873);
nor UO_1207 (O_1207,N_22182,N_21887);
and UO_1208 (O_1208,N_23753,N_23210);
xor UO_1209 (O_1209,N_23865,N_23413);
or UO_1210 (O_1210,N_23113,N_23968);
and UO_1211 (O_1211,N_21916,N_23270);
nor UO_1212 (O_1212,N_22470,N_22853);
nand UO_1213 (O_1213,N_22678,N_24503);
xor UO_1214 (O_1214,N_24933,N_23880);
xor UO_1215 (O_1215,N_22812,N_22888);
nor UO_1216 (O_1216,N_23723,N_23833);
nand UO_1217 (O_1217,N_23192,N_22133);
and UO_1218 (O_1218,N_22156,N_23519);
nand UO_1219 (O_1219,N_21903,N_22650);
and UO_1220 (O_1220,N_23572,N_22562);
or UO_1221 (O_1221,N_23726,N_23040);
xor UO_1222 (O_1222,N_24227,N_24176);
or UO_1223 (O_1223,N_23404,N_24465);
nand UO_1224 (O_1224,N_23527,N_22172);
nor UO_1225 (O_1225,N_24763,N_23762);
or UO_1226 (O_1226,N_22395,N_21904);
xor UO_1227 (O_1227,N_22818,N_23422);
nor UO_1228 (O_1228,N_22191,N_23079);
xnor UO_1229 (O_1229,N_23721,N_24263);
nand UO_1230 (O_1230,N_24187,N_22762);
or UO_1231 (O_1231,N_24424,N_22193);
and UO_1232 (O_1232,N_24576,N_24484);
nand UO_1233 (O_1233,N_22552,N_24988);
or UO_1234 (O_1234,N_22082,N_23897);
nand UO_1235 (O_1235,N_22123,N_24574);
xor UO_1236 (O_1236,N_22232,N_22718);
xor UO_1237 (O_1237,N_24819,N_22227);
and UO_1238 (O_1238,N_22382,N_22460);
nor UO_1239 (O_1239,N_23586,N_23449);
nand UO_1240 (O_1240,N_22947,N_22427);
nand UO_1241 (O_1241,N_24528,N_24550);
nor UO_1242 (O_1242,N_22332,N_24050);
nor UO_1243 (O_1243,N_22728,N_23659);
or UO_1244 (O_1244,N_22591,N_22810);
and UO_1245 (O_1245,N_21983,N_22367);
nand UO_1246 (O_1246,N_23133,N_24833);
nand UO_1247 (O_1247,N_24713,N_22108);
nand UO_1248 (O_1248,N_24336,N_22431);
or UO_1249 (O_1249,N_22139,N_23517);
xnor UO_1250 (O_1250,N_24873,N_24062);
or UO_1251 (O_1251,N_23822,N_22544);
nor UO_1252 (O_1252,N_23758,N_22695);
and UO_1253 (O_1253,N_22668,N_24334);
and UO_1254 (O_1254,N_22308,N_24452);
and UO_1255 (O_1255,N_24110,N_23984);
and UO_1256 (O_1256,N_22969,N_23064);
or UO_1257 (O_1257,N_22629,N_24607);
or UO_1258 (O_1258,N_21899,N_23434);
and UO_1259 (O_1259,N_23167,N_23055);
nand UO_1260 (O_1260,N_22273,N_23071);
xnor UO_1261 (O_1261,N_24127,N_24128);
nand UO_1262 (O_1262,N_23830,N_23237);
nor UO_1263 (O_1263,N_23031,N_24117);
xnor UO_1264 (O_1264,N_23417,N_24055);
nor UO_1265 (O_1265,N_24584,N_21982);
and UO_1266 (O_1266,N_22074,N_23829);
and UO_1267 (O_1267,N_22066,N_22827);
and UO_1268 (O_1268,N_24498,N_24258);
and UO_1269 (O_1269,N_24099,N_24712);
nand UO_1270 (O_1270,N_22782,N_24867);
and UO_1271 (O_1271,N_22293,N_24749);
xnor UO_1272 (O_1272,N_22467,N_23504);
and UO_1273 (O_1273,N_23482,N_22126);
or UO_1274 (O_1274,N_24859,N_23415);
and UO_1275 (O_1275,N_21891,N_23993);
nor UO_1276 (O_1276,N_22923,N_24311);
nand UO_1277 (O_1277,N_22475,N_23116);
or UO_1278 (O_1278,N_22138,N_23945);
nand UO_1279 (O_1279,N_23738,N_22831);
and UO_1280 (O_1280,N_23468,N_23411);
nand UO_1281 (O_1281,N_23484,N_22527);
nand UO_1282 (O_1282,N_22311,N_24196);
nand UO_1283 (O_1283,N_22052,N_23676);
nor UO_1284 (O_1284,N_23409,N_22013);
and UO_1285 (O_1285,N_23427,N_22198);
xnor UO_1286 (O_1286,N_23144,N_23139);
and UO_1287 (O_1287,N_23871,N_23363);
nor UO_1288 (O_1288,N_22739,N_23432);
or UO_1289 (O_1289,N_23246,N_22730);
and UO_1290 (O_1290,N_23682,N_23216);
nand UO_1291 (O_1291,N_24305,N_23292);
xor UO_1292 (O_1292,N_24521,N_23165);
nand UO_1293 (O_1293,N_22215,N_24695);
or UO_1294 (O_1294,N_24809,N_23558);
or UO_1295 (O_1295,N_23299,N_23327);
xor UO_1296 (O_1296,N_23580,N_24962);
nor UO_1297 (O_1297,N_23670,N_23899);
nor UO_1298 (O_1298,N_24043,N_23439);
and UO_1299 (O_1299,N_24435,N_22331);
xor UO_1300 (O_1300,N_23325,N_24272);
nand UO_1301 (O_1301,N_24745,N_22612);
or UO_1302 (O_1302,N_23872,N_22632);
nor UO_1303 (O_1303,N_24277,N_24778);
xnor UO_1304 (O_1304,N_24855,N_24283);
or UO_1305 (O_1305,N_23598,N_23444);
nand UO_1306 (O_1306,N_24249,N_23451);
nor UO_1307 (O_1307,N_22468,N_24877);
nand UO_1308 (O_1308,N_22561,N_23902);
nand UO_1309 (O_1309,N_22075,N_24654);
and UO_1310 (O_1310,N_24581,N_24462);
xnor UO_1311 (O_1311,N_22885,N_24685);
and UO_1312 (O_1312,N_24737,N_24295);
or UO_1313 (O_1313,N_24684,N_22051);
or UO_1314 (O_1314,N_23953,N_24842);
nand UO_1315 (O_1315,N_22915,N_23253);
nor UO_1316 (O_1316,N_23148,N_24348);
xnor UO_1317 (O_1317,N_23333,N_23053);
or UO_1318 (O_1318,N_22815,N_22581);
or UO_1319 (O_1319,N_22148,N_24228);
xor UO_1320 (O_1320,N_24789,N_24823);
or UO_1321 (O_1321,N_22023,N_22372);
and UO_1322 (O_1322,N_24929,N_23943);
nand UO_1323 (O_1323,N_22510,N_23885);
and UO_1324 (O_1324,N_22930,N_23488);
and UO_1325 (O_1325,N_22519,N_22646);
and UO_1326 (O_1326,N_23323,N_23632);
or UO_1327 (O_1327,N_22978,N_22682);
nand UO_1328 (O_1328,N_24910,N_22622);
xor UO_1329 (O_1329,N_23741,N_24185);
xor UO_1330 (O_1330,N_24084,N_23705);
xor UO_1331 (O_1331,N_24287,N_23249);
nor UO_1332 (O_1332,N_23160,N_23999);
and UO_1333 (O_1333,N_22659,N_24335);
and UO_1334 (O_1334,N_22366,N_24113);
xnor UO_1335 (O_1335,N_21979,N_23975);
xor UO_1336 (O_1336,N_22017,N_23219);
and UO_1337 (O_1337,N_23111,N_22983);
or UO_1338 (O_1338,N_22669,N_22410);
or UO_1339 (O_1339,N_23602,N_21878);
xor UO_1340 (O_1340,N_22408,N_22939);
or UO_1341 (O_1341,N_24959,N_23198);
xnor UO_1342 (O_1342,N_22169,N_22749);
xnor UO_1343 (O_1343,N_24014,N_22631);
xor UO_1344 (O_1344,N_23154,N_22745);
nand UO_1345 (O_1345,N_24921,N_23929);
and UO_1346 (O_1346,N_22578,N_23196);
nor UO_1347 (O_1347,N_22458,N_23663);
nor UO_1348 (O_1348,N_23326,N_24376);
or UO_1349 (O_1349,N_24781,N_22495);
nand UO_1350 (O_1350,N_23633,N_23944);
nor UO_1351 (O_1351,N_24772,N_24543);
and UO_1352 (O_1352,N_22173,N_22450);
xor UO_1353 (O_1353,N_21989,N_22608);
nand UO_1354 (O_1354,N_23587,N_23009);
and UO_1355 (O_1355,N_23660,N_23724);
nor UO_1356 (O_1356,N_23152,N_24811);
nor UO_1357 (O_1357,N_22640,N_21913);
xnor UO_1358 (O_1358,N_22472,N_24757);
nor UO_1359 (O_1359,N_21895,N_23734);
nand UO_1360 (O_1360,N_22243,N_24608);
nand UO_1361 (O_1361,N_24549,N_22433);
nor UO_1362 (O_1362,N_22143,N_22579);
nor UO_1363 (O_1363,N_23314,N_22434);
xnor UO_1364 (O_1364,N_22959,N_23454);
and UO_1365 (O_1365,N_24003,N_22511);
nand UO_1366 (O_1366,N_24709,N_23547);
or UO_1367 (O_1367,N_23368,N_22599);
nand UO_1368 (O_1368,N_24419,N_23858);
nor UO_1369 (O_1369,N_24371,N_21961);
nor UO_1370 (O_1370,N_24111,N_23845);
or UO_1371 (O_1371,N_23745,N_23225);
and UO_1372 (O_1372,N_22529,N_23805);
nor UO_1373 (O_1373,N_22914,N_22486);
nor UO_1374 (O_1374,N_24451,N_24996);
or UO_1375 (O_1375,N_22032,N_23903);
nor UO_1376 (O_1376,N_22221,N_24860);
xnor UO_1377 (O_1377,N_23245,N_24090);
nor UO_1378 (O_1378,N_24321,N_24740);
nor UO_1379 (O_1379,N_22253,N_23156);
or UO_1380 (O_1380,N_21958,N_23730);
and UO_1381 (O_1381,N_22814,N_23125);
nand UO_1382 (O_1382,N_22180,N_23437);
nor UO_1383 (O_1383,N_23617,N_24682);
xnor UO_1384 (O_1384,N_22763,N_22557);
nor UO_1385 (O_1385,N_22490,N_23582);
and UO_1386 (O_1386,N_22223,N_23541);
nor UO_1387 (O_1387,N_22340,N_22726);
or UO_1388 (O_1388,N_23289,N_24526);
or UO_1389 (O_1389,N_24769,N_22150);
and UO_1390 (O_1390,N_22747,N_22911);
nor UO_1391 (O_1391,N_23623,N_22954);
xnor UO_1392 (O_1392,N_24425,N_24969);
xnor UO_1393 (O_1393,N_24198,N_24364);
or UO_1394 (O_1394,N_24955,N_24264);
xnor UO_1395 (O_1395,N_22613,N_22484);
nand UO_1396 (O_1396,N_24026,N_22012);
nand UO_1397 (O_1397,N_22025,N_23715);
nor UO_1398 (O_1398,N_21975,N_24444);
nand UO_1399 (O_1399,N_22731,N_23220);
or UO_1400 (O_1400,N_24835,N_24217);
or UO_1401 (O_1401,N_24680,N_23161);
nand UO_1402 (O_1402,N_22166,N_21897);
xnor UO_1403 (O_1403,N_23276,N_22931);
or UO_1404 (O_1404,N_22586,N_22231);
xor UO_1405 (O_1405,N_23460,N_23649);
or UO_1406 (O_1406,N_24971,N_22957);
nor UO_1407 (O_1407,N_22000,N_21905);
or UO_1408 (O_1408,N_24403,N_24653);
and UO_1409 (O_1409,N_23919,N_24868);
nor UO_1410 (O_1410,N_22048,N_23690);
or UO_1411 (O_1411,N_24308,N_23366);
nor UO_1412 (O_1412,N_24542,N_24257);
or UO_1413 (O_1413,N_22649,N_22688);
nand UO_1414 (O_1414,N_24081,N_22457);
xnor UO_1415 (O_1415,N_24686,N_24223);
nand UO_1416 (O_1416,N_22698,N_22299);
nand UO_1417 (O_1417,N_23115,N_22773);
nand UO_1418 (O_1418,N_22524,N_24028);
nand UO_1419 (O_1419,N_24551,N_24074);
or UO_1420 (O_1420,N_21893,N_23162);
nor UO_1421 (O_1421,N_22877,N_24570);
nand UO_1422 (O_1422,N_24579,N_23622);
nand UO_1423 (O_1423,N_22034,N_23669);
nand UO_1424 (O_1424,N_23389,N_23416);
and UO_1425 (O_1425,N_22263,N_22833);
xor UO_1426 (O_1426,N_24356,N_23642);
xnor UO_1427 (O_1427,N_24369,N_23928);
nand UO_1428 (O_1428,N_23043,N_23355);
nor UO_1429 (O_1429,N_24964,N_22010);
nor UO_1430 (O_1430,N_23655,N_24024);
nand UO_1431 (O_1431,N_23608,N_23407);
nor UO_1432 (O_1432,N_23318,N_24524);
xnor UO_1433 (O_1433,N_23746,N_23046);
xor UO_1434 (O_1434,N_22542,N_24284);
and UO_1435 (O_1435,N_22489,N_24232);
nor UO_1436 (O_1436,N_22334,N_22417);
xnor UO_1437 (O_1437,N_23851,N_22950);
and UO_1438 (O_1438,N_22657,N_22113);
nand UO_1439 (O_1439,N_21955,N_24730);
xnor UO_1440 (O_1440,N_22049,N_22251);
nor UO_1441 (O_1441,N_24486,N_24351);
xor UO_1442 (O_1442,N_24603,N_22175);
nor UO_1443 (O_1443,N_24164,N_23367);
or UO_1444 (O_1444,N_24677,N_22894);
nor UO_1445 (O_1445,N_22781,N_24387);
or UO_1446 (O_1446,N_22080,N_24852);
nor UO_1447 (O_1447,N_23478,N_23358);
xnor UO_1448 (O_1448,N_23084,N_24269);
and UO_1449 (O_1449,N_23840,N_22584);
and UO_1450 (O_1450,N_23105,N_23080);
nor UO_1451 (O_1451,N_24560,N_24992);
nor UO_1452 (O_1452,N_22520,N_23074);
nor UO_1453 (O_1453,N_23453,N_22593);
nand UO_1454 (O_1454,N_24838,N_24546);
and UO_1455 (O_1455,N_22114,N_24310);
nand UO_1456 (O_1456,N_24214,N_23114);
or UO_1457 (O_1457,N_22210,N_23699);
or UO_1458 (O_1458,N_22179,N_24747);
nand UO_1459 (O_1459,N_23720,N_22538);
xor UO_1460 (O_1460,N_23567,N_22283);
nor UO_1461 (O_1461,N_22841,N_24440);
nand UO_1462 (O_1462,N_24843,N_24624);
or UO_1463 (O_1463,N_23781,N_23012);
or UO_1464 (O_1464,N_22352,N_22437);
or UO_1465 (O_1465,N_22855,N_22187);
or UO_1466 (O_1466,N_22236,N_24756);
or UO_1467 (O_1467,N_22951,N_22577);
and UO_1468 (O_1468,N_24509,N_24676);
or UO_1469 (O_1469,N_24200,N_22094);
nand UO_1470 (O_1470,N_23242,N_23448);
xor UO_1471 (O_1471,N_24105,N_23988);
or UO_1472 (O_1472,N_24956,N_24822);
or UO_1473 (O_1473,N_23380,N_22881);
nand UO_1474 (O_1474,N_22055,N_23901);
xnor UO_1475 (O_1475,N_21978,N_22335);
nand UO_1476 (O_1476,N_24738,N_23735);
or UO_1477 (O_1477,N_24704,N_24824);
nand UO_1478 (O_1478,N_23896,N_23450);
or UO_1479 (O_1479,N_24286,N_22729);
xnor UO_1480 (O_1480,N_24710,N_22067);
xnor UO_1481 (O_1481,N_23626,N_23965);
nor UO_1482 (O_1482,N_23197,N_22222);
xor UO_1483 (O_1483,N_23912,N_23463);
xnor UO_1484 (O_1484,N_22545,N_24666);
nand UO_1485 (O_1485,N_24627,N_23058);
and UO_1486 (O_1486,N_24947,N_23521);
and UO_1487 (O_1487,N_22097,N_23112);
nand UO_1488 (O_1488,N_24231,N_24592);
nor UO_1489 (O_1489,N_24109,N_21915);
and UO_1490 (O_1490,N_23312,N_22189);
xnor UO_1491 (O_1491,N_23787,N_23518);
and UO_1492 (O_1492,N_24162,N_22309);
xor UO_1493 (O_1493,N_23552,N_22492);
nand UO_1494 (O_1494,N_23477,N_24602);
xnor UO_1495 (O_1495,N_22249,N_22924);
xor UO_1496 (O_1496,N_22893,N_23180);
nand UO_1497 (O_1497,N_24559,N_24188);
or UO_1498 (O_1498,N_22047,N_22439);
or UO_1499 (O_1499,N_22929,N_22503);
or UO_1500 (O_1500,N_21991,N_23436);
nor UO_1501 (O_1501,N_23359,N_22665);
and UO_1502 (O_1502,N_24146,N_21950);
xnor UO_1503 (O_1503,N_22532,N_24136);
and UO_1504 (O_1504,N_22291,N_23251);
nor UO_1505 (O_1505,N_24018,N_22521);
and UO_1506 (O_1506,N_24597,N_22455);
or UO_1507 (O_1507,N_22360,N_22703);
or UO_1508 (O_1508,N_24411,N_24514);
xnor UO_1509 (O_1509,N_24622,N_24385);
nand UO_1510 (O_1510,N_22321,N_23828);
or UO_1511 (O_1511,N_22582,N_22029);
or UO_1512 (O_1512,N_24390,N_22574);
or UO_1513 (O_1513,N_22546,N_21940);
or UO_1514 (O_1514,N_23065,N_24206);
nor UO_1515 (O_1515,N_22513,N_23736);
xor UO_1516 (O_1516,N_24658,N_23321);
nand UO_1517 (O_1517,N_24638,N_22328);
nand UO_1518 (O_1518,N_22871,N_22528);
and UO_1519 (O_1519,N_24170,N_22096);
or UO_1520 (O_1520,N_24398,N_22654);
xnor UO_1521 (O_1521,N_22134,N_22997);
nor UO_1522 (O_1522,N_23991,N_24340);
or UO_1523 (O_1523,N_22225,N_24116);
and UO_1524 (O_1524,N_22935,N_24455);
and UO_1525 (O_1525,N_22008,N_22533);
and UO_1526 (O_1526,N_23190,N_23714);
nor UO_1527 (O_1527,N_22159,N_24053);
or UO_1528 (O_1528,N_23819,N_23492);
nand UO_1529 (O_1529,N_22573,N_23607);
nand UO_1530 (O_1530,N_22943,N_24569);
and UO_1531 (O_1531,N_23636,N_22598);
nand UO_1532 (O_1532,N_22624,N_24098);
nor UO_1533 (O_1533,N_22720,N_23131);
and UO_1534 (O_1534,N_22087,N_22701);
xnor UO_1535 (O_1535,N_22568,N_21993);
nor UO_1536 (O_1536,N_21928,N_23082);
and UO_1537 (O_1537,N_24979,N_23234);
nand UO_1538 (O_1538,N_24609,N_23683);
nor UO_1539 (O_1539,N_24588,N_23638);
nand UO_1540 (O_1540,N_24736,N_24941);
or UO_1541 (O_1541,N_22611,N_24776);
or UO_1542 (O_1542,N_23464,N_24447);
nor UO_1543 (O_1543,N_23770,N_22972);
and UO_1544 (O_1544,N_23336,N_22919);
or UO_1545 (O_1545,N_22936,N_24893);
nand UO_1546 (O_1546,N_24202,N_24052);
and UO_1547 (O_1547,N_23534,N_24825);
nor UO_1548 (O_1548,N_24791,N_24742);
nand UO_1549 (O_1549,N_24265,N_22239);
nor UO_1550 (O_1550,N_22112,N_22093);
and UO_1551 (O_1551,N_22161,N_23228);
and UO_1552 (O_1552,N_22615,N_23614);
or UO_1553 (O_1553,N_24307,N_24463);
xor UO_1554 (O_1554,N_24687,N_23254);
xor UO_1555 (O_1555,N_24301,N_24158);
xor UO_1556 (O_1556,N_23059,N_23784);
nor UO_1557 (O_1557,N_23615,N_22783);
nor UO_1558 (O_1558,N_24631,N_23769);
nand UO_1559 (O_1559,N_24681,N_23791);
xor UO_1560 (O_1560,N_24080,N_24777);
or UO_1561 (O_1561,N_24032,N_21952);
xor UO_1562 (O_1562,N_24861,N_22827);
nand UO_1563 (O_1563,N_24849,N_23965);
or UO_1564 (O_1564,N_23097,N_22082);
or UO_1565 (O_1565,N_24110,N_22865);
nor UO_1566 (O_1566,N_22440,N_23325);
nor UO_1567 (O_1567,N_23312,N_23081);
xnor UO_1568 (O_1568,N_22406,N_24309);
or UO_1569 (O_1569,N_24051,N_23248);
and UO_1570 (O_1570,N_22160,N_24369);
nand UO_1571 (O_1571,N_22130,N_23734);
and UO_1572 (O_1572,N_24825,N_23401);
xnor UO_1573 (O_1573,N_22357,N_24147);
and UO_1574 (O_1574,N_24777,N_24503);
nand UO_1575 (O_1575,N_24860,N_23761);
or UO_1576 (O_1576,N_24993,N_23773);
or UO_1577 (O_1577,N_21952,N_22857);
and UO_1578 (O_1578,N_23733,N_21993);
nor UO_1579 (O_1579,N_22152,N_24540);
nand UO_1580 (O_1580,N_24545,N_22386);
and UO_1581 (O_1581,N_22639,N_21935);
or UO_1582 (O_1582,N_24144,N_24180);
nor UO_1583 (O_1583,N_22805,N_22827);
nand UO_1584 (O_1584,N_23434,N_23022);
nand UO_1585 (O_1585,N_23164,N_22045);
nor UO_1586 (O_1586,N_23573,N_22944);
or UO_1587 (O_1587,N_22457,N_21979);
nand UO_1588 (O_1588,N_21998,N_23185);
nand UO_1589 (O_1589,N_22717,N_22534);
nand UO_1590 (O_1590,N_21905,N_23838);
and UO_1591 (O_1591,N_22053,N_23396);
nor UO_1592 (O_1592,N_22530,N_24138);
nand UO_1593 (O_1593,N_23275,N_23638);
nand UO_1594 (O_1594,N_22462,N_23166);
xnor UO_1595 (O_1595,N_22149,N_23988);
nor UO_1596 (O_1596,N_24514,N_23970);
or UO_1597 (O_1597,N_24427,N_23198);
xnor UO_1598 (O_1598,N_24408,N_24215);
and UO_1599 (O_1599,N_22763,N_24471);
nor UO_1600 (O_1600,N_24250,N_24590);
or UO_1601 (O_1601,N_23959,N_21978);
xor UO_1602 (O_1602,N_24994,N_22767);
and UO_1603 (O_1603,N_22192,N_23404);
nand UO_1604 (O_1604,N_23156,N_22229);
nand UO_1605 (O_1605,N_23828,N_24110);
xor UO_1606 (O_1606,N_22983,N_22278);
nand UO_1607 (O_1607,N_22532,N_24615);
nor UO_1608 (O_1608,N_24114,N_22025);
nor UO_1609 (O_1609,N_23313,N_23643);
xor UO_1610 (O_1610,N_22706,N_23630);
or UO_1611 (O_1611,N_22236,N_21914);
nand UO_1612 (O_1612,N_22735,N_22900);
xor UO_1613 (O_1613,N_22642,N_22513);
or UO_1614 (O_1614,N_23292,N_24934);
xor UO_1615 (O_1615,N_23001,N_24165);
nor UO_1616 (O_1616,N_24916,N_22778);
xnor UO_1617 (O_1617,N_22386,N_24138);
or UO_1618 (O_1618,N_23240,N_22634);
and UO_1619 (O_1619,N_21889,N_23729);
nand UO_1620 (O_1620,N_24667,N_22854);
xor UO_1621 (O_1621,N_23356,N_24278);
nand UO_1622 (O_1622,N_22941,N_22296);
nor UO_1623 (O_1623,N_24239,N_21979);
nor UO_1624 (O_1624,N_22763,N_24362);
nor UO_1625 (O_1625,N_23378,N_22273);
nand UO_1626 (O_1626,N_24342,N_23614);
nand UO_1627 (O_1627,N_24422,N_22299);
or UO_1628 (O_1628,N_22992,N_24365);
and UO_1629 (O_1629,N_22882,N_22852);
or UO_1630 (O_1630,N_22973,N_24802);
nand UO_1631 (O_1631,N_24800,N_24257);
xor UO_1632 (O_1632,N_22088,N_22099);
or UO_1633 (O_1633,N_24416,N_24446);
or UO_1634 (O_1634,N_24054,N_23365);
and UO_1635 (O_1635,N_23725,N_22260);
nor UO_1636 (O_1636,N_22386,N_23216);
nand UO_1637 (O_1637,N_24430,N_22106);
xnor UO_1638 (O_1638,N_24781,N_23377);
xnor UO_1639 (O_1639,N_23664,N_22973);
nand UO_1640 (O_1640,N_22458,N_24655);
xnor UO_1641 (O_1641,N_23469,N_22207);
xnor UO_1642 (O_1642,N_22135,N_22400);
xor UO_1643 (O_1643,N_23956,N_23510);
or UO_1644 (O_1644,N_21898,N_24849);
or UO_1645 (O_1645,N_23064,N_24225);
nand UO_1646 (O_1646,N_21935,N_24710);
nor UO_1647 (O_1647,N_24144,N_24652);
xnor UO_1648 (O_1648,N_23431,N_22218);
and UO_1649 (O_1649,N_24209,N_22712);
xnor UO_1650 (O_1650,N_22683,N_23490);
and UO_1651 (O_1651,N_23850,N_24599);
or UO_1652 (O_1652,N_24554,N_21993);
or UO_1653 (O_1653,N_24070,N_23665);
and UO_1654 (O_1654,N_24369,N_24222);
nor UO_1655 (O_1655,N_22851,N_21893);
xor UO_1656 (O_1656,N_23662,N_24182);
and UO_1657 (O_1657,N_24122,N_23778);
nor UO_1658 (O_1658,N_24155,N_24588);
xor UO_1659 (O_1659,N_22254,N_22316);
nand UO_1660 (O_1660,N_23230,N_23574);
nand UO_1661 (O_1661,N_23044,N_22449);
nand UO_1662 (O_1662,N_24177,N_23877);
and UO_1663 (O_1663,N_23760,N_22635);
or UO_1664 (O_1664,N_23384,N_23969);
or UO_1665 (O_1665,N_22387,N_21939);
nor UO_1666 (O_1666,N_23579,N_21926);
nor UO_1667 (O_1667,N_23831,N_23580);
xor UO_1668 (O_1668,N_23623,N_23264);
and UO_1669 (O_1669,N_24136,N_22868);
and UO_1670 (O_1670,N_23936,N_22188);
xor UO_1671 (O_1671,N_22184,N_24315);
or UO_1672 (O_1672,N_23258,N_24031);
xnor UO_1673 (O_1673,N_22054,N_23381);
and UO_1674 (O_1674,N_24707,N_23176);
xnor UO_1675 (O_1675,N_22690,N_23672);
nand UO_1676 (O_1676,N_23976,N_24330);
xnor UO_1677 (O_1677,N_23240,N_23831);
xor UO_1678 (O_1678,N_24678,N_22241);
nor UO_1679 (O_1679,N_24912,N_22801);
nor UO_1680 (O_1680,N_22381,N_24180);
nand UO_1681 (O_1681,N_23360,N_22777);
or UO_1682 (O_1682,N_24208,N_23564);
xor UO_1683 (O_1683,N_24420,N_23385);
and UO_1684 (O_1684,N_23395,N_23366);
nor UO_1685 (O_1685,N_22666,N_24320);
nor UO_1686 (O_1686,N_22445,N_23877);
xor UO_1687 (O_1687,N_24134,N_21994);
nor UO_1688 (O_1688,N_24929,N_23569);
xnor UO_1689 (O_1689,N_24532,N_23449);
nand UO_1690 (O_1690,N_24715,N_23151);
xor UO_1691 (O_1691,N_22843,N_22293);
or UO_1692 (O_1692,N_22543,N_23275);
or UO_1693 (O_1693,N_24826,N_23763);
nand UO_1694 (O_1694,N_22937,N_24072);
and UO_1695 (O_1695,N_22393,N_24416);
nor UO_1696 (O_1696,N_23362,N_24850);
xnor UO_1697 (O_1697,N_22701,N_22503);
and UO_1698 (O_1698,N_24704,N_24966);
nand UO_1699 (O_1699,N_22329,N_23615);
and UO_1700 (O_1700,N_23766,N_23030);
xnor UO_1701 (O_1701,N_21888,N_24517);
or UO_1702 (O_1702,N_24685,N_23248);
or UO_1703 (O_1703,N_23106,N_24936);
or UO_1704 (O_1704,N_24075,N_22597);
xor UO_1705 (O_1705,N_22392,N_24446);
nand UO_1706 (O_1706,N_22285,N_24675);
nor UO_1707 (O_1707,N_23088,N_24980);
nor UO_1708 (O_1708,N_24682,N_24101);
nor UO_1709 (O_1709,N_22959,N_21883);
or UO_1710 (O_1710,N_24048,N_24448);
nor UO_1711 (O_1711,N_24173,N_24038);
or UO_1712 (O_1712,N_22022,N_23950);
xor UO_1713 (O_1713,N_22190,N_23274);
xnor UO_1714 (O_1714,N_24492,N_23315);
xor UO_1715 (O_1715,N_23218,N_22107);
or UO_1716 (O_1716,N_24656,N_22812);
nor UO_1717 (O_1717,N_24449,N_22633);
and UO_1718 (O_1718,N_22832,N_21929);
or UO_1719 (O_1719,N_24017,N_22184);
or UO_1720 (O_1720,N_22400,N_24704);
nand UO_1721 (O_1721,N_24335,N_22883);
nand UO_1722 (O_1722,N_23185,N_23680);
xor UO_1723 (O_1723,N_24890,N_22753);
xor UO_1724 (O_1724,N_22408,N_23921);
nor UO_1725 (O_1725,N_22708,N_22727);
nand UO_1726 (O_1726,N_23839,N_22867);
xnor UO_1727 (O_1727,N_24156,N_23336);
nor UO_1728 (O_1728,N_23811,N_23947);
xnor UO_1729 (O_1729,N_23288,N_22779);
xor UO_1730 (O_1730,N_23479,N_24583);
nand UO_1731 (O_1731,N_24868,N_22426);
and UO_1732 (O_1732,N_22593,N_22985);
or UO_1733 (O_1733,N_22341,N_24995);
or UO_1734 (O_1734,N_24290,N_24275);
nand UO_1735 (O_1735,N_23881,N_22273);
nor UO_1736 (O_1736,N_23074,N_23165);
nand UO_1737 (O_1737,N_24402,N_23406);
nand UO_1738 (O_1738,N_22014,N_23021);
xor UO_1739 (O_1739,N_22819,N_23803);
xor UO_1740 (O_1740,N_23809,N_24668);
nor UO_1741 (O_1741,N_22755,N_24941);
and UO_1742 (O_1742,N_23832,N_22744);
xnor UO_1743 (O_1743,N_23930,N_22589);
or UO_1744 (O_1744,N_23718,N_24899);
nor UO_1745 (O_1745,N_23307,N_23735);
and UO_1746 (O_1746,N_22486,N_23878);
nor UO_1747 (O_1747,N_24900,N_22089);
xor UO_1748 (O_1748,N_24688,N_24137);
and UO_1749 (O_1749,N_23974,N_24811);
nand UO_1750 (O_1750,N_22014,N_24122);
nor UO_1751 (O_1751,N_23838,N_22083);
xor UO_1752 (O_1752,N_24462,N_22295);
xor UO_1753 (O_1753,N_23256,N_22348);
nand UO_1754 (O_1754,N_24377,N_24565);
or UO_1755 (O_1755,N_23507,N_24046);
nand UO_1756 (O_1756,N_24955,N_24917);
and UO_1757 (O_1757,N_22054,N_24212);
and UO_1758 (O_1758,N_23457,N_22261);
nand UO_1759 (O_1759,N_24950,N_23529);
xnor UO_1760 (O_1760,N_24090,N_24516);
and UO_1761 (O_1761,N_24474,N_21972);
or UO_1762 (O_1762,N_23531,N_24203);
and UO_1763 (O_1763,N_22921,N_24605);
and UO_1764 (O_1764,N_23212,N_24869);
or UO_1765 (O_1765,N_24586,N_24527);
nand UO_1766 (O_1766,N_22678,N_23463);
nor UO_1767 (O_1767,N_24986,N_23478);
and UO_1768 (O_1768,N_23820,N_22224);
nand UO_1769 (O_1769,N_23875,N_24776);
and UO_1770 (O_1770,N_23332,N_23496);
or UO_1771 (O_1771,N_21889,N_22059);
and UO_1772 (O_1772,N_21886,N_23892);
xor UO_1773 (O_1773,N_22668,N_22576);
nor UO_1774 (O_1774,N_22381,N_23929);
xnor UO_1775 (O_1775,N_22450,N_23395);
nor UO_1776 (O_1776,N_23554,N_24013);
nand UO_1777 (O_1777,N_22686,N_21918);
nand UO_1778 (O_1778,N_24511,N_23240);
or UO_1779 (O_1779,N_24020,N_23269);
nand UO_1780 (O_1780,N_22644,N_23253);
or UO_1781 (O_1781,N_22695,N_23878);
nor UO_1782 (O_1782,N_24305,N_23080);
and UO_1783 (O_1783,N_24324,N_23289);
nand UO_1784 (O_1784,N_24204,N_21992);
nor UO_1785 (O_1785,N_23678,N_23227);
nand UO_1786 (O_1786,N_24509,N_21911);
nor UO_1787 (O_1787,N_24210,N_21891);
nor UO_1788 (O_1788,N_23424,N_22319);
or UO_1789 (O_1789,N_23391,N_24357);
nand UO_1790 (O_1790,N_24050,N_23275);
nand UO_1791 (O_1791,N_23130,N_22199);
xor UO_1792 (O_1792,N_22846,N_24360);
nor UO_1793 (O_1793,N_21906,N_23172);
nor UO_1794 (O_1794,N_23579,N_24106);
xor UO_1795 (O_1795,N_22469,N_23510);
xnor UO_1796 (O_1796,N_24038,N_24333);
nor UO_1797 (O_1797,N_24903,N_22619);
and UO_1798 (O_1798,N_22922,N_22009);
nor UO_1799 (O_1799,N_22615,N_22910);
xnor UO_1800 (O_1800,N_23816,N_24808);
and UO_1801 (O_1801,N_23200,N_22379);
or UO_1802 (O_1802,N_23344,N_23670);
or UO_1803 (O_1803,N_23470,N_23373);
or UO_1804 (O_1804,N_23707,N_23045);
or UO_1805 (O_1805,N_22748,N_22785);
nand UO_1806 (O_1806,N_24459,N_22104);
or UO_1807 (O_1807,N_22108,N_22651);
and UO_1808 (O_1808,N_24476,N_24485);
or UO_1809 (O_1809,N_24001,N_24275);
nand UO_1810 (O_1810,N_22341,N_24557);
xor UO_1811 (O_1811,N_23188,N_23124);
nand UO_1812 (O_1812,N_22230,N_22481);
and UO_1813 (O_1813,N_22935,N_22459);
and UO_1814 (O_1814,N_23470,N_23068);
nor UO_1815 (O_1815,N_23671,N_23782);
nand UO_1816 (O_1816,N_24248,N_22461);
nand UO_1817 (O_1817,N_24955,N_24744);
nor UO_1818 (O_1818,N_23300,N_24448);
xor UO_1819 (O_1819,N_22963,N_22759);
xor UO_1820 (O_1820,N_22198,N_22159);
or UO_1821 (O_1821,N_22410,N_22241);
or UO_1822 (O_1822,N_23950,N_23655);
or UO_1823 (O_1823,N_22132,N_23793);
nor UO_1824 (O_1824,N_23990,N_22182);
and UO_1825 (O_1825,N_24585,N_23763);
nor UO_1826 (O_1826,N_23193,N_24456);
or UO_1827 (O_1827,N_22189,N_22069);
xnor UO_1828 (O_1828,N_23531,N_23840);
xor UO_1829 (O_1829,N_21975,N_23423);
nor UO_1830 (O_1830,N_24358,N_23744);
or UO_1831 (O_1831,N_22457,N_22427);
nand UO_1832 (O_1832,N_24503,N_24409);
xor UO_1833 (O_1833,N_24325,N_23983);
or UO_1834 (O_1834,N_23205,N_23748);
or UO_1835 (O_1835,N_23846,N_23312);
nor UO_1836 (O_1836,N_24240,N_23377);
nand UO_1837 (O_1837,N_22553,N_24494);
nor UO_1838 (O_1838,N_23295,N_22201);
nor UO_1839 (O_1839,N_22097,N_24501);
xor UO_1840 (O_1840,N_23956,N_23003);
and UO_1841 (O_1841,N_24455,N_22147);
and UO_1842 (O_1842,N_23798,N_24858);
xor UO_1843 (O_1843,N_22176,N_23144);
xnor UO_1844 (O_1844,N_23885,N_22204);
nand UO_1845 (O_1845,N_22953,N_22441);
or UO_1846 (O_1846,N_22631,N_23435);
xnor UO_1847 (O_1847,N_24338,N_22796);
nor UO_1848 (O_1848,N_24477,N_24867);
nand UO_1849 (O_1849,N_23635,N_23538);
xnor UO_1850 (O_1850,N_23437,N_23538);
and UO_1851 (O_1851,N_24008,N_22543);
nand UO_1852 (O_1852,N_22244,N_24629);
nand UO_1853 (O_1853,N_24438,N_23357);
nor UO_1854 (O_1854,N_21903,N_22345);
and UO_1855 (O_1855,N_23749,N_22221);
xor UO_1856 (O_1856,N_24602,N_23609);
xor UO_1857 (O_1857,N_23226,N_24547);
xnor UO_1858 (O_1858,N_23723,N_22779);
nand UO_1859 (O_1859,N_24308,N_24890);
and UO_1860 (O_1860,N_24412,N_23113);
or UO_1861 (O_1861,N_24215,N_22361);
or UO_1862 (O_1862,N_24029,N_24633);
nor UO_1863 (O_1863,N_22709,N_23493);
nor UO_1864 (O_1864,N_24774,N_22857);
and UO_1865 (O_1865,N_22471,N_24512);
nor UO_1866 (O_1866,N_24585,N_22054);
and UO_1867 (O_1867,N_22379,N_24891);
nor UO_1868 (O_1868,N_23262,N_23773);
and UO_1869 (O_1869,N_22973,N_23981);
and UO_1870 (O_1870,N_22681,N_22168);
nand UO_1871 (O_1871,N_23839,N_22230);
xnor UO_1872 (O_1872,N_22487,N_22168);
and UO_1873 (O_1873,N_22946,N_22521);
nor UO_1874 (O_1874,N_22088,N_21921);
nor UO_1875 (O_1875,N_24125,N_22489);
xnor UO_1876 (O_1876,N_22883,N_24389);
nor UO_1877 (O_1877,N_22610,N_24723);
nor UO_1878 (O_1878,N_24120,N_24687);
or UO_1879 (O_1879,N_22490,N_23231);
xnor UO_1880 (O_1880,N_22605,N_24093);
nor UO_1881 (O_1881,N_23806,N_24260);
or UO_1882 (O_1882,N_24795,N_22749);
nand UO_1883 (O_1883,N_22370,N_21908);
nor UO_1884 (O_1884,N_24165,N_22911);
or UO_1885 (O_1885,N_22396,N_23166);
and UO_1886 (O_1886,N_23784,N_24771);
nand UO_1887 (O_1887,N_24635,N_21888);
nand UO_1888 (O_1888,N_24622,N_23800);
nand UO_1889 (O_1889,N_24023,N_21953);
or UO_1890 (O_1890,N_22812,N_23581);
xnor UO_1891 (O_1891,N_23093,N_22993);
nand UO_1892 (O_1892,N_22972,N_24328);
nand UO_1893 (O_1893,N_24676,N_22048);
nand UO_1894 (O_1894,N_24844,N_21946);
nand UO_1895 (O_1895,N_23286,N_22410);
nor UO_1896 (O_1896,N_23714,N_22847);
or UO_1897 (O_1897,N_24044,N_24697);
nand UO_1898 (O_1898,N_22821,N_22968);
nor UO_1899 (O_1899,N_23024,N_22818);
or UO_1900 (O_1900,N_22783,N_24961);
nand UO_1901 (O_1901,N_24598,N_22252);
xnor UO_1902 (O_1902,N_24471,N_23929);
and UO_1903 (O_1903,N_24403,N_23765);
or UO_1904 (O_1904,N_24561,N_22619);
nand UO_1905 (O_1905,N_23964,N_24119);
and UO_1906 (O_1906,N_22085,N_23178);
xor UO_1907 (O_1907,N_22632,N_24516);
nor UO_1908 (O_1908,N_22665,N_22363);
nor UO_1909 (O_1909,N_24708,N_24360);
xor UO_1910 (O_1910,N_22640,N_24654);
and UO_1911 (O_1911,N_22318,N_24204);
nor UO_1912 (O_1912,N_23667,N_24266);
nand UO_1913 (O_1913,N_24931,N_23939);
and UO_1914 (O_1914,N_23857,N_22437);
nand UO_1915 (O_1915,N_24680,N_22981);
xor UO_1916 (O_1916,N_24045,N_24951);
xor UO_1917 (O_1917,N_24626,N_23364);
xor UO_1918 (O_1918,N_21921,N_23597);
xnor UO_1919 (O_1919,N_24700,N_23854);
and UO_1920 (O_1920,N_24520,N_24852);
nand UO_1921 (O_1921,N_24065,N_24901);
xor UO_1922 (O_1922,N_24176,N_23740);
and UO_1923 (O_1923,N_23023,N_23858);
nand UO_1924 (O_1924,N_22011,N_23055);
xnor UO_1925 (O_1925,N_23856,N_23296);
or UO_1926 (O_1926,N_21932,N_24036);
nand UO_1927 (O_1927,N_24964,N_23784);
and UO_1928 (O_1928,N_22048,N_22813);
and UO_1929 (O_1929,N_22559,N_24798);
and UO_1930 (O_1930,N_22692,N_22606);
and UO_1931 (O_1931,N_24574,N_22972);
or UO_1932 (O_1932,N_23605,N_22090);
and UO_1933 (O_1933,N_22677,N_24824);
and UO_1934 (O_1934,N_22694,N_24382);
nand UO_1935 (O_1935,N_24879,N_24226);
nand UO_1936 (O_1936,N_23084,N_23232);
xnor UO_1937 (O_1937,N_22261,N_22848);
and UO_1938 (O_1938,N_23893,N_24546);
nor UO_1939 (O_1939,N_22766,N_23537);
nor UO_1940 (O_1940,N_22183,N_22381);
or UO_1941 (O_1941,N_23690,N_23086);
nand UO_1942 (O_1942,N_23933,N_23143);
nand UO_1943 (O_1943,N_24355,N_22181);
nand UO_1944 (O_1944,N_24393,N_24024);
nand UO_1945 (O_1945,N_24267,N_24007);
xor UO_1946 (O_1946,N_24436,N_22243);
or UO_1947 (O_1947,N_23509,N_23421);
nor UO_1948 (O_1948,N_24607,N_24931);
xor UO_1949 (O_1949,N_24701,N_22016);
xor UO_1950 (O_1950,N_22633,N_22200);
xnor UO_1951 (O_1951,N_24899,N_24917);
or UO_1952 (O_1952,N_23107,N_23101);
nand UO_1953 (O_1953,N_23875,N_22565);
xor UO_1954 (O_1954,N_23596,N_23675);
xnor UO_1955 (O_1955,N_24793,N_23352);
nor UO_1956 (O_1956,N_22705,N_22980);
nand UO_1957 (O_1957,N_21894,N_22773);
nor UO_1958 (O_1958,N_22594,N_23726);
or UO_1959 (O_1959,N_22588,N_21888);
xor UO_1960 (O_1960,N_24040,N_24668);
nand UO_1961 (O_1961,N_23187,N_24727);
and UO_1962 (O_1962,N_21942,N_23883);
and UO_1963 (O_1963,N_24271,N_22796);
nor UO_1964 (O_1964,N_24121,N_24802);
xnor UO_1965 (O_1965,N_23971,N_22761);
or UO_1966 (O_1966,N_22012,N_22935);
nand UO_1967 (O_1967,N_24849,N_24980);
or UO_1968 (O_1968,N_24884,N_23149);
xor UO_1969 (O_1969,N_23482,N_22863);
or UO_1970 (O_1970,N_22395,N_24305);
or UO_1971 (O_1971,N_24292,N_24372);
nor UO_1972 (O_1972,N_23634,N_24330);
nand UO_1973 (O_1973,N_22735,N_22007);
xor UO_1974 (O_1974,N_24592,N_23762);
and UO_1975 (O_1975,N_22033,N_22094);
and UO_1976 (O_1976,N_24049,N_24138);
xor UO_1977 (O_1977,N_22773,N_24434);
xor UO_1978 (O_1978,N_24587,N_22151);
nand UO_1979 (O_1979,N_23760,N_22695);
nor UO_1980 (O_1980,N_23286,N_24536);
nor UO_1981 (O_1981,N_24525,N_21908);
or UO_1982 (O_1982,N_24436,N_22409);
or UO_1983 (O_1983,N_24053,N_22522);
xnor UO_1984 (O_1984,N_24505,N_24592);
or UO_1985 (O_1985,N_24296,N_21963);
or UO_1986 (O_1986,N_21959,N_22962);
nand UO_1987 (O_1987,N_23199,N_23765);
xnor UO_1988 (O_1988,N_23111,N_24988);
nand UO_1989 (O_1989,N_23741,N_23676);
nor UO_1990 (O_1990,N_22194,N_24912);
or UO_1991 (O_1991,N_23134,N_22187);
or UO_1992 (O_1992,N_24124,N_24174);
nor UO_1993 (O_1993,N_24101,N_21950);
nor UO_1994 (O_1994,N_22859,N_23937);
or UO_1995 (O_1995,N_22024,N_23748);
and UO_1996 (O_1996,N_22040,N_22011);
nor UO_1997 (O_1997,N_22384,N_24208);
or UO_1998 (O_1998,N_23217,N_23004);
xor UO_1999 (O_1999,N_24010,N_21889);
or UO_2000 (O_2000,N_23367,N_23053);
nor UO_2001 (O_2001,N_23684,N_23836);
and UO_2002 (O_2002,N_24967,N_22467);
or UO_2003 (O_2003,N_23013,N_24766);
or UO_2004 (O_2004,N_21899,N_22973);
and UO_2005 (O_2005,N_24139,N_22739);
xor UO_2006 (O_2006,N_24146,N_24720);
nor UO_2007 (O_2007,N_24851,N_22206);
and UO_2008 (O_2008,N_22420,N_24987);
nand UO_2009 (O_2009,N_24524,N_23162);
xor UO_2010 (O_2010,N_22341,N_22551);
nor UO_2011 (O_2011,N_22414,N_22751);
nor UO_2012 (O_2012,N_24199,N_23525);
or UO_2013 (O_2013,N_21928,N_24228);
and UO_2014 (O_2014,N_22399,N_22277);
xnor UO_2015 (O_2015,N_24063,N_22211);
or UO_2016 (O_2016,N_23997,N_22846);
nand UO_2017 (O_2017,N_22181,N_22167);
xor UO_2018 (O_2018,N_22043,N_23238);
nor UO_2019 (O_2019,N_24861,N_23274);
nor UO_2020 (O_2020,N_24647,N_24577);
xor UO_2021 (O_2021,N_24988,N_24198);
nand UO_2022 (O_2022,N_22371,N_22792);
or UO_2023 (O_2023,N_24715,N_23977);
nor UO_2024 (O_2024,N_22775,N_24402);
nand UO_2025 (O_2025,N_22176,N_24430);
or UO_2026 (O_2026,N_24562,N_24838);
and UO_2027 (O_2027,N_23180,N_23138);
nor UO_2028 (O_2028,N_21995,N_23302);
xor UO_2029 (O_2029,N_23308,N_23999);
nand UO_2030 (O_2030,N_24459,N_24109);
xor UO_2031 (O_2031,N_23617,N_24090);
xor UO_2032 (O_2032,N_22123,N_23816);
nor UO_2033 (O_2033,N_21957,N_24143);
nor UO_2034 (O_2034,N_24306,N_24504);
or UO_2035 (O_2035,N_24424,N_24586);
xnor UO_2036 (O_2036,N_24759,N_23443);
xor UO_2037 (O_2037,N_24692,N_22407);
and UO_2038 (O_2038,N_23011,N_22203);
nor UO_2039 (O_2039,N_22063,N_24344);
nand UO_2040 (O_2040,N_23872,N_23480);
and UO_2041 (O_2041,N_23767,N_23574);
xnor UO_2042 (O_2042,N_23741,N_24352);
xor UO_2043 (O_2043,N_24592,N_22512);
and UO_2044 (O_2044,N_22916,N_22303);
xor UO_2045 (O_2045,N_23748,N_23704);
or UO_2046 (O_2046,N_22523,N_23738);
nor UO_2047 (O_2047,N_24626,N_24518);
or UO_2048 (O_2048,N_22310,N_22300);
nand UO_2049 (O_2049,N_24482,N_22609);
nand UO_2050 (O_2050,N_22240,N_22154);
and UO_2051 (O_2051,N_23571,N_22579);
or UO_2052 (O_2052,N_22705,N_24718);
nand UO_2053 (O_2053,N_22765,N_22032);
xnor UO_2054 (O_2054,N_21944,N_24984);
or UO_2055 (O_2055,N_24412,N_23645);
and UO_2056 (O_2056,N_22820,N_24453);
or UO_2057 (O_2057,N_22048,N_24441);
or UO_2058 (O_2058,N_24679,N_22463);
or UO_2059 (O_2059,N_24469,N_22384);
or UO_2060 (O_2060,N_22742,N_23411);
nand UO_2061 (O_2061,N_23297,N_24821);
nand UO_2062 (O_2062,N_22254,N_23610);
nand UO_2063 (O_2063,N_23939,N_21953);
nor UO_2064 (O_2064,N_23153,N_24783);
or UO_2065 (O_2065,N_22866,N_24843);
and UO_2066 (O_2066,N_22425,N_24608);
xor UO_2067 (O_2067,N_23026,N_24730);
xor UO_2068 (O_2068,N_24720,N_22400);
nand UO_2069 (O_2069,N_22612,N_22059);
or UO_2070 (O_2070,N_23965,N_24497);
and UO_2071 (O_2071,N_24515,N_24643);
and UO_2072 (O_2072,N_24815,N_22845);
and UO_2073 (O_2073,N_24906,N_22931);
nand UO_2074 (O_2074,N_21983,N_22333);
and UO_2075 (O_2075,N_24194,N_24840);
nor UO_2076 (O_2076,N_23296,N_22132);
or UO_2077 (O_2077,N_22676,N_22409);
and UO_2078 (O_2078,N_23640,N_24689);
nor UO_2079 (O_2079,N_22161,N_23598);
and UO_2080 (O_2080,N_22982,N_24165);
or UO_2081 (O_2081,N_24141,N_23848);
or UO_2082 (O_2082,N_23834,N_23591);
nand UO_2083 (O_2083,N_23972,N_22844);
or UO_2084 (O_2084,N_24086,N_23672);
nand UO_2085 (O_2085,N_22992,N_23190);
nor UO_2086 (O_2086,N_21975,N_23594);
and UO_2087 (O_2087,N_24090,N_21958);
and UO_2088 (O_2088,N_24078,N_22393);
nand UO_2089 (O_2089,N_23086,N_23660);
and UO_2090 (O_2090,N_24261,N_23852);
or UO_2091 (O_2091,N_22748,N_22532);
nand UO_2092 (O_2092,N_24931,N_23963);
nor UO_2093 (O_2093,N_23040,N_24776);
or UO_2094 (O_2094,N_23678,N_23688);
xor UO_2095 (O_2095,N_23154,N_22497);
nor UO_2096 (O_2096,N_22593,N_22837);
and UO_2097 (O_2097,N_23799,N_22819);
and UO_2098 (O_2098,N_23160,N_22828);
xor UO_2099 (O_2099,N_24671,N_23044);
or UO_2100 (O_2100,N_22988,N_23927);
or UO_2101 (O_2101,N_24430,N_23841);
nor UO_2102 (O_2102,N_23064,N_23765);
nand UO_2103 (O_2103,N_22206,N_22341);
xnor UO_2104 (O_2104,N_22390,N_23820);
or UO_2105 (O_2105,N_22976,N_21977);
nand UO_2106 (O_2106,N_22863,N_22469);
nor UO_2107 (O_2107,N_24359,N_23973);
and UO_2108 (O_2108,N_24778,N_23983);
nand UO_2109 (O_2109,N_22601,N_24418);
xor UO_2110 (O_2110,N_23885,N_24734);
and UO_2111 (O_2111,N_23942,N_24237);
nand UO_2112 (O_2112,N_22839,N_23008);
xor UO_2113 (O_2113,N_24239,N_22690);
xnor UO_2114 (O_2114,N_24614,N_22034);
and UO_2115 (O_2115,N_24158,N_23624);
xor UO_2116 (O_2116,N_24921,N_22262);
nor UO_2117 (O_2117,N_24650,N_23373);
or UO_2118 (O_2118,N_23729,N_24432);
nor UO_2119 (O_2119,N_22860,N_22901);
nand UO_2120 (O_2120,N_24899,N_22542);
and UO_2121 (O_2121,N_23735,N_22329);
or UO_2122 (O_2122,N_22058,N_23106);
and UO_2123 (O_2123,N_22617,N_24091);
and UO_2124 (O_2124,N_23761,N_24269);
nor UO_2125 (O_2125,N_24359,N_24000);
xnor UO_2126 (O_2126,N_23142,N_23768);
or UO_2127 (O_2127,N_22654,N_22732);
and UO_2128 (O_2128,N_24869,N_22267);
nand UO_2129 (O_2129,N_23540,N_23680);
or UO_2130 (O_2130,N_23863,N_23049);
and UO_2131 (O_2131,N_24301,N_23025);
nor UO_2132 (O_2132,N_24365,N_24786);
nor UO_2133 (O_2133,N_23097,N_22363);
or UO_2134 (O_2134,N_22677,N_24474);
or UO_2135 (O_2135,N_24058,N_24045);
nor UO_2136 (O_2136,N_23378,N_24759);
and UO_2137 (O_2137,N_22525,N_24409);
nor UO_2138 (O_2138,N_24056,N_24157);
nand UO_2139 (O_2139,N_24145,N_23205);
or UO_2140 (O_2140,N_24638,N_24072);
and UO_2141 (O_2141,N_24964,N_23502);
nor UO_2142 (O_2142,N_23452,N_24672);
nor UO_2143 (O_2143,N_24658,N_24339);
nor UO_2144 (O_2144,N_22685,N_23339);
or UO_2145 (O_2145,N_23148,N_22316);
or UO_2146 (O_2146,N_24994,N_24141);
and UO_2147 (O_2147,N_23091,N_24351);
xnor UO_2148 (O_2148,N_24871,N_23238);
and UO_2149 (O_2149,N_21985,N_24933);
nor UO_2150 (O_2150,N_24413,N_22026);
xor UO_2151 (O_2151,N_24102,N_22724);
and UO_2152 (O_2152,N_22564,N_22543);
nand UO_2153 (O_2153,N_23658,N_22645);
or UO_2154 (O_2154,N_24597,N_23739);
nor UO_2155 (O_2155,N_22058,N_24161);
and UO_2156 (O_2156,N_24211,N_24688);
xor UO_2157 (O_2157,N_24883,N_23104);
and UO_2158 (O_2158,N_22322,N_22406);
and UO_2159 (O_2159,N_22977,N_23777);
and UO_2160 (O_2160,N_23101,N_24978);
xnor UO_2161 (O_2161,N_22781,N_22886);
or UO_2162 (O_2162,N_24821,N_24092);
and UO_2163 (O_2163,N_24030,N_23914);
xor UO_2164 (O_2164,N_22601,N_22203);
xor UO_2165 (O_2165,N_22555,N_23412);
or UO_2166 (O_2166,N_22187,N_24050);
xor UO_2167 (O_2167,N_22457,N_22006);
and UO_2168 (O_2168,N_23002,N_24256);
nor UO_2169 (O_2169,N_22980,N_24843);
nor UO_2170 (O_2170,N_24041,N_22054);
xnor UO_2171 (O_2171,N_22903,N_23412);
and UO_2172 (O_2172,N_23315,N_24371);
xor UO_2173 (O_2173,N_23201,N_22452);
nand UO_2174 (O_2174,N_24296,N_23401);
nor UO_2175 (O_2175,N_23267,N_22689);
nand UO_2176 (O_2176,N_24196,N_22318);
nor UO_2177 (O_2177,N_24322,N_22649);
or UO_2178 (O_2178,N_22091,N_24543);
or UO_2179 (O_2179,N_23345,N_23976);
nor UO_2180 (O_2180,N_24017,N_21978);
and UO_2181 (O_2181,N_22125,N_22920);
and UO_2182 (O_2182,N_24808,N_23370);
or UO_2183 (O_2183,N_24412,N_22852);
and UO_2184 (O_2184,N_22190,N_22099);
and UO_2185 (O_2185,N_22349,N_22193);
or UO_2186 (O_2186,N_24458,N_24956);
nand UO_2187 (O_2187,N_23382,N_22250);
or UO_2188 (O_2188,N_21993,N_22636);
nand UO_2189 (O_2189,N_23681,N_22218);
nand UO_2190 (O_2190,N_24482,N_24939);
nor UO_2191 (O_2191,N_22205,N_24769);
or UO_2192 (O_2192,N_23682,N_24316);
or UO_2193 (O_2193,N_24859,N_24124);
nor UO_2194 (O_2194,N_22706,N_22466);
and UO_2195 (O_2195,N_23783,N_23644);
nand UO_2196 (O_2196,N_23087,N_24601);
nor UO_2197 (O_2197,N_22448,N_24377);
nor UO_2198 (O_2198,N_22193,N_24567);
xnor UO_2199 (O_2199,N_22052,N_21880);
and UO_2200 (O_2200,N_23851,N_24495);
nor UO_2201 (O_2201,N_22914,N_23431);
and UO_2202 (O_2202,N_23192,N_22593);
nor UO_2203 (O_2203,N_23886,N_23938);
or UO_2204 (O_2204,N_22942,N_22961);
or UO_2205 (O_2205,N_22499,N_23493);
or UO_2206 (O_2206,N_24034,N_23272);
nand UO_2207 (O_2207,N_23120,N_24835);
nand UO_2208 (O_2208,N_22158,N_24585);
xnor UO_2209 (O_2209,N_23476,N_22314);
xnor UO_2210 (O_2210,N_22308,N_22480);
nand UO_2211 (O_2211,N_24489,N_22954);
and UO_2212 (O_2212,N_24914,N_24848);
or UO_2213 (O_2213,N_22091,N_23739);
nand UO_2214 (O_2214,N_22588,N_22152);
xor UO_2215 (O_2215,N_22659,N_23738);
and UO_2216 (O_2216,N_21997,N_24593);
or UO_2217 (O_2217,N_24266,N_24602);
and UO_2218 (O_2218,N_22247,N_22420);
and UO_2219 (O_2219,N_21881,N_24211);
nor UO_2220 (O_2220,N_24381,N_23276);
or UO_2221 (O_2221,N_22577,N_24672);
nand UO_2222 (O_2222,N_23733,N_24533);
nor UO_2223 (O_2223,N_24456,N_24384);
nand UO_2224 (O_2224,N_24080,N_22732);
or UO_2225 (O_2225,N_22842,N_23089);
xnor UO_2226 (O_2226,N_24821,N_23921);
nor UO_2227 (O_2227,N_22707,N_22514);
and UO_2228 (O_2228,N_22273,N_24335);
or UO_2229 (O_2229,N_23116,N_23760);
and UO_2230 (O_2230,N_24399,N_23501);
nand UO_2231 (O_2231,N_24870,N_24766);
nor UO_2232 (O_2232,N_21877,N_23656);
nand UO_2233 (O_2233,N_23165,N_24136);
nand UO_2234 (O_2234,N_23186,N_23914);
or UO_2235 (O_2235,N_24222,N_23409);
nor UO_2236 (O_2236,N_24663,N_22985);
nor UO_2237 (O_2237,N_23187,N_24442);
xnor UO_2238 (O_2238,N_24101,N_22784);
or UO_2239 (O_2239,N_23095,N_23655);
or UO_2240 (O_2240,N_23505,N_23792);
nand UO_2241 (O_2241,N_23347,N_24770);
xor UO_2242 (O_2242,N_23356,N_24656);
or UO_2243 (O_2243,N_22243,N_22190);
nor UO_2244 (O_2244,N_24157,N_24710);
xor UO_2245 (O_2245,N_24683,N_22346);
or UO_2246 (O_2246,N_23874,N_23607);
xor UO_2247 (O_2247,N_23355,N_22747);
nor UO_2248 (O_2248,N_23212,N_22110);
or UO_2249 (O_2249,N_23938,N_23781);
nand UO_2250 (O_2250,N_23481,N_24562);
xnor UO_2251 (O_2251,N_22912,N_23235);
xnor UO_2252 (O_2252,N_24380,N_23523);
and UO_2253 (O_2253,N_23624,N_23024);
or UO_2254 (O_2254,N_24530,N_23474);
and UO_2255 (O_2255,N_24658,N_21970);
or UO_2256 (O_2256,N_22295,N_24896);
and UO_2257 (O_2257,N_22831,N_23048);
xnor UO_2258 (O_2258,N_23983,N_22616);
xor UO_2259 (O_2259,N_22278,N_23934);
nand UO_2260 (O_2260,N_22959,N_22568);
and UO_2261 (O_2261,N_22632,N_23247);
xnor UO_2262 (O_2262,N_23279,N_22332);
and UO_2263 (O_2263,N_22109,N_23287);
and UO_2264 (O_2264,N_23660,N_22259);
and UO_2265 (O_2265,N_23303,N_24731);
nor UO_2266 (O_2266,N_22830,N_22001);
xor UO_2267 (O_2267,N_24332,N_22012);
or UO_2268 (O_2268,N_24656,N_22945);
and UO_2269 (O_2269,N_22265,N_23135);
xnor UO_2270 (O_2270,N_24511,N_23569);
or UO_2271 (O_2271,N_23418,N_23529);
xnor UO_2272 (O_2272,N_24808,N_23959);
xnor UO_2273 (O_2273,N_22887,N_23748);
nor UO_2274 (O_2274,N_24674,N_24928);
nand UO_2275 (O_2275,N_22800,N_24823);
xnor UO_2276 (O_2276,N_24319,N_24988);
nand UO_2277 (O_2277,N_24328,N_23530);
nor UO_2278 (O_2278,N_23039,N_24207);
or UO_2279 (O_2279,N_24335,N_22863);
and UO_2280 (O_2280,N_24201,N_22010);
or UO_2281 (O_2281,N_24010,N_22332);
nor UO_2282 (O_2282,N_23597,N_24746);
and UO_2283 (O_2283,N_23287,N_23684);
or UO_2284 (O_2284,N_24123,N_24250);
or UO_2285 (O_2285,N_21967,N_24162);
and UO_2286 (O_2286,N_24394,N_22727);
nor UO_2287 (O_2287,N_22129,N_23350);
nor UO_2288 (O_2288,N_22831,N_22699);
nor UO_2289 (O_2289,N_24883,N_22057);
and UO_2290 (O_2290,N_23478,N_23581);
nand UO_2291 (O_2291,N_22410,N_23292);
nor UO_2292 (O_2292,N_21879,N_22141);
or UO_2293 (O_2293,N_22514,N_22036);
or UO_2294 (O_2294,N_21955,N_23384);
xor UO_2295 (O_2295,N_21945,N_23048);
nor UO_2296 (O_2296,N_24672,N_24455);
and UO_2297 (O_2297,N_22118,N_23169);
xnor UO_2298 (O_2298,N_22626,N_23430);
xor UO_2299 (O_2299,N_22794,N_22989);
nand UO_2300 (O_2300,N_22497,N_24306);
or UO_2301 (O_2301,N_23905,N_24059);
nand UO_2302 (O_2302,N_23239,N_22734);
nor UO_2303 (O_2303,N_24796,N_23068);
xnor UO_2304 (O_2304,N_23917,N_24394);
nand UO_2305 (O_2305,N_22111,N_22837);
or UO_2306 (O_2306,N_24266,N_23823);
or UO_2307 (O_2307,N_24521,N_21977);
and UO_2308 (O_2308,N_24747,N_21996);
or UO_2309 (O_2309,N_24187,N_24495);
nor UO_2310 (O_2310,N_23820,N_22675);
nand UO_2311 (O_2311,N_23509,N_22991);
or UO_2312 (O_2312,N_22080,N_22647);
and UO_2313 (O_2313,N_22057,N_22956);
xor UO_2314 (O_2314,N_23269,N_23471);
and UO_2315 (O_2315,N_23928,N_22389);
nand UO_2316 (O_2316,N_23751,N_24941);
nor UO_2317 (O_2317,N_22284,N_22932);
xor UO_2318 (O_2318,N_21967,N_24243);
nor UO_2319 (O_2319,N_23573,N_21922);
or UO_2320 (O_2320,N_24999,N_21930);
xnor UO_2321 (O_2321,N_23916,N_23117);
nand UO_2322 (O_2322,N_24189,N_22873);
nor UO_2323 (O_2323,N_21961,N_23250);
nor UO_2324 (O_2324,N_23507,N_22972);
or UO_2325 (O_2325,N_23347,N_24714);
nor UO_2326 (O_2326,N_23059,N_22808);
or UO_2327 (O_2327,N_22547,N_24385);
xnor UO_2328 (O_2328,N_22683,N_23682);
xnor UO_2329 (O_2329,N_22552,N_23444);
nand UO_2330 (O_2330,N_22826,N_23022);
nand UO_2331 (O_2331,N_22676,N_22224);
xnor UO_2332 (O_2332,N_23726,N_24639);
nor UO_2333 (O_2333,N_23260,N_22503);
nor UO_2334 (O_2334,N_23875,N_22367);
nand UO_2335 (O_2335,N_23321,N_23582);
or UO_2336 (O_2336,N_22451,N_22549);
or UO_2337 (O_2337,N_23706,N_23119);
and UO_2338 (O_2338,N_24087,N_24382);
or UO_2339 (O_2339,N_22475,N_24201);
xor UO_2340 (O_2340,N_24772,N_23105);
and UO_2341 (O_2341,N_23970,N_23456);
nand UO_2342 (O_2342,N_23482,N_24209);
nand UO_2343 (O_2343,N_23341,N_24575);
or UO_2344 (O_2344,N_22160,N_24525);
xor UO_2345 (O_2345,N_22928,N_23385);
and UO_2346 (O_2346,N_22676,N_23439);
nand UO_2347 (O_2347,N_23613,N_23392);
or UO_2348 (O_2348,N_22800,N_23561);
or UO_2349 (O_2349,N_24994,N_22440);
nor UO_2350 (O_2350,N_24702,N_22829);
xnor UO_2351 (O_2351,N_23555,N_22048);
nand UO_2352 (O_2352,N_22579,N_22384);
and UO_2353 (O_2353,N_22228,N_23060);
and UO_2354 (O_2354,N_23024,N_24027);
or UO_2355 (O_2355,N_24292,N_22760);
or UO_2356 (O_2356,N_23209,N_22614);
and UO_2357 (O_2357,N_24793,N_22807);
and UO_2358 (O_2358,N_23961,N_23578);
or UO_2359 (O_2359,N_23990,N_24730);
and UO_2360 (O_2360,N_23356,N_22895);
nor UO_2361 (O_2361,N_22316,N_23368);
or UO_2362 (O_2362,N_22705,N_24549);
xor UO_2363 (O_2363,N_24715,N_22321);
xor UO_2364 (O_2364,N_24595,N_22493);
nor UO_2365 (O_2365,N_23670,N_21933);
or UO_2366 (O_2366,N_22196,N_22400);
nor UO_2367 (O_2367,N_22527,N_24055);
nor UO_2368 (O_2368,N_23002,N_24746);
and UO_2369 (O_2369,N_22501,N_23261);
or UO_2370 (O_2370,N_24634,N_22408);
or UO_2371 (O_2371,N_23859,N_24994);
nor UO_2372 (O_2372,N_22124,N_22025);
xnor UO_2373 (O_2373,N_24831,N_24731);
or UO_2374 (O_2374,N_24036,N_22813);
xor UO_2375 (O_2375,N_22867,N_23263);
nor UO_2376 (O_2376,N_22581,N_22124);
and UO_2377 (O_2377,N_24239,N_22472);
nor UO_2378 (O_2378,N_23083,N_22907);
nand UO_2379 (O_2379,N_22833,N_22707);
or UO_2380 (O_2380,N_23304,N_21966);
xor UO_2381 (O_2381,N_22050,N_24759);
and UO_2382 (O_2382,N_23304,N_22610);
and UO_2383 (O_2383,N_22148,N_22284);
nand UO_2384 (O_2384,N_22269,N_23284);
xor UO_2385 (O_2385,N_22688,N_23133);
xor UO_2386 (O_2386,N_22771,N_22735);
xnor UO_2387 (O_2387,N_24133,N_23459);
nand UO_2388 (O_2388,N_24251,N_24853);
and UO_2389 (O_2389,N_24850,N_22747);
nor UO_2390 (O_2390,N_24503,N_23863);
nor UO_2391 (O_2391,N_24438,N_23941);
nor UO_2392 (O_2392,N_22344,N_24410);
nor UO_2393 (O_2393,N_21925,N_23749);
and UO_2394 (O_2394,N_22052,N_23086);
nor UO_2395 (O_2395,N_22873,N_22765);
and UO_2396 (O_2396,N_22842,N_22337);
nor UO_2397 (O_2397,N_23380,N_22519);
nor UO_2398 (O_2398,N_22892,N_22442);
nor UO_2399 (O_2399,N_24694,N_23907);
xor UO_2400 (O_2400,N_24579,N_24291);
nand UO_2401 (O_2401,N_24689,N_23998);
nor UO_2402 (O_2402,N_22141,N_23830);
or UO_2403 (O_2403,N_24881,N_22187);
xnor UO_2404 (O_2404,N_23632,N_22848);
and UO_2405 (O_2405,N_24479,N_24543);
xnor UO_2406 (O_2406,N_23932,N_23427);
nor UO_2407 (O_2407,N_22873,N_24232);
nand UO_2408 (O_2408,N_22570,N_22578);
xor UO_2409 (O_2409,N_22769,N_24803);
xnor UO_2410 (O_2410,N_21913,N_24170);
and UO_2411 (O_2411,N_22244,N_23563);
and UO_2412 (O_2412,N_24513,N_23792);
nand UO_2413 (O_2413,N_24058,N_24286);
or UO_2414 (O_2414,N_24339,N_22865);
or UO_2415 (O_2415,N_24964,N_23664);
and UO_2416 (O_2416,N_23677,N_23297);
nor UO_2417 (O_2417,N_22220,N_23366);
and UO_2418 (O_2418,N_24277,N_21888);
nand UO_2419 (O_2419,N_22989,N_22074);
or UO_2420 (O_2420,N_22454,N_22849);
nand UO_2421 (O_2421,N_24606,N_24364);
nand UO_2422 (O_2422,N_21883,N_21981);
nand UO_2423 (O_2423,N_24616,N_23860);
or UO_2424 (O_2424,N_22569,N_23380);
and UO_2425 (O_2425,N_22510,N_24878);
xor UO_2426 (O_2426,N_23570,N_24424);
nand UO_2427 (O_2427,N_22403,N_22904);
or UO_2428 (O_2428,N_22360,N_22379);
or UO_2429 (O_2429,N_24995,N_22708);
nor UO_2430 (O_2430,N_22906,N_23258);
nand UO_2431 (O_2431,N_22415,N_24318);
or UO_2432 (O_2432,N_24116,N_24226);
nor UO_2433 (O_2433,N_24485,N_22079);
nand UO_2434 (O_2434,N_23989,N_22691);
xnor UO_2435 (O_2435,N_24179,N_22852);
or UO_2436 (O_2436,N_23986,N_24677);
nor UO_2437 (O_2437,N_23198,N_23767);
nor UO_2438 (O_2438,N_22806,N_23490);
nand UO_2439 (O_2439,N_22332,N_24730);
nand UO_2440 (O_2440,N_22586,N_22211);
nand UO_2441 (O_2441,N_24165,N_23220);
and UO_2442 (O_2442,N_24576,N_23577);
or UO_2443 (O_2443,N_24516,N_24660);
and UO_2444 (O_2444,N_23405,N_24512);
xor UO_2445 (O_2445,N_22106,N_22746);
xnor UO_2446 (O_2446,N_23315,N_23193);
xnor UO_2447 (O_2447,N_24380,N_22018);
or UO_2448 (O_2448,N_22789,N_22498);
xnor UO_2449 (O_2449,N_24179,N_23623);
nor UO_2450 (O_2450,N_24034,N_22486);
and UO_2451 (O_2451,N_22870,N_24165);
or UO_2452 (O_2452,N_23308,N_22904);
and UO_2453 (O_2453,N_22196,N_24511);
or UO_2454 (O_2454,N_22224,N_24370);
and UO_2455 (O_2455,N_22262,N_22293);
or UO_2456 (O_2456,N_24035,N_24756);
nand UO_2457 (O_2457,N_23032,N_23712);
nand UO_2458 (O_2458,N_23261,N_22254);
and UO_2459 (O_2459,N_24049,N_22643);
nor UO_2460 (O_2460,N_22553,N_24068);
and UO_2461 (O_2461,N_23381,N_24171);
and UO_2462 (O_2462,N_24732,N_23067);
and UO_2463 (O_2463,N_23308,N_22032);
or UO_2464 (O_2464,N_24087,N_23762);
nor UO_2465 (O_2465,N_23541,N_24988);
and UO_2466 (O_2466,N_24626,N_22079);
xnor UO_2467 (O_2467,N_23431,N_22391);
nor UO_2468 (O_2468,N_22089,N_24801);
or UO_2469 (O_2469,N_22974,N_21941);
nor UO_2470 (O_2470,N_23268,N_24644);
or UO_2471 (O_2471,N_23139,N_23785);
xnor UO_2472 (O_2472,N_24843,N_22259);
and UO_2473 (O_2473,N_22062,N_22076);
or UO_2474 (O_2474,N_24116,N_24566);
or UO_2475 (O_2475,N_23435,N_22141);
and UO_2476 (O_2476,N_24611,N_24237);
nor UO_2477 (O_2477,N_24691,N_24508);
xnor UO_2478 (O_2478,N_24600,N_23086);
nand UO_2479 (O_2479,N_24120,N_22704);
and UO_2480 (O_2480,N_22439,N_24455);
or UO_2481 (O_2481,N_24536,N_24694);
xnor UO_2482 (O_2482,N_23019,N_23130);
xor UO_2483 (O_2483,N_23772,N_22609);
nor UO_2484 (O_2484,N_22027,N_24843);
xnor UO_2485 (O_2485,N_24327,N_24603);
nor UO_2486 (O_2486,N_23882,N_24922);
nand UO_2487 (O_2487,N_22106,N_24023);
and UO_2488 (O_2488,N_24804,N_22403);
nand UO_2489 (O_2489,N_24909,N_24852);
nor UO_2490 (O_2490,N_23457,N_24771);
xor UO_2491 (O_2491,N_23444,N_22755);
or UO_2492 (O_2492,N_23924,N_24907);
or UO_2493 (O_2493,N_23092,N_24021);
nor UO_2494 (O_2494,N_24527,N_23065);
or UO_2495 (O_2495,N_22675,N_22050);
or UO_2496 (O_2496,N_23609,N_22107);
and UO_2497 (O_2497,N_23548,N_23600);
and UO_2498 (O_2498,N_23188,N_22541);
or UO_2499 (O_2499,N_23018,N_23107);
nand UO_2500 (O_2500,N_22892,N_24753);
and UO_2501 (O_2501,N_23125,N_22538);
xor UO_2502 (O_2502,N_23020,N_22825);
nand UO_2503 (O_2503,N_24375,N_22811);
nor UO_2504 (O_2504,N_23897,N_24756);
xor UO_2505 (O_2505,N_24799,N_24165);
nor UO_2506 (O_2506,N_24238,N_24860);
and UO_2507 (O_2507,N_24123,N_23647);
xor UO_2508 (O_2508,N_23963,N_24839);
xor UO_2509 (O_2509,N_22646,N_24668);
and UO_2510 (O_2510,N_24898,N_24784);
nand UO_2511 (O_2511,N_24684,N_23800);
nand UO_2512 (O_2512,N_23526,N_24958);
or UO_2513 (O_2513,N_23895,N_23177);
nand UO_2514 (O_2514,N_23342,N_24858);
and UO_2515 (O_2515,N_24571,N_24007);
xnor UO_2516 (O_2516,N_24982,N_23841);
xnor UO_2517 (O_2517,N_23950,N_21877);
xor UO_2518 (O_2518,N_24336,N_23654);
and UO_2519 (O_2519,N_24923,N_24898);
and UO_2520 (O_2520,N_24635,N_23081);
xnor UO_2521 (O_2521,N_23322,N_21946);
nor UO_2522 (O_2522,N_23277,N_23232);
or UO_2523 (O_2523,N_24602,N_23240);
nor UO_2524 (O_2524,N_22500,N_24273);
and UO_2525 (O_2525,N_23007,N_24960);
or UO_2526 (O_2526,N_22257,N_24684);
or UO_2527 (O_2527,N_24176,N_23773);
or UO_2528 (O_2528,N_24030,N_24414);
nand UO_2529 (O_2529,N_23477,N_24825);
xor UO_2530 (O_2530,N_21928,N_22318);
nor UO_2531 (O_2531,N_24168,N_22364);
xor UO_2532 (O_2532,N_24066,N_24820);
nor UO_2533 (O_2533,N_23996,N_22158);
or UO_2534 (O_2534,N_22759,N_23493);
nor UO_2535 (O_2535,N_22794,N_23627);
nand UO_2536 (O_2536,N_23108,N_23057);
xor UO_2537 (O_2537,N_24779,N_21934);
xor UO_2538 (O_2538,N_22413,N_24517);
nor UO_2539 (O_2539,N_24205,N_24066);
xnor UO_2540 (O_2540,N_24074,N_22629);
and UO_2541 (O_2541,N_22490,N_24135);
or UO_2542 (O_2542,N_23544,N_24518);
nand UO_2543 (O_2543,N_23611,N_23636);
and UO_2544 (O_2544,N_23849,N_24315);
nor UO_2545 (O_2545,N_23123,N_24819);
and UO_2546 (O_2546,N_24913,N_22726);
nor UO_2547 (O_2547,N_22837,N_23232);
xor UO_2548 (O_2548,N_23164,N_23231);
or UO_2549 (O_2549,N_23818,N_24403);
nor UO_2550 (O_2550,N_24283,N_23454);
nor UO_2551 (O_2551,N_24437,N_23427);
nor UO_2552 (O_2552,N_24341,N_22288);
nand UO_2553 (O_2553,N_22320,N_22236);
or UO_2554 (O_2554,N_23454,N_22356);
or UO_2555 (O_2555,N_23577,N_23619);
or UO_2556 (O_2556,N_23790,N_23964);
nor UO_2557 (O_2557,N_24486,N_23820);
xnor UO_2558 (O_2558,N_22639,N_22908);
or UO_2559 (O_2559,N_22016,N_22915);
and UO_2560 (O_2560,N_22166,N_24511);
nand UO_2561 (O_2561,N_23538,N_22146);
nor UO_2562 (O_2562,N_23116,N_24818);
or UO_2563 (O_2563,N_23659,N_24713);
nor UO_2564 (O_2564,N_23353,N_23207);
nand UO_2565 (O_2565,N_22337,N_24271);
or UO_2566 (O_2566,N_24459,N_23586);
nor UO_2567 (O_2567,N_21898,N_23087);
nor UO_2568 (O_2568,N_23040,N_23716);
and UO_2569 (O_2569,N_22220,N_24019);
nand UO_2570 (O_2570,N_23346,N_22560);
xor UO_2571 (O_2571,N_23342,N_23850);
xor UO_2572 (O_2572,N_22585,N_24262);
and UO_2573 (O_2573,N_23359,N_24089);
nor UO_2574 (O_2574,N_23983,N_23505);
or UO_2575 (O_2575,N_22501,N_24360);
nand UO_2576 (O_2576,N_24402,N_23329);
and UO_2577 (O_2577,N_24177,N_24038);
or UO_2578 (O_2578,N_24624,N_22195);
and UO_2579 (O_2579,N_23253,N_24777);
xnor UO_2580 (O_2580,N_22157,N_22659);
and UO_2581 (O_2581,N_23659,N_24254);
xnor UO_2582 (O_2582,N_21907,N_24488);
xnor UO_2583 (O_2583,N_22694,N_22782);
nand UO_2584 (O_2584,N_22889,N_23853);
and UO_2585 (O_2585,N_22180,N_24933);
or UO_2586 (O_2586,N_21984,N_22114);
nor UO_2587 (O_2587,N_22764,N_22876);
xor UO_2588 (O_2588,N_24408,N_24674);
nand UO_2589 (O_2589,N_24506,N_23779);
nor UO_2590 (O_2590,N_24786,N_24002);
or UO_2591 (O_2591,N_23605,N_22976);
nor UO_2592 (O_2592,N_23402,N_24646);
or UO_2593 (O_2593,N_23142,N_22617);
nand UO_2594 (O_2594,N_22355,N_23159);
nor UO_2595 (O_2595,N_22518,N_22937);
xnor UO_2596 (O_2596,N_24902,N_22301);
or UO_2597 (O_2597,N_22717,N_22831);
nor UO_2598 (O_2598,N_23343,N_22297);
nor UO_2599 (O_2599,N_22719,N_23605);
xor UO_2600 (O_2600,N_24955,N_22296);
nor UO_2601 (O_2601,N_24004,N_22058);
or UO_2602 (O_2602,N_23286,N_23898);
nand UO_2603 (O_2603,N_24542,N_22021);
and UO_2604 (O_2604,N_24070,N_23787);
nor UO_2605 (O_2605,N_22055,N_24956);
nor UO_2606 (O_2606,N_21978,N_22528);
xnor UO_2607 (O_2607,N_23353,N_23398);
and UO_2608 (O_2608,N_24089,N_23635);
nand UO_2609 (O_2609,N_23350,N_22709);
or UO_2610 (O_2610,N_24784,N_22324);
xnor UO_2611 (O_2611,N_22181,N_23005);
nor UO_2612 (O_2612,N_23995,N_23365);
nor UO_2613 (O_2613,N_22384,N_23265);
and UO_2614 (O_2614,N_22657,N_22836);
or UO_2615 (O_2615,N_23876,N_22166);
nor UO_2616 (O_2616,N_22027,N_23959);
or UO_2617 (O_2617,N_23384,N_21908);
nand UO_2618 (O_2618,N_24287,N_24835);
or UO_2619 (O_2619,N_24828,N_22128);
and UO_2620 (O_2620,N_23688,N_21925);
and UO_2621 (O_2621,N_23255,N_23266);
xnor UO_2622 (O_2622,N_22254,N_22446);
or UO_2623 (O_2623,N_22662,N_24891);
nor UO_2624 (O_2624,N_23931,N_24782);
nand UO_2625 (O_2625,N_24618,N_23489);
nand UO_2626 (O_2626,N_22679,N_24128);
and UO_2627 (O_2627,N_23642,N_23106);
nand UO_2628 (O_2628,N_21905,N_22287);
xnor UO_2629 (O_2629,N_22339,N_24447);
and UO_2630 (O_2630,N_22936,N_23209);
or UO_2631 (O_2631,N_24744,N_24707);
nand UO_2632 (O_2632,N_23041,N_23637);
xor UO_2633 (O_2633,N_24110,N_22639);
nor UO_2634 (O_2634,N_22661,N_23810);
nand UO_2635 (O_2635,N_23403,N_24475);
nor UO_2636 (O_2636,N_22506,N_24148);
nand UO_2637 (O_2637,N_24795,N_22027);
and UO_2638 (O_2638,N_24423,N_23470);
nor UO_2639 (O_2639,N_23297,N_24965);
and UO_2640 (O_2640,N_24037,N_24637);
nand UO_2641 (O_2641,N_22580,N_22181);
and UO_2642 (O_2642,N_24198,N_21965);
xor UO_2643 (O_2643,N_23284,N_23122);
nand UO_2644 (O_2644,N_22013,N_22740);
xor UO_2645 (O_2645,N_22458,N_24276);
xnor UO_2646 (O_2646,N_23143,N_24014);
and UO_2647 (O_2647,N_23015,N_22645);
nand UO_2648 (O_2648,N_24101,N_24455);
xnor UO_2649 (O_2649,N_22720,N_22985);
and UO_2650 (O_2650,N_23634,N_22352);
and UO_2651 (O_2651,N_22020,N_22884);
xnor UO_2652 (O_2652,N_22629,N_22631);
nor UO_2653 (O_2653,N_22059,N_22102);
nor UO_2654 (O_2654,N_23942,N_22152);
or UO_2655 (O_2655,N_23477,N_24014);
or UO_2656 (O_2656,N_22055,N_24379);
nand UO_2657 (O_2657,N_24532,N_22849);
and UO_2658 (O_2658,N_23755,N_24211);
nor UO_2659 (O_2659,N_23477,N_24044);
xnor UO_2660 (O_2660,N_22664,N_22202);
nor UO_2661 (O_2661,N_24121,N_24033);
and UO_2662 (O_2662,N_22659,N_23719);
and UO_2663 (O_2663,N_24098,N_23819);
nor UO_2664 (O_2664,N_23498,N_24836);
nor UO_2665 (O_2665,N_22330,N_24394);
and UO_2666 (O_2666,N_23508,N_24703);
and UO_2667 (O_2667,N_22713,N_22374);
and UO_2668 (O_2668,N_23600,N_22223);
nand UO_2669 (O_2669,N_24671,N_22423);
nand UO_2670 (O_2670,N_24295,N_24282);
xor UO_2671 (O_2671,N_23226,N_23496);
or UO_2672 (O_2672,N_24338,N_23029);
and UO_2673 (O_2673,N_23296,N_22275);
nor UO_2674 (O_2674,N_23958,N_24731);
nand UO_2675 (O_2675,N_23229,N_23862);
nand UO_2676 (O_2676,N_23688,N_22853);
nand UO_2677 (O_2677,N_22671,N_22446);
and UO_2678 (O_2678,N_24928,N_23281);
and UO_2679 (O_2679,N_24069,N_22106);
or UO_2680 (O_2680,N_22968,N_24588);
and UO_2681 (O_2681,N_22613,N_22446);
xor UO_2682 (O_2682,N_24454,N_23268);
and UO_2683 (O_2683,N_22703,N_23041);
xor UO_2684 (O_2684,N_22113,N_24236);
nand UO_2685 (O_2685,N_22351,N_23859);
and UO_2686 (O_2686,N_22375,N_23354);
or UO_2687 (O_2687,N_22226,N_23978);
xor UO_2688 (O_2688,N_23119,N_22552);
xnor UO_2689 (O_2689,N_24615,N_22993);
nor UO_2690 (O_2690,N_22222,N_24490);
and UO_2691 (O_2691,N_23106,N_23452);
or UO_2692 (O_2692,N_22225,N_22626);
nand UO_2693 (O_2693,N_23200,N_24954);
xor UO_2694 (O_2694,N_24604,N_24214);
and UO_2695 (O_2695,N_23084,N_23012);
xor UO_2696 (O_2696,N_24993,N_22279);
xor UO_2697 (O_2697,N_22995,N_23131);
nand UO_2698 (O_2698,N_24578,N_24562);
nand UO_2699 (O_2699,N_22757,N_23075);
xor UO_2700 (O_2700,N_23399,N_22029);
nor UO_2701 (O_2701,N_22514,N_22958);
nand UO_2702 (O_2702,N_22569,N_24217);
or UO_2703 (O_2703,N_23352,N_24488);
nor UO_2704 (O_2704,N_23909,N_22747);
nand UO_2705 (O_2705,N_22429,N_23547);
nand UO_2706 (O_2706,N_21896,N_24797);
nor UO_2707 (O_2707,N_24072,N_24199);
xor UO_2708 (O_2708,N_24922,N_24736);
and UO_2709 (O_2709,N_22933,N_23644);
and UO_2710 (O_2710,N_23444,N_23071);
or UO_2711 (O_2711,N_22556,N_22835);
and UO_2712 (O_2712,N_22467,N_23667);
and UO_2713 (O_2713,N_24079,N_22798);
and UO_2714 (O_2714,N_23691,N_21906);
and UO_2715 (O_2715,N_23983,N_24521);
nand UO_2716 (O_2716,N_22695,N_24318);
and UO_2717 (O_2717,N_22555,N_23185);
and UO_2718 (O_2718,N_24726,N_24087);
nor UO_2719 (O_2719,N_23781,N_22617);
and UO_2720 (O_2720,N_24420,N_23108);
and UO_2721 (O_2721,N_23884,N_23185);
xnor UO_2722 (O_2722,N_22745,N_21949);
and UO_2723 (O_2723,N_22836,N_24739);
nand UO_2724 (O_2724,N_22807,N_22032);
and UO_2725 (O_2725,N_22638,N_24891);
or UO_2726 (O_2726,N_24054,N_22852);
nand UO_2727 (O_2727,N_24905,N_22252);
nand UO_2728 (O_2728,N_23524,N_24817);
or UO_2729 (O_2729,N_22248,N_22539);
nand UO_2730 (O_2730,N_24700,N_22818);
nand UO_2731 (O_2731,N_23777,N_23221);
and UO_2732 (O_2732,N_24612,N_23581);
and UO_2733 (O_2733,N_23828,N_23469);
xor UO_2734 (O_2734,N_24015,N_22544);
nand UO_2735 (O_2735,N_21932,N_23193);
and UO_2736 (O_2736,N_22630,N_24235);
nand UO_2737 (O_2737,N_22502,N_22466);
nand UO_2738 (O_2738,N_23954,N_24302);
nand UO_2739 (O_2739,N_24908,N_23847);
and UO_2740 (O_2740,N_23608,N_23873);
or UO_2741 (O_2741,N_24819,N_23984);
and UO_2742 (O_2742,N_24002,N_23718);
nor UO_2743 (O_2743,N_24657,N_22307);
xnor UO_2744 (O_2744,N_24882,N_23228);
or UO_2745 (O_2745,N_24820,N_24937);
xnor UO_2746 (O_2746,N_24137,N_24247);
xor UO_2747 (O_2747,N_23547,N_22597);
nor UO_2748 (O_2748,N_24607,N_22494);
xnor UO_2749 (O_2749,N_24576,N_22279);
nor UO_2750 (O_2750,N_22357,N_23974);
or UO_2751 (O_2751,N_23051,N_24587);
xnor UO_2752 (O_2752,N_24782,N_24296);
or UO_2753 (O_2753,N_22439,N_24490);
and UO_2754 (O_2754,N_23462,N_23730);
xnor UO_2755 (O_2755,N_22570,N_24091);
nand UO_2756 (O_2756,N_24891,N_23026);
nor UO_2757 (O_2757,N_23098,N_24379);
xor UO_2758 (O_2758,N_23186,N_23730);
nor UO_2759 (O_2759,N_22118,N_23708);
or UO_2760 (O_2760,N_22093,N_21965);
nor UO_2761 (O_2761,N_22218,N_22020);
xnor UO_2762 (O_2762,N_23502,N_23077);
xnor UO_2763 (O_2763,N_22858,N_23237);
or UO_2764 (O_2764,N_24185,N_22174);
and UO_2765 (O_2765,N_24176,N_22369);
nand UO_2766 (O_2766,N_22628,N_22531);
nor UO_2767 (O_2767,N_24223,N_22196);
nand UO_2768 (O_2768,N_24166,N_22536);
and UO_2769 (O_2769,N_22015,N_24642);
nand UO_2770 (O_2770,N_21902,N_24563);
nor UO_2771 (O_2771,N_22572,N_23381);
nor UO_2772 (O_2772,N_23626,N_23410);
nand UO_2773 (O_2773,N_24310,N_23193);
nor UO_2774 (O_2774,N_23469,N_23126);
nor UO_2775 (O_2775,N_24158,N_22089);
xor UO_2776 (O_2776,N_23919,N_22086);
nor UO_2777 (O_2777,N_22024,N_24364);
nor UO_2778 (O_2778,N_23770,N_24940);
and UO_2779 (O_2779,N_22505,N_24394);
and UO_2780 (O_2780,N_23480,N_24614);
or UO_2781 (O_2781,N_22299,N_24952);
nand UO_2782 (O_2782,N_23340,N_23688);
and UO_2783 (O_2783,N_22393,N_24385);
nor UO_2784 (O_2784,N_24180,N_23100);
nand UO_2785 (O_2785,N_24048,N_22043);
nor UO_2786 (O_2786,N_23785,N_23838);
nor UO_2787 (O_2787,N_24584,N_24377);
xnor UO_2788 (O_2788,N_23910,N_24130);
nor UO_2789 (O_2789,N_24272,N_23457);
nor UO_2790 (O_2790,N_22510,N_23638);
nand UO_2791 (O_2791,N_24217,N_23735);
or UO_2792 (O_2792,N_23560,N_23580);
nor UO_2793 (O_2793,N_21952,N_22667);
xor UO_2794 (O_2794,N_24354,N_24021);
or UO_2795 (O_2795,N_22331,N_24235);
nand UO_2796 (O_2796,N_22044,N_22259);
xor UO_2797 (O_2797,N_23333,N_22681);
nand UO_2798 (O_2798,N_24653,N_23813);
xor UO_2799 (O_2799,N_23998,N_23285);
xnor UO_2800 (O_2800,N_23018,N_23405);
nor UO_2801 (O_2801,N_24581,N_24318);
and UO_2802 (O_2802,N_23635,N_23602);
nor UO_2803 (O_2803,N_22401,N_24627);
nor UO_2804 (O_2804,N_22591,N_23664);
nor UO_2805 (O_2805,N_24930,N_24951);
or UO_2806 (O_2806,N_23999,N_21987);
or UO_2807 (O_2807,N_22652,N_23772);
and UO_2808 (O_2808,N_23689,N_23668);
and UO_2809 (O_2809,N_23638,N_22129);
nand UO_2810 (O_2810,N_23977,N_24250);
xnor UO_2811 (O_2811,N_23038,N_23123);
or UO_2812 (O_2812,N_24746,N_22611);
nand UO_2813 (O_2813,N_22678,N_23604);
or UO_2814 (O_2814,N_23480,N_22455);
or UO_2815 (O_2815,N_23428,N_23390);
and UO_2816 (O_2816,N_23428,N_22513);
nor UO_2817 (O_2817,N_24645,N_22460);
nor UO_2818 (O_2818,N_24137,N_24398);
xor UO_2819 (O_2819,N_24915,N_22924);
xnor UO_2820 (O_2820,N_23105,N_22045);
and UO_2821 (O_2821,N_22636,N_23872);
nand UO_2822 (O_2822,N_23194,N_22146);
nand UO_2823 (O_2823,N_23805,N_22878);
xnor UO_2824 (O_2824,N_23490,N_24193);
and UO_2825 (O_2825,N_23966,N_24244);
or UO_2826 (O_2826,N_22160,N_22742);
nor UO_2827 (O_2827,N_23674,N_23380);
and UO_2828 (O_2828,N_22190,N_23816);
or UO_2829 (O_2829,N_23877,N_23848);
and UO_2830 (O_2830,N_22087,N_22199);
and UO_2831 (O_2831,N_22849,N_24750);
xnor UO_2832 (O_2832,N_23645,N_23678);
nor UO_2833 (O_2833,N_22560,N_23356);
xor UO_2834 (O_2834,N_22237,N_23692);
or UO_2835 (O_2835,N_22566,N_22097);
nor UO_2836 (O_2836,N_22131,N_24453);
xnor UO_2837 (O_2837,N_23605,N_24077);
nand UO_2838 (O_2838,N_24194,N_22135);
or UO_2839 (O_2839,N_23419,N_24979);
nand UO_2840 (O_2840,N_24035,N_22906);
and UO_2841 (O_2841,N_21879,N_23383);
nor UO_2842 (O_2842,N_22298,N_24305);
or UO_2843 (O_2843,N_22777,N_24121);
nor UO_2844 (O_2844,N_24088,N_23236);
nor UO_2845 (O_2845,N_23112,N_22123);
nand UO_2846 (O_2846,N_24219,N_23253);
or UO_2847 (O_2847,N_23889,N_24211);
and UO_2848 (O_2848,N_22106,N_24514);
nor UO_2849 (O_2849,N_23805,N_24967);
or UO_2850 (O_2850,N_21991,N_24117);
or UO_2851 (O_2851,N_24432,N_23691);
and UO_2852 (O_2852,N_24489,N_22466);
nor UO_2853 (O_2853,N_23919,N_23139);
and UO_2854 (O_2854,N_24462,N_24725);
nor UO_2855 (O_2855,N_23411,N_24846);
xor UO_2856 (O_2856,N_23629,N_23807);
and UO_2857 (O_2857,N_24657,N_23950);
xnor UO_2858 (O_2858,N_23316,N_24976);
and UO_2859 (O_2859,N_22043,N_23958);
nand UO_2860 (O_2860,N_24151,N_22072);
nor UO_2861 (O_2861,N_22845,N_24540);
and UO_2862 (O_2862,N_23688,N_24935);
xor UO_2863 (O_2863,N_23084,N_23666);
and UO_2864 (O_2864,N_22160,N_23135);
or UO_2865 (O_2865,N_23709,N_22003);
nor UO_2866 (O_2866,N_22891,N_23230);
or UO_2867 (O_2867,N_22425,N_21921);
and UO_2868 (O_2868,N_23553,N_23370);
xnor UO_2869 (O_2869,N_24191,N_24849);
nand UO_2870 (O_2870,N_22994,N_24965);
or UO_2871 (O_2871,N_24117,N_22327);
nand UO_2872 (O_2872,N_22153,N_24049);
nand UO_2873 (O_2873,N_22055,N_24409);
and UO_2874 (O_2874,N_23672,N_23949);
and UO_2875 (O_2875,N_23098,N_22460);
nor UO_2876 (O_2876,N_23785,N_23314);
nand UO_2877 (O_2877,N_24331,N_22964);
nor UO_2878 (O_2878,N_22964,N_23830);
xnor UO_2879 (O_2879,N_22439,N_22218);
nand UO_2880 (O_2880,N_24536,N_24349);
and UO_2881 (O_2881,N_23246,N_23121);
nor UO_2882 (O_2882,N_22922,N_24595);
and UO_2883 (O_2883,N_21995,N_24652);
xnor UO_2884 (O_2884,N_23572,N_24594);
and UO_2885 (O_2885,N_22406,N_23248);
or UO_2886 (O_2886,N_24599,N_23603);
nor UO_2887 (O_2887,N_23543,N_23998);
nand UO_2888 (O_2888,N_22150,N_22354);
or UO_2889 (O_2889,N_24334,N_24793);
nor UO_2890 (O_2890,N_22091,N_23145);
xnor UO_2891 (O_2891,N_22467,N_22641);
nand UO_2892 (O_2892,N_23492,N_23113);
and UO_2893 (O_2893,N_24850,N_23295);
nand UO_2894 (O_2894,N_22322,N_22720);
and UO_2895 (O_2895,N_21905,N_23066);
xor UO_2896 (O_2896,N_22483,N_24142);
or UO_2897 (O_2897,N_22119,N_23160);
nand UO_2898 (O_2898,N_24792,N_23833);
or UO_2899 (O_2899,N_24991,N_24069);
or UO_2900 (O_2900,N_23883,N_23591);
nor UO_2901 (O_2901,N_24529,N_22596);
xnor UO_2902 (O_2902,N_23617,N_24135);
nand UO_2903 (O_2903,N_22134,N_22451);
nor UO_2904 (O_2904,N_24552,N_23005);
nand UO_2905 (O_2905,N_22322,N_22686);
nor UO_2906 (O_2906,N_22886,N_22555);
or UO_2907 (O_2907,N_22343,N_22112);
and UO_2908 (O_2908,N_23730,N_23971);
and UO_2909 (O_2909,N_24093,N_24549);
nand UO_2910 (O_2910,N_23932,N_24257);
nor UO_2911 (O_2911,N_22581,N_22881);
and UO_2912 (O_2912,N_24085,N_23128);
nand UO_2913 (O_2913,N_24477,N_22596);
xor UO_2914 (O_2914,N_24448,N_24517);
xor UO_2915 (O_2915,N_22177,N_22449);
nand UO_2916 (O_2916,N_21908,N_22055);
and UO_2917 (O_2917,N_22995,N_23555);
nand UO_2918 (O_2918,N_22434,N_24598);
xor UO_2919 (O_2919,N_22263,N_21968);
or UO_2920 (O_2920,N_24814,N_22573);
nor UO_2921 (O_2921,N_23783,N_23406);
nand UO_2922 (O_2922,N_22680,N_22813);
and UO_2923 (O_2923,N_23533,N_23659);
and UO_2924 (O_2924,N_22740,N_22913);
and UO_2925 (O_2925,N_24740,N_23145);
or UO_2926 (O_2926,N_24371,N_22582);
or UO_2927 (O_2927,N_24008,N_24883);
and UO_2928 (O_2928,N_24735,N_23487);
nand UO_2929 (O_2929,N_23536,N_22535);
or UO_2930 (O_2930,N_22152,N_21973);
xnor UO_2931 (O_2931,N_24589,N_24291);
nand UO_2932 (O_2932,N_22121,N_23139);
xor UO_2933 (O_2933,N_23984,N_24934);
nor UO_2934 (O_2934,N_22075,N_23072);
or UO_2935 (O_2935,N_23886,N_23644);
and UO_2936 (O_2936,N_22217,N_22144);
and UO_2937 (O_2937,N_23968,N_21964);
nand UO_2938 (O_2938,N_22907,N_22676);
and UO_2939 (O_2939,N_22745,N_23546);
nand UO_2940 (O_2940,N_23672,N_23916);
xor UO_2941 (O_2941,N_24979,N_24489);
xor UO_2942 (O_2942,N_22756,N_22052);
nor UO_2943 (O_2943,N_21902,N_22492);
xor UO_2944 (O_2944,N_23400,N_24248);
nand UO_2945 (O_2945,N_22505,N_24355);
nand UO_2946 (O_2946,N_24002,N_21954);
xnor UO_2947 (O_2947,N_23290,N_22503);
xor UO_2948 (O_2948,N_24432,N_23789);
nand UO_2949 (O_2949,N_22167,N_24693);
or UO_2950 (O_2950,N_22863,N_22484);
and UO_2951 (O_2951,N_22977,N_24710);
xor UO_2952 (O_2952,N_22609,N_24399);
and UO_2953 (O_2953,N_23515,N_22430);
nor UO_2954 (O_2954,N_23777,N_23444);
xnor UO_2955 (O_2955,N_23568,N_22795);
nand UO_2956 (O_2956,N_24824,N_22389);
or UO_2957 (O_2957,N_22302,N_23415);
xnor UO_2958 (O_2958,N_22894,N_24924);
xnor UO_2959 (O_2959,N_23233,N_21993);
or UO_2960 (O_2960,N_23886,N_22761);
nand UO_2961 (O_2961,N_23378,N_23289);
nand UO_2962 (O_2962,N_23133,N_22401);
xor UO_2963 (O_2963,N_22270,N_23912);
nor UO_2964 (O_2964,N_22901,N_23377);
nand UO_2965 (O_2965,N_23736,N_23200);
nand UO_2966 (O_2966,N_23981,N_24184);
or UO_2967 (O_2967,N_22384,N_22998);
and UO_2968 (O_2968,N_22847,N_24053);
nor UO_2969 (O_2969,N_23704,N_23320);
nor UO_2970 (O_2970,N_24102,N_22878);
and UO_2971 (O_2971,N_22494,N_23649);
and UO_2972 (O_2972,N_23031,N_22332);
and UO_2973 (O_2973,N_22416,N_21928);
and UO_2974 (O_2974,N_22444,N_23964);
or UO_2975 (O_2975,N_22780,N_23303);
nand UO_2976 (O_2976,N_21911,N_24574);
nand UO_2977 (O_2977,N_22012,N_23863);
or UO_2978 (O_2978,N_22441,N_23255);
or UO_2979 (O_2979,N_22643,N_21981);
xnor UO_2980 (O_2980,N_21983,N_24877);
xnor UO_2981 (O_2981,N_22901,N_23926);
and UO_2982 (O_2982,N_21884,N_24654);
and UO_2983 (O_2983,N_22663,N_24942);
or UO_2984 (O_2984,N_24158,N_21884);
nor UO_2985 (O_2985,N_23747,N_24665);
and UO_2986 (O_2986,N_24119,N_22065);
or UO_2987 (O_2987,N_23414,N_22341);
nand UO_2988 (O_2988,N_23450,N_22245);
nand UO_2989 (O_2989,N_22084,N_23620);
nor UO_2990 (O_2990,N_22237,N_24302);
or UO_2991 (O_2991,N_21893,N_23866);
nor UO_2992 (O_2992,N_24670,N_24207);
nand UO_2993 (O_2993,N_24858,N_22189);
and UO_2994 (O_2994,N_24501,N_22760);
xor UO_2995 (O_2995,N_24350,N_24925);
and UO_2996 (O_2996,N_24165,N_22160);
nand UO_2997 (O_2997,N_22860,N_23758);
nand UO_2998 (O_2998,N_22897,N_24004);
nor UO_2999 (O_2999,N_22808,N_23198);
endmodule