module basic_3000_30000_3500_5_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_1572,In_146);
nand U1 (N_1,In_57,In_2000);
nand U2 (N_2,In_2864,In_1505);
xor U3 (N_3,In_2982,In_2813);
nor U4 (N_4,In_1188,In_2312);
and U5 (N_5,In_1109,In_386);
nor U6 (N_6,In_588,In_688);
nand U7 (N_7,In_2193,In_2969);
and U8 (N_8,In_527,In_2138);
nor U9 (N_9,In_2773,In_1361);
nand U10 (N_10,In_149,In_1859);
xor U11 (N_11,In_1267,In_547);
nor U12 (N_12,In_981,In_1062);
nor U13 (N_13,In_2380,In_2103);
or U14 (N_14,In_2277,In_1970);
nor U15 (N_15,In_39,In_2572);
or U16 (N_16,In_2639,In_2266);
or U17 (N_17,In_2025,In_1996);
nor U18 (N_18,In_1264,In_1892);
or U19 (N_19,In_1819,In_1404);
or U20 (N_20,In_2446,In_69);
nor U21 (N_21,In_1373,In_2663);
and U22 (N_22,In_1981,In_1425);
nor U23 (N_23,In_1318,In_179);
or U24 (N_24,In_303,In_2286);
and U25 (N_25,In_1135,In_1215);
or U26 (N_26,In_2698,In_1847);
and U27 (N_27,In_1957,In_2467);
nor U28 (N_28,In_733,In_283);
nor U29 (N_29,In_2192,In_502);
and U30 (N_30,In_1252,In_480);
or U31 (N_31,In_40,In_2665);
nor U32 (N_32,In_1935,In_1219);
xor U33 (N_33,In_1734,In_2974);
nor U34 (N_34,In_2756,In_160);
nor U35 (N_35,In_956,In_2261);
or U36 (N_36,In_1488,In_892);
nand U37 (N_37,In_1469,In_2352);
and U38 (N_38,In_881,In_2462);
and U39 (N_39,In_2166,In_854);
nand U40 (N_40,In_799,In_853);
nand U41 (N_41,In_1484,In_2408);
or U42 (N_42,In_1688,In_1973);
or U43 (N_43,In_1250,In_2280);
nor U44 (N_44,In_1832,In_2476);
nand U45 (N_45,In_319,In_68);
xor U46 (N_46,In_1855,In_47);
nor U47 (N_47,In_2811,In_2056);
and U48 (N_48,In_1416,In_1430);
or U49 (N_49,In_106,In_789);
nor U50 (N_50,In_1100,In_358);
nand U51 (N_51,In_337,In_1339);
nand U52 (N_52,In_1843,In_278);
and U53 (N_53,In_1291,In_1516);
nor U54 (N_54,In_2918,In_56);
nand U55 (N_55,In_1679,In_2851);
or U56 (N_56,In_1966,In_1174);
or U57 (N_57,In_1553,In_394);
nor U58 (N_58,In_2589,In_2976);
and U59 (N_59,In_2066,In_219);
nand U60 (N_60,In_2619,In_66);
nand U61 (N_61,In_1104,In_1084);
and U62 (N_62,In_1586,In_2609);
nor U63 (N_63,In_584,In_1282);
nor U64 (N_64,In_2256,In_776);
nor U65 (N_65,In_510,In_1865);
nand U66 (N_66,In_167,In_1671);
or U67 (N_67,In_1853,In_1313);
nand U68 (N_68,In_2608,In_411);
or U69 (N_69,In_335,In_984);
nand U70 (N_70,In_2559,In_541);
nand U71 (N_71,In_2959,In_388);
nand U72 (N_72,In_1392,In_97);
or U73 (N_73,In_2412,In_828);
and U74 (N_74,In_662,In_2223);
and U75 (N_75,In_1501,In_1414);
nand U76 (N_76,In_624,In_1930);
nand U77 (N_77,In_2059,In_2264);
and U78 (N_78,In_1089,In_427);
xnor U79 (N_79,In_1106,In_157);
and U80 (N_80,In_629,In_1824);
nand U81 (N_81,In_138,In_650);
nand U82 (N_82,In_2506,In_1020);
nand U83 (N_83,In_431,In_1479);
and U84 (N_84,In_867,In_1415);
nor U85 (N_85,In_1003,In_2486);
nand U86 (N_86,In_2791,In_465);
or U87 (N_87,In_2374,In_2510);
nand U88 (N_88,In_1105,In_1461);
nand U89 (N_89,In_1166,In_1682);
nand U90 (N_90,In_875,In_2160);
nand U91 (N_91,In_1569,In_2963);
nand U92 (N_92,In_1451,In_229);
and U93 (N_93,In_1377,In_145);
xor U94 (N_94,In_2719,In_2672);
or U95 (N_95,In_1296,In_1483);
or U96 (N_96,In_1117,In_581);
or U97 (N_97,In_2485,In_131);
or U98 (N_98,In_1093,In_89);
nor U99 (N_99,In_1366,In_2575);
xnor U100 (N_100,In_2675,In_1846);
or U101 (N_101,In_1779,In_1059);
and U102 (N_102,In_2368,In_2202);
nand U103 (N_103,In_834,In_945);
nand U104 (N_104,In_2788,In_2375);
xor U105 (N_105,In_1324,In_509);
nand U106 (N_106,In_2937,In_1199);
or U107 (N_107,In_468,In_2776);
nand U108 (N_108,In_304,In_1011);
nor U109 (N_109,In_1588,In_2117);
or U110 (N_110,In_2095,In_1288);
or U111 (N_111,In_2074,In_2364);
nand U112 (N_112,In_463,In_1295);
nand U113 (N_113,In_320,In_1172);
nand U114 (N_114,In_477,In_1471);
nor U115 (N_115,In_349,In_1090);
xnor U116 (N_116,In_2764,In_2819);
or U117 (N_117,In_1611,In_955);
or U118 (N_118,In_2822,In_762);
and U119 (N_119,In_884,In_2544);
nor U120 (N_120,In_1702,In_125);
nor U121 (N_121,In_2898,In_1103);
nand U122 (N_122,In_2818,In_511);
xor U123 (N_123,In_372,In_2817);
nor U124 (N_124,In_2058,In_330);
nand U125 (N_125,In_185,In_1458);
nor U126 (N_126,In_2883,In_1350);
or U127 (N_127,In_2253,In_2186);
nand U128 (N_128,In_1351,In_1725);
and U129 (N_129,In_603,In_1364);
nor U130 (N_130,In_2617,In_393);
nand U131 (N_131,In_2378,In_2042);
nand U132 (N_132,In_428,In_2112);
or U133 (N_133,In_1085,In_2465);
or U134 (N_134,In_1821,In_1396);
xor U135 (N_135,In_381,In_2371);
nor U136 (N_136,In_1612,In_1420);
or U137 (N_137,In_1137,In_753);
or U138 (N_138,In_1744,In_62);
and U139 (N_139,In_1998,In_1889);
or U140 (N_140,In_2916,In_2793);
and U141 (N_141,In_269,In_1222);
xor U142 (N_142,In_1335,In_748);
or U143 (N_143,In_2697,In_860);
nand U144 (N_144,In_276,In_2988);
nand U145 (N_145,In_1781,In_931);
or U146 (N_146,In_1619,In_247);
nand U147 (N_147,In_2876,In_2020);
xnor U148 (N_148,In_2111,In_1606);
and U149 (N_149,In_437,In_2413);
nor U150 (N_150,In_2523,In_113);
nor U151 (N_151,In_1058,In_134);
or U152 (N_152,In_1573,In_1309);
or U153 (N_153,In_2315,In_870);
and U154 (N_154,In_2552,In_2120);
nor U155 (N_155,In_2322,In_2291);
or U156 (N_156,In_2854,In_470);
nand U157 (N_157,In_245,In_2760);
or U158 (N_158,In_637,In_512);
and U159 (N_159,In_542,In_1258);
and U160 (N_160,In_2005,In_1659);
and U161 (N_161,In_765,In_992);
xnor U162 (N_162,In_1810,In_1359);
and U163 (N_163,In_143,In_432);
nor U164 (N_164,In_1560,In_1475);
nor U165 (N_165,In_362,In_930);
and U166 (N_166,In_744,In_120);
nand U167 (N_167,In_329,In_1876);
nand U168 (N_168,In_2447,In_2231);
and U169 (N_169,In_205,In_2442);
nand U170 (N_170,In_2070,In_48);
nor U171 (N_171,In_1503,In_1861);
and U172 (N_172,In_1535,In_743);
nor U173 (N_173,In_2248,In_2569);
or U174 (N_174,In_2328,In_666);
nand U175 (N_175,In_2068,In_289);
nor U176 (N_176,In_2611,In_1525);
nor U177 (N_177,In_346,In_2757);
and U178 (N_178,In_2037,In_136);
nor U179 (N_179,In_1745,In_1695);
nand U180 (N_180,In_2382,In_310);
and U181 (N_181,In_2782,In_162);
or U182 (N_182,In_1078,In_1526);
nand U183 (N_183,In_2923,In_1774);
nor U184 (N_184,In_475,In_2132);
and U185 (N_185,In_872,In_2955);
and U186 (N_186,In_32,In_2509);
or U187 (N_187,In_10,In_2327);
nand U188 (N_188,In_345,In_2423);
and U189 (N_189,In_2593,In_2420);
nor U190 (N_190,In_1589,In_1620);
nand U191 (N_191,In_922,In_779);
nor U192 (N_192,In_739,In_371);
nand U193 (N_193,In_911,In_2432);
nand U194 (N_194,In_946,In_31);
or U195 (N_195,In_1183,In_67);
nor U196 (N_196,In_2795,In_1086);
or U197 (N_197,In_2054,In_1439);
or U198 (N_198,In_2718,In_771);
nor U199 (N_199,In_2688,In_2389);
nor U200 (N_200,In_2363,In_1294);
nand U201 (N_201,In_1685,In_2499);
or U202 (N_202,In_1253,In_2689);
nand U203 (N_203,In_313,In_667);
or U204 (N_204,In_1205,In_843);
nor U205 (N_205,In_2507,In_116);
nand U206 (N_206,In_985,In_1424);
and U207 (N_207,In_1827,In_101);
xor U208 (N_208,In_2733,In_497);
and U209 (N_209,In_1663,In_1013);
nor U210 (N_210,In_1808,In_1795);
or U211 (N_211,In_2500,In_696);
nand U212 (N_212,In_1585,In_953);
nand U213 (N_213,In_2227,In_1196);
and U214 (N_214,In_2038,In_1382);
nor U215 (N_215,In_77,In_2136);
or U216 (N_216,In_830,In_1527);
or U217 (N_217,In_2388,In_780);
nand U218 (N_218,In_2522,In_807);
nor U219 (N_219,In_1164,In_916);
or U220 (N_220,In_1767,In_2105);
nor U221 (N_221,In_2779,In_1446);
nand U222 (N_222,In_248,In_2449);
xnor U223 (N_223,In_2027,In_1074);
nor U224 (N_224,In_2367,In_1736);
nand U225 (N_225,In_257,In_2536);
and U226 (N_226,In_1480,In_1203);
nor U227 (N_227,In_2177,In_2118);
or U228 (N_228,In_2631,In_2612);
or U229 (N_229,In_1434,In_2743);
nand U230 (N_230,In_2653,In_1593);
nor U231 (N_231,In_2821,In_284);
and U232 (N_232,In_443,In_1951);
nor U233 (N_233,In_2668,In_920);
or U234 (N_234,In_543,In_2796);
and U235 (N_235,In_159,In_2961);
or U236 (N_236,In_615,In_1985);
nand U237 (N_237,In_2513,In_2532);
nor U238 (N_238,In_2100,In_706);
or U239 (N_239,In_2574,In_2910);
nand U240 (N_240,In_2828,In_2621);
nand U241 (N_241,In_2723,In_1642);
or U242 (N_242,In_2339,In_2144);
and U243 (N_243,In_1159,In_453);
nand U244 (N_244,In_260,In_2369);
and U245 (N_245,In_569,In_439);
nor U246 (N_246,In_1257,In_2043);
and U247 (N_247,In_929,In_1750);
nor U248 (N_248,In_684,In_1529);
nor U249 (N_249,In_2094,In_117);
or U250 (N_250,In_1518,In_212);
xnor U251 (N_251,In_2983,In_1707);
nor U252 (N_252,In_261,In_732);
nand U253 (N_253,In_1850,In_561);
nor U254 (N_254,In_2548,In_1374);
or U255 (N_255,In_221,In_2366);
and U256 (N_256,In_1757,In_791);
nand U257 (N_257,In_2155,In_1057);
nor U258 (N_258,In_2474,In_2889);
nand U259 (N_259,In_523,In_2767);
nor U260 (N_260,In_1605,In_2247);
nand U261 (N_261,In_1363,In_363);
nand U262 (N_262,In_2727,In_558);
or U263 (N_263,In_1822,In_2057);
xor U264 (N_264,In_176,In_11);
nor U265 (N_265,In_2754,In_2786);
nor U266 (N_266,In_22,In_1595);
nand U267 (N_267,In_2827,In_719);
nand U268 (N_268,In_1860,In_406);
or U269 (N_269,In_1330,In_2586);
nand U270 (N_270,In_396,In_2659);
or U271 (N_271,In_2929,In_438);
and U272 (N_272,In_2133,In_175);
or U273 (N_273,In_1289,In_1390);
nor U274 (N_274,In_573,In_1928);
or U275 (N_275,In_2625,In_1340);
nand U276 (N_276,In_1036,In_96);
xnor U277 (N_277,In_2069,In_1581);
or U278 (N_278,In_1758,In_49);
and U279 (N_279,In_321,In_530);
and U280 (N_280,In_1095,In_2637);
nand U281 (N_281,In_2064,In_2613);
or U282 (N_282,In_2571,In_677);
xor U283 (N_283,In_2805,In_1844);
and U284 (N_284,In_1706,In_173);
and U285 (N_285,In_75,In_856);
or U286 (N_286,In_1443,In_2207);
or U287 (N_287,In_2694,In_1170);
and U288 (N_288,In_1385,In_354);
nor U289 (N_289,In_2157,In_2319);
nor U290 (N_290,In_1506,In_2201);
and U291 (N_291,In_1438,In_2798);
nor U292 (N_292,In_648,In_1353);
nand U293 (N_293,In_1358,In_426);
xor U294 (N_294,In_378,In_1990);
nand U295 (N_295,In_2334,In_1221);
and U296 (N_296,In_938,In_2568);
nor U297 (N_297,In_1580,In_2902);
xor U298 (N_298,In_2610,In_2416);
or U299 (N_299,In_1919,In_2715);
nand U300 (N_300,In_1091,In_1591);
and U301 (N_301,In_1684,In_1213);
nor U302 (N_302,In_2564,In_1741);
or U303 (N_303,In_2736,In_1532);
nor U304 (N_304,In_2726,In_1198);
or U305 (N_305,In_846,In_1840);
nor U306 (N_306,In_1699,In_92);
nor U307 (N_307,In_452,In_1770);
and U308 (N_308,In_1854,In_1913);
and U309 (N_309,In_1791,In_2224);
nand U310 (N_310,In_1692,In_1356);
nand U311 (N_311,In_1748,In_2320);
nor U312 (N_312,In_2946,In_2336);
nor U313 (N_313,In_130,In_2872);
nand U314 (N_314,In_522,In_2618);
nand U315 (N_315,In_1407,In_1060);
or U316 (N_316,In_2867,In_763);
nand U317 (N_317,In_190,In_1600);
nand U318 (N_318,In_2342,In_647);
and U319 (N_319,In_424,In_1926);
or U320 (N_320,In_960,In_2843);
and U321 (N_321,In_2897,In_1680);
nand U322 (N_322,In_506,In_626);
nor U323 (N_323,In_727,In_1958);
nor U324 (N_324,In_1175,In_1900);
nor U325 (N_325,In_536,In_1557);
and U326 (N_326,In_1670,In_1216);
and U327 (N_327,In_1440,In_832);
nor U328 (N_328,In_2550,In_2826);
nand U329 (N_329,In_232,In_606);
nor U330 (N_330,In_1715,In_366);
and U331 (N_331,In_2932,In_640);
nor U332 (N_332,In_1977,In_2908);
nor U333 (N_333,In_817,In_1035);
xnor U334 (N_334,In_1409,In_2886);
or U335 (N_335,In_1837,In_2497);
or U336 (N_336,In_1485,In_2181);
or U337 (N_337,In_1650,In_2210);
or U338 (N_338,In_1754,In_226);
nand U339 (N_339,In_585,In_1602);
nand U340 (N_340,In_2987,In_118);
and U341 (N_341,In_620,In_1823);
nand U342 (N_342,In_1281,In_1131);
and U343 (N_343,In_2451,In_2478);
or U344 (N_344,In_769,In_2021);
nor U345 (N_345,In_2847,In_1329);
nand U346 (N_346,In_1435,In_27);
nand U347 (N_347,In_2372,In_2079);
or U348 (N_348,In_180,In_1194);
nor U349 (N_349,In_1649,In_713);
nand U350 (N_350,In_1890,In_154);
nand U351 (N_351,In_1422,In_1070);
nand U352 (N_352,In_192,In_2862);
nand U353 (N_353,In_605,In_2833);
nand U354 (N_354,In_2089,In_1676);
and U355 (N_355,In_1631,In_1590);
and U356 (N_356,In_155,In_773);
and U357 (N_357,In_1369,In_2707);
nor U358 (N_358,In_2126,In_794);
or U359 (N_359,In_105,In_2925);
nor U360 (N_360,In_628,In_2525);
or U361 (N_361,In_2404,In_1197);
xor U362 (N_362,In_836,In_1337);
and U363 (N_363,In_350,In_2706);
nand U364 (N_364,In_2134,In_312);
and U365 (N_365,In_1232,In_975);
nand U366 (N_366,In_815,In_781);
nor U367 (N_367,In_989,In_1597);
nor U368 (N_368,In_577,In_1749);
nor U369 (N_369,In_1381,In_2681);
xor U370 (N_370,In_2746,In_2195);
and U371 (N_371,In_1897,In_994);
nor U372 (N_372,In_2724,In_2952);
nor U373 (N_373,In_1974,In_957);
nor U374 (N_374,In_1940,In_2645);
nand U375 (N_375,In_1127,In_2119);
and U376 (N_376,In_360,In_1755);
nor U377 (N_377,In_2236,In_775);
nand U378 (N_378,In_292,In_1120);
or U379 (N_379,In_1955,In_464);
or U380 (N_380,In_58,In_766);
xor U381 (N_381,In_1761,In_1730);
nor U382 (N_382,In_2211,In_395);
and U383 (N_383,In_2104,In_2311);
and U384 (N_384,In_579,In_1261);
nand U385 (N_385,In_2191,In_2762);
and U386 (N_386,In_1561,In_1923);
or U387 (N_387,In_1201,In_908);
nand U388 (N_388,In_2578,In_2942);
and U389 (N_389,In_783,In_2445);
and U390 (N_390,In_2106,In_1675);
or U391 (N_391,In_2588,In_1852);
nand U392 (N_392,In_1010,In_2686);
and U393 (N_393,In_268,In_29);
nand U394 (N_394,In_575,In_2088);
or U395 (N_395,In_897,In_2650);
nor U396 (N_396,In_2953,In_2622);
and U397 (N_397,In_376,In_1703);
nor U398 (N_398,In_413,In_306);
and U399 (N_399,In_1555,In_1255);
nor U400 (N_400,In_135,In_1457);
and U401 (N_401,In_2669,In_2285);
nand U402 (N_402,In_988,In_2071);
nor U403 (N_403,In_1621,In_1541);
or U404 (N_404,In_1660,In_2212);
nor U405 (N_405,In_2390,In_1155);
xor U406 (N_406,In_2329,In_1528);
nor U407 (N_407,In_1136,In_1574);
xnor U408 (N_408,In_2085,In_2199);
and U409 (N_409,In_364,In_2062);
nand U410 (N_410,In_137,In_802);
nor U411 (N_411,In_1584,In_2018);
nor U412 (N_412,In_1302,In_926);
nor U413 (N_413,In_222,In_531);
nor U414 (N_414,In_72,In_215);
and U415 (N_415,In_2415,In_1993);
nor U416 (N_416,In_2855,In_950);
nor U417 (N_417,In_1320,In_2538);
and U418 (N_418,In_2287,In_768);
nor U419 (N_419,In_2794,In_2274);
nor U420 (N_420,In_1956,In_2083);
or U421 (N_421,In_170,In_1021);
or U422 (N_422,In_2182,In_824);
nor U423 (N_423,In_14,In_379);
nor U424 (N_424,In_2091,In_1841);
xnor U425 (N_425,In_1274,In_1793);
xor U426 (N_426,In_2377,In_1980);
nor U427 (N_427,In_2081,In_1220);
nand U428 (N_428,In_2824,In_2951);
nand U429 (N_429,In_2985,In_457);
nor U430 (N_430,In_840,In_2221);
xor U431 (N_431,In_2643,In_1906);
nand U432 (N_432,In_741,In_2906);
and U433 (N_433,In_1231,In_2080);
and U434 (N_434,In_905,In_1907);
xor U435 (N_435,In_1206,In_866);
or U436 (N_436,In_1939,In_652);
nand U437 (N_437,In_545,In_2188);
and U438 (N_438,In_886,In_2147);
nor U439 (N_439,In_38,In_1486);
nor U440 (N_440,In_844,In_1729);
nor U441 (N_441,In_1514,In_2986);
nor U442 (N_442,In_2019,In_2204);
and U443 (N_443,In_2825,In_1144);
nor U444 (N_444,In_1708,In_1018);
and U445 (N_445,In_384,In_2996);
or U446 (N_446,In_1121,In_2479);
nor U447 (N_447,In_1563,In_2852);
nor U448 (N_448,In_1971,In_1798);
and U449 (N_449,In_252,In_1716);
nand U450 (N_450,In_2428,In_1494);
or U451 (N_451,In_1427,In_1613);
and U452 (N_452,In_2711,In_391);
and U453 (N_453,In_2594,In_233);
or U454 (N_454,In_811,In_2849);
and U455 (N_455,In_1604,In_1478);
nor U456 (N_456,In_2678,In_474);
nor U457 (N_457,In_639,In_2321);
nor U458 (N_458,In_951,In_1130);
nor U459 (N_459,In_991,In_1632);
nor U460 (N_460,In_2801,In_1043);
and U461 (N_461,In_2127,In_507);
or U462 (N_462,In_1567,In_1936);
and U463 (N_463,In_710,In_128);
and U464 (N_464,In_2283,In_838);
xor U465 (N_465,In_2272,In_446);
and U466 (N_466,In_322,In_1298);
and U467 (N_467,In_2244,In_2735);
or U468 (N_468,In_2999,In_2587);
and U469 (N_469,In_2721,In_147);
xor U470 (N_470,In_1508,In_847);
xnor U471 (N_471,In_1524,In_976);
xnor U472 (N_472,In_2964,In_2885);
or U473 (N_473,In_977,In_2443);
and U474 (N_474,In_2099,In_2734);
or U475 (N_475,In_1248,In_936);
nor U476 (N_476,In_2324,In_2956);
nor U477 (N_477,In_202,In_2225);
xor U478 (N_478,In_1323,In_961);
or U479 (N_479,In_265,In_2832);
or U480 (N_480,In_534,In_583);
and U481 (N_481,In_2338,In_2815);
xor U482 (N_482,In_1829,In_1107);
and U483 (N_483,In_1497,In_1006);
nor U484 (N_484,In_2573,In_2582);
or U485 (N_485,In_1719,In_728);
xnor U486 (N_486,In_927,In_669);
nand U487 (N_487,In_759,In_2783);
or U488 (N_488,In_1212,In_1635);
nor U489 (N_489,In_2030,In_441);
xor U490 (N_490,In_1234,In_369);
nand U491 (N_491,In_259,In_2419);
and U492 (N_492,In_987,In_1038);
and U493 (N_493,In_1735,In_1881);
and U494 (N_494,In_1163,In_887);
or U495 (N_495,In_1262,In_78);
or U496 (N_496,In_2434,In_2850);
nand U497 (N_497,In_234,In_2973);
and U498 (N_498,In_1110,In_1065);
xnor U499 (N_499,In_2161,In_2029);
nor U500 (N_500,In_286,In_2804);
nand U501 (N_501,In_1646,In_2017);
xor U502 (N_502,In_1153,In_2458);
or U503 (N_503,In_2632,In_2131);
or U504 (N_504,In_1500,In_2935);
xnor U505 (N_505,In_1879,In_334);
or U506 (N_506,In_1720,In_756);
nor U507 (N_507,In_1113,In_2024);
and U508 (N_508,In_643,In_2122);
xnor U509 (N_509,In_852,In_857);
nand U510 (N_510,In_1332,In_1976);
nand U511 (N_511,In_693,In_1418);
nor U512 (N_512,In_150,In_2927);
nand U513 (N_513,In_1717,In_570);
nor U514 (N_514,In_1046,In_2597);
or U515 (N_515,In_642,In_2418);
xnor U516 (N_516,In_1229,In_1016);
nor U517 (N_517,In_1811,In_712);
nor U518 (N_518,In_409,In_2992);
or U519 (N_519,In_2217,In_673);
nand U520 (N_520,In_896,In_1030);
nand U521 (N_521,In_2866,In_20);
nand U522 (N_522,In_2016,In_1972);
and U523 (N_523,In_999,In_2905);
nor U524 (N_524,In_2269,In_1979);
nor U525 (N_525,In_770,In_2863);
nor U526 (N_526,In_1277,In_572);
nor U527 (N_527,In_513,In_932);
and U528 (N_528,In_1538,In_1368);
nand U529 (N_529,In_448,In_385);
nor U530 (N_530,In_1967,In_2333);
nor U531 (N_531,In_1962,In_958);
nand U532 (N_532,In_602,In_2163);
nor U533 (N_533,In_187,In_1347);
and U534 (N_534,In_1934,In_1517);
and U535 (N_535,In_1143,In_1389);
xor U536 (N_536,In_2162,In_736);
and U537 (N_537,In_1417,In_525);
or U538 (N_538,In_1796,In_2421);
or U539 (N_539,In_367,In_1061);
and U540 (N_540,In_627,In_718);
nand U541 (N_541,In_2470,In_1269);
or U542 (N_542,In_355,In_670);
nand U543 (N_543,In_383,In_2781);
xor U544 (N_544,In_1053,In_1807);
and U545 (N_545,In_343,In_2948);
and U546 (N_546,In_1386,In_1047);
or U547 (N_547,In_559,In_754);
and U548 (N_548,In_1815,In_2472);
nand U549 (N_549,In_340,In_1783);
and U550 (N_550,In_469,In_2218);
nand U551 (N_551,In_1097,In_742);
and U552 (N_552,In_244,In_1009);
and U553 (N_553,In_788,In_2841);
or U554 (N_554,In_2279,In_979);
and U555 (N_555,In_1872,In_634);
or U556 (N_556,In_86,In_1942);
nor U557 (N_557,In_1237,In_2417);
or U558 (N_558,In_871,In_102);
and U559 (N_559,In_2528,In_2556);
or U560 (N_560,In_1950,In_1017);
or U561 (N_561,In_1833,In_2926);
nand U562 (N_562,In_2171,In_2975);
nand U563 (N_563,In_2304,In_2243);
and U564 (N_564,In_883,In_392);
and U565 (N_565,In_1738,In_2687);
and U566 (N_566,In_1665,In_2490);
xnor U567 (N_567,In_2701,In_2492);
nor U568 (N_568,In_835,In_503);
xor U569 (N_569,In_1769,In_1968);
or U570 (N_570,In_2049,In_2044);
and U571 (N_571,In_63,In_2289);
xnor U572 (N_572,In_537,In_2962);
nand U573 (N_573,In_1845,In_1804);
nand U574 (N_574,In_2702,In_415);
or U575 (N_575,In_1141,In_539);
and U576 (N_576,In_2012,In_60);
and U577 (N_577,In_1727,In_2607);
and U578 (N_578,In_1656,In_928);
nand U579 (N_579,In_2598,In_2298);
or U580 (N_580,In_2888,In_1304);
nand U581 (N_581,In_2222,In_148);
and U582 (N_582,In_198,In_177);
or U583 (N_583,In_2395,In_2032);
or U584 (N_584,In_1991,In_2400);
or U585 (N_585,In_2696,In_863);
xnor U586 (N_586,In_178,In_2626);
nor U587 (N_587,In_2061,In_996);
nor U588 (N_588,In_1887,In_1603);
or U589 (N_589,In_242,In_1800);
or U590 (N_590,In_1433,In_2228);
nand U591 (N_591,In_1190,In_327);
and U592 (N_592,In_3,In_332);
or U593 (N_593,In_1924,In_2398);
nor U594 (N_594,In_1098,In_560);
nor U595 (N_595,In_1617,In_1673);
xnor U596 (N_596,In_2583,In_1173);
nand U597 (N_597,In_1587,In_211);
and U598 (N_598,In_95,In_5);
nor U599 (N_599,In_263,In_444);
and U600 (N_600,In_2750,In_1630);
nand U601 (N_601,In_1454,In_1700);
and U602 (N_602,In_1915,In_1655);
xnor U603 (N_603,In_2124,In_2214);
nor U604 (N_604,In_2725,In_2229);
and U605 (N_605,In_220,In_1051);
nor U606 (N_606,In_471,In_2958);
nand U607 (N_607,In_882,In_1523);
or U608 (N_608,In_1608,In_2770);
nand U609 (N_609,In_2840,In_2807);
or U610 (N_610,In_2581,In_1666);
nand U611 (N_611,In_2341,In_2011);
nand U612 (N_612,In_664,In_1192);
or U613 (N_613,In_156,In_2993);
nand U614 (N_614,In_2055,In_1096);
and U615 (N_615,In_1482,In_973);
nand U616 (N_616,In_2084,In_2241);
and U617 (N_617,In_939,In_526);
nor U618 (N_618,In_2508,In_282);
and U619 (N_619,In_687,In_401);
nor U620 (N_620,In_1260,In_521);
nor U621 (N_621,In_2634,In_237);
or U622 (N_622,In_656,In_2350);
and U623 (N_623,In_1235,In_2812);
or U624 (N_624,In_2293,In_2455);
or U625 (N_625,In_2331,In_622);
nand U626 (N_626,In_635,In_1088);
nand U627 (N_627,In_73,In_1512);
or U628 (N_628,In_458,In_2337);
nor U629 (N_629,In_2409,In_1786);
nor U630 (N_630,In_571,In_2934);
or U631 (N_631,In_2502,In_1554);
and U632 (N_632,In_954,In_508);
nor U633 (N_633,In_2330,In_966);
nand U634 (N_634,In_1041,In_1112);
nand U635 (N_635,In_1270,In_2325);
xnor U636 (N_636,In_925,In_90);
or U637 (N_637,In_2052,In_1740);
or U638 (N_638,In_704,In_2842);
or U639 (N_639,In_208,In_53);
xor U640 (N_640,In_1125,In_1037);
xor U641 (N_641,In_1836,In_1015);
nor U642 (N_642,In_2433,In_1536);
xnor U643 (N_643,In_230,In_2531);
nor U644 (N_644,In_449,In_864);
or U645 (N_645,In_597,In_41);
nand U646 (N_646,In_1515,In_549);
nor U647 (N_647,In_1867,In_2516);
nor U648 (N_648,In_757,In_858);
nand U649 (N_649,In_2728,In_1148);
nand U650 (N_650,In_112,In_2716);
and U651 (N_651,In_2859,In_1149);
nor U652 (N_652,In_2831,In_2108);
xor U653 (N_653,In_810,In_1691);
nand U654 (N_654,In_419,In_2430);
and U655 (N_655,In_1596,In_2945);
nand U656 (N_656,In_2309,In_2744);
or U657 (N_657,In_1456,In_2766);
or U658 (N_658,In_2994,In_2887);
or U659 (N_659,In_2543,In_1474);
nor U660 (N_660,In_1498,In_404);
and U661 (N_661,In_435,In_2154);
nor U662 (N_662,In_1737,In_2873);
nor U663 (N_663,In_2173,In_611);
and U664 (N_664,In_894,In_1400);
nor U665 (N_665,In_2086,In_816);
nand U666 (N_666,In_1520,In_253);
nand U667 (N_667,In_740,In_1342);
or U668 (N_668,In_88,In_1938);
nand U669 (N_669,In_2628,In_1209);
and U670 (N_670,In_1718,In_1001);
nor U671 (N_671,In_1154,In_1132);
or U672 (N_672,In_2890,In_408);
and U673 (N_673,In_2657,In_2761);
nor U674 (N_674,In_1701,In_1969);
nor U675 (N_675,In_1878,In_2624);
xor U676 (N_676,In_1468,In_174);
and U677 (N_677,In_885,In_344);
nor U678 (N_678,In_1310,In_2635);
nor U679 (N_679,In_1184,In_1470);
nor U680 (N_680,In_1509,In_2967);
or U681 (N_681,In_368,In_555);
nor U682 (N_682,In_2429,In_374);
or U683 (N_683,In_1491,In_2082);
nand U684 (N_684,In_1888,In_1384);
nand U685 (N_685,In_1820,In_660);
and U686 (N_686,In_352,In_2073);
nor U687 (N_687,In_818,In_115);
and U688 (N_688,In_551,In_2780);
and U689 (N_689,In_243,In_933);
nand U690 (N_690,In_1054,In_2263);
nand U691 (N_691,In_2630,In_2565);
nor U692 (N_692,In_983,In_2373);
and U693 (N_693,In_2526,In_514);
or U694 (N_694,In_2674,In_845);
nand U695 (N_695,In_1165,In_1668);
nor U696 (N_696,In_111,In_2356);
nor U697 (N_697,In_1360,In_1731);
nand U698 (N_698,In_964,In_2414);
and U699 (N_699,In_737,In_1378);
nor U700 (N_700,In_665,In_616);
and U701 (N_701,In_701,In_1115);
xnor U702 (N_702,In_2729,In_258);
and U703 (N_703,In_495,In_683);
or U704 (N_704,In_141,In_1025);
or U705 (N_705,In_1007,In_1896);
or U706 (N_706,In_2551,In_1410);
and U707 (N_707,In_2481,In_959);
or U708 (N_708,In_1760,In_275);
nand U709 (N_709,In_1431,In_2242);
nand U710 (N_710,In_2483,In_1490);
nand U711 (N_711,In_655,In_900);
nand U712 (N_712,In_2584,In_418);
and U713 (N_713,In_2047,In_1161);
and U714 (N_714,In_1638,In_2141);
nand U715 (N_715,In_2708,In_2410);
and U716 (N_716,In_808,In_2307);
or U717 (N_717,In_267,In_430);
xor U718 (N_718,In_1654,In_1885);
and U719 (N_719,In_290,In_333);
nor U720 (N_720,In_2051,In_2940);
nor U721 (N_721,In_671,In_891);
and U722 (N_722,In_2128,In_1579);
nand U723 (N_723,In_1771,In_1909);
nor U724 (N_724,In_2644,In_2060);
nand U725 (N_725,In_1200,In_2401);
and U726 (N_726,In_1441,In_224);
and U727 (N_727,In_1773,In_462);
nor U728 (N_728,In_715,In_2406);
or U729 (N_729,In_590,In_2722);
nand U730 (N_730,In_59,In_1949);
or U731 (N_731,In_61,In_1801);
and U732 (N_732,In_601,In_353);
nor U733 (N_733,In_974,In_2187);
and U734 (N_734,In_1898,In_318);
nor U735 (N_735,In_2666,In_481);
nand U736 (N_736,In_921,In_1636);
nand U737 (N_737,In_1448,In_2296);
xnor U738 (N_738,In_142,In_2466);
or U739 (N_739,In_691,In_586);
nor U740 (N_740,In_1556,In_1341);
nand U741 (N_741,In_191,In_1766);
nor U742 (N_742,In_1380,In_336);
nor U743 (N_743,In_2596,In_2640);
nor U744 (N_744,In_1344,In_760);
or U745 (N_745,In_2143,In_971);
nor U746 (N_746,In_1984,In_9);
nand U747 (N_747,In_1129,In_2605);
or U748 (N_748,In_1568,In_2379);
nor U749 (N_749,In_2148,In_1068);
nor U750 (N_750,In_15,In_2966);
nand U751 (N_751,In_274,In_1176);
nand U752 (N_752,In_2660,In_2489);
and U753 (N_753,In_1157,In_2370);
and U754 (N_754,In_400,In_1912);
nor U755 (N_755,In_613,In_1922);
nor U756 (N_756,In_1455,In_1933);
nor U757 (N_757,In_1776,In_467);
or U758 (N_758,In_689,In_793);
or U759 (N_759,In_447,In_1108);
nand U760 (N_760,In_204,In_578);
nand U761 (N_761,In_2130,In_837);
and U762 (N_762,In_1583,In_2457);
xor U763 (N_763,In_2920,In_1601);
or U764 (N_764,In_6,In_2436);
nand U765 (N_765,In_594,In_2200);
or U766 (N_766,In_129,In_144);
nor U767 (N_767,In_1476,In_1899);
nor U768 (N_768,In_2881,In_2899);
nor U769 (N_769,In_235,In_119);
nand U770 (N_770,In_2700,In_382);
nand U771 (N_771,In_1444,In_2979);
nor U772 (N_772,In_1626,In_1780);
nand U773 (N_773,In_982,In_1023);
nor U774 (N_774,In_272,In_1687);
nand U775 (N_775,In_678,In_1238);
and U776 (N_776,In_1367,In_978);
xnor U777 (N_777,In_1462,In_2258);
xnor U778 (N_778,In_1519,In_721);
and U779 (N_779,In_1067,In_2808);
nand U780 (N_780,In_213,In_373);
or U781 (N_781,In_2745,In_7);
or U782 (N_782,In_52,In_492);
nand U783 (N_783,In_2453,In_285);
or U784 (N_784,In_1008,In_1764);
nor U785 (N_785,In_1276,In_1343);
nor U786 (N_786,In_1408,In_2690);
nand U787 (N_787,In_377,In_1751);
nor U788 (N_788,In_1499,In_1187);
nor U789 (N_789,In_2892,In_1321);
nor U790 (N_790,In_1311,In_1179);
nor U791 (N_791,In_1965,In_1228);
nand U792 (N_792,In_288,In_2806);
nor U793 (N_793,In_745,In_1627);
nor U794 (N_794,In_2392,In_827);
nand U795 (N_795,In_1226,In_2753);
nand U796 (N_796,In_564,In_325);
xor U797 (N_797,In_1000,In_2820);
nor U798 (N_798,In_499,In_1978);
and U799 (N_799,In_676,In_2480);
and U800 (N_800,In_2792,In_126);
or U801 (N_801,In_2642,In_1830);
or U802 (N_802,In_2580,In_1217);
nand U803 (N_803,In_2541,In_1624);
nor U804 (N_804,In_2357,In_1652);
or U805 (N_805,In_2759,In_993);
and U806 (N_806,In_2039,In_459);
or U807 (N_807,In_785,In_1704);
or U808 (N_808,In_79,In_255);
or U809 (N_809,In_2870,In_738);
and U810 (N_810,In_1119,In_2747);
nor U811 (N_811,In_1428,In_1640);
nor U812 (N_812,In_2656,In_803);
xnor U813 (N_813,In_1459,In_708);
nor U814 (N_814,In_582,In_2520);
nand U815 (N_815,In_2562,In_2140);
nor U816 (N_816,In_1661,In_1539);
or U817 (N_817,In_2031,In_84);
and U818 (N_818,In_74,In_917);
or U819 (N_819,In_2557,In_869);
or U820 (N_820,In_2614,In_301);
and U821 (N_821,In_488,In_1066);
nor U822 (N_822,In_1902,In_1398);
nor U823 (N_823,In_1319,In_123);
nor U824 (N_824,In_2292,In_962);
and U825 (N_825,In_1880,In_2169);
nand U826 (N_826,In_2695,In_1278);
or U827 (N_827,In_2823,In_1285);
nand U828 (N_828,In_761,In_308);
or U829 (N_829,In_1787,In_2546);
or U830 (N_830,In_153,In_210);
or U831 (N_831,In_1696,In_2809);
nor U832 (N_832,In_1931,In_1835);
nor U833 (N_833,In_2484,In_2814);
nor U834 (N_834,In_2022,In_2950);
nand U835 (N_835,In_1202,In_2033);
and U836 (N_836,In_801,In_307);
and U837 (N_837,In_1426,In_792);
nor U838 (N_838,In_2601,In_1080);
xnor U839 (N_839,In_389,In_2123);
nand U840 (N_840,In_1982,In_705);
xnor U841 (N_841,In_351,In_724);
nand U842 (N_842,In_491,In_2691);
nand U843 (N_843,In_2246,In_414);
and U844 (N_844,In_1251,In_2563);
and U845 (N_845,In_697,In_1102);
and U846 (N_846,In_163,In_326);
xor U847 (N_847,In_702,In_2540);
nor U848 (N_848,In_1423,In_1648);
and U849 (N_849,In_682,In_2168);
nor U850 (N_850,In_716,In_305);
or U851 (N_851,In_1839,In_2250);
nor U852 (N_852,In_707,In_436);
xor U853 (N_853,In_1352,In_342);
nand U854 (N_854,In_1354,In_323);
or U855 (N_855,In_1531,In_1453);
or U856 (N_856,In_19,In_841);
or U857 (N_857,In_2482,In_2535);
nand U858 (N_858,In_2335,In_98);
and U859 (N_859,In_893,In_2121);
nor U860 (N_860,In_1403,In_2682);
xnor U861 (N_861,In_903,In_1331);
and U862 (N_862,In_2768,In_239);
nor U863 (N_863,In_2318,In_1562);
or U864 (N_864,In_1871,In_2471);
and U865 (N_865,In_2461,In_631);
nor U866 (N_866,In_2384,In_2501);
nor U867 (N_867,In_1223,In_2180);
or U868 (N_868,In_2553,In_1405);
nor U869 (N_869,In_1336,In_787);
and U870 (N_870,In_1168,In_797);
nand U871 (N_871,In_80,In_380);
or U872 (N_872,In_2997,In_1709);
nor U873 (N_873,In_1307,In_2172);
and U874 (N_874,In_2717,In_548);
nor U875 (N_875,In_968,In_1079);
nor U876 (N_876,In_2895,In_1992);
nand U877 (N_877,In_13,In_8);
and U878 (N_878,In_520,In_2555);
or U879 (N_879,In_2300,In_1052);
nand U880 (N_880,In_16,In_796);
nand U881 (N_881,In_2288,In_1299);
or U882 (N_882,In_1999,In_207);
nor U883 (N_883,In_679,In_1022);
nand U884 (N_884,In_2463,In_2216);
nand U885 (N_885,In_2542,In_1283);
xnor U886 (N_886,In_2875,In_1712);
nand U887 (N_887,In_2602,In_1834);
nor U888 (N_888,In_341,In_1039);
nor U889 (N_889,In_1905,In_690);
or U890 (N_890,In_1947,In_2784);
nand U891 (N_891,In_1784,In_2184);
nor U892 (N_892,In_2785,In_43);
and U893 (N_893,In_1193,In_1114);
and U894 (N_894,In_649,In_2278);
and U895 (N_895,In_2521,In_658);
xnor U896 (N_896,In_2268,In_703);
nand U897 (N_897,In_947,In_50);
and U898 (N_898,In_1242,In_2765);
or U899 (N_899,In_1452,In_2110);
nor U900 (N_900,In_758,In_152);
or U901 (N_901,In_1044,In_1056);
and U902 (N_902,In_2845,In_2503);
and U903 (N_903,In_1689,In_26);
nand U904 (N_904,In_2196,In_1191);
or U905 (N_905,In_1463,In_2740);
nor U906 (N_906,In_1548,In_2922);
nor U907 (N_907,In_2422,In_196);
or U908 (N_908,In_425,In_2877);
and U909 (N_909,In_668,In_1464);
xnor U910 (N_910,In_410,In_2549);
nor U911 (N_911,In_865,In_2174);
xnor U912 (N_912,In_2703,In_104);
or U913 (N_913,In_2604,In_1763);
nand U914 (N_914,In_822,In_1308);
nor U915 (N_915,In_1785,In_1986);
nor U916 (N_916,In_2590,In_1493);
or U917 (N_917,In_91,In_2175);
xor U918 (N_918,In_2001,In_1678);
and U919 (N_919,In_1249,In_1809);
nor U920 (N_920,In_228,In_599);
and U921 (N_921,In_339,In_1292);
nand U922 (N_922,In_2512,In_1394);
nand U923 (N_923,In_2670,In_2190);
nor U924 (N_924,In_158,In_2775);
nor U925 (N_925,In_1710,In_2924);
nor U926 (N_926,In_183,In_375);
or U927 (N_927,In_2649,In_934);
nand U928 (N_928,In_1948,In_429);
nor U929 (N_929,In_952,In_2301);
and U930 (N_930,In_1399,In_1077);
nor U931 (N_931,In_591,In_1910);
nand U932 (N_932,In_490,In_2459);
nor U933 (N_933,In_1026,In_1698);
nand U934 (N_934,In_2431,In_2456);
or U935 (N_935,In_1634,In_264);
nand U936 (N_936,In_1842,In_246);
nand U937 (N_937,In_18,In_2391);
and U938 (N_938,In_1599,In_1370);
or U939 (N_939,In_0,In_2142);
nand U940 (N_940,In_969,In_2164);
and U941 (N_941,In_1662,In_2323);
and U942 (N_942,In_2145,In_2971);
or U943 (N_943,In_1348,In_193);
or U944 (N_944,In_1891,In_651);
nand U945 (N_945,In_1401,In_825);
and U946 (N_946,In_2093,In_2539);
or U947 (N_947,In_2947,In_1874);
or U948 (N_948,In_1028,In_2858);
nand U949 (N_949,In_1158,In_904);
nor U950 (N_950,In_848,In_2440);
or U951 (N_951,In_1286,In_2230);
or U952 (N_952,In_2226,In_1790);
nor U953 (N_953,In_473,In_2252);
nor U954 (N_954,In_171,In_1609);
nand U955 (N_955,In_2904,In_1686);
nor U956 (N_956,In_795,In_814);
and U957 (N_957,In_2514,In_1816);
nor U958 (N_958,In_714,In_87);
nand U959 (N_959,In_1946,In_1432);
or U960 (N_960,In_2537,In_937);
nand U961 (N_961,In_1802,In_2305);
nor U962 (N_962,In_85,In_1963);
nand U963 (N_963,In_659,In_723);
or U964 (N_964,In_407,In_2063);
and U965 (N_965,In_850,In_914);
and U966 (N_966,In_566,In_940);
or U967 (N_967,In_484,In_1045);
and U968 (N_968,In_296,In_944);
or U969 (N_969,In_434,In_2183);
xor U970 (N_970,In_1777,In_2107);
nand U971 (N_971,In_855,In_1256);
xnor U972 (N_972,In_2758,In_1578);
xor U973 (N_973,In_1544,In_2789);
or U974 (N_974,In_2865,In_1812);
nand U975 (N_975,In_445,In_2464);
or U976 (N_976,In_1797,In_1178);
xnor U977 (N_977,In_1733,In_254);
nor U978 (N_978,In_1657,In_402);
nand U979 (N_979,In_980,In_1357);
nand U980 (N_980,In_2853,In_184);
or U981 (N_981,In_1542,In_2868);
nor U982 (N_982,In_2265,In_574);
nor U983 (N_983,In_1147,In_2314);
nor U984 (N_984,In_1273,In_1094);
nor U985 (N_985,In_1747,In_2684);
and U986 (N_986,In_621,In_2941);
nand U987 (N_987,In_1280,In_151);
or U988 (N_988,In_2469,In_1904);
nand U989 (N_989,In_580,In_2787);
or U990 (N_990,In_2251,In_1075);
and U991 (N_991,In_2076,In_1122);
and U992 (N_992,In_674,In_2673);
nand U993 (N_993,In_2930,In_1362);
nand U994 (N_994,In_472,In_1442);
nor U995 (N_995,In_1988,In_2249);
and U996 (N_996,In_2359,In_1651);
and U997 (N_997,In_2040,In_2448);
and U998 (N_998,In_361,In_2345);
nand U999 (N_999,In_806,In_812);
or U1000 (N_1000,In_2376,In_2615);
nand U1001 (N_1001,In_1050,In_1263);
or U1002 (N_1002,In_1964,In_1598);
or U1003 (N_1003,In_1644,In_2939);
and U1004 (N_1004,In_2498,In_2748);
and U1005 (N_1005,In_2078,In_1772);
nor U1006 (N_1006,In_749,In_1297);
nor U1007 (N_1007,In_2839,In_2606);
nor U1008 (N_1008,In_919,In_314);
nor U1009 (N_1009,In_2454,In_454);
xnor U1010 (N_1010,In_752,In_1920);
nor U1011 (N_1011,In_1543,In_37);
and U1012 (N_1012,In_2344,In_2114);
or U1013 (N_1013,In_2560,In_2648);
nor U1014 (N_1014,In_1169,In_2738);
nor U1015 (N_1015,In_1225,In_2739);
and U1016 (N_1016,In_1607,In_1510);
nor U1017 (N_1017,In_2146,In_2530);
or U1018 (N_1018,In_1372,In_1625);
and U1019 (N_1019,In_94,In_1792);
or U1020 (N_1020,In_2566,In_1653);
and U1021 (N_1021,In_2115,In_2233);
xnor U1022 (N_1022,In_2917,In_2592);
and U1023 (N_1023,In_2267,In_482);
and U1024 (N_1024,In_2830,In_1502);
or U1025 (N_1025,In_2972,In_1945);
nor U1026 (N_1026,In_124,In_2245);
and U1027 (N_1027,In_1116,In_1959);
nand U1028 (N_1028,In_790,In_2907);
nor U1029 (N_1029,In_842,In_2954);
nand U1030 (N_1030,In_1287,In_1477);
and U1031 (N_1031,In_2704,In_1851);
or U1032 (N_1032,In_298,In_214);
xnor U1033 (N_1033,In_127,In_2752);
and U1034 (N_1034,In_2023,In_726);
and U1035 (N_1035,In_1445,In_287);
or U1036 (N_1036,In_1472,In_189);
nor U1037 (N_1037,In_1537,In_1540);
nor U1038 (N_1038,In_1549,In_199);
and U1039 (N_1039,In_1189,In_617);
nand U1040 (N_1040,In_2306,In_2960);
and U1041 (N_1041,In_1411,In_661);
and U1042 (N_1042,In_764,In_209);
nand U1043 (N_1043,In_2585,In_1314);
nor U1044 (N_1044,In_2006,In_935);
and U1045 (N_1045,In_2235,In_1334);
nand U1046 (N_1046,In_317,In_2014);
xnor U1047 (N_1047,In_99,In_1002);
and U1048 (N_1048,In_2387,In_2533);
nor U1049 (N_1049,In_2046,In_587);
nor U1050 (N_1050,In_1447,In_1437);
and U1051 (N_1051,In_2677,In_2928);
or U1052 (N_1052,In_1305,In_2570);
or U1053 (N_1053,In_262,In_2303);
or U1054 (N_1054,In_110,In_2998);
or U1055 (N_1055,In_681,In_1594);
nand U1056 (N_1056,In_2714,In_100);
nor U1057 (N_1057,In_297,In_397);
xor U1058 (N_1058,In_241,In_311);
xnor U1059 (N_1059,In_1713,In_299);
or U1060 (N_1060,In_76,In_2893);
nor U1061 (N_1061,In_36,In_280);
nor U1062 (N_1062,In_2178,In_2989);
nor U1063 (N_1063,In_1099,In_1207);
nand U1064 (N_1064,In_2912,In_2026);
and U1065 (N_1065,In_1610,In_1101);
or U1066 (N_1066,In_476,In_2007);
nand U1067 (N_1067,In_2884,In_1789);
or U1068 (N_1068,In_746,In_2778);
or U1069 (N_1069,In_182,In_505);
or U1070 (N_1070,In_2273,In_2742);
or U1071 (N_1071,In_2741,In_2667);
and U1072 (N_1072,In_2732,In_1856);
nand U1073 (N_1073,In_1254,In_1210);
nand U1074 (N_1074,In_225,In_902);
and U1075 (N_1075,In_1072,In_498);
nand U1076 (N_1076,In_2547,In_813);
and U1077 (N_1077,In_777,In_200);
or U1078 (N_1078,In_2386,In_2977);
or U1079 (N_1079,In_2848,In_1622);
nor U1080 (N_1080,In_2438,In_1997);
and U1081 (N_1081,In_1128,In_1152);
or U1082 (N_1082,In_901,In_331);
nand U1083 (N_1083,In_614,In_370);
or U1084 (N_1084,In_2170,In_619);
and U1085 (N_1085,In_1246,In_2340);
xor U1086 (N_1086,In_2362,In_2435);
and U1087 (N_1087,In_2294,In_493);
nor U1088 (N_1088,In_30,In_2150);
and U1089 (N_1089,In_1504,In_2);
and U1090 (N_1090,In_107,In_33);
and U1091 (N_1091,In_2360,In_2317);
and U1092 (N_1092,In_2710,In_2316);
and U1093 (N_1093,In_2909,In_2072);
or U1094 (N_1094,In_907,In_1577);
nand U1095 (N_1095,In_2004,In_2403);
or U1096 (N_1096,In_1230,In_2036);
and U1097 (N_1097,In_2407,In_1875);
xor U1098 (N_1098,In_593,In_2970);
and U1099 (N_1099,In_700,In_1317);
and U1100 (N_1100,In_1186,In_25);
nor U1101 (N_1101,In_1937,In_1697);
and U1102 (N_1102,In_2913,In_2515);
or U1103 (N_1103,In_2439,In_1863);
or U1104 (N_1104,In_1975,In_1647);
nor U1105 (N_1105,In_71,In_1870);
or U1106 (N_1106,In_636,In_2882);
or U1107 (N_1107,In_1641,In_256);
nor U1108 (N_1108,In_365,In_1076);
or U1109 (N_1109,In_1674,In_2067);
or U1110 (N_1110,In_1882,In_103);
or U1111 (N_1111,In_1869,In_1681);
or U1112 (N_1112,In_1742,In_1914);
or U1113 (N_1113,In_165,In_2441);
or U1114 (N_1114,In_831,In_1857);
and U1115 (N_1115,In_2957,In_2600);
or U1116 (N_1116,In_277,In_483);
or U1117 (N_1117,In_2802,In_2627);
or U1118 (N_1118,In_356,In_1943);
nand U1119 (N_1119,In_729,In_21);
nand U1120 (N_1120,In_2629,In_2116);
nor U1121 (N_1121,In_2332,In_1592);
or U1122 (N_1122,In_2208,In_1412);
nand U1123 (N_1123,In_528,In_2579);
and U1124 (N_1124,In_2203,In_1328);
or U1125 (N_1125,In_2991,In_2984);
nor U1126 (N_1126,In_2452,In_995);
or U1127 (N_1127,In_1303,In_197);
or U1128 (N_1128,In_2260,In_2861);
and U1129 (N_1129,In_2259,In_2397);
or U1130 (N_1130,In_2427,In_873);
and U1131 (N_1131,In_51,In_1953);
or U1132 (N_1132,In_2002,In_625);
nor U1133 (N_1133,In_2308,In_1266);
nor U1134 (N_1134,In_532,In_1419);
nand U1135 (N_1135,In_291,In_2041);
or U1136 (N_1136,In_2534,In_2561);
or U1137 (N_1137,In_1487,In_1496);
nand U1138 (N_1138,In_2914,In_876);
nand U1139 (N_1139,In_1326,In_114);
and U1140 (N_1140,In_1371,In_1284);
or U1141 (N_1141,In_194,In_2349);
or U1142 (N_1142,In_1884,In_1858);
or U1143 (N_1143,In_1628,In_589);
nand U1144 (N_1144,In_1081,In_663);
and U1145 (N_1145,In_1012,In_2623);
and U1146 (N_1146,In_563,In_433);
nor U1147 (N_1147,In_2676,In_535);
and U1148 (N_1148,In_227,In_2679);
nor U1149 (N_1149,In_2257,In_711);
nand U1150 (N_1150,In_1268,In_1788);
nor U1151 (N_1151,In_1171,In_1714);
or U1152 (N_1152,In_1929,In_2699);
and U1153 (N_1153,In_805,In_898);
or U1154 (N_1154,In_2351,In_1643);
and U1155 (N_1155,In_2838,In_963);
or U1156 (N_1156,In_172,In_1614);
xnor U1157 (N_1157,In_81,In_206);
nand U1158 (N_1158,In_1576,In_2641);
and U1159 (N_1159,In_300,In_2013);
nor U1160 (N_1160,In_1546,In_633);
nor U1161 (N_1161,In_1040,In_562);
or U1162 (N_1162,In_2087,In_2900);
nor U1163 (N_1163,In_1224,In_2077);
or U1164 (N_1164,In_1391,In_2576);
nand U1165 (N_1165,In_181,In_755);
or U1166 (N_1166,In_1877,In_1247);
and U1167 (N_1167,In_2943,In_328);
or U1168 (N_1168,In_1315,In_1048);
or U1169 (N_1169,In_2856,In_672);
nand U1170 (N_1170,In_782,In_1768);
nand U1171 (N_1171,In_494,In_1138);
nor U1172 (N_1172,In_2968,In_2921);
or U1173 (N_1173,In_638,In_1732);
nand U1174 (N_1174,In_2777,In_880);
or U1175 (N_1175,In_2949,In_420);
and U1176 (N_1176,In_236,In_948);
and U1177 (N_1177,In_1450,In_1073);
nor U1178 (N_1178,In_778,In_2109);
nand U1179 (N_1179,In_2075,In_2254);
or U1180 (N_1180,In_2477,In_1233);
and U1181 (N_1181,In_2638,In_46);
and U1182 (N_1182,In_293,In_2731);
and U1183 (N_1183,In_496,In_2358);
nor U1184 (N_1184,In_2671,In_608);
xnor U1185 (N_1185,In_2496,In_747);
nand U1186 (N_1186,In_1677,In_2737);
nor U1187 (N_1187,In_1151,In_538);
and U1188 (N_1188,In_2053,In_859);
or U1189 (N_1189,In_2151,In_734);
nor U1190 (N_1190,In_2198,In_1571);
nor U1191 (N_1191,In_70,In_1994);
or U1192 (N_1192,In_833,In_387);
and U1193 (N_1193,In_2799,In_596);
nand U1194 (N_1194,In_1961,In_338);
or U1195 (N_1195,In_2931,In_1866);
nor U1196 (N_1196,In_1327,In_2567);
and U1197 (N_1197,In_2302,In_2343);
xor U1198 (N_1198,In_2213,In_2878);
or U1199 (N_1199,In_774,In_800);
and U1200 (N_1200,In_1279,In_2869);
and U1201 (N_1201,In_2755,In_2652);
and U1202 (N_1202,In_2980,In_1042);
and U1203 (N_1203,In_943,In_623);
nand U1204 (N_1204,In_1817,In_1895);
and U1205 (N_1205,In_804,In_998);
xor U1206 (N_1206,In_2713,In_168);
or U1207 (N_1207,In_1629,In_1014);
nor U1208 (N_1208,In_12,In_1375);
and U1209 (N_1209,In_486,In_986);
nand U1210 (N_1210,In_1306,In_2591);
nor U1211 (N_1211,In_1142,In_1092);
nand U1212 (N_1212,In_2262,In_618);
and U1213 (N_1213,In_2655,In_2730);
nand U1214 (N_1214,In_941,In_1765);
or U1215 (N_1215,In_489,In_654);
or U1216 (N_1216,In_965,In_889);
nor U1217 (N_1217,In_544,In_238);
xor U1218 (N_1218,In_2271,In_324);
and U1219 (N_1219,In_1180,In_504);
nor U1220 (N_1220,In_54,In_2763);
nor U1221 (N_1221,In_918,In_249);
or U1222 (N_1222,In_2518,In_2836);
nand U1223 (N_1223,In_1723,In_1868);
nand U1224 (N_1224,In_2102,In_2297);
nand U1225 (N_1225,In_2129,In_2936);
nand U1226 (N_1226,In_1778,In_1214);
nor U1227 (N_1227,In_915,In_2234);
nor U1228 (N_1228,In_2098,In_1082);
xor U1229 (N_1229,In_1570,In_216);
and U1230 (N_1230,In_1123,In_2034);
nand U1231 (N_1231,In_942,In_2008);
nand U1232 (N_1232,In_720,In_1064);
or U1233 (N_1233,In_4,In_2354);
and U1234 (N_1234,In_2595,In_2662);
nand U1235 (N_1235,In_1393,In_1495);
nor U1236 (N_1236,In_1005,In_188);
nand U1237 (N_1237,In_552,In_1995);
nor U1238 (N_1238,In_1027,In_1004);
or U1239 (N_1239,In_2879,In_1722);
nor U1240 (N_1240,In_1927,In_2661);
nand U1241 (N_1241,In_2167,In_2101);
nand U1242 (N_1242,In_140,In_2402);
nor U1243 (N_1243,In_1775,In_487);
xnor U1244 (N_1244,In_1828,In_34);
and U1245 (N_1245,In_1245,In_2545);
nand U1246 (N_1246,In_65,In_735);
nand U1247 (N_1247,In_1160,In_250);
or U1248 (N_1248,In_2749,In_2837);
nand U1249 (N_1249,In_17,In_1633);
nor U1250 (N_1250,In_281,In_767);
and U1251 (N_1251,In_1893,In_890);
nor U1252 (N_1252,In_1150,In_1421);
or U1253 (N_1253,In_2797,In_2355);
nor U1254 (N_1254,In_2460,In_1290);
xnor U1255 (N_1255,In_2774,In_861);
nor U1256 (N_1256,In_399,In_1124);
and U1257 (N_1257,In_2771,In_390);
and U1258 (N_1258,In_1726,In_1240);
nand U1259 (N_1259,In_348,In_109);
xor U1260 (N_1260,In_240,In_1782);
nor U1261 (N_1261,In_967,In_1185);
or U1262 (N_1262,In_2511,In_1134);
xnor U1263 (N_1263,In_1181,In_2473);
or U1264 (N_1264,In_1521,In_2860);
xor U1265 (N_1265,In_2880,In_1145);
xor U1266 (N_1266,In_519,In_2664);
nand U1267 (N_1267,In_1300,In_592);
or U1268 (N_1268,In_1492,In_2720);
nand U1269 (N_1269,In_1873,In_2045);
and U1270 (N_1270,In_709,In_565);
nand U1271 (N_1271,In_568,In_1275);
nand U1272 (N_1272,In_1069,In_1111);
nor U1273 (N_1273,In_1312,In_2381);
and U1274 (N_1274,In_604,In_2646);
nand U1275 (N_1275,In_2938,In_2803);
and U1276 (N_1276,In_1346,In_913);
xor U1277 (N_1277,In_1397,In_2270);
nor U1278 (N_1278,In_906,In_271);
nor U1279 (N_1279,In_1322,In_2284);
or U1280 (N_1280,In_108,In_518);
nand U1281 (N_1281,In_1031,In_451);
and U1282 (N_1282,In_839,In_1071);
nor U1283 (N_1283,In_2651,In_2194);
nand U1284 (N_1284,In_1436,In_1534);
or U1285 (N_1285,In_1752,In_357);
nand U1286 (N_1286,In_1024,In_1271);
nand U1287 (N_1287,In_546,In_295);
nand U1288 (N_1288,In_2295,In_2411);
and U1289 (N_1289,In_2310,In_2009);
nor U1290 (N_1290,In_2156,In_2189);
nand U1291 (N_1291,In_1376,In_1672);
xnor U1292 (N_1292,In_1467,In_2209);
nand U1293 (N_1293,In_1917,In_2981);
and U1294 (N_1294,In_2834,In_2835);
nor U1295 (N_1295,In_2113,In_2028);
xnor U1296 (N_1296,In_24,In_1481);
nand U1297 (N_1297,In_1429,In_1615);
nand U1298 (N_1298,In_924,In_2276);
nor U1299 (N_1299,In_2857,In_2353);
xnor U1300 (N_1300,In_1954,In_2450);
or U1301 (N_1301,In_731,In_1513);
and U1302 (N_1302,In_2519,In_1195);
nand U1303 (N_1303,In_851,In_2705);
nor U1304 (N_1304,In_1806,In_2529);
nor U1305 (N_1305,In_1658,In_2517);
nand U1306 (N_1306,In_1831,In_456);
or U1307 (N_1307,In_1133,In_2348);
or U1308 (N_1308,In_641,In_1908);
nand U1309 (N_1309,In_1813,In_1379);
or U1310 (N_1310,In_2383,In_405);
or U1311 (N_1311,In_1551,In_680);
or U1312 (N_1312,In_2468,In_2197);
or U1313 (N_1313,In_2185,In_1349);
nand U1314 (N_1314,In_1,In_1916);
xnor U1315 (N_1315,In_1218,In_485);
and U1316 (N_1316,In_1575,In_1618);
and U1317 (N_1317,In_2176,In_2990);
and U1318 (N_1318,In_1259,In_2978);
and U1319 (N_1319,In_524,In_1989);
and U1320 (N_1320,In_2220,In_2313);
nand U1321 (N_1321,In_1558,In_1552);
or U1322 (N_1322,In_1033,In_316);
and U1323 (N_1323,In_1272,In_2299);
and U1324 (N_1324,In_64,In_2437);
nand U1325 (N_1325,In_2290,In_2394);
and U1326 (N_1326,In_2425,In_829);
or U1327 (N_1327,In_2527,In_169);
or U1328 (N_1328,In_600,In_2139);
and U1329 (N_1329,In_1616,In_1522);
nand U1330 (N_1330,In_2894,In_2125);
and U1331 (N_1331,In_1055,In_1029);
or U1332 (N_1332,In_772,In_2424);
or U1333 (N_1333,In_823,In_201);
xnor U1334 (N_1334,In_2240,In_1645);
and U1335 (N_1335,In_2709,In_1241);
nand U1336 (N_1336,In_895,In_1683);
nor U1337 (N_1337,In_1083,In_2846);
nand U1338 (N_1338,In_2232,In_1639);
nand U1339 (N_1339,In_2015,In_1146);
nand U1340 (N_1340,In_877,In_1063);
nor U1341 (N_1341,In_2159,In_2504);
nand U1342 (N_1342,In_2647,In_1489);
nand U1343 (N_1343,In_868,In_195);
xor U1344 (N_1344,In_1739,In_699);
nand U1345 (N_1345,In_557,In_2237);
xor U1346 (N_1346,In_412,In_1338);
or U1347 (N_1347,In_1208,In_442);
xor U1348 (N_1348,In_422,In_309);
and U1349 (N_1349,In_1236,In_515);
xor U1350 (N_1350,In_2524,In_2346);
nor U1351 (N_1351,In_423,In_1156);
or U1352 (N_1352,In_1803,In_598);
or U1353 (N_1353,In_1049,In_862);
xor U1354 (N_1354,In_2800,In_2152);
and U1355 (N_1355,In_646,In_359);
xor U1356 (N_1356,In_550,In_657);
nand U1357 (N_1357,In_231,In_2347);
or U1358 (N_1358,In_1034,In_2693);
or U1359 (N_1359,In_2944,In_1894);
nor U1360 (N_1360,In_612,In_1449);
and U1361 (N_1361,In_970,In_479);
nand U1362 (N_1362,In_2255,In_2239);
and U1363 (N_1363,In_2558,In_553);
nor U1364 (N_1364,In_139,In_1547);
nand U1365 (N_1365,In_2050,In_1406);
and U1366 (N_1366,In_2048,In_2603);
nand U1367 (N_1367,In_1799,In_2326);
nand U1368 (N_1368,In_1559,In_2158);
or U1369 (N_1369,In_2487,In_460);
or U1370 (N_1370,In_2396,In_2385);
and U1371 (N_1371,In_1565,In_1667);
nor U1372 (N_1372,In_2090,In_1211);
nor U1373 (N_1373,In_1826,In_1862);
nand U1374 (N_1374,In_809,In_2616);
and U1375 (N_1375,In_1623,In_784);
or U1376 (N_1376,In_1473,In_1465);
xor U1377 (N_1377,In_1511,In_1345);
or U1378 (N_1378,In_1711,In_2891);
xnor U1379 (N_1379,In_1886,In_266);
and U1380 (N_1380,In_132,In_686);
nor U1381 (N_1381,In_1669,In_1903);
and U1382 (N_1382,In_888,In_2965);
nand U1383 (N_1383,In_730,In_1983);
nand U1384 (N_1384,In_1087,In_2219);
nor U1385 (N_1385,In_1243,In_1325);
or U1386 (N_1386,In_1032,In_2097);
or U1387 (N_1387,In_55,In_2712);
or U1388 (N_1388,In_1694,In_1204);
nand U1389 (N_1389,In_1402,In_923);
xor U1390 (N_1390,In_1118,In_1126);
nor U1391 (N_1391,In_122,In_821);
xnor U1392 (N_1392,In_653,In_302);
nor U1393 (N_1393,In_1724,In_440);
or U1394 (N_1394,In_1759,In_500);
xnor U1395 (N_1395,In_478,In_529);
or U1396 (N_1396,In_1460,In_909);
and U1397 (N_1397,In_2829,In_2633);
nand U1398 (N_1398,In_217,In_2399);
and U1399 (N_1399,In_1721,In_218);
and U1400 (N_1400,In_2772,In_2692);
nor U1401 (N_1401,In_2683,In_1413);
or U1402 (N_1402,In_2281,In_461);
nor U1403 (N_1403,In_315,In_1746);
nor U1404 (N_1404,In_949,In_203);
nand U1405 (N_1405,In_990,In_694);
and U1406 (N_1406,In_1825,In_23);
and U1407 (N_1407,In_83,In_972);
xnor U1408 (N_1408,In_1814,In_1533);
or U1409 (N_1409,In_540,In_2901);
or U1410 (N_1410,In_2871,In_750);
xor U1411 (N_1411,In_2405,In_644);
nor U1412 (N_1412,In_632,In_161);
or U1413 (N_1413,In_1293,In_2165);
nor U1414 (N_1414,In_1921,In_2275);
and U1415 (N_1415,In_2426,In_273);
or U1416 (N_1416,In_403,In_186);
nand U1417 (N_1417,In_630,In_910);
nand U1418 (N_1418,In_1849,In_1848);
or U1419 (N_1419,In_685,In_1743);
and U1420 (N_1420,In_2685,In_786);
or U1421 (N_1421,In_2475,In_610);
and U1422 (N_1422,In_2577,In_819);
or U1423 (N_1423,In_2206,In_698);
or U1424 (N_1424,In_164,In_2933);
nor U1425 (N_1425,In_1387,In_1818);
nand U1426 (N_1426,In_899,In_1265);
nand U1427 (N_1427,In_2751,In_1944);
and U1428 (N_1428,In_82,In_1960);
nand U1429 (N_1429,In_294,In_2205);
or U1430 (N_1430,In_1333,In_1952);
nor U1431 (N_1431,In_1355,In_1805);
xor U1432 (N_1432,In_2444,In_1794);
or U1433 (N_1433,In_270,In_609);
nor U1434 (N_1434,In_2035,In_1911);
or U1435 (N_1435,In_1987,In_1728);
and U1436 (N_1436,In_1693,In_1177);
xnor U1437 (N_1437,In_2361,In_2816);
and U1438 (N_1438,In_2282,In_279);
and U1439 (N_1439,In_2096,In_1566);
and U1440 (N_1440,In_997,In_1864);
and U1441 (N_1441,In_1705,In_533);
and U1442 (N_1442,In_645,In_2654);
nor U1443 (N_1443,In_751,In_849);
or U1444 (N_1444,In_1838,In_347);
nand U1445 (N_1445,In_1530,In_1918);
nand U1446 (N_1446,In_607,In_692);
nor U1447 (N_1447,In_2636,In_2554);
and U1448 (N_1448,In_556,In_2769);
and U1449 (N_1449,In_1182,In_121);
and U1450 (N_1450,In_251,In_2896);
nor U1451 (N_1451,In_421,In_1383);
or U1452 (N_1452,In_1690,In_466);
nor U1453 (N_1453,In_166,In_874);
nand U1454 (N_1454,In_1883,In_2092);
nor U1455 (N_1455,In_2215,In_1395);
nor U1456 (N_1456,In_826,In_455);
xnor U1457 (N_1457,In_1244,In_722);
nand U1458 (N_1458,In_516,In_1162);
and U1459 (N_1459,In_2488,In_2003);
nand U1460 (N_1460,In_1582,In_675);
nand U1461 (N_1461,In_1365,In_45);
or U1462 (N_1462,In_576,In_42);
and U1463 (N_1463,In_2810,In_2493);
and U1464 (N_1464,In_517,In_2680);
and U1465 (N_1465,In_1637,In_417);
and U1466 (N_1466,In_1545,In_2599);
or U1467 (N_1467,In_725,In_93);
or U1468 (N_1468,In_595,In_1756);
or U1469 (N_1469,In_2505,In_879);
nand U1470 (N_1470,In_450,In_2995);
or U1471 (N_1471,In_2153,In_2844);
or U1472 (N_1472,In_1239,In_2915);
nand U1473 (N_1473,In_1301,In_1550);
nand U1474 (N_1474,In_695,In_1316);
or U1475 (N_1475,In_2365,In_1564);
and U1476 (N_1476,In_2179,In_1466);
nor U1477 (N_1477,In_1941,In_398);
nor U1478 (N_1478,In_1901,In_1753);
or U1479 (N_1479,In_878,In_2494);
nand U1480 (N_1480,In_28,In_133);
and U1481 (N_1481,In_2238,In_1932);
and U1482 (N_1482,In_2620,In_1762);
and U1483 (N_1483,In_820,In_2658);
nand U1484 (N_1484,In_2495,In_2135);
nor U1485 (N_1485,In_2065,In_2874);
and U1486 (N_1486,In_2149,In_1664);
nor U1487 (N_1487,In_2393,In_1388);
xnor U1488 (N_1488,In_501,In_1140);
nor U1489 (N_1489,In_717,In_2491);
nor U1490 (N_1490,In_2137,In_798);
or U1491 (N_1491,In_1139,In_2911);
nand U1492 (N_1492,In_44,In_223);
xnor U1493 (N_1493,In_1925,In_2010);
or U1494 (N_1494,In_1019,In_1227);
or U1495 (N_1495,In_912,In_2919);
and U1496 (N_1496,In_1507,In_416);
nand U1497 (N_1497,In_554,In_2903);
or U1498 (N_1498,In_567,In_1167);
nor U1499 (N_1499,In_35,In_2790);
or U1500 (N_1500,In_180,In_1213);
and U1501 (N_1501,In_1242,In_1488);
or U1502 (N_1502,In_1316,In_1776);
or U1503 (N_1503,In_881,In_2518);
or U1504 (N_1504,In_2951,In_2417);
nand U1505 (N_1505,In_510,In_1532);
nand U1506 (N_1506,In_1205,In_191);
or U1507 (N_1507,In_927,In_2472);
and U1508 (N_1508,In_2433,In_2659);
and U1509 (N_1509,In_1488,In_1755);
or U1510 (N_1510,In_1513,In_165);
and U1511 (N_1511,In_1444,In_2757);
or U1512 (N_1512,In_339,In_738);
and U1513 (N_1513,In_2513,In_2160);
or U1514 (N_1514,In_2465,In_915);
or U1515 (N_1515,In_1619,In_1302);
nor U1516 (N_1516,In_1102,In_1898);
nand U1517 (N_1517,In_507,In_223);
nand U1518 (N_1518,In_816,In_2339);
or U1519 (N_1519,In_825,In_326);
nor U1520 (N_1520,In_804,In_1715);
or U1521 (N_1521,In_2843,In_895);
nor U1522 (N_1522,In_1071,In_2353);
and U1523 (N_1523,In_1392,In_533);
or U1524 (N_1524,In_2982,In_1760);
nand U1525 (N_1525,In_2869,In_456);
or U1526 (N_1526,In_576,In_1404);
nor U1527 (N_1527,In_1914,In_2268);
xnor U1528 (N_1528,In_1807,In_1396);
nand U1529 (N_1529,In_1503,In_1740);
or U1530 (N_1530,In_2638,In_319);
and U1531 (N_1531,In_1887,In_2143);
nand U1532 (N_1532,In_2299,In_2515);
xnor U1533 (N_1533,In_2294,In_1304);
nand U1534 (N_1534,In_1161,In_2954);
or U1535 (N_1535,In_1014,In_817);
nand U1536 (N_1536,In_2158,In_1428);
xnor U1537 (N_1537,In_2985,In_224);
and U1538 (N_1538,In_2950,In_2865);
and U1539 (N_1539,In_2790,In_1861);
or U1540 (N_1540,In_130,In_1908);
nand U1541 (N_1541,In_638,In_2080);
xor U1542 (N_1542,In_26,In_1322);
or U1543 (N_1543,In_1578,In_1447);
nor U1544 (N_1544,In_1391,In_563);
nand U1545 (N_1545,In_1455,In_191);
nand U1546 (N_1546,In_1606,In_1626);
nand U1547 (N_1547,In_2393,In_404);
xor U1548 (N_1548,In_2879,In_1129);
xor U1549 (N_1549,In_977,In_110);
xnor U1550 (N_1550,In_1836,In_1324);
or U1551 (N_1551,In_236,In_2623);
and U1552 (N_1552,In_2825,In_1262);
and U1553 (N_1553,In_1469,In_1310);
and U1554 (N_1554,In_1977,In_2658);
or U1555 (N_1555,In_511,In_1111);
and U1556 (N_1556,In_2161,In_2265);
nand U1557 (N_1557,In_862,In_2686);
nor U1558 (N_1558,In_1386,In_2748);
and U1559 (N_1559,In_2088,In_520);
nand U1560 (N_1560,In_479,In_2208);
nor U1561 (N_1561,In_1172,In_562);
or U1562 (N_1562,In_2962,In_2500);
and U1563 (N_1563,In_448,In_868);
nor U1564 (N_1564,In_1812,In_684);
and U1565 (N_1565,In_2124,In_2928);
nor U1566 (N_1566,In_1963,In_2197);
and U1567 (N_1567,In_17,In_1214);
nand U1568 (N_1568,In_1082,In_2930);
nor U1569 (N_1569,In_712,In_648);
and U1570 (N_1570,In_2891,In_2156);
nand U1571 (N_1571,In_153,In_213);
nand U1572 (N_1572,In_2237,In_2534);
nor U1573 (N_1573,In_736,In_274);
nor U1574 (N_1574,In_2069,In_398);
xnor U1575 (N_1575,In_22,In_2349);
nor U1576 (N_1576,In_2531,In_675);
and U1577 (N_1577,In_400,In_2680);
nand U1578 (N_1578,In_1188,In_2021);
xnor U1579 (N_1579,In_1174,In_2332);
xor U1580 (N_1580,In_1201,In_892);
and U1581 (N_1581,In_1501,In_61);
nor U1582 (N_1582,In_1522,In_1253);
or U1583 (N_1583,In_564,In_1215);
nand U1584 (N_1584,In_203,In_746);
xnor U1585 (N_1585,In_1450,In_192);
xnor U1586 (N_1586,In_1452,In_2263);
xnor U1587 (N_1587,In_99,In_2524);
and U1588 (N_1588,In_1152,In_237);
nand U1589 (N_1589,In_283,In_1843);
xnor U1590 (N_1590,In_2421,In_506);
nor U1591 (N_1591,In_365,In_2316);
or U1592 (N_1592,In_1729,In_638);
nor U1593 (N_1593,In_657,In_1741);
nor U1594 (N_1594,In_902,In_383);
and U1595 (N_1595,In_2983,In_512);
and U1596 (N_1596,In_2346,In_786);
nor U1597 (N_1597,In_2228,In_1790);
or U1598 (N_1598,In_1658,In_1404);
and U1599 (N_1599,In_2366,In_1208);
and U1600 (N_1600,In_449,In_642);
or U1601 (N_1601,In_1581,In_1407);
nor U1602 (N_1602,In_2931,In_1535);
or U1603 (N_1603,In_886,In_2776);
xor U1604 (N_1604,In_335,In_1846);
nand U1605 (N_1605,In_519,In_2957);
or U1606 (N_1606,In_1906,In_354);
and U1607 (N_1607,In_440,In_741);
or U1608 (N_1608,In_2572,In_521);
nand U1609 (N_1609,In_2606,In_1177);
nand U1610 (N_1610,In_2965,In_2340);
or U1611 (N_1611,In_457,In_2460);
or U1612 (N_1612,In_1777,In_2502);
nand U1613 (N_1613,In_1396,In_2978);
xor U1614 (N_1614,In_1651,In_632);
nand U1615 (N_1615,In_22,In_1399);
or U1616 (N_1616,In_2146,In_783);
and U1617 (N_1617,In_386,In_1062);
nor U1618 (N_1618,In_2066,In_1320);
xor U1619 (N_1619,In_611,In_1256);
and U1620 (N_1620,In_2909,In_1876);
nand U1621 (N_1621,In_1410,In_399);
nor U1622 (N_1622,In_2821,In_491);
nor U1623 (N_1623,In_1217,In_567);
or U1624 (N_1624,In_66,In_2065);
and U1625 (N_1625,In_303,In_701);
nand U1626 (N_1626,In_916,In_416);
nor U1627 (N_1627,In_1944,In_1409);
nand U1628 (N_1628,In_2858,In_853);
nor U1629 (N_1629,In_2370,In_1456);
or U1630 (N_1630,In_1587,In_2784);
nor U1631 (N_1631,In_2312,In_2049);
or U1632 (N_1632,In_1292,In_1024);
or U1633 (N_1633,In_2664,In_2488);
nor U1634 (N_1634,In_2000,In_492);
and U1635 (N_1635,In_2000,In_84);
and U1636 (N_1636,In_1904,In_341);
nor U1637 (N_1637,In_1556,In_1397);
or U1638 (N_1638,In_1308,In_2539);
or U1639 (N_1639,In_2169,In_540);
nor U1640 (N_1640,In_1669,In_1193);
and U1641 (N_1641,In_781,In_1630);
xnor U1642 (N_1642,In_302,In_124);
and U1643 (N_1643,In_2225,In_1483);
nor U1644 (N_1644,In_2414,In_1436);
and U1645 (N_1645,In_2703,In_204);
or U1646 (N_1646,In_2822,In_143);
nor U1647 (N_1647,In_269,In_572);
and U1648 (N_1648,In_913,In_1168);
xnor U1649 (N_1649,In_1332,In_1680);
nor U1650 (N_1650,In_1220,In_1079);
nor U1651 (N_1651,In_1602,In_1494);
xor U1652 (N_1652,In_1617,In_2973);
nor U1653 (N_1653,In_1650,In_1908);
nand U1654 (N_1654,In_2476,In_2583);
or U1655 (N_1655,In_2786,In_2306);
xnor U1656 (N_1656,In_1047,In_2243);
and U1657 (N_1657,In_2573,In_905);
nand U1658 (N_1658,In_829,In_1407);
and U1659 (N_1659,In_2817,In_2560);
nand U1660 (N_1660,In_2143,In_2352);
or U1661 (N_1661,In_1593,In_2745);
and U1662 (N_1662,In_809,In_1363);
nand U1663 (N_1663,In_2951,In_1285);
or U1664 (N_1664,In_1833,In_1037);
nand U1665 (N_1665,In_2177,In_612);
nand U1666 (N_1666,In_2544,In_2775);
or U1667 (N_1667,In_1620,In_610);
nor U1668 (N_1668,In_2666,In_755);
or U1669 (N_1669,In_1212,In_831);
nor U1670 (N_1670,In_502,In_196);
nand U1671 (N_1671,In_2851,In_161);
nand U1672 (N_1672,In_2307,In_2778);
nor U1673 (N_1673,In_1119,In_2924);
and U1674 (N_1674,In_2948,In_1240);
nand U1675 (N_1675,In_2441,In_369);
and U1676 (N_1676,In_1452,In_723);
nor U1677 (N_1677,In_2780,In_1892);
nand U1678 (N_1678,In_2671,In_122);
or U1679 (N_1679,In_1467,In_1787);
or U1680 (N_1680,In_2728,In_122);
nor U1681 (N_1681,In_1004,In_2027);
nor U1682 (N_1682,In_800,In_2506);
nand U1683 (N_1683,In_1522,In_808);
nor U1684 (N_1684,In_2300,In_2583);
nand U1685 (N_1685,In_2161,In_2417);
or U1686 (N_1686,In_2705,In_1817);
and U1687 (N_1687,In_647,In_2124);
and U1688 (N_1688,In_853,In_11);
and U1689 (N_1689,In_1073,In_433);
nor U1690 (N_1690,In_544,In_2050);
nand U1691 (N_1691,In_2382,In_2907);
and U1692 (N_1692,In_1176,In_983);
nand U1693 (N_1693,In_2852,In_796);
and U1694 (N_1694,In_1175,In_1041);
nand U1695 (N_1695,In_23,In_1536);
or U1696 (N_1696,In_552,In_2348);
nor U1697 (N_1697,In_220,In_448);
nand U1698 (N_1698,In_1971,In_38);
nor U1699 (N_1699,In_2098,In_1408);
or U1700 (N_1700,In_440,In_519);
and U1701 (N_1701,In_919,In_175);
nand U1702 (N_1702,In_1654,In_1377);
xor U1703 (N_1703,In_1835,In_2096);
nand U1704 (N_1704,In_2167,In_1561);
xnor U1705 (N_1705,In_2661,In_399);
and U1706 (N_1706,In_2606,In_712);
or U1707 (N_1707,In_843,In_2714);
and U1708 (N_1708,In_780,In_1281);
and U1709 (N_1709,In_1843,In_734);
nor U1710 (N_1710,In_1377,In_1153);
xor U1711 (N_1711,In_2148,In_1106);
xor U1712 (N_1712,In_765,In_2851);
nor U1713 (N_1713,In_557,In_1253);
and U1714 (N_1714,In_129,In_2071);
nor U1715 (N_1715,In_34,In_427);
nand U1716 (N_1716,In_1415,In_709);
nand U1717 (N_1717,In_2767,In_621);
nor U1718 (N_1718,In_385,In_2162);
and U1719 (N_1719,In_2495,In_774);
or U1720 (N_1720,In_1521,In_1616);
nand U1721 (N_1721,In_2347,In_2027);
and U1722 (N_1722,In_1695,In_2560);
or U1723 (N_1723,In_2745,In_2055);
or U1724 (N_1724,In_1501,In_1341);
and U1725 (N_1725,In_2760,In_2103);
or U1726 (N_1726,In_2894,In_1072);
or U1727 (N_1727,In_188,In_190);
nor U1728 (N_1728,In_1401,In_1498);
or U1729 (N_1729,In_1415,In_27);
or U1730 (N_1730,In_2699,In_1054);
or U1731 (N_1731,In_516,In_2307);
xnor U1732 (N_1732,In_1912,In_1695);
nand U1733 (N_1733,In_1972,In_1214);
and U1734 (N_1734,In_1850,In_1101);
or U1735 (N_1735,In_1274,In_2398);
nand U1736 (N_1736,In_47,In_713);
or U1737 (N_1737,In_465,In_816);
and U1738 (N_1738,In_167,In_391);
nand U1739 (N_1739,In_680,In_2306);
nor U1740 (N_1740,In_2402,In_2436);
and U1741 (N_1741,In_881,In_1063);
nand U1742 (N_1742,In_1223,In_66);
nor U1743 (N_1743,In_434,In_2960);
and U1744 (N_1744,In_1008,In_1304);
nor U1745 (N_1745,In_90,In_1321);
and U1746 (N_1746,In_2660,In_104);
or U1747 (N_1747,In_2042,In_1168);
nand U1748 (N_1748,In_2306,In_1060);
or U1749 (N_1749,In_1595,In_711);
or U1750 (N_1750,In_2896,In_564);
nor U1751 (N_1751,In_2438,In_701);
and U1752 (N_1752,In_1995,In_643);
and U1753 (N_1753,In_1441,In_2297);
and U1754 (N_1754,In_2852,In_1746);
and U1755 (N_1755,In_2118,In_82);
or U1756 (N_1756,In_1538,In_1074);
or U1757 (N_1757,In_891,In_1657);
and U1758 (N_1758,In_2635,In_494);
and U1759 (N_1759,In_2224,In_2691);
or U1760 (N_1760,In_727,In_1101);
nor U1761 (N_1761,In_1806,In_676);
or U1762 (N_1762,In_279,In_705);
nand U1763 (N_1763,In_2070,In_1015);
nor U1764 (N_1764,In_443,In_111);
or U1765 (N_1765,In_2564,In_2783);
and U1766 (N_1766,In_600,In_441);
and U1767 (N_1767,In_1626,In_2801);
nand U1768 (N_1768,In_1925,In_215);
nor U1769 (N_1769,In_1450,In_883);
and U1770 (N_1770,In_1711,In_2835);
or U1771 (N_1771,In_896,In_2550);
nor U1772 (N_1772,In_486,In_2995);
nor U1773 (N_1773,In_2028,In_882);
or U1774 (N_1774,In_147,In_2940);
nor U1775 (N_1775,In_1711,In_2170);
and U1776 (N_1776,In_356,In_577);
and U1777 (N_1777,In_279,In_2412);
and U1778 (N_1778,In_462,In_2551);
xnor U1779 (N_1779,In_2265,In_1975);
and U1780 (N_1780,In_1307,In_2129);
nand U1781 (N_1781,In_2898,In_82);
xor U1782 (N_1782,In_1049,In_69);
and U1783 (N_1783,In_2687,In_705);
or U1784 (N_1784,In_1830,In_198);
and U1785 (N_1785,In_934,In_534);
or U1786 (N_1786,In_74,In_1174);
nor U1787 (N_1787,In_2993,In_1260);
nand U1788 (N_1788,In_850,In_201);
nor U1789 (N_1789,In_1844,In_2376);
and U1790 (N_1790,In_2072,In_872);
nand U1791 (N_1791,In_1163,In_211);
or U1792 (N_1792,In_959,In_1267);
nor U1793 (N_1793,In_1831,In_2857);
and U1794 (N_1794,In_1245,In_698);
xnor U1795 (N_1795,In_1156,In_1047);
nand U1796 (N_1796,In_1461,In_2119);
nor U1797 (N_1797,In_2440,In_2346);
nor U1798 (N_1798,In_1436,In_1864);
xor U1799 (N_1799,In_2096,In_2485);
and U1800 (N_1800,In_622,In_345);
nand U1801 (N_1801,In_1021,In_1887);
nor U1802 (N_1802,In_569,In_1876);
nor U1803 (N_1803,In_2245,In_1833);
nor U1804 (N_1804,In_1256,In_2991);
nand U1805 (N_1805,In_2659,In_564);
or U1806 (N_1806,In_384,In_2448);
and U1807 (N_1807,In_2638,In_1470);
or U1808 (N_1808,In_1577,In_2896);
nor U1809 (N_1809,In_1974,In_897);
nor U1810 (N_1810,In_476,In_361);
xor U1811 (N_1811,In_2053,In_2433);
or U1812 (N_1812,In_2991,In_2535);
and U1813 (N_1813,In_632,In_2258);
or U1814 (N_1814,In_2235,In_94);
and U1815 (N_1815,In_252,In_27);
nand U1816 (N_1816,In_2601,In_2437);
and U1817 (N_1817,In_1598,In_1987);
nand U1818 (N_1818,In_1366,In_721);
nand U1819 (N_1819,In_2159,In_2326);
xor U1820 (N_1820,In_55,In_1826);
and U1821 (N_1821,In_2099,In_1821);
nand U1822 (N_1822,In_1314,In_1457);
and U1823 (N_1823,In_37,In_1648);
or U1824 (N_1824,In_1054,In_2723);
nand U1825 (N_1825,In_593,In_2849);
nor U1826 (N_1826,In_2865,In_457);
nand U1827 (N_1827,In_2580,In_1724);
or U1828 (N_1828,In_2882,In_2490);
and U1829 (N_1829,In_614,In_2699);
and U1830 (N_1830,In_1110,In_64);
and U1831 (N_1831,In_41,In_472);
nand U1832 (N_1832,In_1487,In_1764);
and U1833 (N_1833,In_1588,In_1074);
or U1834 (N_1834,In_2694,In_417);
nor U1835 (N_1835,In_810,In_1484);
or U1836 (N_1836,In_161,In_95);
nor U1837 (N_1837,In_2952,In_2730);
and U1838 (N_1838,In_1712,In_2786);
nand U1839 (N_1839,In_2710,In_916);
nand U1840 (N_1840,In_663,In_2122);
nand U1841 (N_1841,In_2495,In_903);
nor U1842 (N_1842,In_299,In_1572);
nor U1843 (N_1843,In_677,In_30);
xnor U1844 (N_1844,In_1332,In_1608);
xnor U1845 (N_1845,In_2787,In_736);
xor U1846 (N_1846,In_133,In_969);
xnor U1847 (N_1847,In_1598,In_1438);
or U1848 (N_1848,In_2571,In_2285);
nor U1849 (N_1849,In_30,In_1175);
or U1850 (N_1850,In_1347,In_2182);
or U1851 (N_1851,In_362,In_787);
nor U1852 (N_1852,In_912,In_2208);
nor U1853 (N_1853,In_1580,In_574);
or U1854 (N_1854,In_249,In_2207);
and U1855 (N_1855,In_1970,In_2066);
nor U1856 (N_1856,In_2715,In_6);
and U1857 (N_1857,In_1736,In_2921);
and U1858 (N_1858,In_2776,In_1763);
nand U1859 (N_1859,In_2629,In_95);
and U1860 (N_1860,In_2640,In_464);
and U1861 (N_1861,In_2686,In_1925);
nand U1862 (N_1862,In_2482,In_579);
or U1863 (N_1863,In_1594,In_1287);
or U1864 (N_1864,In_2867,In_499);
nand U1865 (N_1865,In_545,In_1102);
xor U1866 (N_1866,In_2160,In_2760);
and U1867 (N_1867,In_878,In_1155);
or U1868 (N_1868,In_954,In_866);
nor U1869 (N_1869,In_277,In_781);
nand U1870 (N_1870,In_1593,In_704);
nor U1871 (N_1871,In_530,In_2333);
or U1872 (N_1872,In_1143,In_1344);
or U1873 (N_1873,In_1527,In_1282);
nand U1874 (N_1874,In_1184,In_1891);
or U1875 (N_1875,In_1145,In_2546);
nor U1876 (N_1876,In_341,In_682);
nand U1877 (N_1877,In_238,In_2785);
xor U1878 (N_1878,In_126,In_733);
xnor U1879 (N_1879,In_355,In_1833);
nor U1880 (N_1880,In_136,In_2915);
nand U1881 (N_1881,In_2826,In_1307);
nand U1882 (N_1882,In_96,In_1994);
xnor U1883 (N_1883,In_741,In_2499);
xnor U1884 (N_1884,In_1581,In_2021);
nor U1885 (N_1885,In_2557,In_2683);
nand U1886 (N_1886,In_2570,In_2750);
or U1887 (N_1887,In_2538,In_239);
nor U1888 (N_1888,In_2831,In_478);
nor U1889 (N_1889,In_2385,In_492);
nor U1890 (N_1890,In_584,In_208);
xor U1891 (N_1891,In_383,In_1192);
nor U1892 (N_1892,In_2595,In_1894);
xor U1893 (N_1893,In_1034,In_2663);
or U1894 (N_1894,In_2875,In_584);
nor U1895 (N_1895,In_96,In_536);
nand U1896 (N_1896,In_2056,In_766);
or U1897 (N_1897,In_1503,In_676);
nor U1898 (N_1898,In_2551,In_1620);
nor U1899 (N_1899,In_2178,In_1033);
nand U1900 (N_1900,In_2189,In_2755);
or U1901 (N_1901,In_2230,In_1538);
nand U1902 (N_1902,In_562,In_2371);
or U1903 (N_1903,In_280,In_1899);
nand U1904 (N_1904,In_2754,In_2327);
and U1905 (N_1905,In_2655,In_217);
nand U1906 (N_1906,In_927,In_859);
or U1907 (N_1907,In_1027,In_314);
nand U1908 (N_1908,In_2878,In_1111);
nand U1909 (N_1909,In_2450,In_2089);
nor U1910 (N_1910,In_2954,In_1514);
nor U1911 (N_1911,In_2575,In_2952);
or U1912 (N_1912,In_2548,In_516);
or U1913 (N_1913,In_2120,In_920);
nand U1914 (N_1914,In_351,In_1984);
nor U1915 (N_1915,In_2,In_1);
nor U1916 (N_1916,In_2435,In_1400);
or U1917 (N_1917,In_1002,In_1625);
nor U1918 (N_1918,In_2777,In_2820);
nor U1919 (N_1919,In_2211,In_154);
or U1920 (N_1920,In_1865,In_262);
or U1921 (N_1921,In_2802,In_673);
and U1922 (N_1922,In_1455,In_1857);
or U1923 (N_1923,In_2483,In_1096);
or U1924 (N_1924,In_751,In_1324);
xor U1925 (N_1925,In_181,In_2264);
nand U1926 (N_1926,In_1941,In_1356);
xnor U1927 (N_1927,In_2682,In_263);
nand U1928 (N_1928,In_2736,In_2303);
and U1929 (N_1929,In_2763,In_992);
or U1930 (N_1930,In_2857,In_2122);
and U1931 (N_1931,In_2530,In_2039);
nor U1932 (N_1932,In_1671,In_478);
nand U1933 (N_1933,In_749,In_556);
nand U1934 (N_1934,In_1902,In_1644);
nand U1935 (N_1935,In_25,In_1054);
nor U1936 (N_1936,In_627,In_2567);
or U1937 (N_1937,In_1717,In_2788);
xor U1938 (N_1938,In_1497,In_2136);
xor U1939 (N_1939,In_2331,In_120);
or U1940 (N_1940,In_254,In_2918);
nand U1941 (N_1941,In_2363,In_2029);
nand U1942 (N_1942,In_2811,In_2335);
and U1943 (N_1943,In_275,In_1754);
nand U1944 (N_1944,In_1873,In_1725);
and U1945 (N_1945,In_2204,In_1879);
and U1946 (N_1946,In_1550,In_1517);
nor U1947 (N_1947,In_1600,In_1628);
and U1948 (N_1948,In_2575,In_636);
nand U1949 (N_1949,In_111,In_2860);
nor U1950 (N_1950,In_500,In_1030);
and U1951 (N_1951,In_2356,In_614);
and U1952 (N_1952,In_1487,In_811);
nand U1953 (N_1953,In_1966,In_2794);
and U1954 (N_1954,In_2729,In_534);
nand U1955 (N_1955,In_1781,In_714);
xor U1956 (N_1956,In_1362,In_130);
xnor U1957 (N_1957,In_876,In_1888);
or U1958 (N_1958,In_2396,In_1193);
nor U1959 (N_1959,In_1184,In_1552);
nand U1960 (N_1960,In_326,In_1746);
nor U1961 (N_1961,In_2213,In_96);
or U1962 (N_1962,In_374,In_2348);
or U1963 (N_1963,In_2186,In_177);
nand U1964 (N_1964,In_1130,In_996);
nand U1965 (N_1965,In_1128,In_1379);
nand U1966 (N_1966,In_1690,In_1509);
nor U1967 (N_1967,In_2035,In_1426);
nor U1968 (N_1968,In_2528,In_1344);
nand U1969 (N_1969,In_1134,In_1116);
xnor U1970 (N_1970,In_2990,In_2501);
nand U1971 (N_1971,In_329,In_2593);
xor U1972 (N_1972,In_1498,In_2109);
or U1973 (N_1973,In_2646,In_2632);
nor U1974 (N_1974,In_1269,In_316);
or U1975 (N_1975,In_2099,In_1958);
nor U1976 (N_1976,In_2505,In_2898);
nor U1977 (N_1977,In_2400,In_831);
and U1978 (N_1978,In_2020,In_2854);
xnor U1979 (N_1979,In_2545,In_2334);
nor U1980 (N_1980,In_2397,In_2132);
nand U1981 (N_1981,In_56,In_1191);
or U1982 (N_1982,In_54,In_1214);
or U1983 (N_1983,In_167,In_1203);
or U1984 (N_1984,In_243,In_1369);
nand U1985 (N_1985,In_2829,In_1755);
or U1986 (N_1986,In_2971,In_2401);
and U1987 (N_1987,In_1145,In_2735);
nor U1988 (N_1988,In_1964,In_1388);
nor U1989 (N_1989,In_1312,In_2287);
or U1990 (N_1990,In_2357,In_2908);
or U1991 (N_1991,In_2731,In_200);
and U1992 (N_1992,In_2996,In_2884);
and U1993 (N_1993,In_2208,In_2599);
xor U1994 (N_1994,In_1260,In_2716);
nand U1995 (N_1995,In_1306,In_1799);
nor U1996 (N_1996,In_1533,In_1334);
nor U1997 (N_1997,In_830,In_955);
nor U1998 (N_1998,In_1886,In_848);
and U1999 (N_1999,In_2661,In_2943);
or U2000 (N_2000,In_1535,In_1522);
and U2001 (N_2001,In_506,In_503);
or U2002 (N_2002,In_385,In_1471);
xor U2003 (N_2003,In_1691,In_2546);
xnor U2004 (N_2004,In_2134,In_923);
nand U2005 (N_2005,In_819,In_1063);
or U2006 (N_2006,In_1344,In_2759);
nand U2007 (N_2007,In_1125,In_1549);
and U2008 (N_2008,In_2392,In_1704);
and U2009 (N_2009,In_892,In_1092);
and U2010 (N_2010,In_386,In_2091);
or U2011 (N_2011,In_377,In_781);
nand U2012 (N_2012,In_2950,In_68);
xnor U2013 (N_2013,In_1890,In_2299);
nand U2014 (N_2014,In_1259,In_1191);
nor U2015 (N_2015,In_2993,In_2402);
or U2016 (N_2016,In_542,In_1935);
nor U2017 (N_2017,In_2393,In_313);
nand U2018 (N_2018,In_2350,In_737);
xnor U2019 (N_2019,In_488,In_1918);
nand U2020 (N_2020,In_1486,In_61);
and U2021 (N_2021,In_1554,In_1511);
nor U2022 (N_2022,In_2274,In_2233);
or U2023 (N_2023,In_1857,In_362);
nand U2024 (N_2024,In_363,In_182);
nor U2025 (N_2025,In_2670,In_682);
or U2026 (N_2026,In_2993,In_1590);
xnor U2027 (N_2027,In_1953,In_922);
or U2028 (N_2028,In_1456,In_2110);
xnor U2029 (N_2029,In_234,In_857);
nand U2030 (N_2030,In_2087,In_2697);
nand U2031 (N_2031,In_958,In_1196);
or U2032 (N_2032,In_2387,In_1964);
and U2033 (N_2033,In_483,In_161);
or U2034 (N_2034,In_2332,In_2158);
nand U2035 (N_2035,In_150,In_199);
nor U2036 (N_2036,In_1269,In_505);
nor U2037 (N_2037,In_1848,In_142);
and U2038 (N_2038,In_404,In_2710);
nor U2039 (N_2039,In_2249,In_2451);
nor U2040 (N_2040,In_1999,In_2154);
or U2041 (N_2041,In_2587,In_1421);
and U2042 (N_2042,In_1491,In_1049);
and U2043 (N_2043,In_2313,In_1613);
nand U2044 (N_2044,In_1367,In_1836);
and U2045 (N_2045,In_2461,In_2167);
and U2046 (N_2046,In_1343,In_1016);
nand U2047 (N_2047,In_2396,In_505);
nor U2048 (N_2048,In_1092,In_2414);
nand U2049 (N_2049,In_2716,In_2703);
nor U2050 (N_2050,In_1100,In_1874);
or U2051 (N_2051,In_47,In_768);
or U2052 (N_2052,In_1358,In_64);
xnor U2053 (N_2053,In_167,In_2683);
nand U2054 (N_2054,In_2447,In_606);
or U2055 (N_2055,In_2706,In_2616);
or U2056 (N_2056,In_651,In_2886);
or U2057 (N_2057,In_2405,In_2793);
nand U2058 (N_2058,In_2356,In_1804);
nand U2059 (N_2059,In_721,In_1405);
nand U2060 (N_2060,In_1430,In_2969);
or U2061 (N_2061,In_251,In_1656);
xnor U2062 (N_2062,In_2727,In_355);
or U2063 (N_2063,In_226,In_944);
nand U2064 (N_2064,In_875,In_1154);
nor U2065 (N_2065,In_2463,In_2122);
and U2066 (N_2066,In_1021,In_815);
and U2067 (N_2067,In_2859,In_369);
nand U2068 (N_2068,In_1536,In_542);
or U2069 (N_2069,In_2342,In_2461);
nand U2070 (N_2070,In_1096,In_1929);
and U2071 (N_2071,In_1503,In_235);
or U2072 (N_2072,In_2377,In_1065);
or U2073 (N_2073,In_240,In_2233);
nor U2074 (N_2074,In_2218,In_2728);
and U2075 (N_2075,In_2326,In_633);
or U2076 (N_2076,In_860,In_866);
nand U2077 (N_2077,In_42,In_2443);
nand U2078 (N_2078,In_1702,In_753);
or U2079 (N_2079,In_2376,In_1524);
and U2080 (N_2080,In_2088,In_859);
and U2081 (N_2081,In_404,In_1786);
or U2082 (N_2082,In_1439,In_1538);
xnor U2083 (N_2083,In_917,In_2611);
and U2084 (N_2084,In_1665,In_386);
nor U2085 (N_2085,In_686,In_1254);
and U2086 (N_2086,In_1175,In_58);
and U2087 (N_2087,In_888,In_2025);
xor U2088 (N_2088,In_1221,In_2165);
nor U2089 (N_2089,In_298,In_1358);
nand U2090 (N_2090,In_1639,In_515);
nor U2091 (N_2091,In_141,In_590);
and U2092 (N_2092,In_1680,In_75);
nand U2093 (N_2093,In_901,In_2682);
or U2094 (N_2094,In_1568,In_1829);
and U2095 (N_2095,In_2371,In_211);
nand U2096 (N_2096,In_2012,In_2052);
nor U2097 (N_2097,In_2294,In_1400);
nand U2098 (N_2098,In_664,In_530);
or U2099 (N_2099,In_247,In_2952);
nor U2100 (N_2100,In_2295,In_2228);
or U2101 (N_2101,In_791,In_2057);
or U2102 (N_2102,In_1628,In_1942);
nor U2103 (N_2103,In_2823,In_2901);
or U2104 (N_2104,In_1264,In_2839);
xnor U2105 (N_2105,In_864,In_2382);
or U2106 (N_2106,In_917,In_2180);
xor U2107 (N_2107,In_1557,In_1628);
or U2108 (N_2108,In_429,In_531);
and U2109 (N_2109,In_557,In_1978);
or U2110 (N_2110,In_1441,In_678);
or U2111 (N_2111,In_948,In_1545);
or U2112 (N_2112,In_1719,In_1562);
and U2113 (N_2113,In_265,In_204);
nor U2114 (N_2114,In_1684,In_1165);
nor U2115 (N_2115,In_1189,In_2965);
and U2116 (N_2116,In_741,In_2577);
nand U2117 (N_2117,In_2747,In_1289);
nor U2118 (N_2118,In_1961,In_2206);
nor U2119 (N_2119,In_466,In_503);
nand U2120 (N_2120,In_1066,In_2915);
nor U2121 (N_2121,In_796,In_1851);
xor U2122 (N_2122,In_644,In_1467);
nand U2123 (N_2123,In_2109,In_1476);
nor U2124 (N_2124,In_2514,In_283);
nor U2125 (N_2125,In_2302,In_373);
xnor U2126 (N_2126,In_2092,In_1932);
nor U2127 (N_2127,In_2226,In_1326);
nand U2128 (N_2128,In_717,In_436);
xor U2129 (N_2129,In_551,In_239);
xnor U2130 (N_2130,In_2876,In_1824);
nand U2131 (N_2131,In_2064,In_1764);
and U2132 (N_2132,In_2367,In_2049);
and U2133 (N_2133,In_2718,In_2210);
nor U2134 (N_2134,In_2091,In_2179);
xnor U2135 (N_2135,In_2158,In_2882);
xor U2136 (N_2136,In_1744,In_1021);
and U2137 (N_2137,In_1780,In_1130);
nor U2138 (N_2138,In_2293,In_16);
and U2139 (N_2139,In_1066,In_1017);
and U2140 (N_2140,In_2155,In_1040);
and U2141 (N_2141,In_1997,In_1243);
and U2142 (N_2142,In_1669,In_2920);
nor U2143 (N_2143,In_1596,In_1656);
or U2144 (N_2144,In_2309,In_311);
nand U2145 (N_2145,In_1334,In_774);
and U2146 (N_2146,In_1472,In_2638);
nor U2147 (N_2147,In_484,In_417);
xnor U2148 (N_2148,In_2755,In_2076);
and U2149 (N_2149,In_741,In_2507);
and U2150 (N_2150,In_637,In_2539);
nand U2151 (N_2151,In_2934,In_1637);
nand U2152 (N_2152,In_1867,In_1134);
or U2153 (N_2153,In_1703,In_1737);
and U2154 (N_2154,In_803,In_905);
xor U2155 (N_2155,In_437,In_1008);
and U2156 (N_2156,In_2742,In_2662);
and U2157 (N_2157,In_210,In_2642);
or U2158 (N_2158,In_2148,In_2618);
or U2159 (N_2159,In_2848,In_1766);
nand U2160 (N_2160,In_479,In_2335);
and U2161 (N_2161,In_2829,In_2945);
and U2162 (N_2162,In_1902,In_2077);
nand U2163 (N_2163,In_947,In_515);
xnor U2164 (N_2164,In_1586,In_2419);
and U2165 (N_2165,In_1055,In_93);
and U2166 (N_2166,In_601,In_1394);
or U2167 (N_2167,In_189,In_1414);
or U2168 (N_2168,In_528,In_97);
nor U2169 (N_2169,In_2768,In_650);
nand U2170 (N_2170,In_165,In_699);
and U2171 (N_2171,In_836,In_1040);
nor U2172 (N_2172,In_950,In_2494);
nand U2173 (N_2173,In_619,In_2723);
or U2174 (N_2174,In_1036,In_1413);
and U2175 (N_2175,In_1681,In_2860);
or U2176 (N_2176,In_156,In_2999);
nand U2177 (N_2177,In_2693,In_1016);
and U2178 (N_2178,In_616,In_606);
nand U2179 (N_2179,In_159,In_830);
nor U2180 (N_2180,In_2356,In_2923);
nor U2181 (N_2181,In_1605,In_2486);
and U2182 (N_2182,In_538,In_1971);
nand U2183 (N_2183,In_2119,In_920);
nor U2184 (N_2184,In_377,In_2266);
nor U2185 (N_2185,In_585,In_146);
or U2186 (N_2186,In_837,In_486);
xor U2187 (N_2187,In_340,In_2092);
nor U2188 (N_2188,In_2088,In_2572);
and U2189 (N_2189,In_2830,In_1334);
nand U2190 (N_2190,In_2741,In_2465);
or U2191 (N_2191,In_169,In_1179);
nand U2192 (N_2192,In_1789,In_2001);
or U2193 (N_2193,In_168,In_1271);
nor U2194 (N_2194,In_47,In_772);
or U2195 (N_2195,In_69,In_121);
nand U2196 (N_2196,In_1645,In_1932);
or U2197 (N_2197,In_2264,In_1819);
or U2198 (N_2198,In_1656,In_750);
nand U2199 (N_2199,In_399,In_2621);
nor U2200 (N_2200,In_1599,In_364);
nand U2201 (N_2201,In_2524,In_7);
and U2202 (N_2202,In_1732,In_2444);
and U2203 (N_2203,In_2290,In_2879);
and U2204 (N_2204,In_1151,In_212);
nand U2205 (N_2205,In_1367,In_1196);
or U2206 (N_2206,In_1602,In_2344);
xnor U2207 (N_2207,In_880,In_815);
or U2208 (N_2208,In_2810,In_955);
and U2209 (N_2209,In_2005,In_2040);
and U2210 (N_2210,In_1535,In_198);
or U2211 (N_2211,In_510,In_1084);
or U2212 (N_2212,In_1480,In_2125);
nor U2213 (N_2213,In_2674,In_1857);
nand U2214 (N_2214,In_2998,In_163);
nor U2215 (N_2215,In_1779,In_2708);
and U2216 (N_2216,In_1382,In_842);
nand U2217 (N_2217,In_155,In_1927);
nor U2218 (N_2218,In_1513,In_858);
xnor U2219 (N_2219,In_2399,In_1440);
and U2220 (N_2220,In_2854,In_2231);
nor U2221 (N_2221,In_1911,In_2354);
xnor U2222 (N_2222,In_2134,In_1871);
nand U2223 (N_2223,In_1008,In_2792);
or U2224 (N_2224,In_857,In_2808);
or U2225 (N_2225,In_2798,In_843);
or U2226 (N_2226,In_38,In_1020);
and U2227 (N_2227,In_1467,In_1649);
nand U2228 (N_2228,In_1111,In_2514);
nor U2229 (N_2229,In_1363,In_2665);
and U2230 (N_2230,In_467,In_2705);
nor U2231 (N_2231,In_713,In_2958);
and U2232 (N_2232,In_930,In_2578);
xnor U2233 (N_2233,In_1563,In_844);
or U2234 (N_2234,In_850,In_542);
and U2235 (N_2235,In_2173,In_839);
nand U2236 (N_2236,In_2837,In_347);
nand U2237 (N_2237,In_2607,In_2609);
and U2238 (N_2238,In_88,In_1749);
or U2239 (N_2239,In_2664,In_2828);
or U2240 (N_2240,In_2031,In_641);
or U2241 (N_2241,In_1359,In_1943);
nand U2242 (N_2242,In_1658,In_2604);
or U2243 (N_2243,In_829,In_1277);
nand U2244 (N_2244,In_2619,In_2641);
and U2245 (N_2245,In_1299,In_568);
or U2246 (N_2246,In_2380,In_1239);
and U2247 (N_2247,In_2251,In_1119);
nor U2248 (N_2248,In_2989,In_587);
or U2249 (N_2249,In_611,In_259);
nor U2250 (N_2250,In_917,In_588);
nand U2251 (N_2251,In_47,In_549);
nor U2252 (N_2252,In_2443,In_268);
and U2253 (N_2253,In_876,In_658);
or U2254 (N_2254,In_1700,In_2670);
nor U2255 (N_2255,In_33,In_2636);
nor U2256 (N_2256,In_1280,In_1215);
and U2257 (N_2257,In_1806,In_2832);
and U2258 (N_2258,In_1431,In_857);
nor U2259 (N_2259,In_310,In_635);
nor U2260 (N_2260,In_2612,In_706);
nand U2261 (N_2261,In_812,In_496);
nand U2262 (N_2262,In_1728,In_2773);
nor U2263 (N_2263,In_2423,In_2287);
or U2264 (N_2264,In_1801,In_1408);
nand U2265 (N_2265,In_919,In_2339);
and U2266 (N_2266,In_2804,In_1231);
and U2267 (N_2267,In_1913,In_681);
or U2268 (N_2268,In_1556,In_1627);
nand U2269 (N_2269,In_2326,In_693);
and U2270 (N_2270,In_1465,In_243);
nand U2271 (N_2271,In_2981,In_2714);
nor U2272 (N_2272,In_1130,In_714);
nor U2273 (N_2273,In_2592,In_342);
nor U2274 (N_2274,In_602,In_291);
xor U2275 (N_2275,In_1731,In_2806);
nand U2276 (N_2276,In_2239,In_195);
nand U2277 (N_2277,In_506,In_149);
and U2278 (N_2278,In_1414,In_288);
xor U2279 (N_2279,In_35,In_2066);
and U2280 (N_2280,In_1652,In_1256);
nor U2281 (N_2281,In_255,In_2583);
nor U2282 (N_2282,In_2100,In_1039);
nand U2283 (N_2283,In_814,In_1103);
and U2284 (N_2284,In_2800,In_1585);
xor U2285 (N_2285,In_2297,In_2147);
and U2286 (N_2286,In_317,In_2154);
nor U2287 (N_2287,In_2542,In_1328);
xnor U2288 (N_2288,In_168,In_2249);
and U2289 (N_2289,In_768,In_1955);
nor U2290 (N_2290,In_1508,In_1834);
nand U2291 (N_2291,In_1251,In_2486);
nand U2292 (N_2292,In_2821,In_891);
and U2293 (N_2293,In_710,In_387);
or U2294 (N_2294,In_125,In_1680);
or U2295 (N_2295,In_583,In_1611);
or U2296 (N_2296,In_2027,In_105);
xnor U2297 (N_2297,In_436,In_2855);
nand U2298 (N_2298,In_2761,In_1919);
and U2299 (N_2299,In_1164,In_1671);
nor U2300 (N_2300,In_2641,In_844);
nand U2301 (N_2301,In_1574,In_789);
nand U2302 (N_2302,In_143,In_2045);
or U2303 (N_2303,In_217,In_2765);
and U2304 (N_2304,In_2171,In_1886);
nand U2305 (N_2305,In_624,In_1553);
nor U2306 (N_2306,In_707,In_1618);
nor U2307 (N_2307,In_1943,In_2301);
or U2308 (N_2308,In_2487,In_2193);
xor U2309 (N_2309,In_927,In_2024);
nand U2310 (N_2310,In_1430,In_12);
nor U2311 (N_2311,In_1047,In_1286);
and U2312 (N_2312,In_605,In_800);
nand U2313 (N_2313,In_226,In_442);
nor U2314 (N_2314,In_1079,In_2959);
xnor U2315 (N_2315,In_2987,In_1455);
and U2316 (N_2316,In_1853,In_380);
and U2317 (N_2317,In_1452,In_2506);
xor U2318 (N_2318,In_947,In_2186);
nor U2319 (N_2319,In_1750,In_2521);
nor U2320 (N_2320,In_2105,In_2167);
nand U2321 (N_2321,In_2805,In_1597);
xnor U2322 (N_2322,In_1138,In_1974);
nand U2323 (N_2323,In_2034,In_1659);
nor U2324 (N_2324,In_1031,In_2312);
or U2325 (N_2325,In_2972,In_914);
nor U2326 (N_2326,In_1582,In_2265);
nand U2327 (N_2327,In_348,In_2429);
nor U2328 (N_2328,In_1341,In_658);
and U2329 (N_2329,In_2818,In_777);
or U2330 (N_2330,In_2368,In_1542);
nor U2331 (N_2331,In_1709,In_467);
and U2332 (N_2332,In_1181,In_1857);
nand U2333 (N_2333,In_886,In_352);
nor U2334 (N_2334,In_445,In_1449);
nor U2335 (N_2335,In_2821,In_85);
or U2336 (N_2336,In_1916,In_549);
and U2337 (N_2337,In_2827,In_438);
or U2338 (N_2338,In_390,In_33);
or U2339 (N_2339,In_1805,In_364);
nand U2340 (N_2340,In_31,In_502);
and U2341 (N_2341,In_1052,In_2718);
nor U2342 (N_2342,In_269,In_546);
nand U2343 (N_2343,In_2240,In_1335);
nand U2344 (N_2344,In_399,In_2903);
or U2345 (N_2345,In_821,In_1492);
xnor U2346 (N_2346,In_2862,In_1214);
nor U2347 (N_2347,In_1711,In_1660);
or U2348 (N_2348,In_2444,In_772);
nor U2349 (N_2349,In_2194,In_896);
or U2350 (N_2350,In_1505,In_2536);
nand U2351 (N_2351,In_1015,In_484);
nor U2352 (N_2352,In_1826,In_1596);
or U2353 (N_2353,In_435,In_1007);
nand U2354 (N_2354,In_2903,In_1951);
nor U2355 (N_2355,In_1409,In_2089);
nor U2356 (N_2356,In_2569,In_2908);
nor U2357 (N_2357,In_320,In_2231);
nand U2358 (N_2358,In_1265,In_809);
and U2359 (N_2359,In_2894,In_108);
and U2360 (N_2360,In_1063,In_1793);
or U2361 (N_2361,In_1661,In_2108);
xnor U2362 (N_2362,In_2014,In_236);
and U2363 (N_2363,In_2152,In_110);
nor U2364 (N_2364,In_1658,In_2315);
nor U2365 (N_2365,In_2079,In_51);
or U2366 (N_2366,In_1584,In_1609);
nor U2367 (N_2367,In_1212,In_2696);
and U2368 (N_2368,In_2196,In_2420);
or U2369 (N_2369,In_376,In_135);
or U2370 (N_2370,In_2234,In_436);
or U2371 (N_2371,In_738,In_1570);
and U2372 (N_2372,In_1417,In_1535);
nand U2373 (N_2373,In_741,In_1616);
or U2374 (N_2374,In_2125,In_1123);
or U2375 (N_2375,In_203,In_2524);
and U2376 (N_2376,In_272,In_2888);
nor U2377 (N_2377,In_2574,In_939);
or U2378 (N_2378,In_59,In_2153);
or U2379 (N_2379,In_1345,In_1675);
nor U2380 (N_2380,In_816,In_1928);
and U2381 (N_2381,In_2698,In_801);
and U2382 (N_2382,In_1996,In_1780);
nand U2383 (N_2383,In_424,In_602);
and U2384 (N_2384,In_2025,In_2987);
or U2385 (N_2385,In_2315,In_185);
nand U2386 (N_2386,In_2576,In_1929);
nor U2387 (N_2387,In_970,In_530);
or U2388 (N_2388,In_2207,In_1512);
or U2389 (N_2389,In_2564,In_1456);
and U2390 (N_2390,In_812,In_181);
xnor U2391 (N_2391,In_28,In_849);
xnor U2392 (N_2392,In_2379,In_2567);
nand U2393 (N_2393,In_2959,In_779);
nor U2394 (N_2394,In_2704,In_2010);
nor U2395 (N_2395,In_911,In_527);
and U2396 (N_2396,In_2910,In_905);
nor U2397 (N_2397,In_22,In_230);
or U2398 (N_2398,In_1225,In_1046);
or U2399 (N_2399,In_479,In_1327);
nand U2400 (N_2400,In_1268,In_1903);
or U2401 (N_2401,In_1581,In_2008);
or U2402 (N_2402,In_663,In_881);
nand U2403 (N_2403,In_2281,In_318);
and U2404 (N_2404,In_2499,In_1862);
nand U2405 (N_2405,In_934,In_1449);
nand U2406 (N_2406,In_2874,In_2379);
or U2407 (N_2407,In_2062,In_1609);
and U2408 (N_2408,In_1499,In_1464);
nand U2409 (N_2409,In_2340,In_2990);
nand U2410 (N_2410,In_987,In_2697);
nor U2411 (N_2411,In_394,In_744);
and U2412 (N_2412,In_824,In_1498);
and U2413 (N_2413,In_2663,In_400);
and U2414 (N_2414,In_2039,In_2171);
nor U2415 (N_2415,In_857,In_1103);
and U2416 (N_2416,In_122,In_2321);
xnor U2417 (N_2417,In_237,In_1900);
and U2418 (N_2418,In_1495,In_1681);
and U2419 (N_2419,In_606,In_1014);
and U2420 (N_2420,In_73,In_2611);
and U2421 (N_2421,In_2780,In_1778);
and U2422 (N_2422,In_2185,In_2874);
xor U2423 (N_2423,In_212,In_609);
nand U2424 (N_2424,In_1910,In_969);
and U2425 (N_2425,In_2008,In_346);
and U2426 (N_2426,In_311,In_1878);
and U2427 (N_2427,In_2207,In_179);
and U2428 (N_2428,In_422,In_797);
nand U2429 (N_2429,In_542,In_2112);
xnor U2430 (N_2430,In_2078,In_2229);
nand U2431 (N_2431,In_2051,In_1581);
or U2432 (N_2432,In_1562,In_1556);
or U2433 (N_2433,In_1149,In_747);
and U2434 (N_2434,In_2917,In_730);
nor U2435 (N_2435,In_606,In_1004);
and U2436 (N_2436,In_99,In_518);
nor U2437 (N_2437,In_1721,In_2970);
nor U2438 (N_2438,In_2959,In_1778);
nor U2439 (N_2439,In_2276,In_2112);
nor U2440 (N_2440,In_1814,In_217);
nand U2441 (N_2441,In_2636,In_1868);
nor U2442 (N_2442,In_211,In_2654);
nand U2443 (N_2443,In_1566,In_52);
and U2444 (N_2444,In_773,In_2333);
or U2445 (N_2445,In_632,In_421);
xnor U2446 (N_2446,In_1604,In_1479);
nor U2447 (N_2447,In_1157,In_31);
and U2448 (N_2448,In_2182,In_2534);
xnor U2449 (N_2449,In_968,In_2947);
nand U2450 (N_2450,In_1158,In_2703);
nand U2451 (N_2451,In_899,In_1999);
xor U2452 (N_2452,In_1242,In_1333);
and U2453 (N_2453,In_1899,In_2828);
nor U2454 (N_2454,In_746,In_2941);
nand U2455 (N_2455,In_1670,In_447);
nand U2456 (N_2456,In_217,In_2343);
and U2457 (N_2457,In_1363,In_2121);
xor U2458 (N_2458,In_1263,In_1268);
or U2459 (N_2459,In_1149,In_133);
nor U2460 (N_2460,In_2444,In_2654);
and U2461 (N_2461,In_1046,In_1416);
nand U2462 (N_2462,In_2105,In_1720);
and U2463 (N_2463,In_2080,In_945);
xnor U2464 (N_2464,In_533,In_1711);
and U2465 (N_2465,In_480,In_1112);
and U2466 (N_2466,In_1445,In_2848);
nor U2467 (N_2467,In_1549,In_2345);
nor U2468 (N_2468,In_2975,In_1787);
nand U2469 (N_2469,In_1510,In_1168);
and U2470 (N_2470,In_2409,In_2026);
nand U2471 (N_2471,In_2317,In_2868);
and U2472 (N_2472,In_1143,In_949);
nand U2473 (N_2473,In_2855,In_1665);
or U2474 (N_2474,In_2652,In_1065);
and U2475 (N_2475,In_584,In_380);
nand U2476 (N_2476,In_1036,In_1479);
nand U2477 (N_2477,In_1028,In_1367);
nor U2478 (N_2478,In_233,In_2199);
or U2479 (N_2479,In_2509,In_734);
or U2480 (N_2480,In_1178,In_2762);
xnor U2481 (N_2481,In_665,In_1503);
and U2482 (N_2482,In_2110,In_1832);
nand U2483 (N_2483,In_2710,In_2309);
or U2484 (N_2484,In_408,In_1927);
nor U2485 (N_2485,In_827,In_940);
and U2486 (N_2486,In_1825,In_145);
nor U2487 (N_2487,In_317,In_1318);
xnor U2488 (N_2488,In_1814,In_2902);
or U2489 (N_2489,In_591,In_1517);
or U2490 (N_2490,In_1668,In_1648);
nand U2491 (N_2491,In_655,In_1945);
or U2492 (N_2492,In_844,In_1278);
nand U2493 (N_2493,In_2236,In_1436);
or U2494 (N_2494,In_726,In_1057);
and U2495 (N_2495,In_900,In_1261);
nand U2496 (N_2496,In_2454,In_1724);
nor U2497 (N_2497,In_1004,In_2080);
nor U2498 (N_2498,In_2972,In_1635);
nor U2499 (N_2499,In_936,In_212);
nor U2500 (N_2500,In_2688,In_1686);
and U2501 (N_2501,In_2286,In_596);
nand U2502 (N_2502,In_1965,In_353);
or U2503 (N_2503,In_2951,In_604);
nor U2504 (N_2504,In_2783,In_1575);
xnor U2505 (N_2505,In_2098,In_2867);
nand U2506 (N_2506,In_2828,In_1019);
nor U2507 (N_2507,In_799,In_385);
nor U2508 (N_2508,In_530,In_2912);
nor U2509 (N_2509,In_1131,In_2917);
nor U2510 (N_2510,In_610,In_2186);
nor U2511 (N_2511,In_2904,In_1558);
nor U2512 (N_2512,In_373,In_1753);
xor U2513 (N_2513,In_2997,In_677);
nand U2514 (N_2514,In_2805,In_1376);
nand U2515 (N_2515,In_2440,In_1266);
xnor U2516 (N_2516,In_142,In_2061);
or U2517 (N_2517,In_1014,In_554);
or U2518 (N_2518,In_1451,In_471);
nor U2519 (N_2519,In_477,In_1752);
nand U2520 (N_2520,In_700,In_1058);
nand U2521 (N_2521,In_643,In_2233);
and U2522 (N_2522,In_37,In_2741);
or U2523 (N_2523,In_1023,In_2975);
xor U2524 (N_2524,In_13,In_2340);
nor U2525 (N_2525,In_2722,In_1823);
and U2526 (N_2526,In_447,In_2914);
nor U2527 (N_2527,In_2944,In_220);
and U2528 (N_2528,In_531,In_2309);
and U2529 (N_2529,In_1005,In_336);
or U2530 (N_2530,In_141,In_996);
or U2531 (N_2531,In_1680,In_1997);
and U2532 (N_2532,In_2631,In_2504);
and U2533 (N_2533,In_880,In_695);
nand U2534 (N_2534,In_345,In_15);
nor U2535 (N_2535,In_1768,In_1526);
xor U2536 (N_2536,In_1059,In_183);
nand U2537 (N_2537,In_2258,In_1860);
or U2538 (N_2538,In_1071,In_18);
and U2539 (N_2539,In_1918,In_557);
nand U2540 (N_2540,In_1038,In_1213);
nor U2541 (N_2541,In_741,In_1051);
or U2542 (N_2542,In_871,In_1252);
nand U2543 (N_2543,In_1874,In_2015);
nor U2544 (N_2544,In_1213,In_1727);
and U2545 (N_2545,In_1639,In_1293);
xnor U2546 (N_2546,In_641,In_2939);
or U2547 (N_2547,In_1869,In_2553);
or U2548 (N_2548,In_952,In_799);
or U2549 (N_2549,In_1609,In_744);
and U2550 (N_2550,In_2276,In_2064);
nand U2551 (N_2551,In_809,In_1982);
nor U2552 (N_2552,In_1641,In_1011);
nor U2553 (N_2553,In_12,In_2493);
and U2554 (N_2554,In_749,In_2869);
nand U2555 (N_2555,In_402,In_1590);
nand U2556 (N_2556,In_1966,In_426);
or U2557 (N_2557,In_2397,In_2362);
or U2558 (N_2558,In_1754,In_1303);
and U2559 (N_2559,In_1242,In_2668);
nand U2560 (N_2560,In_1736,In_651);
xor U2561 (N_2561,In_1721,In_1906);
nor U2562 (N_2562,In_2256,In_1326);
xnor U2563 (N_2563,In_1662,In_1698);
nor U2564 (N_2564,In_2855,In_2508);
and U2565 (N_2565,In_179,In_1183);
and U2566 (N_2566,In_2613,In_386);
nor U2567 (N_2567,In_133,In_1883);
nand U2568 (N_2568,In_1803,In_2991);
or U2569 (N_2569,In_1960,In_2868);
nor U2570 (N_2570,In_109,In_1128);
or U2571 (N_2571,In_2180,In_1139);
or U2572 (N_2572,In_1807,In_2830);
and U2573 (N_2573,In_2691,In_2781);
and U2574 (N_2574,In_425,In_2893);
and U2575 (N_2575,In_1902,In_1477);
and U2576 (N_2576,In_632,In_557);
nand U2577 (N_2577,In_730,In_1503);
or U2578 (N_2578,In_1518,In_505);
and U2579 (N_2579,In_534,In_1696);
xor U2580 (N_2580,In_2561,In_1798);
or U2581 (N_2581,In_1118,In_69);
and U2582 (N_2582,In_2158,In_1398);
or U2583 (N_2583,In_1181,In_549);
nor U2584 (N_2584,In_2478,In_1576);
and U2585 (N_2585,In_579,In_31);
or U2586 (N_2586,In_2602,In_756);
xnor U2587 (N_2587,In_1998,In_1539);
nand U2588 (N_2588,In_1733,In_175);
nor U2589 (N_2589,In_1130,In_854);
nand U2590 (N_2590,In_413,In_455);
and U2591 (N_2591,In_1238,In_2401);
nor U2592 (N_2592,In_2122,In_1580);
nor U2593 (N_2593,In_2696,In_1808);
and U2594 (N_2594,In_302,In_2);
or U2595 (N_2595,In_2371,In_2643);
nor U2596 (N_2596,In_2950,In_2069);
nand U2597 (N_2597,In_1585,In_1536);
xnor U2598 (N_2598,In_886,In_1064);
nor U2599 (N_2599,In_415,In_309);
nand U2600 (N_2600,In_839,In_953);
xor U2601 (N_2601,In_1473,In_137);
nand U2602 (N_2602,In_1777,In_1682);
nor U2603 (N_2603,In_2655,In_2834);
xor U2604 (N_2604,In_2026,In_2900);
or U2605 (N_2605,In_2508,In_896);
nand U2606 (N_2606,In_1575,In_695);
or U2607 (N_2607,In_2923,In_2877);
nand U2608 (N_2608,In_1378,In_2162);
nand U2609 (N_2609,In_2245,In_2985);
xnor U2610 (N_2610,In_529,In_1102);
or U2611 (N_2611,In_662,In_2494);
nand U2612 (N_2612,In_588,In_1153);
nand U2613 (N_2613,In_1977,In_2942);
or U2614 (N_2614,In_2894,In_2832);
nor U2615 (N_2615,In_484,In_1609);
and U2616 (N_2616,In_2817,In_2566);
nor U2617 (N_2617,In_43,In_1717);
nand U2618 (N_2618,In_1475,In_981);
xnor U2619 (N_2619,In_2873,In_1078);
xor U2620 (N_2620,In_397,In_2814);
or U2621 (N_2621,In_297,In_2185);
nand U2622 (N_2622,In_921,In_1028);
and U2623 (N_2623,In_1810,In_850);
nand U2624 (N_2624,In_2507,In_760);
nor U2625 (N_2625,In_991,In_675);
nand U2626 (N_2626,In_1679,In_2127);
nor U2627 (N_2627,In_701,In_1333);
and U2628 (N_2628,In_110,In_768);
and U2629 (N_2629,In_591,In_2261);
nor U2630 (N_2630,In_2363,In_2467);
nor U2631 (N_2631,In_504,In_2762);
and U2632 (N_2632,In_2774,In_1433);
and U2633 (N_2633,In_979,In_27);
nor U2634 (N_2634,In_2205,In_1075);
or U2635 (N_2635,In_1404,In_865);
and U2636 (N_2636,In_594,In_512);
nand U2637 (N_2637,In_529,In_2109);
nand U2638 (N_2638,In_67,In_1301);
or U2639 (N_2639,In_394,In_1455);
nor U2640 (N_2640,In_2506,In_2905);
nand U2641 (N_2641,In_1930,In_2118);
or U2642 (N_2642,In_1880,In_1191);
and U2643 (N_2643,In_1044,In_1000);
xor U2644 (N_2644,In_2227,In_2940);
xnor U2645 (N_2645,In_1585,In_1095);
nor U2646 (N_2646,In_775,In_1151);
and U2647 (N_2647,In_1599,In_2478);
and U2648 (N_2648,In_2246,In_1646);
nor U2649 (N_2649,In_2924,In_1225);
and U2650 (N_2650,In_226,In_2094);
nand U2651 (N_2651,In_1249,In_1563);
and U2652 (N_2652,In_1956,In_2878);
xnor U2653 (N_2653,In_30,In_230);
and U2654 (N_2654,In_523,In_1470);
nor U2655 (N_2655,In_2523,In_1696);
nor U2656 (N_2656,In_1754,In_1054);
nand U2657 (N_2657,In_1401,In_2687);
nor U2658 (N_2658,In_1675,In_1503);
xnor U2659 (N_2659,In_2274,In_282);
and U2660 (N_2660,In_1081,In_2059);
nand U2661 (N_2661,In_1644,In_736);
nor U2662 (N_2662,In_2324,In_1284);
or U2663 (N_2663,In_2222,In_2518);
nor U2664 (N_2664,In_1251,In_296);
nand U2665 (N_2665,In_560,In_1785);
nor U2666 (N_2666,In_2214,In_1291);
nand U2667 (N_2667,In_427,In_1993);
xor U2668 (N_2668,In_1346,In_2554);
or U2669 (N_2669,In_2830,In_2379);
nor U2670 (N_2670,In_689,In_340);
nand U2671 (N_2671,In_1301,In_2874);
nor U2672 (N_2672,In_2982,In_2567);
nand U2673 (N_2673,In_2056,In_2886);
nand U2674 (N_2674,In_2239,In_1242);
and U2675 (N_2675,In_2189,In_593);
and U2676 (N_2676,In_639,In_1394);
nor U2677 (N_2677,In_2514,In_0);
and U2678 (N_2678,In_1652,In_467);
or U2679 (N_2679,In_1992,In_258);
nor U2680 (N_2680,In_2957,In_2859);
and U2681 (N_2681,In_167,In_1387);
nor U2682 (N_2682,In_367,In_157);
and U2683 (N_2683,In_2807,In_838);
xnor U2684 (N_2684,In_2959,In_2586);
nor U2685 (N_2685,In_510,In_197);
and U2686 (N_2686,In_611,In_162);
nor U2687 (N_2687,In_2417,In_1314);
nand U2688 (N_2688,In_1685,In_2466);
and U2689 (N_2689,In_1698,In_1961);
or U2690 (N_2690,In_87,In_2599);
nand U2691 (N_2691,In_19,In_2732);
xnor U2692 (N_2692,In_1486,In_2097);
nand U2693 (N_2693,In_711,In_2306);
nand U2694 (N_2694,In_2271,In_2559);
nand U2695 (N_2695,In_1553,In_253);
and U2696 (N_2696,In_1609,In_2880);
nand U2697 (N_2697,In_1839,In_2596);
and U2698 (N_2698,In_487,In_2092);
and U2699 (N_2699,In_528,In_2361);
xnor U2700 (N_2700,In_537,In_981);
xor U2701 (N_2701,In_208,In_2012);
nor U2702 (N_2702,In_2382,In_2081);
xnor U2703 (N_2703,In_236,In_1096);
nor U2704 (N_2704,In_429,In_1072);
nand U2705 (N_2705,In_1081,In_1793);
nor U2706 (N_2706,In_1758,In_2380);
and U2707 (N_2707,In_2165,In_2596);
nor U2708 (N_2708,In_2618,In_2661);
nand U2709 (N_2709,In_1728,In_56);
or U2710 (N_2710,In_2096,In_555);
nor U2711 (N_2711,In_1992,In_1020);
or U2712 (N_2712,In_1889,In_1305);
nor U2713 (N_2713,In_513,In_345);
nor U2714 (N_2714,In_2396,In_1804);
nor U2715 (N_2715,In_1871,In_1507);
nor U2716 (N_2716,In_859,In_14);
xnor U2717 (N_2717,In_1915,In_1163);
nand U2718 (N_2718,In_587,In_2404);
nor U2719 (N_2719,In_2271,In_2677);
nand U2720 (N_2720,In_54,In_2722);
or U2721 (N_2721,In_1504,In_264);
or U2722 (N_2722,In_753,In_1558);
nand U2723 (N_2723,In_250,In_2928);
nor U2724 (N_2724,In_2354,In_1985);
nand U2725 (N_2725,In_606,In_2920);
nor U2726 (N_2726,In_122,In_1715);
nand U2727 (N_2727,In_1208,In_1544);
or U2728 (N_2728,In_2056,In_2036);
or U2729 (N_2729,In_2971,In_668);
and U2730 (N_2730,In_2877,In_457);
nor U2731 (N_2731,In_2815,In_366);
and U2732 (N_2732,In_1341,In_297);
nor U2733 (N_2733,In_1485,In_417);
and U2734 (N_2734,In_2302,In_117);
nor U2735 (N_2735,In_1062,In_260);
nor U2736 (N_2736,In_2585,In_709);
nor U2737 (N_2737,In_1417,In_970);
xor U2738 (N_2738,In_221,In_417);
or U2739 (N_2739,In_427,In_1430);
and U2740 (N_2740,In_1814,In_2920);
xnor U2741 (N_2741,In_2215,In_1002);
or U2742 (N_2742,In_1646,In_2218);
nand U2743 (N_2743,In_1475,In_2813);
nor U2744 (N_2744,In_1079,In_2893);
and U2745 (N_2745,In_2049,In_1620);
or U2746 (N_2746,In_2819,In_484);
or U2747 (N_2747,In_1378,In_1396);
nor U2748 (N_2748,In_496,In_1461);
or U2749 (N_2749,In_2752,In_2448);
nand U2750 (N_2750,In_2595,In_605);
or U2751 (N_2751,In_2238,In_2184);
xor U2752 (N_2752,In_2661,In_295);
nand U2753 (N_2753,In_274,In_1651);
or U2754 (N_2754,In_1475,In_500);
or U2755 (N_2755,In_2295,In_542);
nor U2756 (N_2756,In_1420,In_1764);
or U2757 (N_2757,In_1209,In_1720);
or U2758 (N_2758,In_1845,In_1483);
and U2759 (N_2759,In_2650,In_2819);
or U2760 (N_2760,In_816,In_1725);
nor U2761 (N_2761,In_2794,In_520);
or U2762 (N_2762,In_1567,In_100);
xor U2763 (N_2763,In_1971,In_1794);
and U2764 (N_2764,In_241,In_631);
and U2765 (N_2765,In_855,In_729);
nand U2766 (N_2766,In_272,In_72);
xnor U2767 (N_2767,In_1325,In_2633);
or U2768 (N_2768,In_167,In_2908);
or U2769 (N_2769,In_1791,In_1761);
and U2770 (N_2770,In_1141,In_445);
or U2771 (N_2771,In_1549,In_446);
nor U2772 (N_2772,In_2070,In_2582);
nor U2773 (N_2773,In_1154,In_2437);
xor U2774 (N_2774,In_609,In_1926);
nor U2775 (N_2775,In_158,In_107);
nor U2776 (N_2776,In_204,In_1988);
nand U2777 (N_2777,In_2012,In_853);
or U2778 (N_2778,In_465,In_1904);
or U2779 (N_2779,In_928,In_2934);
or U2780 (N_2780,In_2612,In_1537);
nand U2781 (N_2781,In_2904,In_168);
nor U2782 (N_2782,In_334,In_1564);
or U2783 (N_2783,In_2852,In_1029);
or U2784 (N_2784,In_1505,In_1838);
nor U2785 (N_2785,In_1216,In_765);
and U2786 (N_2786,In_2708,In_1321);
or U2787 (N_2787,In_2043,In_795);
xnor U2788 (N_2788,In_1455,In_1212);
nand U2789 (N_2789,In_353,In_2368);
and U2790 (N_2790,In_2629,In_269);
or U2791 (N_2791,In_2091,In_627);
or U2792 (N_2792,In_2568,In_905);
nand U2793 (N_2793,In_1918,In_427);
or U2794 (N_2794,In_2289,In_2890);
nor U2795 (N_2795,In_1040,In_1779);
and U2796 (N_2796,In_1926,In_247);
and U2797 (N_2797,In_544,In_2888);
and U2798 (N_2798,In_2626,In_1726);
nand U2799 (N_2799,In_503,In_2496);
and U2800 (N_2800,In_2501,In_791);
or U2801 (N_2801,In_512,In_234);
or U2802 (N_2802,In_1155,In_1863);
xor U2803 (N_2803,In_1408,In_2138);
nand U2804 (N_2804,In_1102,In_2997);
or U2805 (N_2805,In_1124,In_1106);
nor U2806 (N_2806,In_1708,In_2675);
or U2807 (N_2807,In_1087,In_408);
or U2808 (N_2808,In_2132,In_1820);
nand U2809 (N_2809,In_137,In_1293);
or U2810 (N_2810,In_855,In_2895);
and U2811 (N_2811,In_640,In_259);
nand U2812 (N_2812,In_1770,In_1714);
nand U2813 (N_2813,In_1625,In_1465);
and U2814 (N_2814,In_420,In_2469);
or U2815 (N_2815,In_930,In_2594);
nand U2816 (N_2816,In_715,In_2979);
nand U2817 (N_2817,In_2187,In_491);
and U2818 (N_2818,In_1286,In_117);
or U2819 (N_2819,In_1134,In_122);
nor U2820 (N_2820,In_1538,In_2515);
or U2821 (N_2821,In_2608,In_1990);
or U2822 (N_2822,In_1029,In_1147);
nor U2823 (N_2823,In_143,In_2176);
nor U2824 (N_2824,In_213,In_1751);
or U2825 (N_2825,In_2344,In_1135);
and U2826 (N_2826,In_2810,In_1118);
xnor U2827 (N_2827,In_1414,In_2760);
and U2828 (N_2828,In_1143,In_2717);
or U2829 (N_2829,In_1243,In_1580);
or U2830 (N_2830,In_996,In_129);
xnor U2831 (N_2831,In_808,In_1457);
or U2832 (N_2832,In_2759,In_1082);
xnor U2833 (N_2833,In_544,In_473);
xnor U2834 (N_2834,In_893,In_2201);
nor U2835 (N_2835,In_2828,In_2502);
and U2836 (N_2836,In_2974,In_1662);
nor U2837 (N_2837,In_511,In_503);
nor U2838 (N_2838,In_1833,In_1568);
nand U2839 (N_2839,In_2237,In_1879);
nand U2840 (N_2840,In_2774,In_329);
nand U2841 (N_2841,In_2750,In_1437);
xnor U2842 (N_2842,In_1622,In_1771);
or U2843 (N_2843,In_1074,In_254);
and U2844 (N_2844,In_2410,In_2887);
xor U2845 (N_2845,In_1820,In_619);
nor U2846 (N_2846,In_361,In_2765);
nand U2847 (N_2847,In_2822,In_694);
or U2848 (N_2848,In_2885,In_1840);
xor U2849 (N_2849,In_2036,In_1558);
or U2850 (N_2850,In_2982,In_234);
nand U2851 (N_2851,In_516,In_1673);
or U2852 (N_2852,In_2953,In_2062);
nor U2853 (N_2853,In_283,In_345);
and U2854 (N_2854,In_2909,In_1436);
nand U2855 (N_2855,In_1500,In_2174);
xor U2856 (N_2856,In_2762,In_408);
nand U2857 (N_2857,In_2981,In_1887);
nand U2858 (N_2858,In_1594,In_2061);
nand U2859 (N_2859,In_1059,In_2588);
or U2860 (N_2860,In_1720,In_1573);
nand U2861 (N_2861,In_1957,In_491);
and U2862 (N_2862,In_2220,In_1989);
nor U2863 (N_2863,In_1587,In_1263);
nor U2864 (N_2864,In_1845,In_1012);
nand U2865 (N_2865,In_2155,In_1752);
and U2866 (N_2866,In_1765,In_2066);
xnor U2867 (N_2867,In_1203,In_1329);
nor U2868 (N_2868,In_2304,In_2995);
nand U2869 (N_2869,In_2828,In_2007);
nand U2870 (N_2870,In_75,In_1902);
or U2871 (N_2871,In_2475,In_1990);
nand U2872 (N_2872,In_718,In_125);
nand U2873 (N_2873,In_1290,In_2862);
nor U2874 (N_2874,In_643,In_2577);
nor U2875 (N_2875,In_935,In_1158);
or U2876 (N_2876,In_593,In_1872);
nand U2877 (N_2877,In_2156,In_130);
nand U2878 (N_2878,In_2908,In_1163);
or U2879 (N_2879,In_557,In_960);
or U2880 (N_2880,In_239,In_1266);
nand U2881 (N_2881,In_1892,In_2576);
nor U2882 (N_2882,In_815,In_2736);
and U2883 (N_2883,In_1985,In_2397);
nor U2884 (N_2884,In_406,In_929);
nor U2885 (N_2885,In_745,In_1055);
nor U2886 (N_2886,In_1858,In_355);
and U2887 (N_2887,In_2454,In_1006);
or U2888 (N_2888,In_1744,In_112);
xor U2889 (N_2889,In_2118,In_654);
xnor U2890 (N_2890,In_1746,In_1092);
nand U2891 (N_2891,In_1938,In_1359);
or U2892 (N_2892,In_1202,In_2587);
nand U2893 (N_2893,In_2300,In_1226);
nand U2894 (N_2894,In_1042,In_2648);
or U2895 (N_2895,In_840,In_2233);
and U2896 (N_2896,In_485,In_2763);
nor U2897 (N_2897,In_642,In_1152);
and U2898 (N_2898,In_1600,In_1691);
or U2899 (N_2899,In_192,In_2358);
nand U2900 (N_2900,In_110,In_2671);
nor U2901 (N_2901,In_2219,In_265);
and U2902 (N_2902,In_170,In_2794);
or U2903 (N_2903,In_2271,In_1328);
and U2904 (N_2904,In_1960,In_2054);
or U2905 (N_2905,In_835,In_1680);
or U2906 (N_2906,In_660,In_573);
and U2907 (N_2907,In_2552,In_355);
and U2908 (N_2908,In_1794,In_2924);
and U2909 (N_2909,In_623,In_763);
and U2910 (N_2910,In_949,In_2313);
nor U2911 (N_2911,In_945,In_1969);
or U2912 (N_2912,In_1494,In_887);
nand U2913 (N_2913,In_33,In_1331);
or U2914 (N_2914,In_2093,In_787);
nand U2915 (N_2915,In_1923,In_584);
nor U2916 (N_2916,In_1770,In_1148);
nand U2917 (N_2917,In_2647,In_2970);
or U2918 (N_2918,In_2092,In_2406);
or U2919 (N_2919,In_835,In_2922);
xor U2920 (N_2920,In_772,In_881);
and U2921 (N_2921,In_1427,In_975);
or U2922 (N_2922,In_2987,In_2304);
nor U2923 (N_2923,In_1177,In_1790);
or U2924 (N_2924,In_2392,In_2515);
and U2925 (N_2925,In_946,In_704);
and U2926 (N_2926,In_2974,In_2475);
or U2927 (N_2927,In_1046,In_2362);
nor U2928 (N_2928,In_2024,In_850);
nand U2929 (N_2929,In_2094,In_1538);
nand U2930 (N_2930,In_2434,In_1997);
nand U2931 (N_2931,In_2317,In_1814);
nor U2932 (N_2932,In_697,In_545);
and U2933 (N_2933,In_1577,In_2096);
nor U2934 (N_2934,In_239,In_1198);
or U2935 (N_2935,In_2787,In_2652);
and U2936 (N_2936,In_89,In_1143);
nor U2937 (N_2937,In_2331,In_1927);
xor U2938 (N_2938,In_71,In_1046);
or U2939 (N_2939,In_1776,In_1378);
nor U2940 (N_2940,In_2270,In_2032);
or U2941 (N_2941,In_1014,In_809);
nor U2942 (N_2942,In_670,In_1161);
or U2943 (N_2943,In_2983,In_1983);
nor U2944 (N_2944,In_2714,In_2296);
nand U2945 (N_2945,In_740,In_967);
xor U2946 (N_2946,In_2136,In_2748);
nand U2947 (N_2947,In_109,In_2012);
or U2948 (N_2948,In_2960,In_1915);
xor U2949 (N_2949,In_454,In_1223);
nand U2950 (N_2950,In_1338,In_2457);
or U2951 (N_2951,In_2982,In_223);
or U2952 (N_2952,In_538,In_2584);
and U2953 (N_2953,In_1678,In_2594);
nand U2954 (N_2954,In_1916,In_2051);
nand U2955 (N_2955,In_2429,In_2471);
and U2956 (N_2956,In_1567,In_2411);
nor U2957 (N_2957,In_1006,In_1715);
nand U2958 (N_2958,In_521,In_259);
or U2959 (N_2959,In_2524,In_1113);
nor U2960 (N_2960,In_2799,In_2525);
nor U2961 (N_2961,In_1461,In_476);
nor U2962 (N_2962,In_2818,In_870);
nor U2963 (N_2963,In_1079,In_2093);
nand U2964 (N_2964,In_1567,In_1663);
nand U2965 (N_2965,In_313,In_2615);
nor U2966 (N_2966,In_1031,In_2420);
nand U2967 (N_2967,In_1338,In_1712);
nor U2968 (N_2968,In_1415,In_2565);
and U2969 (N_2969,In_556,In_1614);
nor U2970 (N_2970,In_1488,In_2305);
and U2971 (N_2971,In_2222,In_166);
nor U2972 (N_2972,In_2734,In_987);
and U2973 (N_2973,In_1641,In_1538);
and U2974 (N_2974,In_2992,In_1430);
or U2975 (N_2975,In_787,In_1926);
nor U2976 (N_2976,In_332,In_2418);
or U2977 (N_2977,In_2829,In_2475);
nor U2978 (N_2978,In_1610,In_2771);
nor U2979 (N_2979,In_2500,In_531);
and U2980 (N_2980,In_2671,In_2449);
nand U2981 (N_2981,In_644,In_301);
xnor U2982 (N_2982,In_2521,In_750);
or U2983 (N_2983,In_1280,In_1852);
nand U2984 (N_2984,In_1359,In_1431);
or U2985 (N_2985,In_2603,In_2361);
nand U2986 (N_2986,In_468,In_22);
nand U2987 (N_2987,In_2899,In_2657);
xor U2988 (N_2988,In_2502,In_6);
nand U2989 (N_2989,In_1921,In_1633);
nand U2990 (N_2990,In_1131,In_2920);
and U2991 (N_2991,In_2979,In_7);
or U2992 (N_2992,In_1675,In_1250);
and U2993 (N_2993,In_733,In_378);
nand U2994 (N_2994,In_2643,In_1026);
and U2995 (N_2995,In_1540,In_2989);
nor U2996 (N_2996,In_568,In_2369);
nand U2997 (N_2997,In_1597,In_182);
xor U2998 (N_2998,In_1093,In_2075);
nand U2999 (N_2999,In_1499,In_2201);
nor U3000 (N_3000,In_2452,In_1356);
or U3001 (N_3001,In_1323,In_2302);
xor U3002 (N_3002,In_464,In_824);
and U3003 (N_3003,In_432,In_2764);
or U3004 (N_3004,In_2176,In_200);
nand U3005 (N_3005,In_2322,In_2674);
nor U3006 (N_3006,In_1819,In_2808);
nor U3007 (N_3007,In_2953,In_2721);
and U3008 (N_3008,In_1070,In_252);
or U3009 (N_3009,In_2250,In_2472);
or U3010 (N_3010,In_2564,In_670);
or U3011 (N_3011,In_2212,In_555);
nor U3012 (N_3012,In_1257,In_1199);
nor U3013 (N_3013,In_2377,In_2402);
nand U3014 (N_3014,In_842,In_2690);
xor U3015 (N_3015,In_1341,In_1786);
and U3016 (N_3016,In_2400,In_1367);
and U3017 (N_3017,In_2899,In_849);
or U3018 (N_3018,In_1068,In_232);
nor U3019 (N_3019,In_2671,In_2768);
nand U3020 (N_3020,In_2097,In_2204);
nor U3021 (N_3021,In_1359,In_1563);
nor U3022 (N_3022,In_249,In_2539);
or U3023 (N_3023,In_962,In_204);
or U3024 (N_3024,In_2569,In_285);
nand U3025 (N_3025,In_1624,In_2359);
or U3026 (N_3026,In_2901,In_298);
or U3027 (N_3027,In_2603,In_2142);
nor U3028 (N_3028,In_924,In_2103);
nor U3029 (N_3029,In_454,In_277);
and U3030 (N_3030,In_1963,In_2796);
or U3031 (N_3031,In_1765,In_2191);
nor U3032 (N_3032,In_1200,In_576);
or U3033 (N_3033,In_1200,In_1270);
or U3034 (N_3034,In_1402,In_1685);
nand U3035 (N_3035,In_225,In_642);
xor U3036 (N_3036,In_1766,In_1876);
xor U3037 (N_3037,In_981,In_2624);
nor U3038 (N_3038,In_2886,In_1786);
nor U3039 (N_3039,In_2988,In_1680);
or U3040 (N_3040,In_1393,In_970);
and U3041 (N_3041,In_1292,In_2415);
nand U3042 (N_3042,In_2225,In_1256);
and U3043 (N_3043,In_2006,In_709);
nor U3044 (N_3044,In_2631,In_200);
nor U3045 (N_3045,In_313,In_903);
nor U3046 (N_3046,In_726,In_2200);
or U3047 (N_3047,In_1229,In_367);
nor U3048 (N_3048,In_2176,In_1788);
nand U3049 (N_3049,In_2801,In_352);
nor U3050 (N_3050,In_655,In_642);
or U3051 (N_3051,In_2653,In_363);
nor U3052 (N_3052,In_620,In_2239);
nand U3053 (N_3053,In_2493,In_1964);
or U3054 (N_3054,In_130,In_1073);
nand U3055 (N_3055,In_1660,In_605);
and U3056 (N_3056,In_2301,In_1601);
nand U3057 (N_3057,In_1368,In_1593);
nand U3058 (N_3058,In_2034,In_1068);
nand U3059 (N_3059,In_1179,In_1161);
nor U3060 (N_3060,In_2013,In_1504);
or U3061 (N_3061,In_550,In_1819);
nand U3062 (N_3062,In_96,In_2470);
or U3063 (N_3063,In_2900,In_277);
and U3064 (N_3064,In_2093,In_137);
nor U3065 (N_3065,In_187,In_1757);
nor U3066 (N_3066,In_1494,In_692);
or U3067 (N_3067,In_1681,In_170);
nor U3068 (N_3068,In_1596,In_243);
nand U3069 (N_3069,In_1792,In_1224);
nand U3070 (N_3070,In_2847,In_799);
nor U3071 (N_3071,In_1662,In_2706);
and U3072 (N_3072,In_737,In_390);
nand U3073 (N_3073,In_1182,In_1351);
nand U3074 (N_3074,In_945,In_2297);
nand U3075 (N_3075,In_2033,In_746);
or U3076 (N_3076,In_1237,In_2407);
nand U3077 (N_3077,In_2933,In_2019);
and U3078 (N_3078,In_2916,In_498);
and U3079 (N_3079,In_365,In_2106);
and U3080 (N_3080,In_1065,In_568);
xnor U3081 (N_3081,In_2387,In_985);
or U3082 (N_3082,In_800,In_590);
and U3083 (N_3083,In_2503,In_371);
nand U3084 (N_3084,In_1361,In_7);
or U3085 (N_3085,In_2172,In_982);
nor U3086 (N_3086,In_1567,In_1371);
and U3087 (N_3087,In_2740,In_1796);
and U3088 (N_3088,In_1016,In_956);
nand U3089 (N_3089,In_1609,In_492);
nor U3090 (N_3090,In_2313,In_1233);
nand U3091 (N_3091,In_1453,In_537);
nor U3092 (N_3092,In_1401,In_1317);
or U3093 (N_3093,In_1952,In_2809);
and U3094 (N_3094,In_748,In_2538);
nor U3095 (N_3095,In_604,In_1458);
nand U3096 (N_3096,In_576,In_767);
or U3097 (N_3097,In_894,In_2956);
and U3098 (N_3098,In_1425,In_2628);
or U3099 (N_3099,In_1230,In_2726);
nor U3100 (N_3100,In_438,In_1820);
nand U3101 (N_3101,In_263,In_1684);
nor U3102 (N_3102,In_968,In_2053);
nand U3103 (N_3103,In_2710,In_1096);
xnor U3104 (N_3104,In_240,In_1232);
nor U3105 (N_3105,In_568,In_2277);
xor U3106 (N_3106,In_767,In_2624);
and U3107 (N_3107,In_1030,In_2112);
nand U3108 (N_3108,In_1696,In_2580);
and U3109 (N_3109,In_1429,In_2008);
or U3110 (N_3110,In_100,In_1370);
xor U3111 (N_3111,In_2202,In_2086);
xnor U3112 (N_3112,In_383,In_2411);
nor U3113 (N_3113,In_888,In_2175);
and U3114 (N_3114,In_2637,In_1639);
nand U3115 (N_3115,In_1041,In_2164);
nor U3116 (N_3116,In_382,In_92);
nor U3117 (N_3117,In_2122,In_1011);
nor U3118 (N_3118,In_680,In_2876);
or U3119 (N_3119,In_1492,In_2460);
and U3120 (N_3120,In_1854,In_976);
or U3121 (N_3121,In_2306,In_1519);
nor U3122 (N_3122,In_1662,In_911);
nor U3123 (N_3123,In_1465,In_1022);
and U3124 (N_3124,In_1829,In_2457);
nand U3125 (N_3125,In_2860,In_839);
and U3126 (N_3126,In_2147,In_487);
nor U3127 (N_3127,In_1770,In_1578);
nand U3128 (N_3128,In_939,In_1389);
xor U3129 (N_3129,In_537,In_1297);
nor U3130 (N_3130,In_2389,In_2358);
xor U3131 (N_3131,In_796,In_2954);
or U3132 (N_3132,In_2056,In_781);
xor U3133 (N_3133,In_1769,In_2870);
nor U3134 (N_3134,In_1248,In_2362);
nor U3135 (N_3135,In_2394,In_1333);
and U3136 (N_3136,In_2084,In_447);
nor U3137 (N_3137,In_1470,In_2612);
nor U3138 (N_3138,In_710,In_1299);
nor U3139 (N_3139,In_628,In_2838);
nand U3140 (N_3140,In_1946,In_2375);
and U3141 (N_3141,In_1938,In_1088);
nor U3142 (N_3142,In_1537,In_546);
or U3143 (N_3143,In_381,In_1995);
or U3144 (N_3144,In_2149,In_272);
nor U3145 (N_3145,In_1382,In_832);
and U3146 (N_3146,In_2360,In_1825);
and U3147 (N_3147,In_744,In_716);
or U3148 (N_3148,In_537,In_1077);
or U3149 (N_3149,In_811,In_2783);
and U3150 (N_3150,In_562,In_2311);
nand U3151 (N_3151,In_663,In_2143);
nand U3152 (N_3152,In_645,In_1707);
nor U3153 (N_3153,In_2329,In_2139);
xor U3154 (N_3154,In_1867,In_415);
nor U3155 (N_3155,In_841,In_1197);
nor U3156 (N_3156,In_60,In_2565);
or U3157 (N_3157,In_2065,In_1758);
nor U3158 (N_3158,In_662,In_970);
nand U3159 (N_3159,In_974,In_234);
and U3160 (N_3160,In_1444,In_511);
and U3161 (N_3161,In_894,In_283);
or U3162 (N_3162,In_903,In_1902);
and U3163 (N_3163,In_1659,In_1083);
nand U3164 (N_3164,In_515,In_996);
nand U3165 (N_3165,In_2148,In_939);
nand U3166 (N_3166,In_1347,In_2609);
and U3167 (N_3167,In_854,In_2919);
nor U3168 (N_3168,In_1506,In_1844);
nand U3169 (N_3169,In_2417,In_2305);
or U3170 (N_3170,In_1747,In_2524);
or U3171 (N_3171,In_2336,In_2634);
nand U3172 (N_3172,In_1400,In_2076);
nand U3173 (N_3173,In_199,In_291);
or U3174 (N_3174,In_2248,In_2153);
nand U3175 (N_3175,In_1485,In_1729);
nor U3176 (N_3176,In_629,In_2193);
nand U3177 (N_3177,In_2797,In_163);
nor U3178 (N_3178,In_570,In_687);
nor U3179 (N_3179,In_2493,In_2148);
nand U3180 (N_3180,In_426,In_2024);
xor U3181 (N_3181,In_257,In_135);
nand U3182 (N_3182,In_2448,In_2702);
and U3183 (N_3183,In_406,In_157);
or U3184 (N_3184,In_2031,In_2702);
and U3185 (N_3185,In_966,In_1394);
and U3186 (N_3186,In_1011,In_2105);
nor U3187 (N_3187,In_2182,In_2247);
nor U3188 (N_3188,In_507,In_2763);
or U3189 (N_3189,In_1200,In_1495);
nand U3190 (N_3190,In_1472,In_2621);
nor U3191 (N_3191,In_1005,In_355);
nor U3192 (N_3192,In_2777,In_1887);
nor U3193 (N_3193,In_1460,In_1758);
and U3194 (N_3194,In_1449,In_2694);
nor U3195 (N_3195,In_2011,In_1507);
and U3196 (N_3196,In_2952,In_2528);
and U3197 (N_3197,In_198,In_1164);
and U3198 (N_3198,In_1846,In_567);
and U3199 (N_3199,In_1918,In_2451);
nand U3200 (N_3200,In_1127,In_768);
and U3201 (N_3201,In_2676,In_580);
nor U3202 (N_3202,In_898,In_778);
and U3203 (N_3203,In_1136,In_14);
xnor U3204 (N_3204,In_2106,In_2153);
and U3205 (N_3205,In_1078,In_1664);
nand U3206 (N_3206,In_116,In_923);
and U3207 (N_3207,In_2670,In_2856);
nor U3208 (N_3208,In_525,In_2375);
or U3209 (N_3209,In_1953,In_663);
nor U3210 (N_3210,In_1987,In_1397);
and U3211 (N_3211,In_2691,In_2245);
xor U3212 (N_3212,In_2197,In_1524);
xor U3213 (N_3213,In_118,In_2019);
nor U3214 (N_3214,In_945,In_1373);
nor U3215 (N_3215,In_741,In_438);
nor U3216 (N_3216,In_947,In_82);
and U3217 (N_3217,In_566,In_2181);
nand U3218 (N_3218,In_717,In_884);
nor U3219 (N_3219,In_427,In_1640);
nand U3220 (N_3220,In_148,In_2961);
nor U3221 (N_3221,In_1206,In_1220);
nor U3222 (N_3222,In_183,In_1466);
and U3223 (N_3223,In_954,In_284);
and U3224 (N_3224,In_920,In_2958);
nand U3225 (N_3225,In_1711,In_1380);
nand U3226 (N_3226,In_2278,In_213);
nor U3227 (N_3227,In_1085,In_1841);
or U3228 (N_3228,In_386,In_1974);
or U3229 (N_3229,In_2837,In_2630);
or U3230 (N_3230,In_1720,In_619);
xnor U3231 (N_3231,In_1481,In_401);
and U3232 (N_3232,In_1859,In_573);
xor U3233 (N_3233,In_511,In_1709);
and U3234 (N_3234,In_1155,In_902);
nand U3235 (N_3235,In_2067,In_516);
or U3236 (N_3236,In_958,In_2688);
and U3237 (N_3237,In_2455,In_2410);
nand U3238 (N_3238,In_2137,In_417);
and U3239 (N_3239,In_285,In_189);
and U3240 (N_3240,In_2362,In_829);
or U3241 (N_3241,In_1499,In_1148);
nor U3242 (N_3242,In_2002,In_834);
or U3243 (N_3243,In_277,In_22);
nand U3244 (N_3244,In_1279,In_2255);
or U3245 (N_3245,In_2742,In_314);
or U3246 (N_3246,In_2307,In_780);
nand U3247 (N_3247,In_2232,In_1109);
and U3248 (N_3248,In_1400,In_27);
nor U3249 (N_3249,In_1952,In_472);
nand U3250 (N_3250,In_51,In_1761);
and U3251 (N_3251,In_491,In_57);
and U3252 (N_3252,In_2403,In_255);
nor U3253 (N_3253,In_2386,In_1638);
and U3254 (N_3254,In_744,In_2383);
nand U3255 (N_3255,In_2788,In_1310);
nor U3256 (N_3256,In_1692,In_298);
nor U3257 (N_3257,In_2731,In_833);
or U3258 (N_3258,In_50,In_406);
nor U3259 (N_3259,In_833,In_909);
nand U3260 (N_3260,In_1334,In_816);
nor U3261 (N_3261,In_2208,In_1632);
or U3262 (N_3262,In_322,In_1840);
nor U3263 (N_3263,In_1787,In_468);
nor U3264 (N_3264,In_1274,In_1682);
nand U3265 (N_3265,In_1967,In_770);
or U3266 (N_3266,In_2713,In_1544);
or U3267 (N_3267,In_1156,In_7);
or U3268 (N_3268,In_806,In_274);
nand U3269 (N_3269,In_2702,In_1276);
or U3270 (N_3270,In_275,In_1749);
or U3271 (N_3271,In_23,In_2214);
nor U3272 (N_3272,In_669,In_1968);
or U3273 (N_3273,In_2985,In_1646);
nand U3274 (N_3274,In_1191,In_2437);
xor U3275 (N_3275,In_2633,In_838);
nor U3276 (N_3276,In_1645,In_2762);
nand U3277 (N_3277,In_1262,In_296);
or U3278 (N_3278,In_945,In_1605);
or U3279 (N_3279,In_1648,In_669);
xor U3280 (N_3280,In_1112,In_1439);
nand U3281 (N_3281,In_1712,In_1472);
nand U3282 (N_3282,In_2746,In_2038);
nor U3283 (N_3283,In_1722,In_2178);
and U3284 (N_3284,In_560,In_1549);
or U3285 (N_3285,In_1383,In_2634);
xnor U3286 (N_3286,In_2490,In_609);
or U3287 (N_3287,In_583,In_1025);
nor U3288 (N_3288,In_504,In_1877);
or U3289 (N_3289,In_2989,In_365);
nor U3290 (N_3290,In_1617,In_1277);
nor U3291 (N_3291,In_2529,In_291);
and U3292 (N_3292,In_1891,In_2612);
nand U3293 (N_3293,In_1836,In_1032);
nand U3294 (N_3294,In_1041,In_2151);
nor U3295 (N_3295,In_353,In_2825);
or U3296 (N_3296,In_1947,In_1821);
and U3297 (N_3297,In_289,In_223);
nor U3298 (N_3298,In_383,In_2009);
nor U3299 (N_3299,In_2114,In_1803);
nor U3300 (N_3300,In_1554,In_819);
nor U3301 (N_3301,In_1722,In_2857);
nor U3302 (N_3302,In_808,In_2302);
nand U3303 (N_3303,In_802,In_1822);
or U3304 (N_3304,In_2539,In_1176);
nor U3305 (N_3305,In_497,In_2447);
nand U3306 (N_3306,In_2432,In_1684);
xnor U3307 (N_3307,In_1617,In_445);
xnor U3308 (N_3308,In_2571,In_2678);
xor U3309 (N_3309,In_2459,In_2318);
and U3310 (N_3310,In_1536,In_1128);
nand U3311 (N_3311,In_492,In_2801);
and U3312 (N_3312,In_1640,In_2573);
nand U3313 (N_3313,In_186,In_2550);
or U3314 (N_3314,In_1404,In_945);
nand U3315 (N_3315,In_374,In_2270);
xor U3316 (N_3316,In_1643,In_449);
nand U3317 (N_3317,In_1938,In_1990);
or U3318 (N_3318,In_2927,In_2829);
and U3319 (N_3319,In_593,In_1387);
or U3320 (N_3320,In_11,In_1007);
and U3321 (N_3321,In_931,In_2926);
nor U3322 (N_3322,In_2583,In_1715);
nand U3323 (N_3323,In_182,In_883);
or U3324 (N_3324,In_287,In_2257);
nor U3325 (N_3325,In_965,In_235);
nor U3326 (N_3326,In_1233,In_2754);
nor U3327 (N_3327,In_2861,In_2487);
nand U3328 (N_3328,In_2929,In_1261);
xnor U3329 (N_3329,In_1799,In_2417);
nand U3330 (N_3330,In_1432,In_840);
nand U3331 (N_3331,In_2664,In_1506);
or U3332 (N_3332,In_882,In_99);
nor U3333 (N_3333,In_705,In_1691);
nand U3334 (N_3334,In_2187,In_1924);
xnor U3335 (N_3335,In_1145,In_485);
and U3336 (N_3336,In_2936,In_763);
nor U3337 (N_3337,In_955,In_1498);
or U3338 (N_3338,In_116,In_651);
nand U3339 (N_3339,In_1671,In_1141);
and U3340 (N_3340,In_1350,In_1440);
nand U3341 (N_3341,In_2270,In_2757);
nand U3342 (N_3342,In_560,In_496);
nor U3343 (N_3343,In_395,In_1027);
xnor U3344 (N_3344,In_1030,In_2286);
nand U3345 (N_3345,In_1788,In_2565);
nor U3346 (N_3346,In_2036,In_1134);
or U3347 (N_3347,In_1378,In_1966);
nand U3348 (N_3348,In_987,In_2866);
or U3349 (N_3349,In_261,In_766);
nor U3350 (N_3350,In_2090,In_952);
nand U3351 (N_3351,In_869,In_1027);
or U3352 (N_3352,In_1296,In_193);
nand U3353 (N_3353,In_1046,In_138);
nand U3354 (N_3354,In_415,In_1941);
xnor U3355 (N_3355,In_1189,In_166);
and U3356 (N_3356,In_132,In_2731);
nor U3357 (N_3357,In_1942,In_1115);
nor U3358 (N_3358,In_2151,In_626);
nor U3359 (N_3359,In_1803,In_2400);
xor U3360 (N_3360,In_2445,In_2596);
xnor U3361 (N_3361,In_16,In_2647);
nor U3362 (N_3362,In_1274,In_2305);
nand U3363 (N_3363,In_71,In_347);
xor U3364 (N_3364,In_1793,In_2511);
nand U3365 (N_3365,In_503,In_1998);
nand U3366 (N_3366,In_2703,In_2993);
or U3367 (N_3367,In_2869,In_136);
xnor U3368 (N_3368,In_2797,In_1963);
and U3369 (N_3369,In_2675,In_540);
or U3370 (N_3370,In_2473,In_1967);
nor U3371 (N_3371,In_1128,In_1390);
nor U3372 (N_3372,In_1262,In_646);
nand U3373 (N_3373,In_803,In_1949);
nor U3374 (N_3374,In_2571,In_1162);
or U3375 (N_3375,In_2934,In_161);
nand U3376 (N_3376,In_2693,In_702);
nor U3377 (N_3377,In_1812,In_935);
xor U3378 (N_3378,In_848,In_1624);
xnor U3379 (N_3379,In_648,In_2942);
nand U3380 (N_3380,In_980,In_984);
nor U3381 (N_3381,In_1566,In_783);
or U3382 (N_3382,In_2867,In_561);
nor U3383 (N_3383,In_1513,In_2542);
and U3384 (N_3384,In_2565,In_1948);
or U3385 (N_3385,In_856,In_2420);
and U3386 (N_3386,In_1400,In_192);
nand U3387 (N_3387,In_2346,In_845);
xor U3388 (N_3388,In_935,In_2113);
and U3389 (N_3389,In_422,In_1114);
or U3390 (N_3390,In_1499,In_1383);
and U3391 (N_3391,In_73,In_538);
nand U3392 (N_3392,In_347,In_1127);
or U3393 (N_3393,In_544,In_400);
and U3394 (N_3394,In_553,In_2361);
and U3395 (N_3395,In_535,In_1880);
or U3396 (N_3396,In_1370,In_2323);
nor U3397 (N_3397,In_1540,In_1444);
nor U3398 (N_3398,In_884,In_259);
or U3399 (N_3399,In_2832,In_481);
nor U3400 (N_3400,In_739,In_788);
and U3401 (N_3401,In_2774,In_2249);
or U3402 (N_3402,In_2175,In_936);
nor U3403 (N_3403,In_805,In_1278);
and U3404 (N_3404,In_622,In_2469);
nor U3405 (N_3405,In_2440,In_1294);
xor U3406 (N_3406,In_1703,In_1038);
and U3407 (N_3407,In_2342,In_1779);
and U3408 (N_3408,In_2498,In_1401);
nand U3409 (N_3409,In_1889,In_517);
nor U3410 (N_3410,In_1624,In_705);
nand U3411 (N_3411,In_206,In_144);
and U3412 (N_3412,In_2505,In_330);
and U3413 (N_3413,In_1541,In_2001);
nand U3414 (N_3414,In_537,In_531);
nor U3415 (N_3415,In_1223,In_1993);
nor U3416 (N_3416,In_796,In_239);
and U3417 (N_3417,In_1268,In_2123);
or U3418 (N_3418,In_1668,In_527);
and U3419 (N_3419,In_1168,In_2407);
xor U3420 (N_3420,In_2800,In_1475);
and U3421 (N_3421,In_1992,In_1829);
nor U3422 (N_3422,In_760,In_970);
xor U3423 (N_3423,In_889,In_2559);
and U3424 (N_3424,In_327,In_1532);
or U3425 (N_3425,In_1821,In_2548);
or U3426 (N_3426,In_2271,In_572);
and U3427 (N_3427,In_2184,In_1507);
nand U3428 (N_3428,In_1407,In_2209);
nor U3429 (N_3429,In_1155,In_1720);
or U3430 (N_3430,In_2359,In_382);
or U3431 (N_3431,In_657,In_914);
or U3432 (N_3432,In_2511,In_1884);
and U3433 (N_3433,In_2229,In_1420);
nor U3434 (N_3434,In_2669,In_19);
nand U3435 (N_3435,In_2703,In_2598);
nand U3436 (N_3436,In_1188,In_354);
nor U3437 (N_3437,In_59,In_1503);
or U3438 (N_3438,In_1805,In_618);
or U3439 (N_3439,In_344,In_2176);
nor U3440 (N_3440,In_1352,In_2193);
and U3441 (N_3441,In_2378,In_2181);
and U3442 (N_3442,In_59,In_1476);
nand U3443 (N_3443,In_483,In_1098);
and U3444 (N_3444,In_1190,In_492);
nor U3445 (N_3445,In_460,In_932);
nand U3446 (N_3446,In_2078,In_500);
or U3447 (N_3447,In_613,In_680);
nand U3448 (N_3448,In_127,In_2777);
and U3449 (N_3449,In_704,In_145);
nand U3450 (N_3450,In_205,In_2747);
or U3451 (N_3451,In_348,In_1598);
or U3452 (N_3452,In_816,In_2329);
and U3453 (N_3453,In_2272,In_2960);
or U3454 (N_3454,In_487,In_995);
or U3455 (N_3455,In_2373,In_408);
nor U3456 (N_3456,In_1424,In_2100);
nand U3457 (N_3457,In_1845,In_1237);
nor U3458 (N_3458,In_652,In_2632);
nor U3459 (N_3459,In_398,In_2764);
and U3460 (N_3460,In_211,In_1583);
and U3461 (N_3461,In_140,In_345);
or U3462 (N_3462,In_1631,In_552);
and U3463 (N_3463,In_941,In_1018);
and U3464 (N_3464,In_2467,In_2949);
nand U3465 (N_3465,In_1997,In_721);
nor U3466 (N_3466,In_1826,In_1312);
or U3467 (N_3467,In_1861,In_1524);
xnor U3468 (N_3468,In_2974,In_2176);
and U3469 (N_3469,In_2794,In_2483);
or U3470 (N_3470,In_2644,In_1484);
nor U3471 (N_3471,In_1411,In_2451);
and U3472 (N_3472,In_1467,In_383);
and U3473 (N_3473,In_375,In_1242);
or U3474 (N_3474,In_1733,In_700);
or U3475 (N_3475,In_2358,In_810);
xor U3476 (N_3476,In_2045,In_306);
nor U3477 (N_3477,In_1867,In_2012);
and U3478 (N_3478,In_1439,In_1674);
nor U3479 (N_3479,In_1166,In_2647);
xnor U3480 (N_3480,In_1773,In_382);
or U3481 (N_3481,In_2193,In_658);
or U3482 (N_3482,In_1251,In_678);
xor U3483 (N_3483,In_1091,In_1261);
nand U3484 (N_3484,In_2241,In_932);
or U3485 (N_3485,In_1863,In_882);
or U3486 (N_3486,In_2899,In_475);
and U3487 (N_3487,In_1277,In_2616);
nor U3488 (N_3488,In_2449,In_2119);
nor U3489 (N_3489,In_803,In_1638);
nor U3490 (N_3490,In_2037,In_1685);
and U3491 (N_3491,In_2691,In_2378);
or U3492 (N_3492,In_1067,In_1362);
nor U3493 (N_3493,In_1492,In_2610);
nor U3494 (N_3494,In_1094,In_2067);
nand U3495 (N_3495,In_1585,In_2318);
or U3496 (N_3496,In_196,In_1899);
nand U3497 (N_3497,In_269,In_2326);
and U3498 (N_3498,In_859,In_1292);
nand U3499 (N_3499,In_2897,In_2457);
nand U3500 (N_3500,In_413,In_2375);
nand U3501 (N_3501,In_1781,In_1807);
nand U3502 (N_3502,In_2133,In_1030);
and U3503 (N_3503,In_767,In_2167);
or U3504 (N_3504,In_841,In_301);
nor U3505 (N_3505,In_1227,In_627);
nand U3506 (N_3506,In_2221,In_2401);
or U3507 (N_3507,In_1647,In_1175);
nand U3508 (N_3508,In_2349,In_825);
nor U3509 (N_3509,In_98,In_78);
nor U3510 (N_3510,In_626,In_1012);
nand U3511 (N_3511,In_533,In_658);
nand U3512 (N_3512,In_1857,In_2716);
or U3513 (N_3513,In_330,In_994);
nor U3514 (N_3514,In_356,In_1608);
or U3515 (N_3515,In_225,In_122);
or U3516 (N_3516,In_2532,In_2367);
or U3517 (N_3517,In_1235,In_823);
or U3518 (N_3518,In_2180,In_784);
and U3519 (N_3519,In_1847,In_669);
nor U3520 (N_3520,In_2630,In_193);
and U3521 (N_3521,In_1382,In_76);
nand U3522 (N_3522,In_2235,In_2342);
nor U3523 (N_3523,In_2212,In_1450);
and U3524 (N_3524,In_1845,In_194);
nor U3525 (N_3525,In_1741,In_1225);
nor U3526 (N_3526,In_1384,In_683);
or U3527 (N_3527,In_1365,In_2653);
and U3528 (N_3528,In_1025,In_1557);
nor U3529 (N_3529,In_2161,In_1944);
nor U3530 (N_3530,In_2739,In_192);
or U3531 (N_3531,In_1982,In_572);
nand U3532 (N_3532,In_315,In_1288);
or U3533 (N_3533,In_732,In_1699);
nor U3534 (N_3534,In_2132,In_501);
and U3535 (N_3535,In_2750,In_1412);
nand U3536 (N_3536,In_143,In_1553);
nand U3537 (N_3537,In_65,In_1565);
and U3538 (N_3538,In_456,In_2246);
or U3539 (N_3539,In_213,In_989);
and U3540 (N_3540,In_816,In_54);
xnor U3541 (N_3541,In_447,In_2742);
nand U3542 (N_3542,In_2276,In_1515);
nand U3543 (N_3543,In_2138,In_2883);
and U3544 (N_3544,In_496,In_1654);
nor U3545 (N_3545,In_115,In_305);
xor U3546 (N_3546,In_1232,In_907);
and U3547 (N_3547,In_2309,In_680);
or U3548 (N_3548,In_168,In_671);
or U3549 (N_3549,In_856,In_500);
and U3550 (N_3550,In_2665,In_359);
and U3551 (N_3551,In_1680,In_762);
or U3552 (N_3552,In_1013,In_690);
and U3553 (N_3553,In_2333,In_2920);
and U3554 (N_3554,In_2417,In_670);
and U3555 (N_3555,In_1880,In_2797);
or U3556 (N_3556,In_2758,In_1726);
or U3557 (N_3557,In_1894,In_1417);
or U3558 (N_3558,In_197,In_2914);
nor U3559 (N_3559,In_1362,In_1925);
nor U3560 (N_3560,In_470,In_986);
and U3561 (N_3561,In_2903,In_935);
nor U3562 (N_3562,In_1100,In_1593);
nand U3563 (N_3563,In_477,In_1264);
or U3564 (N_3564,In_1341,In_481);
or U3565 (N_3565,In_367,In_1997);
nor U3566 (N_3566,In_534,In_1116);
and U3567 (N_3567,In_2280,In_1799);
nand U3568 (N_3568,In_2396,In_437);
and U3569 (N_3569,In_1968,In_1340);
and U3570 (N_3570,In_100,In_2091);
or U3571 (N_3571,In_271,In_1840);
and U3572 (N_3572,In_206,In_2312);
and U3573 (N_3573,In_2045,In_2861);
nor U3574 (N_3574,In_2212,In_2964);
or U3575 (N_3575,In_1809,In_1199);
and U3576 (N_3576,In_2723,In_628);
xnor U3577 (N_3577,In_1114,In_676);
nand U3578 (N_3578,In_1270,In_2750);
and U3579 (N_3579,In_2368,In_1551);
nand U3580 (N_3580,In_2473,In_614);
and U3581 (N_3581,In_1185,In_2821);
or U3582 (N_3582,In_2172,In_2232);
nor U3583 (N_3583,In_226,In_499);
nor U3584 (N_3584,In_951,In_2455);
xor U3585 (N_3585,In_1055,In_1231);
nand U3586 (N_3586,In_1301,In_2431);
nor U3587 (N_3587,In_2855,In_417);
or U3588 (N_3588,In_1709,In_719);
nor U3589 (N_3589,In_1126,In_1731);
xnor U3590 (N_3590,In_2846,In_1706);
and U3591 (N_3591,In_2689,In_1215);
and U3592 (N_3592,In_1942,In_2095);
or U3593 (N_3593,In_488,In_2027);
nand U3594 (N_3594,In_1803,In_1003);
nand U3595 (N_3595,In_893,In_1619);
or U3596 (N_3596,In_2216,In_1253);
and U3597 (N_3597,In_1242,In_1253);
or U3598 (N_3598,In_432,In_1253);
or U3599 (N_3599,In_554,In_648);
nor U3600 (N_3600,In_1135,In_285);
nor U3601 (N_3601,In_1665,In_2619);
and U3602 (N_3602,In_1069,In_31);
xnor U3603 (N_3603,In_103,In_1619);
nand U3604 (N_3604,In_2119,In_175);
nor U3605 (N_3605,In_2164,In_2069);
nand U3606 (N_3606,In_1388,In_729);
nand U3607 (N_3607,In_1593,In_2659);
or U3608 (N_3608,In_571,In_2983);
xnor U3609 (N_3609,In_2796,In_2450);
and U3610 (N_3610,In_112,In_11);
nor U3611 (N_3611,In_1794,In_2042);
nand U3612 (N_3612,In_754,In_2233);
nor U3613 (N_3613,In_7,In_221);
or U3614 (N_3614,In_54,In_803);
xor U3615 (N_3615,In_2470,In_2778);
or U3616 (N_3616,In_2185,In_641);
or U3617 (N_3617,In_576,In_1474);
xnor U3618 (N_3618,In_2908,In_2297);
nor U3619 (N_3619,In_2736,In_310);
xnor U3620 (N_3620,In_1455,In_2289);
nand U3621 (N_3621,In_1113,In_1324);
or U3622 (N_3622,In_2693,In_1673);
or U3623 (N_3623,In_1213,In_2387);
nor U3624 (N_3624,In_2465,In_2490);
and U3625 (N_3625,In_32,In_2660);
xnor U3626 (N_3626,In_2210,In_356);
or U3627 (N_3627,In_2373,In_2543);
or U3628 (N_3628,In_1379,In_1662);
and U3629 (N_3629,In_1194,In_1169);
and U3630 (N_3630,In_63,In_771);
nand U3631 (N_3631,In_1016,In_1019);
and U3632 (N_3632,In_1083,In_1453);
or U3633 (N_3633,In_880,In_1725);
xor U3634 (N_3634,In_1566,In_2592);
nand U3635 (N_3635,In_2960,In_2303);
or U3636 (N_3636,In_2497,In_1574);
or U3637 (N_3637,In_2563,In_1402);
and U3638 (N_3638,In_929,In_2046);
and U3639 (N_3639,In_366,In_2635);
xnor U3640 (N_3640,In_2591,In_2767);
or U3641 (N_3641,In_1266,In_2265);
and U3642 (N_3642,In_439,In_281);
xnor U3643 (N_3643,In_950,In_2482);
or U3644 (N_3644,In_1712,In_1166);
nand U3645 (N_3645,In_1832,In_377);
nand U3646 (N_3646,In_476,In_2623);
and U3647 (N_3647,In_1835,In_2662);
xnor U3648 (N_3648,In_1376,In_3);
nor U3649 (N_3649,In_720,In_1499);
or U3650 (N_3650,In_2961,In_1231);
nor U3651 (N_3651,In_2731,In_1704);
and U3652 (N_3652,In_1389,In_368);
nor U3653 (N_3653,In_81,In_895);
nor U3654 (N_3654,In_882,In_2305);
nand U3655 (N_3655,In_1284,In_2253);
xor U3656 (N_3656,In_620,In_368);
nand U3657 (N_3657,In_1179,In_1031);
and U3658 (N_3658,In_2605,In_2625);
nand U3659 (N_3659,In_303,In_2526);
nor U3660 (N_3660,In_2847,In_311);
and U3661 (N_3661,In_1816,In_316);
nand U3662 (N_3662,In_319,In_1087);
nand U3663 (N_3663,In_1747,In_443);
nor U3664 (N_3664,In_2637,In_1081);
or U3665 (N_3665,In_4,In_427);
or U3666 (N_3666,In_1031,In_2858);
nand U3667 (N_3667,In_643,In_1528);
nor U3668 (N_3668,In_2519,In_66);
nor U3669 (N_3669,In_1167,In_1055);
and U3670 (N_3670,In_896,In_2697);
nor U3671 (N_3671,In_804,In_1952);
nor U3672 (N_3672,In_2930,In_978);
xnor U3673 (N_3673,In_2828,In_148);
nand U3674 (N_3674,In_1063,In_919);
nand U3675 (N_3675,In_1829,In_247);
nand U3676 (N_3676,In_2587,In_1431);
and U3677 (N_3677,In_1106,In_396);
and U3678 (N_3678,In_2440,In_1517);
or U3679 (N_3679,In_65,In_299);
nand U3680 (N_3680,In_2511,In_1834);
xnor U3681 (N_3681,In_1483,In_2027);
or U3682 (N_3682,In_2044,In_1045);
or U3683 (N_3683,In_444,In_2452);
nor U3684 (N_3684,In_880,In_1265);
xor U3685 (N_3685,In_1461,In_2051);
or U3686 (N_3686,In_590,In_1870);
and U3687 (N_3687,In_328,In_2293);
nand U3688 (N_3688,In_1059,In_1383);
nand U3689 (N_3689,In_2305,In_215);
nand U3690 (N_3690,In_90,In_1375);
or U3691 (N_3691,In_459,In_1237);
xor U3692 (N_3692,In_46,In_596);
or U3693 (N_3693,In_24,In_2552);
nand U3694 (N_3694,In_443,In_2975);
nand U3695 (N_3695,In_414,In_212);
or U3696 (N_3696,In_2229,In_2216);
nor U3697 (N_3697,In_2213,In_547);
and U3698 (N_3698,In_231,In_75);
xnor U3699 (N_3699,In_362,In_570);
nor U3700 (N_3700,In_1393,In_830);
or U3701 (N_3701,In_1085,In_2593);
nand U3702 (N_3702,In_1937,In_1071);
or U3703 (N_3703,In_2514,In_509);
or U3704 (N_3704,In_512,In_151);
xnor U3705 (N_3705,In_2295,In_2168);
nand U3706 (N_3706,In_137,In_1901);
or U3707 (N_3707,In_1009,In_2106);
and U3708 (N_3708,In_193,In_1176);
nor U3709 (N_3709,In_24,In_2708);
and U3710 (N_3710,In_586,In_2566);
and U3711 (N_3711,In_216,In_919);
and U3712 (N_3712,In_1180,In_1889);
nor U3713 (N_3713,In_1917,In_1283);
nand U3714 (N_3714,In_2502,In_2739);
or U3715 (N_3715,In_526,In_2118);
nor U3716 (N_3716,In_964,In_718);
or U3717 (N_3717,In_484,In_1036);
nand U3718 (N_3718,In_816,In_108);
nand U3719 (N_3719,In_2315,In_1743);
or U3720 (N_3720,In_781,In_549);
and U3721 (N_3721,In_732,In_2296);
and U3722 (N_3722,In_1760,In_901);
and U3723 (N_3723,In_2304,In_96);
and U3724 (N_3724,In_2508,In_2878);
and U3725 (N_3725,In_1126,In_509);
nand U3726 (N_3726,In_2958,In_2130);
nand U3727 (N_3727,In_2367,In_2861);
or U3728 (N_3728,In_124,In_782);
nor U3729 (N_3729,In_2747,In_2032);
or U3730 (N_3730,In_2492,In_37);
nor U3731 (N_3731,In_2022,In_867);
nand U3732 (N_3732,In_814,In_740);
or U3733 (N_3733,In_2022,In_1908);
or U3734 (N_3734,In_2843,In_1533);
nand U3735 (N_3735,In_1448,In_989);
nor U3736 (N_3736,In_2572,In_913);
nor U3737 (N_3737,In_2787,In_20);
nor U3738 (N_3738,In_206,In_300);
nand U3739 (N_3739,In_651,In_1376);
nor U3740 (N_3740,In_450,In_745);
and U3741 (N_3741,In_2021,In_2518);
nand U3742 (N_3742,In_1812,In_1816);
nand U3743 (N_3743,In_638,In_846);
or U3744 (N_3744,In_948,In_433);
nor U3745 (N_3745,In_1464,In_979);
nor U3746 (N_3746,In_2235,In_2565);
nand U3747 (N_3747,In_2700,In_786);
and U3748 (N_3748,In_225,In_1842);
and U3749 (N_3749,In_2879,In_1516);
nor U3750 (N_3750,In_1269,In_2540);
nor U3751 (N_3751,In_2964,In_2566);
nand U3752 (N_3752,In_2258,In_2699);
and U3753 (N_3753,In_2696,In_687);
and U3754 (N_3754,In_2396,In_2753);
and U3755 (N_3755,In_1588,In_1438);
and U3756 (N_3756,In_627,In_863);
xnor U3757 (N_3757,In_2786,In_2443);
or U3758 (N_3758,In_1860,In_2683);
xnor U3759 (N_3759,In_1758,In_541);
nand U3760 (N_3760,In_1966,In_2049);
and U3761 (N_3761,In_1824,In_1602);
nand U3762 (N_3762,In_457,In_2612);
nand U3763 (N_3763,In_1135,In_202);
nor U3764 (N_3764,In_564,In_1654);
and U3765 (N_3765,In_616,In_1144);
and U3766 (N_3766,In_1102,In_1367);
nand U3767 (N_3767,In_590,In_834);
or U3768 (N_3768,In_2977,In_1111);
or U3769 (N_3769,In_2870,In_1215);
or U3770 (N_3770,In_20,In_479);
and U3771 (N_3771,In_1920,In_1108);
and U3772 (N_3772,In_2283,In_2741);
and U3773 (N_3773,In_1017,In_641);
nor U3774 (N_3774,In_537,In_240);
or U3775 (N_3775,In_1435,In_989);
or U3776 (N_3776,In_663,In_559);
and U3777 (N_3777,In_2287,In_1205);
or U3778 (N_3778,In_2549,In_1755);
xnor U3779 (N_3779,In_2355,In_2459);
and U3780 (N_3780,In_2113,In_1201);
nand U3781 (N_3781,In_904,In_1150);
xnor U3782 (N_3782,In_2857,In_772);
xor U3783 (N_3783,In_444,In_2400);
xnor U3784 (N_3784,In_1183,In_922);
nor U3785 (N_3785,In_661,In_2707);
and U3786 (N_3786,In_2108,In_1584);
or U3787 (N_3787,In_1,In_1361);
nand U3788 (N_3788,In_474,In_670);
nor U3789 (N_3789,In_114,In_1974);
nor U3790 (N_3790,In_848,In_2829);
or U3791 (N_3791,In_2869,In_999);
xor U3792 (N_3792,In_18,In_574);
or U3793 (N_3793,In_735,In_129);
nor U3794 (N_3794,In_1718,In_1907);
nor U3795 (N_3795,In_1984,In_1940);
or U3796 (N_3796,In_2217,In_2616);
nor U3797 (N_3797,In_2192,In_420);
nor U3798 (N_3798,In_2543,In_1473);
nor U3799 (N_3799,In_1474,In_1341);
xor U3800 (N_3800,In_209,In_2615);
or U3801 (N_3801,In_868,In_61);
nand U3802 (N_3802,In_1120,In_2532);
xnor U3803 (N_3803,In_907,In_822);
nor U3804 (N_3804,In_753,In_1538);
xnor U3805 (N_3805,In_1356,In_1060);
or U3806 (N_3806,In_2427,In_406);
or U3807 (N_3807,In_2308,In_1255);
and U3808 (N_3808,In_876,In_2039);
or U3809 (N_3809,In_15,In_1954);
or U3810 (N_3810,In_2990,In_284);
or U3811 (N_3811,In_1399,In_2413);
and U3812 (N_3812,In_2411,In_299);
and U3813 (N_3813,In_667,In_2949);
nand U3814 (N_3814,In_2374,In_2977);
nor U3815 (N_3815,In_1406,In_358);
nor U3816 (N_3816,In_93,In_2936);
or U3817 (N_3817,In_2507,In_1657);
and U3818 (N_3818,In_1579,In_211);
and U3819 (N_3819,In_2273,In_1929);
nor U3820 (N_3820,In_787,In_1006);
or U3821 (N_3821,In_390,In_2623);
or U3822 (N_3822,In_2765,In_357);
xnor U3823 (N_3823,In_16,In_2321);
nand U3824 (N_3824,In_239,In_1611);
or U3825 (N_3825,In_2354,In_171);
and U3826 (N_3826,In_2319,In_1731);
or U3827 (N_3827,In_2758,In_2875);
nor U3828 (N_3828,In_570,In_2254);
nand U3829 (N_3829,In_288,In_912);
nand U3830 (N_3830,In_2954,In_714);
or U3831 (N_3831,In_1121,In_1268);
xnor U3832 (N_3832,In_2216,In_1122);
or U3833 (N_3833,In_2434,In_1641);
nand U3834 (N_3834,In_7,In_641);
xor U3835 (N_3835,In_2582,In_1371);
nand U3836 (N_3836,In_1951,In_2060);
or U3837 (N_3837,In_1383,In_331);
nand U3838 (N_3838,In_2726,In_325);
and U3839 (N_3839,In_1512,In_661);
nor U3840 (N_3840,In_942,In_535);
and U3841 (N_3841,In_2850,In_977);
or U3842 (N_3842,In_2535,In_695);
nand U3843 (N_3843,In_1350,In_550);
nor U3844 (N_3844,In_333,In_2798);
nand U3845 (N_3845,In_1719,In_935);
nand U3846 (N_3846,In_302,In_2278);
nor U3847 (N_3847,In_2084,In_2733);
xnor U3848 (N_3848,In_2893,In_2064);
nor U3849 (N_3849,In_646,In_2938);
and U3850 (N_3850,In_137,In_1514);
nand U3851 (N_3851,In_1957,In_1918);
nand U3852 (N_3852,In_1754,In_1776);
xnor U3853 (N_3853,In_2839,In_665);
nor U3854 (N_3854,In_1309,In_586);
nor U3855 (N_3855,In_1585,In_1414);
xnor U3856 (N_3856,In_1539,In_623);
nand U3857 (N_3857,In_127,In_1671);
xnor U3858 (N_3858,In_1952,In_2853);
and U3859 (N_3859,In_2047,In_1953);
or U3860 (N_3860,In_1498,In_2151);
xor U3861 (N_3861,In_1847,In_1823);
nor U3862 (N_3862,In_221,In_218);
nand U3863 (N_3863,In_2613,In_2922);
nor U3864 (N_3864,In_578,In_1942);
or U3865 (N_3865,In_597,In_901);
nand U3866 (N_3866,In_2838,In_645);
or U3867 (N_3867,In_232,In_468);
or U3868 (N_3868,In_2017,In_706);
or U3869 (N_3869,In_385,In_1692);
and U3870 (N_3870,In_2565,In_2849);
and U3871 (N_3871,In_1936,In_806);
nand U3872 (N_3872,In_1280,In_1935);
and U3873 (N_3873,In_2707,In_2727);
nor U3874 (N_3874,In_2070,In_2128);
nand U3875 (N_3875,In_1667,In_2609);
nor U3876 (N_3876,In_104,In_2685);
nand U3877 (N_3877,In_546,In_2615);
or U3878 (N_3878,In_2195,In_2932);
or U3879 (N_3879,In_2693,In_2470);
nor U3880 (N_3880,In_2494,In_2376);
nor U3881 (N_3881,In_703,In_2605);
nor U3882 (N_3882,In_1770,In_2162);
or U3883 (N_3883,In_1094,In_404);
nand U3884 (N_3884,In_2736,In_2020);
nand U3885 (N_3885,In_2193,In_1723);
nand U3886 (N_3886,In_2814,In_696);
nor U3887 (N_3887,In_2209,In_2089);
nor U3888 (N_3888,In_1400,In_2133);
xor U3889 (N_3889,In_1634,In_431);
nor U3890 (N_3890,In_1942,In_2936);
nand U3891 (N_3891,In_2604,In_1326);
xor U3892 (N_3892,In_1967,In_1859);
or U3893 (N_3893,In_2534,In_2416);
nand U3894 (N_3894,In_1228,In_395);
nor U3895 (N_3895,In_604,In_1038);
nor U3896 (N_3896,In_2601,In_2388);
nand U3897 (N_3897,In_1456,In_2041);
nand U3898 (N_3898,In_50,In_993);
or U3899 (N_3899,In_2338,In_2907);
nand U3900 (N_3900,In_1007,In_2925);
xor U3901 (N_3901,In_1067,In_1249);
nand U3902 (N_3902,In_1302,In_324);
nor U3903 (N_3903,In_1258,In_1227);
nor U3904 (N_3904,In_1487,In_827);
or U3905 (N_3905,In_2705,In_2891);
and U3906 (N_3906,In_2643,In_2700);
nand U3907 (N_3907,In_2112,In_1774);
nor U3908 (N_3908,In_2807,In_2514);
and U3909 (N_3909,In_1415,In_1787);
nor U3910 (N_3910,In_1502,In_639);
nor U3911 (N_3911,In_1535,In_347);
nor U3912 (N_3912,In_2289,In_523);
nand U3913 (N_3913,In_700,In_744);
nor U3914 (N_3914,In_1882,In_2286);
nor U3915 (N_3915,In_2003,In_1955);
nor U3916 (N_3916,In_2061,In_2717);
nor U3917 (N_3917,In_2315,In_683);
and U3918 (N_3918,In_973,In_1142);
or U3919 (N_3919,In_1127,In_2947);
or U3920 (N_3920,In_801,In_669);
nor U3921 (N_3921,In_1653,In_596);
nor U3922 (N_3922,In_491,In_946);
and U3923 (N_3923,In_584,In_2521);
nand U3924 (N_3924,In_1756,In_457);
nor U3925 (N_3925,In_1813,In_1401);
nand U3926 (N_3926,In_730,In_618);
xor U3927 (N_3927,In_494,In_305);
nand U3928 (N_3928,In_2691,In_778);
nor U3929 (N_3929,In_775,In_597);
and U3930 (N_3930,In_2233,In_2520);
nor U3931 (N_3931,In_618,In_777);
and U3932 (N_3932,In_2699,In_2195);
or U3933 (N_3933,In_1590,In_2459);
and U3934 (N_3934,In_969,In_178);
or U3935 (N_3935,In_43,In_1321);
nand U3936 (N_3936,In_1882,In_52);
or U3937 (N_3937,In_132,In_103);
nor U3938 (N_3938,In_1445,In_464);
and U3939 (N_3939,In_2715,In_2168);
and U3940 (N_3940,In_1576,In_757);
nor U3941 (N_3941,In_2011,In_2369);
nor U3942 (N_3942,In_55,In_1510);
xor U3943 (N_3943,In_269,In_2559);
or U3944 (N_3944,In_1108,In_643);
nor U3945 (N_3945,In_102,In_1754);
nor U3946 (N_3946,In_2524,In_1504);
nor U3947 (N_3947,In_1440,In_1229);
nand U3948 (N_3948,In_2695,In_1722);
nor U3949 (N_3949,In_916,In_1062);
nor U3950 (N_3950,In_1320,In_506);
nand U3951 (N_3951,In_2806,In_1284);
nor U3952 (N_3952,In_1107,In_2296);
nor U3953 (N_3953,In_1117,In_2465);
nor U3954 (N_3954,In_2962,In_589);
and U3955 (N_3955,In_1291,In_2786);
and U3956 (N_3956,In_366,In_2247);
and U3957 (N_3957,In_1555,In_1498);
or U3958 (N_3958,In_125,In_1334);
nand U3959 (N_3959,In_1685,In_167);
nand U3960 (N_3960,In_1766,In_1032);
and U3961 (N_3961,In_1427,In_693);
or U3962 (N_3962,In_2497,In_955);
nor U3963 (N_3963,In_2501,In_1060);
or U3964 (N_3964,In_337,In_1199);
nor U3965 (N_3965,In_338,In_1934);
xnor U3966 (N_3966,In_2339,In_2080);
nand U3967 (N_3967,In_605,In_1020);
nor U3968 (N_3968,In_2846,In_2437);
nand U3969 (N_3969,In_1587,In_2056);
or U3970 (N_3970,In_2099,In_1842);
nor U3971 (N_3971,In_2390,In_768);
xnor U3972 (N_3972,In_1065,In_9);
nand U3973 (N_3973,In_1156,In_102);
nand U3974 (N_3974,In_83,In_673);
or U3975 (N_3975,In_1983,In_1757);
nand U3976 (N_3976,In_2969,In_2415);
or U3977 (N_3977,In_1566,In_278);
and U3978 (N_3978,In_2047,In_1382);
nand U3979 (N_3979,In_2078,In_2065);
nand U3980 (N_3980,In_2370,In_2057);
or U3981 (N_3981,In_1411,In_1479);
nand U3982 (N_3982,In_2541,In_308);
xor U3983 (N_3983,In_942,In_2616);
and U3984 (N_3984,In_646,In_2350);
or U3985 (N_3985,In_649,In_2550);
and U3986 (N_3986,In_165,In_1812);
nor U3987 (N_3987,In_1765,In_2311);
nand U3988 (N_3988,In_893,In_1649);
nand U3989 (N_3989,In_1536,In_794);
and U3990 (N_3990,In_322,In_575);
and U3991 (N_3991,In_2375,In_2825);
and U3992 (N_3992,In_603,In_644);
xnor U3993 (N_3993,In_66,In_1419);
xnor U3994 (N_3994,In_847,In_535);
or U3995 (N_3995,In_1537,In_143);
nand U3996 (N_3996,In_554,In_1365);
or U3997 (N_3997,In_2230,In_317);
and U3998 (N_3998,In_562,In_957);
or U3999 (N_3999,In_2079,In_2695);
nand U4000 (N_4000,In_2638,In_1184);
and U4001 (N_4001,In_2899,In_2102);
nor U4002 (N_4002,In_309,In_1887);
nand U4003 (N_4003,In_295,In_2663);
or U4004 (N_4004,In_553,In_928);
nor U4005 (N_4005,In_2486,In_2075);
nand U4006 (N_4006,In_1721,In_2519);
and U4007 (N_4007,In_1516,In_960);
or U4008 (N_4008,In_2934,In_1367);
and U4009 (N_4009,In_1700,In_1973);
nand U4010 (N_4010,In_2428,In_2136);
and U4011 (N_4011,In_197,In_250);
and U4012 (N_4012,In_2727,In_797);
nor U4013 (N_4013,In_2888,In_889);
and U4014 (N_4014,In_1646,In_1368);
nand U4015 (N_4015,In_2379,In_2052);
nand U4016 (N_4016,In_354,In_356);
or U4017 (N_4017,In_1954,In_1303);
nand U4018 (N_4018,In_806,In_1886);
and U4019 (N_4019,In_1945,In_2686);
and U4020 (N_4020,In_200,In_2884);
nor U4021 (N_4021,In_1091,In_2484);
nor U4022 (N_4022,In_2558,In_205);
or U4023 (N_4023,In_1764,In_1854);
and U4024 (N_4024,In_1648,In_2007);
nor U4025 (N_4025,In_2425,In_2783);
or U4026 (N_4026,In_161,In_1296);
nor U4027 (N_4027,In_1255,In_1230);
and U4028 (N_4028,In_129,In_108);
and U4029 (N_4029,In_2131,In_2845);
and U4030 (N_4030,In_2376,In_188);
or U4031 (N_4031,In_1377,In_2046);
nor U4032 (N_4032,In_410,In_91);
nand U4033 (N_4033,In_2987,In_1996);
or U4034 (N_4034,In_655,In_852);
nor U4035 (N_4035,In_1171,In_2091);
nand U4036 (N_4036,In_781,In_2927);
and U4037 (N_4037,In_2917,In_1500);
xnor U4038 (N_4038,In_2254,In_2093);
and U4039 (N_4039,In_1980,In_2130);
nor U4040 (N_4040,In_1487,In_2498);
or U4041 (N_4041,In_482,In_2768);
nor U4042 (N_4042,In_2655,In_1518);
nand U4043 (N_4043,In_2489,In_2664);
nor U4044 (N_4044,In_946,In_2894);
or U4045 (N_4045,In_2867,In_1282);
nand U4046 (N_4046,In_550,In_2540);
nand U4047 (N_4047,In_2761,In_1271);
and U4048 (N_4048,In_2168,In_2205);
or U4049 (N_4049,In_1778,In_769);
nand U4050 (N_4050,In_2389,In_552);
nand U4051 (N_4051,In_130,In_174);
nor U4052 (N_4052,In_1745,In_1571);
or U4053 (N_4053,In_1576,In_2487);
or U4054 (N_4054,In_998,In_1762);
or U4055 (N_4055,In_1000,In_2645);
xor U4056 (N_4056,In_2883,In_2713);
nand U4057 (N_4057,In_2403,In_2544);
nor U4058 (N_4058,In_1430,In_1559);
and U4059 (N_4059,In_1693,In_1600);
and U4060 (N_4060,In_1513,In_464);
and U4061 (N_4061,In_876,In_1039);
xor U4062 (N_4062,In_1130,In_375);
nor U4063 (N_4063,In_1006,In_703);
and U4064 (N_4064,In_2027,In_875);
nand U4065 (N_4065,In_2038,In_1883);
or U4066 (N_4066,In_1872,In_1224);
or U4067 (N_4067,In_796,In_2871);
nor U4068 (N_4068,In_327,In_1090);
and U4069 (N_4069,In_1631,In_769);
nor U4070 (N_4070,In_2775,In_1194);
xor U4071 (N_4071,In_518,In_2137);
or U4072 (N_4072,In_2501,In_2561);
or U4073 (N_4073,In_2355,In_1952);
nand U4074 (N_4074,In_1211,In_1717);
nand U4075 (N_4075,In_1111,In_850);
nor U4076 (N_4076,In_451,In_1016);
nor U4077 (N_4077,In_2767,In_1583);
nor U4078 (N_4078,In_307,In_2556);
and U4079 (N_4079,In_1589,In_2233);
nor U4080 (N_4080,In_2745,In_902);
nand U4081 (N_4081,In_188,In_2947);
and U4082 (N_4082,In_1006,In_535);
nor U4083 (N_4083,In_1497,In_2313);
nor U4084 (N_4084,In_1160,In_1268);
nand U4085 (N_4085,In_973,In_2285);
nand U4086 (N_4086,In_2871,In_987);
nand U4087 (N_4087,In_654,In_1372);
xor U4088 (N_4088,In_1932,In_433);
and U4089 (N_4089,In_1061,In_1954);
and U4090 (N_4090,In_325,In_2412);
nor U4091 (N_4091,In_520,In_970);
nor U4092 (N_4092,In_2612,In_54);
or U4093 (N_4093,In_2128,In_769);
or U4094 (N_4094,In_1238,In_1933);
and U4095 (N_4095,In_1019,In_1646);
or U4096 (N_4096,In_368,In_768);
xor U4097 (N_4097,In_2884,In_1380);
nor U4098 (N_4098,In_2129,In_2136);
and U4099 (N_4099,In_612,In_111);
nand U4100 (N_4100,In_47,In_1726);
nor U4101 (N_4101,In_1518,In_2422);
and U4102 (N_4102,In_780,In_847);
and U4103 (N_4103,In_926,In_609);
or U4104 (N_4104,In_2622,In_879);
or U4105 (N_4105,In_2735,In_659);
nor U4106 (N_4106,In_953,In_913);
or U4107 (N_4107,In_1117,In_1030);
and U4108 (N_4108,In_2304,In_2476);
or U4109 (N_4109,In_539,In_2937);
nand U4110 (N_4110,In_2423,In_1721);
nor U4111 (N_4111,In_159,In_1415);
and U4112 (N_4112,In_2716,In_1882);
nand U4113 (N_4113,In_2736,In_567);
xor U4114 (N_4114,In_1553,In_115);
nor U4115 (N_4115,In_558,In_165);
or U4116 (N_4116,In_2051,In_1758);
or U4117 (N_4117,In_331,In_189);
nor U4118 (N_4118,In_767,In_543);
and U4119 (N_4119,In_580,In_89);
nor U4120 (N_4120,In_971,In_1062);
nand U4121 (N_4121,In_347,In_525);
or U4122 (N_4122,In_2794,In_1660);
and U4123 (N_4123,In_1927,In_1940);
nor U4124 (N_4124,In_2037,In_2649);
nor U4125 (N_4125,In_1898,In_1224);
xor U4126 (N_4126,In_1536,In_886);
and U4127 (N_4127,In_2494,In_2234);
or U4128 (N_4128,In_1435,In_2692);
nand U4129 (N_4129,In_657,In_1472);
and U4130 (N_4130,In_290,In_1053);
nand U4131 (N_4131,In_2304,In_1373);
or U4132 (N_4132,In_180,In_750);
nor U4133 (N_4133,In_792,In_420);
and U4134 (N_4134,In_2989,In_2386);
and U4135 (N_4135,In_304,In_1198);
xor U4136 (N_4136,In_2963,In_2352);
nor U4137 (N_4137,In_64,In_1023);
nand U4138 (N_4138,In_502,In_1328);
and U4139 (N_4139,In_430,In_2922);
nor U4140 (N_4140,In_807,In_1559);
or U4141 (N_4141,In_415,In_447);
nor U4142 (N_4142,In_1678,In_1040);
xor U4143 (N_4143,In_1850,In_2746);
and U4144 (N_4144,In_817,In_386);
and U4145 (N_4145,In_2201,In_2703);
nor U4146 (N_4146,In_2666,In_1948);
or U4147 (N_4147,In_2123,In_1322);
nand U4148 (N_4148,In_478,In_2648);
nor U4149 (N_4149,In_2149,In_2678);
xnor U4150 (N_4150,In_1063,In_775);
nor U4151 (N_4151,In_2195,In_277);
or U4152 (N_4152,In_2406,In_2642);
or U4153 (N_4153,In_145,In_1715);
xnor U4154 (N_4154,In_62,In_1342);
or U4155 (N_4155,In_965,In_2869);
nor U4156 (N_4156,In_89,In_2228);
nor U4157 (N_4157,In_642,In_718);
and U4158 (N_4158,In_1182,In_2760);
nand U4159 (N_4159,In_803,In_430);
and U4160 (N_4160,In_2024,In_2467);
nand U4161 (N_4161,In_1887,In_604);
and U4162 (N_4162,In_2379,In_999);
and U4163 (N_4163,In_1887,In_477);
nand U4164 (N_4164,In_296,In_218);
nand U4165 (N_4165,In_2825,In_789);
or U4166 (N_4166,In_2353,In_2119);
nor U4167 (N_4167,In_1041,In_2579);
xor U4168 (N_4168,In_865,In_285);
or U4169 (N_4169,In_137,In_2630);
or U4170 (N_4170,In_1298,In_97);
nor U4171 (N_4171,In_2803,In_2073);
and U4172 (N_4172,In_2942,In_2042);
and U4173 (N_4173,In_2641,In_1452);
and U4174 (N_4174,In_554,In_2709);
or U4175 (N_4175,In_2489,In_2552);
xor U4176 (N_4176,In_2029,In_88);
and U4177 (N_4177,In_156,In_2429);
and U4178 (N_4178,In_2037,In_1361);
nand U4179 (N_4179,In_501,In_968);
nand U4180 (N_4180,In_958,In_2156);
and U4181 (N_4181,In_2594,In_1150);
and U4182 (N_4182,In_114,In_1985);
nor U4183 (N_4183,In_2947,In_927);
xor U4184 (N_4184,In_1131,In_1927);
nor U4185 (N_4185,In_254,In_467);
or U4186 (N_4186,In_96,In_633);
nor U4187 (N_4187,In_2126,In_2413);
nand U4188 (N_4188,In_915,In_1397);
nand U4189 (N_4189,In_718,In_2546);
nand U4190 (N_4190,In_1194,In_2940);
and U4191 (N_4191,In_839,In_923);
nor U4192 (N_4192,In_74,In_759);
nand U4193 (N_4193,In_148,In_1047);
nor U4194 (N_4194,In_2176,In_878);
xor U4195 (N_4195,In_1749,In_1334);
and U4196 (N_4196,In_2071,In_275);
nor U4197 (N_4197,In_2617,In_2038);
and U4198 (N_4198,In_2293,In_2176);
nand U4199 (N_4199,In_1556,In_1533);
nor U4200 (N_4200,In_1949,In_965);
or U4201 (N_4201,In_725,In_1738);
nor U4202 (N_4202,In_2005,In_700);
nor U4203 (N_4203,In_1582,In_1816);
xor U4204 (N_4204,In_461,In_2628);
and U4205 (N_4205,In_2255,In_1516);
nor U4206 (N_4206,In_886,In_1101);
xnor U4207 (N_4207,In_734,In_2307);
xor U4208 (N_4208,In_1961,In_468);
xnor U4209 (N_4209,In_2298,In_2834);
nor U4210 (N_4210,In_905,In_2750);
or U4211 (N_4211,In_2581,In_2311);
or U4212 (N_4212,In_2349,In_1652);
or U4213 (N_4213,In_2914,In_1085);
and U4214 (N_4214,In_1369,In_1668);
or U4215 (N_4215,In_2785,In_1245);
nand U4216 (N_4216,In_1385,In_741);
nand U4217 (N_4217,In_1776,In_143);
nor U4218 (N_4218,In_2555,In_2086);
or U4219 (N_4219,In_98,In_107);
xnor U4220 (N_4220,In_2317,In_1381);
nor U4221 (N_4221,In_161,In_259);
and U4222 (N_4222,In_1915,In_488);
and U4223 (N_4223,In_1553,In_2131);
or U4224 (N_4224,In_2056,In_2063);
nor U4225 (N_4225,In_895,In_1039);
and U4226 (N_4226,In_429,In_1637);
xor U4227 (N_4227,In_2073,In_2070);
xnor U4228 (N_4228,In_2884,In_1964);
nand U4229 (N_4229,In_2796,In_2848);
nand U4230 (N_4230,In_2955,In_2056);
or U4231 (N_4231,In_1786,In_489);
xor U4232 (N_4232,In_1589,In_483);
nand U4233 (N_4233,In_1506,In_843);
nor U4234 (N_4234,In_851,In_736);
nor U4235 (N_4235,In_1990,In_2857);
and U4236 (N_4236,In_2549,In_1690);
or U4237 (N_4237,In_1343,In_1413);
or U4238 (N_4238,In_499,In_1450);
or U4239 (N_4239,In_1773,In_2039);
nand U4240 (N_4240,In_2809,In_2686);
nor U4241 (N_4241,In_2920,In_1955);
nor U4242 (N_4242,In_2928,In_2443);
nor U4243 (N_4243,In_1309,In_2813);
nand U4244 (N_4244,In_1927,In_2699);
and U4245 (N_4245,In_2984,In_91);
and U4246 (N_4246,In_2314,In_2577);
nor U4247 (N_4247,In_2516,In_2457);
nor U4248 (N_4248,In_1686,In_637);
xnor U4249 (N_4249,In_1375,In_2633);
or U4250 (N_4250,In_1637,In_2139);
or U4251 (N_4251,In_2739,In_709);
or U4252 (N_4252,In_2653,In_2027);
or U4253 (N_4253,In_1593,In_1165);
nand U4254 (N_4254,In_1459,In_671);
nand U4255 (N_4255,In_1483,In_2167);
nand U4256 (N_4256,In_72,In_1265);
or U4257 (N_4257,In_977,In_637);
and U4258 (N_4258,In_1158,In_719);
or U4259 (N_4259,In_2760,In_1452);
or U4260 (N_4260,In_69,In_1921);
xnor U4261 (N_4261,In_2327,In_1613);
and U4262 (N_4262,In_1726,In_425);
and U4263 (N_4263,In_2091,In_368);
and U4264 (N_4264,In_1338,In_1654);
nor U4265 (N_4265,In_1644,In_2360);
or U4266 (N_4266,In_2153,In_40);
nor U4267 (N_4267,In_1056,In_1496);
nor U4268 (N_4268,In_1918,In_2208);
or U4269 (N_4269,In_2406,In_2719);
nor U4270 (N_4270,In_1925,In_297);
nand U4271 (N_4271,In_2994,In_2256);
and U4272 (N_4272,In_2163,In_1195);
or U4273 (N_4273,In_1778,In_761);
nor U4274 (N_4274,In_1973,In_823);
or U4275 (N_4275,In_655,In_519);
nor U4276 (N_4276,In_1079,In_1197);
xnor U4277 (N_4277,In_73,In_1913);
nand U4278 (N_4278,In_2371,In_686);
xor U4279 (N_4279,In_2179,In_1930);
and U4280 (N_4280,In_1162,In_1755);
or U4281 (N_4281,In_2742,In_1840);
nor U4282 (N_4282,In_476,In_2951);
nand U4283 (N_4283,In_1690,In_2166);
and U4284 (N_4284,In_1378,In_2120);
and U4285 (N_4285,In_207,In_2053);
nand U4286 (N_4286,In_2113,In_701);
and U4287 (N_4287,In_845,In_1607);
and U4288 (N_4288,In_1720,In_487);
nor U4289 (N_4289,In_1554,In_2578);
nand U4290 (N_4290,In_1404,In_1006);
nand U4291 (N_4291,In_2603,In_1521);
and U4292 (N_4292,In_1675,In_2598);
nor U4293 (N_4293,In_2429,In_1298);
xor U4294 (N_4294,In_2699,In_1215);
nand U4295 (N_4295,In_1106,In_804);
and U4296 (N_4296,In_1467,In_349);
nand U4297 (N_4297,In_1955,In_2459);
nand U4298 (N_4298,In_1358,In_2418);
nor U4299 (N_4299,In_1459,In_689);
nand U4300 (N_4300,In_848,In_2224);
nand U4301 (N_4301,In_2675,In_1568);
xnor U4302 (N_4302,In_1048,In_2410);
or U4303 (N_4303,In_2851,In_1193);
nand U4304 (N_4304,In_386,In_2685);
nand U4305 (N_4305,In_736,In_963);
nor U4306 (N_4306,In_2745,In_57);
nor U4307 (N_4307,In_775,In_2199);
and U4308 (N_4308,In_886,In_1541);
and U4309 (N_4309,In_2356,In_2206);
and U4310 (N_4310,In_589,In_938);
xor U4311 (N_4311,In_1842,In_1297);
nor U4312 (N_4312,In_1227,In_1916);
nand U4313 (N_4313,In_1839,In_1079);
and U4314 (N_4314,In_1830,In_24);
or U4315 (N_4315,In_712,In_125);
xor U4316 (N_4316,In_2739,In_200);
nand U4317 (N_4317,In_543,In_537);
nand U4318 (N_4318,In_1529,In_1901);
or U4319 (N_4319,In_1296,In_2747);
nand U4320 (N_4320,In_556,In_1633);
nand U4321 (N_4321,In_2932,In_1368);
nand U4322 (N_4322,In_1615,In_736);
and U4323 (N_4323,In_1056,In_2208);
nor U4324 (N_4324,In_1611,In_243);
or U4325 (N_4325,In_1963,In_2260);
nor U4326 (N_4326,In_2859,In_2850);
and U4327 (N_4327,In_1503,In_2662);
or U4328 (N_4328,In_1073,In_2553);
nand U4329 (N_4329,In_1179,In_95);
nor U4330 (N_4330,In_1272,In_164);
nor U4331 (N_4331,In_16,In_423);
xnor U4332 (N_4332,In_2758,In_553);
nor U4333 (N_4333,In_2893,In_2636);
nor U4334 (N_4334,In_2417,In_867);
or U4335 (N_4335,In_2662,In_2183);
and U4336 (N_4336,In_2812,In_2276);
or U4337 (N_4337,In_2631,In_2959);
xor U4338 (N_4338,In_2851,In_2749);
or U4339 (N_4339,In_2916,In_955);
or U4340 (N_4340,In_296,In_2948);
or U4341 (N_4341,In_2800,In_1212);
or U4342 (N_4342,In_1735,In_1455);
xnor U4343 (N_4343,In_1176,In_666);
nor U4344 (N_4344,In_317,In_1871);
and U4345 (N_4345,In_916,In_1797);
and U4346 (N_4346,In_1677,In_1621);
nand U4347 (N_4347,In_2651,In_2611);
nor U4348 (N_4348,In_1623,In_962);
and U4349 (N_4349,In_1150,In_111);
xor U4350 (N_4350,In_1991,In_1620);
or U4351 (N_4351,In_2900,In_1722);
nor U4352 (N_4352,In_105,In_1078);
and U4353 (N_4353,In_2723,In_2276);
and U4354 (N_4354,In_2009,In_677);
or U4355 (N_4355,In_2232,In_1867);
nand U4356 (N_4356,In_1222,In_426);
nor U4357 (N_4357,In_2172,In_1953);
nand U4358 (N_4358,In_122,In_2294);
nand U4359 (N_4359,In_1731,In_2136);
xnor U4360 (N_4360,In_1616,In_797);
nor U4361 (N_4361,In_1278,In_1908);
nor U4362 (N_4362,In_502,In_2403);
nand U4363 (N_4363,In_360,In_1280);
and U4364 (N_4364,In_780,In_854);
or U4365 (N_4365,In_135,In_879);
or U4366 (N_4366,In_2452,In_1896);
nand U4367 (N_4367,In_934,In_2468);
and U4368 (N_4368,In_2159,In_1596);
and U4369 (N_4369,In_20,In_1309);
and U4370 (N_4370,In_1145,In_1855);
xor U4371 (N_4371,In_2043,In_1905);
nor U4372 (N_4372,In_854,In_2672);
nor U4373 (N_4373,In_2373,In_2255);
xnor U4374 (N_4374,In_2027,In_2111);
nor U4375 (N_4375,In_695,In_1524);
and U4376 (N_4376,In_558,In_990);
or U4377 (N_4377,In_2644,In_1413);
nor U4378 (N_4378,In_2171,In_922);
nand U4379 (N_4379,In_1018,In_2214);
or U4380 (N_4380,In_1093,In_2082);
and U4381 (N_4381,In_2380,In_2744);
and U4382 (N_4382,In_757,In_1649);
and U4383 (N_4383,In_362,In_1764);
nand U4384 (N_4384,In_1950,In_2992);
nand U4385 (N_4385,In_1651,In_1523);
nor U4386 (N_4386,In_1901,In_1972);
or U4387 (N_4387,In_931,In_2385);
or U4388 (N_4388,In_2530,In_1070);
xor U4389 (N_4389,In_1204,In_42);
and U4390 (N_4390,In_1862,In_2693);
and U4391 (N_4391,In_202,In_2890);
nand U4392 (N_4392,In_1644,In_2920);
nand U4393 (N_4393,In_1417,In_1015);
nand U4394 (N_4394,In_803,In_70);
nand U4395 (N_4395,In_832,In_741);
and U4396 (N_4396,In_1878,In_710);
nor U4397 (N_4397,In_1626,In_1432);
or U4398 (N_4398,In_1108,In_2591);
or U4399 (N_4399,In_568,In_1572);
and U4400 (N_4400,In_733,In_159);
or U4401 (N_4401,In_2542,In_2120);
nor U4402 (N_4402,In_2160,In_849);
or U4403 (N_4403,In_1324,In_2805);
nor U4404 (N_4404,In_1696,In_2658);
and U4405 (N_4405,In_1031,In_1159);
and U4406 (N_4406,In_1090,In_931);
nand U4407 (N_4407,In_2276,In_821);
nor U4408 (N_4408,In_840,In_2421);
nor U4409 (N_4409,In_2673,In_324);
nand U4410 (N_4410,In_470,In_361);
nand U4411 (N_4411,In_287,In_1436);
or U4412 (N_4412,In_1653,In_1227);
nor U4413 (N_4413,In_1864,In_369);
nand U4414 (N_4414,In_1702,In_881);
and U4415 (N_4415,In_1779,In_2490);
and U4416 (N_4416,In_1448,In_501);
nor U4417 (N_4417,In_1695,In_1261);
or U4418 (N_4418,In_2173,In_323);
and U4419 (N_4419,In_2957,In_1230);
xor U4420 (N_4420,In_567,In_1806);
nand U4421 (N_4421,In_367,In_1528);
nor U4422 (N_4422,In_1285,In_1807);
nand U4423 (N_4423,In_993,In_2339);
and U4424 (N_4424,In_2897,In_1412);
and U4425 (N_4425,In_1637,In_160);
nor U4426 (N_4426,In_2819,In_310);
or U4427 (N_4427,In_1386,In_847);
or U4428 (N_4428,In_829,In_1079);
or U4429 (N_4429,In_2276,In_1874);
or U4430 (N_4430,In_1745,In_433);
and U4431 (N_4431,In_2157,In_2782);
and U4432 (N_4432,In_703,In_45);
or U4433 (N_4433,In_2900,In_506);
nand U4434 (N_4434,In_825,In_1266);
or U4435 (N_4435,In_519,In_904);
nor U4436 (N_4436,In_825,In_996);
or U4437 (N_4437,In_316,In_1856);
and U4438 (N_4438,In_1618,In_2935);
nor U4439 (N_4439,In_2473,In_2177);
and U4440 (N_4440,In_499,In_1161);
or U4441 (N_4441,In_2427,In_444);
nand U4442 (N_4442,In_2988,In_460);
or U4443 (N_4443,In_2141,In_1463);
nand U4444 (N_4444,In_2809,In_41);
or U4445 (N_4445,In_1657,In_2395);
or U4446 (N_4446,In_677,In_767);
nor U4447 (N_4447,In_2331,In_1420);
or U4448 (N_4448,In_1498,In_2087);
and U4449 (N_4449,In_2627,In_830);
xor U4450 (N_4450,In_940,In_918);
nand U4451 (N_4451,In_1281,In_1024);
nand U4452 (N_4452,In_2512,In_2067);
nor U4453 (N_4453,In_1629,In_1336);
nand U4454 (N_4454,In_2673,In_691);
nor U4455 (N_4455,In_1580,In_1177);
xnor U4456 (N_4456,In_1321,In_160);
and U4457 (N_4457,In_1163,In_1536);
nor U4458 (N_4458,In_2902,In_2430);
and U4459 (N_4459,In_213,In_809);
or U4460 (N_4460,In_557,In_2712);
and U4461 (N_4461,In_1189,In_1689);
nor U4462 (N_4462,In_762,In_1371);
and U4463 (N_4463,In_2410,In_1386);
nor U4464 (N_4464,In_925,In_850);
or U4465 (N_4465,In_30,In_1899);
nand U4466 (N_4466,In_2891,In_19);
nor U4467 (N_4467,In_554,In_1578);
nor U4468 (N_4468,In_421,In_1937);
and U4469 (N_4469,In_2867,In_1294);
nor U4470 (N_4470,In_1040,In_254);
or U4471 (N_4471,In_231,In_2883);
and U4472 (N_4472,In_432,In_1995);
and U4473 (N_4473,In_1506,In_1770);
or U4474 (N_4474,In_354,In_2656);
nand U4475 (N_4475,In_338,In_351);
or U4476 (N_4476,In_2248,In_2350);
and U4477 (N_4477,In_2032,In_1133);
nor U4478 (N_4478,In_2441,In_2021);
or U4479 (N_4479,In_2893,In_727);
and U4480 (N_4480,In_1122,In_1624);
nor U4481 (N_4481,In_778,In_427);
or U4482 (N_4482,In_484,In_2066);
xnor U4483 (N_4483,In_2741,In_742);
nor U4484 (N_4484,In_1438,In_1703);
or U4485 (N_4485,In_1742,In_415);
nor U4486 (N_4486,In_62,In_593);
nor U4487 (N_4487,In_1762,In_2642);
nand U4488 (N_4488,In_1857,In_2995);
or U4489 (N_4489,In_2344,In_2376);
nand U4490 (N_4490,In_2526,In_1759);
nor U4491 (N_4491,In_525,In_2786);
nor U4492 (N_4492,In_1031,In_568);
or U4493 (N_4493,In_1989,In_2732);
and U4494 (N_4494,In_1380,In_1237);
nand U4495 (N_4495,In_661,In_2059);
nor U4496 (N_4496,In_1742,In_2434);
nand U4497 (N_4497,In_1946,In_1903);
and U4498 (N_4498,In_1489,In_2841);
and U4499 (N_4499,In_332,In_731);
nand U4500 (N_4500,In_2682,In_2254);
nand U4501 (N_4501,In_2827,In_2547);
nor U4502 (N_4502,In_2392,In_2357);
nor U4503 (N_4503,In_1184,In_1609);
nand U4504 (N_4504,In_2744,In_2413);
nor U4505 (N_4505,In_563,In_2949);
nor U4506 (N_4506,In_2784,In_2598);
nand U4507 (N_4507,In_227,In_2658);
nand U4508 (N_4508,In_1743,In_2617);
xor U4509 (N_4509,In_2046,In_2685);
and U4510 (N_4510,In_1561,In_1176);
nor U4511 (N_4511,In_948,In_1489);
nor U4512 (N_4512,In_113,In_15);
nor U4513 (N_4513,In_639,In_1517);
nand U4514 (N_4514,In_1191,In_1427);
or U4515 (N_4515,In_1359,In_1065);
nand U4516 (N_4516,In_1767,In_224);
xnor U4517 (N_4517,In_1808,In_943);
and U4518 (N_4518,In_2272,In_42);
nand U4519 (N_4519,In_142,In_586);
and U4520 (N_4520,In_2003,In_392);
nor U4521 (N_4521,In_2093,In_2471);
nand U4522 (N_4522,In_1008,In_697);
nor U4523 (N_4523,In_2160,In_1395);
nor U4524 (N_4524,In_1315,In_242);
nor U4525 (N_4525,In_2092,In_289);
and U4526 (N_4526,In_1877,In_964);
nor U4527 (N_4527,In_2500,In_1748);
nand U4528 (N_4528,In_162,In_2988);
and U4529 (N_4529,In_394,In_1098);
or U4530 (N_4530,In_2375,In_714);
or U4531 (N_4531,In_2905,In_925);
xnor U4532 (N_4532,In_1245,In_1793);
nor U4533 (N_4533,In_574,In_2146);
nor U4534 (N_4534,In_887,In_1080);
nand U4535 (N_4535,In_23,In_1182);
and U4536 (N_4536,In_1038,In_1400);
or U4537 (N_4537,In_2781,In_1051);
or U4538 (N_4538,In_2351,In_2025);
or U4539 (N_4539,In_1089,In_2417);
or U4540 (N_4540,In_2921,In_1818);
or U4541 (N_4541,In_1670,In_2215);
xnor U4542 (N_4542,In_1732,In_869);
nand U4543 (N_4543,In_538,In_714);
and U4544 (N_4544,In_174,In_1660);
nor U4545 (N_4545,In_727,In_2402);
or U4546 (N_4546,In_1684,In_1313);
and U4547 (N_4547,In_1021,In_1513);
nor U4548 (N_4548,In_2957,In_1337);
and U4549 (N_4549,In_487,In_175);
xor U4550 (N_4550,In_576,In_1767);
or U4551 (N_4551,In_2644,In_282);
or U4552 (N_4552,In_2644,In_2422);
nor U4553 (N_4553,In_1939,In_2083);
and U4554 (N_4554,In_798,In_1611);
xnor U4555 (N_4555,In_1462,In_1714);
or U4556 (N_4556,In_2001,In_2916);
nand U4557 (N_4557,In_884,In_2999);
nor U4558 (N_4558,In_2413,In_2007);
xor U4559 (N_4559,In_1855,In_875);
nand U4560 (N_4560,In_2490,In_515);
nor U4561 (N_4561,In_1240,In_941);
nand U4562 (N_4562,In_2648,In_2438);
xnor U4563 (N_4563,In_2484,In_817);
or U4564 (N_4564,In_2238,In_998);
and U4565 (N_4565,In_2690,In_352);
or U4566 (N_4566,In_1105,In_1101);
or U4567 (N_4567,In_772,In_2148);
and U4568 (N_4568,In_2605,In_2751);
xnor U4569 (N_4569,In_1082,In_564);
or U4570 (N_4570,In_1464,In_248);
nor U4571 (N_4571,In_624,In_2315);
and U4572 (N_4572,In_1807,In_89);
and U4573 (N_4573,In_2622,In_752);
nand U4574 (N_4574,In_1339,In_793);
xor U4575 (N_4575,In_1344,In_1536);
or U4576 (N_4576,In_1651,In_872);
xor U4577 (N_4577,In_585,In_2897);
xnor U4578 (N_4578,In_2865,In_153);
xnor U4579 (N_4579,In_1690,In_2532);
or U4580 (N_4580,In_135,In_2564);
nand U4581 (N_4581,In_1120,In_684);
or U4582 (N_4582,In_2117,In_571);
xnor U4583 (N_4583,In_919,In_2601);
nand U4584 (N_4584,In_1405,In_2197);
and U4585 (N_4585,In_2371,In_1794);
nand U4586 (N_4586,In_2836,In_1179);
xnor U4587 (N_4587,In_131,In_562);
or U4588 (N_4588,In_396,In_847);
and U4589 (N_4589,In_1528,In_619);
or U4590 (N_4590,In_317,In_724);
or U4591 (N_4591,In_678,In_329);
nand U4592 (N_4592,In_1453,In_1993);
or U4593 (N_4593,In_357,In_1314);
nor U4594 (N_4594,In_1680,In_2451);
nor U4595 (N_4595,In_1159,In_1171);
or U4596 (N_4596,In_808,In_1991);
and U4597 (N_4597,In_2637,In_1359);
and U4598 (N_4598,In_485,In_2713);
nand U4599 (N_4599,In_1953,In_1827);
nor U4600 (N_4600,In_1194,In_1388);
nor U4601 (N_4601,In_1804,In_2701);
xor U4602 (N_4602,In_1032,In_2120);
nand U4603 (N_4603,In_2918,In_301);
nand U4604 (N_4604,In_184,In_1115);
nand U4605 (N_4605,In_691,In_169);
nand U4606 (N_4606,In_929,In_232);
and U4607 (N_4607,In_394,In_1969);
and U4608 (N_4608,In_560,In_1213);
nand U4609 (N_4609,In_505,In_992);
or U4610 (N_4610,In_1938,In_2503);
nand U4611 (N_4611,In_1996,In_1144);
and U4612 (N_4612,In_847,In_2254);
or U4613 (N_4613,In_2648,In_1494);
nor U4614 (N_4614,In_2636,In_1463);
nand U4615 (N_4615,In_1385,In_2806);
nand U4616 (N_4616,In_290,In_999);
nand U4617 (N_4617,In_2312,In_1820);
nor U4618 (N_4618,In_1320,In_2019);
nor U4619 (N_4619,In_1465,In_1005);
or U4620 (N_4620,In_949,In_1252);
nor U4621 (N_4621,In_2277,In_741);
and U4622 (N_4622,In_806,In_2569);
nor U4623 (N_4623,In_1081,In_2606);
nand U4624 (N_4624,In_423,In_276);
or U4625 (N_4625,In_2122,In_1155);
nand U4626 (N_4626,In_1408,In_2593);
xor U4627 (N_4627,In_1767,In_1127);
and U4628 (N_4628,In_2088,In_481);
or U4629 (N_4629,In_2167,In_387);
nand U4630 (N_4630,In_407,In_1786);
or U4631 (N_4631,In_1562,In_2208);
nand U4632 (N_4632,In_2394,In_633);
and U4633 (N_4633,In_201,In_2565);
or U4634 (N_4634,In_2191,In_2228);
nand U4635 (N_4635,In_396,In_781);
and U4636 (N_4636,In_87,In_1483);
xnor U4637 (N_4637,In_85,In_1365);
and U4638 (N_4638,In_2254,In_1689);
nor U4639 (N_4639,In_2234,In_1660);
and U4640 (N_4640,In_2953,In_2103);
nor U4641 (N_4641,In_929,In_2938);
nand U4642 (N_4642,In_1576,In_855);
nand U4643 (N_4643,In_922,In_2606);
nand U4644 (N_4644,In_2278,In_2525);
xnor U4645 (N_4645,In_1896,In_1360);
xor U4646 (N_4646,In_2777,In_146);
xnor U4647 (N_4647,In_2297,In_1726);
nor U4648 (N_4648,In_298,In_606);
nand U4649 (N_4649,In_2995,In_326);
or U4650 (N_4650,In_1733,In_2596);
nand U4651 (N_4651,In_668,In_2822);
nor U4652 (N_4652,In_789,In_1723);
nand U4653 (N_4653,In_2923,In_1838);
nand U4654 (N_4654,In_1592,In_2624);
nor U4655 (N_4655,In_529,In_1292);
or U4656 (N_4656,In_1833,In_2384);
nor U4657 (N_4657,In_2950,In_1453);
nand U4658 (N_4658,In_1231,In_1876);
and U4659 (N_4659,In_1034,In_1448);
nand U4660 (N_4660,In_1843,In_1671);
xor U4661 (N_4661,In_594,In_2768);
and U4662 (N_4662,In_1799,In_2584);
and U4663 (N_4663,In_2374,In_2444);
nor U4664 (N_4664,In_508,In_183);
nand U4665 (N_4665,In_1573,In_346);
nand U4666 (N_4666,In_373,In_996);
or U4667 (N_4667,In_455,In_829);
and U4668 (N_4668,In_1813,In_1284);
and U4669 (N_4669,In_2669,In_1889);
or U4670 (N_4670,In_2701,In_1186);
or U4671 (N_4671,In_2497,In_2294);
xnor U4672 (N_4672,In_769,In_1311);
nand U4673 (N_4673,In_2311,In_1199);
nor U4674 (N_4674,In_1626,In_290);
nand U4675 (N_4675,In_1180,In_2849);
xnor U4676 (N_4676,In_2122,In_4);
or U4677 (N_4677,In_421,In_1314);
nand U4678 (N_4678,In_1981,In_1379);
and U4679 (N_4679,In_1168,In_1191);
nand U4680 (N_4680,In_2935,In_1430);
nand U4681 (N_4681,In_1370,In_2467);
or U4682 (N_4682,In_1742,In_1137);
or U4683 (N_4683,In_2207,In_2018);
and U4684 (N_4684,In_2644,In_746);
nor U4685 (N_4685,In_1581,In_1186);
xnor U4686 (N_4686,In_1231,In_1164);
or U4687 (N_4687,In_233,In_911);
nor U4688 (N_4688,In_2438,In_1948);
nor U4689 (N_4689,In_2106,In_2052);
nor U4690 (N_4690,In_1099,In_773);
and U4691 (N_4691,In_1370,In_1329);
nand U4692 (N_4692,In_1878,In_246);
or U4693 (N_4693,In_544,In_2951);
nor U4694 (N_4694,In_726,In_77);
nor U4695 (N_4695,In_46,In_2992);
nor U4696 (N_4696,In_1590,In_421);
and U4697 (N_4697,In_570,In_2591);
nand U4698 (N_4698,In_1983,In_2972);
nor U4699 (N_4699,In_1314,In_71);
and U4700 (N_4700,In_1418,In_423);
or U4701 (N_4701,In_2634,In_409);
or U4702 (N_4702,In_2531,In_1304);
nor U4703 (N_4703,In_623,In_1989);
nand U4704 (N_4704,In_1940,In_1223);
or U4705 (N_4705,In_2353,In_1404);
and U4706 (N_4706,In_2797,In_1539);
xnor U4707 (N_4707,In_1635,In_1774);
nor U4708 (N_4708,In_627,In_2860);
or U4709 (N_4709,In_557,In_674);
xnor U4710 (N_4710,In_1464,In_1201);
or U4711 (N_4711,In_437,In_2185);
xnor U4712 (N_4712,In_763,In_2734);
nand U4713 (N_4713,In_1132,In_158);
nor U4714 (N_4714,In_1354,In_2247);
nand U4715 (N_4715,In_496,In_980);
nor U4716 (N_4716,In_2210,In_921);
nor U4717 (N_4717,In_115,In_16);
and U4718 (N_4718,In_292,In_206);
nand U4719 (N_4719,In_6,In_1830);
xor U4720 (N_4720,In_1983,In_2133);
nand U4721 (N_4721,In_81,In_181);
or U4722 (N_4722,In_614,In_547);
nand U4723 (N_4723,In_2219,In_1947);
nor U4724 (N_4724,In_2081,In_1293);
or U4725 (N_4725,In_169,In_1304);
and U4726 (N_4726,In_2610,In_1993);
nand U4727 (N_4727,In_894,In_2864);
nand U4728 (N_4728,In_235,In_1014);
and U4729 (N_4729,In_2154,In_1551);
nor U4730 (N_4730,In_34,In_673);
nor U4731 (N_4731,In_2707,In_2790);
or U4732 (N_4732,In_929,In_2469);
or U4733 (N_4733,In_409,In_427);
and U4734 (N_4734,In_2104,In_2472);
nand U4735 (N_4735,In_2428,In_2702);
nand U4736 (N_4736,In_1581,In_2790);
nor U4737 (N_4737,In_321,In_2694);
nand U4738 (N_4738,In_2045,In_1216);
or U4739 (N_4739,In_2739,In_396);
nor U4740 (N_4740,In_1806,In_1025);
nor U4741 (N_4741,In_1876,In_2851);
nor U4742 (N_4742,In_1861,In_12);
and U4743 (N_4743,In_861,In_444);
nand U4744 (N_4744,In_791,In_2974);
or U4745 (N_4745,In_2600,In_1853);
and U4746 (N_4746,In_1084,In_2469);
nor U4747 (N_4747,In_2574,In_2982);
nor U4748 (N_4748,In_1735,In_473);
nand U4749 (N_4749,In_965,In_2655);
nand U4750 (N_4750,In_209,In_675);
and U4751 (N_4751,In_1094,In_49);
xnor U4752 (N_4752,In_794,In_2772);
nand U4753 (N_4753,In_622,In_1363);
and U4754 (N_4754,In_1461,In_1366);
nand U4755 (N_4755,In_2760,In_2989);
nor U4756 (N_4756,In_2383,In_21);
nand U4757 (N_4757,In_828,In_1246);
nand U4758 (N_4758,In_681,In_1908);
or U4759 (N_4759,In_640,In_19);
nand U4760 (N_4760,In_1242,In_1082);
or U4761 (N_4761,In_2123,In_2391);
or U4762 (N_4762,In_1803,In_849);
nand U4763 (N_4763,In_2667,In_1686);
nand U4764 (N_4764,In_1383,In_1762);
nor U4765 (N_4765,In_1683,In_89);
and U4766 (N_4766,In_10,In_1295);
nand U4767 (N_4767,In_1947,In_2604);
nand U4768 (N_4768,In_895,In_1215);
or U4769 (N_4769,In_202,In_800);
nand U4770 (N_4770,In_157,In_2928);
or U4771 (N_4771,In_1944,In_117);
nor U4772 (N_4772,In_2299,In_2993);
or U4773 (N_4773,In_1920,In_2180);
and U4774 (N_4774,In_634,In_2236);
nor U4775 (N_4775,In_2430,In_2087);
nor U4776 (N_4776,In_462,In_2304);
and U4777 (N_4777,In_2570,In_2090);
xnor U4778 (N_4778,In_1942,In_2980);
nand U4779 (N_4779,In_1450,In_2325);
nor U4780 (N_4780,In_2796,In_2351);
or U4781 (N_4781,In_1056,In_1431);
nand U4782 (N_4782,In_1824,In_2103);
nor U4783 (N_4783,In_1184,In_686);
or U4784 (N_4784,In_2768,In_2267);
and U4785 (N_4785,In_1628,In_1136);
and U4786 (N_4786,In_2385,In_440);
and U4787 (N_4787,In_207,In_2159);
nor U4788 (N_4788,In_182,In_256);
nand U4789 (N_4789,In_1014,In_2804);
nor U4790 (N_4790,In_329,In_323);
or U4791 (N_4791,In_1763,In_932);
xor U4792 (N_4792,In_812,In_2695);
or U4793 (N_4793,In_2615,In_2390);
xor U4794 (N_4794,In_41,In_986);
nand U4795 (N_4795,In_1175,In_2551);
or U4796 (N_4796,In_534,In_2031);
or U4797 (N_4797,In_1945,In_136);
or U4798 (N_4798,In_2494,In_188);
or U4799 (N_4799,In_951,In_2041);
nand U4800 (N_4800,In_2867,In_2818);
and U4801 (N_4801,In_426,In_2627);
or U4802 (N_4802,In_621,In_728);
nor U4803 (N_4803,In_1259,In_765);
nor U4804 (N_4804,In_1285,In_2916);
nand U4805 (N_4805,In_1017,In_2659);
nand U4806 (N_4806,In_1898,In_2356);
and U4807 (N_4807,In_362,In_308);
nor U4808 (N_4808,In_1329,In_1747);
or U4809 (N_4809,In_903,In_2202);
nor U4810 (N_4810,In_218,In_1457);
and U4811 (N_4811,In_1506,In_2454);
and U4812 (N_4812,In_116,In_323);
and U4813 (N_4813,In_1697,In_2981);
or U4814 (N_4814,In_777,In_1792);
nor U4815 (N_4815,In_2179,In_2375);
nor U4816 (N_4816,In_990,In_1291);
nor U4817 (N_4817,In_513,In_1723);
xor U4818 (N_4818,In_1243,In_1753);
nand U4819 (N_4819,In_863,In_609);
and U4820 (N_4820,In_1110,In_1052);
nand U4821 (N_4821,In_1831,In_1932);
nand U4822 (N_4822,In_1696,In_552);
and U4823 (N_4823,In_2276,In_2015);
nand U4824 (N_4824,In_2620,In_2183);
and U4825 (N_4825,In_739,In_1499);
and U4826 (N_4826,In_1038,In_707);
and U4827 (N_4827,In_542,In_745);
nor U4828 (N_4828,In_2332,In_1705);
nor U4829 (N_4829,In_2205,In_1092);
nand U4830 (N_4830,In_1157,In_180);
nor U4831 (N_4831,In_1410,In_1779);
nor U4832 (N_4832,In_1389,In_2819);
and U4833 (N_4833,In_471,In_2598);
nand U4834 (N_4834,In_890,In_560);
nand U4835 (N_4835,In_914,In_2179);
or U4836 (N_4836,In_2145,In_2667);
and U4837 (N_4837,In_2452,In_1888);
nor U4838 (N_4838,In_1969,In_1644);
nand U4839 (N_4839,In_633,In_1545);
nand U4840 (N_4840,In_242,In_2196);
nor U4841 (N_4841,In_736,In_562);
or U4842 (N_4842,In_858,In_2700);
or U4843 (N_4843,In_2877,In_1836);
xor U4844 (N_4844,In_2486,In_1313);
nor U4845 (N_4845,In_246,In_878);
or U4846 (N_4846,In_2665,In_2490);
and U4847 (N_4847,In_2146,In_2155);
or U4848 (N_4848,In_472,In_1644);
nor U4849 (N_4849,In_2041,In_896);
or U4850 (N_4850,In_1008,In_2431);
or U4851 (N_4851,In_2700,In_2912);
nand U4852 (N_4852,In_104,In_1533);
and U4853 (N_4853,In_2252,In_2374);
nand U4854 (N_4854,In_2281,In_618);
nand U4855 (N_4855,In_1317,In_2923);
or U4856 (N_4856,In_90,In_208);
and U4857 (N_4857,In_2496,In_900);
and U4858 (N_4858,In_2039,In_1737);
nand U4859 (N_4859,In_576,In_372);
or U4860 (N_4860,In_1976,In_1413);
nand U4861 (N_4861,In_239,In_184);
and U4862 (N_4862,In_1031,In_2662);
xnor U4863 (N_4863,In_671,In_2690);
xnor U4864 (N_4864,In_2080,In_717);
nand U4865 (N_4865,In_1566,In_2361);
and U4866 (N_4866,In_455,In_1527);
and U4867 (N_4867,In_1966,In_1696);
nor U4868 (N_4868,In_251,In_73);
nor U4869 (N_4869,In_1314,In_444);
xnor U4870 (N_4870,In_208,In_481);
and U4871 (N_4871,In_696,In_1268);
nand U4872 (N_4872,In_565,In_2643);
and U4873 (N_4873,In_1625,In_2517);
and U4874 (N_4874,In_29,In_2999);
and U4875 (N_4875,In_366,In_1035);
and U4876 (N_4876,In_601,In_2173);
and U4877 (N_4877,In_2610,In_2635);
nand U4878 (N_4878,In_492,In_2847);
nand U4879 (N_4879,In_1806,In_1068);
nand U4880 (N_4880,In_2689,In_886);
or U4881 (N_4881,In_1917,In_2405);
nand U4882 (N_4882,In_1053,In_2609);
nor U4883 (N_4883,In_2355,In_2503);
nand U4884 (N_4884,In_80,In_2879);
or U4885 (N_4885,In_1510,In_2132);
nand U4886 (N_4886,In_87,In_2368);
and U4887 (N_4887,In_2357,In_98);
xor U4888 (N_4888,In_1973,In_308);
or U4889 (N_4889,In_31,In_859);
or U4890 (N_4890,In_1029,In_1305);
and U4891 (N_4891,In_471,In_1677);
nor U4892 (N_4892,In_1316,In_505);
and U4893 (N_4893,In_2222,In_384);
or U4894 (N_4894,In_231,In_51);
nand U4895 (N_4895,In_438,In_1680);
nand U4896 (N_4896,In_759,In_2034);
and U4897 (N_4897,In_519,In_1567);
or U4898 (N_4898,In_379,In_2664);
and U4899 (N_4899,In_2815,In_1575);
nor U4900 (N_4900,In_1244,In_1558);
and U4901 (N_4901,In_2845,In_893);
xnor U4902 (N_4902,In_64,In_589);
nand U4903 (N_4903,In_2172,In_1270);
and U4904 (N_4904,In_948,In_2423);
or U4905 (N_4905,In_2391,In_1061);
nand U4906 (N_4906,In_1805,In_505);
nand U4907 (N_4907,In_830,In_1317);
or U4908 (N_4908,In_445,In_813);
nand U4909 (N_4909,In_224,In_1702);
or U4910 (N_4910,In_491,In_987);
or U4911 (N_4911,In_781,In_362);
xor U4912 (N_4912,In_2789,In_1665);
and U4913 (N_4913,In_1001,In_1408);
xor U4914 (N_4914,In_1265,In_61);
and U4915 (N_4915,In_301,In_1774);
or U4916 (N_4916,In_1468,In_2864);
nand U4917 (N_4917,In_27,In_1350);
or U4918 (N_4918,In_978,In_1155);
or U4919 (N_4919,In_2001,In_1126);
and U4920 (N_4920,In_2330,In_1274);
nor U4921 (N_4921,In_1595,In_2647);
or U4922 (N_4922,In_2385,In_401);
nand U4923 (N_4923,In_953,In_340);
nor U4924 (N_4924,In_2726,In_627);
and U4925 (N_4925,In_227,In_747);
nor U4926 (N_4926,In_903,In_1608);
nand U4927 (N_4927,In_1395,In_2078);
or U4928 (N_4928,In_1553,In_2950);
or U4929 (N_4929,In_879,In_1040);
nand U4930 (N_4930,In_2688,In_2332);
or U4931 (N_4931,In_2852,In_1567);
nor U4932 (N_4932,In_48,In_2404);
nor U4933 (N_4933,In_389,In_831);
or U4934 (N_4934,In_499,In_677);
and U4935 (N_4935,In_743,In_2372);
nor U4936 (N_4936,In_344,In_1791);
or U4937 (N_4937,In_1309,In_941);
nand U4938 (N_4938,In_2014,In_821);
or U4939 (N_4939,In_1734,In_2564);
nand U4940 (N_4940,In_1642,In_1709);
or U4941 (N_4941,In_95,In_2521);
nand U4942 (N_4942,In_1397,In_2842);
or U4943 (N_4943,In_2447,In_1334);
or U4944 (N_4944,In_395,In_2735);
and U4945 (N_4945,In_565,In_618);
or U4946 (N_4946,In_616,In_65);
and U4947 (N_4947,In_1037,In_757);
nor U4948 (N_4948,In_1982,In_1243);
xor U4949 (N_4949,In_1133,In_1867);
nor U4950 (N_4950,In_510,In_902);
nand U4951 (N_4951,In_2082,In_1669);
and U4952 (N_4952,In_1703,In_2507);
or U4953 (N_4953,In_1333,In_2469);
nor U4954 (N_4954,In_316,In_2554);
and U4955 (N_4955,In_2555,In_2859);
and U4956 (N_4956,In_116,In_1358);
or U4957 (N_4957,In_283,In_1702);
or U4958 (N_4958,In_1328,In_135);
nand U4959 (N_4959,In_434,In_2816);
nor U4960 (N_4960,In_1390,In_2297);
nor U4961 (N_4961,In_29,In_2935);
and U4962 (N_4962,In_350,In_109);
nand U4963 (N_4963,In_2510,In_1164);
and U4964 (N_4964,In_2064,In_1219);
nand U4965 (N_4965,In_2179,In_2260);
and U4966 (N_4966,In_2990,In_1389);
or U4967 (N_4967,In_464,In_1618);
nand U4968 (N_4968,In_147,In_1324);
and U4969 (N_4969,In_2055,In_2819);
and U4970 (N_4970,In_2739,In_2789);
nand U4971 (N_4971,In_1918,In_1542);
nor U4972 (N_4972,In_2475,In_2241);
nand U4973 (N_4973,In_1084,In_42);
or U4974 (N_4974,In_2649,In_1416);
nor U4975 (N_4975,In_2999,In_2770);
nand U4976 (N_4976,In_1806,In_2481);
nor U4977 (N_4977,In_798,In_963);
nor U4978 (N_4978,In_1516,In_1469);
or U4979 (N_4979,In_1020,In_2766);
or U4980 (N_4980,In_1870,In_1144);
and U4981 (N_4981,In_2300,In_1447);
or U4982 (N_4982,In_1831,In_1891);
and U4983 (N_4983,In_733,In_1083);
and U4984 (N_4984,In_526,In_151);
nor U4985 (N_4985,In_1651,In_2820);
and U4986 (N_4986,In_2053,In_2876);
nand U4987 (N_4987,In_2508,In_2200);
nor U4988 (N_4988,In_1845,In_2809);
or U4989 (N_4989,In_2476,In_17);
xnor U4990 (N_4990,In_1230,In_242);
or U4991 (N_4991,In_1540,In_2636);
nor U4992 (N_4992,In_2241,In_1335);
nor U4993 (N_4993,In_14,In_1626);
and U4994 (N_4994,In_1619,In_1019);
nor U4995 (N_4995,In_1208,In_188);
and U4996 (N_4996,In_926,In_2562);
xnor U4997 (N_4997,In_2995,In_2933);
nor U4998 (N_4998,In_495,In_1913);
or U4999 (N_4999,In_1366,In_2190);
nor U5000 (N_5000,In_546,In_61);
nor U5001 (N_5001,In_331,In_140);
nand U5002 (N_5002,In_945,In_2033);
nand U5003 (N_5003,In_383,In_2056);
and U5004 (N_5004,In_784,In_1452);
nand U5005 (N_5005,In_1295,In_55);
xor U5006 (N_5006,In_1445,In_1358);
nand U5007 (N_5007,In_27,In_328);
xor U5008 (N_5008,In_392,In_2175);
nand U5009 (N_5009,In_2257,In_2077);
or U5010 (N_5010,In_2168,In_1274);
nor U5011 (N_5011,In_1626,In_1183);
or U5012 (N_5012,In_1114,In_1840);
nor U5013 (N_5013,In_2714,In_692);
nor U5014 (N_5014,In_1208,In_1228);
xor U5015 (N_5015,In_837,In_1114);
xnor U5016 (N_5016,In_2915,In_1712);
xor U5017 (N_5017,In_2558,In_2624);
nor U5018 (N_5018,In_90,In_706);
and U5019 (N_5019,In_792,In_991);
nor U5020 (N_5020,In_2617,In_192);
nand U5021 (N_5021,In_2895,In_2427);
xnor U5022 (N_5022,In_2406,In_1581);
and U5023 (N_5023,In_142,In_2594);
nor U5024 (N_5024,In_1557,In_697);
nor U5025 (N_5025,In_981,In_1056);
nor U5026 (N_5026,In_144,In_149);
nand U5027 (N_5027,In_2125,In_2570);
or U5028 (N_5028,In_2725,In_2180);
xnor U5029 (N_5029,In_1292,In_2597);
and U5030 (N_5030,In_2047,In_2187);
nand U5031 (N_5031,In_1320,In_1926);
nand U5032 (N_5032,In_686,In_842);
or U5033 (N_5033,In_595,In_2274);
and U5034 (N_5034,In_1178,In_2788);
or U5035 (N_5035,In_2936,In_1674);
and U5036 (N_5036,In_1020,In_754);
nor U5037 (N_5037,In_929,In_2371);
or U5038 (N_5038,In_2408,In_307);
or U5039 (N_5039,In_1976,In_323);
and U5040 (N_5040,In_1501,In_1010);
and U5041 (N_5041,In_1677,In_1071);
and U5042 (N_5042,In_1430,In_599);
and U5043 (N_5043,In_2654,In_555);
or U5044 (N_5044,In_1180,In_1131);
nand U5045 (N_5045,In_320,In_1541);
xor U5046 (N_5046,In_194,In_1288);
nand U5047 (N_5047,In_118,In_1625);
and U5048 (N_5048,In_588,In_561);
nor U5049 (N_5049,In_945,In_1224);
xnor U5050 (N_5050,In_1403,In_1537);
nor U5051 (N_5051,In_106,In_387);
and U5052 (N_5052,In_2360,In_906);
nand U5053 (N_5053,In_134,In_2720);
nor U5054 (N_5054,In_552,In_2916);
nor U5055 (N_5055,In_2583,In_2907);
and U5056 (N_5056,In_2042,In_2134);
and U5057 (N_5057,In_137,In_2839);
nand U5058 (N_5058,In_1930,In_2541);
nand U5059 (N_5059,In_2935,In_1321);
nand U5060 (N_5060,In_2325,In_1353);
nand U5061 (N_5061,In_1479,In_2570);
and U5062 (N_5062,In_1129,In_2568);
nand U5063 (N_5063,In_2483,In_2590);
and U5064 (N_5064,In_1226,In_1356);
nor U5065 (N_5065,In_2435,In_2511);
nand U5066 (N_5066,In_362,In_57);
nand U5067 (N_5067,In_1067,In_1474);
and U5068 (N_5068,In_2852,In_2226);
or U5069 (N_5069,In_2742,In_853);
xor U5070 (N_5070,In_1022,In_1456);
xor U5071 (N_5071,In_2409,In_1546);
nor U5072 (N_5072,In_2020,In_2654);
nor U5073 (N_5073,In_599,In_1022);
xor U5074 (N_5074,In_2567,In_748);
or U5075 (N_5075,In_1898,In_31);
nor U5076 (N_5076,In_168,In_2791);
or U5077 (N_5077,In_140,In_2560);
nor U5078 (N_5078,In_801,In_1750);
nand U5079 (N_5079,In_2251,In_2980);
and U5080 (N_5080,In_679,In_1628);
and U5081 (N_5081,In_90,In_420);
and U5082 (N_5082,In_1187,In_1193);
nor U5083 (N_5083,In_2292,In_744);
and U5084 (N_5084,In_1144,In_1102);
nand U5085 (N_5085,In_1945,In_1258);
nor U5086 (N_5086,In_359,In_1132);
nor U5087 (N_5087,In_2287,In_78);
nor U5088 (N_5088,In_1216,In_814);
and U5089 (N_5089,In_2586,In_420);
nand U5090 (N_5090,In_1665,In_1400);
nand U5091 (N_5091,In_2770,In_308);
xor U5092 (N_5092,In_2194,In_853);
nand U5093 (N_5093,In_1200,In_505);
nand U5094 (N_5094,In_1517,In_2997);
and U5095 (N_5095,In_1147,In_1405);
nand U5096 (N_5096,In_621,In_1814);
or U5097 (N_5097,In_2990,In_985);
nand U5098 (N_5098,In_820,In_660);
nor U5099 (N_5099,In_2744,In_2245);
or U5100 (N_5100,In_2096,In_1627);
or U5101 (N_5101,In_344,In_1792);
and U5102 (N_5102,In_1247,In_2314);
xor U5103 (N_5103,In_190,In_956);
or U5104 (N_5104,In_1730,In_2292);
nor U5105 (N_5105,In_596,In_1051);
nor U5106 (N_5106,In_1140,In_385);
nand U5107 (N_5107,In_1010,In_2723);
and U5108 (N_5108,In_2438,In_372);
xnor U5109 (N_5109,In_980,In_1664);
nor U5110 (N_5110,In_1425,In_385);
nand U5111 (N_5111,In_2227,In_2851);
nor U5112 (N_5112,In_1830,In_473);
and U5113 (N_5113,In_2988,In_1290);
nand U5114 (N_5114,In_1028,In_445);
nand U5115 (N_5115,In_217,In_2606);
and U5116 (N_5116,In_606,In_2976);
nor U5117 (N_5117,In_1523,In_1211);
and U5118 (N_5118,In_1720,In_636);
nand U5119 (N_5119,In_480,In_1522);
or U5120 (N_5120,In_459,In_1902);
nor U5121 (N_5121,In_419,In_134);
nor U5122 (N_5122,In_1014,In_1178);
xnor U5123 (N_5123,In_140,In_248);
and U5124 (N_5124,In_1496,In_2281);
nand U5125 (N_5125,In_2508,In_1729);
and U5126 (N_5126,In_686,In_2564);
nand U5127 (N_5127,In_27,In_2260);
nor U5128 (N_5128,In_1890,In_908);
nor U5129 (N_5129,In_2818,In_997);
nand U5130 (N_5130,In_364,In_561);
xor U5131 (N_5131,In_2585,In_674);
nor U5132 (N_5132,In_2192,In_1790);
or U5133 (N_5133,In_2268,In_2344);
and U5134 (N_5134,In_216,In_1243);
and U5135 (N_5135,In_1980,In_2385);
xnor U5136 (N_5136,In_2232,In_1372);
nor U5137 (N_5137,In_389,In_2046);
nand U5138 (N_5138,In_1212,In_443);
or U5139 (N_5139,In_2679,In_2653);
or U5140 (N_5140,In_590,In_677);
or U5141 (N_5141,In_195,In_2734);
nand U5142 (N_5142,In_395,In_1759);
or U5143 (N_5143,In_1883,In_2665);
nor U5144 (N_5144,In_27,In_2441);
xor U5145 (N_5145,In_2910,In_1319);
or U5146 (N_5146,In_2835,In_2380);
and U5147 (N_5147,In_2553,In_598);
nand U5148 (N_5148,In_1284,In_2673);
nor U5149 (N_5149,In_2877,In_2404);
or U5150 (N_5150,In_2615,In_1749);
and U5151 (N_5151,In_2825,In_2288);
nand U5152 (N_5152,In_393,In_1973);
and U5153 (N_5153,In_1397,In_621);
nor U5154 (N_5154,In_2927,In_901);
and U5155 (N_5155,In_2720,In_1334);
and U5156 (N_5156,In_866,In_1365);
nand U5157 (N_5157,In_1007,In_2188);
nand U5158 (N_5158,In_2567,In_2221);
or U5159 (N_5159,In_1278,In_2468);
or U5160 (N_5160,In_1510,In_51);
and U5161 (N_5161,In_103,In_1369);
and U5162 (N_5162,In_857,In_869);
xnor U5163 (N_5163,In_1405,In_1359);
nand U5164 (N_5164,In_1449,In_1750);
and U5165 (N_5165,In_2806,In_729);
nand U5166 (N_5166,In_2112,In_899);
nand U5167 (N_5167,In_723,In_858);
xor U5168 (N_5168,In_910,In_397);
or U5169 (N_5169,In_1687,In_1849);
nand U5170 (N_5170,In_1782,In_965);
xnor U5171 (N_5171,In_98,In_1335);
and U5172 (N_5172,In_1452,In_983);
nor U5173 (N_5173,In_409,In_313);
nand U5174 (N_5174,In_2645,In_1754);
nand U5175 (N_5175,In_195,In_2717);
nor U5176 (N_5176,In_2633,In_2785);
or U5177 (N_5177,In_2960,In_505);
or U5178 (N_5178,In_736,In_1824);
or U5179 (N_5179,In_2748,In_1397);
nor U5180 (N_5180,In_84,In_1205);
nand U5181 (N_5181,In_1079,In_751);
nand U5182 (N_5182,In_1159,In_1053);
or U5183 (N_5183,In_2538,In_1948);
or U5184 (N_5184,In_852,In_2398);
nor U5185 (N_5185,In_1518,In_442);
or U5186 (N_5186,In_859,In_2252);
or U5187 (N_5187,In_2040,In_577);
and U5188 (N_5188,In_2412,In_2290);
nand U5189 (N_5189,In_1727,In_1055);
xor U5190 (N_5190,In_1353,In_565);
or U5191 (N_5191,In_1459,In_1878);
nand U5192 (N_5192,In_2772,In_1087);
nor U5193 (N_5193,In_63,In_2834);
and U5194 (N_5194,In_121,In_315);
xnor U5195 (N_5195,In_685,In_1515);
nor U5196 (N_5196,In_1265,In_859);
or U5197 (N_5197,In_2816,In_2442);
and U5198 (N_5198,In_624,In_2501);
and U5199 (N_5199,In_1269,In_321);
or U5200 (N_5200,In_1885,In_2600);
or U5201 (N_5201,In_2255,In_312);
or U5202 (N_5202,In_123,In_1602);
xnor U5203 (N_5203,In_1899,In_2532);
nor U5204 (N_5204,In_2713,In_1543);
or U5205 (N_5205,In_1570,In_980);
and U5206 (N_5206,In_1916,In_2236);
nand U5207 (N_5207,In_1078,In_234);
or U5208 (N_5208,In_341,In_2975);
and U5209 (N_5209,In_1620,In_1018);
or U5210 (N_5210,In_2553,In_751);
nand U5211 (N_5211,In_2918,In_1593);
or U5212 (N_5212,In_2077,In_1245);
nand U5213 (N_5213,In_1080,In_671);
nor U5214 (N_5214,In_1644,In_2819);
nor U5215 (N_5215,In_2712,In_48);
nand U5216 (N_5216,In_2154,In_467);
nor U5217 (N_5217,In_730,In_22);
nand U5218 (N_5218,In_2185,In_1220);
or U5219 (N_5219,In_1892,In_928);
and U5220 (N_5220,In_1716,In_1355);
or U5221 (N_5221,In_872,In_2966);
or U5222 (N_5222,In_161,In_1646);
nor U5223 (N_5223,In_199,In_653);
and U5224 (N_5224,In_440,In_207);
or U5225 (N_5225,In_1325,In_120);
or U5226 (N_5226,In_975,In_2752);
nand U5227 (N_5227,In_1798,In_2342);
xnor U5228 (N_5228,In_1427,In_2265);
nand U5229 (N_5229,In_2190,In_2801);
nor U5230 (N_5230,In_214,In_139);
and U5231 (N_5231,In_1728,In_391);
and U5232 (N_5232,In_1852,In_134);
nor U5233 (N_5233,In_2983,In_2720);
nor U5234 (N_5234,In_1428,In_2953);
nand U5235 (N_5235,In_2769,In_1542);
and U5236 (N_5236,In_2404,In_2021);
xnor U5237 (N_5237,In_749,In_2027);
nor U5238 (N_5238,In_170,In_2199);
nor U5239 (N_5239,In_1819,In_2652);
nor U5240 (N_5240,In_799,In_2081);
nand U5241 (N_5241,In_2437,In_1857);
or U5242 (N_5242,In_1260,In_2325);
and U5243 (N_5243,In_1072,In_1430);
and U5244 (N_5244,In_117,In_822);
and U5245 (N_5245,In_1995,In_1794);
nand U5246 (N_5246,In_1672,In_1058);
nand U5247 (N_5247,In_2989,In_555);
and U5248 (N_5248,In_801,In_82);
nand U5249 (N_5249,In_441,In_1842);
and U5250 (N_5250,In_488,In_1950);
and U5251 (N_5251,In_2779,In_2321);
or U5252 (N_5252,In_733,In_2068);
nor U5253 (N_5253,In_1477,In_802);
nor U5254 (N_5254,In_467,In_1735);
xor U5255 (N_5255,In_2522,In_2621);
or U5256 (N_5256,In_159,In_2627);
or U5257 (N_5257,In_805,In_2328);
and U5258 (N_5258,In_1601,In_1140);
nand U5259 (N_5259,In_643,In_8);
or U5260 (N_5260,In_2116,In_1672);
nand U5261 (N_5261,In_1101,In_27);
nand U5262 (N_5262,In_1431,In_2468);
nor U5263 (N_5263,In_2680,In_2507);
nor U5264 (N_5264,In_1427,In_805);
and U5265 (N_5265,In_1804,In_2931);
nand U5266 (N_5266,In_1540,In_548);
nand U5267 (N_5267,In_2566,In_757);
nor U5268 (N_5268,In_1840,In_109);
nand U5269 (N_5269,In_2609,In_917);
nand U5270 (N_5270,In_2765,In_1603);
or U5271 (N_5271,In_1113,In_1957);
nand U5272 (N_5272,In_1994,In_1741);
nand U5273 (N_5273,In_1879,In_750);
or U5274 (N_5274,In_1630,In_854);
or U5275 (N_5275,In_100,In_250);
or U5276 (N_5276,In_2183,In_905);
and U5277 (N_5277,In_281,In_1913);
or U5278 (N_5278,In_2287,In_1168);
nand U5279 (N_5279,In_1328,In_2294);
nor U5280 (N_5280,In_2037,In_814);
nor U5281 (N_5281,In_41,In_233);
nand U5282 (N_5282,In_2881,In_1866);
xor U5283 (N_5283,In_1457,In_2964);
and U5284 (N_5284,In_1289,In_1600);
and U5285 (N_5285,In_1353,In_2655);
nor U5286 (N_5286,In_726,In_269);
nand U5287 (N_5287,In_1008,In_1164);
nor U5288 (N_5288,In_1110,In_1718);
nand U5289 (N_5289,In_2758,In_2656);
and U5290 (N_5290,In_24,In_1567);
or U5291 (N_5291,In_528,In_374);
or U5292 (N_5292,In_2823,In_1485);
xor U5293 (N_5293,In_316,In_2044);
and U5294 (N_5294,In_2722,In_112);
nor U5295 (N_5295,In_1773,In_893);
or U5296 (N_5296,In_866,In_2534);
nor U5297 (N_5297,In_1524,In_1133);
nand U5298 (N_5298,In_2126,In_2500);
and U5299 (N_5299,In_2643,In_2778);
or U5300 (N_5300,In_92,In_417);
and U5301 (N_5301,In_1736,In_1813);
or U5302 (N_5302,In_221,In_1490);
and U5303 (N_5303,In_2007,In_734);
nand U5304 (N_5304,In_265,In_51);
or U5305 (N_5305,In_302,In_2601);
and U5306 (N_5306,In_1992,In_2741);
or U5307 (N_5307,In_1908,In_2164);
or U5308 (N_5308,In_2362,In_1671);
nor U5309 (N_5309,In_1326,In_2433);
nand U5310 (N_5310,In_851,In_518);
and U5311 (N_5311,In_2478,In_1536);
and U5312 (N_5312,In_1506,In_591);
and U5313 (N_5313,In_448,In_369);
nor U5314 (N_5314,In_840,In_108);
nand U5315 (N_5315,In_1439,In_1845);
and U5316 (N_5316,In_1715,In_1403);
or U5317 (N_5317,In_1972,In_1563);
xnor U5318 (N_5318,In_60,In_1486);
nand U5319 (N_5319,In_1402,In_1082);
nand U5320 (N_5320,In_147,In_2558);
nand U5321 (N_5321,In_307,In_880);
nor U5322 (N_5322,In_2143,In_1293);
xnor U5323 (N_5323,In_905,In_1533);
or U5324 (N_5324,In_166,In_788);
or U5325 (N_5325,In_2629,In_71);
or U5326 (N_5326,In_2840,In_1309);
nor U5327 (N_5327,In_688,In_297);
or U5328 (N_5328,In_1813,In_2710);
nor U5329 (N_5329,In_141,In_746);
or U5330 (N_5330,In_1891,In_866);
xor U5331 (N_5331,In_1708,In_1484);
xnor U5332 (N_5332,In_966,In_1375);
and U5333 (N_5333,In_2742,In_2043);
and U5334 (N_5334,In_2103,In_12);
nor U5335 (N_5335,In_756,In_1766);
nand U5336 (N_5336,In_1779,In_594);
nand U5337 (N_5337,In_1394,In_2719);
or U5338 (N_5338,In_503,In_25);
nor U5339 (N_5339,In_1599,In_2620);
nor U5340 (N_5340,In_2515,In_643);
and U5341 (N_5341,In_214,In_1117);
xor U5342 (N_5342,In_1430,In_1111);
and U5343 (N_5343,In_2215,In_1158);
and U5344 (N_5344,In_1307,In_2464);
nand U5345 (N_5345,In_2694,In_2512);
and U5346 (N_5346,In_1041,In_2843);
nor U5347 (N_5347,In_1528,In_542);
or U5348 (N_5348,In_2130,In_2205);
xnor U5349 (N_5349,In_2505,In_1596);
or U5350 (N_5350,In_806,In_2522);
or U5351 (N_5351,In_2501,In_2032);
nor U5352 (N_5352,In_2529,In_77);
or U5353 (N_5353,In_1862,In_541);
xnor U5354 (N_5354,In_1292,In_421);
and U5355 (N_5355,In_1817,In_1912);
nor U5356 (N_5356,In_869,In_777);
or U5357 (N_5357,In_1026,In_657);
nor U5358 (N_5358,In_484,In_2126);
and U5359 (N_5359,In_2341,In_765);
and U5360 (N_5360,In_464,In_567);
nand U5361 (N_5361,In_96,In_2201);
or U5362 (N_5362,In_170,In_2531);
nand U5363 (N_5363,In_302,In_2796);
xnor U5364 (N_5364,In_576,In_2936);
nor U5365 (N_5365,In_2037,In_245);
nand U5366 (N_5366,In_864,In_2195);
nor U5367 (N_5367,In_2748,In_303);
nand U5368 (N_5368,In_567,In_2459);
or U5369 (N_5369,In_2254,In_694);
nor U5370 (N_5370,In_470,In_2065);
or U5371 (N_5371,In_2707,In_2184);
nand U5372 (N_5372,In_291,In_170);
or U5373 (N_5373,In_1964,In_2520);
nand U5374 (N_5374,In_855,In_2835);
and U5375 (N_5375,In_1389,In_873);
xor U5376 (N_5376,In_2787,In_174);
nor U5377 (N_5377,In_2668,In_1183);
or U5378 (N_5378,In_2913,In_2663);
and U5379 (N_5379,In_963,In_2370);
or U5380 (N_5380,In_1124,In_1367);
nand U5381 (N_5381,In_1050,In_1563);
or U5382 (N_5382,In_2487,In_2242);
or U5383 (N_5383,In_86,In_1459);
or U5384 (N_5384,In_2189,In_2644);
nand U5385 (N_5385,In_1427,In_299);
and U5386 (N_5386,In_998,In_2659);
and U5387 (N_5387,In_2501,In_2808);
nor U5388 (N_5388,In_1867,In_2530);
nor U5389 (N_5389,In_434,In_349);
and U5390 (N_5390,In_2970,In_2103);
and U5391 (N_5391,In_2709,In_2144);
and U5392 (N_5392,In_1401,In_2379);
nor U5393 (N_5393,In_2236,In_882);
and U5394 (N_5394,In_2132,In_1577);
and U5395 (N_5395,In_473,In_2866);
nor U5396 (N_5396,In_881,In_1584);
or U5397 (N_5397,In_938,In_1981);
or U5398 (N_5398,In_1867,In_1211);
xor U5399 (N_5399,In_156,In_1414);
and U5400 (N_5400,In_2713,In_2604);
nor U5401 (N_5401,In_1825,In_2681);
and U5402 (N_5402,In_2520,In_2705);
or U5403 (N_5403,In_2257,In_1015);
nor U5404 (N_5404,In_1213,In_1905);
nor U5405 (N_5405,In_1409,In_2529);
or U5406 (N_5406,In_341,In_187);
nand U5407 (N_5407,In_2086,In_1838);
xnor U5408 (N_5408,In_1306,In_1757);
xor U5409 (N_5409,In_2016,In_1235);
nand U5410 (N_5410,In_1285,In_941);
and U5411 (N_5411,In_1675,In_805);
or U5412 (N_5412,In_184,In_1971);
or U5413 (N_5413,In_1792,In_1390);
and U5414 (N_5414,In_1657,In_902);
and U5415 (N_5415,In_2513,In_2207);
or U5416 (N_5416,In_2519,In_2571);
and U5417 (N_5417,In_2989,In_151);
or U5418 (N_5418,In_2065,In_1795);
or U5419 (N_5419,In_1418,In_201);
nand U5420 (N_5420,In_2018,In_2796);
or U5421 (N_5421,In_2160,In_271);
or U5422 (N_5422,In_2529,In_2138);
nand U5423 (N_5423,In_1925,In_1473);
nor U5424 (N_5424,In_2770,In_1025);
nand U5425 (N_5425,In_407,In_2877);
nor U5426 (N_5426,In_1293,In_847);
or U5427 (N_5427,In_703,In_1143);
and U5428 (N_5428,In_1789,In_422);
or U5429 (N_5429,In_529,In_2067);
or U5430 (N_5430,In_758,In_1526);
nor U5431 (N_5431,In_2352,In_1415);
or U5432 (N_5432,In_737,In_63);
or U5433 (N_5433,In_41,In_2461);
or U5434 (N_5434,In_1931,In_118);
or U5435 (N_5435,In_883,In_2516);
nand U5436 (N_5436,In_2482,In_273);
xor U5437 (N_5437,In_1719,In_1531);
and U5438 (N_5438,In_1742,In_1941);
and U5439 (N_5439,In_696,In_2584);
nor U5440 (N_5440,In_1077,In_193);
nor U5441 (N_5441,In_1660,In_197);
and U5442 (N_5442,In_2402,In_1089);
or U5443 (N_5443,In_1302,In_1918);
and U5444 (N_5444,In_720,In_2070);
nand U5445 (N_5445,In_602,In_1234);
xor U5446 (N_5446,In_632,In_1260);
nand U5447 (N_5447,In_272,In_1829);
nor U5448 (N_5448,In_407,In_1448);
and U5449 (N_5449,In_1727,In_2053);
or U5450 (N_5450,In_2818,In_2061);
xnor U5451 (N_5451,In_834,In_1866);
or U5452 (N_5452,In_1579,In_2226);
nor U5453 (N_5453,In_2849,In_2738);
nand U5454 (N_5454,In_543,In_94);
xnor U5455 (N_5455,In_1291,In_779);
xor U5456 (N_5456,In_1426,In_2706);
nand U5457 (N_5457,In_1106,In_676);
nand U5458 (N_5458,In_2066,In_2447);
nor U5459 (N_5459,In_1426,In_40);
nand U5460 (N_5460,In_2579,In_1393);
and U5461 (N_5461,In_501,In_2476);
and U5462 (N_5462,In_72,In_416);
nor U5463 (N_5463,In_34,In_1799);
or U5464 (N_5464,In_2714,In_1715);
or U5465 (N_5465,In_791,In_94);
and U5466 (N_5466,In_2742,In_659);
nand U5467 (N_5467,In_922,In_1989);
nor U5468 (N_5468,In_142,In_1076);
nor U5469 (N_5469,In_2775,In_1207);
xor U5470 (N_5470,In_616,In_1331);
or U5471 (N_5471,In_1007,In_1037);
nand U5472 (N_5472,In_1983,In_1569);
or U5473 (N_5473,In_2020,In_1225);
or U5474 (N_5474,In_506,In_2164);
nor U5475 (N_5475,In_2911,In_912);
xnor U5476 (N_5476,In_2763,In_1874);
nand U5477 (N_5477,In_2010,In_2690);
or U5478 (N_5478,In_2581,In_2823);
and U5479 (N_5479,In_2420,In_2376);
or U5480 (N_5480,In_1947,In_1507);
nand U5481 (N_5481,In_1964,In_29);
and U5482 (N_5482,In_276,In_299);
xnor U5483 (N_5483,In_2883,In_1376);
and U5484 (N_5484,In_1801,In_582);
and U5485 (N_5485,In_1483,In_1218);
nand U5486 (N_5486,In_492,In_1654);
and U5487 (N_5487,In_2891,In_215);
nor U5488 (N_5488,In_2622,In_2706);
xor U5489 (N_5489,In_104,In_2342);
nand U5490 (N_5490,In_402,In_2811);
and U5491 (N_5491,In_2887,In_2881);
nor U5492 (N_5492,In_2342,In_653);
nand U5493 (N_5493,In_2598,In_2354);
and U5494 (N_5494,In_2055,In_372);
nand U5495 (N_5495,In_1550,In_1736);
xnor U5496 (N_5496,In_47,In_148);
nand U5497 (N_5497,In_1019,In_1473);
and U5498 (N_5498,In_1566,In_437);
or U5499 (N_5499,In_1610,In_1909);
nor U5500 (N_5500,In_586,In_534);
xor U5501 (N_5501,In_1826,In_2717);
or U5502 (N_5502,In_2313,In_442);
nor U5503 (N_5503,In_2379,In_486);
nor U5504 (N_5504,In_2469,In_2063);
nand U5505 (N_5505,In_1967,In_723);
nand U5506 (N_5506,In_976,In_1060);
or U5507 (N_5507,In_712,In_538);
nand U5508 (N_5508,In_689,In_2217);
or U5509 (N_5509,In_1021,In_2198);
or U5510 (N_5510,In_1181,In_2743);
and U5511 (N_5511,In_1001,In_2406);
nand U5512 (N_5512,In_1709,In_140);
and U5513 (N_5513,In_2869,In_1640);
nor U5514 (N_5514,In_806,In_2659);
or U5515 (N_5515,In_1618,In_2986);
xor U5516 (N_5516,In_1117,In_929);
nand U5517 (N_5517,In_1237,In_1088);
or U5518 (N_5518,In_382,In_2064);
xnor U5519 (N_5519,In_2665,In_2420);
or U5520 (N_5520,In_1884,In_731);
and U5521 (N_5521,In_1982,In_61);
nand U5522 (N_5522,In_199,In_794);
or U5523 (N_5523,In_2297,In_239);
or U5524 (N_5524,In_1287,In_464);
or U5525 (N_5525,In_380,In_2063);
nor U5526 (N_5526,In_112,In_2042);
or U5527 (N_5527,In_2837,In_2202);
and U5528 (N_5528,In_1011,In_62);
or U5529 (N_5529,In_2385,In_2655);
and U5530 (N_5530,In_1425,In_2681);
or U5531 (N_5531,In_319,In_802);
or U5532 (N_5532,In_1573,In_1760);
and U5533 (N_5533,In_1351,In_2421);
nor U5534 (N_5534,In_1608,In_1479);
or U5535 (N_5535,In_1111,In_237);
and U5536 (N_5536,In_745,In_2717);
nor U5537 (N_5537,In_1284,In_597);
nor U5538 (N_5538,In_2107,In_764);
and U5539 (N_5539,In_1918,In_2731);
nor U5540 (N_5540,In_58,In_713);
and U5541 (N_5541,In_579,In_2543);
and U5542 (N_5542,In_1297,In_2580);
or U5543 (N_5543,In_2836,In_1190);
and U5544 (N_5544,In_2343,In_2882);
nand U5545 (N_5545,In_686,In_2688);
nor U5546 (N_5546,In_81,In_999);
or U5547 (N_5547,In_286,In_2041);
nor U5548 (N_5548,In_535,In_384);
nand U5549 (N_5549,In_2911,In_2511);
nor U5550 (N_5550,In_2861,In_1334);
nor U5551 (N_5551,In_2155,In_1526);
or U5552 (N_5552,In_921,In_1337);
or U5553 (N_5553,In_425,In_1578);
nand U5554 (N_5554,In_2941,In_2587);
nor U5555 (N_5555,In_2142,In_1177);
and U5556 (N_5556,In_1394,In_1687);
nand U5557 (N_5557,In_274,In_1602);
nor U5558 (N_5558,In_881,In_837);
xnor U5559 (N_5559,In_176,In_758);
nor U5560 (N_5560,In_1479,In_1069);
nor U5561 (N_5561,In_2051,In_397);
or U5562 (N_5562,In_692,In_805);
or U5563 (N_5563,In_301,In_904);
and U5564 (N_5564,In_732,In_2552);
xnor U5565 (N_5565,In_1129,In_2105);
nand U5566 (N_5566,In_1363,In_1313);
nand U5567 (N_5567,In_808,In_1838);
nor U5568 (N_5568,In_704,In_1512);
xnor U5569 (N_5569,In_769,In_2471);
nand U5570 (N_5570,In_2967,In_1228);
nand U5571 (N_5571,In_2694,In_472);
nand U5572 (N_5572,In_332,In_1906);
nor U5573 (N_5573,In_1341,In_407);
or U5574 (N_5574,In_1643,In_266);
nand U5575 (N_5575,In_70,In_645);
or U5576 (N_5576,In_986,In_2117);
nand U5577 (N_5577,In_608,In_1289);
xor U5578 (N_5578,In_1561,In_574);
nor U5579 (N_5579,In_672,In_2376);
nor U5580 (N_5580,In_2116,In_2621);
xor U5581 (N_5581,In_1464,In_1173);
and U5582 (N_5582,In_1219,In_2896);
and U5583 (N_5583,In_2606,In_215);
and U5584 (N_5584,In_334,In_2851);
or U5585 (N_5585,In_2037,In_724);
and U5586 (N_5586,In_2176,In_1692);
nand U5587 (N_5587,In_1858,In_1740);
or U5588 (N_5588,In_1988,In_1580);
nand U5589 (N_5589,In_1866,In_2050);
or U5590 (N_5590,In_1085,In_1733);
and U5591 (N_5591,In_1059,In_1606);
nand U5592 (N_5592,In_982,In_2796);
nand U5593 (N_5593,In_816,In_2707);
and U5594 (N_5594,In_722,In_662);
or U5595 (N_5595,In_2680,In_2345);
or U5596 (N_5596,In_1327,In_575);
nor U5597 (N_5597,In_2195,In_651);
nor U5598 (N_5598,In_1187,In_982);
xor U5599 (N_5599,In_785,In_2440);
and U5600 (N_5600,In_868,In_605);
and U5601 (N_5601,In_5,In_2667);
nor U5602 (N_5602,In_324,In_17);
nor U5603 (N_5603,In_2602,In_2840);
and U5604 (N_5604,In_2730,In_417);
or U5605 (N_5605,In_212,In_1635);
nand U5606 (N_5606,In_2871,In_1246);
or U5607 (N_5607,In_2228,In_769);
nand U5608 (N_5608,In_2911,In_2256);
nor U5609 (N_5609,In_1608,In_2864);
nand U5610 (N_5610,In_709,In_2147);
nand U5611 (N_5611,In_1086,In_672);
nor U5612 (N_5612,In_823,In_1401);
nand U5613 (N_5613,In_161,In_2579);
nor U5614 (N_5614,In_2765,In_935);
or U5615 (N_5615,In_708,In_1858);
xor U5616 (N_5616,In_70,In_2364);
nand U5617 (N_5617,In_836,In_502);
and U5618 (N_5618,In_633,In_1380);
nor U5619 (N_5619,In_1545,In_2548);
nor U5620 (N_5620,In_2272,In_1546);
xnor U5621 (N_5621,In_1901,In_1719);
and U5622 (N_5622,In_978,In_2061);
nand U5623 (N_5623,In_1832,In_785);
nand U5624 (N_5624,In_1365,In_558);
and U5625 (N_5625,In_2040,In_861);
and U5626 (N_5626,In_2583,In_1019);
xor U5627 (N_5627,In_1322,In_1772);
nand U5628 (N_5628,In_1572,In_404);
xor U5629 (N_5629,In_844,In_2432);
xnor U5630 (N_5630,In_1643,In_2168);
or U5631 (N_5631,In_2987,In_1411);
nor U5632 (N_5632,In_837,In_2550);
nand U5633 (N_5633,In_2537,In_2500);
and U5634 (N_5634,In_2478,In_2476);
nor U5635 (N_5635,In_1351,In_779);
or U5636 (N_5636,In_2837,In_59);
nand U5637 (N_5637,In_1764,In_2912);
or U5638 (N_5638,In_1081,In_2549);
xnor U5639 (N_5639,In_2944,In_1734);
or U5640 (N_5640,In_2801,In_1373);
nand U5641 (N_5641,In_313,In_222);
nor U5642 (N_5642,In_1867,In_2472);
nor U5643 (N_5643,In_832,In_2752);
nand U5644 (N_5644,In_696,In_2108);
or U5645 (N_5645,In_2858,In_1248);
nand U5646 (N_5646,In_1578,In_2724);
nor U5647 (N_5647,In_2651,In_436);
nand U5648 (N_5648,In_1065,In_1216);
or U5649 (N_5649,In_542,In_2303);
nor U5650 (N_5650,In_1226,In_1977);
nand U5651 (N_5651,In_571,In_2837);
nand U5652 (N_5652,In_1387,In_322);
and U5653 (N_5653,In_2201,In_122);
nor U5654 (N_5654,In_2184,In_1683);
and U5655 (N_5655,In_320,In_507);
and U5656 (N_5656,In_851,In_1592);
and U5657 (N_5657,In_2126,In_2821);
nor U5658 (N_5658,In_1824,In_2177);
nand U5659 (N_5659,In_876,In_391);
and U5660 (N_5660,In_1926,In_2526);
nor U5661 (N_5661,In_283,In_2818);
or U5662 (N_5662,In_270,In_1582);
and U5663 (N_5663,In_2978,In_634);
and U5664 (N_5664,In_755,In_2022);
or U5665 (N_5665,In_1682,In_2231);
nor U5666 (N_5666,In_506,In_1539);
or U5667 (N_5667,In_1589,In_351);
nand U5668 (N_5668,In_970,In_1162);
nor U5669 (N_5669,In_1342,In_1764);
nand U5670 (N_5670,In_1113,In_2978);
or U5671 (N_5671,In_99,In_1402);
and U5672 (N_5672,In_1986,In_1140);
nand U5673 (N_5673,In_644,In_113);
nor U5674 (N_5674,In_953,In_796);
and U5675 (N_5675,In_2005,In_2986);
xor U5676 (N_5676,In_2366,In_1);
and U5677 (N_5677,In_2465,In_1223);
xnor U5678 (N_5678,In_990,In_1578);
nand U5679 (N_5679,In_1523,In_1063);
nor U5680 (N_5680,In_893,In_1100);
or U5681 (N_5681,In_927,In_1421);
nor U5682 (N_5682,In_981,In_1144);
xor U5683 (N_5683,In_404,In_1809);
nor U5684 (N_5684,In_1166,In_743);
or U5685 (N_5685,In_913,In_2492);
nand U5686 (N_5686,In_2864,In_2840);
and U5687 (N_5687,In_1956,In_800);
xor U5688 (N_5688,In_690,In_2720);
and U5689 (N_5689,In_2133,In_1236);
nand U5690 (N_5690,In_1496,In_2900);
or U5691 (N_5691,In_2559,In_689);
xnor U5692 (N_5692,In_359,In_2642);
or U5693 (N_5693,In_1826,In_68);
nor U5694 (N_5694,In_2119,In_2194);
nor U5695 (N_5695,In_1882,In_745);
nand U5696 (N_5696,In_1175,In_2115);
nor U5697 (N_5697,In_2869,In_2542);
nand U5698 (N_5698,In_37,In_937);
xor U5699 (N_5699,In_789,In_420);
nor U5700 (N_5700,In_919,In_2158);
or U5701 (N_5701,In_444,In_2069);
nor U5702 (N_5702,In_1523,In_2948);
nor U5703 (N_5703,In_2037,In_18);
and U5704 (N_5704,In_1960,In_2344);
and U5705 (N_5705,In_1820,In_2580);
or U5706 (N_5706,In_2128,In_2490);
xor U5707 (N_5707,In_1718,In_2408);
or U5708 (N_5708,In_1646,In_1176);
nand U5709 (N_5709,In_37,In_523);
nand U5710 (N_5710,In_25,In_203);
nand U5711 (N_5711,In_1793,In_342);
and U5712 (N_5712,In_504,In_2201);
and U5713 (N_5713,In_749,In_935);
nor U5714 (N_5714,In_2709,In_2218);
and U5715 (N_5715,In_2547,In_1867);
nor U5716 (N_5716,In_2532,In_1694);
and U5717 (N_5717,In_1954,In_2583);
nor U5718 (N_5718,In_1923,In_1363);
or U5719 (N_5719,In_1160,In_1281);
nor U5720 (N_5720,In_1455,In_2123);
or U5721 (N_5721,In_2030,In_889);
nand U5722 (N_5722,In_2396,In_1912);
nor U5723 (N_5723,In_2898,In_552);
and U5724 (N_5724,In_382,In_1105);
or U5725 (N_5725,In_571,In_2503);
or U5726 (N_5726,In_1596,In_2234);
and U5727 (N_5727,In_2433,In_180);
nor U5728 (N_5728,In_1113,In_1497);
xnor U5729 (N_5729,In_1653,In_2655);
and U5730 (N_5730,In_541,In_2192);
and U5731 (N_5731,In_1228,In_1863);
nand U5732 (N_5732,In_1133,In_2134);
nand U5733 (N_5733,In_2779,In_362);
nand U5734 (N_5734,In_2974,In_2024);
nand U5735 (N_5735,In_2895,In_2445);
and U5736 (N_5736,In_2565,In_2856);
nand U5737 (N_5737,In_1568,In_2874);
nand U5738 (N_5738,In_375,In_1371);
nand U5739 (N_5739,In_2930,In_631);
nand U5740 (N_5740,In_679,In_145);
nor U5741 (N_5741,In_2013,In_1808);
nor U5742 (N_5742,In_1649,In_52);
or U5743 (N_5743,In_1667,In_2228);
and U5744 (N_5744,In_2808,In_251);
nand U5745 (N_5745,In_2028,In_2484);
or U5746 (N_5746,In_2292,In_106);
nand U5747 (N_5747,In_1525,In_2968);
nand U5748 (N_5748,In_1299,In_1276);
nor U5749 (N_5749,In_2409,In_2845);
and U5750 (N_5750,In_249,In_2185);
nand U5751 (N_5751,In_1927,In_1793);
xor U5752 (N_5752,In_2106,In_589);
nor U5753 (N_5753,In_2192,In_2143);
and U5754 (N_5754,In_967,In_1221);
and U5755 (N_5755,In_2660,In_2890);
nor U5756 (N_5756,In_875,In_2586);
nor U5757 (N_5757,In_430,In_85);
and U5758 (N_5758,In_1998,In_116);
nor U5759 (N_5759,In_244,In_1445);
nand U5760 (N_5760,In_1632,In_1728);
and U5761 (N_5761,In_1830,In_1076);
xor U5762 (N_5762,In_650,In_468);
or U5763 (N_5763,In_2800,In_808);
xnor U5764 (N_5764,In_2923,In_393);
or U5765 (N_5765,In_2492,In_2037);
and U5766 (N_5766,In_383,In_307);
nand U5767 (N_5767,In_1776,In_2250);
or U5768 (N_5768,In_2455,In_2204);
or U5769 (N_5769,In_2530,In_1762);
nand U5770 (N_5770,In_2077,In_571);
and U5771 (N_5771,In_1605,In_2253);
xor U5772 (N_5772,In_1927,In_9);
nand U5773 (N_5773,In_197,In_1694);
nand U5774 (N_5774,In_1210,In_2967);
nor U5775 (N_5775,In_1307,In_2279);
nand U5776 (N_5776,In_1097,In_2307);
and U5777 (N_5777,In_1334,In_674);
and U5778 (N_5778,In_2807,In_186);
xnor U5779 (N_5779,In_1040,In_1948);
or U5780 (N_5780,In_1869,In_1835);
nand U5781 (N_5781,In_2345,In_2244);
and U5782 (N_5782,In_1366,In_805);
xor U5783 (N_5783,In_1700,In_1881);
and U5784 (N_5784,In_818,In_2678);
nand U5785 (N_5785,In_1919,In_373);
or U5786 (N_5786,In_2592,In_860);
or U5787 (N_5787,In_1889,In_1419);
or U5788 (N_5788,In_2006,In_1284);
nor U5789 (N_5789,In_867,In_1597);
or U5790 (N_5790,In_2696,In_2776);
xnor U5791 (N_5791,In_2242,In_2838);
nand U5792 (N_5792,In_2725,In_2629);
or U5793 (N_5793,In_2112,In_1955);
nor U5794 (N_5794,In_2501,In_1908);
nand U5795 (N_5795,In_64,In_2221);
or U5796 (N_5796,In_978,In_2990);
and U5797 (N_5797,In_2386,In_486);
xor U5798 (N_5798,In_426,In_2591);
or U5799 (N_5799,In_1205,In_2813);
nand U5800 (N_5800,In_1999,In_1061);
xnor U5801 (N_5801,In_1183,In_2428);
xnor U5802 (N_5802,In_1695,In_2179);
nor U5803 (N_5803,In_320,In_2825);
or U5804 (N_5804,In_2834,In_1273);
and U5805 (N_5805,In_2170,In_1534);
or U5806 (N_5806,In_2493,In_970);
nor U5807 (N_5807,In_1072,In_1610);
nor U5808 (N_5808,In_932,In_1525);
nand U5809 (N_5809,In_819,In_1638);
nor U5810 (N_5810,In_1393,In_1093);
nor U5811 (N_5811,In_1970,In_1173);
or U5812 (N_5812,In_876,In_1929);
and U5813 (N_5813,In_423,In_1222);
nand U5814 (N_5814,In_2150,In_1316);
nor U5815 (N_5815,In_1034,In_2181);
and U5816 (N_5816,In_2244,In_1408);
nand U5817 (N_5817,In_1398,In_1369);
and U5818 (N_5818,In_1624,In_1272);
and U5819 (N_5819,In_787,In_47);
nor U5820 (N_5820,In_1641,In_2113);
nor U5821 (N_5821,In_2707,In_2649);
nor U5822 (N_5822,In_1069,In_2681);
nor U5823 (N_5823,In_165,In_128);
and U5824 (N_5824,In_2886,In_2846);
nor U5825 (N_5825,In_1695,In_1610);
and U5826 (N_5826,In_1517,In_2436);
and U5827 (N_5827,In_2426,In_170);
or U5828 (N_5828,In_1145,In_1644);
or U5829 (N_5829,In_915,In_1684);
nand U5830 (N_5830,In_743,In_2191);
or U5831 (N_5831,In_2465,In_796);
and U5832 (N_5832,In_452,In_2991);
nand U5833 (N_5833,In_1009,In_533);
or U5834 (N_5834,In_2099,In_2021);
nor U5835 (N_5835,In_336,In_935);
nand U5836 (N_5836,In_491,In_106);
and U5837 (N_5837,In_2911,In_1504);
nand U5838 (N_5838,In_1322,In_854);
or U5839 (N_5839,In_794,In_257);
and U5840 (N_5840,In_681,In_1936);
nor U5841 (N_5841,In_2601,In_2849);
or U5842 (N_5842,In_1836,In_2676);
nand U5843 (N_5843,In_2196,In_2987);
nand U5844 (N_5844,In_1413,In_132);
nor U5845 (N_5845,In_2858,In_2896);
nand U5846 (N_5846,In_334,In_160);
nand U5847 (N_5847,In_754,In_2382);
nor U5848 (N_5848,In_332,In_1930);
nand U5849 (N_5849,In_2485,In_1423);
or U5850 (N_5850,In_829,In_2326);
nand U5851 (N_5851,In_1422,In_1102);
or U5852 (N_5852,In_2537,In_601);
and U5853 (N_5853,In_1250,In_2627);
xor U5854 (N_5854,In_196,In_156);
and U5855 (N_5855,In_1520,In_1772);
nand U5856 (N_5856,In_1142,In_170);
xor U5857 (N_5857,In_2073,In_1823);
nor U5858 (N_5858,In_945,In_2474);
and U5859 (N_5859,In_203,In_482);
nor U5860 (N_5860,In_1241,In_46);
or U5861 (N_5861,In_1639,In_2538);
nor U5862 (N_5862,In_354,In_2254);
nor U5863 (N_5863,In_1917,In_2966);
nand U5864 (N_5864,In_1531,In_1184);
nor U5865 (N_5865,In_56,In_2574);
or U5866 (N_5866,In_1623,In_1543);
nand U5867 (N_5867,In_1281,In_908);
nand U5868 (N_5868,In_1145,In_2063);
nor U5869 (N_5869,In_435,In_460);
nor U5870 (N_5870,In_2423,In_2043);
and U5871 (N_5871,In_2655,In_123);
xnor U5872 (N_5872,In_2780,In_537);
nand U5873 (N_5873,In_2984,In_2779);
nor U5874 (N_5874,In_340,In_1449);
nand U5875 (N_5875,In_887,In_167);
and U5876 (N_5876,In_802,In_1872);
and U5877 (N_5877,In_295,In_2738);
xnor U5878 (N_5878,In_2991,In_2954);
and U5879 (N_5879,In_267,In_711);
nand U5880 (N_5880,In_123,In_369);
or U5881 (N_5881,In_751,In_517);
or U5882 (N_5882,In_2345,In_571);
and U5883 (N_5883,In_796,In_935);
or U5884 (N_5884,In_2354,In_997);
xnor U5885 (N_5885,In_1484,In_481);
and U5886 (N_5886,In_673,In_1489);
xnor U5887 (N_5887,In_1411,In_2052);
nand U5888 (N_5888,In_1719,In_1497);
or U5889 (N_5889,In_1508,In_1824);
or U5890 (N_5890,In_2075,In_186);
and U5891 (N_5891,In_2697,In_132);
xnor U5892 (N_5892,In_359,In_2872);
nor U5893 (N_5893,In_2560,In_2477);
nor U5894 (N_5894,In_1840,In_2455);
nor U5895 (N_5895,In_1576,In_1781);
nor U5896 (N_5896,In_1404,In_286);
or U5897 (N_5897,In_359,In_1204);
and U5898 (N_5898,In_1677,In_2113);
or U5899 (N_5899,In_1714,In_197);
or U5900 (N_5900,In_2148,In_1903);
and U5901 (N_5901,In_319,In_2641);
or U5902 (N_5902,In_1025,In_1681);
or U5903 (N_5903,In_2958,In_624);
xor U5904 (N_5904,In_1355,In_140);
nor U5905 (N_5905,In_782,In_1254);
nor U5906 (N_5906,In_2109,In_1679);
nand U5907 (N_5907,In_1421,In_1548);
and U5908 (N_5908,In_1542,In_723);
xnor U5909 (N_5909,In_2575,In_1855);
nor U5910 (N_5910,In_19,In_2098);
nor U5911 (N_5911,In_2829,In_1903);
nand U5912 (N_5912,In_388,In_480);
nor U5913 (N_5913,In_2943,In_414);
xnor U5914 (N_5914,In_233,In_101);
nor U5915 (N_5915,In_39,In_2073);
nand U5916 (N_5916,In_435,In_1082);
nand U5917 (N_5917,In_2007,In_1840);
xnor U5918 (N_5918,In_2237,In_1194);
nand U5919 (N_5919,In_1748,In_144);
nand U5920 (N_5920,In_1138,In_1258);
and U5921 (N_5921,In_2568,In_588);
nand U5922 (N_5922,In_2293,In_841);
xor U5923 (N_5923,In_1602,In_645);
and U5924 (N_5924,In_1958,In_255);
nand U5925 (N_5925,In_1702,In_1257);
nand U5926 (N_5926,In_1116,In_1777);
xnor U5927 (N_5927,In_2403,In_829);
xor U5928 (N_5928,In_2494,In_1233);
or U5929 (N_5929,In_2440,In_544);
xnor U5930 (N_5930,In_808,In_175);
nand U5931 (N_5931,In_1352,In_1953);
xor U5932 (N_5932,In_2235,In_2978);
xnor U5933 (N_5933,In_701,In_1328);
nand U5934 (N_5934,In_2068,In_2515);
or U5935 (N_5935,In_1144,In_428);
or U5936 (N_5936,In_1244,In_2131);
nand U5937 (N_5937,In_406,In_1249);
nand U5938 (N_5938,In_586,In_1031);
nand U5939 (N_5939,In_1447,In_1739);
nand U5940 (N_5940,In_1040,In_99);
and U5941 (N_5941,In_294,In_432);
nor U5942 (N_5942,In_2425,In_563);
nand U5943 (N_5943,In_856,In_1489);
and U5944 (N_5944,In_2076,In_2805);
and U5945 (N_5945,In_1530,In_2121);
nor U5946 (N_5946,In_2863,In_2395);
or U5947 (N_5947,In_603,In_2120);
and U5948 (N_5948,In_1641,In_2438);
and U5949 (N_5949,In_4,In_2250);
or U5950 (N_5950,In_2027,In_1599);
xnor U5951 (N_5951,In_2581,In_1038);
nand U5952 (N_5952,In_2060,In_891);
xor U5953 (N_5953,In_2258,In_2311);
or U5954 (N_5954,In_1921,In_2665);
or U5955 (N_5955,In_177,In_50);
nor U5956 (N_5956,In_418,In_1192);
nor U5957 (N_5957,In_1715,In_488);
nand U5958 (N_5958,In_957,In_889);
nand U5959 (N_5959,In_2028,In_504);
or U5960 (N_5960,In_488,In_2735);
nor U5961 (N_5961,In_2587,In_690);
or U5962 (N_5962,In_636,In_1356);
xor U5963 (N_5963,In_647,In_1366);
or U5964 (N_5964,In_1901,In_2756);
nor U5965 (N_5965,In_1750,In_334);
nand U5966 (N_5966,In_990,In_1596);
nor U5967 (N_5967,In_880,In_1140);
nand U5968 (N_5968,In_2806,In_1225);
or U5969 (N_5969,In_1027,In_148);
and U5970 (N_5970,In_312,In_2342);
or U5971 (N_5971,In_1053,In_743);
and U5972 (N_5972,In_2171,In_648);
xor U5973 (N_5973,In_2110,In_1572);
nor U5974 (N_5974,In_1717,In_539);
nor U5975 (N_5975,In_2299,In_536);
nor U5976 (N_5976,In_282,In_1293);
nor U5977 (N_5977,In_915,In_2747);
and U5978 (N_5978,In_2178,In_930);
nand U5979 (N_5979,In_1091,In_2761);
xor U5980 (N_5980,In_2213,In_339);
or U5981 (N_5981,In_2793,In_713);
xnor U5982 (N_5982,In_753,In_1849);
or U5983 (N_5983,In_1281,In_2983);
xor U5984 (N_5984,In_2433,In_954);
nand U5985 (N_5985,In_2768,In_1872);
nand U5986 (N_5986,In_2945,In_28);
or U5987 (N_5987,In_1128,In_2559);
or U5988 (N_5988,In_1362,In_1231);
xor U5989 (N_5989,In_1366,In_1168);
nor U5990 (N_5990,In_1278,In_1015);
xor U5991 (N_5991,In_2176,In_1471);
or U5992 (N_5992,In_669,In_1997);
xnor U5993 (N_5993,In_706,In_2606);
nor U5994 (N_5994,In_1420,In_1749);
nand U5995 (N_5995,In_2242,In_627);
or U5996 (N_5996,In_115,In_1746);
or U5997 (N_5997,In_1414,In_157);
and U5998 (N_5998,In_2435,In_503);
or U5999 (N_5999,In_1786,In_462);
nand U6000 (N_6000,N_2774,N_3569);
xnor U6001 (N_6001,N_2968,N_5155);
and U6002 (N_6002,N_5816,N_4982);
xor U6003 (N_6003,N_1887,N_2770);
nand U6004 (N_6004,N_4257,N_3379);
or U6005 (N_6005,N_3499,N_1951);
nor U6006 (N_6006,N_2105,N_4395);
or U6007 (N_6007,N_3907,N_3700);
nand U6008 (N_6008,N_508,N_2451);
or U6009 (N_6009,N_5096,N_1561);
and U6010 (N_6010,N_4442,N_4373);
xnor U6011 (N_6011,N_324,N_3781);
xor U6012 (N_6012,N_261,N_4151);
xnor U6013 (N_6013,N_5344,N_245);
nor U6014 (N_6014,N_4631,N_3215);
nor U6015 (N_6015,N_4954,N_4902);
nor U6016 (N_6016,N_1944,N_3234);
xnor U6017 (N_6017,N_513,N_711);
xor U6018 (N_6018,N_1822,N_5480);
and U6019 (N_6019,N_3971,N_672);
and U6020 (N_6020,N_370,N_3484);
or U6021 (N_6021,N_4052,N_5970);
and U6022 (N_6022,N_489,N_3862);
or U6023 (N_6023,N_3718,N_1515);
or U6024 (N_6024,N_506,N_4076);
and U6025 (N_6025,N_2398,N_2741);
or U6026 (N_6026,N_4108,N_3985);
xnor U6027 (N_6027,N_2038,N_2169);
or U6028 (N_6028,N_3029,N_1262);
and U6029 (N_6029,N_1149,N_1734);
and U6030 (N_6030,N_2193,N_154);
xnor U6031 (N_6031,N_1024,N_956);
nor U6032 (N_6032,N_4859,N_1701);
nand U6033 (N_6033,N_1147,N_3799);
or U6034 (N_6034,N_93,N_1236);
xnor U6035 (N_6035,N_1600,N_3310);
and U6036 (N_6036,N_2997,N_1512);
nor U6037 (N_6037,N_2118,N_697);
nand U6038 (N_6038,N_4718,N_1835);
and U6039 (N_6039,N_5527,N_5929);
nor U6040 (N_6040,N_1911,N_1322);
and U6041 (N_6041,N_1736,N_3595);
or U6042 (N_6042,N_1391,N_1837);
nor U6043 (N_6043,N_4586,N_4966);
and U6044 (N_6044,N_1195,N_5773);
nor U6045 (N_6045,N_5073,N_4223);
nand U6046 (N_6046,N_5758,N_5931);
nand U6047 (N_6047,N_2361,N_4126);
and U6048 (N_6048,N_2493,N_3691);
xnor U6049 (N_6049,N_671,N_4240);
and U6050 (N_6050,N_2656,N_4087);
nor U6051 (N_6051,N_1796,N_2221);
and U6052 (N_6052,N_1498,N_3976);
nand U6053 (N_6053,N_3301,N_2295);
nor U6054 (N_6054,N_4561,N_2133);
nor U6055 (N_6055,N_1163,N_838);
nor U6056 (N_6056,N_275,N_1888);
or U6057 (N_6057,N_186,N_4577);
nor U6058 (N_6058,N_2478,N_5168);
nand U6059 (N_6059,N_2257,N_3184);
and U6060 (N_6060,N_2313,N_5319);
or U6061 (N_6061,N_4740,N_2387);
nor U6062 (N_6062,N_754,N_1042);
nor U6063 (N_6063,N_880,N_5616);
or U6064 (N_6064,N_5276,N_3317);
or U6065 (N_6065,N_1665,N_440);
nand U6066 (N_6066,N_2114,N_5373);
xnor U6067 (N_6067,N_4035,N_771);
or U6068 (N_6068,N_2297,N_906);
xnor U6069 (N_6069,N_2877,N_4206);
and U6070 (N_6070,N_3536,N_3399);
nand U6071 (N_6071,N_1965,N_5347);
and U6072 (N_6072,N_2823,N_4285);
or U6073 (N_6073,N_3991,N_929);
xor U6074 (N_6074,N_528,N_3303);
nor U6075 (N_6075,N_5998,N_3954);
nor U6076 (N_6076,N_4433,N_2423);
and U6077 (N_6077,N_4043,N_5224);
or U6078 (N_6078,N_3992,N_5165);
or U6079 (N_6079,N_2164,N_5464);
or U6080 (N_6080,N_1064,N_410);
or U6081 (N_6081,N_2380,N_4644);
nand U6082 (N_6082,N_2690,N_1811);
xor U6083 (N_6083,N_4999,N_4268);
nand U6084 (N_6084,N_5129,N_848);
nor U6085 (N_6085,N_156,N_5380);
or U6086 (N_6086,N_1778,N_5580);
nor U6087 (N_6087,N_195,N_2068);
nand U6088 (N_6088,N_120,N_2177);
nand U6089 (N_6089,N_1553,N_2476);
and U6090 (N_6090,N_3256,N_428);
or U6091 (N_6091,N_4283,N_2559);
nor U6092 (N_6092,N_3441,N_1999);
nor U6093 (N_6093,N_5561,N_2132);
or U6094 (N_6094,N_3151,N_1641);
nand U6095 (N_6095,N_3863,N_5353);
nand U6096 (N_6096,N_5338,N_586);
nand U6097 (N_6097,N_3274,N_5571);
xnor U6098 (N_6098,N_3012,N_3244);
nand U6099 (N_6099,N_3933,N_4178);
nand U6100 (N_6100,N_4830,N_5633);
or U6101 (N_6101,N_4014,N_218);
nand U6102 (N_6102,N_2332,N_3621);
and U6103 (N_6103,N_243,N_4416);
nor U6104 (N_6104,N_2383,N_3989);
nand U6105 (N_6105,N_4272,N_2874);
nor U6106 (N_6106,N_137,N_5667);
xnor U6107 (N_6107,N_4277,N_4389);
or U6108 (N_6108,N_4393,N_5010);
nor U6109 (N_6109,N_607,N_3706);
nor U6110 (N_6110,N_95,N_2236);
nor U6111 (N_6111,N_2319,N_5268);
and U6112 (N_6112,N_4513,N_5292);
and U6113 (N_6113,N_5585,N_2856);
or U6114 (N_6114,N_2722,N_4004);
or U6115 (N_6115,N_3305,N_3028);
or U6116 (N_6116,N_5107,N_994);
nand U6117 (N_6117,N_1976,N_1052);
and U6118 (N_6118,N_5932,N_3020);
nand U6119 (N_6119,N_4689,N_3808);
xor U6120 (N_6120,N_16,N_4048);
nor U6121 (N_6121,N_1463,N_3771);
nand U6122 (N_6122,N_64,N_5671);
nor U6123 (N_6123,N_1536,N_1000);
nor U6124 (N_6124,N_3659,N_5649);
nand U6125 (N_6125,N_2106,N_5574);
and U6126 (N_6126,N_2063,N_5367);
xnor U6127 (N_6127,N_2778,N_5974);
and U6128 (N_6128,N_866,N_2944);
or U6129 (N_6129,N_1510,N_2702);
and U6130 (N_6130,N_1291,N_4308);
xnor U6131 (N_6131,N_5050,N_5769);
and U6132 (N_6132,N_5053,N_290);
and U6133 (N_6133,N_3173,N_2458);
and U6134 (N_6134,N_1191,N_2090);
xnor U6135 (N_6135,N_5074,N_1547);
nor U6136 (N_6136,N_3607,N_1281);
nor U6137 (N_6137,N_4419,N_3883);
nor U6138 (N_6138,N_2216,N_4782);
nand U6139 (N_6139,N_3237,N_2397);
nor U6140 (N_6140,N_5166,N_4520);
nand U6141 (N_6141,N_669,N_2125);
nor U6142 (N_6142,N_5676,N_3372);
and U6143 (N_6143,N_1789,N_4376);
or U6144 (N_6144,N_5781,N_222);
nor U6145 (N_6145,N_2178,N_1856);
xnor U6146 (N_6146,N_437,N_1678);
or U6147 (N_6147,N_91,N_259);
nor U6148 (N_6148,N_4017,N_3642);
nor U6149 (N_6149,N_3362,N_656);
xnor U6150 (N_6150,N_3331,N_3852);
nor U6151 (N_6151,N_5807,N_3913);
xnor U6152 (N_6152,N_2291,N_279);
xor U6153 (N_6153,N_1632,N_1174);
nor U6154 (N_6154,N_2697,N_1823);
xor U6155 (N_6155,N_3214,N_901);
or U6156 (N_6156,N_152,N_232);
and U6157 (N_6157,N_1494,N_4305);
or U6158 (N_6158,N_2678,N_1915);
and U6159 (N_6159,N_2223,N_5337);
nand U6160 (N_6160,N_4614,N_2735);
nor U6161 (N_6161,N_2886,N_1245);
or U6162 (N_6162,N_515,N_5288);
or U6163 (N_6163,N_2718,N_5463);
or U6164 (N_6164,N_3397,N_5919);
or U6165 (N_6165,N_1263,N_1090);
and U6166 (N_6166,N_2645,N_1253);
nor U6167 (N_6167,N_3754,N_449);
or U6168 (N_6168,N_2440,N_971);
or U6169 (N_6169,N_4665,N_5994);
xnor U6170 (N_6170,N_3377,N_4224);
nand U6171 (N_6171,N_185,N_1629);
or U6172 (N_6172,N_3597,N_2467);
and U6173 (N_6173,N_1587,N_5468);
xor U6174 (N_6174,N_2173,N_1862);
xor U6175 (N_6175,N_2660,N_3473);
nand U6176 (N_6176,N_383,N_5721);
xnor U6177 (N_6177,N_1220,N_2315);
or U6178 (N_6178,N_2468,N_4836);
nand U6179 (N_6179,N_1098,N_1389);
nand U6180 (N_6180,N_2352,N_5806);
nor U6181 (N_6181,N_1443,N_2519);
and U6182 (N_6182,N_5724,N_3627);
nor U6183 (N_6183,N_1797,N_3326);
or U6184 (N_6184,N_433,N_3601);
nor U6185 (N_6185,N_720,N_2055);
nor U6186 (N_6186,N_4526,N_1084);
or U6187 (N_6187,N_3292,N_1320);
or U6188 (N_6188,N_381,N_102);
xnor U6189 (N_6189,N_2996,N_447);
nand U6190 (N_6190,N_1208,N_2160);
nand U6191 (N_6191,N_2547,N_3955);
and U6192 (N_6192,N_1673,N_4077);
or U6193 (N_6193,N_4845,N_3636);
nand U6194 (N_6194,N_5392,N_1182);
or U6195 (N_6195,N_4847,N_3118);
and U6196 (N_6196,N_3919,N_902);
or U6197 (N_6197,N_3130,N_2862);
xnor U6198 (N_6198,N_2681,N_2542);
nor U6199 (N_6199,N_655,N_4085);
or U6200 (N_6200,N_4487,N_2564);
nand U6201 (N_6201,N_1524,N_1286);
nor U6202 (N_6202,N_1214,N_1584);
nor U6203 (N_6203,N_5350,N_1046);
nand U6204 (N_6204,N_5264,N_3894);
nor U6205 (N_6205,N_89,N_4167);
and U6206 (N_6206,N_4230,N_446);
xor U6207 (N_6207,N_2769,N_594);
and U6208 (N_6208,N_4121,N_925);
nand U6209 (N_6209,N_3015,N_1941);
nor U6210 (N_6210,N_764,N_1590);
and U6211 (N_6211,N_373,N_5871);
and U6212 (N_6212,N_4949,N_5613);
and U6213 (N_6213,N_2835,N_1066);
and U6214 (N_6214,N_5051,N_3916);
nor U6215 (N_6215,N_556,N_3680);
or U6216 (N_6216,N_3364,N_1407);
or U6217 (N_6217,N_2158,N_2616);
and U6218 (N_6218,N_530,N_1522);
or U6219 (N_6219,N_219,N_2203);
nand U6220 (N_6220,N_3671,N_3175);
and U6221 (N_6221,N_5853,N_2736);
and U6222 (N_6222,N_4371,N_5301);
xnor U6223 (N_6223,N_3177,N_1851);
nand U6224 (N_6224,N_3103,N_661);
and U6225 (N_6225,N_5248,N_98);
nand U6226 (N_6226,N_2095,N_5785);
nand U6227 (N_6227,N_3327,N_3287);
and U6228 (N_6228,N_3267,N_3747);
and U6229 (N_6229,N_2435,N_5735);
nor U6230 (N_6230,N_3762,N_3199);
nor U6231 (N_6231,N_2930,N_3942);
or U6232 (N_6232,N_4838,N_3587);
and U6233 (N_6233,N_5489,N_972);
or U6234 (N_6234,N_517,N_1015);
nor U6235 (N_6235,N_2958,N_5918);
nand U6236 (N_6236,N_5397,N_5928);
or U6237 (N_6237,N_5855,N_5954);
nor U6238 (N_6238,N_496,N_1907);
or U6239 (N_6239,N_1259,N_5500);
and U6240 (N_6240,N_574,N_3937);
nand U6241 (N_6241,N_1966,N_5425);
and U6242 (N_6242,N_1767,N_4539);
and U6243 (N_6243,N_4199,N_1696);
and U6244 (N_6244,N_307,N_5626);
or U6245 (N_6245,N_2641,N_2649);
xor U6246 (N_6246,N_2721,N_4327);
and U6247 (N_6247,N_898,N_1857);
and U6248 (N_6248,N_341,N_1591);
nand U6249 (N_6249,N_2781,N_634);
or U6250 (N_6250,N_1981,N_5535);
nor U6251 (N_6251,N_1959,N_3092);
nand U6252 (N_6252,N_4291,N_3926);
xor U6253 (N_6253,N_5587,N_2911);
or U6254 (N_6254,N_3498,N_5450);
nor U6255 (N_6255,N_5222,N_418);
nand U6256 (N_6256,N_4320,N_5056);
nor U6257 (N_6257,N_2929,N_4863);
and U6258 (N_6258,N_3827,N_1809);
xnor U6259 (N_6259,N_724,N_4955);
nand U6260 (N_6260,N_1520,N_4338);
or U6261 (N_6261,N_4464,N_4959);
and U6262 (N_6262,N_5543,N_419);
xnor U6263 (N_6263,N_4325,N_651);
and U6264 (N_6264,N_984,N_317);
or U6265 (N_6265,N_1563,N_738);
nor U6266 (N_6266,N_1631,N_3519);
and U6267 (N_6267,N_1717,N_1481);
xor U6268 (N_6268,N_4703,N_12);
and U6269 (N_6269,N_4720,N_3152);
or U6270 (N_6270,N_1122,N_1283);
or U6271 (N_6271,N_4647,N_2019);
nand U6272 (N_6272,N_945,N_2142);
nor U6273 (N_6273,N_5790,N_2524);
nand U6274 (N_6274,N_4624,N_3133);
and U6275 (N_6275,N_2964,N_2923);
or U6276 (N_6276,N_930,N_3759);
and U6277 (N_6277,N_2138,N_2116);
or U6278 (N_6278,N_4792,N_2648);
and U6279 (N_6279,N_361,N_2516);
nor U6280 (N_6280,N_1307,N_3067);
nand U6281 (N_6281,N_2231,N_3162);
nor U6282 (N_6282,N_1244,N_3163);
nand U6283 (N_6283,N_1518,N_4580);
or U6284 (N_6284,N_286,N_4221);
nor U6285 (N_6285,N_3577,N_5739);
or U6286 (N_6286,N_118,N_3651);
nand U6287 (N_6287,N_3227,N_2786);
xnor U6288 (N_6288,N_5369,N_3285);
or U6289 (N_6289,N_4364,N_3102);
xnor U6290 (N_6290,N_5095,N_3840);
and U6291 (N_6291,N_3279,N_4552);
nand U6292 (N_6292,N_783,N_2717);
nand U6293 (N_6293,N_1499,N_2359);
or U6294 (N_6294,N_2746,N_2633);
and U6295 (N_6295,N_4073,N_179);
and U6296 (N_6296,N_1628,N_4686);
xnor U6297 (N_6297,N_2758,N_2011);
xnor U6298 (N_6298,N_728,N_3570);
or U6299 (N_6299,N_2634,N_5726);
xor U6300 (N_6300,N_5779,N_3145);
and U6301 (N_6301,N_991,N_97);
nor U6302 (N_6302,N_125,N_1788);
or U6303 (N_6303,N_1771,N_694);
nor U6304 (N_6304,N_2002,N_4040);
and U6305 (N_6305,N_2224,N_453);
or U6306 (N_6306,N_675,N_1432);
xnor U6307 (N_6307,N_2909,N_3996);
nor U6308 (N_6308,N_5081,N_426);
nor U6309 (N_6309,N_1740,N_5737);
nand U6310 (N_6310,N_2,N_2321);
xor U6311 (N_6311,N_3861,N_3746);
nand U6312 (N_6312,N_2395,N_4738);
or U6313 (N_6313,N_4994,N_4544);
xnor U6314 (N_6314,N_1721,N_1990);
or U6315 (N_6315,N_490,N_3450);
nand U6316 (N_6316,N_2671,N_4569);
nand U6317 (N_6317,N_5239,N_4839);
nand U6318 (N_6318,N_1511,N_5317);
xor U6319 (N_6319,N_5219,N_4033);
or U6320 (N_6320,N_4091,N_4555);
nand U6321 (N_6321,N_438,N_2829);
nor U6322 (N_6322,N_1528,N_3668);
and U6323 (N_6323,N_4719,N_313);
nor U6324 (N_6324,N_699,N_1836);
nand U6325 (N_6325,N_157,N_1424);
or U6326 (N_6326,N_1593,N_1056);
nand U6327 (N_6327,N_5874,N_3442);
nor U6328 (N_6328,N_2016,N_3334);
nand U6329 (N_6329,N_3692,N_3393);
and U6330 (N_6330,N_4542,N_5206);
or U6331 (N_6331,N_105,N_2014);
xor U6332 (N_6332,N_3705,N_209);
nor U6333 (N_6333,N_595,N_3972);
nor U6334 (N_6334,N_4559,N_4797);
or U6335 (N_6335,N_1950,N_4940);
nand U6336 (N_6336,N_534,N_4791);
and U6337 (N_6337,N_1114,N_4412);
nor U6338 (N_6338,N_2333,N_1685);
nor U6339 (N_6339,N_3282,N_284);
and U6340 (N_6340,N_5304,N_2851);
nand U6341 (N_6341,N_1640,N_2639);
xnor U6342 (N_6342,N_4896,N_5348);
or U6343 (N_6343,N_1725,N_1359);
xor U6344 (N_6344,N_849,N_2327);
and U6345 (N_6345,N_619,N_4913);
or U6346 (N_6346,N_4801,N_3887);
and U6347 (N_6347,N_1843,N_4);
or U6348 (N_6348,N_584,N_3774);
xnor U6349 (N_6349,N_5287,N_5009);
xnor U6350 (N_6350,N_4168,N_5223);
nor U6351 (N_6351,N_2689,N_5329);
nand U6352 (N_6352,N_5914,N_5523);
nor U6353 (N_6353,N_5154,N_4022);
xor U6354 (N_6354,N_3854,N_1746);
and U6355 (N_6355,N_363,N_2370);
or U6356 (N_6356,N_2674,N_4027);
or U6357 (N_6357,N_737,N_958);
or U6358 (N_6358,N_226,N_3660);
and U6359 (N_6359,N_431,N_3245);
and U6360 (N_6360,N_5831,N_1068);
and U6361 (N_6361,N_2554,N_1844);
nand U6362 (N_6362,N_524,N_890);
nor U6363 (N_6363,N_2187,N_487);
nand U6364 (N_6364,N_2442,N_5236);
nand U6365 (N_6365,N_2783,N_2777);
and U6366 (N_6366,N_4106,N_1394);
nand U6367 (N_6367,N_1410,N_4591);
xnor U6368 (N_6368,N_5457,N_1850);
and U6369 (N_6369,N_3206,N_1526);
nand U6370 (N_6370,N_5267,N_2831);
and U6371 (N_6371,N_356,N_1702);
and U6372 (N_6372,N_4177,N_2948);
and U6373 (N_6373,N_4273,N_1110);
or U6374 (N_6374,N_1660,N_4629);
nor U6375 (N_6375,N_1969,N_5185);
and U6376 (N_6376,N_1830,N_4758);
xor U6377 (N_6377,N_4165,N_2131);
nor U6378 (N_6378,N_2389,N_2740);
or U6379 (N_6379,N_4554,N_4226);
or U6380 (N_6380,N_4096,N_2161);
or U6381 (N_6381,N_3154,N_2157);
and U6382 (N_6382,N_4140,N_2136);
or U6383 (N_6383,N_2506,N_1032);
or U6384 (N_6384,N_3786,N_597);
nor U6385 (N_6385,N_1689,N_5621);
nand U6386 (N_6386,N_71,N_3134);
xor U6387 (N_6387,N_4438,N_1560);
nand U6388 (N_6388,N_1842,N_2119);
and U6389 (N_6389,N_4279,N_1081);
or U6390 (N_6390,N_3731,N_2284);
nor U6391 (N_6391,N_109,N_633);
nand U6392 (N_6392,N_626,N_5844);
nand U6393 (N_6393,N_5557,N_3348);
nand U6394 (N_6394,N_384,N_3796);
or U6395 (N_6395,N_1403,N_5151);
nor U6396 (N_6396,N_4060,N_1080);
nor U6397 (N_6397,N_3611,N_1412);
and U6398 (N_6398,N_5340,N_3449);
nor U6399 (N_6399,N_5474,N_3192);
or U6400 (N_6400,N_4095,N_2710);
nor U6401 (N_6401,N_3221,N_1203);
and U6402 (N_6402,N_2898,N_5765);
or U6403 (N_6403,N_2447,N_5092);
nand U6404 (N_6404,N_1930,N_5868);
and U6405 (N_6405,N_4590,N_5537);
and U6406 (N_6406,N_3249,N_5659);
nand U6407 (N_6407,N_1974,N_1742);
xnor U6408 (N_6408,N_3204,N_1482);
nand U6409 (N_6409,N_5182,N_2043);
and U6410 (N_6410,N_910,N_5840);
nor U6411 (N_6411,N_2679,N_5863);
or U6412 (N_6412,N_368,N_1272);
nand U6413 (N_6413,N_1460,N_935);
and U6414 (N_6414,N_5406,N_294);
nor U6415 (N_6415,N_2743,N_562);
nand U6416 (N_6416,N_5478,N_962);
and U6417 (N_6417,N_2238,N_2797);
xnor U6418 (N_6418,N_5157,N_3620);
nand U6419 (N_6419,N_5709,N_1910);
nand U6420 (N_6420,N_3727,N_3023);
nand U6421 (N_6421,N_4734,N_570);
nor U6422 (N_6422,N_2446,N_2403);
xnor U6423 (N_6423,N_141,N_4485);
nand U6424 (N_6424,N_1365,N_3444);
xnor U6425 (N_6425,N_4039,N_1293);
xor U6426 (N_6426,N_3782,N_283);
or U6427 (N_6427,N_772,N_3041);
and U6428 (N_6428,N_4363,N_2842);
xor U6429 (N_6429,N_4957,N_2659);
nand U6430 (N_6430,N_3375,N_1353);
or U6431 (N_6431,N_3522,N_2404);
and U6432 (N_6432,N_4680,N_3784);
nand U6433 (N_6433,N_3385,N_571);
or U6434 (N_6434,N_5303,N_2704);
nor U6435 (N_6435,N_150,N_11);
and U6436 (N_6436,N_4079,N_808);
nand U6437 (N_6437,N_3349,N_1366);
and U6438 (N_6438,N_3477,N_4050);
and U6439 (N_6439,N_638,N_2381);
and U6440 (N_6440,N_2599,N_5699);
or U6441 (N_6441,N_4993,N_740);
nor U6442 (N_6442,N_3612,N_2727);
nand U6443 (N_6443,N_1176,N_4191);
or U6444 (N_6444,N_3286,N_5714);
nand U6445 (N_6445,N_3936,N_2215);
nand U6446 (N_6446,N_3157,N_189);
nor U6447 (N_6447,N_2347,N_5240);
and U6448 (N_6448,N_2903,N_2271);
and U6449 (N_6449,N_602,N_3677);
xor U6450 (N_6450,N_457,N_2809);
or U6451 (N_6451,N_2076,N_2578);
and U6452 (N_6452,N_2981,N_338);
nand U6453 (N_6453,N_5112,N_2812);
and U6454 (N_6454,N_4075,N_2501);
and U6455 (N_6455,N_436,N_3277);
and U6456 (N_6456,N_2957,N_1417);
nor U6457 (N_6457,N_4548,N_4944);
nor U6458 (N_6458,N_3436,N_5972);
nand U6459 (N_6459,N_3432,N_4046);
and U6460 (N_6460,N_2179,N_2220);
nand U6461 (N_6461,N_5087,N_5901);
nor U6462 (N_6462,N_2463,N_4744);
or U6463 (N_6463,N_5647,N_1817);
xor U6464 (N_6464,N_4349,N_642);
xor U6465 (N_6465,N_2392,N_2228);
nand U6466 (N_6466,N_4258,N_3054);
or U6467 (N_6467,N_2343,N_5801);
or U6468 (N_6468,N_2026,N_2646);
nor U6469 (N_6469,N_4546,N_2785);
nand U6470 (N_6470,N_2162,N_4960);
nand U6471 (N_6471,N_4390,N_2642);
nand U6472 (N_6472,N_3521,N_2844);
nor U6473 (N_6473,N_566,N_5221);
or U6474 (N_6474,N_163,N_1221);
nand U6475 (N_6475,N_3914,N_4294);
or U6476 (N_6476,N_1962,N_4741);
nand U6477 (N_6477,N_927,N_1855);
nand U6478 (N_6478,N_1312,N_107);
and U6479 (N_6479,N_3859,N_588);
nand U6480 (N_6480,N_1783,N_3243);
and U6481 (N_6481,N_405,N_3117);
or U6482 (N_6482,N_1405,N_4746);
nand U6483 (N_6483,N_1300,N_550);
nand U6484 (N_6484,N_5387,N_1464);
or U6485 (N_6485,N_76,N_5124);
or U6486 (N_6486,N_3688,N_300);
or U6487 (N_6487,N_1813,N_4385);
nor U6488 (N_6488,N_1202,N_2569);
nor U6489 (N_6489,N_1519,N_4187);
and U6490 (N_6490,N_3230,N_4301);
nor U6491 (N_6491,N_3033,N_5728);
and U6492 (N_6492,N_4831,N_2412);
and U6493 (N_6493,N_18,N_2018);
nand U6494 (N_6494,N_5141,N_2061);
or U6495 (N_6495,N_51,N_208);
nor U6496 (N_6496,N_4372,N_4929);
nor U6497 (N_6497,N_1853,N_640);
nor U6498 (N_6498,N_4074,N_5685);
nor U6499 (N_6499,N_158,N_576);
and U6500 (N_6500,N_1765,N_4775);
nor U6501 (N_6501,N_3401,N_666);
or U6502 (N_6502,N_1358,N_860);
nand U6503 (N_6503,N_5725,N_1957);
and U6504 (N_6504,N_2023,N_3143);
or U6505 (N_6505,N_5183,N_4426);
nand U6506 (N_6506,N_1328,N_1825);
nand U6507 (N_6507,N_2062,N_2239);
nand U6508 (N_6508,N_1532,N_27);
nor U6509 (N_6509,N_4638,N_5456);
or U6510 (N_6510,N_2730,N_5983);
xnor U6511 (N_6511,N_1728,N_520);
nand U6512 (N_6512,N_1497,N_2635);
xnor U6513 (N_6513,N_3482,N_790);
nor U6514 (N_6514,N_1785,N_4933);
nor U6515 (N_6515,N_493,N_2008);
nand U6516 (N_6516,N_2184,N_3783);
xnor U6517 (N_6517,N_2950,N_657);
nor U6518 (N_6518,N_1034,N_519);
and U6519 (N_6519,N_4653,N_1192);
nor U6520 (N_6520,N_1917,N_1050);
nor U6521 (N_6521,N_2512,N_5388);
or U6522 (N_6522,N_2492,N_4890);
and U6523 (N_6523,N_575,N_3407);
nor U6524 (N_6524,N_70,N_2796);
nand U6525 (N_6525,N_2310,N_5390);
nor U6526 (N_6526,N_2692,N_5110);
or U6527 (N_6527,N_5153,N_5933);
xnor U6528 (N_6528,N_4018,N_1798);
nor U6529 (N_6529,N_4784,N_4306);
nor U6530 (N_6530,N_5532,N_999);
xnor U6531 (N_6531,N_2604,N_4229);
and U6532 (N_6532,N_2110,N_5436);
or U6533 (N_6533,N_2762,N_5608);
nand U6534 (N_6534,N_820,N_3107);
nand U6535 (N_6535,N_3193,N_3088);
nand U6536 (N_6536,N_913,N_5357);
and U6537 (N_6537,N_2059,N_5672);
or U6538 (N_6538,N_4934,N_475);
nor U6539 (N_6539,N_4522,N_5910);
and U6540 (N_6540,N_4783,N_1228);
nor U6541 (N_6541,N_1466,N_5911);
and U6542 (N_6542,N_5627,N_5798);
xnor U6543 (N_6543,N_686,N_3584);
and U6544 (N_6544,N_2300,N_4967);
or U6545 (N_6545,N_2498,N_4440);
or U6546 (N_6546,N_5383,N_2643);
or U6547 (N_6547,N_2305,N_5916);
nand U6548 (N_6548,N_3613,N_2414);
xor U6549 (N_6549,N_630,N_2376);
xnor U6550 (N_6550,N_3608,N_4058);
or U6551 (N_6551,N_4418,N_4000);
nor U6552 (N_6552,N_3344,N_2871);
nor U6553 (N_6553,N_1691,N_623);
nand U6554 (N_6554,N_5604,N_1495);
nor U6555 (N_6555,N_775,N_231);
nand U6556 (N_6556,N_5760,N_1883);
nand U6557 (N_6557,N_643,N_422);
or U6558 (N_6558,N_5443,N_4458);
nor U6559 (N_6559,N_4928,N_5615);
nand U6560 (N_6560,N_5515,N_2406);
and U6561 (N_6561,N_4563,N_3342);
or U6562 (N_6562,N_522,N_4492);
nor U6563 (N_6563,N_767,N_1304);
or U6564 (N_6564,N_2920,N_3864);
xor U6565 (N_6565,N_1155,N_14);
or U6566 (N_6566,N_3022,N_5651);
or U6567 (N_6567,N_1653,N_3106);
and U6568 (N_6568,N_1093,N_563);
or U6569 (N_6569,N_2808,N_1535);
nor U6570 (N_6570,N_451,N_5597);
nand U6571 (N_6571,N_4297,N_59);
nand U6572 (N_6572,N_1077,N_5046);
and U6573 (N_6573,N_1427,N_2227);
xor U6574 (N_6574,N_985,N_3891);
or U6575 (N_6575,N_5506,N_1709);
nor U6576 (N_6576,N_782,N_2413);
or U6577 (N_6577,N_4460,N_2103);
nand U6578 (N_6578,N_5265,N_3845);
nor U6579 (N_6579,N_5898,N_4357);
nand U6580 (N_6580,N_4904,N_1994);
and U6581 (N_6581,N_1525,N_1014);
and U6582 (N_6582,N_1544,N_3670);
nor U6583 (N_6583,N_3046,N_4883);
or U6584 (N_6584,N_230,N_1662);
and U6585 (N_6585,N_5942,N_5360);
or U6586 (N_6586,N_133,N_5925);
nor U6587 (N_6587,N_1606,N_289);
nor U6588 (N_6588,N_3361,N_5078);
xor U6589 (N_6589,N_1543,N_4807);
and U6590 (N_6590,N_2866,N_1661);
or U6591 (N_6591,N_2682,N_806);
nand U6592 (N_6592,N_974,N_3160);
nor U6593 (N_6593,N_648,N_2594);
nand U6594 (N_6594,N_5404,N_4402);
nor U6595 (N_6595,N_1980,N_5987);
nor U6596 (N_6596,N_5565,N_4164);
nor U6597 (N_6597,N_2003,N_74);
and U6598 (N_6598,N_5936,N_2453);
and U6599 (N_6599,N_302,N_4732);
nand U6600 (N_6600,N_3412,N_4553);
or U6601 (N_6601,N_5125,N_5487);
and U6602 (N_6602,N_2077,N_3171);
or U6603 (N_6603,N_4341,N_1916);
nor U6604 (N_6604,N_4612,N_1877);
or U6605 (N_6605,N_2320,N_2089);
nand U6606 (N_6606,N_3363,N_1972);
and U6607 (N_6607,N_5405,N_3185);
nor U6608 (N_6608,N_1036,N_5072);
nand U6609 (N_6609,N_884,N_58);
or U6610 (N_6610,N_1308,N_4626);
and U6611 (N_6611,N_1880,N_509);
nor U6612 (N_6612,N_4843,N_4988);
and U6613 (N_6613,N_4105,N_4617);
or U6614 (N_6614,N_50,N_3146);
nand U6615 (N_6615,N_2840,N_5733);
and U6616 (N_6616,N_5690,N_4215);
nand U6617 (N_6617,N_1819,N_796);
nor U6618 (N_6618,N_2431,N_3250);
and U6619 (N_6619,N_3599,N_4868);
and U6620 (N_6620,N_3910,N_4640);
or U6621 (N_6621,N_1112,N_5917);
nor U6622 (N_6622,N_4218,N_2240);
and U6623 (N_6623,N_579,N_3126);
nor U6624 (N_6624,N_1285,N_2028);
nand U6625 (N_6625,N_4366,N_3801);
nor U6626 (N_6626,N_2256,N_3018);
nor U6627 (N_6627,N_2979,N_5269);
xor U6628 (N_6628,N_3367,N_3918);
or U6629 (N_6629,N_2280,N_5943);
nor U6630 (N_6630,N_3507,N_2655);
nand U6631 (N_6631,N_1373,N_1380);
nand U6632 (N_6632,N_5862,N_4420);
nand U6633 (N_6633,N_4434,N_2113);
or U6634 (N_6634,N_1292,N_4670);
nand U6635 (N_6635,N_4854,N_4701);
nor U6636 (N_6636,N_5213,N_65);
nand U6637 (N_6637,N_4015,N_5511);
nor U6638 (N_6638,N_435,N_1889);
nor U6639 (N_6639,N_3920,N_3195);
or U6640 (N_6640,N_5803,N_964);
or U6641 (N_6641,N_2044,N_4533);
or U6642 (N_6642,N_3896,N_1967);
xnor U6643 (N_6643,N_1755,N_5115);
nand U6644 (N_6644,N_4750,N_254);
xnor U6645 (N_6645,N_303,N_2530);
xnor U6646 (N_6646,N_1751,N_2081);
nor U6647 (N_6647,N_3109,N_3780);
xor U6648 (N_6648,N_5655,N_2181);
and U6649 (N_6649,N_2553,N_3880);
and U6650 (N_6650,N_5924,N_2854);
nand U6651 (N_6651,N_3948,N_177);
or U6652 (N_6652,N_4619,N_5605);
or U6653 (N_6653,N_2074,N_3673);
or U6654 (N_6654,N_4962,N_22);
nor U6655 (N_6655,N_1329,N_1804);
and U6656 (N_6656,N_2150,N_5832);
nand U6657 (N_6657,N_5630,N_2358);
and U6658 (N_6658,N_3386,N_2189);
nor U6659 (N_6659,N_5491,N_4871);
nand U6660 (N_6660,N_1763,N_5002);
or U6661 (N_6661,N_2205,N_1573);
nor U6662 (N_6662,N_4945,N_3419);
xnor U6663 (N_6663,N_5237,N_5503);
nor U6664 (N_6664,N_2601,N_4785);
nand U6665 (N_6665,N_3455,N_4964);
and U6666 (N_6666,N_4139,N_5743);
or U6667 (N_6667,N_4984,N_5795);
or U6668 (N_6668,N_5652,N_4163);
nor U6669 (N_6669,N_1548,N_5498);
nand U6670 (N_6670,N_5016,N_5603);
nand U6671 (N_6671,N_4660,N_4131);
and U6672 (N_6672,N_4672,N_4175);
nor U6673 (N_6673,N_2523,N_5071);
nand U6674 (N_6674,N_73,N_5981);
or U6675 (N_6675,N_3500,N_5330);
nor U6676 (N_6676,N_3857,N_2867);
or U6677 (N_6677,N_1026,N_3949);
and U6678 (N_6678,N_4400,N_1599);
nor U6679 (N_6679,N_1171,N_3403);
and U6680 (N_6680,N_1169,N_3332);
nand U6681 (N_6681,N_4380,N_4138);
nor U6682 (N_6682,N_3652,N_5575);
and U6683 (N_6683,N_3641,N_3544);
nor U6684 (N_6684,N_80,N_4739);
or U6685 (N_6685,N_950,N_2505);
or U6686 (N_6686,N_5376,N_912);
and U6687 (N_6687,N_5300,N_5400);
or U6688 (N_6688,N_392,N_4571);
nor U6689 (N_6689,N_5920,N_3462);
or U6690 (N_6690,N_2470,N_5207);
nand U6691 (N_6691,N_1027,N_1800);
and U6692 (N_6692,N_3236,N_2377);
or U6693 (N_6693,N_2657,N_3728);
or U6694 (N_6694,N_3311,N_1626);
or U6695 (N_6695,N_5377,N_5018);
nand U6696 (N_6696,N_4528,N_2124);
nor U6697 (N_6697,N_4693,N_194);
xor U6698 (N_6698,N_5008,N_577);
or U6699 (N_6699,N_863,N_2533);
nand U6700 (N_6700,N_1782,N_4551);
and U6701 (N_6701,N_922,N_1603);
and U6702 (N_6702,N_115,N_130);
nand U6703 (N_6703,N_3202,N_3268);
nand U6704 (N_6704,N_3042,N_5501);
and U6705 (N_6705,N_2037,N_2885);
xor U6706 (N_6706,N_3514,N_2888);
or U6707 (N_6707,N_1318,N_3312);
and U6708 (N_6708,N_3591,N_1987);
nand U6709 (N_6709,N_5545,N_4472);
nor U6710 (N_6710,N_5421,N_1241);
nand U6711 (N_6711,N_5711,N_4155);
nand U6712 (N_6712,N_5108,N_2773);
xnor U6713 (N_6713,N_2820,N_327);
nand U6714 (N_6714,N_5114,N_4810);
xnor U6715 (N_6715,N_667,N_387);
nand U6716 (N_6716,N_4322,N_4697);
or U6717 (N_6717,N_4698,N_5513);
and U6718 (N_6718,N_3838,N_5416);
or U6719 (N_6719,N_2572,N_4562);
nand U6720 (N_6720,N_5045,N_2573);
xnor U6721 (N_6721,N_362,N_3368);
nor U6722 (N_6722,N_4196,N_379);
and U6723 (N_6723,N_5961,N_206);
xor U6724 (N_6724,N_3615,N_888);
or U6725 (N_6725,N_5740,N_5227);
xor U6726 (N_6726,N_2560,N_4529);
or U6727 (N_6727,N_55,N_3351);
xor U6728 (N_6728,N_3925,N_620);
nor U6729 (N_6729,N_2611,N_858);
nor U6730 (N_6730,N_982,N_2353);
or U6731 (N_6731,N_2494,N_1072);
or U6732 (N_6732,N_2894,N_4176);
and U6733 (N_6733,N_1549,N_2782);
and U6734 (N_6734,N_4655,N_2534);
or U6735 (N_6735,N_82,N_873);
nand U6736 (N_6736,N_2354,N_755);
and U6737 (N_6737,N_646,N_3336);
nor U6738 (N_6738,N_3998,N_3137);
xor U6739 (N_6739,N_823,N_1805);
or U6740 (N_6740,N_3322,N_350);
and U6741 (N_6741,N_104,N_617);
and U6742 (N_6742,N_345,N_5512);
and U6743 (N_6743,N_5459,N_3935);
nor U6744 (N_6744,N_2356,N_2970);
and U6745 (N_6745,N_1743,N_4054);
or U6746 (N_6746,N_2437,N_5451);
xor U6747 (N_6747,N_3490,N_2384);
or U6748 (N_6748,N_4880,N_5593);
and U6749 (N_6749,N_3240,N_4030);
or U6750 (N_6750,N_1646,N_3520);
and U6751 (N_6751,N_3076,N_3253);
xnor U6752 (N_6752,N_512,N_5452);
nor U6753 (N_6753,N_5231,N_2863);
nor U6754 (N_6754,N_366,N_2790);
and U6755 (N_6755,N_5976,N_5680);
or U6756 (N_6756,N_459,N_4245);
and U6757 (N_6757,N_4252,N_5355);
nor U6758 (N_6758,N_5715,N_4021);
nor U6759 (N_6759,N_3672,N_3908);
nand U6760 (N_6760,N_3543,N_1423);
or U6761 (N_6761,N_1485,N_2264);
and U6762 (N_6762,N_3353,N_4715);
and U6763 (N_6763,N_5650,N_3275);
nand U6764 (N_6764,N_4484,N_3260);
and U6765 (N_6765,N_2355,N_4692);
nor U6766 (N_6766,N_3000,N_2570);
and U6767 (N_6767,N_2230,N_2531);
nand U6768 (N_6768,N_4545,N_1866);
nor U6769 (N_6769,N_4809,N_2086);
xnor U6770 (N_6770,N_647,N_4527);
nand U6771 (N_6771,N_3389,N_2703);
nor U6772 (N_6772,N_5879,N_99);
nor U6773 (N_6773,N_2628,N_1126);
nor U6774 (N_6774,N_567,N_2571);
and U6775 (N_6775,N_5858,N_3259);
nand U6776 (N_6776,N_5278,N_639);
nand U6777 (N_6777,N_3729,N_4486);
nand U6778 (N_6778,N_1477,N_691);
xor U6779 (N_6779,N_4067,N_3205);
or U6780 (N_6780,N_321,N_3528);
nand U6781 (N_6781,N_5767,N_2612);
or U6782 (N_6782,N_3357,N_4020);
nor U6783 (N_6783,N_3469,N_5670);
nand U6784 (N_6784,N_4930,N_2924);
nor U6785 (N_6785,N_5027,N_3538);
nand U6786 (N_6786,N_1097,N_2748);
and U6787 (N_6787,N_1420,N_5006);
or U6788 (N_6788,N_5433,N_1872);
and U6789 (N_6789,N_268,N_1227);
xor U6790 (N_6790,N_5752,N_4923);
and U6791 (N_6791,N_1005,N_297);
nand U6792 (N_6792,N_3806,N_4833);
and U6793 (N_6793,N_2739,N_977);
nand U6794 (N_6794,N_3633,N_4748);
and U6795 (N_6795,N_5149,N_2800);
nor U6796 (N_6796,N_4001,N_5837);
xor U6797 (N_6797,N_5639,N_1153);
nor U6798 (N_6798,N_2791,N_1676);
xnor U6799 (N_6799,N_473,N_578);
xnor U6800 (N_6800,N_4694,N_2669);
nand U6801 (N_6801,N_4536,N_844);
and U6802 (N_6802,N_5426,N_4445);
nor U6803 (N_6803,N_2488,N_4323);
and U6804 (N_6804,N_5768,N_1486);
and U6805 (N_6805,N_1937,N_5657);
nor U6806 (N_6806,N_4303,N_4399);
xor U6807 (N_6807,N_561,N_5960);
xnor U6808 (N_6808,N_2245,N_255);
nand U6809 (N_6809,N_1780,N_892);
nor U6810 (N_6810,N_5375,N_4659);
nand U6811 (N_6811,N_3339,N_1834);
nor U6812 (N_6812,N_5306,N_3515);
or U6813 (N_6813,N_2972,N_5540);
nand U6814 (N_6814,N_5441,N_2580);
and U6815 (N_6815,N_3704,N_2434);
xnor U6816 (N_6816,N_1886,N_5363);
and U6817 (N_6817,N_1418,N_3049);
and U6818 (N_6818,N_1791,N_3545);
or U6819 (N_6819,N_833,N_5986);
or U6820 (N_6820,N_2848,N_3956);
nand U6821 (N_6821,N_4699,N_3075);
nand U6822 (N_6822,N_966,N_2935);
or U6823 (N_6823,N_3083,N_499);
nand U6824 (N_6824,N_1503,N_292);
nand U6825 (N_6825,N_2799,N_5281);
and U6826 (N_6826,N_3617,N_2852);
or U6827 (N_6827,N_1975,N_5461);
or U6828 (N_6828,N_5966,N_2609);
or U6829 (N_6829,N_4857,N_2734);
nor U6830 (N_6830,N_4903,N_1554);
and U6831 (N_6831,N_5746,N_1047);
nand U6832 (N_6832,N_2042,N_5823);
and U6833 (N_6833,N_5408,N_1713);
or U6834 (N_6834,N_4673,N_5555);
or U6835 (N_6835,N_4494,N_1297);
and U6836 (N_6836,N_5754,N_3431);
xnor U6837 (N_6837,N_535,N_747);
nor U6838 (N_6838,N_182,N_1513);
and U6839 (N_6839,N_5900,N_2582);
nand U6840 (N_6840,N_751,N_1294);
xor U6841 (N_6841,N_1637,N_3820);
and U6842 (N_6842,N_5275,N_1766);
or U6843 (N_6843,N_5607,N_1447);
nand U6844 (N_6844,N_914,N_90);
or U6845 (N_6845,N_4097,N_859);
nor U6846 (N_6846,N_116,N_5722);
nor U6847 (N_6847,N_2544,N_3238);
and U6848 (N_6848,N_4633,N_658);
or U6849 (N_6849,N_1508,N_1345);
xor U6850 (N_6850,N_3724,N_5747);
nand U6851 (N_6851,N_4972,N_5205);
xnor U6852 (N_6852,N_788,N_5399);
or U6853 (N_6853,N_3439,N_2091);
or U6854 (N_6854,N_3833,N_3176);
nor U6855 (N_6855,N_5395,N_1315);
or U6856 (N_6856,N_4056,N_5049);
nor U6857 (N_6857,N_3777,N_5720);
xor U6858 (N_6858,N_3219,N_1250);
and U6859 (N_6859,N_4028,N_4534);
nand U6860 (N_6860,N_5398,N_4049);
nand U6861 (N_6861,N_4401,N_2126);
nand U6862 (N_6862,N_2452,N_5203);
nor U6863 (N_6863,N_876,N_172);
or U6864 (N_6864,N_3929,N_707);
xnor U6865 (N_6865,N_4152,N_28);
nand U6866 (N_6866,N_937,N_1004);
or U6867 (N_6867,N_3610,N_126);
nand U6868 (N_6868,N_3213,N_1213);
or U6869 (N_6869,N_1677,N_1828);
nand U6870 (N_6870,N_3369,N_1453);
and U6871 (N_6871,N_5894,N_3849);
nand U6872 (N_6872,N_4574,N_3382);
nand U6873 (N_6873,N_2386,N_2869);
and U6874 (N_6874,N_5980,N_1964);
and U6875 (N_6875,N_2916,N_5530);
or U6876 (N_6876,N_3773,N_3628);
nor U6877 (N_6877,N_2031,N_2005);
nand U6878 (N_6878,N_822,N_2259);
and U6879 (N_6879,N_1159,N_1741);
xor U6880 (N_6880,N_153,N_4985);
or U6881 (N_6881,N_1807,N_5780);
nor U6882 (N_6882,N_1664,N_5508);
and U6883 (N_6883,N_2337,N_4425);
nand U6884 (N_6884,N_4772,N_1489);
or U6885 (N_6885,N_4771,N_1978);
nand U6886 (N_6886,N_3457,N_4866);
or U6887 (N_6887,N_2499,N_3040);
nand U6888 (N_6888,N_2010,N_1467);
nand U6889 (N_6889,N_2497,N_4795);
or U6890 (N_6890,N_1468,N_3060);
nor U6891 (N_6891,N_2507,N_4233);
or U6892 (N_6892,N_1089,N_5882);
or U6893 (N_6893,N_1963,N_1092);
nand U6894 (N_6894,N_5058,N_5396);
nand U6895 (N_6895,N_5903,N_5885);
and U6896 (N_6896,N_2368,N_3921);
nand U6897 (N_6897,N_463,N_1616);
xor U6898 (N_6898,N_2969,N_2015);
and U6899 (N_6899,N_365,N_200);
nor U6900 (N_6900,N_4708,N_5791);
nand U6901 (N_6901,N_951,N_598);
nand U6902 (N_6902,N_5946,N_4754);
nand U6903 (N_6903,N_253,N_4840);
or U6904 (N_6904,N_2836,N_1663);
nand U6905 (N_6905,N_1530,N_4970);
nand U6906 (N_6906,N_320,N_5028);
nand U6907 (N_6907,N_1956,N_4024);
xnor U6908 (N_6908,N_1175,N_5723);
xor U6909 (N_6909,N_920,N_66);
xnor U6910 (N_6910,N_1473,N_5055);
nand U6911 (N_6911,N_5849,N_483);
nand U6912 (N_6912,N_5794,N_188);
nor U6913 (N_6913,N_4585,N_868);
nor U6914 (N_6914,N_3743,N_3848);
or U6915 (N_6915,N_2075,N_2610);
and U6916 (N_6916,N_3846,N_1870);
or U6917 (N_6917,N_5505,N_5820);
or U6918 (N_6918,N_2861,N_336);
nor U6919 (N_6919,N_3614,N_3594);
nor U6920 (N_6920,N_2614,N_1180);
nand U6921 (N_6921,N_4184,N_1177);
nand U6922 (N_6922,N_4337,N_2511);
nor U6923 (N_6923,N_3557,N_5385);
nor U6924 (N_6924,N_2613,N_1927);
nor U6925 (N_6925,N_5323,N_5600);
or U6926 (N_6926,N_2590,N_1968);
xnor U6927 (N_6927,N_1162,N_980);
or U6928 (N_6928,N_491,N_3464);
and U6929 (N_6929,N_1142,N_3053);
and U6930 (N_6930,N_5040,N_3752);
nand U6931 (N_6931,N_4927,N_1609);
and U6932 (N_6932,N_4343,N_1799);
and U6933 (N_6933,N_2457,N_1472);
xor U6934 (N_6934,N_2443,N_3869);
nand U6935 (N_6935,N_5331,N_220);
or U6936 (N_6936,N_4505,N_1428);
nor U6937 (N_6937,N_3217,N_897);
nor U6938 (N_6938,N_5063,N_5069);
or U6939 (N_6939,N_1306,N_4281);
xor U6940 (N_6940,N_1865,N_3155);
or U6941 (N_6941,N_3818,N_2870);
nand U6942 (N_6942,N_789,N_3559);
nand U6943 (N_6943,N_4848,N_467);
or U6944 (N_6944,N_4466,N_5440);
or U6945 (N_6945,N_2185,N_3593);
nor U6946 (N_6946,N_511,N_2252);
and U6947 (N_6947,N_2139,N_1643);
nand U6948 (N_6948,N_1382,N_4700);
or U6949 (N_6949,N_5136,N_2363);
nor U6950 (N_6950,N_3009,N_3308);
and U6951 (N_6951,N_1374,N_4711);
or U6952 (N_6952,N_3218,N_5088);
or U6953 (N_6953,N_4803,N_3050);
nand U6954 (N_6954,N_2514,N_481);
xnor U6955 (N_6955,N_1343,N_2306);
nand U6956 (N_6956,N_4581,N_1988);
nor U6957 (N_6957,N_5877,N_5100);
xnor U6958 (N_6958,N_1605,N_4455);
nor U6959 (N_6959,N_2990,N_2508);
nor U6960 (N_6960,N_4350,N_621);
and U6961 (N_6961,N_3745,N_1029);
or U6962 (N_6962,N_4584,N_441);
and U6963 (N_6963,N_2651,N_2827);
nor U6964 (N_6964,N_2892,N_4278);
and U6965 (N_6965,N_1784,N_785);
or U6966 (N_6966,N_2893,N_3306);
or U6967 (N_6967,N_3629,N_2908);
nor U6968 (N_6968,N_2933,N_2811);
or U6969 (N_6969,N_1317,N_4968);
or U6970 (N_6970,N_2627,N_2294);
nor U6971 (N_6971,N_2426,N_3950);
and U6972 (N_6972,N_885,N_1864);
nor U6973 (N_6973,N_1470,N_221);
nand U6974 (N_6974,N_3737,N_314);
nand U6975 (N_6975,N_3823,N_700);
and U6976 (N_6976,N_611,N_4995);
nand U6977 (N_6977,N_5321,N_779);
nand U6978 (N_6978,N_983,N_1737);
nor U6979 (N_6979,N_5014,N_2041);
xnor U6980 (N_6980,N_963,N_4799);
nor U6981 (N_6981,N_1654,N_1270);
nand U6982 (N_6982,N_2001,N_5786);
or U6983 (N_6983,N_1938,N_2475);
nor U6984 (N_6984,N_2640,N_2936);
or U6985 (N_6985,N_5978,N_2344);
xnor U6986 (N_6986,N_1614,N_1776);
xnor U6987 (N_6987,N_355,N_4387);
or U6988 (N_6988,N_1902,N_5620);
nand U6989 (N_6989,N_1565,N_538);
nor U6990 (N_6990,N_2552,N_4424);
or U6991 (N_6991,N_2653,N_4549);
nand U6992 (N_6992,N_0,N_698);
nor U6993 (N_6993,N_1913,N_310);
and U6994 (N_6994,N_5738,N_5251);
and U6995 (N_6995,N_1185,N_1096);
and U6996 (N_6996,N_347,N_1890);
or U6997 (N_6997,N_3839,N_5834);
xor U6998 (N_6998,N_1222,N_765);
nor U6999 (N_6999,N_1361,N_3307);
nand U7000 (N_7000,N_1557,N_3501);
nor U7001 (N_7001,N_2056,N_2302);
or U7002 (N_7002,N_5296,N_2938);
and U7003 (N_7003,N_3632,N_168);
or U7004 (N_7004,N_5244,N_4862);
nor U7005 (N_7005,N_4921,N_2159);
or U7006 (N_7006,N_4286,N_3043);
and U7007 (N_7007,N_3084,N_2400);
and U7008 (N_7008,N_3048,N_1669);
or U7009 (N_7009,N_2818,N_4119);
nor U7010 (N_7010,N_4432,N_5345);
xor U7011 (N_7011,N_318,N_3537);
xor U7012 (N_7012,N_3297,N_1492);
xor U7013 (N_7013,N_2107,N_32);
nand U7014 (N_7014,N_1961,N_3829);
or U7015 (N_7015,N_1949,N_3979);
or U7016 (N_7016,N_4573,N_5167);
and U7017 (N_7017,N_3148,N_1408);
nor U7018 (N_7018,N_2804,N_3191);
or U7019 (N_7019,N_4222,N_399);
nand U7020 (N_7020,N_4274,N_946);
and U7021 (N_7021,N_2998,N_2725);
nor U7022 (N_7022,N_1216,N_708);
and U7023 (N_7023,N_3815,N_5959);
nand U7024 (N_7024,N_2487,N_1971);
nor U7025 (N_7025,N_5812,N_840);
or U7026 (N_7026,N_2705,N_3696);
or U7027 (N_7027,N_883,N_2154);
or U7028 (N_7028,N_3578,N_3036);
and U7029 (N_7029,N_2549,N_5951);
and U7030 (N_7030,N_308,N_4328);
nor U7031 (N_7031,N_1397,N_5775);
nor U7032 (N_7032,N_79,N_2518);
nand U7033 (N_7033,N_4600,N_2766);
or U7034 (N_7034,N_3087,N_1445);
and U7035 (N_7035,N_5934,N_1523);
or U7036 (N_7036,N_4065,N_1948);
nor U7037 (N_7037,N_3740,N_5429);
nand U7038 (N_7038,N_7,N_1693);
and U7039 (N_7039,N_3634,N_2723);
or U7040 (N_7040,N_4763,N_1900);
or U7041 (N_7041,N_1371,N_5159);
or U7042 (N_7042,N_3422,N_2502);
nor U7043 (N_7043,N_454,N_5996);
nor U7044 (N_7044,N_3793,N_353);
and U7045 (N_7045,N_3150,N_3055);
nor U7046 (N_7046,N_1772,N_3035);
and U7047 (N_7047,N_3553,N_1986);
or U7048 (N_7048,N_818,N_1009);
or U7049 (N_7049,N_2749,N_240);
nand U7050 (N_7050,N_5787,N_1083);
xor U7051 (N_7051,N_3573,N_4507);
nor U7052 (N_7052,N_777,N_2027);
or U7053 (N_7053,N_5864,N_242);
and U7054 (N_7054,N_2939,N_761);
and U7055 (N_7055,N_1762,N_2535);
nand U7056 (N_7056,N_1229,N_3890);
nor U7057 (N_7057,N_1186,N_3086);
or U7058 (N_7058,N_3969,N_4778);
nor U7059 (N_7059,N_1501,N_5466);
or U7060 (N_7060,N_743,N_3911);
xor U7061 (N_7061,N_3161,N_703);
xor U7062 (N_7062,N_2024,N_2373);
and U7063 (N_7063,N_4461,N_5592);
xnor U7064 (N_7064,N_5389,N_5876);
nand U7065 (N_7065,N_502,N_3093);
xnor U7066 (N_7066,N_397,N_3679);
and U7067 (N_7067,N_5562,N_3899);
nand U7068 (N_7068,N_4410,N_1534);
xnor U7069 (N_7069,N_3390,N_5310);
nand U7070 (N_7070,N_4707,N_3529);
and U7071 (N_7071,N_2350,N_3517);
nand U7072 (N_7072,N_3744,N_4452);
xor U7073 (N_7073,N_443,N_3502);
nor U7074 (N_7074,N_3158,N_5896);
or U7075 (N_7075,N_110,N_1650);
and U7076 (N_7076,N_3551,N_3939);
nand U7077 (N_7077,N_1111,N_2810);
and U7078 (N_7078,N_4289,N_5646);
or U7079 (N_7079,N_2441,N_4892);
xor U7080 (N_7080,N_210,N_760);
nand U7081 (N_7081,N_492,N_2152);
xnor U7082 (N_7082,N_1054,N_165);
or U7083 (N_7083,N_3512,N_1517);
or U7084 (N_7084,N_769,N_4508);
and U7085 (N_7085,N_1493,N_5526);
or U7086 (N_7086,N_249,N_5687);
nand U7087 (N_7087,N_5609,N_5349);
xnor U7088 (N_7088,N_4465,N_4493);
xnor U7089 (N_7089,N_996,N_1892);
and U7090 (N_7090,N_1935,N_1652);
and U7091 (N_7091,N_4437,N_1254);
and U7092 (N_7092,N_2807,N_2706);
xor U7093 (N_7093,N_2839,N_836);
nand U7094 (N_7094,N_1161,N_5490);
and U7095 (N_7095,N_4397,N_1055);
nor U7096 (N_7096,N_654,N_961);
nand U7097 (N_7097,N_710,N_5542);
and U7098 (N_7098,N_5623,N_3105);
and U7099 (N_7099,N_3138,N_1752);
or U7100 (N_7100,N_1267,N_299);
or U7101 (N_7101,N_3198,N_1699);
or U7102 (N_7102,N_5431,N_1757);
and U7103 (N_7103,N_1076,N_3461);
and U7104 (N_7104,N_2455,N_3922);
or U7105 (N_7105,N_3296,N_791);
or U7106 (N_7106,N_4777,N_251);
or U7107 (N_7107,N_3354,N_670);
xnor U7108 (N_7108,N_3565,N_3897);
xor U7109 (N_7109,N_5683,N_1895);
or U7110 (N_7110,N_3860,N_4755);
nor U7111 (N_7111,N_938,N_4417);
and U7112 (N_7112,N_1120,N_3002);
nor U7113 (N_7113,N_4873,N_3071);
nand U7114 (N_7114,N_5113,N_3278);
nand U7115 (N_7115,N_2621,N_2521);
nor U7116 (N_7116,N_2219,N_3711);
nor U7117 (N_7117,N_1379,N_1115);
and U7118 (N_7118,N_4375,N_1506);
xnor U7119 (N_7119,N_1923,N_3812);
or U7120 (N_7120,N_5822,N_5469);
xor U7121 (N_7121,N_2815,N_2206);
and U7122 (N_7122,N_2630,N_2802);
nand U7123 (N_7123,N_3426,N_5521);
nand U7124 (N_7124,N_1367,N_5784);
nand U7125 (N_7125,N_2274,N_3153);
xnor U7126 (N_7126,N_3947,N_386);
nand U7127 (N_7127,N_4068,N_1989);
nor U7128 (N_7128,N_5707,N_993);
nand U7129 (N_7129,N_4195,N_52);
or U7130 (N_7130,N_3059,N_2825);
nor U7131 (N_7131,N_998,N_5866);
or U7132 (N_7132,N_5424,N_4459);
nand U7133 (N_7133,N_4550,N_199);
nand U7134 (N_7134,N_4894,N_3643);
xor U7135 (N_7135,N_311,N_5922);
and U7136 (N_7136,N_1158,N_138);
nor U7137 (N_7137,N_4246,N_4214);
nor U7138 (N_7138,N_3058,N_1826);
and U7139 (N_7139,N_4099,N_4531);
nor U7140 (N_7140,N_3766,N_5854);
xnor U7141 (N_7141,N_2849,N_2254);
nor U7142 (N_7142,N_2890,N_1611);
nand U7143 (N_7143,N_3639,N_5284);
nand U7144 (N_7144,N_5938,N_5899);
nor U7145 (N_7145,N_3125,N_464);
nand U7146 (N_7146,N_4045,N_5904);
nand U7147 (N_7147,N_4726,N_53);
and U7148 (N_7148,N_5907,N_4118);
and U7149 (N_7149,N_5897,N_2584);
and U7150 (N_7150,N_413,N_5544);
nor U7151 (N_7151,N_5247,N_4136);
and U7152 (N_7152,N_465,N_3924);
and U7153 (N_7153,N_4247,N_262);
and U7154 (N_7154,N_5805,N_4265);
nand U7155 (N_7155,N_5079,N_4669);
or U7156 (N_7156,N_319,N_1440);
and U7157 (N_7157,N_636,N_4666);
or U7158 (N_7158,N_3063,N_1001);
nand U7159 (N_7159,N_5473,N_5949);
and U7160 (N_7160,N_4203,N_223);
nor U7161 (N_7161,N_1885,N_2562);
or U7162 (N_7162,N_4041,N_5548);
and U7163 (N_7163,N_4566,N_706);
and U7164 (N_7164,N_1324,N_735);
and U7165 (N_7165,N_1779,N_3725);
nor U7166 (N_7166,N_2199,N_312);
and U7167 (N_7167,N_2273,N_2821);
or U7168 (N_7168,N_5279,N_5572);
or U7169 (N_7169,N_1720,N_1690);
and U7170 (N_7170,N_4557,N_5235);
nor U7171 (N_7171,N_2341,N_2445);
nand U7172 (N_7172,N_3415,N_4869);
or U7173 (N_7173,N_2960,N_1129);
or U7174 (N_7174,N_505,N_4378);
nor U7175 (N_7175,N_1479,N_1021);
xor U7176 (N_7176,N_1249,N_3980);
and U7177 (N_7177,N_1277,N_2013);
or U7178 (N_7178,N_5830,N_2565);
nand U7179 (N_7179,N_3589,N_4865);
and U7180 (N_7180,N_1952,N_3345);
nor U7181 (N_7181,N_4012,N_5742);
or U7182 (N_7182,N_3798,N_3554);
or U7183 (N_7183,N_257,N_1604);
and U7184 (N_7184,N_3826,N_3468);
or U7185 (N_7185,N_5188,N_5438);
or U7186 (N_7186,N_4946,N_5216);
nor U7187 (N_7187,N_4500,N_420);
or U7188 (N_7188,N_404,N_5679);
nor U7189 (N_7189,N_2575,N_1514);
and U7190 (N_7190,N_5048,N_4834);
or U7191 (N_7191,N_3836,N_4300);
and U7192 (N_7192,N_3370,N_1362);
or U7193 (N_7193,N_2687,N_4942);
and U7194 (N_7194,N_488,N_3967);
nor U7195 (N_7195,N_4275,N_3271);
and U7196 (N_7196,N_4183,N_744);
and U7197 (N_7197,N_5529,N_388);
and U7198 (N_7198,N_5169,N_1332);
and U7199 (N_7199,N_1732,N_3755);
and U7200 (N_7200,N_3165,N_2536);
nand U7201 (N_7201,N_1483,N_770);
or U7202 (N_7202,N_1314,N_2277);
nor U7203 (N_7203,N_306,N_3903);
nor U7204 (N_7204,N_3592,N_3623);
xor U7205 (N_7205,N_187,N_1814);
nor U7206 (N_7206,N_3983,N_5895);
and U7207 (N_7207,N_2450,N_3765);
nand U7208 (N_7208,N_1251,N_3844);
nand U7209 (N_7209,N_4663,N_5285);
nor U7210 (N_7210,N_5316,N_717);
nor U7211 (N_7211,N_5068,N_375);
nor U7212 (N_7212,N_3156,N_5170);
nor U7213 (N_7213,N_5052,N_4588);
or U7214 (N_7214,N_4158,N_1898);
and U7215 (N_7215,N_3721,N_969);
nand U7216 (N_7216,N_4808,N_5736);
and U7217 (N_7217,N_559,N_622);
nor U7218 (N_7218,N_29,N_4824);
or U7219 (N_7219,N_3224,N_1469);
and U7220 (N_7220,N_768,N_1926);
nor U7221 (N_7221,N_2328,N_5788);
xnor U7222 (N_7222,N_2137,N_4540);
and U7223 (N_7223,N_5272,N_5665);
or U7224 (N_7224,N_5686,N_4632);
nand U7225 (N_7225,N_1260,N_1416);
or U7226 (N_7226,N_33,N_1003);
nand U7227 (N_7227,N_3843,N_36);
or U7228 (N_7228,N_5432,N_4724);
and U7229 (N_7229,N_4262,N_3095);
xor U7230 (N_7230,N_5706,N_5085);
nor U7231 (N_7231,N_5643,N_2269);
nor U7232 (N_7232,N_2393,N_4449);
and U7233 (N_7233,N_1067,N_2293);
and U7234 (N_7234,N_5467,N_2545);
nor U7235 (N_7235,N_3847,N_4780);
nor U7236 (N_7236,N_1712,N_1698);
or U7237 (N_7237,N_5037,N_5881);
nor U7238 (N_7238,N_2226,N_1521);
or U7239 (N_7239,N_5940,N_5558);
nor U7240 (N_7240,N_3451,N_406);
and U7241 (N_7241,N_1039,N_2995);
nor U7242 (N_7242,N_4153,N_2096);
or U7243 (N_7243,N_773,N_2989);
or U7244 (N_7244,N_1552,N_298);
nand U7245 (N_7245,N_3665,N_2676);
nor U7246 (N_7246,N_3376,N_4114);
xor U7247 (N_7247,N_1533,N_3791);
xor U7248 (N_7248,N_5635,N_5410);
or U7249 (N_7249,N_3435,N_2408);
nand U7250 (N_7250,N_5869,N_4037);
nand U7251 (N_7251,N_4990,N_5838);
nor U7252 (N_7252,N_4832,N_3540);
or U7253 (N_7253,N_5312,N_2522);
and U7254 (N_7254,N_911,N_5122);
nand U7255 (N_7255,N_1205,N_5796);
nor U7256 (N_7256,N_3056,N_4762);
xnor U7257 (N_7257,N_5927,N_3885);
nand U7258 (N_7258,N_4876,N_1759);
xor U7259 (N_7259,N_3768,N_3600);
xnor U7260 (N_7260,N_3794,N_1058);
nor U7261 (N_7261,N_1509,N_162);
nor U7262 (N_7262,N_832,N_2700);
or U7263 (N_7263,N_2902,N_1792);
nand U7264 (N_7264,N_2817,N_2999);
and U7265 (N_7265,N_4379,N_3934);
xor U7266 (N_7266,N_1808,N_3073);
or U7267 (N_7267,N_1157,N_5152);
or U7268 (N_7268,N_2814,N_5552);
nand U7269 (N_7269,N_5271,N_2490);
nand U7270 (N_7270,N_1556,N_2415);
nor U7271 (N_7271,N_503,N_2182);
nand U7272 (N_7272,N_4462,N_4874);
xnor U7273 (N_7273,N_1444,N_5232);
or U7274 (N_7274,N_2992,N_2728);
nor U7275 (N_7275,N_3423,N_4730);
nand U7276 (N_7276,N_2675,N_1426);
and U7277 (N_7277,N_1874,N_1671);
nor U7278 (N_7278,N_5004,N_1011);
and U7279 (N_7279,N_921,N_3346);
nand U7280 (N_7280,N_845,N_2726);
and U7281 (N_7281,N_2004,N_3004);
nand U7282 (N_7282,N_3552,N_5119);
or U7283 (N_7283,N_4084,N_86);
or U7284 (N_7284,N_750,N_2966);
nor U7285 (N_7285,N_1983,N_5067);
xnor U7286 (N_7286,N_100,N_47);
nand U7287 (N_7287,N_4975,N_4648);
or U7288 (N_7288,N_1290,N_2737);
or U7289 (N_7289,N_1025,N_3726);
nor U7290 (N_7290,N_5277,N_2325);
xnor U7291 (N_7291,N_337,N_4344);
xor U7292 (N_7292,N_2049,N_2065);
and U7293 (N_7293,N_2048,N_19);
nor U7294 (N_7294,N_4535,N_3409);
nor U7295 (N_7295,N_872,N_4881);
nand U7296 (N_7296,N_2961,N_1770);
nand U7297 (N_7297,N_5525,N_2047);
and U7298 (N_7298,N_731,N_2261);
and U7299 (N_7299,N_2129,N_2978);
nand U7300 (N_7300,N_96,N_3066);
or U7301 (N_7301,N_5827,N_4925);
and U7302 (N_7302,N_516,N_1350);
and U7303 (N_7303,N_734,N_599);
and U7304 (N_7304,N_4204,N_3877);
or U7305 (N_7305,N_1284,N_1128);
or U7306 (N_7306,N_1031,N_1134);
or U7307 (N_7307,N_1037,N_948);
nor U7308 (N_7308,N_5674,N_2993);
nand U7309 (N_7309,N_3814,N_4595);
nand U7310 (N_7310,N_2012,N_5610);
nor U7311 (N_7311,N_1079,N_3338);
nor U7312 (N_7312,N_2436,N_4369);
xor U7313 (N_7313,N_585,N_954);
xor U7314 (N_7314,N_817,N_1947);
nand U7315 (N_7315,N_3182,N_2225);
nor U7316 (N_7316,N_893,N_3915);
or U7317 (N_7317,N_85,N_5873);
nand U7318 (N_7318,N_3006,N_4490);
nor U7319 (N_7319,N_3209,N_5648);
or U7320 (N_7320,N_3488,N_1409);
and U7321 (N_7321,N_3981,N_5759);
xnor U7322 (N_7322,N_5848,N_4443);
and U7323 (N_7323,N_5968,N_5591);
nor U7324 (N_7324,N_2504,N_3990);
xor U7325 (N_7325,N_3486,N_4066);
or U7326 (N_7326,N_5859,N_1644);
xnor U7327 (N_7327,N_5611,N_3662);
nor U7328 (N_7328,N_722,N_1333);
and U7329 (N_7329,N_4481,N_3769);
nor U7330 (N_7330,N_2064,N_1592);
nand U7331 (N_7331,N_4716,N_2054);
nor U7332 (N_7332,N_4317,N_5226);
xor U7333 (N_7333,N_5257,N_3051);
nand U7334 (N_7334,N_3964,N_1248);
nand U7335 (N_7335,N_3889,N_4912);
or U7336 (N_7336,N_1675,N_3027);
xnor U7337 (N_7337,N_1041,N_2974);
nor U7338 (N_7338,N_2365,N_3247);
xnor U7339 (N_7339,N_5036,N_1433);
nor U7340 (N_7340,N_5618,N_1617);
or U7341 (N_7341,N_4134,N_4983);
and U7342 (N_7342,N_461,N_3454);
nand U7343 (N_7343,N_2805,N_3108);
xnor U7344 (N_7344,N_1413,N_1922);
or U7345 (N_7345,N_5047,N_333);
nor U7346 (N_7346,N_727,N_4639);
nand U7347 (N_7347,N_2067,N_2838);
and U7348 (N_7348,N_2311,N_295);
and U7349 (N_7349,N_1302,N_4889);
xor U7350 (N_7350,N_403,N_4948);
nand U7351 (N_7351,N_482,N_21);
and U7352 (N_7352,N_5826,N_3973);
or U7353 (N_7353,N_736,N_5034);
and U7354 (N_7354,N_5083,N_4667);
nor U7355 (N_7355,N_2694,N_896);
nand U7356 (N_7356,N_4594,N_4237);
nor U7357 (N_7357,N_1833,N_4025);
nand U7358 (N_7358,N_907,N_5080);
xor U7359 (N_7359,N_2603,N_4078);
nor U7360 (N_7360,N_5470,N_184);
or U7361 (N_7361,N_4302,N_3487);
or U7362 (N_7362,N_3094,N_3220);
nand U7363 (N_7363,N_3693,N_4888);
nand U7364 (N_7364,N_641,N_4360);
nand U7365 (N_7365,N_3622,N_1946);
or U7366 (N_7366,N_1487,N_4788);
nand U7367 (N_7367,N_2751,N_5133);
nand U7368 (N_7368,N_4760,N_5971);
and U7369 (N_7369,N_396,N_5007);
and U7370 (N_7370,N_4266,N_2942);
nor U7371 (N_7371,N_3590,N_3347);
nand U7372 (N_7372,N_4254,N_2263);
or U7373 (N_7373,N_3596,N_455);
or U7374 (N_7374,N_864,N_5177);
nor U7375 (N_7375,N_3865,N_5534);
xnor U7376 (N_7376,N_4181,N_4310);
or U7377 (N_7377,N_2503,N_536);
and U7378 (N_7378,N_500,N_5800);
and U7379 (N_7379,N_637,N_3810);
or U7380 (N_7380,N_3115,N_4144);
nor U7381 (N_7381,N_2058,N_3210);
or U7382 (N_7382,N_423,N_4468);
nor U7383 (N_7383,N_2595,N_136);
nor U7384 (N_7384,N_5835,N_1316);
or U7385 (N_7385,N_5578,N_2432);
nand U7386 (N_7386,N_3638,N_2299);
nand U7387 (N_7387,N_5673,N_5218);
nor U7388 (N_7388,N_3241,N_5988);
or U7389 (N_7389,N_714,N_1845);
or U7390 (N_7390,N_1588,N_1160);
nand U7391 (N_7391,N_4475,N_3266);
or U7392 (N_7392,N_2029,N_5494);
and U7393 (N_7393,N_5499,N_4499);
and U7394 (N_7394,N_2021,N_3961);
nor U7395 (N_7395,N_587,N_2994);
nor U7396 (N_7396,N_1275,N_610);
nor U7397 (N_7397,N_3406,N_4312);
or U7398 (N_7398,N_4664,N_3291);
nor U7399 (N_7399,N_2050,N_4069);
xor U7400 (N_7400,N_5150,N_2952);
and U7401 (N_7401,N_3646,N_3682);
or U7402 (N_7402,N_2427,N_4451);
nand U7403 (N_7403,N_3471,N_5789);
nand U7404 (N_7404,N_1991,N_5013);
and U7405 (N_7405,N_3440,N_4351);
nor U7406 (N_7406,N_3356,N_1237);
and U7407 (N_7407,N_4706,N_3294);
nor U7408 (N_7408,N_1840,N_3136);
xor U7409 (N_7409,N_2949,N_4367);
or U7410 (N_7410,N_3072,N_4811);
and U7411 (N_7411,N_4875,N_414);
and U7412 (N_7412,N_5336,N_5700);
and U7413 (N_7413,N_227,N_2787);
nor U7414 (N_7414,N_5293,N_4661);
or U7415 (N_7415,N_1094,N_3506);
nor U7416 (N_7416,N_827,N_159);
nor U7417 (N_7417,N_4538,N_5148);
xor U7418 (N_7418,N_1006,N_5641);
or U7419 (N_7419,N_1727,N_2374);
or U7420 (N_7420,N_2312,N_1750);
and U7421 (N_7421,N_278,N_629);
and U7422 (N_7422,N_5550,N_239);
or U7423 (N_7423,N_5845,N_4924);
nor U7424 (N_7424,N_1596,N_2190);
and U7425 (N_7425,N_1579,N_2865);
nand U7426 (N_7426,N_5164,N_4690);
and U7427 (N_7427,N_2586,N_5201);
nand U7428 (N_7428,N_1057,N_867);
and U7429 (N_7429,N_147,N_1985);
xor U7430 (N_7430,N_5504,N_3384);
nand U7431 (N_7431,N_5024,N_1363);
nand U7432 (N_7432,N_635,N_4217);
or U7433 (N_7433,N_3644,N_2528);
nand U7434 (N_7434,N_1165,N_4146);
and U7435 (N_7435,N_2822,N_2448);
or U7436 (N_7436,N_4235,N_3932);
or U7437 (N_7437,N_322,N_1695);
or U7438 (N_7438,N_4013,N_1091);
nor U7439 (N_7439,N_5220,N_4298);
nand U7440 (N_7440,N_4238,N_5341);
nor U7441 (N_7441,N_4684,N_2428);
nand U7442 (N_7442,N_4313,N_1069);
or U7443 (N_7443,N_891,N_3988);
nor U7444 (N_7444,N_5939,N_3476);
nand U7445 (N_7445,N_3695,N_957);
nand U7446 (N_7446,N_2864,N_719);
or U7447 (N_7447,N_1760,N_3207);
and U7448 (N_7448,N_4646,N_2855);
and U7449 (N_7449,N_4409,N_3365);
nor U7450 (N_7450,N_225,N_398);
nand U7451 (N_7451,N_4603,N_1002);
nor U7452 (N_7452,N_1625,N_4886);
and U7453 (N_7453,N_4406,N_4111);
and U7454 (N_7454,N_5209,N_2342);
and U7455 (N_7455,N_2629,N_1849);
nand U7456 (N_7456,N_5401,N_3975);
nand U7457 (N_7457,N_1977,N_5070);
nor U7458 (N_7458,N_4556,N_2529);
or U7459 (N_7459,N_198,N_4829);
or U7460 (N_7460,N_3568,N_5761);
or U7461 (N_7461,N_3524,N_5870);
and U7462 (N_7462,N_1829,N_1303);
or U7463 (N_7463,N_1349,N_5262);
xor U7464 (N_7464,N_628,N_4261);
or U7465 (N_7465,N_4849,N_5549);
nor U7466 (N_7466,N_2093,N_2006);
xor U7467 (N_7467,N_2806,N_3624);
and U7468 (N_7468,N_3395,N_3797);
and U7469 (N_7469,N_3280,N_3433);
and U7470 (N_7470,N_1370,N_5270);
nor U7471 (N_7471,N_3941,N_933);
nand U7472 (N_7472,N_5912,N_3556);
and U7473 (N_7473,N_2382,N_3647);
and U7474 (N_7474,N_4583,N_3764);
and U7475 (N_7475,N_2673,N_4709);
nand U7476 (N_7476,N_4362,N_1125);
nand U7477 (N_7477,N_3909,N_2680);
nor U7478 (N_7478,N_645,N_3359);
or U7479 (N_7479,N_3564,N_5824);
nor U7480 (N_7480,N_5249,N_293);
and U7481 (N_7481,N_201,N_5668);
or U7482 (N_7482,N_5886,N_4851);
xor U7483 (N_7483,N_5198,N_5241);
nand U7484 (N_7484,N_1141,N_5339);
nor U7485 (N_7485,N_2020,N_5692);
nor U7486 (N_7486,N_1786,N_4170);
or U7487 (N_7487,N_1348,N_4180);
or U7488 (N_7488,N_3653,N_5109);
or U7489 (N_7489,N_792,N_5678);
or U7490 (N_7490,N_5731,N_5792);
and U7491 (N_7491,N_4610,N_4609);
and U7492 (N_7492,N_1612,N_4630);
nor U7493 (N_7493,N_39,N_4213);
and U7494 (N_7494,N_427,N_1130);
and U7495 (N_7495,N_469,N_4756);
and U7496 (N_7496,N_1334,N_5691);
nor U7497 (N_7497,N_3366,N_1106);
nand U7498 (N_7498,N_4161,N_2598);
or U7499 (N_7499,N_5640,N_1225);
or U7500 (N_7500,N_2232,N_2172);
nor U7501 (N_7501,N_4088,N_4284);
nand U7502 (N_7502,N_5327,N_5520);
and U7503 (N_7503,N_5802,N_2469);
and U7504 (N_7504,N_5729,N_3685);
and U7505 (N_7505,N_2577,N_31);
and U7506 (N_7506,N_5734,N_5825);
and U7507 (N_7507,N_997,N_13);
xor U7508 (N_7508,N_2388,N_1569);
nand U7509 (N_7509,N_1731,N_4002);
nand U7510 (N_7510,N_5766,N_5274);
or U7511 (N_7511,N_5583,N_821);
nor U7512 (N_7512,N_5419,N_3178);
nor U7513 (N_7513,N_1296,N_3159);
and U7514 (N_7514,N_1555,N_466);
xnor U7515 (N_7515,N_2955,N_1639);
nand U7516 (N_7516,N_3170,N_5533);
nor U7517 (N_7517,N_988,N_970);
nor U7518 (N_7518,N_2759,N_2155);
nand U7519 (N_7519,N_1313,N_504);
nand U7520 (N_7520,N_30,N_3868);
and U7521 (N_7521,N_918,N_5409);
or U7522 (N_7522,N_357,N_4906);
nor U7523 (N_7523,N_2593,N_5041);
or U7524 (N_7524,N_4333,N_2592);
or U7525 (N_7525,N_3841,N_973);
nor U7526 (N_7526,N_3039,N_393);
nand U7527 (N_7527,N_5351,N_5948);
and U7528 (N_7528,N_3070,N_2985);
nor U7529 (N_7529,N_4421,N_4260);
nand U7530 (N_7530,N_3478,N_3572);
or U7531 (N_7531,N_3141,N_1033);
nand U7532 (N_7532,N_2688,N_452);
nor U7533 (N_7533,N_3456,N_2121);
and U7534 (N_7534,N_42,N_3563);
or U7535 (N_7535,N_2229,N_3834);
nor U7536 (N_7536,N_5865,N_5111);
nor U7537 (N_7537,N_3341,N_4023);
xnor U7538 (N_7538,N_1073,N_3770);
and U7539 (N_7539,N_1993,N_2922);
nand U7540 (N_7540,N_3940,N_5160);
xor U7541 (N_7541,N_171,N_2322);
and U7542 (N_7542,N_4806,N_2214);
or U7543 (N_7543,N_3532,N_417);
nor U7544 (N_7544,N_5025,N_1576);
or U7545 (N_7545,N_2197,N_3803);
xnor U7546 (N_7546,N_442,N_4160);
xor U7547 (N_7547,N_1931,N_4723);
and U7548 (N_7548,N_1235,N_2767);
and U7549 (N_7549,N_4413,N_5741);
nand U7550 (N_7550,N_4062,N_5098);
and U7551 (N_7551,N_4931,N_4587);
nor U7552 (N_7552,N_3946,N_3438);
and U7553 (N_7553,N_2889,N_5704);
nand U7554 (N_7554,N_2092,N_1906);
xnor U7555 (N_7555,N_2828,N_4977);
and U7556 (N_7556,N_2837,N_5225);
or U7557 (N_7557,N_681,N_5763);
nor U7558 (N_7558,N_701,N_4342);
nor U7559 (N_7559,N_1138,N_591);
xnor U7560 (N_7560,N_4248,N_5590);
and U7561 (N_7561,N_3875,N_739);
xnor U7562 (N_7562,N_5573,N_2605);
and U7563 (N_7563,N_1787,N_3174);
or U7564 (N_7564,N_759,N_3421);
and U7565 (N_7565,N_4821,N_2366);
xor U7566 (N_7566,N_5957,N_5653);
or U7567 (N_7567,N_721,N_4853);
nand U7568 (N_7568,N_5324,N_2464);
or U7569 (N_7569,N_1697,N_4496);
or U7570 (N_7570,N_2039,N_815);
or U7571 (N_7571,N_4456,N_2071);
xnor U7572 (N_7572,N_2776,N_1442);
nor U7573 (N_7573,N_2795,N_3223);
and U7574 (N_7574,N_5745,N_3637);
nor U7575 (N_7575,N_2747,N_4447);
and U7576 (N_7576,N_3101,N_1568);
and U7577 (N_7577,N_5243,N_1894);
nor U7578 (N_7578,N_2875,N_3525);
nor U7579 (N_7579,N_5210,N_4159);
or U7580 (N_7580,N_3180,N_3586);
nor U7581 (N_7581,N_936,N_2439);
and U7582 (N_7582,N_4100,N_3140);
xor U7583 (N_7583,N_4251,N_514);
nand U7584 (N_7584,N_4564,N_5174);
and U7585 (N_7585,N_4129,N_5730);
or U7586 (N_7586,N_3531,N_5872);
or U7587 (N_7587,N_5147,N_4996);
xor U7588 (N_7588,N_425,N_787);
xor U7589 (N_7589,N_2250,N_2847);
nor U7590 (N_7590,N_2175,N_4905);
nand U7591 (N_7591,N_2880,N_3447);
nand U7592 (N_7592,N_4007,N_685);
nor U7593 (N_7593,N_5146,N_1030);
nand U7594 (N_7594,N_3966,N_1683);
or U7595 (N_7595,N_2527,N_5776);
nor U7596 (N_7596,N_61,N_4491);
nand U7597 (N_7597,N_1795,N_1201);
nand U7598 (N_7598,N_1878,N_1266);
nor U7599 (N_7599,N_4828,N_2618);
nor U7600 (N_7600,N_1914,N_4695);
and U7601 (N_7601,N_742,N_498);
and U7602 (N_7602,N_1360,N_2638);
and U7603 (N_7603,N_1434,N_959);
and U7604 (N_7604,N_4582,N_1196);
nand U7605 (N_7605,N_4501,N_4844);
nand U7606 (N_7606,N_3997,N_1674);
nor U7607 (N_7607,N_4509,N_25);
xor U7608 (N_7608,N_2953,N_3837);
xnor U7609 (N_7609,N_1958,N_3977);
and U7610 (N_7610,N_816,N_2101);
and U7611 (N_7611,N_5595,N_4752);
nand U7612 (N_7612,N_2194,N_416);
nand U7613 (N_7613,N_2496,N_5893);
and U7614 (N_7614,N_2275,N_4127);
nor U7615 (N_7615,N_688,N_3580);
xnor U7616 (N_7616,N_582,N_2647);
nand U7617 (N_7617,N_352,N_3763);
nor U7618 (N_7618,N_3866,N_2367);
nand U7619 (N_7619,N_1749,N_272);
nand U7620 (N_7620,N_904,N_3113);
and U7621 (N_7621,N_181,N_752);
nor U7622 (N_7622,N_4044,N_2596);
or U7623 (N_7623,N_2208,N_2788);
and U7624 (N_7624,N_4415,N_3052);
xnor U7625 (N_7625,N_2128,N_3930);
or U7626 (N_7626,N_3807,N_5479);
xor U7627 (N_7627,N_1295,N_5402);
nor U7628 (N_7628,N_4149,N_3315);
or U7629 (N_7629,N_371,N_2242);
nand U7630 (N_7630,N_478,N_359);
or U7631 (N_7631,N_3458,N_1189);
or U7632 (N_7632,N_851,N_5000);
nand U7633 (N_7633,N_2597,N_4242);
nand U7634 (N_7634,N_1516,N_5181);
or U7635 (N_7635,N_24,N_5694);
nor U7636 (N_7636,N_4745,N_987);
nand U7637 (N_7637,N_1562,N_564);
nand U7638 (N_7638,N_2371,N_2744);
nand U7639 (N_7639,N_2724,N_3149);
nand U7640 (N_7640,N_1346,N_1392);
or U7641 (N_7641,N_4518,N_2729);
nand U7642 (N_7642,N_3561,N_3410);
and U7643 (N_7643,N_4568,N_2210);
nor U7644 (N_7644,N_3124,N_1062);
nor U7645 (N_7645,N_4790,N_604);
nand U7646 (N_7646,N_3135,N_2973);
xnor U7647 (N_7647,N_5567,N_1622);
nand U7648 (N_7648,N_716,N_4495);
and U7649 (N_7649,N_5364,N_3411);
nand U7650 (N_7650,N_4729,N_1567);
or U7651 (N_7651,N_3398,N_3761);
xor U7652 (N_7652,N_660,N_5471);
nor U7653 (N_7653,N_5568,N_4282);
nand U7654 (N_7654,N_3273,N_1139);
nand U7655 (N_7655,N_2568,N_5744);
or U7656 (N_7656,N_5955,N_4781);
or U7657 (N_7657,N_1940,N_542);
or U7658 (N_7658,N_875,N_4137);
nor U7659 (N_7659,N_3694,N_2084);
xnor U7660 (N_7660,N_521,N_4019);
or U7661 (N_7661,N_4083,N_1119);
nor U7662 (N_7662,N_1010,N_2906);
and U7663 (N_7663,N_1739,N_2167);
and U7664 (N_7664,N_5952,N_1621);
and U7665 (N_7665,N_4773,N_1630);
and U7666 (N_7666,N_5612,N_5250);
and U7667 (N_7667,N_3655,N_1385);
nand U7668 (N_7668,N_1022,N_693);
nand U7669 (N_7669,N_5842,N_4979);
nand U7670 (N_7670,N_5191,N_4992);
or U7671 (N_7671,N_5012,N_4963);
or U7672 (N_7672,N_830,N_5412);
nand U7673 (N_7673,N_857,N_3116);
and U7674 (N_7674,N_5428,N_916);
nor U7675 (N_7675,N_2650,N_3079);
nand U7676 (N_7676,N_4264,N_2449);
and U7677 (N_7677,N_949,N_784);
nand U7678 (N_7678,N_3129,N_5140);
or U7679 (N_7679,N_4798,N_5366);
or U7680 (N_7680,N_1597,N_878);
and U7681 (N_7681,N_1247,N_601);
and U7682 (N_7682,N_4332,N_819);
nor U7683 (N_7683,N_1801,N_1301);
and U7684 (N_7684,N_3031,N_1546);
xnor U7685 (N_7685,N_501,N_1623);
nand U7686 (N_7686,N_680,N_5307);
nand U7687 (N_7687,N_5065,N_3319);
nor U7688 (N_7688,N_2561,N_2391);
or U7689 (N_7689,N_4860,N_1309);
nand U7690 (N_7690,N_3320,N_2789);
nand U7691 (N_7691,N_4687,N_3555);
or U7692 (N_7692,N_2033,N_4658);
nand U7693 (N_7693,N_4976,N_4616);
nor U7694 (N_7694,N_4802,N_5774);
nor U7695 (N_7695,N_4381,N_2034);
nand U7696 (N_7696,N_3703,N_624);
xnor U7697 (N_7697,N_339,N_5963);
xor U7698 (N_7698,N_1681,N_1330);
nor U7699 (N_7699,N_1500,N_2120);
or U7700 (N_7700,N_903,N_4190);
and U7701 (N_7701,N_3360,N_4269);
xnor U7702 (N_7702,N_3074,N_1905);
nor U7703 (N_7703,N_4742,N_304);
nor U7704 (N_7704,N_5342,N_2244);
or U7705 (N_7705,N_2479,N_4042);
or U7706 (N_7706,N_4951,N_1903);
and U7707 (N_7707,N_5732,N_4053);
or U7708 (N_7708,N_3030,N_5887);
and U7709 (N_7709,N_2394,N_2904);
nand U7710 (N_7710,N_1818,N_4953);
xnor U7711 (N_7711,N_1384,N_2243);
and U7712 (N_7712,N_3299,N_5783);
nand U7713 (N_7713,N_250,N_3222);
and U7714 (N_7714,N_2632,N_5857);
or U7715 (N_7715,N_2335,N_3254);
or U7716 (N_7716,N_5001,N_3090);
or U7717 (N_7717,N_939,N_3082);
and U7718 (N_7718,N_4241,N_3751);
and U7719 (N_7719,N_4914,N_3167);
nand U7720 (N_7720,N_4547,N_2832);
and U7721 (N_7721,N_88,N_401);
nor U7722 (N_7722,N_4225,N_3945);
or U7723 (N_7723,N_1326,N_2209);
nand U7724 (N_7724,N_1341,N_395);
nand U7725 (N_7725,N_798,N_2699);
nand U7726 (N_7726,N_4572,N_5828);
xor U7727 (N_7727,N_5371,N_4112);
and U7728 (N_7728,N_3825,N_877);
nor U7729 (N_7729,N_1852,N_1694);
and U7730 (N_7730,N_3325,N_3656);
xor U7731 (N_7731,N_3912,N_3951);
nand U7732 (N_7732,N_5162,N_4205);
and U7733 (N_7733,N_3472,N_5962);
or U7734 (N_7734,N_3189,N_1280);
nor U7735 (N_7735,N_1288,N_5212);
nand U7736 (N_7736,N_5030,N_3);
and U7737 (N_7737,N_5809,N_4599);
and U7738 (N_7738,N_5702,N_2424);
nand U7739 (N_7739,N_5138,N_608);
nor U7740 (N_7740,N_2845,N_2665);
xor U7741 (N_7741,N_5861,N_4961);
nor U7742 (N_7742,N_3943,N_1781);
or U7743 (N_7743,N_4971,N_2340);
or U7744 (N_7744,N_3119,N_5);
and U7745 (N_7745,N_894,N_4722);
and U7746 (N_7746,N_2022,N_4219);
nor U7747 (N_7747,N_4120,N_4842);
nor U7748 (N_7748,N_2402,N_1429);
xor U7749 (N_7749,N_4643,N_129);
nor U7750 (N_7750,N_1670,N_2620);
nand U7751 (N_7751,N_211,N_5356);
nor U7752 (N_7752,N_4800,N_192);
and U7753 (N_7753,N_2937,N_236);
nand U7754 (N_7754,N_5846,N_1178);
and U7755 (N_7755,N_4143,N_4256);
nand U7756 (N_7756,N_2716,N_1105);
and U7757 (N_7757,N_2122,N_3541);
or U7758 (N_7758,N_2289,N_486);
and U7759 (N_7759,N_5202,N_62);
nand U7760 (N_7760,N_3381,N_3343);
and U7761 (N_7761,N_5362,N_870);
xor U7762 (N_7762,N_1207,N_1200);
nor U7763 (N_7763,N_3068,N_3927);
or U7764 (N_7764,N_2462,N_4973);
or U7765 (N_7765,N_4761,N_1137);
nor U7766 (N_7766,N_329,N_2304);
nand U7767 (N_7767,N_3496,N_5453);
nand U7768 (N_7768,N_241,N_2693);
and U7769 (N_7769,N_3309,N_3371);
and U7770 (N_7770,N_4436,N_2066);
and U7771 (N_7771,N_2588,N_2684);
and U7772 (N_7772,N_1257,N_1710);
nor U7773 (N_7773,N_3792,N_246);
and U7774 (N_7774,N_5075,N_1400);
nand U7775 (N_7775,N_753,N_2168);
and U7776 (N_7776,N_1074,N_3738);
and U7777 (N_7777,N_3701,N_3197);
nor U7778 (N_7778,N_1145,N_484);
or U7779 (N_7779,N_2526,N_2677);
nor U7780 (N_7780,N_3878,N_718);
and U7781 (N_7781,N_886,N_931);
and U7782 (N_7782,N_3867,N_3602);
nor U7783 (N_7783,N_1337,N_4974);
nand U7784 (N_7784,N_5117,N_3497);
and U7785 (N_7785,N_5086,N_4525);
nand U7786 (N_7786,N_5753,N_5204);
and U7787 (N_7787,N_3008,N_5531);
nand U7788 (N_7788,N_2357,N_955);
nor U7789 (N_7789,N_1687,N_2060);
and U7790 (N_7790,N_2895,N_4314);
nor U7791 (N_7791,N_1061,N_4431);
nor U7792 (N_7792,N_2385,N_3504);
nand U7793 (N_7793,N_1881,N_142);
nand U7794 (N_7794,N_1268,N_2540);
nor U7795 (N_7795,N_5891,N_2881);
nand U7796 (N_7796,N_1539,N_1502);
nor U7797 (N_7797,N_5658,N_3962);
or U7798 (N_7798,N_2143,N_529);
nor U7799 (N_7799,N_5492,N_5260);
or U7800 (N_7800,N_5192,N_652);
or U7801 (N_7801,N_2631,N_3111);
nor U7802 (N_7802,N_2369,N_555);
xor U7803 (N_7803,N_2430,N_5042);
or U7804 (N_7804,N_1018,N_990);
or U7805 (N_7805,N_2251,N_3734);
nor U7806 (N_7806,N_2606,N_2696);
or U7807 (N_7807,N_4627,N_2919);
nor U7808 (N_7808,N_5104,N_408);
and U7809 (N_7809,N_4657,N_5984);
nor U7810 (N_7810,N_2798,N_4288);
nand U7811 (N_7811,N_360,N_3650);
and U7812 (N_7812,N_4597,N_145);
nand U7813 (N_7813,N_1387,N_1645);
nand U7814 (N_7814,N_5038,N_4124);
or U7815 (N_7815,N_5909,N_1575);
nand U7816 (N_7816,N_5821,N_5175);
nor U7817 (N_7817,N_2135,N_3474);
and U7818 (N_7818,N_2658,N_2962);
nor U7819 (N_7819,N_1998,N_3418);
nor U7820 (N_7820,N_4009,N_3505);
and U7821 (N_7821,N_4346,N_3034);
and U7822 (N_7822,N_5524,N_1718);
nor U7823 (N_7823,N_1059,N_1708);
nand U7824 (N_7824,N_5368,N_445);
and U7825 (N_7825,N_5184,N_2253);
and U7826 (N_7826,N_4404,N_37);
or U7827 (N_7827,N_38,N_2069);
nand U7828 (N_7828,N_1692,N_3383);
nand U7829 (N_7829,N_2176,N_2876);
xor U7830 (N_7830,N_1212,N_87);
nand U7831 (N_7831,N_4920,N_1131);
and U7832 (N_7832,N_3481,N_4135);
and U7833 (N_7833,N_4649,N_2543);
and U7834 (N_7834,N_3904,N_49);
nand U7835 (N_7835,N_354,N_4820);
nand U7836 (N_7836,N_3898,N_1439);
nor U7837 (N_7837,N_5121,N_1421);
and U7838 (N_7838,N_4651,N_547);
nor U7839 (N_7839,N_5636,N_135);
nor U7840 (N_7840,N_1053,N_523);
nor U7841 (N_7841,N_5696,N_4331);
xnor U7842 (N_7842,N_5143,N_1868);
nand U7843 (N_7843,N_4374,N_476);
nand U7844 (N_7844,N_1619,N_2109);
xnor U7845 (N_7845,N_3678,N_3821);
or U7846 (N_7846,N_730,N_5322);
nor U7847 (N_7847,N_2070,N_4825);
or U7848 (N_7848,N_1143,N_678);
nand U7849 (N_7849,N_5632,N_614);
xnor U7850 (N_7850,N_5228,N_3131);
nand U7851 (N_7851,N_4489,N_3231);
and U7852 (N_7852,N_5553,N_4743);
or U7853 (N_7853,N_3226,N_1875);
nand U7854 (N_7854,N_1537,N_1929);
and U7855 (N_7855,N_5793,N_5346);
or U7856 (N_7856,N_2282,N_5569);
nand U7857 (N_7857,N_1744,N_1282);
xnor U7858 (N_7858,N_382,N_35);
or U7859 (N_7859,N_1133,N_5628);
nand U7860 (N_7860,N_6,N_3978);
and U7861 (N_7861,N_3011,N_2591);
xnor U7862 (N_7862,N_4216,N_301);
nand U7863 (N_7863,N_2316,N_1920);
nor U7864 (N_7864,N_3516,N_4885);
and U7865 (N_7865,N_3666,N_4384);
or U7866 (N_7866,N_1151,N_4125);
nand U7867 (N_7867,N_2846,N_3938);
nor U7868 (N_7868,N_1594,N_1891);
or U7869 (N_7869,N_4321,N_3019);
and U7870 (N_7870,N_346,N_3100);
and U7871 (N_7871,N_5712,N_1634);
and U7872 (N_7872,N_2713,N_1893);
nor U7873 (N_7873,N_5455,N_549);
and U7874 (N_7874,N_1924,N_4299);
and U7875 (N_7875,N_4736,N_2279);
or U7876 (N_7876,N_3645,N_5454);
nor U7877 (N_7877,N_4319,N_2954);
and U7878 (N_7878,N_3830,N_573);
or U7879 (N_7879,N_43,N_4006);
nand U7880 (N_7880,N_1230,N_5818);
nor U7881 (N_7881,N_5992,N_63);
or U7882 (N_7882,N_1331,N_2546);
nor U7883 (N_7883,N_3619,N_593);
or U7884 (N_7884,N_1319,N_5695);
xnor U7885 (N_7885,N_2491,N_2087);
nor U7886 (N_7886,N_4867,N_3753);
or U7887 (N_7887,N_1867,N_2698);
and U7888 (N_7888,N_376,N_3314);
and U7889 (N_7889,N_2292,N_3588);
and U7890 (N_7890,N_5698,N_5645);
nand U7891 (N_7891,N_3575,N_3562);
or U7892 (N_7892,N_1383,N_3463);
or U7893 (N_7893,N_4365,N_668);
or U7894 (N_7894,N_3186,N_2147);
and U7895 (N_7895,N_2515,N_2082);
nor U7896 (N_7896,N_4596,N_3900);
and U7897 (N_7897,N_84,N_2416);
nand U7898 (N_7898,N_2390,N_4937);
or U7899 (N_7899,N_4345,N_2266);
or U7900 (N_7900,N_2644,N_3870);
and U7901 (N_7901,N_4483,N_4916);
nor U7902 (N_7902,N_5128,N_4101);
nand U7903 (N_7903,N_3400,N_696);
or U7904 (N_7904,N_1325,N_4786);
or U7905 (N_7905,N_342,N_5662);
nand U7906 (N_7906,N_2334,N_1934);
or U7907 (N_7907,N_3021,N_3003);
nor U7908 (N_7908,N_3530,N_3404);
or U7909 (N_7909,N_4032,N_2899);
or U7910 (N_7910,N_2314,N_5581);
xor U7911 (N_7911,N_1197,N_5519);
nor U7912 (N_7912,N_5560,N_5965);
and U7913 (N_7913,N_4668,N_3518);
nor U7914 (N_7914,N_2399,N_673);
xor U7915 (N_7915,N_5163,N_1871);
and U7916 (N_7916,N_3681,N_1154);
and U7917 (N_7917,N_266,N_1960);
nand U7918 (N_7918,N_5617,N_4098);
and U7919 (N_7919,N_5799,N_687);
nor U7920 (N_7920,N_4082,N_843);
or U7921 (N_7921,N_1104,N_627);
or U7922 (N_7922,N_2932,N_527);
or U7923 (N_7923,N_2548,N_5884);
nand U7924 (N_7924,N_3335,N_3269);
or U7925 (N_7925,N_124,N_531);
nand U7926 (N_7926,N_612,N_4898);
nor U7927 (N_7927,N_140,N_5179);
nor U7928 (N_7928,N_3723,N_2421);
nand U7929 (N_7929,N_282,N_229);
nor U7930 (N_7930,N_4090,N_4909);
nor U7931 (N_7931,N_887,N_92);
xor U7932 (N_7932,N_3242,N_3892);
nand U7933 (N_7933,N_2537,N_5510);
or U7934 (N_7934,N_287,N_2500);
nand U7935 (N_7935,N_3778,N_3037);
nand U7936 (N_7936,N_1336,N_5031);
or U7937 (N_7937,N_5254,N_2662);
or U7938 (N_7938,N_4804,N_315);
nor U7939 (N_7939,N_5814,N_4835);
nand U7940 (N_7940,N_1085,N_2664);
nor U7941 (N_7941,N_1049,N_54);
nand U7942 (N_7942,N_4234,N_3188);
xor U7943 (N_7943,N_4685,N_213);
nor U7944 (N_7944,N_3475,N_3960);
or U7945 (N_7945,N_4368,N_3121);
nand U7946 (N_7946,N_4171,N_5689);
and U7947 (N_7947,N_2401,N_4864);
nand U7948 (N_7948,N_1773,N_1764);
nor U7949 (N_7949,N_1327,N_2123);
nor U7950 (N_7950,N_193,N_4936);
nand U7951 (N_7951,N_4815,N_4339);
nor U7952 (N_7952,N_605,N_5200);
xnor U7953 (N_7953,N_4911,N_5333);
nor U7954 (N_7954,N_2754,N_3625);
and U7955 (N_7955,N_4036,N_248);
xor U7956 (N_7956,N_3229,N_2652);
and U7957 (N_7957,N_1745,N_852);
nand U7958 (N_7958,N_2032,N_5554);
and U7959 (N_7959,N_2731,N_4315);
nand U7960 (N_7960,N_824,N_40);
nor U7961 (N_7961,N_1724,N_3748);
nand U7962 (N_7962,N_3190,N_1879);
and U7963 (N_7963,N_4197,N_1446);
xor U7964 (N_7964,N_4939,N_5305);
nor U7965 (N_7965,N_3722,N_615);
xor U7966 (N_7966,N_1278,N_1082);
nand U7967 (N_7967,N_1,N_429);
and U7968 (N_7968,N_4228,N_1340);
and U7969 (N_7969,N_757,N_3408);
nand U7970 (N_7970,N_335,N_3560);
nor U7971 (N_7971,N_4047,N_4192);
nor U7972 (N_7972,N_3535,N_1909);
nor U7973 (N_7973,N_4884,N_5343);
nand U7974 (N_7974,N_3790,N_5043);
nand U7975 (N_7975,N_4081,N_2438);
nor U7976 (N_7976,N_1323,N_3995);
nand U7977 (N_7977,N_1118,N_4947);
nand U7978 (N_7978,N_5945,N_2695);
nand U7979 (N_7979,N_4656,N_2146);
or U7980 (N_7980,N_839,N_3424);
nand U7981 (N_7981,N_3982,N_4253);
xor U7982 (N_7982,N_2153,N_989);
or U7983 (N_7983,N_5843,N_4878);
nand U7984 (N_7984,N_4682,N_1455);
and U7985 (N_7985,N_330,N_4579);
nand U7986 (N_7986,N_5717,N_4759);
or U7987 (N_7987,N_123,N_2112);
and U7988 (N_7988,N_5975,N_2615);
and U7989 (N_7989,N_5437,N_267);
or U7990 (N_7990,N_5584,N_1824);
nor U7991 (N_7991,N_5435,N_4987);
nand U7992 (N_7992,N_4064,N_3779);
or U7993 (N_7993,N_1344,N_1846);
nand U7994 (N_7994,N_4521,N_3788);
nand U7995 (N_7995,N_889,N_5422);
xnor U7996 (N_7996,N_3965,N_3427);
and U7997 (N_7997,N_1038,N_113);
xnor U7998 (N_7998,N_161,N_5482);
and U7999 (N_7999,N_4244,N_316);
and U8000 (N_8000,N_3168,N_3566);
nor U8001 (N_8001,N_5208,N_3080);
or U8002 (N_8002,N_3225,N_2480);
or U8003 (N_8003,N_4683,N_1425);
or U8004 (N_8004,N_166,N_5019);
and U8005 (N_8005,N_1020,N_2878);
xor U8006 (N_8006,N_928,N_1815);
nor U8007 (N_8007,N_5462,N_128);
or U8008 (N_8008,N_3631,N_3181);
and U8009 (N_8009,N_3216,N_2378);
nand U8010 (N_8010,N_114,N_5311);
xor U8011 (N_8011,N_5020,N_4589);
and U8012 (N_8012,N_477,N_149);
and U8013 (N_8013,N_1375,N_4774);
and U8014 (N_8014,N_4010,N_4812);
or U8015 (N_8015,N_45,N_2986);
and U8016 (N_8016,N_4712,N_4926);
or U8017 (N_8017,N_3120,N_216);
and U8018 (N_8018,N_5495,N_5003);
or U8019 (N_8019,N_5566,N_5215);
nor U8020 (N_8020,N_1719,N_5594);
nand U8021 (N_8021,N_853,N_960);
nor U8022 (N_8022,N_2149,N_592);
nor U8023 (N_8023,N_4676,N_942);
or U8024 (N_8024,N_1932,N_4611);
nand U8025 (N_8025,N_3276,N_3986);
nand U8026 (N_8026,N_5867,N_2482);
or U8027 (N_8027,N_2141,N_4476);
and U8028 (N_8028,N_332,N_1704);
or U8029 (N_8029,N_5094,N_1869);
and U8030 (N_8030,N_2258,N_3776);
or U8031 (N_8031,N_4607,N_4405);
and U8032 (N_8032,N_1179,N_196);
or U8033 (N_8033,N_2100,N_3549);
or U8034 (N_8034,N_78,N_1921);
xor U8035 (N_8035,N_1378,N_4725);
or U8036 (N_8036,N_3064,N_2410);
nor U8037 (N_8037,N_4255,N_943);
nor U8038 (N_8038,N_865,N_5654);
and U8039 (N_8039,N_197,N_650);
and U8040 (N_8040,N_3324,N_3203);
and U8041 (N_8041,N_4358,N_2764);
nor U8042 (N_8042,N_1102,N_2988);
or U8043 (N_8043,N_4593,N_5320);
nor U8044 (N_8044,N_4128,N_5134);
nor U8045 (N_8045,N_1310,N_1217);
or U8046 (N_8046,N_5379,N_5777);
and U8047 (N_8047,N_5084,N_1726);
nor U8048 (N_8048,N_2532,N_5171);
nand U8049 (N_8049,N_155,N_409);
and U8050 (N_8050,N_3289,N_369);
nand U8051 (N_8051,N_3445,N_4826);
or U8052 (N_8052,N_967,N_2247);
nand U8053 (N_8053,N_2285,N_5403);
and U8054 (N_8054,N_2934,N_799);
xnor U8055 (N_8055,N_2581,N_5559);
and U8056 (N_8056,N_68,N_5958);
or U8057 (N_8057,N_5602,N_1827);
or U8058 (N_8058,N_3654,N_325);
nor U8059 (N_8059,N_2574,N_2857);
xnor U8060 (N_8060,N_4537,N_4210);
nor U8061 (N_8061,N_4092,N_2079);
nand U8062 (N_8062,N_676,N_1854);
nor U8063 (N_8063,N_1716,N_5764);
and U8064 (N_8064,N_3785,N_4768);
nor U8065 (N_8065,N_1992,N_1242);
nor U8066 (N_8066,N_2241,N_663);
or U8067 (N_8067,N_4850,N_3061);
nor U8068 (N_8068,N_5596,N_5234);
xor U8069 (N_8069,N_5944,N_3396);
and U8070 (N_8070,N_1402,N_2873);
and U8071 (N_8071,N_1044,N_3352);
or U8072 (N_8072,N_495,N_3211);
nor U8073 (N_8073,N_811,N_4232);
or U8074 (N_8074,N_5990,N_4110);
nor U8075 (N_8075,N_148,N_4457);
and U8076 (N_8076,N_4897,N_4511);
or U8077 (N_8077,N_5297,N_5908);
nor U8078 (N_8078,N_119,N_4497);
and U8079 (N_8079,N_2897,N_2483);
nand U8080 (N_8080,N_1655,N_2088);
nand U8081 (N_8081,N_5407,N_3316);
nor U8082 (N_8082,N_603,N_3758);
or U8083 (N_8083,N_402,N_5688);
and U8084 (N_8084,N_1436,N_296);
xnor U8085 (N_8085,N_2489,N_828);
nand U8086 (N_8086,N_4997,N_3416);
xnor U8087 (N_8087,N_83,N_3452);
nand U8088 (N_8088,N_762,N_67);
xor U8089 (N_8089,N_4958,N_3953);
and U8090 (N_8090,N_1942,N_850);
xor U8091 (N_8091,N_4733,N_5762);
nor U8092 (N_8092,N_23,N_4714);
or U8093 (N_8093,N_763,N_1414);
and U8094 (N_8094,N_1711,N_48);
and U8095 (N_8095,N_4398,N_2330);
or U8096 (N_8096,N_2192,N_4613);
or U8097 (N_8097,N_5060,N_2983);
and U8098 (N_8098,N_2585,N_3264);
or U8099 (N_8099,N_411,N_541);
nand U8100 (N_8100,N_4057,N_1368);
and U8101 (N_8101,N_4470,N_4735);
and U8102 (N_8102,N_5582,N_1435);
or U8103 (N_8103,N_5139,N_20);
nand U8104 (N_8104,N_3710,N_4407);
nand U8105 (N_8105,N_4575,N_2346);
nor U8106 (N_8106,N_2262,N_5102);
and U8107 (N_8107,N_3974,N_1598);
nor U8108 (N_8108,N_3663,N_2486);
nor U8109 (N_8109,N_537,N_238);
nor U8110 (N_8110,N_3713,N_5137);
xnor U8111 (N_8111,N_1070,N_952);
nor U8112 (N_8112,N_4391,N_5677);
or U8113 (N_8113,N_1150,N_1672);
and U8114 (N_8114,N_554,N_713);
nand U8115 (N_8115,N_3510,N_745);
nor U8116 (N_8116,N_2260,N_683);
and U8117 (N_8117,N_1918,N_3233);
nor U8118 (N_8118,N_2683,N_1761);
nor U8119 (N_8119,N_2917,N_3690);
nor U8120 (N_8120,N_1271,N_214);
and U8121 (N_8121,N_879,N_632);
and U8122 (N_8122,N_2472,N_846);
nor U8123 (N_8123,N_1936,N_1876);
xor U8124 (N_8124,N_5313,N_1527);
or U8125 (N_8125,N_5029,N_3200);
nand U8126 (N_8126,N_4688,N_4473);
and U8127 (N_8127,N_1793,N_2830);
and U8128 (N_8128,N_1457,N_3819);
and U8129 (N_8129,N_1456,N_2144);
or U8130 (N_8130,N_1193,N_5411);
nand U8131 (N_8131,N_1415,N_1858);
and U8132 (N_8132,N_5576,N_2287);
nand U8133 (N_8133,N_4450,N_2017);
nand U8134 (N_8134,N_5445,N_2035);
or U8135 (N_8135,N_5427,N_3467);
and U8136 (N_8136,N_3828,N_2466);
nor U8137 (N_8137,N_5131,N_5979);
nand U8138 (N_8138,N_2444,N_280);
nand U8139 (N_8139,N_2715,N_4270);
nand U8140 (N_8140,N_5599,N_5703);
and U8141 (N_8141,N_3835,N_2474);
nand U8142 (N_8142,N_1602,N_3127);
and U8143 (N_8143,N_3757,N_4408);
nor U8144 (N_8144,N_1649,N_4173);
and U8145 (N_8145,N_1831,N_5097);
or U8146 (N_8146,N_2977,N_1839);
nor U8147 (N_8147,N_5033,N_4969);
or U8148 (N_8148,N_2918,N_4145);
and U8149 (N_8149,N_2211,N_4154);
or U8150 (N_8150,N_733,N_3831);
or U8151 (N_8151,N_932,N_2711);
and U8152 (N_8152,N_2709,N_1943);
and U8153 (N_8153,N_5103,N_3045);
nor U8154 (N_8154,N_1258,N_3123);
or U8155 (N_8155,N_2984,N_4622);
or U8156 (N_8156,N_1656,N_1364);
or U8157 (N_8157,N_1841,N_2967);
nor U8158 (N_8158,N_4295,N_1570);
or U8159 (N_8159,N_1899,N_3144);
and U8160 (N_8160,N_2007,N_5579);
and U8161 (N_8161,N_4236,N_2345);
or U8162 (N_8162,N_1127,N_4093);
xnor U8163 (N_8163,N_895,N_5782);
nand U8164 (N_8164,N_674,N_364);
and U8165 (N_8165,N_5693,N_4186);
and U8166 (N_8166,N_3984,N_5178);
nand U8167 (N_8167,N_1347,N_4113);
or U8168 (N_8168,N_1144,N_3775);
nor U8169 (N_8169,N_2237,N_5261);
xor U8170 (N_8170,N_5413,N_2098);
xor U8171 (N_8171,N_4189,N_1226);
or U8172 (N_8172,N_5197,N_5325);
and U8173 (N_8173,N_4570,N_4749);
xnor U8174 (N_8174,N_5066,N_2051);
or U8175 (N_8175,N_41,N_5021);
and U8176 (N_8176,N_1386,N_3895);
or U8177 (N_8177,N_944,N_3527);
nor U8178 (N_8178,N_5172,N_471);
nand U8179 (N_8179,N_1276,N_127);
xnor U8180 (N_8180,N_758,N_1529);
and U8181 (N_8181,N_5642,N_3795);
and U8182 (N_8182,N_3550,N_917);
and U8183 (N_8183,N_1305,N_4123);
nand U8184 (N_8184,N_3122,N_112);
xor U8185 (N_8185,N_2707,N_5035);
nand U8186 (N_8186,N_625,N_3443);
nand U8187 (N_8187,N_4115,N_385);
nor U8188 (N_8188,N_3047,N_202);
nand U8189 (N_8189,N_121,N_4813);
or U8190 (N_8190,N_1484,N_458);
nand U8191 (N_8191,N_3760,N_5286);
nand U8192 (N_8192,N_164,N_4104);
nor U8193 (N_8193,N_2460,N_2801);
and U8194 (N_8194,N_3603,N_3526);
or U8195 (N_8195,N_3606,N_2896);
nand U8196 (N_8196,N_2323,N_4818);
and U8197 (N_8197,N_3492,N_1608);
and U8198 (N_8198,N_1040,N_3689);
and U8199 (N_8199,N_1164,N_919);
xor U8200 (N_8200,N_3902,N_2945);
and U8201 (N_8201,N_5614,N_3466);
nand U8202 (N_8202,N_1973,N_4287);
nor U8203 (N_8203,N_4439,N_175);
nand U8204 (N_8204,N_4899,N_3480);
and U8205 (N_8205,N_4765,N_3513);
nor U8206 (N_8206,N_1088,N_778);
and U8207 (N_8207,N_746,N_2134);
and U8208 (N_8208,N_4879,N_285);
nand U8209 (N_8209,N_4467,N_5280);
nor U8210 (N_8210,N_3558,N_4789);
and U8211 (N_8211,N_421,N_4411);
nand U8212 (N_8212,N_4541,N_3251);
and U8213 (N_8213,N_3858,N_2661);
and U8214 (N_8214,N_518,N_5811);
and U8215 (N_8215,N_274,N_1722);
nand U8216 (N_8216,N_3856,N_2975);
and U8217 (N_8217,N_3313,N_3298);
or U8218 (N_8218,N_5808,N_5194);
and U8219 (N_8219,N_829,N_3007);
and U8220 (N_8220,N_77,N_1507);
nand U8221 (N_8221,N_3425,N_4354);
or U8222 (N_8222,N_3712,N_5969);
nor U8223 (N_8223,N_237,N_3489);
or U8224 (N_8224,N_4728,N_1583);
nor U8225 (N_8225,N_649,N_2780);
nor U8226 (N_8226,N_1279,N_1863);
nor U8227 (N_8227,N_4793,N_5481);
xnor U8228 (N_8228,N_2667,N_2104);
nand U8229 (N_8229,N_348,N_2626);
or U8230 (N_8230,N_882,N_5365);
nand U8231 (N_8231,N_2156,N_3699);
and U8232 (N_8232,N_75,N_2654);
and U8233 (N_8233,N_756,N_539);
or U8234 (N_8234,N_3816,N_3465);
xnor U8235 (N_8235,N_2760,N_46);
nand U8236 (N_8236,N_430,N_3010);
nor U8237 (N_8237,N_4188,N_3906);
and U8238 (N_8238,N_328,N_1686);
xnor U8239 (N_8239,N_2551,N_3038);
or U8240 (N_8240,N_4361,N_203);
nand U8241 (N_8241,N_5158,N_3542);
and U8242 (N_8242,N_4316,N_34);
nand U8243 (N_8243,N_207,N_1265);
nand U8244 (N_8244,N_5256,N_644);
nor U8245 (N_8245,N_344,N_4377);
nor U8246 (N_8246,N_1471,N_581);
nand U8247 (N_8247,N_2196,N_1458);
and U8248 (N_8248,N_1715,N_546);
and U8249 (N_8249,N_3805,N_2218);
xnor U8250 (N_8250,N_5629,N_986);
or U8251 (N_8251,N_2286,N_3104);
or U8252 (N_8252,N_1339,N_616);
nand U8253 (N_8253,N_2784,N_4386);
and U8254 (N_8254,N_1571,N_1335);
xor U8255 (N_8255,N_947,N_4621);
nand U8256 (N_8256,N_606,N_4602);
nor U8257 (N_8257,N_3508,N_3374);
nand U8258 (N_8258,N_2907,N_479);
nand U8259 (N_8259,N_2195,N_4510);
nand U8260 (N_8260,N_1224,N_3091);
xnor U8261 (N_8261,N_4855,N_2379);
nor U8262 (N_8262,N_1181,N_3546);
nand U8263 (N_8263,N_786,N_5921);
nor U8264 (N_8264,N_1577,N_1667);
and U8265 (N_8265,N_3667,N_178);
and U8266 (N_8266,N_1729,N_5778);
or U8267 (N_8267,N_424,N_4157);
and U8268 (N_8268,N_4634,N_3923);
or U8269 (N_8269,N_5258,N_3098);
and U8270 (N_8270,N_4016,N_4448);
and U8271 (N_8271,N_2959,N_1406);
and U8272 (N_8272,N_3609,N_4029);
xor U8273 (N_8273,N_975,N_2636);
xnor U8274 (N_8274,N_4827,N_5551);
nor U8275 (N_8275,N_1218,N_3720);
or U8276 (N_8276,N_5180,N_4478);
nand U8277 (N_8277,N_2148,N_5190);
nor U8278 (N_8278,N_5434,N_4816);
nor U8279 (N_8279,N_2339,N_3255);
and U8280 (N_8280,N_69,N_5118);
and U8281 (N_8281,N_4200,N_3001);
nor U8282 (N_8282,N_1441,N_3928);
nor U8283 (N_8283,N_5105,N_5701);
nor U8284 (N_8284,N_871,N_995);
nor U8285 (N_8285,N_5710,N_4211);
nand U8286 (N_8286,N_3832,N_2234);
or U8287 (N_8287,N_3533,N_367);
and U8288 (N_8288,N_1794,N_1919);
or U8289 (N_8289,N_3648,N_1103);
nand U8290 (N_8290,N_2080,N_2407);
or U8291 (N_8291,N_2140,N_234);
nand U8292 (N_8292,N_2461,N_1610);
and U8293 (N_8293,N_3618,N_1684);
and U8294 (N_8294,N_2183,N_1707);
nand U8295 (N_8295,N_5032,N_2174);
xor U8296 (N_8296,N_3585,N_3716);
xnor U8297 (N_8297,N_3142,N_1008);
nand U8298 (N_8298,N_1945,N_5439);
or U8299 (N_8299,N_3963,N_3851);
nand U8300 (N_8300,N_4915,N_117);
nand U8301 (N_8301,N_526,N_3574);
and U8302 (N_8302,N_3232,N_2910);
or U8303 (N_8303,N_5797,N_5564);
nor U8304 (N_8304,N_1013,N_794);
nor U8305 (N_8305,N_1680,N_1682);
nor U8306 (N_8306,N_5598,N_5282);
nor U8307 (N_8307,N_4721,N_4805);
nor U8308 (N_8308,N_4026,N_557);
and U8309 (N_8309,N_5847,N_2745);
nor U8310 (N_8310,N_4637,N_252);
nand U8311 (N_8311,N_968,N_1395);
nand U8312 (N_8312,N_2976,N_5199);
nand U8313 (N_8313,N_5448,N_4598);
nand U8314 (N_8314,N_5361,N_2348);
and U8315 (N_8315,N_4292,N_3999);
xor U8316 (N_8316,N_552,N_57);
nand U8317 (N_8317,N_3635,N_3958);
xor U8318 (N_8318,N_2756,N_1735);
and U8319 (N_8319,N_3333,N_1215);
nand U8320 (N_8320,N_2000,N_3005);
nor U8321 (N_8321,N_2102,N_2927);
and U8322 (N_8322,N_1595,N_2887);
or U8323 (N_8323,N_5242,N_4005);
nand U8324 (N_8324,N_4935,N_5950);
nor U8325 (N_8325,N_3265,N_4267);
or U8326 (N_8326,N_4172,N_4169);
xnor U8327 (N_8327,N_3503,N_5130);
xnor U8328 (N_8328,N_1666,N_4823);
nor U8329 (N_8329,N_340,N_2212);
xnor U8330 (N_8330,N_2853,N_5507);
or U8331 (N_8331,N_908,N_5913);
nor U8332 (N_8332,N_4089,N_802);
or U8333 (N_8333,N_1582,N_4063);
nor U8334 (N_8334,N_4463,N_3676);
or U8335 (N_8335,N_5977,N_1861);
nand U8336 (N_8336,N_4220,N_1100);
nor U8337 (N_8337,N_856,N_2921);
and U8338 (N_8338,N_3201,N_776);
or U8339 (N_8339,N_5488,N_3717);
or U8340 (N_8340,N_5684,N_4182);
or U8341 (N_8341,N_3281,N_143);
xor U8342 (N_8342,N_4293,N_3388);
nor U8343 (N_8343,N_2538,N_1063);
nor U8344 (N_8344,N_814,N_5902);
or U8345 (N_8345,N_774,N_4469);
and U8346 (N_8346,N_5420,N_2045);
nor U8347 (N_8347,N_3328,N_3739);
xnor U8348 (N_8348,N_589,N_1476);
nand U8349 (N_8349,N_3881,N_460);
xnor U8350 (N_8350,N_271,N_926);
or U8351 (N_8351,N_1256,N_5539);
xor U8352 (N_8352,N_5589,N_3571);
or U8353 (N_8353,N_4605,N_2078);
xor U8354 (N_8354,N_2637,N_132);
nor U8355 (N_8355,N_1234,N_3257);
nor U8356 (N_8356,N_4194,N_4662);
nand U8357 (N_8357,N_5999,N_4403);
and U8358 (N_8358,N_2914,N_4141);
nor U8359 (N_8359,N_2826,N_2563);
or U8360 (N_8360,N_5444,N_3479);
nand U8361 (N_8361,N_3420,N_4592);
xnor U8362 (N_8362,N_2755,N_2265);
or U8363 (N_8363,N_5299,N_1023);
and U8364 (N_8364,N_807,N_1984);
and U8365 (N_8365,N_3318,N_533);
and U8366 (N_8366,N_5619,N_2520);
nand U8367 (N_8367,N_1449,N_174);
nand U8368 (N_8368,N_1806,N_1541);
nand U8369 (N_8369,N_2235,N_2579);
nand U8370 (N_8370,N_2859,N_2362);
or U8371 (N_8371,N_1706,N_3302);
nand U8372 (N_8372,N_4396,N_2188);
nor U8373 (N_8373,N_3686,N_247);
and U8374 (N_8374,N_5253,N_3702);
nor U8375 (N_8375,N_4122,N_715);
and U8376 (N_8376,N_3736,N_4981);
xor U8377 (N_8377,N_1803,N_3132);
nand U8378 (N_8378,N_4757,N_2165);
and U8379 (N_8379,N_3453,N_1658);
xor U8380 (N_8380,N_56,N_1953);
or U8381 (N_8381,N_5517,N_5484);
nand U8382 (N_8382,N_5606,N_44);
and U8383 (N_8383,N_3355,N_5502);
or U8384 (N_8384,N_8,N_4764);
and U8385 (N_8385,N_276,N_2550);
nor U8386 (N_8386,N_665,N_3873);
nand U8387 (N_8387,N_3077,N_3017);
and U8388 (N_8388,N_1060,N_5076);
or U8389 (N_8389,N_5475,N_3387);
nor U8390 (N_8390,N_378,N_5378);
nand U8391 (N_8391,N_1775,N_1071);
and U8392 (N_8392,N_5675,N_1388);
nor U8393 (N_8393,N_4618,N_3112);
and U8394 (N_8394,N_5810,N_1928);
xnor U8395 (N_8395,N_3756,N_4394);
or U8396 (N_8396,N_5669,N_5460);
or U8397 (N_8397,N_1101,N_5091);
xor U8398 (N_8398,N_4166,N_5308);
or U8399 (N_8399,N_2602,N_3824);
or U8400 (N_8400,N_2115,N_1117);
nand U8401 (N_8401,N_2757,N_3874);
and U8402 (N_8402,N_3179,N_2281);
or U8403 (N_8403,N_2872,N_5546);
or U8404 (N_8404,N_2947,N_1465);
or U8405 (N_8405,N_5315,N_5120);
nand U8406 (N_8406,N_3604,N_3732);
nand U8407 (N_8407,N_1657,N_4625);
or U8408 (N_8408,N_3708,N_2943);
nor U8409 (N_8409,N_4207,N_3687);
and U8410 (N_8410,N_2555,N_5101);
nor U8411 (N_8411,N_2670,N_4751);
and U8412 (N_8412,N_3169,N_5964);
or U8413 (N_8413,N_2127,N_497);
nor U8414 (N_8414,N_1659,N_1816);
and U8415 (N_8415,N_3534,N_1821);
or U8416 (N_8416,N_288,N_4212);
or U8417 (N_8417,N_2557,N_3024);
and U8418 (N_8418,N_2268,N_343);
nor U8419 (N_8419,N_1121,N_5255);
or U8420 (N_8420,N_3032,N_269);
nor U8421 (N_8421,N_3196,N_5982);
and U8422 (N_8422,N_1095,N_3582);
and U8423 (N_8423,N_3187,N_5705);
or U8424 (N_8424,N_1167,N_1204);
and U8425 (N_8425,N_4051,N_2794);
nor U8426 (N_8426,N_2771,N_3888);
nor U8427 (N_8427,N_847,N_111);
and U8428 (N_8428,N_3069,N_3649);
nor U8429 (N_8429,N_3917,N_5829);
and U8430 (N_8430,N_723,N_510);
or U8431 (N_8431,N_5358,N_795);
or U8432 (N_8432,N_2915,N_5839);
or U8433 (N_8433,N_4910,N_2622);
and U8434 (N_8434,N_4388,N_2425);
or U8435 (N_8435,N_2283,N_900);
and U8436 (N_8436,N_2465,N_5856);
and U8437 (N_8437,N_4837,N_1287);
nor U8438 (N_8438,N_3321,N_5833);
xnor U8439 (N_8439,N_854,N_3987);
nor U8440 (N_8440,N_1714,N_4311);
and U8441 (N_8441,N_5195,N_5023);
nor U8442 (N_8442,N_3437,N_2296);
nor U8443 (N_8443,N_5941,N_265);
and U8444 (N_8444,N_3483,N_1996);
and U8445 (N_8445,N_5995,N_1396);
nand U8446 (N_8446,N_1585,N_2558);
nand U8447 (N_8447,N_1633,N_108);
and U8448 (N_8448,N_741,N_3872);
or U8449 (N_8449,N_5283,N_3968);
nand U8450 (N_8450,N_2913,N_3414);
nand U8451 (N_8451,N_4318,N_3804);
nand U8452 (N_8452,N_4578,N_3081);
nand U8453 (N_8453,N_4677,N_861);
nor U8454 (N_8454,N_2925,N_3664);
nor U8455 (N_8455,N_2882,N_3640);
nor U8456 (N_8456,N_5906,N_3089);
or U8457 (N_8457,N_1810,N_4753);
nor U8458 (N_8458,N_4558,N_2738);
and U8459 (N_8459,N_3730,N_2608);
nor U8460 (N_8460,N_4150,N_5997);
and U8461 (N_8461,N_3402,N_4887);
or U8462 (N_8462,N_4604,N_434);
or U8463 (N_8463,N_4482,N_749);
or U8464 (N_8464,N_5486,N_689);
and U8465 (N_8465,N_2307,N_180);
nor U8466 (N_8466,N_235,N_3630);
nand U8467 (N_8467,N_507,N_26);
and U8468 (N_8468,N_5187,N_4986);
or U8469 (N_8469,N_5430,N_4950);
or U8470 (N_8470,N_1019,N_2217);
xnor U8471 (N_8471,N_1802,N_5751);
or U8472 (N_8472,N_5883,N_1859);
nor U8473 (N_8473,N_2186,N_5090);
and U8474 (N_8474,N_1488,N_2040);
or U8475 (N_8475,N_4952,N_4822);
nand U8476 (N_8476,N_4635,N_1393);
or U8477 (N_8477,N_4383,N_831);
nor U8478 (N_8478,N_4576,N_264);
and U8479 (N_8479,N_4796,N_1925);
nor U8480 (N_8480,N_1580,N_2459);
or U8481 (N_8481,N_4209,N_580);
nor U8482 (N_8482,N_1636,N_5263);
and U8483 (N_8483,N_2099,N_1356);
or U8484 (N_8484,N_2364,N_3110);
or U8485 (N_8485,N_4560,N_5077);
nor U8486 (N_8486,N_5093,N_4814);
nand U8487 (N_8487,N_1401,N_5748);
nand U8488 (N_8488,N_1651,N_167);
nand U8489 (N_8489,N_2714,N_4070);
and U8490 (N_8490,N_5334,N_3583);
nor U8491 (N_8491,N_5391,N_2301);
or U8492 (N_8492,N_548,N_4250);
nand U8493 (N_8493,N_2349,N_256);
and U8494 (N_8494,N_2288,N_224);
nor U8495 (N_8495,N_2987,N_244);
and U8496 (N_8496,N_4846,N_1299);
xnor U8497 (N_8497,N_2509,N_5661);
xnor U8498 (N_8498,N_215,N_726);
or U8499 (N_8499,N_1620,N_4103);
nor U8500 (N_8500,N_2733,N_4201);
nand U8501 (N_8501,N_1756,N_2926);
and U8502 (N_8502,N_5266,N_1578);
nand U8503 (N_8503,N_1904,N_1172);
nand U8504 (N_8504,N_258,N_5718);
nor U8505 (N_8505,N_3491,N_60);
nand U8506 (N_8506,N_415,N_5193);
and U8507 (N_8507,N_3605,N_1542);
or U8508 (N_8508,N_3448,N_5638);
or U8509 (N_8509,N_1545,N_4908);
nor U8510 (N_8510,N_5386,N_3993);
xnor U8511 (N_8511,N_101,N_4498);
nand U8512 (N_8512,N_3944,N_4713);
nor U8513 (N_8513,N_4142,N_5176);
and U8514 (N_8514,N_2589,N_3380);
or U8515 (N_8515,N_3548,N_2052);
nand U8516 (N_8516,N_5892,N_3329);
nor U8517 (N_8517,N_5442,N_2517);
nor U8518 (N_8518,N_5314,N_2485);
xnor U8519 (N_8519,N_4650,N_1188);
or U8520 (N_8520,N_474,N_1016);
nand U8521 (N_8521,N_940,N_1140);
or U8522 (N_8522,N_2248,N_1551);
nand U8523 (N_8523,N_3749,N_4008);
nand U8524 (N_8524,N_4179,N_2222);
or U8525 (N_8525,N_4193,N_134);
and U8526 (N_8526,N_3539,N_1452);
nand U8527 (N_8527,N_1146,N_173);
nor U8528 (N_8528,N_532,N_151);
nor U8529 (N_8529,N_677,N_1087);
and U8530 (N_8530,N_4304,N_3697);
nor U8531 (N_8531,N_5493,N_377);
nand U8532 (N_8532,N_1148,N_2170);
and U8533 (N_8533,N_3252,N_3459);
nor U8534 (N_8534,N_1474,N_291);
nand U8535 (N_8535,N_2539,N_456);
and U8536 (N_8536,N_4109,N_5813);
nand U8537 (N_8537,N_3579,N_2843);
nor U8538 (N_8538,N_2270,N_1357);
and U8539 (N_8539,N_5393,N_5217);
and U8540 (N_8540,N_1748,N_1376);
nand U8541 (N_8541,N_1390,N_3661);
and U8542 (N_8542,N_2249,N_5230);
and U8543 (N_8543,N_4488,N_5556);
and U8544 (N_8544,N_4819,N_3772);
nor U8545 (N_8545,N_3598,N_139);
and U8546 (N_8546,N_480,N_4530);
or U8547 (N_8547,N_702,N_5394);
or U8548 (N_8548,N_5352,N_543);
and U8549 (N_8549,N_1051,N_1354);
nand U8550 (N_8550,N_1450,N_1638);
and U8551 (N_8551,N_3657,N_3750);
nand U8552 (N_8552,N_3096,N_5915);
or U8553 (N_8553,N_1589,N_1123);
nand U8554 (N_8554,N_2772,N_3261);
or U8555 (N_8555,N_1586,N_1618);
nand U8556 (N_8556,N_941,N_5328);
and U8557 (N_8557,N_1116,N_544);
and U8558 (N_8558,N_3430,N_835);
nand U8559 (N_8559,N_2338,N_2083);
nor U8560 (N_8560,N_4679,N_5656);
nand U8561 (N_8561,N_2750,N_5229);
and U8562 (N_8562,N_1099,N_358);
and U8563 (N_8563,N_4031,N_1352);
and U8564 (N_8564,N_5062,N_5099);
xor U8565 (N_8565,N_1774,N_4678);
xnor U8566 (N_8566,N_5935,N_4414);
nand U8567 (N_8567,N_5372,N_4208);
and U8568 (N_8568,N_3085,N_2298);
nor U8569 (N_8569,N_934,N_3789);
and U8570 (N_8570,N_190,N_5622);
nor U8571 (N_8571,N_3057,N_4296);
and U8572 (N_8572,N_2928,N_5815);
nor U8573 (N_8573,N_5189,N_191);
and U8574 (N_8574,N_2691,N_2329);
xnor U8575 (N_8575,N_4642,N_583);
xor U8576 (N_8576,N_281,N_2278);
or U8577 (N_8577,N_4532,N_4919);
nor U8578 (N_8578,N_2824,N_5246);
nor U8579 (N_8579,N_4606,N_1411);
nand U8580 (N_8580,N_3495,N_1045);
nor U8581 (N_8581,N_81,N_4918);
nand U8582 (N_8582,N_5196,N_1777);
nand U8583 (N_8583,N_323,N_5354);
nand U8584 (N_8584,N_618,N_5326);
or U8585 (N_8585,N_525,N_5634);
and U8586 (N_8586,N_4943,N_3194);
nor U8587 (N_8587,N_1790,N_2761);
nor U8588 (N_8588,N_1078,N_5547);
or U8589 (N_8589,N_979,N_4856);
or U8590 (N_8590,N_4731,N_1574);
or U8591 (N_8591,N_4922,N_3228);
nor U8592 (N_8592,N_160,N_3434);
and U8593 (N_8593,N_5850,N_3931);
nand U8594 (N_8594,N_3684,N_2668);
or U8595 (N_8595,N_3719,N_4681);
or U8596 (N_8596,N_4877,N_5382);
or U8597 (N_8597,N_5082,N_4133);
nand U8598 (N_8598,N_2663,N_1896);
or U8599 (N_8599,N_1679,N_372);
nand U8600 (N_8600,N_5384,N_4132);
or U8601 (N_8601,N_1210,N_3378);
xor U8602 (N_8602,N_3959,N_1848);
nor U8603 (N_8603,N_3802,N_1648);
xor U8604 (N_8604,N_5211,N_2712);
and U8605 (N_8605,N_1199,N_2418);
or U8606 (N_8606,N_4198,N_5252);
and U8607 (N_8607,N_5586,N_1223);
and U8608 (N_8608,N_5186,N_1183);
nand U8609 (N_8609,N_2481,N_263);
xor U8610 (N_8610,N_4147,N_2879);
nor U8611 (N_8611,N_1198,N_4259);
and U8612 (N_8612,N_3014,N_5804);
or U8613 (N_8613,N_1703,N_5750);
xor U8614 (N_8614,N_1232,N_2163);
nor U8615 (N_8615,N_3139,N_2036);
nor U8616 (N_8616,N_810,N_1321);
and U8617 (N_8617,N_2556,N_1901);
nor U8618 (N_8618,N_5836,N_4779);
or U8619 (N_8619,N_412,N_4003);
and U8620 (N_8620,N_2326,N_2276);
nand U8621 (N_8621,N_2046,N_4356);
or U8622 (N_8622,N_4515,N_1274);
and U8623 (N_8623,N_3065,N_3485);
or U8624 (N_8624,N_4704,N_5302);
or U8625 (N_8625,N_4249,N_4747);
xor U8626 (N_8626,N_2813,N_3013);
and U8627 (N_8627,N_5156,N_3581);
and U8628 (N_8628,N_5106,N_1613);
nor U8629 (N_8629,N_2763,N_2858);
nand U8630 (N_8630,N_3208,N_1108);
or U8631 (N_8631,N_1908,N_5973);
and U8632 (N_8632,N_1723,N_4917);
nor U8633 (N_8633,N_4907,N_3787);
nor U8634 (N_8634,N_3853,N_1132);
and U8635 (N_8635,N_2484,N_1668);
or U8636 (N_8636,N_2708,N_1007);
xnor U8637 (N_8637,N_1211,N_2201);
or U8638 (N_8638,N_837,N_389);
and U8639 (N_8639,N_825,N_1995);
nor U8640 (N_8640,N_4932,N_4059);
or U8641 (N_8641,N_1954,N_4353);
or U8642 (N_8642,N_4717,N_4608);
or U8643 (N_8643,N_1298,N_2779);
or U8644 (N_8644,N_3078,N_1166);
and U8645 (N_8645,N_812,N_2513);
or U8646 (N_8646,N_122,N_2097);
nand U8647 (N_8647,N_5289,N_1454);
nand U8648 (N_8648,N_3576,N_4330);
nor U8649 (N_8649,N_4565,N_494);
or U8650 (N_8650,N_4430,N_432);
or U8651 (N_8651,N_1113,N_5476);
and U8652 (N_8652,N_5449,N_1912);
and U8653 (N_8653,N_2471,N_4517);
nor U8654 (N_8654,N_3493,N_1238);
or U8655 (N_8655,N_5477,N_2850);
or U8656 (N_8656,N_5713,N_3147);
nand U8657 (N_8657,N_217,N_3800);
nand U8658 (N_8658,N_3842,N_1173);
xnor U8659 (N_8659,N_273,N_4061);
nor U8660 (N_8660,N_5985,N_1075);
and U8661 (N_8661,N_1311,N_5415);
or U8662 (N_8662,N_3811,N_1430);
nand U8663 (N_8663,N_874,N_2429);
and U8664 (N_8664,N_1231,N_468);
and U8665 (N_8665,N_690,N_4474);
nand U8666 (N_8666,N_3026,N_1372);
and U8667 (N_8667,N_1369,N_3884);
nor U8668 (N_8668,N_5991,N_4861);
xnor U8669 (N_8669,N_5681,N_1124);
nor U8670 (N_8670,N_3290,N_899);
nand U8671 (N_8671,N_1419,N_1754);
nor U8672 (N_8672,N_1240,N_1769);
xnor U8673 (N_8673,N_4335,N_5624);
or U8674 (N_8674,N_2411,N_5214);
or U8675 (N_8675,N_1190,N_391);
nand U8676 (N_8676,N_4978,N_5273);
nand U8677 (N_8677,N_5509,N_2419);
or U8678 (N_8678,N_485,N_205);
xnor U8679 (N_8679,N_978,N_664);
or U8680 (N_8680,N_5989,N_212);
nor U8681 (N_8681,N_1505,N_1448);
xor U8682 (N_8682,N_394,N_1136);
nor U8683 (N_8683,N_5514,N_5017);
or U8684 (N_8684,N_1860,N_729);
or U8685 (N_8685,N_3882,N_1832);
nand U8686 (N_8686,N_5414,N_4852);
xor U8687 (N_8687,N_2686,N_170);
nor U8688 (N_8688,N_5132,N_1738);
or U8689 (N_8689,N_103,N_3547);
xor U8690 (N_8690,N_1206,N_780);
nand U8691 (N_8691,N_4340,N_5770);
or U8692 (N_8692,N_2901,N_1269);
and U8693 (N_8693,N_2701,N_712);
or U8694 (N_8694,N_2111,N_4900);
nor U8695 (N_8695,N_3246,N_2309);
xnor U8696 (N_8696,N_881,N_5145);
xnor U8697 (N_8697,N_3674,N_3097);
and U8698 (N_8698,N_2931,N_600);
and U8699 (N_8699,N_797,N_5064);
nand U8700 (N_8700,N_1997,N_5852);
or U8701 (N_8701,N_4441,N_5536);
and U8702 (N_8702,N_4435,N_2360);
and U8703 (N_8703,N_1615,N_1135);
nand U8704 (N_8704,N_1437,N_3263);
xor U8705 (N_8705,N_1753,N_1564);
and U8706 (N_8706,N_4524,N_1351);
nand U8707 (N_8707,N_1490,N_905);
nand U8708 (N_8708,N_2819,N_2841);
and U8709 (N_8709,N_3901,N_3698);
nand U8710 (N_8710,N_662,N_5126);
nand U8711 (N_8711,N_439,N_4428);
nor U8712 (N_8712,N_4870,N_3417);
xnor U8713 (N_8713,N_4991,N_732);
or U8714 (N_8714,N_2971,N_2587);
xnor U8715 (N_8715,N_2720,N_2073);
nand U8716 (N_8716,N_2057,N_2009);
nand U8717 (N_8717,N_4504,N_5116);
nor U8718 (N_8718,N_2868,N_705);
or U8719 (N_8719,N_2030,N_804);
nor U8720 (N_8720,N_4480,N_1747);
nand U8721 (N_8721,N_682,N_3707);
and U8722 (N_8722,N_4938,N_1422);
or U8723 (N_8723,N_4094,N_4347);
or U8724 (N_8724,N_834,N_4956);
or U8725 (N_8725,N_4336,N_568);
or U8726 (N_8726,N_4671,N_4329);
nor U8727 (N_8727,N_5644,N_2202);
nand U8728 (N_8728,N_1451,N_3494);
and U8729 (N_8729,N_2372,N_5905);
nor U8730 (N_8730,N_1012,N_4290);
and U8731 (N_8731,N_3373,N_965);
nor U8732 (N_8732,N_5880,N_3970);
or U8733 (N_8733,N_596,N_631);
and U8734 (N_8734,N_3172,N_5756);
or U8735 (N_8735,N_390,N_5875);
nand U8736 (N_8736,N_3809,N_5588);
nor U8737 (N_8737,N_4117,N_3994);
nand U8738 (N_8738,N_2617,N_4162);
nand U8739 (N_8739,N_5772,N_2473);
nand U8740 (N_8740,N_331,N_3876);
nand U8741 (N_8741,N_5771,N_3683);
and U8742 (N_8742,N_5123,N_4477);
nor U8743 (N_8743,N_3392,N_3879);
nor U8744 (N_8744,N_2719,N_2318);
or U8745 (N_8745,N_2566,N_4280);
or U8746 (N_8746,N_976,N_5930);
nor U8747 (N_8747,N_260,N_2417);
nand U8748 (N_8748,N_4453,N_3742);
or U8749 (N_8749,N_5664,N_3767);
xor U8750 (N_8750,N_3239,N_1399);
or U8751 (N_8751,N_4086,N_1540);
xnor U8752 (N_8752,N_5817,N_4471);
nor U8753 (N_8753,N_5472,N_5719);
nor U8754 (N_8754,N_3340,N_3957);
xnor U8755 (N_8755,N_4696,N_5381);
and U8756 (N_8756,N_2510,N_1705);
nand U8757 (N_8757,N_277,N_793);
or U8758 (N_8758,N_4675,N_4055);
nor U8759 (N_8759,N_4479,N_2965);
nand U8760 (N_8760,N_5039,N_4901);
nand U8761 (N_8761,N_3413,N_2180);
xor U8762 (N_8762,N_684,N_3394);
xor U8763 (N_8763,N_2233,N_2324);
or U8764 (N_8764,N_5291,N_590);
nor U8765 (N_8765,N_3358,N_5446);
nor U8766 (N_8766,N_4348,N_5026);
nand U8767 (N_8767,N_1733,N_462);
or U8768 (N_8768,N_2912,N_2768);
nor U8769 (N_8769,N_470,N_803);
and U8770 (N_8770,N_5057,N_183);
or U8771 (N_8771,N_569,N_5465);
nand U8772 (N_8772,N_4965,N_3733);
xor U8773 (N_8773,N_5727,N_5374);
or U8774 (N_8774,N_4641,N_5233);
nor U8775 (N_8775,N_1264,N_1355);
nor U8776 (N_8776,N_862,N_1933);
nor U8777 (N_8777,N_1627,N_400);
or U8778 (N_8778,N_472,N_2951);
nor U8779 (N_8779,N_3509,N_725);
nor U8780 (N_8780,N_4454,N_3272);
or U8781 (N_8781,N_5418,N_2207);
nor U8782 (N_8782,N_2025,N_4601);
or U8783 (N_8783,N_801,N_3813);
and U8784 (N_8784,N_709,N_1273);
and U8785 (N_8785,N_1065,N_1459);
and U8786 (N_8786,N_1261,N_3323);
and U8787 (N_8787,N_1882,N_309);
or U8788 (N_8788,N_5370,N_915);
or U8789 (N_8789,N_3270,N_326);
or U8790 (N_8790,N_1688,N_2130);
nor U8791 (N_8791,N_3822,N_981);
or U8792 (N_8792,N_695,N_1289);
nor U8793 (N_8793,N_1170,N_4702);
nand U8794 (N_8794,N_5697,N_334);
or U8795 (N_8795,N_2405,N_1246);
and U8796 (N_8796,N_3709,N_4543);
xor U8797 (N_8797,N_3114,N_4620);
or U8798 (N_8798,N_4422,N_3428);
xor U8799 (N_8799,N_2336,N_305);
xnor U8800 (N_8800,N_1812,N_2883);
and U8801 (N_8801,N_3675,N_1156);
or U8802 (N_8802,N_4148,N_1939);
or U8803 (N_8803,N_2982,N_841);
nand U8804 (N_8804,N_558,N_4674);
or U8805 (N_8805,N_4872,N_1478);
and U8806 (N_8806,N_2255,N_4239);
nor U8807 (N_8807,N_3905,N_131);
and U8808 (N_8808,N_1381,N_3429);
xor U8809 (N_8809,N_2477,N_4998);
nor U8810 (N_8810,N_2576,N_4352);
nor U8811 (N_8811,N_3567,N_2420);
nand U8812 (N_8812,N_4102,N_2980);
and U8813 (N_8813,N_855,N_2433);
nand U8814 (N_8814,N_1730,N_4506);
or U8815 (N_8815,N_1873,N_551);
or U8816 (N_8816,N_3183,N_3164);
nor U8817 (N_8817,N_4787,N_3330);
or U8818 (N_8818,N_2834,N_2454);
nand U8819 (N_8819,N_3350,N_5926);
and U8820 (N_8820,N_4567,N_5295);
nor U8821 (N_8821,N_2290,N_3886);
nor U8822 (N_8822,N_5889,N_613);
nor U8823 (N_8823,N_2094,N_4072);
and U8824 (N_8824,N_3405,N_748);
nand U8825 (N_8825,N_1635,N_5332);
or U8826 (N_8826,N_5135,N_1168);
or U8827 (N_8827,N_2685,N_3262);
xnor U8828 (N_8828,N_5878,N_1475);
and U8829 (N_8829,N_2303,N_1209);
xor U8830 (N_8830,N_5888,N_4615);
nand U8831 (N_8831,N_2792,N_4227);
xnor U8832 (N_8832,N_5890,N_2191);
nor U8833 (N_8833,N_444,N_3511);
or U8834 (N_8834,N_2946,N_2625);
nor U8835 (N_8835,N_565,N_2422);
nand U8836 (N_8836,N_5749,N_766);
nand U8837 (N_8837,N_4107,N_4770);
nand U8838 (N_8838,N_2567,N_4628);
nand U8839 (N_8839,N_2666,N_5716);
and U8840 (N_8840,N_4263,N_2171);
or U8841 (N_8841,N_5335,N_3248);
nor U8842 (N_8842,N_1239,N_2108);
nor U8843 (N_8843,N_2905,N_1048);
or U8844 (N_8844,N_2583,N_4011);
nor U8845 (N_8845,N_3235,N_5485);
and U8846 (N_8846,N_5059,N_3817);
or U8847 (N_8847,N_553,N_4705);
xnor U8848 (N_8848,N_5682,N_3626);
nand U8849 (N_8849,N_1607,N_4071);
or U8850 (N_8850,N_3044,N_1538);
nor U8851 (N_8851,N_800,N_5953);
nand U8852 (N_8852,N_1184,N_2793);
and U8853 (N_8853,N_2624,N_2860);
nor U8854 (N_8854,N_3212,N_2940);
nand U8855 (N_8855,N_4202,N_659);
and U8856 (N_8856,N_270,N_3283);
nand U8857 (N_8857,N_4645,N_4941);
xnor U8858 (N_8858,N_3669,N_4516);
or U8859 (N_8859,N_2600,N_4503);
nor U8860 (N_8860,N_4623,N_4691);
and U8861 (N_8861,N_4767,N_5127);
nand U8862 (N_8862,N_1504,N_2495);
and U8863 (N_8863,N_4519,N_5841);
xnor U8864 (N_8864,N_5161,N_5144);
nand U8865 (N_8865,N_106,N_5497);
nand U8866 (N_8866,N_1838,N_4309);
or U8867 (N_8867,N_692,N_4174);
and U8868 (N_8868,N_3952,N_1572);
nand U8869 (N_8869,N_5309,N_351);
xor U8870 (N_8870,N_1979,N_380);
and U8871 (N_8871,N_2166,N_5423);
and U8872 (N_8872,N_349,N_3293);
nand U8873 (N_8873,N_5005,N_2396);
nor U8874 (N_8874,N_1233,N_1642);
xnor U8875 (N_8875,N_1624,N_1086);
or U8876 (N_8876,N_4514,N_4038);
and U8877 (N_8877,N_3300,N_5947);
and U8878 (N_8878,N_4427,N_2375);
nor U8879 (N_8879,N_144,N_2072);
or U8880 (N_8880,N_5570,N_2956);
or U8881 (N_8881,N_1398,N_1187);
nor U8882 (N_8882,N_1109,N_1601);
or U8883 (N_8883,N_4895,N_2833);
nor U8884 (N_8884,N_3295,N_2991);
nor U8885 (N_8885,N_2145,N_10);
nand U8886 (N_8886,N_3893,N_5458);
and U8887 (N_8887,N_2204,N_2742);
nand U8888 (N_8888,N_3714,N_4370);
and U8889 (N_8889,N_5015,N_17);
nand U8890 (N_8890,N_4766,N_609);
and U8891 (N_8891,N_1252,N_1955);
nand U8892 (N_8892,N_4130,N_3025);
xor U8893 (N_8893,N_5054,N_1897);
and U8894 (N_8894,N_5142,N_1480);
and U8895 (N_8895,N_5666,N_204);
nand U8896 (N_8896,N_448,N_233);
nand U8897 (N_8897,N_3166,N_4444);
and U8898 (N_8898,N_3871,N_2525);
nor U8899 (N_8899,N_5967,N_2607);
nor U8900 (N_8900,N_3850,N_909);
nor U8901 (N_8901,N_4769,N_2900);
nor U8902 (N_8902,N_924,N_805);
nand U8903 (N_8903,N_1847,N_2200);
or U8904 (N_8904,N_1758,N_4891);
or U8905 (N_8905,N_9,N_5923);
nor U8906 (N_8906,N_5483,N_5755);
or U8907 (N_8907,N_3446,N_2752);
nor U8908 (N_8908,N_5245,N_1491);
and U8909 (N_8909,N_5528,N_4446);
or U8910 (N_8910,N_1970,N_3391);
nor U8911 (N_8911,N_1581,N_4737);
and U8912 (N_8912,N_5061,N_3337);
nand U8913 (N_8913,N_1647,N_5516);
and U8914 (N_8914,N_4636,N_4654);
and U8915 (N_8915,N_1982,N_2619);
xnor U8916 (N_8916,N_4156,N_5518);
xnor U8917 (N_8917,N_2151,N_2456);
and U8918 (N_8918,N_3616,N_2308);
or U8919 (N_8919,N_1377,N_1431);
or U8920 (N_8920,N_4989,N_572);
and U8921 (N_8921,N_869,N_1496);
xnor U8922 (N_8922,N_1243,N_5541);
or U8923 (N_8923,N_2816,N_3304);
nor U8924 (N_8924,N_2541,N_1531);
nand U8925 (N_8925,N_2117,N_3658);
nand U8926 (N_8926,N_4727,N_5993);
or U8927 (N_8927,N_4512,N_2351);
or U8928 (N_8928,N_813,N_653);
nor U8929 (N_8929,N_4231,N_5819);
nor U8930 (N_8930,N_1461,N_4324);
xnor U8931 (N_8931,N_169,N_5011);
or U8932 (N_8932,N_176,N_3016);
or U8933 (N_8933,N_4710,N_1884);
or U8934 (N_8934,N_2331,N_5318);
nand U8935 (N_8935,N_1820,N_1219);
or U8936 (N_8936,N_228,N_450);
or U8937 (N_8937,N_4980,N_923);
nand U8938 (N_8938,N_1342,N_2891);
and U8939 (N_8939,N_4429,N_2963);
and U8940 (N_8940,N_4326,N_407);
nand U8941 (N_8941,N_5298,N_4359);
and U8942 (N_8942,N_2753,N_4776);
or U8943 (N_8943,N_3470,N_2317);
or U8944 (N_8944,N_1700,N_3741);
nand U8945 (N_8945,N_1028,N_1255);
or U8946 (N_8946,N_3284,N_2884);
nand U8947 (N_8947,N_5660,N_4893);
nand U8948 (N_8948,N_5631,N_809);
or U8949 (N_8949,N_146,N_2672);
xnor U8950 (N_8950,N_5538,N_2213);
nand U8951 (N_8951,N_1404,N_5637);
nand U8952 (N_8952,N_4882,N_5860);
nor U8953 (N_8953,N_5238,N_5663);
or U8954 (N_8954,N_5294,N_5044);
and U8955 (N_8955,N_15,N_4841);
nand U8956 (N_8956,N_3523,N_3062);
xor U8957 (N_8957,N_2941,N_2085);
nand U8958 (N_8958,N_2272,N_4652);
nand U8959 (N_8959,N_2765,N_4307);
and U8960 (N_8960,N_2623,N_1462);
xnor U8961 (N_8961,N_5937,N_953);
and U8962 (N_8962,N_5522,N_3855);
nor U8963 (N_8963,N_2732,N_2409);
nor U8964 (N_8964,N_4423,N_5447);
nand U8965 (N_8965,N_2198,N_4116);
nand U8966 (N_8966,N_3715,N_3460);
nor U8967 (N_8967,N_4034,N_4080);
or U8968 (N_8968,N_4858,N_1438);
nor U8969 (N_8969,N_5417,N_5496);
nand U8970 (N_8970,N_1558,N_5359);
nand U8971 (N_8971,N_540,N_1194);
xnor U8972 (N_8972,N_4382,N_1017);
and U8973 (N_8973,N_4271,N_3258);
nor U8974 (N_8974,N_2267,N_4817);
and U8975 (N_8975,N_5259,N_5577);
xnor U8976 (N_8976,N_4523,N_5601);
nand U8977 (N_8977,N_4334,N_781);
nor U8978 (N_8978,N_5022,N_842);
and U8979 (N_8979,N_4502,N_94);
and U8980 (N_8980,N_545,N_2775);
and U8981 (N_8981,N_1566,N_2053);
and U8982 (N_8982,N_4794,N_679);
xor U8983 (N_8983,N_1043,N_4185);
nand U8984 (N_8984,N_5173,N_992);
xor U8985 (N_8985,N_4276,N_3288);
and U8986 (N_8986,N_374,N_2803);
or U8987 (N_8987,N_1559,N_4355);
and U8988 (N_8988,N_2246,N_1338);
or U8989 (N_8989,N_704,N_5563);
nand U8990 (N_8990,N_1152,N_3735);
nor U8991 (N_8991,N_72,N_5851);
nor U8992 (N_8992,N_5708,N_1107);
and U8993 (N_8993,N_5757,N_5089);
and U8994 (N_8994,N_5290,N_3099);
nand U8995 (N_8995,N_560,N_826);
nand U8996 (N_8996,N_5625,N_1768);
and U8997 (N_8997,N_5956,N_3128);
and U8998 (N_8998,N_4392,N_4243);
and U8999 (N_8999,N_1035,N_1550);
nor U9000 (N_9000,N_1827,N_4682);
xor U9001 (N_9001,N_5478,N_2715);
nor U9002 (N_9002,N_3956,N_2115);
nand U9003 (N_9003,N_3399,N_4145);
nand U9004 (N_9004,N_1585,N_959);
nand U9005 (N_9005,N_1121,N_483);
and U9006 (N_9006,N_4402,N_1913);
nand U9007 (N_9007,N_3755,N_4438);
nand U9008 (N_9008,N_5481,N_5207);
nor U9009 (N_9009,N_3751,N_5673);
and U9010 (N_9010,N_4489,N_4942);
nand U9011 (N_9011,N_4937,N_3265);
or U9012 (N_9012,N_2794,N_5302);
nor U9013 (N_9013,N_634,N_3556);
and U9014 (N_9014,N_4979,N_3656);
xnor U9015 (N_9015,N_2841,N_5980);
or U9016 (N_9016,N_2498,N_4685);
nand U9017 (N_9017,N_1271,N_5520);
and U9018 (N_9018,N_4344,N_5280);
and U9019 (N_9019,N_5524,N_3280);
xor U9020 (N_9020,N_3893,N_2261);
nand U9021 (N_9021,N_2203,N_3904);
nand U9022 (N_9022,N_5930,N_3603);
and U9023 (N_9023,N_5468,N_3020);
nor U9024 (N_9024,N_216,N_2792);
and U9025 (N_9025,N_1241,N_5429);
and U9026 (N_9026,N_5738,N_813);
or U9027 (N_9027,N_4256,N_3256);
nor U9028 (N_9028,N_3337,N_4227);
or U9029 (N_9029,N_4606,N_2341);
nand U9030 (N_9030,N_5404,N_5691);
nor U9031 (N_9031,N_5098,N_4149);
and U9032 (N_9032,N_1649,N_3258);
nand U9033 (N_9033,N_5355,N_3685);
xor U9034 (N_9034,N_3713,N_5424);
nand U9035 (N_9035,N_5213,N_1996);
and U9036 (N_9036,N_1372,N_448);
or U9037 (N_9037,N_5941,N_3506);
nor U9038 (N_9038,N_4046,N_1605);
nor U9039 (N_9039,N_2822,N_347);
nand U9040 (N_9040,N_1550,N_944);
or U9041 (N_9041,N_526,N_3569);
nand U9042 (N_9042,N_710,N_4746);
or U9043 (N_9043,N_975,N_5464);
and U9044 (N_9044,N_2655,N_1082);
nand U9045 (N_9045,N_3460,N_4615);
xor U9046 (N_9046,N_2287,N_1375);
and U9047 (N_9047,N_5282,N_2671);
or U9048 (N_9048,N_2456,N_2224);
or U9049 (N_9049,N_3916,N_2244);
nand U9050 (N_9050,N_4404,N_2644);
nand U9051 (N_9051,N_740,N_1845);
and U9052 (N_9052,N_344,N_5715);
or U9053 (N_9053,N_5124,N_1164);
or U9054 (N_9054,N_204,N_5258);
nand U9055 (N_9055,N_3672,N_2359);
nor U9056 (N_9056,N_4484,N_2494);
nor U9057 (N_9057,N_563,N_30);
or U9058 (N_9058,N_1127,N_1101);
nor U9059 (N_9059,N_141,N_1416);
nand U9060 (N_9060,N_4124,N_237);
xnor U9061 (N_9061,N_2152,N_2144);
nand U9062 (N_9062,N_842,N_1402);
or U9063 (N_9063,N_3722,N_668);
nor U9064 (N_9064,N_4519,N_665);
or U9065 (N_9065,N_4260,N_3810);
or U9066 (N_9066,N_1916,N_1861);
and U9067 (N_9067,N_4546,N_4197);
nand U9068 (N_9068,N_3403,N_3486);
or U9069 (N_9069,N_4082,N_2694);
nand U9070 (N_9070,N_2310,N_3591);
or U9071 (N_9071,N_1774,N_5039);
nor U9072 (N_9072,N_2821,N_2878);
nor U9073 (N_9073,N_3358,N_3133);
xnor U9074 (N_9074,N_2203,N_844);
and U9075 (N_9075,N_3751,N_4678);
xnor U9076 (N_9076,N_3423,N_4026);
nand U9077 (N_9077,N_4760,N_2816);
and U9078 (N_9078,N_5502,N_3282);
nor U9079 (N_9079,N_4710,N_5988);
nand U9080 (N_9080,N_4514,N_1825);
nand U9081 (N_9081,N_3172,N_3557);
and U9082 (N_9082,N_928,N_3766);
and U9083 (N_9083,N_4683,N_1783);
nand U9084 (N_9084,N_2363,N_4480);
nor U9085 (N_9085,N_4921,N_5584);
nand U9086 (N_9086,N_5872,N_5394);
nand U9087 (N_9087,N_3298,N_908);
nand U9088 (N_9088,N_4878,N_5696);
or U9089 (N_9089,N_5237,N_2302);
nor U9090 (N_9090,N_3384,N_4219);
and U9091 (N_9091,N_421,N_4435);
and U9092 (N_9092,N_3199,N_529);
nand U9093 (N_9093,N_1453,N_4051);
and U9094 (N_9094,N_5978,N_571);
or U9095 (N_9095,N_5359,N_3653);
nor U9096 (N_9096,N_1009,N_1115);
or U9097 (N_9097,N_3878,N_2412);
xor U9098 (N_9098,N_4797,N_566);
and U9099 (N_9099,N_4454,N_683);
or U9100 (N_9100,N_1921,N_4974);
or U9101 (N_9101,N_4244,N_1880);
nor U9102 (N_9102,N_5877,N_3807);
xnor U9103 (N_9103,N_2728,N_823);
nor U9104 (N_9104,N_3565,N_1794);
and U9105 (N_9105,N_1816,N_3845);
nand U9106 (N_9106,N_4819,N_304);
nand U9107 (N_9107,N_3773,N_3);
nor U9108 (N_9108,N_867,N_282);
nor U9109 (N_9109,N_94,N_4117);
and U9110 (N_9110,N_4900,N_4348);
nand U9111 (N_9111,N_2586,N_5565);
nor U9112 (N_9112,N_3224,N_564);
or U9113 (N_9113,N_2437,N_5150);
xor U9114 (N_9114,N_866,N_2603);
or U9115 (N_9115,N_13,N_57);
nand U9116 (N_9116,N_5847,N_2591);
and U9117 (N_9117,N_3114,N_136);
and U9118 (N_9118,N_3677,N_1661);
nor U9119 (N_9119,N_3038,N_2377);
or U9120 (N_9120,N_504,N_3439);
and U9121 (N_9121,N_5011,N_1082);
nand U9122 (N_9122,N_2706,N_3138);
nand U9123 (N_9123,N_863,N_566);
and U9124 (N_9124,N_4341,N_4738);
nor U9125 (N_9125,N_2024,N_2937);
nand U9126 (N_9126,N_5339,N_1493);
nand U9127 (N_9127,N_4471,N_682);
and U9128 (N_9128,N_3279,N_4344);
and U9129 (N_9129,N_2105,N_2551);
xor U9130 (N_9130,N_3346,N_5357);
or U9131 (N_9131,N_2272,N_5312);
or U9132 (N_9132,N_1309,N_2434);
nor U9133 (N_9133,N_1309,N_845);
nand U9134 (N_9134,N_5293,N_5119);
or U9135 (N_9135,N_5175,N_5107);
nor U9136 (N_9136,N_167,N_4759);
nand U9137 (N_9137,N_5223,N_5556);
xnor U9138 (N_9138,N_5820,N_2195);
or U9139 (N_9139,N_1137,N_5657);
xnor U9140 (N_9140,N_4764,N_2019);
nand U9141 (N_9141,N_2145,N_461);
nor U9142 (N_9142,N_137,N_4679);
or U9143 (N_9143,N_5833,N_2991);
xnor U9144 (N_9144,N_4712,N_5610);
nand U9145 (N_9145,N_4201,N_4757);
and U9146 (N_9146,N_48,N_5430);
and U9147 (N_9147,N_2726,N_2553);
nand U9148 (N_9148,N_791,N_1211);
nand U9149 (N_9149,N_5821,N_1288);
xor U9150 (N_9150,N_4531,N_869);
nand U9151 (N_9151,N_3042,N_3324);
and U9152 (N_9152,N_2195,N_3941);
nor U9153 (N_9153,N_2432,N_2428);
or U9154 (N_9154,N_1944,N_1218);
nand U9155 (N_9155,N_1531,N_4422);
or U9156 (N_9156,N_3176,N_4695);
and U9157 (N_9157,N_596,N_1091);
nor U9158 (N_9158,N_2149,N_3137);
nor U9159 (N_9159,N_4508,N_4092);
nor U9160 (N_9160,N_190,N_1643);
nand U9161 (N_9161,N_5579,N_2341);
and U9162 (N_9162,N_1280,N_791);
or U9163 (N_9163,N_5401,N_1597);
or U9164 (N_9164,N_1082,N_4330);
nor U9165 (N_9165,N_519,N_2088);
nor U9166 (N_9166,N_5632,N_4480);
nand U9167 (N_9167,N_3754,N_4753);
nand U9168 (N_9168,N_280,N_399);
nor U9169 (N_9169,N_5027,N_1918);
nand U9170 (N_9170,N_3643,N_1565);
and U9171 (N_9171,N_708,N_112);
nand U9172 (N_9172,N_5538,N_4752);
and U9173 (N_9173,N_2912,N_1590);
or U9174 (N_9174,N_5105,N_5942);
nand U9175 (N_9175,N_1032,N_4266);
and U9176 (N_9176,N_3901,N_1511);
or U9177 (N_9177,N_1449,N_2808);
nor U9178 (N_9178,N_4500,N_4873);
nand U9179 (N_9179,N_2292,N_4153);
nand U9180 (N_9180,N_2645,N_3509);
nor U9181 (N_9181,N_5800,N_3220);
and U9182 (N_9182,N_1500,N_1906);
and U9183 (N_9183,N_5218,N_5193);
or U9184 (N_9184,N_3714,N_948);
xnor U9185 (N_9185,N_4625,N_5782);
nand U9186 (N_9186,N_917,N_2935);
xor U9187 (N_9187,N_3684,N_1317);
and U9188 (N_9188,N_4069,N_4183);
nor U9189 (N_9189,N_1332,N_5902);
or U9190 (N_9190,N_4052,N_4004);
xor U9191 (N_9191,N_3715,N_1438);
and U9192 (N_9192,N_3976,N_1751);
and U9193 (N_9193,N_5247,N_3577);
and U9194 (N_9194,N_1408,N_3026);
nand U9195 (N_9195,N_3696,N_4433);
or U9196 (N_9196,N_2993,N_5363);
or U9197 (N_9197,N_113,N_1464);
and U9198 (N_9198,N_4355,N_5980);
and U9199 (N_9199,N_5259,N_75);
nand U9200 (N_9200,N_1219,N_5456);
or U9201 (N_9201,N_960,N_5110);
nand U9202 (N_9202,N_4998,N_611);
xnor U9203 (N_9203,N_605,N_567);
or U9204 (N_9204,N_5928,N_5894);
and U9205 (N_9205,N_608,N_3799);
or U9206 (N_9206,N_1123,N_3321);
nand U9207 (N_9207,N_1501,N_2690);
nor U9208 (N_9208,N_3745,N_4300);
and U9209 (N_9209,N_5029,N_1026);
nand U9210 (N_9210,N_5337,N_5398);
and U9211 (N_9211,N_3137,N_2395);
nor U9212 (N_9212,N_3772,N_2568);
nor U9213 (N_9213,N_3821,N_1326);
and U9214 (N_9214,N_3550,N_1894);
nor U9215 (N_9215,N_2865,N_5824);
nor U9216 (N_9216,N_435,N_3612);
nor U9217 (N_9217,N_2659,N_2184);
and U9218 (N_9218,N_4197,N_4510);
and U9219 (N_9219,N_2714,N_5714);
nor U9220 (N_9220,N_3640,N_29);
xnor U9221 (N_9221,N_2081,N_3917);
or U9222 (N_9222,N_5073,N_1668);
and U9223 (N_9223,N_2344,N_3941);
nor U9224 (N_9224,N_1265,N_4346);
nand U9225 (N_9225,N_685,N_495);
or U9226 (N_9226,N_2834,N_3684);
or U9227 (N_9227,N_1385,N_1599);
and U9228 (N_9228,N_3827,N_5343);
nor U9229 (N_9229,N_4056,N_3088);
and U9230 (N_9230,N_4584,N_158);
nor U9231 (N_9231,N_5898,N_697);
nand U9232 (N_9232,N_1422,N_3785);
or U9233 (N_9233,N_272,N_3982);
nand U9234 (N_9234,N_5464,N_5412);
and U9235 (N_9235,N_5964,N_2206);
and U9236 (N_9236,N_3677,N_3342);
nand U9237 (N_9237,N_4130,N_3080);
or U9238 (N_9238,N_1331,N_5810);
nand U9239 (N_9239,N_202,N_3098);
or U9240 (N_9240,N_1012,N_5316);
nand U9241 (N_9241,N_3950,N_814);
or U9242 (N_9242,N_3330,N_2988);
nand U9243 (N_9243,N_1555,N_4362);
xnor U9244 (N_9244,N_1959,N_2694);
nor U9245 (N_9245,N_5990,N_3165);
nor U9246 (N_9246,N_3287,N_845);
and U9247 (N_9247,N_1146,N_5835);
nand U9248 (N_9248,N_763,N_3618);
nand U9249 (N_9249,N_5143,N_182);
xor U9250 (N_9250,N_3474,N_918);
or U9251 (N_9251,N_3539,N_1122);
nand U9252 (N_9252,N_5444,N_5151);
or U9253 (N_9253,N_5125,N_3713);
nor U9254 (N_9254,N_3875,N_4358);
or U9255 (N_9255,N_2436,N_2825);
nor U9256 (N_9256,N_1777,N_1277);
nand U9257 (N_9257,N_498,N_2210);
nor U9258 (N_9258,N_5892,N_1442);
nor U9259 (N_9259,N_4363,N_5220);
nand U9260 (N_9260,N_4150,N_3429);
and U9261 (N_9261,N_3857,N_1774);
and U9262 (N_9262,N_5680,N_5503);
nor U9263 (N_9263,N_2022,N_4852);
or U9264 (N_9264,N_4198,N_3340);
and U9265 (N_9265,N_1439,N_3083);
or U9266 (N_9266,N_937,N_2396);
xor U9267 (N_9267,N_4991,N_1696);
nor U9268 (N_9268,N_1673,N_2738);
xnor U9269 (N_9269,N_5036,N_315);
nor U9270 (N_9270,N_3842,N_5945);
nor U9271 (N_9271,N_41,N_4028);
nor U9272 (N_9272,N_390,N_288);
nor U9273 (N_9273,N_5844,N_625);
and U9274 (N_9274,N_2773,N_752);
or U9275 (N_9275,N_2859,N_473);
or U9276 (N_9276,N_2675,N_3490);
or U9277 (N_9277,N_176,N_1974);
nand U9278 (N_9278,N_2520,N_1650);
and U9279 (N_9279,N_5475,N_136);
or U9280 (N_9280,N_4541,N_1352);
nand U9281 (N_9281,N_1524,N_5161);
nand U9282 (N_9282,N_5942,N_2801);
nor U9283 (N_9283,N_1055,N_4446);
or U9284 (N_9284,N_4866,N_692);
nand U9285 (N_9285,N_2496,N_5183);
nand U9286 (N_9286,N_4812,N_666);
and U9287 (N_9287,N_5873,N_646);
nor U9288 (N_9288,N_5423,N_315);
nand U9289 (N_9289,N_2702,N_3210);
or U9290 (N_9290,N_3902,N_1559);
or U9291 (N_9291,N_4786,N_3701);
and U9292 (N_9292,N_1373,N_174);
or U9293 (N_9293,N_1594,N_470);
nor U9294 (N_9294,N_2487,N_3013);
nand U9295 (N_9295,N_2749,N_706);
or U9296 (N_9296,N_455,N_1393);
or U9297 (N_9297,N_5732,N_4352);
nand U9298 (N_9298,N_77,N_331);
nor U9299 (N_9299,N_3904,N_5330);
xor U9300 (N_9300,N_5587,N_4688);
or U9301 (N_9301,N_1136,N_586);
or U9302 (N_9302,N_4217,N_4671);
or U9303 (N_9303,N_5356,N_2871);
and U9304 (N_9304,N_4447,N_1694);
and U9305 (N_9305,N_1830,N_1972);
and U9306 (N_9306,N_4420,N_4514);
xor U9307 (N_9307,N_3054,N_3008);
nor U9308 (N_9308,N_5082,N_5573);
nor U9309 (N_9309,N_508,N_324);
or U9310 (N_9310,N_878,N_844);
or U9311 (N_9311,N_4793,N_634);
xnor U9312 (N_9312,N_166,N_4767);
nor U9313 (N_9313,N_4323,N_4752);
or U9314 (N_9314,N_4958,N_2604);
nor U9315 (N_9315,N_2175,N_3363);
nor U9316 (N_9316,N_459,N_1984);
nand U9317 (N_9317,N_3548,N_270);
nand U9318 (N_9318,N_2682,N_1032);
nor U9319 (N_9319,N_3730,N_2751);
nor U9320 (N_9320,N_5970,N_4660);
nand U9321 (N_9321,N_4447,N_1419);
nand U9322 (N_9322,N_5211,N_5660);
and U9323 (N_9323,N_2683,N_1795);
or U9324 (N_9324,N_1024,N_647);
or U9325 (N_9325,N_4231,N_4247);
nand U9326 (N_9326,N_289,N_4717);
nand U9327 (N_9327,N_4514,N_3088);
nand U9328 (N_9328,N_1477,N_4602);
nor U9329 (N_9329,N_3905,N_4432);
nand U9330 (N_9330,N_3728,N_1925);
nand U9331 (N_9331,N_2695,N_3288);
xnor U9332 (N_9332,N_3264,N_2215);
nand U9333 (N_9333,N_5558,N_2922);
xor U9334 (N_9334,N_2090,N_598);
or U9335 (N_9335,N_5996,N_1067);
nand U9336 (N_9336,N_4704,N_1653);
and U9337 (N_9337,N_5193,N_900);
xor U9338 (N_9338,N_5855,N_660);
nor U9339 (N_9339,N_1281,N_2363);
xor U9340 (N_9340,N_2182,N_2216);
nand U9341 (N_9341,N_1490,N_919);
nand U9342 (N_9342,N_2321,N_173);
and U9343 (N_9343,N_4526,N_4767);
or U9344 (N_9344,N_3980,N_2040);
nor U9345 (N_9345,N_2423,N_5635);
nand U9346 (N_9346,N_1802,N_211);
nor U9347 (N_9347,N_5338,N_5618);
nor U9348 (N_9348,N_4054,N_851);
xnor U9349 (N_9349,N_5386,N_4772);
or U9350 (N_9350,N_3520,N_516);
or U9351 (N_9351,N_3137,N_5808);
nand U9352 (N_9352,N_3575,N_4955);
and U9353 (N_9353,N_4395,N_3499);
xnor U9354 (N_9354,N_1235,N_2219);
nand U9355 (N_9355,N_5447,N_887);
and U9356 (N_9356,N_245,N_4487);
or U9357 (N_9357,N_2534,N_5426);
nor U9358 (N_9358,N_5528,N_1017);
xor U9359 (N_9359,N_756,N_5808);
nand U9360 (N_9360,N_4480,N_186);
or U9361 (N_9361,N_5449,N_1526);
or U9362 (N_9362,N_4527,N_359);
nand U9363 (N_9363,N_2966,N_202);
nor U9364 (N_9364,N_3868,N_5449);
or U9365 (N_9365,N_2364,N_1152);
nand U9366 (N_9366,N_5823,N_3046);
or U9367 (N_9367,N_5652,N_1341);
or U9368 (N_9368,N_3987,N_1877);
and U9369 (N_9369,N_360,N_166);
and U9370 (N_9370,N_5085,N_4173);
nand U9371 (N_9371,N_1130,N_1783);
or U9372 (N_9372,N_4844,N_5528);
nor U9373 (N_9373,N_1471,N_4653);
or U9374 (N_9374,N_857,N_5014);
nor U9375 (N_9375,N_2225,N_640);
or U9376 (N_9376,N_1016,N_5264);
or U9377 (N_9377,N_795,N_3393);
or U9378 (N_9378,N_2645,N_1513);
nor U9379 (N_9379,N_678,N_4471);
xor U9380 (N_9380,N_2491,N_1062);
and U9381 (N_9381,N_821,N_5741);
and U9382 (N_9382,N_3864,N_4128);
nand U9383 (N_9383,N_2713,N_2201);
xor U9384 (N_9384,N_5166,N_3818);
nand U9385 (N_9385,N_1496,N_463);
or U9386 (N_9386,N_5390,N_2331);
and U9387 (N_9387,N_2150,N_3458);
nor U9388 (N_9388,N_3687,N_5380);
or U9389 (N_9389,N_5834,N_4284);
nor U9390 (N_9390,N_353,N_201);
or U9391 (N_9391,N_2763,N_4220);
nor U9392 (N_9392,N_336,N_3536);
nand U9393 (N_9393,N_4142,N_1377);
nor U9394 (N_9394,N_3561,N_1352);
nor U9395 (N_9395,N_4674,N_3658);
and U9396 (N_9396,N_5939,N_4270);
or U9397 (N_9397,N_5381,N_5205);
or U9398 (N_9398,N_4447,N_1114);
and U9399 (N_9399,N_620,N_2783);
or U9400 (N_9400,N_5491,N_545);
nand U9401 (N_9401,N_2665,N_348);
nor U9402 (N_9402,N_1507,N_2524);
nor U9403 (N_9403,N_3779,N_5841);
nor U9404 (N_9404,N_4350,N_5189);
nor U9405 (N_9405,N_4699,N_2585);
and U9406 (N_9406,N_2581,N_4371);
nand U9407 (N_9407,N_4301,N_856);
xnor U9408 (N_9408,N_9,N_2612);
and U9409 (N_9409,N_1839,N_142);
or U9410 (N_9410,N_4890,N_446);
nor U9411 (N_9411,N_4234,N_5951);
or U9412 (N_9412,N_2680,N_923);
or U9413 (N_9413,N_1638,N_1306);
or U9414 (N_9414,N_2642,N_3902);
nand U9415 (N_9415,N_5557,N_4485);
nand U9416 (N_9416,N_4625,N_4585);
or U9417 (N_9417,N_1564,N_4810);
and U9418 (N_9418,N_2059,N_3775);
nand U9419 (N_9419,N_3292,N_2915);
nand U9420 (N_9420,N_1616,N_597);
and U9421 (N_9421,N_2071,N_1591);
xnor U9422 (N_9422,N_2706,N_535);
and U9423 (N_9423,N_4705,N_4976);
nand U9424 (N_9424,N_5551,N_2118);
or U9425 (N_9425,N_5699,N_3855);
nand U9426 (N_9426,N_2625,N_693);
nand U9427 (N_9427,N_4135,N_469);
and U9428 (N_9428,N_2081,N_909);
nand U9429 (N_9429,N_1592,N_2183);
or U9430 (N_9430,N_3784,N_1517);
or U9431 (N_9431,N_143,N_5871);
and U9432 (N_9432,N_3264,N_3790);
nor U9433 (N_9433,N_5112,N_36);
and U9434 (N_9434,N_2888,N_3720);
and U9435 (N_9435,N_1147,N_3448);
nor U9436 (N_9436,N_1668,N_104);
nor U9437 (N_9437,N_2475,N_4416);
nor U9438 (N_9438,N_2150,N_1207);
nor U9439 (N_9439,N_558,N_1376);
nor U9440 (N_9440,N_3009,N_587);
nor U9441 (N_9441,N_5502,N_2863);
or U9442 (N_9442,N_1520,N_3621);
and U9443 (N_9443,N_668,N_1200);
nor U9444 (N_9444,N_790,N_4392);
nor U9445 (N_9445,N_1171,N_4556);
or U9446 (N_9446,N_5065,N_2819);
or U9447 (N_9447,N_881,N_298);
nand U9448 (N_9448,N_2441,N_5430);
and U9449 (N_9449,N_4020,N_2656);
xnor U9450 (N_9450,N_4872,N_2724);
nor U9451 (N_9451,N_1513,N_5512);
nand U9452 (N_9452,N_3704,N_5975);
and U9453 (N_9453,N_2421,N_397);
or U9454 (N_9454,N_2606,N_1012);
nor U9455 (N_9455,N_2914,N_85);
or U9456 (N_9456,N_4223,N_3702);
nand U9457 (N_9457,N_4654,N_5094);
nor U9458 (N_9458,N_4929,N_900);
nand U9459 (N_9459,N_1396,N_2966);
nand U9460 (N_9460,N_5114,N_1474);
or U9461 (N_9461,N_3269,N_5920);
or U9462 (N_9462,N_5698,N_3563);
nor U9463 (N_9463,N_5528,N_2476);
and U9464 (N_9464,N_4287,N_2337);
nand U9465 (N_9465,N_3759,N_4683);
and U9466 (N_9466,N_4117,N_3208);
and U9467 (N_9467,N_5588,N_5886);
or U9468 (N_9468,N_4919,N_1964);
and U9469 (N_9469,N_1719,N_2011);
nor U9470 (N_9470,N_995,N_2676);
nor U9471 (N_9471,N_4354,N_3765);
nor U9472 (N_9472,N_952,N_3971);
and U9473 (N_9473,N_3319,N_3579);
or U9474 (N_9474,N_856,N_5468);
or U9475 (N_9475,N_3862,N_1953);
or U9476 (N_9476,N_5012,N_5176);
xnor U9477 (N_9477,N_5287,N_3777);
and U9478 (N_9478,N_4434,N_4636);
or U9479 (N_9479,N_4971,N_3678);
and U9480 (N_9480,N_2587,N_519);
or U9481 (N_9481,N_1394,N_5863);
nor U9482 (N_9482,N_3816,N_4071);
nor U9483 (N_9483,N_3293,N_3150);
nor U9484 (N_9484,N_1114,N_4256);
nor U9485 (N_9485,N_5504,N_1548);
xor U9486 (N_9486,N_295,N_573);
nand U9487 (N_9487,N_1096,N_1429);
nor U9488 (N_9488,N_1084,N_5491);
nand U9489 (N_9489,N_2752,N_2559);
nor U9490 (N_9490,N_2132,N_1241);
or U9491 (N_9491,N_1592,N_3384);
xnor U9492 (N_9492,N_5539,N_1417);
or U9493 (N_9493,N_5866,N_5852);
nand U9494 (N_9494,N_4280,N_3076);
and U9495 (N_9495,N_558,N_1735);
nor U9496 (N_9496,N_4197,N_5007);
or U9497 (N_9497,N_3082,N_5165);
and U9498 (N_9498,N_2296,N_3323);
nand U9499 (N_9499,N_5749,N_2853);
nor U9500 (N_9500,N_2329,N_5069);
nand U9501 (N_9501,N_2835,N_4575);
nor U9502 (N_9502,N_1767,N_920);
nor U9503 (N_9503,N_4263,N_80);
nand U9504 (N_9504,N_4397,N_5276);
or U9505 (N_9505,N_3453,N_5227);
and U9506 (N_9506,N_1051,N_1794);
nor U9507 (N_9507,N_3923,N_3035);
nand U9508 (N_9508,N_5862,N_995);
nand U9509 (N_9509,N_3988,N_3469);
or U9510 (N_9510,N_4587,N_5844);
and U9511 (N_9511,N_617,N_2422);
or U9512 (N_9512,N_5938,N_2252);
and U9513 (N_9513,N_5417,N_3112);
or U9514 (N_9514,N_4582,N_4012);
nor U9515 (N_9515,N_2913,N_4298);
xor U9516 (N_9516,N_5791,N_1463);
nand U9517 (N_9517,N_2785,N_2805);
nand U9518 (N_9518,N_1126,N_4773);
or U9519 (N_9519,N_27,N_1063);
nor U9520 (N_9520,N_969,N_1152);
and U9521 (N_9521,N_2654,N_264);
or U9522 (N_9522,N_1988,N_1414);
and U9523 (N_9523,N_5771,N_807);
and U9524 (N_9524,N_3836,N_281);
nand U9525 (N_9525,N_827,N_603);
and U9526 (N_9526,N_669,N_4394);
nor U9527 (N_9527,N_4666,N_339);
or U9528 (N_9528,N_711,N_5694);
or U9529 (N_9529,N_2333,N_1644);
and U9530 (N_9530,N_1248,N_5924);
nand U9531 (N_9531,N_3440,N_672);
or U9532 (N_9532,N_5869,N_4512);
nor U9533 (N_9533,N_1815,N_4381);
or U9534 (N_9534,N_1020,N_2909);
and U9535 (N_9535,N_490,N_4437);
and U9536 (N_9536,N_5423,N_2328);
nand U9537 (N_9537,N_4026,N_5762);
nor U9538 (N_9538,N_5521,N_220);
or U9539 (N_9539,N_897,N_4459);
nand U9540 (N_9540,N_3197,N_4272);
and U9541 (N_9541,N_300,N_3485);
nor U9542 (N_9542,N_1140,N_51);
nor U9543 (N_9543,N_867,N_4730);
nand U9544 (N_9544,N_267,N_4928);
xor U9545 (N_9545,N_2056,N_5153);
nor U9546 (N_9546,N_3587,N_4466);
or U9547 (N_9547,N_4255,N_3339);
nor U9548 (N_9548,N_1054,N_5595);
nand U9549 (N_9549,N_4108,N_2196);
nand U9550 (N_9550,N_2469,N_4944);
xor U9551 (N_9551,N_1942,N_2916);
nand U9552 (N_9552,N_3008,N_3298);
and U9553 (N_9553,N_2260,N_2632);
or U9554 (N_9554,N_861,N_2050);
nand U9555 (N_9555,N_909,N_4304);
or U9556 (N_9556,N_390,N_1079);
nor U9557 (N_9557,N_770,N_1235);
and U9558 (N_9558,N_3121,N_3725);
and U9559 (N_9559,N_4028,N_3254);
nand U9560 (N_9560,N_2409,N_3397);
or U9561 (N_9561,N_5952,N_3427);
and U9562 (N_9562,N_1147,N_1366);
or U9563 (N_9563,N_4670,N_5045);
and U9564 (N_9564,N_1849,N_5378);
nor U9565 (N_9565,N_5373,N_1393);
and U9566 (N_9566,N_704,N_1176);
nor U9567 (N_9567,N_3632,N_4949);
nor U9568 (N_9568,N_1407,N_4254);
and U9569 (N_9569,N_3579,N_4461);
xnor U9570 (N_9570,N_2520,N_546);
and U9571 (N_9571,N_545,N_3192);
or U9572 (N_9572,N_5898,N_1814);
nor U9573 (N_9573,N_3972,N_4200);
or U9574 (N_9574,N_18,N_1955);
nor U9575 (N_9575,N_5297,N_1900);
nor U9576 (N_9576,N_1469,N_4974);
and U9577 (N_9577,N_175,N_4962);
nor U9578 (N_9578,N_4067,N_5001);
nor U9579 (N_9579,N_2124,N_4346);
nor U9580 (N_9580,N_4452,N_3208);
nor U9581 (N_9581,N_1480,N_4534);
nor U9582 (N_9582,N_131,N_597);
nand U9583 (N_9583,N_3600,N_3312);
and U9584 (N_9584,N_1084,N_5810);
xnor U9585 (N_9585,N_3737,N_5300);
nor U9586 (N_9586,N_2200,N_5287);
nor U9587 (N_9587,N_4700,N_2715);
and U9588 (N_9588,N_5119,N_5116);
or U9589 (N_9589,N_2287,N_4751);
and U9590 (N_9590,N_2999,N_2631);
nand U9591 (N_9591,N_2808,N_5632);
nor U9592 (N_9592,N_487,N_550);
xnor U9593 (N_9593,N_446,N_664);
nand U9594 (N_9594,N_2717,N_1973);
or U9595 (N_9595,N_632,N_5835);
and U9596 (N_9596,N_3573,N_2188);
and U9597 (N_9597,N_4370,N_4449);
xnor U9598 (N_9598,N_5257,N_761);
or U9599 (N_9599,N_4101,N_1249);
nor U9600 (N_9600,N_2279,N_4829);
and U9601 (N_9601,N_5120,N_3393);
and U9602 (N_9602,N_607,N_555);
nor U9603 (N_9603,N_2781,N_2958);
and U9604 (N_9604,N_5550,N_4869);
and U9605 (N_9605,N_5610,N_4973);
and U9606 (N_9606,N_4802,N_51);
or U9607 (N_9607,N_3106,N_2988);
or U9608 (N_9608,N_2647,N_4268);
or U9609 (N_9609,N_4152,N_3380);
or U9610 (N_9610,N_2474,N_5455);
nand U9611 (N_9611,N_3483,N_3894);
or U9612 (N_9612,N_5423,N_5246);
nor U9613 (N_9613,N_4088,N_4578);
or U9614 (N_9614,N_1459,N_5491);
or U9615 (N_9615,N_1088,N_5211);
and U9616 (N_9616,N_2899,N_942);
nor U9617 (N_9617,N_4204,N_5529);
nor U9618 (N_9618,N_5141,N_1546);
nand U9619 (N_9619,N_1432,N_158);
or U9620 (N_9620,N_5165,N_383);
nor U9621 (N_9621,N_474,N_5820);
nor U9622 (N_9622,N_1236,N_2364);
xor U9623 (N_9623,N_4240,N_5240);
and U9624 (N_9624,N_2371,N_3229);
or U9625 (N_9625,N_4234,N_3546);
and U9626 (N_9626,N_4193,N_1559);
or U9627 (N_9627,N_3485,N_2852);
nor U9628 (N_9628,N_20,N_5952);
nor U9629 (N_9629,N_4077,N_1983);
nand U9630 (N_9630,N_4922,N_4034);
and U9631 (N_9631,N_4818,N_5335);
nor U9632 (N_9632,N_92,N_565);
nor U9633 (N_9633,N_3722,N_182);
nand U9634 (N_9634,N_1327,N_2933);
or U9635 (N_9635,N_2139,N_3263);
or U9636 (N_9636,N_738,N_2462);
and U9637 (N_9637,N_486,N_3671);
nand U9638 (N_9638,N_3648,N_4087);
nand U9639 (N_9639,N_2130,N_3912);
xnor U9640 (N_9640,N_3302,N_3100);
nor U9641 (N_9641,N_5529,N_1178);
xor U9642 (N_9642,N_5845,N_498);
nor U9643 (N_9643,N_4331,N_5876);
nand U9644 (N_9644,N_1627,N_2295);
and U9645 (N_9645,N_3852,N_3023);
nor U9646 (N_9646,N_3326,N_4385);
or U9647 (N_9647,N_33,N_1567);
or U9648 (N_9648,N_1260,N_3589);
xnor U9649 (N_9649,N_2360,N_3154);
nand U9650 (N_9650,N_4502,N_3575);
nand U9651 (N_9651,N_2025,N_632);
nand U9652 (N_9652,N_4162,N_1111);
and U9653 (N_9653,N_4098,N_5176);
nor U9654 (N_9654,N_4766,N_4873);
nand U9655 (N_9655,N_1581,N_5654);
nand U9656 (N_9656,N_4806,N_5669);
and U9657 (N_9657,N_1031,N_4811);
nor U9658 (N_9658,N_1981,N_1949);
and U9659 (N_9659,N_2558,N_3488);
nand U9660 (N_9660,N_4008,N_5060);
nand U9661 (N_9661,N_4331,N_531);
nor U9662 (N_9662,N_2426,N_366);
or U9663 (N_9663,N_5982,N_853);
nor U9664 (N_9664,N_162,N_381);
nand U9665 (N_9665,N_4525,N_2175);
or U9666 (N_9666,N_4810,N_862);
xnor U9667 (N_9667,N_5053,N_5397);
nor U9668 (N_9668,N_4240,N_4064);
and U9669 (N_9669,N_1962,N_311);
nor U9670 (N_9670,N_5537,N_4042);
and U9671 (N_9671,N_2582,N_4189);
or U9672 (N_9672,N_2935,N_303);
xor U9673 (N_9673,N_2178,N_1735);
nor U9674 (N_9674,N_3181,N_4711);
nor U9675 (N_9675,N_3291,N_5708);
nand U9676 (N_9676,N_2432,N_2845);
nor U9677 (N_9677,N_4221,N_3262);
and U9678 (N_9678,N_550,N_1403);
nand U9679 (N_9679,N_727,N_974);
and U9680 (N_9680,N_5734,N_1278);
nor U9681 (N_9681,N_3620,N_2173);
or U9682 (N_9682,N_1866,N_2648);
and U9683 (N_9683,N_5055,N_5850);
and U9684 (N_9684,N_1616,N_2499);
nand U9685 (N_9685,N_21,N_2876);
or U9686 (N_9686,N_5290,N_3041);
or U9687 (N_9687,N_438,N_5148);
xor U9688 (N_9688,N_882,N_5756);
nand U9689 (N_9689,N_2869,N_4131);
and U9690 (N_9690,N_4558,N_1758);
nand U9691 (N_9691,N_518,N_2474);
nand U9692 (N_9692,N_1796,N_783);
or U9693 (N_9693,N_5398,N_927);
nor U9694 (N_9694,N_3256,N_2295);
and U9695 (N_9695,N_4479,N_3174);
xnor U9696 (N_9696,N_1681,N_2399);
or U9697 (N_9697,N_3632,N_3956);
or U9698 (N_9698,N_4711,N_3600);
xor U9699 (N_9699,N_4908,N_5664);
nor U9700 (N_9700,N_4097,N_311);
nand U9701 (N_9701,N_2607,N_3377);
or U9702 (N_9702,N_3332,N_3137);
nor U9703 (N_9703,N_3473,N_649);
nand U9704 (N_9704,N_1454,N_4152);
nand U9705 (N_9705,N_1926,N_2651);
and U9706 (N_9706,N_770,N_1086);
and U9707 (N_9707,N_1827,N_1986);
and U9708 (N_9708,N_1601,N_205);
or U9709 (N_9709,N_1959,N_5924);
nor U9710 (N_9710,N_5797,N_3820);
xor U9711 (N_9711,N_5907,N_2506);
or U9712 (N_9712,N_5504,N_3557);
and U9713 (N_9713,N_1929,N_550);
or U9714 (N_9714,N_3020,N_1322);
nor U9715 (N_9715,N_2552,N_4868);
nor U9716 (N_9716,N_3964,N_4899);
nor U9717 (N_9717,N_3151,N_1432);
or U9718 (N_9718,N_4836,N_3160);
and U9719 (N_9719,N_3672,N_4917);
nand U9720 (N_9720,N_2881,N_1042);
nor U9721 (N_9721,N_3809,N_2461);
or U9722 (N_9722,N_2678,N_907);
and U9723 (N_9723,N_4039,N_5277);
and U9724 (N_9724,N_3927,N_3062);
nor U9725 (N_9725,N_2901,N_197);
and U9726 (N_9726,N_678,N_4498);
or U9727 (N_9727,N_4346,N_5875);
or U9728 (N_9728,N_1820,N_4490);
nor U9729 (N_9729,N_2784,N_1328);
nand U9730 (N_9730,N_3969,N_2264);
nor U9731 (N_9731,N_4349,N_3977);
or U9732 (N_9732,N_1654,N_386);
or U9733 (N_9733,N_5306,N_2597);
or U9734 (N_9734,N_4304,N_1071);
or U9735 (N_9735,N_1606,N_3218);
nor U9736 (N_9736,N_1135,N_3975);
or U9737 (N_9737,N_2502,N_3496);
or U9738 (N_9738,N_4787,N_4363);
and U9739 (N_9739,N_1432,N_3495);
nand U9740 (N_9740,N_3107,N_4964);
and U9741 (N_9741,N_4868,N_5220);
or U9742 (N_9742,N_5853,N_386);
and U9743 (N_9743,N_4680,N_4263);
and U9744 (N_9744,N_2781,N_446);
nand U9745 (N_9745,N_632,N_2768);
or U9746 (N_9746,N_3308,N_707);
and U9747 (N_9747,N_4585,N_5421);
xor U9748 (N_9748,N_5455,N_5435);
nand U9749 (N_9749,N_34,N_3620);
nand U9750 (N_9750,N_5341,N_2677);
nor U9751 (N_9751,N_3283,N_3389);
and U9752 (N_9752,N_4130,N_1331);
xnor U9753 (N_9753,N_2211,N_1395);
or U9754 (N_9754,N_699,N_3067);
and U9755 (N_9755,N_3249,N_1526);
nand U9756 (N_9756,N_194,N_4999);
nor U9757 (N_9757,N_1301,N_2260);
nand U9758 (N_9758,N_5711,N_4549);
xnor U9759 (N_9759,N_1468,N_4643);
and U9760 (N_9760,N_5237,N_470);
nor U9761 (N_9761,N_2512,N_2081);
xnor U9762 (N_9762,N_4233,N_1755);
and U9763 (N_9763,N_5521,N_1702);
nor U9764 (N_9764,N_4552,N_5821);
or U9765 (N_9765,N_2990,N_2096);
or U9766 (N_9766,N_4644,N_3612);
or U9767 (N_9767,N_4295,N_348);
or U9768 (N_9768,N_1925,N_1607);
nand U9769 (N_9769,N_2325,N_3792);
nor U9770 (N_9770,N_735,N_138);
and U9771 (N_9771,N_1423,N_2919);
and U9772 (N_9772,N_333,N_1665);
nor U9773 (N_9773,N_4289,N_3065);
xnor U9774 (N_9774,N_3902,N_3735);
and U9775 (N_9775,N_468,N_4154);
and U9776 (N_9776,N_1376,N_179);
nand U9777 (N_9777,N_3615,N_1641);
nand U9778 (N_9778,N_5804,N_1713);
nor U9779 (N_9779,N_4058,N_1305);
and U9780 (N_9780,N_5240,N_790);
and U9781 (N_9781,N_1571,N_1584);
and U9782 (N_9782,N_1074,N_2542);
nor U9783 (N_9783,N_1440,N_809);
nor U9784 (N_9784,N_4356,N_493);
or U9785 (N_9785,N_4333,N_1223);
nor U9786 (N_9786,N_2000,N_3166);
nor U9787 (N_9787,N_4646,N_4651);
nand U9788 (N_9788,N_2110,N_896);
and U9789 (N_9789,N_1162,N_3229);
xnor U9790 (N_9790,N_1947,N_1377);
or U9791 (N_9791,N_2166,N_5702);
nor U9792 (N_9792,N_5555,N_2184);
nor U9793 (N_9793,N_3574,N_1436);
nand U9794 (N_9794,N_778,N_4325);
and U9795 (N_9795,N_4794,N_4137);
xnor U9796 (N_9796,N_876,N_2351);
or U9797 (N_9797,N_157,N_887);
or U9798 (N_9798,N_1285,N_169);
nand U9799 (N_9799,N_1660,N_44);
or U9800 (N_9800,N_807,N_3798);
nor U9801 (N_9801,N_3681,N_1818);
or U9802 (N_9802,N_5846,N_4832);
and U9803 (N_9803,N_3135,N_2937);
nor U9804 (N_9804,N_2544,N_5878);
nand U9805 (N_9805,N_5650,N_1457);
and U9806 (N_9806,N_1384,N_721);
or U9807 (N_9807,N_2354,N_607);
nand U9808 (N_9808,N_4458,N_3424);
nor U9809 (N_9809,N_4512,N_382);
nand U9810 (N_9810,N_5882,N_3595);
nor U9811 (N_9811,N_4471,N_5432);
or U9812 (N_9812,N_2149,N_4162);
and U9813 (N_9813,N_820,N_185);
or U9814 (N_9814,N_5276,N_2566);
and U9815 (N_9815,N_990,N_5587);
and U9816 (N_9816,N_1549,N_2683);
nand U9817 (N_9817,N_1213,N_3648);
and U9818 (N_9818,N_5355,N_1865);
nand U9819 (N_9819,N_5163,N_297);
or U9820 (N_9820,N_5948,N_3187);
and U9821 (N_9821,N_4022,N_2879);
and U9822 (N_9822,N_3138,N_4519);
nand U9823 (N_9823,N_1420,N_4349);
nand U9824 (N_9824,N_2549,N_158);
and U9825 (N_9825,N_2304,N_5785);
nand U9826 (N_9826,N_3633,N_3315);
nand U9827 (N_9827,N_5847,N_661);
or U9828 (N_9828,N_5274,N_4098);
xor U9829 (N_9829,N_598,N_5217);
nand U9830 (N_9830,N_662,N_2891);
nand U9831 (N_9831,N_2206,N_849);
and U9832 (N_9832,N_909,N_2499);
nor U9833 (N_9833,N_3022,N_647);
nand U9834 (N_9834,N_302,N_1494);
xor U9835 (N_9835,N_5814,N_3111);
nand U9836 (N_9836,N_1252,N_2730);
nor U9837 (N_9837,N_1834,N_3801);
and U9838 (N_9838,N_3937,N_3627);
nand U9839 (N_9839,N_220,N_2160);
or U9840 (N_9840,N_5975,N_40);
nor U9841 (N_9841,N_2011,N_2790);
and U9842 (N_9842,N_1522,N_923);
or U9843 (N_9843,N_4189,N_3303);
xor U9844 (N_9844,N_5630,N_5916);
or U9845 (N_9845,N_1052,N_5789);
or U9846 (N_9846,N_1914,N_3325);
and U9847 (N_9847,N_1610,N_5027);
xnor U9848 (N_9848,N_326,N_3659);
nor U9849 (N_9849,N_2755,N_91);
and U9850 (N_9850,N_4328,N_1748);
nand U9851 (N_9851,N_1178,N_1645);
or U9852 (N_9852,N_180,N_5857);
and U9853 (N_9853,N_631,N_4391);
or U9854 (N_9854,N_4687,N_849);
and U9855 (N_9855,N_1960,N_5699);
nand U9856 (N_9856,N_4611,N_3502);
nand U9857 (N_9857,N_5105,N_5935);
and U9858 (N_9858,N_4418,N_3630);
and U9859 (N_9859,N_4854,N_3009);
nand U9860 (N_9860,N_5876,N_563);
or U9861 (N_9861,N_1392,N_3723);
nand U9862 (N_9862,N_3948,N_72);
or U9863 (N_9863,N_1633,N_5497);
and U9864 (N_9864,N_2051,N_5953);
xnor U9865 (N_9865,N_782,N_2474);
and U9866 (N_9866,N_1919,N_4350);
nor U9867 (N_9867,N_1080,N_4211);
or U9868 (N_9868,N_779,N_519);
nor U9869 (N_9869,N_795,N_5433);
nand U9870 (N_9870,N_4070,N_2000);
or U9871 (N_9871,N_4794,N_5189);
nor U9872 (N_9872,N_388,N_716);
or U9873 (N_9873,N_3187,N_1678);
xnor U9874 (N_9874,N_4920,N_5128);
and U9875 (N_9875,N_3746,N_531);
and U9876 (N_9876,N_1821,N_2939);
nand U9877 (N_9877,N_4236,N_4194);
and U9878 (N_9878,N_5259,N_2246);
nor U9879 (N_9879,N_4088,N_565);
xor U9880 (N_9880,N_3531,N_3968);
or U9881 (N_9881,N_21,N_2543);
nor U9882 (N_9882,N_235,N_2378);
or U9883 (N_9883,N_276,N_2926);
nand U9884 (N_9884,N_3327,N_3093);
and U9885 (N_9885,N_429,N_4467);
nand U9886 (N_9886,N_3249,N_506);
and U9887 (N_9887,N_1655,N_101);
or U9888 (N_9888,N_1338,N_3709);
or U9889 (N_9889,N_2912,N_2773);
nand U9890 (N_9890,N_4629,N_2705);
nand U9891 (N_9891,N_3263,N_5979);
and U9892 (N_9892,N_3064,N_5843);
or U9893 (N_9893,N_1615,N_5669);
xor U9894 (N_9894,N_424,N_208);
or U9895 (N_9895,N_1040,N_1212);
xor U9896 (N_9896,N_2363,N_2480);
nand U9897 (N_9897,N_5177,N_5392);
nor U9898 (N_9898,N_3048,N_4392);
nor U9899 (N_9899,N_2308,N_849);
or U9900 (N_9900,N_1102,N_4928);
nand U9901 (N_9901,N_1226,N_1795);
nand U9902 (N_9902,N_4849,N_4966);
nor U9903 (N_9903,N_2935,N_4912);
nand U9904 (N_9904,N_2513,N_856);
and U9905 (N_9905,N_2018,N_3083);
and U9906 (N_9906,N_4237,N_1104);
nor U9907 (N_9907,N_1570,N_2909);
or U9908 (N_9908,N_510,N_4034);
xnor U9909 (N_9909,N_5623,N_4706);
or U9910 (N_9910,N_4007,N_2725);
or U9911 (N_9911,N_826,N_2431);
and U9912 (N_9912,N_4849,N_101);
and U9913 (N_9913,N_2929,N_1568);
nand U9914 (N_9914,N_2264,N_4069);
nor U9915 (N_9915,N_3569,N_1290);
or U9916 (N_9916,N_5153,N_2239);
and U9917 (N_9917,N_4701,N_4186);
or U9918 (N_9918,N_5521,N_2207);
nand U9919 (N_9919,N_5659,N_3552);
and U9920 (N_9920,N_5356,N_2870);
or U9921 (N_9921,N_2017,N_1457);
nor U9922 (N_9922,N_2911,N_1335);
or U9923 (N_9923,N_2776,N_1976);
nand U9924 (N_9924,N_754,N_2681);
nor U9925 (N_9925,N_2057,N_5304);
or U9926 (N_9926,N_3150,N_5238);
or U9927 (N_9927,N_4873,N_4353);
or U9928 (N_9928,N_4175,N_962);
and U9929 (N_9929,N_2982,N_3807);
xnor U9930 (N_9930,N_4883,N_1135);
and U9931 (N_9931,N_662,N_2856);
nor U9932 (N_9932,N_4435,N_1623);
or U9933 (N_9933,N_3448,N_374);
or U9934 (N_9934,N_3788,N_1872);
nand U9935 (N_9935,N_5525,N_1926);
or U9936 (N_9936,N_5219,N_1578);
nand U9937 (N_9937,N_4224,N_5253);
and U9938 (N_9938,N_5356,N_22);
nor U9939 (N_9939,N_2884,N_4082);
nor U9940 (N_9940,N_4002,N_3111);
or U9941 (N_9941,N_5730,N_5216);
and U9942 (N_9942,N_1528,N_4840);
nor U9943 (N_9943,N_2136,N_2185);
and U9944 (N_9944,N_131,N_5581);
or U9945 (N_9945,N_2919,N_4577);
xor U9946 (N_9946,N_3891,N_772);
nand U9947 (N_9947,N_2077,N_2407);
nand U9948 (N_9948,N_4701,N_4440);
nor U9949 (N_9949,N_671,N_3772);
or U9950 (N_9950,N_2810,N_5773);
nand U9951 (N_9951,N_3143,N_5651);
and U9952 (N_9952,N_2133,N_2175);
or U9953 (N_9953,N_1690,N_3220);
and U9954 (N_9954,N_1105,N_1664);
nand U9955 (N_9955,N_924,N_5907);
xnor U9956 (N_9956,N_1625,N_1139);
nand U9957 (N_9957,N_4370,N_4061);
and U9958 (N_9958,N_2558,N_4028);
nor U9959 (N_9959,N_3824,N_5834);
nand U9960 (N_9960,N_390,N_5617);
nand U9961 (N_9961,N_695,N_3828);
nand U9962 (N_9962,N_5526,N_1164);
xor U9963 (N_9963,N_5474,N_5208);
or U9964 (N_9964,N_1073,N_2709);
xor U9965 (N_9965,N_2840,N_4488);
or U9966 (N_9966,N_4656,N_5778);
xor U9967 (N_9967,N_2304,N_5369);
nand U9968 (N_9968,N_2250,N_4264);
nand U9969 (N_9969,N_4331,N_2347);
xnor U9970 (N_9970,N_491,N_4531);
nand U9971 (N_9971,N_4326,N_3679);
and U9972 (N_9972,N_1120,N_4999);
or U9973 (N_9973,N_3472,N_1958);
nand U9974 (N_9974,N_628,N_1128);
and U9975 (N_9975,N_3031,N_4983);
nor U9976 (N_9976,N_5263,N_244);
nand U9977 (N_9977,N_4655,N_4532);
nand U9978 (N_9978,N_2820,N_1512);
nand U9979 (N_9979,N_2319,N_1683);
or U9980 (N_9980,N_3516,N_5423);
and U9981 (N_9981,N_1650,N_2308);
xnor U9982 (N_9982,N_4450,N_2037);
nand U9983 (N_9983,N_5198,N_2457);
or U9984 (N_9984,N_2800,N_4179);
and U9985 (N_9985,N_3354,N_4507);
or U9986 (N_9986,N_4487,N_5273);
nor U9987 (N_9987,N_62,N_3982);
nand U9988 (N_9988,N_4849,N_2688);
xor U9989 (N_9989,N_2958,N_1452);
nor U9990 (N_9990,N_1077,N_839);
and U9991 (N_9991,N_570,N_4764);
xor U9992 (N_9992,N_1510,N_2742);
and U9993 (N_9993,N_168,N_5917);
nor U9994 (N_9994,N_5840,N_3306);
xor U9995 (N_9995,N_1257,N_1741);
nor U9996 (N_9996,N_908,N_677);
nor U9997 (N_9997,N_3473,N_2997);
or U9998 (N_9998,N_2059,N_5759);
xnor U9999 (N_9999,N_4751,N_4409);
and U10000 (N_10000,N_3912,N_2709);
nor U10001 (N_10001,N_4856,N_5190);
nor U10002 (N_10002,N_666,N_5884);
or U10003 (N_10003,N_2646,N_3865);
and U10004 (N_10004,N_3529,N_4041);
nor U10005 (N_10005,N_5629,N_2116);
and U10006 (N_10006,N_592,N_4757);
nor U10007 (N_10007,N_338,N_1353);
and U10008 (N_10008,N_5755,N_4159);
nor U10009 (N_10009,N_1335,N_5982);
or U10010 (N_10010,N_271,N_4711);
nor U10011 (N_10011,N_543,N_3094);
nor U10012 (N_10012,N_1841,N_4892);
or U10013 (N_10013,N_69,N_5747);
nor U10014 (N_10014,N_2001,N_1752);
and U10015 (N_10015,N_5440,N_23);
or U10016 (N_10016,N_4947,N_521);
nand U10017 (N_10017,N_3371,N_2068);
or U10018 (N_10018,N_2302,N_1609);
or U10019 (N_10019,N_906,N_5530);
and U10020 (N_10020,N_264,N_5480);
nand U10021 (N_10021,N_316,N_2819);
nand U10022 (N_10022,N_3513,N_534);
or U10023 (N_10023,N_5016,N_4385);
or U10024 (N_10024,N_3307,N_1739);
or U10025 (N_10025,N_1647,N_5470);
nand U10026 (N_10026,N_202,N_1823);
and U10027 (N_10027,N_4464,N_3489);
nor U10028 (N_10028,N_4537,N_5107);
and U10029 (N_10029,N_3201,N_3795);
nor U10030 (N_10030,N_3217,N_5202);
or U10031 (N_10031,N_1966,N_2024);
nand U10032 (N_10032,N_4716,N_395);
xnor U10033 (N_10033,N_5285,N_1122);
or U10034 (N_10034,N_2878,N_3878);
nor U10035 (N_10035,N_4847,N_1494);
and U10036 (N_10036,N_3644,N_1425);
and U10037 (N_10037,N_4699,N_544);
or U10038 (N_10038,N_2421,N_5964);
or U10039 (N_10039,N_2547,N_5049);
nand U10040 (N_10040,N_3248,N_1206);
xor U10041 (N_10041,N_3384,N_5610);
or U10042 (N_10042,N_67,N_2127);
and U10043 (N_10043,N_3094,N_4825);
or U10044 (N_10044,N_405,N_567);
nor U10045 (N_10045,N_4628,N_639);
nand U10046 (N_10046,N_262,N_4533);
and U10047 (N_10047,N_2299,N_3034);
nand U10048 (N_10048,N_4228,N_5740);
or U10049 (N_10049,N_4380,N_2880);
xor U10050 (N_10050,N_1810,N_1081);
and U10051 (N_10051,N_765,N_5658);
nor U10052 (N_10052,N_1474,N_3545);
nand U10053 (N_10053,N_5368,N_5406);
nor U10054 (N_10054,N_4533,N_2898);
nor U10055 (N_10055,N_5703,N_664);
nor U10056 (N_10056,N_2386,N_5154);
nor U10057 (N_10057,N_606,N_5017);
or U10058 (N_10058,N_641,N_284);
nor U10059 (N_10059,N_467,N_231);
xnor U10060 (N_10060,N_3257,N_1663);
xor U10061 (N_10061,N_958,N_4090);
xor U10062 (N_10062,N_3276,N_5315);
nor U10063 (N_10063,N_4965,N_1876);
nand U10064 (N_10064,N_114,N_2564);
nand U10065 (N_10065,N_5445,N_2242);
or U10066 (N_10066,N_4060,N_5556);
and U10067 (N_10067,N_4915,N_4637);
nand U10068 (N_10068,N_4155,N_3216);
nand U10069 (N_10069,N_2485,N_4518);
and U10070 (N_10070,N_5721,N_5254);
or U10071 (N_10071,N_4465,N_1288);
or U10072 (N_10072,N_5564,N_4835);
nand U10073 (N_10073,N_947,N_3388);
nand U10074 (N_10074,N_4777,N_4922);
and U10075 (N_10075,N_3933,N_3034);
nand U10076 (N_10076,N_5344,N_5894);
or U10077 (N_10077,N_5355,N_4619);
nand U10078 (N_10078,N_5784,N_3378);
and U10079 (N_10079,N_4532,N_5056);
nand U10080 (N_10080,N_4981,N_5960);
or U10081 (N_10081,N_2031,N_2884);
and U10082 (N_10082,N_224,N_1531);
nor U10083 (N_10083,N_5354,N_5824);
or U10084 (N_10084,N_299,N_1235);
or U10085 (N_10085,N_2822,N_3525);
nand U10086 (N_10086,N_4058,N_3230);
and U10087 (N_10087,N_56,N_173);
or U10088 (N_10088,N_5131,N_5159);
and U10089 (N_10089,N_564,N_605);
and U10090 (N_10090,N_4828,N_2723);
or U10091 (N_10091,N_2094,N_3432);
and U10092 (N_10092,N_1714,N_4095);
or U10093 (N_10093,N_3718,N_1959);
or U10094 (N_10094,N_1483,N_4126);
nand U10095 (N_10095,N_451,N_3640);
nor U10096 (N_10096,N_5146,N_5319);
nor U10097 (N_10097,N_5251,N_1002);
and U10098 (N_10098,N_3703,N_2619);
nor U10099 (N_10099,N_5384,N_4626);
nor U10100 (N_10100,N_1710,N_1223);
and U10101 (N_10101,N_733,N_2238);
or U10102 (N_10102,N_4653,N_2358);
xnor U10103 (N_10103,N_1505,N_4802);
and U10104 (N_10104,N_2344,N_3410);
or U10105 (N_10105,N_3867,N_3032);
nor U10106 (N_10106,N_2307,N_2404);
nand U10107 (N_10107,N_2493,N_1582);
nor U10108 (N_10108,N_231,N_3251);
and U10109 (N_10109,N_5332,N_683);
xnor U10110 (N_10110,N_5514,N_3017);
and U10111 (N_10111,N_1560,N_829);
or U10112 (N_10112,N_236,N_1158);
nand U10113 (N_10113,N_1385,N_2369);
nand U10114 (N_10114,N_5749,N_2916);
xnor U10115 (N_10115,N_4601,N_1736);
nor U10116 (N_10116,N_4600,N_2431);
nor U10117 (N_10117,N_4423,N_3372);
and U10118 (N_10118,N_373,N_5354);
or U10119 (N_10119,N_605,N_1751);
or U10120 (N_10120,N_1459,N_3750);
and U10121 (N_10121,N_590,N_3806);
nand U10122 (N_10122,N_2910,N_4826);
or U10123 (N_10123,N_5822,N_4240);
or U10124 (N_10124,N_4582,N_2342);
nor U10125 (N_10125,N_3183,N_3381);
nand U10126 (N_10126,N_5858,N_3106);
and U10127 (N_10127,N_754,N_5698);
nor U10128 (N_10128,N_2960,N_2254);
or U10129 (N_10129,N_2681,N_1482);
or U10130 (N_10130,N_2707,N_2652);
nor U10131 (N_10131,N_370,N_2184);
and U10132 (N_10132,N_1966,N_5153);
nand U10133 (N_10133,N_3683,N_3020);
or U10134 (N_10134,N_5823,N_4220);
and U10135 (N_10135,N_5751,N_4776);
and U10136 (N_10136,N_118,N_1956);
or U10137 (N_10137,N_676,N_3413);
nand U10138 (N_10138,N_3360,N_4921);
or U10139 (N_10139,N_630,N_4897);
or U10140 (N_10140,N_182,N_4468);
nor U10141 (N_10141,N_1308,N_1764);
and U10142 (N_10142,N_812,N_5553);
or U10143 (N_10143,N_5725,N_4437);
or U10144 (N_10144,N_320,N_1715);
or U10145 (N_10145,N_4607,N_1493);
nand U10146 (N_10146,N_4855,N_4101);
or U10147 (N_10147,N_5180,N_3687);
xor U10148 (N_10148,N_3089,N_3516);
nor U10149 (N_10149,N_894,N_3084);
nor U10150 (N_10150,N_431,N_287);
nand U10151 (N_10151,N_2729,N_2159);
nor U10152 (N_10152,N_2203,N_5358);
nor U10153 (N_10153,N_1392,N_3731);
nor U10154 (N_10154,N_4053,N_364);
or U10155 (N_10155,N_2517,N_2595);
nor U10156 (N_10156,N_2492,N_4023);
xor U10157 (N_10157,N_1873,N_491);
or U10158 (N_10158,N_1724,N_4147);
nand U10159 (N_10159,N_373,N_4359);
and U10160 (N_10160,N_484,N_4566);
nand U10161 (N_10161,N_4084,N_677);
nand U10162 (N_10162,N_842,N_818);
nor U10163 (N_10163,N_2139,N_3640);
or U10164 (N_10164,N_2210,N_1682);
and U10165 (N_10165,N_4041,N_1517);
nor U10166 (N_10166,N_2790,N_1706);
nand U10167 (N_10167,N_3165,N_92);
nand U10168 (N_10168,N_5699,N_2041);
or U10169 (N_10169,N_4028,N_3516);
nand U10170 (N_10170,N_2535,N_3302);
and U10171 (N_10171,N_5201,N_1126);
nor U10172 (N_10172,N_2619,N_3247);
nor U10173 (N_10173,N_5796,N_1072);
nor U10174 (N_10174,N_2805,N_3092);
and U10175 (N_10175,N_5901,N_4782);
nor U10176 (N_10176,N_5444,N_3247);
and U10177 (N_10177,N_1118,N_3029);
and U10178 (N_10178,N_4160,N_444);
and U10179 (N_10179,N_4679,N_4636);
nor U10180 (N_10180,N_4512,N_5317);
nor U10181 (N_10181,N_4364,N_154);
and U10182 (N_10182,N_4727,N_1481);
nand U10183 (N_10183,N_2734,N_3060);
nand U10184 (N_10184,N_3531,N_2116);
or U10185 (N_10185,N_4680,N_2985);
nor U10186 (N_10186,N_3739,N_2453);
xnor U10187 (N_10187,N_1342,N_4914);
and U10188 (N_10188,N_2239,N_5640);
and U10189 (N_10189,N_5582,N_4424);
nand U10190 (N_10190,N_3895,N_3848);
or U10191 (N_10191,N_4008,N_4796);
nand U10192 (N_10192,N_4863,N_5156);
or U10193 (N_10193,N_3780,N_1414);
or U10194 (N_10194,N_1255,N_1157);
nor U10195 (N_10195,N_5676,N_2689);
nor U10196 (N_10196,N_5209,N_4708);
xor U10197 (N_10197,N_2211,N_3016);
nor U10198 (N_10198,N_3518,N_5229);
and U10199 (N_10199,N_5724,N_3012);
xnor U10200 (N_10200,N_2809,N_3500);
and U10201 (N_10201,N_42,N_1218);
nor U10202 (N_10202,N_5250,N_5087);
nor U10203 (N_10203,N_811,N_3990);
nor U10204 (N_10204,N_5562,N_1970);
nor U10205 (N_10205,N_1991,N_2452);
and U10206 (N_10206,N_1537,N_4086);
nand U10207 (N_10207,N_291,N_1621);
nand U10208 (N_10208,N_5465,N_1516);
nand U10209 (N_10209,N_2762,N_2204);
nand U10210 (N_10210,N_434,N_2469);
nand U10211 (N_10211,N_4172,N_5231);
nand U10212 (N_10212,N_267,N_4425);
nand U10213 (N_10213,N_2894,N_1939);
nor U10214 (N_10214,N_1020,N_189);
nand U10215 (N_10215,N_5930,N_5056);
and U10216 (N_10216,N_1743,N_729);
or U10217 (N_10217,N_5410,N_2056);
xor U10218 (N_10218,N_5802,N_428);
nand U10219 (N_10219,N_790,N_2142);
nor U10220 (N_10220,N_2370,N_1257);
nand U10221 (N_10221,N_2264,N_2471);
xnor U10222 (N_10222,N_5233,N_3338);
and U10223 (N_10223,N_2197,N_2136);
or U10224 (N_10224,N_5853,N_2626);
nand U10225 (N_10225,N_1977,N_3999);
or U10226 (N_10226,N_1598,N_5253);
or U10227 (N_10227,N_5075,N_4691);
nand U10228 (N_10228,N_1635,N_2386);
xnor U10229 (N_10229,N_22,N_5283);
nand U10230 (N_10230,N_1261,N_5088);
nand U10231 (N_10231,N_986,N_2685);
and U10232 (N_10232,N_2823,N_1801);
nor U10233 (N_10233,N_5927,N_3920);
xor U10234 (N_10234,N_5582,N_5160);
and U10235 (N_10235,N_3021,N_5894);
nor U10236 (N_10236,N_3972,N_4114);
or U10237 (N_10237,N_2061,N_3170);
and U10238 (N_10238,N_3253,N_5491);
nand U10239 (N_10239,N_1116,N_3680);
and U10240 (N_10240,N_2112,N_2581);
or U10241 (N_10241,N_4339,N_5864);
and U10242 (N_10242,N_3749,N_753);
and U10243 (N_10243,N_4300,N_223);
and U10244 (N_10244,N_1358,N_2198);
or U10245 (N_10245,N_4048,N_1980);
nor U10246 (N_10246,N_2464,N_156);
or U10247 (N_10247,N_804,N_1466);
nor U10248 (N_10248,N_1052,N_3719);
nor U10249 (N_10249,N_3404,N_5452);
nor U10250 (N_10250,N_235,N_4037);
or U10251 (N_10251,N_3420,N_3565);
and U10252 (N_10252,N_656,N_3894);
and U10253 (N_10253,N_5694,N_3817);
nand U10254 (N_10254,N_4949,N_1811);
nor U10255 (N_10255,N_4012,N_38);
and U10256 (N_10256,N_105,N_4776);
or U10257 (N_10257,N_1757,N_5753);
and U10258 (N_10258,N_4939,N_4761);
nor U10259 (N_10259,N_229,N_1973);
and U10260 (N_10260,N_5975,N_2221);
nand U10261 (N_10261,N_282,N_4104);
or U10262 (N_10262,N_1903,N_2480);
or U10263 (N_10263,N_3926,N_774);
and U10264 (N_10264,N_4669,N_2260);
nand U10265 (N_10265,N_2795,N_4634);
nor U10266 (N_10266,N_2789,N_5923);
nor U10267 (N_10267,N_2255,N_5001);
xnor U10268 (N_10268,N_694,N_1379);
nand U10269 (N_10269,N_3506,N_4197);
or U10270 (N_10270,N_714,N_5865);
nand U10271 (N_10271,N_3513,N_2993);
or U10272 (N_10272,N_1821,N_1162);
and U10273 (N_10273,N_1777,N_3014);
nor U10274 (N_10274,N_3667,N_4396);
and U10275 (N_10275,N_403,N_2451);
or U10276 (N_10276,N_1513,N_1859);
nor U10277 (N_10277,N_5298,N_5021);
nand U10278 (N_10278,N_5413,N_5806);
or U10279 (N_10279,N_394,N_5251);
xor U10280 (N_10280,N_2207,N_3771);
nand U10281 (N_10281,N_2546,N_2043);
nor U10282 (N_10282,N_4907,N_4180);
nand U10283 (N_10283,N_1579,N_5226);
nor U10284 (N_10284,N_2101,N_1291);
nand U10285 (N_10285,N_986,N_839);
xor U10286 (N_10286,N_4500,N_3915);
and U10287 (N_10287,N_5017,N_3027);
nor U10288 (N_10288,N_5133,N_1487);
and U10289 (N_10289,N_2496,N_3592);
nand U10290 (N_10290,N_3362,N_5611);
and U10291 (N_10291,N_5031,N_1972);
and U10292 (N_10292,N_3422,N_2707);
nor U10293 (N_10293,N_5562,N_5215);
and U10294 (N_10294,N_165,N_3495);
and U10295 (N_10295,N_2271,N_1779);
or U10296 (N_10296,N_4232,N_1452);
nor U10297 (N_10297,N_3607,N_1335);
nand U10298 (N_10298,N_3000,N_5883);
nor U10299 (N_10299,N_2716,N_2910);
or U10300 (N_10300,N_1199,N_4589);
xnor U10301 (N_10301,N_3261,N_5283);
nor U10302 (N_10302,N_1758,N_5654);
xor U10303 (N_10303,N_4546,N_1564);
nand U10304 (N_10304,N_5742,N_2351);
or U10305 (N_10305,N_1898,N_309);
or U10306 (N_10306,N_5097,N_311);
or U10307 (N_10307,N_5466,N_1887);
and U10308 (N_10308,N_5919,N_2038);
nor U10309 (N_10309,N_1192,N_5375);
nor U10310 (N_10310,N_5937,N_2190);
or U10311 (N_10311,N_4899,N_1187);
or U10312 (N_10312,N_5,N_1803);
xor U10313 (N_10313,N_3623,N_3284);
nand U10314 (N_10314,N_4819,N_3386);
or U10315 (N_10315,N_3721,N_3176);
or U10316 (N_10316,N_5995,N_1338);
nand U10317 (N_10317,N_2333,N_4827);
and U10318 (N_10318,N_3616,N_561);
or U10319 (N_10319,N_537,N_4419);
nand U10320 (N_10320,N_5912,N_4926);
and U10321 (N_10321,N_3904,N_2705);
or U10322 (N_10322,N_3946,N_2602);
nand U10323 (N_10323,N_5274,N_5409);
and U10324 (N_10324,N_803,N_3669);
nor U10325 (N_10325,N_1753,N_1674);
nor U10326 (N_10326,N_2256,N_142);
or U10327 (N_10327,N_1015,N_5484);
nand U10328 (N_10328,N_86,N_2928);
or U10329 (N_10329,N_2575,N_1804);
or U10330 (N_10330,N_5633,N_4326);
or U10331 (N_10331,N_3546,N_2360);
or U10332 (N_10332,N_2953,N_2785);
nand U10333 (N_10333,N_4024,N_1195);
xnor U10334 (N_10334,N_1131,N_2899);
and U10335 (N_10335,N_2679,N_4796);
and U10336 (N_10336,N_3627,N_3768);
nand U10337 (N_10337,N_3185,N_2968);
xnor U10338 (N_10338,N_687,N_4369);
and U10339 (N_10339,N_3202,N_3741);
and U10340 (N_10340,N_4479,N_1658);
and U10341 (N_10341,N_405,N_4650);
nor U10342 (N_10342,N_2295,N_4740);
and U10343 (N_10343,N_4577,N_2183);
or U10344 (N_10344,N_307,N_482);
nor U10345 (N_10345,N_3971,N_1942);
nor U10346 (N_10346,N_1043,N_3642);
nand U10347 (N_10347,N_532,N_999);
nor U10348 (N_10348,N_5661,N_1830);
or U10349 (N_10349,N_3625,N_1360);
and U10350 (N_10350,N_2465,N_3874);
or U10351 (N_10351,N_5838,N_5845);
or U10352 (N_10352,N_2747,N_5764);
and U10353 (N_10353,N_3843,N_5850);
nor U10354 (N_10354,N_4020,N_3583);
nand U10355 (N_10355,N_4833,N_3162);
nand U10356 (N_10356,N_1620,N_5632);
or U10357 (N_10357,N_4989,N_2908);
xnor U10358 (N_10358,N_3368,N_3197);
nand U10359 (N_10359,N_2862,N_1039);
or U10360 (N_10360,N_5825,N_4254);
and U10361 (N_10361,N_1445,N_1046);
nand U10362 (N_10362,N_2943,N_477);
or U10363 (N_10363,N_229,N_5108);
or U10364 (N_10364,N_5706,N_1079);
and U10365 (N_10365,N_1804,N_2570);
nor U10366 (N_10366,N_3904,N_4030);
and U10367 (N_10367,N_2867,N_4618);
nor U10368 (N_10368,N_5487,N_1605);
or U10369 (N_10369,N_803,N_550);
and U10370 (N_10370,N_1294,N_5451);
xor U10371 (N_10371,N_3176,N_2195);
or U10372 (N_10372,N_2189,N_824);
and U10373 (N_10373,N_3437,N_3687);
nand U10374 (N_10374,N_527,N_5602);
or U10375 (N_10375,N_3655,N_4235);
and U10376 (N_10376,N_2366,N_4371);
or U10377 (N_10377,N_5059,N_2567);
nand U10378 (N_10378,N_2798,N_2780);
or U10379 (N_10379,N_4015,N_2906);
or U10380 (N_10380,N_1378,N_3903);
nor U10381 (N_10381,N_5193,N_604);
and U10382 (N_10382,N_458,N_4549);
or U10383 (N_10383,N_3038,N_1194);
nor U10384 (N_10384,N_1514,N_651);
nor U10385 (N_10385,N_1905,N_1274);
nand U10386 (N_10386,N_2308,N_5299);
nand U10387 (N_10387,N_4634,N_5644);
or U10388 (N_10388,N_4580,N_1681);
xor U10389 (N_10389,N_4003,N_4807);
and U10390 (N_10390,N_263,N_92);
or U10391 (N_10391,N_2748,N_2608);
and U10392 (N_10392,N_2127,N_94);
xor U10393 (N_10393,N_4948,N_195);
nor U10394 (N_10394,N_2970,N_2037);
and U10395 (N_10395,N_5514,N_2210);
and U10396 (N_10396,N_2974,N_4173);
xor U10397 (N_10397,N_2353,N_4128);
xnor U10398 (N_10398,N_5877,N_1853);
xor U10399 (N_10399,N_3558,N_1286);
or U10400 (N_10400,N_2622,N_1654);
xnor U10401 (N_10401,N_1030,N_3090);
and U10402 (N_10402,N_4303,N_5834);
and U10403 (N_10403,N_3816,N_3149);
and U10404 (N_10404,N_4744,N_4065);
nand U10405 (N_10405,N_4449,N_145);
nor U10406 (N_10406,N_1829,N_5498);
nand U10407 (N_10407,N_151,N_3880);
and U10408 (N_10408,N_4105,N_4223);
and U10409 (N_10409,N_4254,N_4592);
xor U10410 (N_10410,N_2677,N_1665);
nor U10411 (N_10411,N_3457,N_5474);
nand U10412 (N_10412,N_4175,N_4929);
and U10413 (N_10413,N_2750,N_5987);
or U10414 (N_10414,N_1864,N_4651);
or U10415 (N_10415,N_1850,N_5190);
and U10416 (N_10416,N_295,N_345);
and U10417 (N_10417,N_2906,N_3458);
nor U10418 (N_10418,N_1310,N_5939);
or U10419 (N_10419,N_3,N_3492);
and U10420 (N_10420,N_2334,N_5617);
nor U10421 (N_10421,N_5167,N_1316);
and U10422 (N_10422,N_1014,N_3467);
nand U10423 (N_10423,N_4696,N_1503);
nor U10424 (N_10424,N_535,N_430);
nand U10425 (N_10425,N_494,N_1080);
nor U10426 (N_10426,N_4513,N_4629);
and U10427 (N_10427,N_3637,N_4397);
nand U10428 (N_10428,N_2056,N_2548);
or U10429 (N_10429,N_1530,N_752);
nand U10430 (N_10430,N_2671,N_1575);
nor U10431 (N_10431,N_2245,N_3708);
and U10432 (N_10432,N_2489,N_1614);
nand U10433 (N_10433,N_1267,N_274);
nor U10434 (N_10434,N_2049,N_2728);
or U10435 (N_10435,N_1006,N_646);
nor U10436 (N_10436,N_5105,N_3431);
or U10437 (N_10437,N_599,N_3488);
nor U10438 (N_10438,N_4464,N_1553);
xnor U10439 (N_10439,N_705,N_3721);
nor U10440 (N_10440,N_1693,N_458);
xnor U10441 (N_10441,N_954,N_1980);
nor U10442 (N_10442,N_4368,N_3849);
nor U10443 (N_10443,N_2205,N_1586);
and U10444 (N_10444,N_1791,N_276);
nor U10445 (N_10445,N_2095,N_1414);
xnor U10446 (N_10446,N_5141,N_1941);
nand U10447 (N_10447,N_4239,N_2188);
or U10448 (N_10448,N_3521,N_857);
nand U10449 (N_10449,N_3194,N_1575);
and U10450 (N_10450,N_3818,N_333);
or U10451 (N_10451,N_1649,N_1171);
or U10452 (N_10452,N_5964,N_1786);
nor U10453 (N_10453,N_5720,N_2880);
nor U10454 (N_10454,N_761,N_5333);
nor U10455 (N_10455,N_578,N_3544);
nor U10456 (N_10456,N_3662,N_270);
nand U10457 (N_10457,N_1562,N_3274);
nor U10458 (N_10458,N_2763,N_315);
nand U10459 (N_10459,N_4392,N_2263);
xnor U10460 (N_10460,N_3166,N_5869);
xor U10461 (N_10461,N_729,N_2112);
nor U10462 (N_10462,N_5431,N_401);
and U10463 (N_10463,N_2245,N_5316);
nand U10464 (N_10464,N_3482,N_4165);
nor U10465 (N_10465,N_3974,N_2525);
nor U10466 (N_10466,N_3956,N_294);
nand U10467 (N_10467,N_422,N_2614);
and U10468 (N_10468,N_5652,N_436);
nand U10469 (N_10469,N_2823,N_1128);
xor U10470 (N_10470,N_105,N_2836);
nor U10471 (N_10471,N_2314,N_3697);
nor U10472 (N_10472,N_4020,N_4682);
nand U10473 (N_10473,N_1443,N_1995);
nand U10474 (N_10474,N_5263,N_4141);
nor U10475 (N_10475,N_2738,N_4242);
xnor U10476 (N_10476,N_4476,N_5653);
and U10477 (N_10477,N_3117,N_4597);
and U10478 (N_10478,N_1467,N_4658);
and U10479 (N_10479,N_1322,N_1827);
nand U10480 (N_10480,N_416,N_1224);
nor U10481 (N_10481,N_1228,N_765);
nand U10482 (N_10482,N_3559,N_1367);
and U10483 (N_10483,N_3161,N_606);
and U10484 (N_10484,N_4178,N_273);
xor U10485 (N_10485,N_1467,N_990);
nor U10486 (N_10486,N_3035,N_1127);
or U10487 (N_10487,N_277,N_1648);
nand U10488 (N_10488,N_5723,N_2115);
nor U10489 (N_10489,N_970,N_3290);
nor U10490 (N_10490,N_2310,N_3230);
or U10491 (N_10491,N_2432,N_3353);
or U10492 (N_10492,N_3104,N_188);
nand U10493 (N_10493,N_4531,N_788);
nand U10494 (N_10494,N_5740,N_2214);
nor U10495 (N_10495,N_901,N_5348);
and U10496 (N_10496,N_5071,N_3062);
nor U10497 (N_10497,N_2730,N_604);
or U10498 (N_10498,N_777,N_334);
and U10499 (N_10499,N_2380,N_5310);
or U10500 (N_10500,N_2695,N_5448);
nand U10501 (N_10501,N_2925,N_5004);
or U10502 (N_10502,N_5992,N_102);
nand U10503 (N_10503,N_431,N_3439);
nand U10504 (N_10504,N_1558,N_55);
nand U10505 (N_10505,N_681,N_4865);
nor U10506 (N_10506,N_2698,N_5196);
nand U10507 (N_10507,N_1534,N_3803);
and U10508 (N_10508,N_4795,N_2749);
xor U10509 (N_10509,N_4933,N_2316);
nor U10510 (N_10510,N_5960,N_4170);
nand U10511 (N_10511,N_2143,N_5522);
nand U10512 (N_10512,N_5923,N_607);
and U10513 (N_10513,N_5895,N_486);
nand U10514 (N_10514,N_2449,N_5513);
and U10515 (N_10515,N_1263,N_210);
nor U10516 (N_10516,N_5688,N_3385);
or U10517 (N_10517,N_4041,N_971);
nand U10518 (N_10518,N_1587,N_2666);
nor U10519 (N_10519,N_3845,N_2612);
nand U10520 (N_10520,N_1771,N_498);
nand U10521 (N_10521,N_2752,N_5446);
nor U10522 (N_10522,N_2232,N_4244);
nand U10523 (N_10523,N_1113,N_4546);
or U10524 (N_10524,N_180,N_2771);
and U10525 (N_10525,N_15,N_2091);
or U10526 (N_10526,N_4359,N_5500);
and U10527 (N_10527,N_431,N_5767);
or U10528 (N_10528,N_1183,N_5563);
nand U10529 (N_10529,N_3061,N_5299);
or U10530 (N_10530,N_233,N_914);
nor U10531 (N_10531,N_5699,N_4948);
nand U10532 (N_10532,N_1608,N_1392);
xor U10533 (N_10533,N_3169,N_2404);
and U10534 (N_10534,N_5917,N_2208);
nor U10535 (N_10535,N_267,N_3417);
nor U10536 (N_10536,N_5371,N_5875);
nand U10537 (N_10537,N_947,N_3225);
and U10538 (N_10538,N_1721,N_3361);
nand U10539 (N_10539,N_2445,N_1485);
nor U10540 (N_10540,N_1101,N_344);
or U10541 (N_10541,N_4720,N_3195);
or U10542 (N_10542,N_2143,N_1424);
nand U10543 (N_10543,N_2986,N_1757);
nand U10544 (N_10544,N_320,N_3706);
nand U10545 (N_10545,N_4622,N_5075);
and U10546 (N_10546,N_4109,N_166);
nor U10547 (N_10547,N_5960,N_4609);
or U10548 (N_10548,N_3839,N_1294);
or U10549 (N_10549,N_5146,N_1423);
nor U10550 (N_10550,N_4288,N_2104);
nand U10551 (N_10551,N_5148,N_722);
or U10552 (N_10552,N_1711,N_5290);
nand U10553 (N_10553,N_5766,N_4006);
and U10554 (N_10554,N_3146,N_1014);
xor U10555 (N_10555,N_5941,N_351);
nor U10556 (N_10556,N_3174,N_1810);
and U10557 (N_10557,N_2116,N_3313);
nand U10558 (N_10558,N_228,N_3235);
or U10559 (N_10559,N_46,N_4956);
or U10560 (N_10560,N_843,N_5973);
nand U10561 (N_10561,N_5755,N_4760);
xnor U10562 (N_10562,N_55,N_1164);
nor U10563 (N_10563,N_2452,N_1193);
nor U10564 (N_10564,N_343,N_2076);
and U10565 (N_10565,N_4492,N_3082);
nand U10566 (N_10566,N_108,N_2810);
nor U10567 (N_10567,N_3685,N_5484);
nand U10568 (N_10568,N_4436,N_1486);
nand U10569 (N_10569,N_5678,N_5591);
xnor U10570 (N_10570,N_4953,N_2635);
nand U10571 (N_10571,N_4544,N_2424);
nand U10572 (N_10572,N_4490,N_5878);
and U10573 (N_10573,N_2150,N_2055);
xor U10574 (N_10574,N_3081,N_972);
xor U10575 (N_10575,N_1145,N_2796);
and U10576 (N_10576,N_5934,N_4710);
and U10577 (N_10577,N_1767,N_1225);
or U10578 (N_10578,N_661,N_4101);
nor U10579 (N_10579,N_5632,N_2720);
nand U10580 (N_10580,N_5090,N_725);
and U10581 (N_10581,N_4866,N_844);
xor U10582 (N_10582,N_183,N_646);
xnor U10583 (N_10583,N_3512,N_4685);
nor U10584 (N_10584,N_67,N_3235);
and U10585 (N_10585,N_1867,N_455);
nand U10586 (N_10586,N_4863,N_1426);
or U10587 (N_10587,N_4333,N_5197);
or U10588 (N_10588,N_2024,N_3067);
nor U10589 (N_10589,N_5969,N_5147);
and U10590 (N_10590,N_631,N_4134);
and U10591 (N_10591,N_1858,N_2910);
and U10592 (N_10592,N_1866,N_2356);
nor U10593 (N_10593,N_177,N_2582);
and U10594 (N_10594,N_2861,N_5507);
and U10595 (N_10595,N_5680,N_1510);
nor U10596 (N_10596,N_1327,N_5209);
or U10597 (N_10597,N_1563,N_4064);
nor U10598 (N_10598,N_5746,N_32);
nor U10599 (N_10599,N_1757,N_1007);
nor U10600 (N_10600,N_4318,N_1316);
and U10601 (N_10601,N_4848,N_3706);
nand U10602 (N_10602,N_2631,N_5047);
or U10603 (N_10603,N_2355,N_3732);
and U10604 (N_10604,N_2938,N_5662);
or U10605 (N_10605,N_2804,N_107);
and U10606 (N_10606,N_5325,N_1733);
and U10607 (N_10607,N_3932,N_2919);
nor U10608 (N_10608,N_3083,N_4507);
nand U10609 (N_10609,N_2045,N_5575);
nor U10610 (N_10610,N_14,N_4702);
xor U10611 (N_10611,N_3385,N_4903);
nor U10612 (N_10612,N_1976,N_242);
and U10613 (N_10613,N_3297,N_5916);
nand U10614 (N_10614,N_1223,N_673);
nor U10615 (N_10615,N_3496,N_1419);
xor U10616 (N_10616,N_3549,N_2929);
nand U10617 (N_10617,N_521,N_2797);
or U10618 (N_10618,N_5444,N_3130);
and U10619 (N_10619,N_4646,N_687);
xnor U10620 (N_10620,N_1101,N_5097);
nand U10621 (N_10621,N_5860,N_5880);
nor U10622 (N_10622,N_3822,N_5244);
nor U10623 (N_10623,N_1001,N_5788);
nor U10624 (N_10624,N_3076,N_2810);
nand U10625 (N_10625,N_3457,N_5571);
nand U10626 (N_10626,N_799,N_4994);
and U10627 (N_10627,N_1931,N_2472);
and U10628 (N_10628,N_650,N_5777);
and U10629 (N_10629,N_2996,N_2520);
nand U10630 (N_10630,N_5680,N_5459);
or U10631 (N_10631,N_426,N_4702);
nor U10632 (N_10632,N_4242,N_3593);
nand U10633 (N_10633,N_5458,N_1877);
nand U10634 (N_10634,N_562,N_4133);
nand U10635 (N_10635,N_3091,N_2224);
nor U10636 (N_10636,N_854,N_2907);
or U10637 (N_10637,N_4860,N_4739);
nand U10638 (N_10638,N_3639,N_2601);
nand U10639 (N_10639,N_1077,N_5512);
or U10640 (N_10640,N_5238,N_1430);
and U10641 (N_10641,N_2310,N_855);
nand U10642 (N_10642,N_4201,N_5190);
nor U10643 (N_10643,N_0,N_2648);
nor U10644 (N_10644,N_4867,N_2359);
and U10645 (N_10645,N_5347,N_2930);
nand U10646 (N_10646,N_4272,N_3001);
nor U10647 (N_10647,N_4915,N_5947);
nand U10648 (N_10648,N_1575,N_146);
or U10649 (N_10649,N_4941,N_4477);
and U10650 (N_10650,N_376,N_3574);
or U10651 (N_10651,N_5127,N_718);
and U10652 (N_10652,N_4895,N_3475);
nand U10653 (N_10653,N_5092,N_4839);
nand U10654 (N_10654,N_277,N_5299);
or U10655 (N_10655,N_1266,N_215);
or U10656 (N_10656,N_4285,N_2794);
or U10657 (N_10657,N_15,N_2495);
nor U10658 (N_10658,N_5976,N_5573);
or U10659 (N_10659,N_5361,N_4598);
or U10660 (N_10660,N_1616,N_2069);
and U10661 (N_10661,N_4522,N_5213);
or U10662 (N_10662,N_593,N_3485);
nor U10663 (N_10663,N_653,N_3684);
nand U10664 (N_10664,N_4210,N_3794);
xnor U10665 (N_10665,N_1151,N_4653);
nand U10666 (N_10666,N_3784,N_3761);
or U10667 (N_10667,N_2143,N_3047);
xor U10668 (N_10668,N_3768,N_1877);
nand U10669 (N_10669,N_3469,N_787);
nand U10670 (N_10670,N_358,N_676);
nand U10671 (N_10671,N_3675,N_5552);
or U10672 (N_10672,N_4660,N_1943);
nand U10673 (N_10673,N_3120,N_5238);
and U10674 (N_10674,N_1164,N_4020);
nor U10675 (N_10675,N_2059,N_2449);
and U10676 (N_10676,N_239,N_5991);
and U10677 (N_10677,N_4633,N_1076);
and U10678 (N_10678,N_114,N_4742);
and U10679 (N_10679,N_1246,N_4138);
nand U10680 (N_10680,N_2594,N_2228);
or U10681 (N_10681,N_4872,N_565);
and U10682 (N_10682,N_2361,N_5583);
nand U10683 (N_10683,N_595,N_4654);
nor U10684 (N_10684,N_191,N_1824);
xor U10685 (N_10685,N_482,N_4059);
and U10686 (N_10686,N_5657,N_2996);
nor U10687 (N_10687,N_1875,N_1892);
nand U10688 (N_10688,N_5232,N_383);
and U10689 (N_10689,N_2883,N_5107);
or U10690 (N_10690,N_3718,N_2766);
or U10691 (N_10691,N_2056,N_3346);
nor U10692 (N_10692,N_3886,N_5527);
nor U10693 (N_10693,N_3562,N_4178);
nor U10694 (N_10694,N_1983,N_2869);
nor U10695 (N_10695,N_4758,N_5136);
and U10696 (N_10696,N_3782,N_2287);
nor U10697 (N_10697,N_5545,N_1471);
nor U10698 (N_10698,N_4500,N_2893);
xnor U10699 (N_10699,N_3600,N_1378);
nand U10700 (N_10700,N_3995,N_1113);
nand U10701 (N_10701,N_1010,N_3712);
nand U10702 (N_10702,N_3015,N_4654);
nand U10703 (N_10703,N_5744,N_5568);
nand U10704 (N_10704,N_3983,N_1531);
and U10705 (N_10705,N_1364,N_4833);
and U10706 (N_10706,N_3873,N_2465);
nand U10707 (N_10707,N_419,N_5255);
nand U10708 (N_10708,N_1261,N_3154);
nor U10709 (N_10709,N_4568,N_4023);
xor U10710 (N_10710,N_1705,N_709);
nand U10711 (N_10711,N_1312,N_5247);
and U10712 (N_10712,N_3294,N_5593);
nor U10713 (N_10713,N_2002,N_3285);
and U10714 (N_10714,N_4789,N_382);
nand U10715 (N_10715,N_1004,N_5297);
and U10716 (N_10716,N_3413,N_976);
nand U10717 (N_10717,N_3834,N_4628);
nand U10718 (N_10718,N_2025,N_427);
nand U10719 (N_10719,N_1545,N_765);
and U10720 (N_10720,N_741,N_2901);
or U10721 (N_10721,N_5545,N_1756);
and U10722 (N_10722,N_1932,N_565);
or U10723 (N_10723,N_2567,N_2226);
and U10724 (N_10724,N_724,N_2656);
and U10725 (N_10725,N_3245,N_970);
or U10726 (N_10726,N_3807,N_876);
xnor U10727 (N_10727,N_96,N_32);
nand U10728 (N_10728,N_5064,N_1161);
nand U10729 (N_10729,N_3139,N_2843);
nand U10730 (N_10730,N_316,N_3250);
nand U10731 (N_10731,N_4678,N_1000);
nand U10732 (N_10732,N_4451,N_4902);
or U10733 (N_10733,N_1096,N_5041);
or U10734 (N_10734,N_204,N_1262);
and U10735 (N_10735,N_3912,N_1592);
nand U10736 (N_10736,N_1217,N_5949);
nor U10737 (N_10737,N_1539,N_1829);
and U10738 (N_10738,N_4218,N_4234);
xnor U10739 (N_10739,N_171,N_3767);
xnor U10740 (N_10740,N_289,N_457);
and U10741 (N_10741,N_1734,N_1991);
or U10742 (N_10742,N_2831,N_1495);
nand U10743 (N_10743,N_775,N_5600);
nor U10744 (N_10744,N_5453,N_2727);
and U10745 (N_10745,N_3722,N_1653);
nor U10746 (N_10746,N_2947,N_3118);
nor U10747 (N_10747,N_2531,N_5656);
nor U10748 (N_10748,N_4386,N_4856);
nor U10749 (N_10749,N_2484,N_2111);
or U10750 (N_10750,N_5842,N_4758);
and U10751 (N_10751,N_5432,N_1336);
nor U10752 (N_10752,N_2308,N_5752);
nand U10753 (N_10753,N_4650,N_3841);
nand U10754 (N_10754,N_5030,N_5462);
nand U10755 (N_10755,N_3436,N_230);
xnor U10756 (N_10756,N_5385,N_2803);
xor U10757 (N_10757,N_2639,N_4903);
or U10758 (N_10758,N_4638,N_2808);
nand U10759 (N_10759,N_2197,N_2515);
or U10760 (N_10760,N_565,N_2889);
or U10761 (N_10761,N_4337,N_5762);
nand U10762 (N_10762,N_5884,N_4952);
and U10763 (N_10763,N_4876,N_3041);
xor U10764 (N_10764,N_3654,N_1739);
and U10765 (N_10765,N_5274,N_1227);
nor U10766 (N_10766,N_364,N_2026);
nor U10767 (N_10767,N_2222,N_2526);
nand U10768 (N_10768,N_5626,N_4112);
nor U10769 (N_10769,N_1266,N_4302);
nor U10770 (N_10770,N_1767,N_2142);
xor U10771 (N_10771,N_660,N_4909);
or U10772 (N_10772,N_2463,N_1068);
nand U10773 (N_10773,N_5220,N_5075);
nand U10774 (N_10774,N_3598,N_4471);
or U10775 (N_10775,N_2340,N_649);
nand U10776 (N_10776,N_3478,N_2240);
xnor U10777 (N_10777,N_2087,N_2661);
and U10778 (N_10778,N_3015,N_1328);
and U10779 (N_10779,N_5907,N_369);
nand U10780 (N_10780,N_549,N_5331);
nand U10781 (N_10781,N_2735,N_5988);
nor U10782 (N_10782,N_0,N_1787);
xor U10783 (N_10783,N_581,N_4986);
xnor U10784 (N_10784,N_5996,N_1406);
or U10785 (N_10785,N_4215,N_395);
nand U10786 (N_10786,N_4668,N_3715);
and U10787 (N_10787,N_2957,N_2573);
nor U10788 (N_10788,N_4499,N_2846);
nand U10789 (N_10789,N_3880,N_4308);
nand U10790 (N_10790,N_3712,N_53);
or U10791 (N_10791,N_5321,N_2113);
xor U10792 (N_10792,N_3763,N_4451);
and U10793 (N_10793,N_4713,N_1369);
or U10794 (N_10794,N_2819,N_5188);
or U10795 (N_10795,N_4713,N_418);
xor U10796 (N_10796,N_1332,N_1175);
or U10797 (N_10797,N_2681,N_562);
nand U10798 (N_10798,N_3724,N_837);
and U10799 (N_10799,N_4689,N_2604);
and U10800 (N_10800,N_2562,N_5447);
xnor U10801 (N_10801,N_2122,N_3684);
or U10802 (N_10802,N_1385,N_4562);
and U10803 (N_10803,N_5162,N_4828);
and U10804 (N_10804,N_4116,N_3346);
and U10805 (N_10805,N_5999,N_3336);
nor U10806 (N_10806,N_176,N_868);
and U10807 (N_10807,N_4722,N_5097);
nor U10808 (N_10808,N_2836,N_3417);
nor U10809 (N_10809,N_219,N_1226);
nand U10810 (N_10810,N_5942,N_420);
nand U10811 (N_10811,N_5054,N_3654);
and U10812 (N_10812,N_2218,N_2203);
or U10813 (N_10813,N_4746,N_5759);
or U10814 (N_10814,N_3891,N_232);
nand U10815 (N_10815,N_2377,N_4219);
and U10816 (N_10816,N_758,N_4657);
and U10817 (N_10817,N_330,N_2503);
nor U10818 (N_10818,N_3627,N_2323);
nand U10819 (N_10819,N_1546,N_3974);
nor U10820 (N_10820,N_3732,N_3685);
and U10821 (N_10821,N_2078,N_212);
nor U10822 (N_10822,N_2666,N_4673);
or U10823 (N_10823,N_4350,N_3754);
nor U10824 (N_10824,N_5124,N_2393);
and U10825 (N_10825,N_1127,N_973);
nand U10826 (N_10826,N_126,N_2523);
or U10827 (N_10827,N_2298,N_2371);
xnor U10828 (N_10828,N_3626,N_3085);
or U10829 (N_10829,N_741,N_3932);
and U10830 (N_10830,N_1635,N_4004);
and U10831 (N_10831,N_5202,N_2170);
nor U10832 (N_10832,N_5637,N_4017);
nor U10833 (N_10833,N_1165,N_5909);
or U10834 (N_10834,N_1824,N_1255);
or U10835 (N_10835,N_4790,N_1078);
nor U10836 (N_10836,N_4229,N_276);
xor U10837 (N_10837,N_1233,N_475);
nor U10838 (N_10838,N_5823,N_5311);
xnor U10839 (N_10839,N_1644,N_2796);
or U10840 (N_10840,N_3116,N_1961);
nand U10841 (N_10841,N_3257,N_3437);
or U10842 (N_10842,N_3363,N_1755);
nor U10843 (N_10843,N_1997,N_4616);
or U10844 (N_10844,N_3538,N_952);
nand U10845 (N_10845,N_3364,N_1227);
or U10846 (N_10846,N_92,N_2287);
and U10847 (N_10847,N_5197,N_5366);
or U10848 (N_10848,N_4553,N_809);
or U10849 (N_10849,N_4114,N_4465);
or U10850 (N_10850,N_3605,N_3414);
nor U10851 (N_10851,N_153,N_3349);
xnor U10852 (N_10852,N_3809,N_5750);
nand U10853 (N_10853,N_1194,N_2489);
xor U10854 (N_10854,N_5290,N_3245);
nand U10855 (N_10855,N_4849,N_913);
and U10856 (N_10856,N_4015,N_3172);
xor U10857 (N_10857,N_2294,N_4756);
or U10858 (N_10858,N_5531,N_1291);
nor U10859 (N_10859,N_4544,N_4254);
and U10860 (N_10860,N_786,N_229);
nor U10861 (N_10861,N_2128,N_4824);
or U10862 (N_10862,N_1254,N_1407);
or U10863 (N_10863,N_4919,N_574);
and U10864 (N_10864,N_1210,N_1840);
or U10865 (N_10865,N_5391,N_1398);
or U10866 (N_10866,N_2303,N_459);
nand U10867 (N_10867,N_761,N_1121);
or U10868 (N_10868,N_1631,N_5719);
nand U10869 (N_10869,N_3844,N_5577);
xnor U10870 (N_10870,N_318,N_384);
nand U10871 (N_10871,N_3755,N_403);
nand U10872 (N_10872,N_4885,N_649);
or U10873 (N_10873,N_4286,N_552);
nand U10874 (N_10874,N_905,N_794);
nand U10875 (N_10875,N_3188,N_2400);
nand U10876 (N_10876,N_1049,N_1678);
and U10877 (N_10877,N_5320,N_2087);
and U10878 (N_10878,N_1903,N_3318);
or U10879 (N_10879,N_308,N_2376);
xor U10880 (N_10880,N_2519,N_2201);
nor U10881 (N_10881,N_5404,N_1218);
xnor U10882 (N_10882,N_3150,N_1718);
nand U10883 (N_10883,N_1380,N_5539);
xnor U10884 (N_10884,N_4928,N_1546);
nand U10885 (N_10885,N_568,N_4827);
nand U10886 (N_10886,N_2682,N_3545);
or U10887 (N_10887,N_4639,N_2713);
nor U10888 (N_10888,N_4699,N_5056);
or U10889 (N_10889,N_975,N_4394);
and U10890 (N_10890,N_713,N_5175);
nand U10891 (N_10891,N_5954,N_3387);
and U10892 (N_10892,N_4843,N_2845);
or U10893 (N_10893,N_1342,N_339);
nand U10894 (N_10894,N_5645,N_5558);
or U10895 (N_10895,N_405,N_5403);
nand U10896 (N_10896,N_5247,N_5813);
and U10897 (N_10897,N_2126,N_4079);
or U10898 (N_10898,N_1874,N_3170);
or U10899 (N_10899,N_4062,N_3787);
nand U10900 (N_10900,N_701,N_3035);
nand U10901 (N_10901,N_5389,N_1521);
nor U10902 (N_10902,N_2383,N_1220);
nor U10903 (N_10903,N_3870,N_1185);
and U10904 (N_10904,N_5785,N_3874);
nor U10905 (N_10905,N_1848,N_471);
nand U10906 (N_10906,N_5711,N_2322);
and U10907 (N_10907,N_984,N_5588);
nand U10908 (N_10908,N_5485,N_3170);
nor U10909 (N_10909,N_1385,N_5740);
nand U10910 (N_10910,N_1904,N_2843);
or U10911 (N_10911,N_1033,N_2324);
nor U10912 (N_10912,N_5862,N_3422);
nor U10913 (N_10913,N_4202,N_3427);
nand U10914 (N_10914,N_2758,N_5151);
nand U10915 (N_10915,N_5382,N_2505);
or U10916 (N_10916,N_1145,N_4237);
and U10917 (N_10917,N_456,N_5650);
nand U10918 (N_10918,N_898,N_1188);
and U10919 (N_10919,N_4491,N_4134);
and U10920 (N_10920,N_4588,N_5845);
or U10921 (N_10921,N_3598,N_261);
nand U10922 (N_10922,N_713,N_81);
nand U10923 (N_10923,N_4093,N_3946);
nand U10924 (N_10924,N_4083,N_667);
nor U10925 (N_10925,N_1169,N_1798);
and U10926 (N_10926,N_2112,N_5381);
and U10927 (N_10927,N_1112,N_4074);
and U10928 (N_10928,N_2592,N_916);
and U10929 (N_10929,N_5175,N_3664);
or U10930 (N_10930,N_1672,N_652);
and U10931 (N_10931,N_113,N_2051);
nand U10932 (N_10932,N_5282,N_1446);
and U10933 (N_10933,N_5092,N_3712);
or U10934 (N_10934,N_65,N_561);
and U10935 (N_10935,N_80,N_106);
nand U10936 (N_10936,N_5909,N_423);
or U10937 (N_10937,N_1130,N_992);
xnor U10938 (N_10938,N_5589,N_5673);
or U10939 (N_10939,N_2628,N_2690);
nand U10940 (N_10940,N_4149,N_1228);
nand U10941 (N_10941,N_4538,N_5668);
nor U10942 (N_10942,N_2041,N_772);
or U10943 (N_10943,N_5810,N_4354);
xor U10944 (N_10944,N_2185,N_4020);
nor U10945 (N_10945,N_4730,N_357);
and U10946 (N_10946,N_5237,N_3119);
nor U10947 (N_10947,N_4218,N_703);
and U10948 (N_10948,N_4329,N_2590);
nor U10949 (N_10949,N_55,N_1993);
nor U10950 (N_10950,N_4234,N_1451);
xnor U10951 (N_10951,N_1643,N_3164);
or U10952 (N_10952,N_3418,N_364);
and U10953 (N_10953,N_731,N_4079);
or U10954 (N_10954,N_3454,N_3475);
or U10955 (N_10955,N_1877,N_4786);
xnor U10956 (N_10956,N_4602,N_2004);
or U10957 (N_10957,N_2291,N_1075);
nand U10958 (N_10958,N_2756,N_1891);
and U10959 (N_10959,N_4226,N_4798);
and U10960 (N_10960,N_4179,N_99);
or U10961 (N_10961,N_3251,N_3865);
nor U10962 (N_10962,N_3542,N_2679);
xor U10963 (N_10963,N_2094,N_5289);
nand U10964 (N_10964,N_2526,N_100);
and U10965 (N_10965,N_5372,N_1943);
nor U10966 (N_10966,N_5103,N_5718);
or U10967 (N_10967,N_5943,N_5261);
xnor U10968 (N_10968,N_5345,N_5659);
xnor U10969 (N_10969,N_147,N_1091);
xor U10970 (N_10970,N_5169,N_4956);
or U10971 (N_10971,N_1701,N_428);
nor U10972 (N_10972,N_11,N_661);
nor U10973 (N_10973,N_582,N_4520);
nor U10974 (N_10974,N_744,N_1839);
nor U10975 (N_10975,N_3080,N_136);
or U10976 (N_10976,N_5628,N_1264);
or U10977 (N_10977,N_3197,N_3760);
or U10978 (N_10978,N_3463,N_717);
nor U10979 (N_10979,N_855,N_3663);
or U10980 (N_10980,N_1026,N_1841);
or U10981 (N_10981,N_2266,N_4271);
and U10982 (N_10982,N_5443,N_52);
nand U10983 (N_10983,N_3163,N_3027);
and U10984 (N_10984,N_5205,N_2755);
nor U10985 (N_10985,N_3424,N_1778);
nand U10986 (N_10986,N_1008,N_2618);
nor U10987 (N_10987,N_4836,N_3560);
and U10988 (N_10988,N_2151,N_2942);
and U10989 (N_10989,N_4216,N_5682);
nand U10990 (N_10990,N_4032,N_4906);
or U10991 (N_10991,N_2597,N_2135);
and U10992 (N_10992,N_3256,N_3669);
and U10993 (N_10993,N_2445,N_1133);
and U10994 (N_10994,N_3567,N_1259);
or U10995 (N_10995,N_5233,N_3424);
or U10996 (N_10996,N_280,N_1593);
nand U10997 (N_10997,N_2325,N_5145);
xnor U10998 (N_10998,N_253,N_2860);
and U10999 (N_10999,N_2138,N_5459);
or U11000 (N_11000,N_708,N_3327);
and U11001 (N_11001,N_3752,N_3285);
or U11002 (N_11002,N_2274,N_5888);
and U11003 (N_11003,N_3760,N_777);
or U11004 (N_11004,N_5447,N_1600);
and U11005 (N_11005,N_76,N_2404);
nor U11006 (N_11006,N_4021,N_1053);
or U11007 (N_11007,N_977,N_4768);
or U11008 (N_11008,N_4031,N_2735);
and U11009 (N_11009,N_2020,N_5092);
nor U11010 (N_11010,N_2831,N_4402);
xor U11011 (N_11011,N_3440,N_5525);
or U11012 (N_11012,N_5255,N_4111);
nor U11013 (N_11013,N_2461,N_220);
nor U11014 (N_11014,N_2414,N_2182);
and U11015 (N_11015,N_2326,N_5295);
and U11016 (N_11016,N_851,N_4615);
nor U11017 (N_11017,N_5567,N_4213);
xor U11018 (N_11018,N_5049,N_1676);
xnor U11019 (N_11019,N_2162,N_790);
xor U11020 (N_11020,N_915,N_2507);
or U11021 (N_11021,N_193,N_1294);
and U11022 (N_11022,N_4190,N_3798);
nor U11023 (N_11023,N_5398,N_1163);
and U11024 (N_11024,N_4946,N_1818);
and U11025 (N_11025,N_5929,N_1254);
nand U11026 (N_11026,N_3062,N_2908);
and U11027 (N_11027,N_1652,N_4345);
nor U11028 (N_11028,N_4874,N_883);
and U11029 (N_11029,N_4885,N_4681);
nand U11030 (N_11030,N_5175,N_2962);
and U11031 (N_11031,N_5969,N_5401);
and U11032 (N_11032,N_3620,N_1146);
nor U11033 (N_11033,N_5362,N_5920);
nand U11034 (N_11034,N_3826,N_2161);
or U11035 (N_11035,N_3042,N_3398);
nor U11036 (N_11036,N_1210,N_609);
or U11037 (N_11037,N_4097,N_1144);
and U11038 (N_11038,N_4191,N_3042);
nand U11039 (N_11039,N_2149,N_2192);
xor U11040 (N_11040,N_4865,N_5645);
xnor U11041 (N_11041,N_5132,N_1789);
and U11042 (N_11042,N_5794,N_5633);
nor U11043 (N_11043,N_5572,N_4728);
xnor U11044 (N_11044,N_1865,N_3984);
nand U11045 (N_11045,N_5615,N_4862);
nor U11046 (N_11046,N_4533,N_3652);
nor U11047 (N_11047,N_1305,N_4235);
and U11048 (N_11048,N_4069,N_214);
nor U11049 (N_11049,N_1661,N_977);
or U11050 (N_11050,N_4106,N_4279);
and U11051 (N_11051,N_2290,N_3588);
nor U11052 (N_11052,N_435,N_468);
xnor U11053 (N_11053,N_2769,N_400);
nor U11054 (N_11054,N_1787,N_2179);
and U11055 (N_11055,N_4515,N_2530);
xnor U11056 (N_11056,N_4054,N_3777);
and U11057 (N_11057,N_2484,N_979);
or U11058 (N_11058,N_5128,N_2375);
nand U11059 (N_11059,N_2462,N_177);
or U11060 (N_11060,N_1717,N_836);
nor U11061 (N_11061,N_532,N_721);
or U11062 (N_11062,N_3584,N_1839);
nor U11063 (N_11063,N_3455,N_4912);
or U11064 (N_11064,N_951,N_2351);
nor U11065 (N_11065,N_5819,N_571);
and U11066 (N_11066,N_2710,N_4733);
or U11067 (N_11067,N_2382,N_4299);
nand U11068 (N_11068,N_612,N_2128);
or U11069 (N_11069,N_513,N_764);
nor U11070 (N_11070,N_5160,N_44);
and U11071 (N_11071,N_5944,N_3912);
xor U11072 (N_11072,N_4754,N_1790);
or U11073 (N_11073,N_3898,N_543);
and U11074 (N_11074,N_5227,N_4844);
nor U11075 (N_11075,N_5740,N_3858);
nand U11076 (N_11076,N_157,N_132);
nand U11077 (N_11077,N_913,N_2991);
nor U11078 (N_11078,N_3837,N_3955);
or U11079 (N_11079,N_3186,N_5969);
nor U11080 (N_11080,N_4273,N_3119);
nor U11081 (N_11081,N_1820,N_2144);
or U11082 (N_11082,N_3761,N_238);
xor U11083 (N_11083,N_4325,N_1505);
or U11084 (N_11084,N_5986,N_1974);
nor U11085 (N_11085,N_5383,N_3383);
nand U11086 (N_11086,N_4390,N_426);
or U11087 (N_11087,N_5842,N_3450);
and U11088 (N_11088,N_289,N_4679);
or U11089 (N_11089,N_4231,N_894);
nor U11090 (N_11090,N_923,N_54);
nand U11091 (N_11091,N_1302,N_1388);
or U11092 (N_11092,N_697,N_4565);
nor U11093 (N_11093,N_1286,N_1687);
nand U11094 (N_11094,N_3873,N_3834);
and U11095 (N_11095,N_110,N_2645);
and U11096 (N_11096,N_3231,N_286);
nor U11097 (N_11097,N_2789,N_1085);
nor U11098 (N_11098,N_3735,N_2022);
xor U11099 (N_11099,N_1596,N_5079);
xor U11100 (N_11100,N_2587,N_3276);
nor U11101 (N_11101,N_3450,N_444);
or U11102 (N_11102,N_5869,N_2374);
nand U11103 (N_11103,N_529,N_5642);
nand U11104 (N_11104,N_1452,N_5908);
or U11105 (N_11105,N_1765,N_2671);
nand U11106 (N_11106,N_1162,N_2312);
and U11107 (N_11107,N_5859,N_314);
xor U11108 (N_11108,N_2601,N_4617);
and U11109 (N_11109,N_471,N_4499);
nand U11110 (N_11110,N_202,N_3146);
nor U11111 (N_11111,N_358,N_2467);
nor U11112 (N_11112,N_753,N_4124);
nand U11113 (N_11113,N_4504,N_1627);
nor U11114 (N_11114,N_3227,N_1326);
nor U11115 (N_11115,N_3778,N_364);
or U11116 (N_11116,N_3904,N_3633);
and U11117 (N_11117,N_1559,N_919);
or U11118 (N_11118,N_4153,N_2186);
or U11119 (N_11119,N_2242,N_5230);
and U11120 (N_11120,N_2018,N_419);
nand U11121 (N_11121,N_3574,N_733);
nand U11122 (N_11122,N_3732,N_615);
or U11123 (N_11123,N_3104,N_2562);
nand U11124 (N_11124,N_2246,N_5886);
and U11125 (N_11125,N_1458,N_3184);
or U11126 (N_11126,N_2062,N_338);
or U11127 (N_11127,N_546,N_2897);
nand U11128 (N_11128,N_4187,N_5959);
and U11129 (N_11129,N_4028,N_3237);
or U11130 (N_11130,N_2439,N_3538);
or U11131 (N_11131,N_3795,N_748);
nor U11132 (N_11132,N_3539,N_5476);
and U11133 (N_11133,N_125,N_4884);
and U11134 (N_11134,N_493,N_4006);
nor U11135 (N_11135,N_2265,N_2689);
and U11136 (N_11136,N_1899,N_2146);
or U11137 (N_11137,N_4386,N_4613);
nor U11138 (N_11138,N_5581,N_5052);
nor U11139 (N_11139,N_5224,N_4123);
or U11140 (N_11140,N_4750,N_4245);
nor U11141 (N_11141,N_935,N_53);
or U11142 (N_11142,N_5594,N_2458);
and U11143 (N_11143,N_96,N_2853);
nand U11144 (N_11144,N_3251,N_5508);
nor U11145 (N_11145,N_1378,N_5359);
or U11146 (N_11146,N_1491,N_3251);
and U11147 (N_11147,N_3517,N_5861);
or U11148 (N_11148,N_1892,N_3669);
or U11149 (N_11149,N_4321,N_5656);
or U11150 (N_11150,N_3463,N_1117);
or U11151 (N_11151,N_768,N_1801);
nand U11152 (N_11152,N_5903,N_94);
and U11153 (N_11153,N_2386,N_3652);
xnor U11154 (N_11154,N_5872,N_4589);
or U11155 (N_11155,N_4091,N_736);
or U11156 (N_11156,N_774,N_1409);
nand U11157 (N_11157,N_5579,N_5978);
and U11158 (N_11158,N_2230,N_823);
xor U11159 (N_11159,N_4829,N_4555);
nand U11160 (N_11160,N_5104,N_670);
xnor U11161 (N_11161,N_3661,N_4097);
and U11162 (N_11162,N_465,N_3600);
nand U11163 (N_11163,N_5945,N_87);
and U11164 (N_11164,N_2580,N_1798);
nor U11165 (N_11165,N_1921,N_1290);
nand U11166 (N_11166,N_4077,N_4146);
nor U11167 (N_11167,N_3466,N_4169);
nor U11168 (N_11168,N_3279,N_1389);
nor U11169 (N_11169,N_4007,N_2794);
or U11170 (N_11170,N_792,N_5413);
nand U11171 (N_11171,N_2718,N_805);
and U11172 (N_11172,N_191,N_675);
nor U11173 (N_11173,N_840,N_1838);
nand U11174 (N_11174,N_2851,N_5305);
and U11175 (N_11175,N_1273,N_1498);
nand U11176 (N_11176,N_4296,N_3801);
nor U11177 (N_11177,N_655,N_1397);
and U11178 (N_11178,N_2620,N_2248);
or U11179 (N_11179,N_3297,N_2076);
xnor U11180 (N_11180,N_166,N_2654);
nand U11181 (N_11181,N_5707,N_4082);
and U11182 (N_11182,N_3628,N_3854);
and U11183 (N_11183,N_1341,N_4888);
or U11184 (N_11184,N_2793,N_5908);
nor U11185 (N_11185,N_1093,N_5630);
xor U11186 (N_11186,N_5348,N_616);
or U11187 (N_11187,N_5276,N_237);
or U11188 (N_11188,N_4438,N_402);
nand U11189 (N_11189,N_1747,N_2983);
and U11190 (N_11190,N_1786,N_919);
nor U11191 (N_11191,N_725,N_4220);
nor U11192 (N_11192,N_1749,N_4375);
nor U11193 (N_11193,N_4104,N_2591);
nand U11194 (N_11194,N_4233,N_2373);
nor U11195 (N_11195,N_2613,N_4459);
nand U11196 (N_11196,N_1600,N_1715);
and U11197 (N_11197,N_4696,N_3919);
or U11198 (N_11198,N_5431,N_5169);
and U11199 (N_11199,N_4057,N_334);
nand U11200 (N_11200,N_1994,N_1355);
or U11201 (N_11201,N_5094,N_673);
or U11202 (N_11202,N_5692,N_1318);
or U11203 (N_11203,N_3097,N_3180);
or U11204 (N_11204,N_3526,N_5574);
xnor U11205 (N_11205,N_5786,N_3720);
nand U11206 (N_11206,N_1442,N_2600);
or U11207 (N_11207,N_5454,N_3679);
nand U11208 (N_11208,N_2577,N_3966);
xnor U11209 (N_11209,N_2283,N_1176);
xnor U11210 (N_11210,N_5194,N_1424);
and U11211 (N_11211,N_3162,N_738);
and U11212 (N_11212,N_621,N_5127);
xnor U11213 (N_11213,N_3233,N_2408);
nor U11214 (N_11214,N_4310,N_3643);
or U11215 (N_11215,N_4360,N_2341);
and U11216 (N_11216,N_5867,N_3967);
nand U11217 (N_11217,N_995,N_1857);
nor U11218 (N_11218,N_2238,N_2108);
xnor U11219 (N_11219,N_1588,N_1898);
and U11220 (N_11220,N_5606,N_5675);
and U11221 (N_11221,N_4405,N_1143);
and U11222 (N_11222,N_4782,N_321);
nand U11223 (N_11223,N_3331,N_1282);
or U11224 (N_11224,N_4725,N_2782);
and U11225 (N_11225,N_5902,N_1961);
nand U11226 (N_11226,N_2911,N_4354);
or U11227 (N_11227,N_5513,N_3552);
or U11228 (N_11228,N_948,N_1036);
and U11229 (N_11229,N_2001,N_1965);
and U11230 (N_11230,N_3133,N_107);
and U11231 (N_11231,N_3774,N_5764);
xor U11232 (N_11232,N_2563,N_3411);
nand U11233 (N_11233,N_3357,N_5571);
nand U11234 (N_11234,N_5721,N_286);
xor U11235 (N_11235,N_2302,N_3871);
and U11236 (N_11236,N_2196,N_1130);
or U11237 (N_11237,N_3702,N_1205);
and U11238 (N_11238,N_3331,N_2340);
or U11239 (N_11239,N_3002,N_492);
nand U11240 (N_11240,N_3035,N_5175);
xnor U11241 (N_11241,N_3013,N_2528);
and U11242 (N_11242,N_2508,N_3046);
nand U11243 (N_11243,N_5365,N_4713);
xor U11244 (N_11244,N_4568,N_4044);
nor U11245 (N_11245,N_814,N_2101);
and U11246 (N_11246,N_626,N_4410);
or U11247 (N_11247,N_3242,N_4714);
nand U11248 (N_11248,N_4486,N_4348);
or U11249 (N_11249,N_2941,N_5256);
nand U11250 (N_11250,N_4083,N_797);
nor U11251 (N_11251,N_2253,N_1601);
or U11252 (N_11252,N_438,N_1042);
and U11253 (N_11253,N_1279,N_3908);
nor U11254 (N_11254,N_499,N_4433);
and U11255 (N_11255,N_3778,N_115);
nand U11256 (N_11256,N_4165,N_892);
and U11257 (N_11257,N_2090,N_1591);
nand U11258 (N_11258,N_1014,N_388);
or U11259 (N_11259,N_1678,N_2);
and U11260 (N_11260,N_1075,N_5079);
nor U11261 (N_11261,N_3473,N_5731);
or U11262 (N_11262,N_5446,N_4567);
and U11263 (N_11263,N_3139,N_5964);
xor U11264 (N_11264,N_3545,N_3275);
nand U11265 (N_11265,N_150,N_2869);
nor U11266 (N_11266,N_1663,N_1693);
and U11267 (N_11267,N_3870,N_1804);
and U11268 (N_11268,N_1400,N_1331);
and U11269 (N_11269,N_3992,N_5157);
nor U11270 (N_11270,N_1567,N_2572);
nand U11271 (N_11271,N_1503,N_5389);
nand U11272 (N_11272,N_1494,N_4139);
or U11273 (N_11273,N_3990,N_1202);
nand U11274 (N_11274,N_5897,N_3035);
xnor U11275 (N_11275,N_205,N_3138);
nand U11276 (N_11276,N_2511,N_398);
nand U11277 (N_11277,N_562,N_5844);
and U11278 (N_11278,N_3090,N_357);
xnor U11279 (N_11279,N_2320,N_2339);
nand U11280 (N_11280,N_4697,N_4804);
xor U11281 (N_11281,N_455,N_2032);
nor U11282 (N_11282,N_5072,N_3292);
nor U11283 (N_11283,N_20,N_1602);
nor U11284 (N_11284,N_3822,N_5889);
and U11285 (N_11285,N_5460,N_4626);
nand U11286 (N_11286,N_2640,N_1193);
or U11287 (N_11287,N_3190,N_2347);
or U11288 (N_11288,N_1474,N_46);
nor U11289 (N_11289,N_3772,N_2846);
xnor U11290 (N_11290,N_3259,N_133);
nor U11291 (N_11291,N_3607,N_2825);
and U11292 (N_11292,N_4979,N_946);
nor U11293 (N_11293,N_450,N_1278);
xor U11294 (N_11294,N_4458,N_4679);
nand U11295 (N_11295,N_5023,N_3404);
nor U11296 (N_11296,N_577,N_4779);
and U11297 (N_11297,N_5522,N_1051);
nor U11298 (N_11298,N_88,N_865);
and U11299 (N_11299,N_5655,N_461);
nor U11300 (N_11300,N_972,N_3503);
and U11301 (N_11301,N_3600,N_2406);
nor U11302 (N_11302,N_208,N_4917);
xnor U11303 (N_11303,N_2740,N_2732);
nor U11304 (N_11304,N_34,N_4895);
nand U11305 (N_11305,N_3291,N_4895);
and U11306 (N_11306,N_4098,N_253);
xnor U11307 (N_11307,N_5910,N_185);
or U11308 (N_11308,N_5949,N_1817);
and U11309 (N_11309,N_1740,N_184);
xor U11310 (N_11310,N_3539,N_5630);
nand U11311 (N_11311,N_5994,N_4019);
nor U11312 (N_11312,N_1796,N_4303);
and U11313 (N_11313,N_558,N_1477);
or U11314 (N_11314,N_3313,N_5370);
nor U11315 (N_11315,N_1646,N_1287);
nand U11316 (N_11316,N_973,N_3366);
nor U11317 (N_11317,N_1228,N_1334);
or U11318 (N_11318,N_4188,N_129);
xnor U11319 (N_11319,N_1841,N_1256);
or U11320 (N_11320,N_3551,N_4204);
and U11321 (N_11321,N_3213,N_3345);
nor U11322 (N_11322,N_219,N_3573);
or U11323 (N_11323,N_1946,N_4526);
nor U11324 (N_11324,N_1840,N_2331);
or U11325 (N_11325,N_3433,N_5918);
and U11326 (N_11326,N_3800,N_1431);
or U11327 (N_11327,N_4935,N_3812);
and U11328 (N_11328,N_4135,N_743);
nor U11329 (N_11329,N_2144,N_5843);
xnor U11330 (N_11330,N_1686,N_4896);
or U11331 (N_11331,N_5830,N_1174);
or U11332 (N_11332,N_1965,N_2273);
and U11333 (N_11333,N_2219,N_411);
or U11334 (N_11334,N_3471,N_353);
and U11335 (N_11335,N_4266,N_420);
or U11336 (N_11336,N_1293,N_1247);
and U11337 (N_11337,N_2922,N_3749);
nand U11338 (N_11338,N_2886,N_4237);
nor U11339 (N_11339,N_4040,N_3172);
xor U11340 (N_11340,N_1571,N_2284);
and U11341 (N_11341,N_2986,N_5472);
nand U11342 (N_11342,N_3457,N_3884);
and U11343 (N_11343,N_5981,N_3369);
or U11344 (N_11344,N_1150,N_5706);
and U11345 (N_11345,N_5493,N_4331);
nor U11346 (N_11346,N_658,N_3366);
and U11347 (N_11347,N_2537,N_2096);
or U11348 (N_11348,N_350,N_4219);
nor U11349 (N_11349,N_1606,N_3000);
xnor U11350 (N_11350,N_5367,N_14);
or U11351 (N_11351,N_2300,N_5102);
nand U11352 (N_11352,N_974,N_5423);
nand U11353 (N_11353,N_4083,N_1738);
nand U11354 (N_11354,N_5028,N_4722);
and U11355 (N_11355,N_1846,N_5122);
nor U11356 (N_11356,N_223,N_5022);
xnor U11357 (N_11357,N_2430,N_5943);
nor U11358 (N_11358,N_1892,N_5155);
or U11359 (N_11359,N_1775,N_2357);
nor U11360 (N_11360,N_5489,N_5368);
or U11361 (N_11361,N_2544,N_5581);
nor U11362 (N_11362,N_2396,N_418);
nand U11363 (N_11363,N_1272,N_4216);
and U11364 (N_11364,N_2024,N_4366);
and U11365 (N_11365,N_1209,N_5335);
xnor U11366 (N_11366,N_3055,N_3029);
or U11367 (N_11367,N_4308,N_4503);
or U11368 (N_11368,N_2064,N_1408);
or U11369 (N_11369,N_480,N_700);
and U11370 (N_11370,N_3118,N_2326);
nor U11371 (N_11371,N_1187,N_4340);
xor U11372 (N_11372,N_520,N_1544);
and U11373 (N_11373,N_3965,N_3791);
and U11374 (N_11374,N_2642,N_5229);
nand U11375 (N_11375,N_1123,N_4127);
nand U11376 (N_11376,N_2241,N_878);
nand U11377 (N_11377,N_2883,N_445);
or U11378 (N_11378,N_1055,N_4251);
and U11379 (N_11379,N_3293,N_5837);
nor U11380 (N_11380,N_2599,N_1633);
nand U11381 (N_11381,N_5760,N_5301);
or U11382 (N_11382,N_2472,N_4375);
xnor U11383 (N_11383,N_3378,N_5728);
or U11384 (N_11384,N_4501,N_5278);
nand U11385 (N_11385,N_1088,N_386);
or U11386 (N_11386,N_4086,N_5311);
and U11387 (N_11387,N_3878,N_4179);
xnor U11388 (N_11388,N_2699,N_3822);
nand U11389 (N_11389,N_3366,N_4978);
xor U11390 (N_11390,N_4803,N_2148);
nand U11391 (N_11391,N_4334,N_3289);
xnor U11392 (N_11392,N_3443,N_4818);
xnor U11393 (N_11393,N_4935,N_4917);
nor U11394 (N_11394,N_1317,N_5384);
nor U11395 (N_11395,N_4712,N_1620);
nor U11396 (N_11396,N_2385,N_1087);
nor U11397 (N_11397,N_3598,N_4947);
nor U11398 (N_11398,N_4749,N_3358);
xnor U11399 (N_11399,N_1430,N_2252);
xor U11400 (N_11400,N_5988,N_3358);
xor U11401 (N_11401,N_1540,N_397);
and U11402 (N_11402,N_1201,N_5749);
and U11403 (N_11403,N_4665,N_3114);
and U11404 (N_11404,N_3156,N_4723);
xnor U11405 (N_11405,N_1482,N_78);
nor U11406 (N_11406,N_1816,N_2283);
or U11407 (N_11407,N_5998,N_705);
and U11408 (N_11408,N_5724,N_775);
xnor U11409 (N_11409,N_4331,N_369);
or U11410 (N_11410,N_751,N_5221);
nor U11411 (N_11411,N_3239,N_3752);
nand U11412 (N_11412,N_2238,N_2107);
xor U11413 (N_11413,N_1827,N_906);
nand U11414 (N_11414,N_5775,N_4543);
or U11415 (N_11415,N_5933,N_1893);
or U11416 (N_11416,N_2503,N_1926);
nand U11417 (N_11417,N_3284,N_4134);
nand U11418 (N_11418,N_1649,N_1348);
and U11419 (N_11419,N_1443,N_1338);
nand U11420 (N_11420,N_3748,N_2504);
xnor U11421 (N_11421,N_3604,N_5478);
xnor U11422 (N_11422,N_2123,N_4246);
and U11423 (N_11423,N_5269,N_300);
or U11424 (N_11424,N_3806,N_414);
nor U11425 (N_11425,N_5362,N_1571);
nor U11426 (N_11426,N_1250,N_438);
or U11427 (N_11427,N_443,N_3362);
and U11428 (N_11428,N_3216,N_754);
nand U11429 (N_11429,N_1443,N_758);
or U11430 (N_11430,N_3764,N_3942);
and U11431 (N_11431,N_3059,N_5925);
and U11432 (N_11432,N_350,N_4390);
or U11433 (N_11433,N_1431,N_4007);
or U11434 (N_11434,N_2499,N_1540);
or U11435 (N_11435,N_830,N_4036);
and U11436 (N_11436,N_5849,N_5378);
or U11437 (N_11437,N_2899,N_2132);
nor U11438 (N_11438,N_4910,N_5614);
or U11439 (N_11439,N_1448,N_4531);
nand U11440 (N_11440,N_1886,N_216);
and U11441 (N_11441,N_392,N_5144);
and U11442 (N_11442,N_4702,N_4089);
and U11443 (N_11443,N_1299,N_828);
xnor U11444 (N_11444,N_3613,N_935);
nor U11445 (N_11445,N_888,N_895);
nor U11446 (N_11446,N_5427,N_2613);
nand U11447 (N_11447,N_3821,N_314);
nor U11448 (N_11448,N_1269,N_5876);
nor U11449 (N_11449,N_2391,N_4698);
and U11450 (N_11450,N_1893,N_4914);
nand U11451 (N_11451,N_3823,N_1734);
or U11452 (N_11452,N_3778,N_1649);
or U11453 (N_11453,N_1298,N_5603);
nand U11454 (N_11454,N_2910,N_3746);
nor U11455 (N_11455,N_2066,N_2522);
and U11456 (N_11456,N_5386,N_5846);
or U11457 (N_11457,N_1532,N_4851);
nor U11458 (N_11458,N_556,N_909);
and U11459 (N_11459,N_3292,N_5678);
and U11460 (N_11460,N_5075,N_4408);
xor U11461 (N_11461,N_3277,N_3662);
nor U11462 (N_11462,N_3070,N_3566);
and U11463 (N_11463,N_4331,N_3456);
or U11464 (N_11464,N_2339,N_5824);
xor U11465 (N_11465,N_4006,N_5504);
and U11466 (N_11466,N_4363,N_2834);
and U11467 (N_11467,N_2803,N_1281);
or U11468 (N_11468,N_2177,N_1711);
nand U11469 (N_11469,N_4946,N_2206);
and U11470 (N_11470,N_4137,N_5811);
nor U11471 (N_11471,N_4501,N_5836);
nor U11472 (N_11472,N_4568,N_2127);
xor U11473 (N_11473,N_3046,N_1627);
or U11474 (N_11474,N_4777,N_2968);
or U11475 (N_11475,N_489,N_2177);
and U11476 (N_11476,N_3862,N_4016);
nor U11477 (N_11477,N_2715,N_1401);
nand U11478 (N_11478,N_968,N_3966);
or U11479 (N_11479,N_1832,N_4946);
or U11480 (N_11480,N_31,N_1707);
nand U11481 (N_11481,N_1908,N_3074);
xor U11482 (N_11482,N_774,N_2453);
nor U11483 (N_11483,N_3343,N_4061);
or U11484 (N_11484,N_3565,N_2558);
nand U11485 (N_11485,N_1813,N_1056);
nor U11486 (N_11486,N_1230,N_1511);
and U11487 (N_11487,N_3157,N_3492);
or U11488 (N_11488,N_1164,N_3185);
and U11489 (N_11489,N_1259,N_3135);
nor U11490 (N_11490,N_192,N_2199);
or U11491 (N_11491,N_166,N_1828);
or U11492 (N_11492,N_4849,N_256);
and U11493 (N_11493,N_1415,N_4219);
or U11494 (N_11494,N_4050,N_4011);
xor U11495 (N_11495,N_1160,N_1882);
nand U11496 (N_11496,N_2508,N_4427);
and U11497 (N_11497,N_5689,N_2463);
nand U11498 (N_11498,N_1648,N_5612);
nand U11499 (N_11499,N_4800,N_2298);
nor U11500 (N_11500,N_2889,N_1743);
and U11501 (N_11501,N_4681,N_4842);
nor U11502 (N_11502,N_3719,N_5831);
or U11503 (N_11503,N_908,N_2110);
and U11504 (N_11504,N_3212,N_3615);
nand U11505 (N_11505,N_940,N_4166);
nor U11506 (N_11506,N_5780,N_4108);
xor U11507 (N_11507,N_2776,N_2324);
and U11508 (N_11508,N_4260,N_2382);
xor U11509 (N_11509,N_4039,N_466);
nor U11510 (N_11510,N_3451,N_3401);
and U11511 (N_11511,N_352,N_1007);
or U11512 (N_11512,N_2826,N_157);
or U11513 (N_11513,N_5470,N_650);
and U11514 (N_11514,N_2925,N_714);
and U11515 (N_11515,N_1400,N_3862);
nor U11516 (N_11516,N_639,N_3243);
xnor U11517 (N_11517,N_2717,N_4099);
nand U11518 (N_11518,N_1957,N_1361);
or U11519 (N_11519,N_1641,N_513);
nor U11520 (N_11520,N_2476,N_5517);
nor U11521 (N_11521,N_832,N_2108);
nand U11522 (N_11522,N_4999,N_985);
nand U11523 (N_11523,N_4926,N_1899);
and U11524 (N_11524,N_90,N_5692);
or U11525 (N_11525,N_5477,N_3033);
and U11526 (N_11526,N_5362,N_3880);
nor U11527 (N_11527,N_5030,N_732);
or U11528 (N_11528,N_5608,N_4194);
nor U11529 (N_11529,N_3304,N_2395);
or U11530 (N_11530,N_2844,N_1184);
nor U11531 (N_11531,N_5407,N_655);
xnor U11532 (N_11532,N_1339,N_2261);
nand U11533 (N_11533,N_4613,N_509);
or U11534 (N_11534,N_5146,N_1573);
and U11535 (N_11535,N_1032,N_2281);
nor U11536 (N_11536,N_5914,N_2238);
xor U11537 (N_11537,N_4253,N_3572);
and U11538 (N_11538,N_53,N_5349);
nand U11539 (N_11539,N_1525,N_2688);
or U11540 (N_11540,N_5895,N_3753);
nand U11541 (N_11541,N_3190,N_5650);
nor U11542 (N_11542,N_3693,N_3805);
nor U11543 (N_11543,N_624,N_2038);
nand U11544 (N_11544,N_1640,N_1905);
xnor U11545 (N_11545,N_3089,N_5871);
nand U11546 (N_11546,N_4687,N_475);
nand U11547 (N_11547,N_5270,N_4017);
nand U11548 (N_11548,N_1248,N_1522);
nor U11549 (N_11549,N_2504,N_4704);
nor U11550 (N_11550,N_5061,N_2981);
or U11551 (N_11551,N_1388,N_4495);
and U11552 (N_11552,N_648,N_3638);
nor U11553 (N_11553,N_5363,N_5954);
nand U11554 (N_11554,N_4449,N_3185);
nand U11555 (N_11555,N_138,N_4845);
nand U11556 (N_11556,N_3917,N_3585);
nand U11557 (N_11557,N_2303,N_3302);
nand U11558 (N_11558,N_2961,N_5314);
and U11559 (N_11559,N_4257,N_5754);
or U11560 (N_11560,N_2351,N_5855);
or U11561 (N_11561,N_3405,N_5319);
or U11562 (N_11562,N_475,N_4963);
nor U11563 (N_11563,N_314,N_270);
nand U11564 (N_11564,N_539,N_703);
or U11565 (N_11565,N_5433,N_5656);
nand U11566 (N_11566,N_5377,N_1179);
nand U11567 (N_11567,N_978,N_307);
or U11568 (N_11568,N_1873,N_3388);
and U11569 (N_11569,N_337,N_1495);
nor U11570 (N_11570,N_2391,N_5799);
or U11571 (N_11571,N_3048,N_2403);
or U11572 (N_11572,N_3587,N_4482);
xor U11573 (N_11573,N_5413,N_4513);
nor U11574 (N_11574,N_5213,N_519);
nor U11575 (N_11575,N_3219,N_5981);
or U11576 (N_11576,N_1546,N_5027);
or U11577 (N_11577,N_4673,N_2198);
and U11578 (N_11578,N_5866,N_2116);
and U11579 (N_11579,N_5810,N_5391);
or U11580 (N_11580,N_4768,N_1610);
or U11581 (N_11581,N_833,N_2561);
nand U11582 (N_11582,N_1858,N_4553);
nand U11583 (N_11583,N_1901,N_3352);
and U11584 (N_11584,N_2683,N_5370);
and U11585 (N_11585,N_4679,N_5903);
and U11586 (N_11586,N_3973,N_279);
nand U11587 (N_11587,N_3169,N_4752);
and U11588 (N_11588,N_4439,N_631);
nor U11589 (N_11589,N_3731,N_2001);
and U11590 (N_11590,N_3336,N_321);
nand U11591 (N_11591,N_2184,N_5167);
nor U11592 (N_11592,N_1039,N_2761);
nor U11593 (N_11593,N_4427,N_524);
and U11594 (N_11594,N_3073,N_1610);
nor U11595 (N_11595,N_1562,N_3783);
or U11596 (N_11596,N_5609,N_4992);
and U11597 (N_11597,N_1042,N_4048);
nand U11598 (N_11598,N_4878,N_2465);
nand U11599 (N_11599,N_955,N_3170);
nand U11600 (N_11600,N_1835,N_4701);
or U11601 (N_11601,N_4861,N_548);
and U11602 (N_11602,N_3599,N_4238);
and U11603 (N_11603,N_1486,N_4295);
or U11604 (N_11604,N_254,N_3473);
nand U11605 (N_11605,N_2161,N_2913);
nand U11606 (N_11606,N_1047,N_2006);
nor U11607 (N_11607,N_4871,N_3235);
or U11608 (N_11608,N_1494,N_4483);
nand U11609 (N_11609,N_3499,N_845);
or U11610 (N_11610,N_5589,N_5061);
nand U11611 (N_11611,N_5338,N_4425);
or U11612 (N_11612,N_1216,N_2826);
nor U11613 (N_11613,N_2438,N_2191);
or U11614 (N_11614,N_808,N_5142);
nor U11615 (N_11615,N_3462,N_4913);
and U11616 (N_11616,N_797,N_357);
or U11617 (N_11617,N_391,N_4235);
nor U11618 (N_11618,N_2448,N_5591);
nand U11619 (N_11619,N_2294,N_4770);
and U11620 (N_11620,N_2694,N_4274);
xnor U11621 (N_11621,N_653,N_4763);
nand U11622 (N_11622,N_671,N_682);
nand U11623 (N_11623,N_1333,N_1109);
nor U11624 (N_11624,N_882,N_686);
or U11625 (N_11625,N_5296,N_1623);
nand U11626 (N_11626,N_5388,N_1891);
nand U11627 (N_11627,N_885,N_2243);
or U11628 (N_11628,N_862,N_1106);
and U11629 (N_11629,N_1424,N_3451);
and U11630 (N_11630,N_692,N_1209);
xor U11631 (N_11631,N_440,N_5397);
xor U11632 (N_11632,N_4497,N_182);
nor U11633 (N_11633,N_2199,N_583);
nor U11634 (N_11634,N_3559,N_2681);
xnor U11635 (N_11635,N_4490,N_660);
or U11636 (N_11636,N_5205,N_2174);
nor U11637 (N_11637,N_5008,N_5282);
nand U11638 (N_11638,N_3475,N_4922);
nand U11639 (N_11639,N_1378,N_4194);
and U11640 (N_11640,N_206,N_5185);
or U11641 (N_11641,N_4165,N_5694);
nor U11642 (N_11642,N_4008,N_5475);
and U11643 (N_11643,N_4172,N_2716);
and U11644 (N_11644,N_1758,N_2546);
or U11645 (N_11645,N_1237,N_5708);
nand U11646 (N_11646,N_2248,N_2797);
nor U11647 (N_11647,N_5853,N_3757);
nand U11648 (N_11648,N_2637,N_2598);
nand U11649 (N_11649,N_3566,N_5651);
nor U11650 (N_11650,N_2202,N_4608);
and U11651 (N_11651,N_5851,N_826);
or U11652 (N_11652,N_1585,N_5492);
and U11653 (N_11653,N_1495,N_2596);
nor U11654 (N_11654,N_3681,N_5220);
nand U11655 (N_11655,N_2307,N_5622);
and U11656 (N_11656,N_3003,N_2466);
or U11657 (N_11657,N_908,N_1834);
nor U11658 (N_11658,N_3276,N_3637);
xnor U11659 (N_11659,N_3895,N_1371);
and U11660 (N_11660,N_23,N_3916);
and U11661 (N_11661,N_2293,N_1787);
or U11662 (N_11662,N_602,N_5498);
and U11663 (N_11663,N_2810,N_1972);
nand U11664 (N_11664,N_5366,N_3922);
xor U11665 (N_11665,N_4675,N_3778);
nor U11666 (N_11666,N_4335,N_3299);
nand U11667 (N_11667,N_5935,N_926);
or U11668 (N_11668,N_5828,N_703);
and U11669 (N_11669,N_2732,N_1298);
or U11670 (N_11670,N_3894,N_918);
and U11671 (N_11671,N_5326,N_1531);
or U11672 (N_11672,N_899,N_3985);
xnor U11673 (N_11673,N_2997,N_2875);
and U11674 (N_11674,N_3908,N_789);
xnor U11675 (N_11675,N_5362,N_3023);
nor U11676 (N_11676,N_4296,N_3471);
nand U11677 (N_11677,N_1742,N_4155);
and U11678 (N_11678,N_2195,N_4901);
or U11679 (N_11679,N_4316,N_5902);
nand U11680 (N_11680,N_451,N_2463);
and U11681 (N_11681,N_3733,N_2525);
and U11682 (N_11682,N_1831,N_4777);
xor U11683 (N_11683,N_1766,N_5737);
and U11684 (N_11684,N_1131,N_1851);
and U11685 (N_11685,N_700,N_4908);
nor U11686 (N_11686,N_4435,N_1891);
or U11687 (N_11687,N_3759,N_539);
xor U11688 (N_11688,N_5622,N_775);
xor U11689 (N_11689,N_667,N_2492);
nor U11690 (N_11690,N_4708,N_5262);
xor U11691 (N_11691,N_678,N_5719);
nand U11692 (N_11692,N_2247,N_1911);
nand U11693 (N_11693,N_125,N_5204);
nand U11694 (N_11694,N_3030,N_4639);
nor U11695 (N_11695,N_882,N_879);
and U11696 (N_11696,N_2118,N_1668);
or U11697 (N_11697,N_409,N_2248);
and U11698 (N_11698,N_5473,N_4439);
xor U11699 (N_11699,N_780,N_862);
nor U11700 (N_11700,N_2950,N_2115);
nor U11701 (N_11701,N_2396,N_1997);
or U11702 (N_11702,N_3565,N_538);
nand U11703 (N_11703,N_3176,N_5228);
or U11704 (N_11704,N_228,N_5262);
nand U11705 (N_11705,N_2990,N_2200);
or U11706 (N_11706,N_4411,N_2921);
nand U11707 (N_11707,N_5545,N_1383);
and U11708 (N_11708,N_3954,N_928);
and U11709 (N_11709,N_672,N_471);
nand U11710 (N_11710,N_3353,N_5999);
or U11711 (N_11711,N_2310,N_2142);
and U11712 (N_11712,N_1128,N_300);
nor U11713 (N_11713,N_5550,N_1036);
nand U11714 (N_11714,N_2302,N_5351);
nor U11715 (N_11715,N_2975,N_4995);
and U11716 (N_11716,N_2980,N_844);
nand U11717 (N_11717,N_1246,N_1363);
nand U11718 (N_11718,N_4065,N_3583);
nand U11719 (N_11719,N_1718,N_2446);
and U11720 (N_11720,N_3948,N_4854);
nor U11721 (N_11721,N_2756,N_5554);
nand U11722 (N_11722,N_1186,N_1538);
and U11723 (N_11723,N_3593,N_2923);
nand U11724 (N_11724,N_259,N_1684);
nand U11725 (N_11725,N_723,N_4150);
nor U11726 (N_11726,N_4466,N_1375);
or U11727 (N_11727,N_4005,N_1689);
and U11728 (N_11728,N_813,N_2118);
xnor U11729 (N_11729,N_5194,N_3524);
nor U11730 (N_11730,N_2846,N_726);
nor U11731 (N_11731,N_1402,N_3410);
or U11732 (N_11732,N_4933,N_2603);
nor U11733 (N_11733,N_3428,N_4488);
and U11734 (N_11734,N_3486,N_4264);
nor U11735 (N_11735,N_2054,N_2742);
nand U11736 (N_11736,N_3186,N_3507);
and U11737 (N_11737,N_1564,N_3775);
and U11738 (N_11738,N_5862,N_2575);
nand U11739 (N_11739,N_2457,N_4074);
or U11740 (N_11740,N_3363,N_3102);
xor U11741 (N_11741,N_4333,N_4759);
or U11742 (N_11742,N_1760,N_1264);
nand U11743 (N_11743,N_1962,N_1471);
nor U11744 (N_11744,N_195,N_5513);
or U11745 (N_11745,N_1877,N_1254);
or U11746 (N_11746,N_3746,N_352);
nand U11747 (N_11747,N_2751,N_393);
and U11748 (N_11748,N_2211,N_1886);
and U11749 (N_11749,N_1416,N_5598);
and U11750 (N_11750,N_1707,N_2905);
and U11751 (N_11751,N_5266,N_5008);
nor U11752 (N_11752,N_1464,N_5252);
or U11753 (N_11753,N_3014,N_3565);
and U11754 (N_11754,N_1497,N_2057);
nand U11755 (N_11755,N_3121,N_2770);
xor U11756 (N_11756,N_280,N_1191);
xnor U11757 (N_11757,N_2244,N_2037);
or U11758 (N_11758,N_2690,N_87);
xnor U11759 (N_11759,N_1351,N_4338);
and U11760 (N_11760,N_4540,N_711);
and U11761 (N_11761,N_2848,N_5908);
nor U11762 (N_11762,N_2425,N_3080);
nand U11763 (N_11763,N_5665,N_5581);
nor U11764 (N_11764,N_2373,N_1187);
nor U11765 (N_11765,N_633,N_5674);
nand U11766 (N_11766,N_2335,N_2149);
or U11767 (N_11767,N_5862,N_1269);
xnor U11768 (N_11768,N_5434,N_1451);
nor U11769 (N_11769,N_2227,N_3939);
nand U11770 (N_11770,N_5507,N_4327);
nand U11771 (N_11771,N_4760,N_724);
xnor U11772 (N_11772,N_4465,N_2863);
and U11773 (N_11773,N_1177,N_2546);
nor U11774 (N_11774,N_4711,N_2865);
and U11775 (N_11775,N_2186,N_1815);
nor U11776 (N_11776,N_1613,N_5884);
nor U11777 (N_11777,N_2419,N_1925);
nor U11778 (N_11778,N_876,N_4920);
nand U11779 (N_11779,N_4042,N_3365);
xor U11780 (N_11780,N_1291,N_4255);
or U11781 (N_11781,N_5042,N_4037);
nor U11782 (N_11782,N_3417,N_1064);
and U11783 (N_11783,N_2686,N_1411);
nor U11784 (N_11784,N_3118,N_2637);
nand U11785 (N_11785,N_2971,N_4394);
nor U11786 (N_11786,N_212,N_1495);
nor U11787 (N_11787,N_2784,N_220);
and U11788 (N_11788,N_1751,N_3267);
nand U11789 (N_11789,N_1148,N_1182);
nor U11790 (N_11790,N_976,N_2507);
nor U11791 (N_11791,N_1757,N_293);
or U11792 (N_11792,N_3882,N_1622);
and U11793 (N_11793,N_5346,N_1366);
or U11794 (N_11794,N_4344,N_5148);
xor U11795 (N_11795,N_646,N_3534);
nand U11796 (N_11796,N_3379,N_4081);
or U11797 (N_11797,N_270,N_2650);
and U11798 (N_11798,N_5137,N_4540);
xnor U11799 (N_11799,N_5138,N_5258);
nand U11800 (N_11800,N_3932,N_566);
nor U11801 (N_11801,N_1387,N_3988);
nor U11802 (N_11802,N_1534,N_2052);
nor U11803 (N_11803,N_3803,N_3589);
and U11804 (N_11804,N_1100,N_2270);
nor U11805 (N_11805,N_2465,N_5852);
xnor U11806 (N_11806,N_2748,N_5326);
nand U11807 (N_11807,N_3747,N_4159);
nand U11808 (N_11808,N_2868,N_4674);
and U11809 (N_11809,N_1900,N_5325);
or U11810 (N_11810,N_4841,N_5883);
nor U11811 (N_11811,N_4538,N_1423);
nor U11812 (N_11812,N_3095,N_1748);
and U11813 (N_11813,N_3582,N_1274);
nor U11814 (N_11814,N_2646,N_670);
nand U11815 (N_11815,N_4312,N_5137);
nor U11816 (N_11816,N_2396,N_125);
and U11817 (N_11817,N_4229,N_2476);
or U11818 (N_11818,N_5241,N_5939);
and U11819 (N_11819,N_3115,N_5217);
nand U11820 (N_11820,N_4301,N_5324);
nand U11821 (N_11821,N_3255,N_3449);
xor U11822 (N_11822,N_2167,N_624);
nand U11823 (N_11823,N_4447,N_790);
and U11824 (N_11824,N_3315,N_5184);
nand U11825 (N_11825,N_1108,N_153);
nor U11826 (N_11826,N_5557,N_2673);
nand U11827 (N_11827,N_5476,N_1932);
and U11828 (N_11828,N_2561,N_5360);
or U11829 (N_11829,N_721,N_5171);
nor U11830 (N_11830,N_3031,N_5001);
xnor U11831 (N_11831,N_5938,N_5868);
and U11832 (N_11832,N_5288,N_5148);
nand U11833 (N_11833,N_235,N_2536);
or U11834 (N_11834,N_5612,N_3362);
nor U11835 (N_11835,N_3076,N_1011);
and U11836 (N_11836,N_2514,N_2127);
nor U11837 (N_11837,N_599,N_1713);
nor U11838 (N_11838,N_4580,N_1516);
and U11839 (N_11839,N_3473,N_3358);
and U11840 (N_11840,N_438,N_1755);
nand U11841 (N_11841,N_2520,N_948);
or U11842 (N_11842,N_734,N_4547);
and U11843 (N_11843,N_3227,N_1003);
or U11844 (N_11844,N_287,N_2624);
xor U11845 (N_11845,N_3350,N_2543);
and U11846 (N_11846,N_1816,N_5738);
nor U11847 (N_11847,N_5276,N_3139);
or U11848 (N_11848,N_230,N_5994);
and U11849 (N_11849,N_5060,N_3949);
or U11850 (N_11850,N_1072,N_2448);
nor U11851 (N_11851,N_4289,N_1791);
nand U11852 (N_11852,N_4007,N_4272);
and U11853 (N_11853,N_2032,N_3354);
nand U11854 (N_11854,N_1809,N_3982);
or U11855 (N_11855,N_2409,N_3086);
and U11856 (N_11856,N_1729,N_5812);
or U11857 (N_11857,N_629,N_1710);
and U11858 (N_11858,N_1293,N_4004);
xnor U11859 (N_11859,N_3392,N_2523);
or U11860 (N_11860,N_4064,N_3235);
nor U11861 (N_11861,N_4980,N_964);
nand U11862 (N_11862,N_4024,N_2992);
or U11863 (N_11863,N_2886,N_1655);
or U11864 (N_11864,N_1960,N_2543);
nor U11865 (N_11865,N_4950,N_4313);
nand U11866 (N_11866,N_3034,N_4616);
nand U11867 (N_11867,N_5827,N_3058);
and U11868 (N_11868,N_605,N_4569);
nand U11869 (N_11869,N_3671,N_2461);
and U11870 (N_11870,N_3260,N_4990);
or U11871 (N_11871,N_4426,N_1846);
nand U11872 (N_11872,N_1586,N_341);
nor U11873 (N_11873,N_2463,N_639);
or U11874 (N_11874,N_5120,N_299);
nor U11875 (N_11875,N_3684,N_5008);
and U11876 (N_11876,N_2447,N_3044);
nor U11877 (N_11877,N_4980,N_3845);
nand U11878 (N_11878,N_1543,N_3094);
xor U11879 (N_11879,N_2689,N_2571);
nor U11880 (N_11880,N_1216,N_5184);
or U11881 (N_11881,N_5915,N_3237);
nor U11882 (N_11882,N_4810,N_3680);
and U11883 (N_11883,N_4374,N_1100);
nand U11884 (N_11884,N_3446,N_2348);
nand U11885 (N_11885,N_1599,N_730);
nand U11886 (N_11886,N_4840,N_1617);
nor U11887 (N_11887,N_2140,N_4028);
or U11888 (N_11888,N_4060,N_2561);
nor U11889 (N_11889,N_2192,N_413);
nor U11890 (N_11890,N_3473,N_521);
and U11891 (N_11891,N_1126,N_3632);
nand U11892 (N_11892,N_5401,N_5932);
xor U11893 (N_11893,N_4238,N_2452);
nor U11894 (N_11894,N_5271,N_144);
or U11895 (N_11895,N_4052,N_5721);
or U11896 (N_11896,N_4172,N_5182);
and U11897 (N_11897,N_5284,N_5750);
and U11898 (N_11898,N_2097,N_822);
nand U11899 (N_11899,N_1066,N_4537);
nand U11900 (N_11900,N_4703,N_2932);
nand U11901 (N_11901,N_2647,N_448);
and U11902 (N_11902,N_2086,N_633);
and U11903 (N_11903,N_487,N_2426);
nand U11904 (N_11904,N_1634,N_4384);
xnor U11905 (N_11905,N_5401,N_5200);
and U11906 (N_11906,N_514,N_3740);
or U11907 (N_11907,N_5916,N_2573);
nand U11908 (N_11908,N_2974,N_2522);
and U11909 (N_11909,N_5924,N_4194);
nor U11910 (N_11910,N_3231,N_3917);
nor U11911 (N_11911,N_2191,N_1760);
nand U11912 (N_11912,N_3409,N_1354);
nand U11913 (N_11913,N_1232,N_2314);
and U11914 (N_11914,N_4260,N_4703);
xor U11915 (N_11915,N_1476,N_685);
xor U11916 (N_11916,N_749,N_600);
xor U11917 (N_11917,N_3268,N_2239);
nor U11918 (N_11918,N_3861,N_3256);
nand U11919 (N_11919,N_2907,N_5055);
nor U11920 (N_11920,N_2490,N_1921);
or U11921 (N_11921,N_5510,N_3788);
and U11922 (N_11922,N_4102,N_256);
and U11923 (N_11923,N_1404,N_5741);
and U11924 (N_11924,N_812,N_3005);
nand U11925 (N_11925,N_3472,N_4899);
or U11926 (N_11926,N_903,N_5556);
xnor U11927 (N_11927,N_5013,N_937);
nand U11928 (N_11928,N_388,N_3441);
and U11929 (N_11929,N_558,N_5294);
nor U11930 (N_11930,N_3401,N_5999);
and U11931 (N_11931,N_5767,N_3067);
nand U11932 (N_11932,N_478,N_625);
nand U11933 (N_11933,N_4956,N_3368);
and U11934 (N_11934,N_4671,N_2902);
or U11935 (N_11935,N_5171,N_3575);
and U11936 (N_11936,N_3433,N_2385);
and U11937 (N_11937,N_2124,N_5374);
nor U11938 (N_11938,N_162,N_1649);
or U11939 (N_11939,N_2088,N_3763);
nor U11940 (N_11940,N_5864,N_812);
nand U11941 (N_11941,N_334,N_4837);
and U11942 (N_11942,N_2249,N_5182);
and U11943 (N_11943,N_2403,N_2105);
xnor U11944 (N_11944,N_2686,N_4483);
and U11945 (N_11945,N_1090,N_5626);
nand U11946 (N_11946,N_260,N_3470);
or U11947 (N_11947,N_732,N_2246);
or U11948 (N_11948,N_5149,N_4402);
nor U11949 (N_11949,N_3373,N_4069);
and U11950 (N_11950,N_3869,N_5607);
nand U11951 (N_11951,N_300,N_5953);
nand U11952 (N_11952,N_955,N_661);
nand U11953 (N_11953,N_5795,N_4286);
nand U11954 (N_11954,N_4896,N_3204);
and U11955 (N_11955,N_4165,N_4134);
nor U11956 (N_11956,N_5534,N_1441);
or U11957 (N_11957,N_5172,N_5715);
nor U11958 (N_11958,N_4645,N_1394);
nor U11959 (N_11959,N_4051,N_2383);
nor U11960 (N_11960,N_3332,N_3968);
nand U11961 (N_11961,N_2742,N_316);
xnor U11962 (N_11962,N_3459,N_226);
or U11963 (N_11963,N_2998,N_5035);
and U11964 (N_11964,N_349,N_5446);
nand U11965 (N_11965,N_4253,N_5374);
or U11966 (N_11966,N_3437,N_4766);
or U11967 (N_11967,N_5319,N_1902);
or U11968 (N_11968,N_4066,N_321);
or U11969 (N_11969,N_5596,N_4832);
nand U11970 (N_11970,N_2720,N_4356);
and U11971 (N_11971,N_4058,N_4442);
nor U11972 (N_11972,N_4055,N_1632);
and U11973 (N_11973,N_1557,N_2419);
nand U11974 (N_11974,N_1573,N_1321);
nor U11975 (N_11975,N_361,N_5723);
and U11976 (N_11976,N_3102,N_947);
nand U11977 (N_11977,N_4573,N_2800);
nand U11978 (N_11978,N_1863,N_5903);
or U11979 (N_11979,N_5016,N_2352);
nand U11980 (N_11980,N_1571,N_5400);
nand U11981 (N_11981,N_3226,N_3010);
and U11982 (N_11982,N_1432,N_954);
and U11983 (N_11983,N_3465,N_5989);
or U11984 (N_11984,N_2898,N_2498);
nor U11985 (N_11985,N_372,N_139);
nor U11986 (N_11986,N_4146,N_2481);
nand U11987 (N_11987,N_2822,N_1046);
nand U11988 (N_11988,N_5195,N_2397);
or U11989 (N_11989,N_908,N_448);
nand U11990 (N_11990,N_1219,N_651);
nand U11991 (N_11991,N_3327,N_5325);
nor U11992 (N_11992,N_3880,N_5962);
or U11993 (N_11993,N_63,N_2905);
nand U11994 (N_11994,N_1733,N_710);
and U11995 (N_11995,N_4296,N_5623);
xnor U11996 (N_11996,N_5212,N_2515);
and U11997 (N_11997,N_1432,N_2094);
and U11998 (N_11998,N_1958,N_3158);
and U11999 (N_11999,N_1244,N_1370);
or U12000 (N_12000,N_7195,N_9426);
nor U12001 (N_12001,N_11937,N_9485);
or U12002 (N_12002,N_10183,N_9462);
and U12003 (N_12003,N_10250,N_8999);
nor U12004 (N_12004,N_10205,N_9716);
nor U12005 (N_12005,N_7849,N_8431);
and U12006 (N_12006,N_7880,N_6106);
or U12007 (N_12007,N_6493,N_11014);
nor U12008 (N_12008,N_7026,N_7708);
and U12009 (N_12009,N_7683,N_7095);
or U12010 (N_12010,N_10115,N_9264);
xnor U12011 (N_12011,N_10261,N_8923);
nand U12012 (N_12012,N_7379,N_7561);
xnor U12013 (N_12013,N_9576,N_11095);
nand U12014 (N_12014,N_8264,N_8505);
xor U12015 (N_12015,N_6701,N_8063);
nor U12016 (N_12016,N_10876,N_6559);
nor U12017 (N_12017,N_10139,N_10248);
nor U12018 (N_12018,N_6786,N_9945);
and U12019 (N_12019,N_8219,N_7784);
xor U12020 (N_12020,N_7121,N_6274);
and U12021 (N_12021,N_7721,N_10522);
xor U12022 (N_12022,N_10993,N_10703);
and U12023 (N_12023,N_8201,N_9282);
or U12024 (N_12024,N_10288,N_9536);
nand U12025 (N_12025,N_7272,N_11549);
nand U12026 (N_12026,N_6119,N_8997);
or U12027 (N_12027,N_8274,N_8676);
nor U12028 (N_12028,N_8231,N_8159);
nor U12029 (N_12029,N_9567,N_7553);
nor U12030 (N_12030,N_8919,N_8446);
nor U12031 (N_12031,N_8820,N_7088);
nor U12032 (N_12032,N_11788,N_7404);
nand U12033 (N_12033,N_10696,N_11860);
nand U12034 (N_12034,N_10566,N_11565);
or U12035 (N_12035,N_10521,N_10832);
nor U12036 (N_12036,N_11468,N_7429);
and U12037 (N_12037,N_7521,N_7264);
nand U12038 (N_12038,N_10618,N_9774);
nor U12039 (N_12039,N_9408,N_8704);
nand U12040 (N_12040,N_9957,N_9074);
nand U12041 (N_12041,N_6341,N_10901);
and U12042 (N_12042,N_10594,N_7356);
nand U12043 (N_12043,N_10553,N_8612);
or U12044 (N_12044,N_8510,N_8598);
nand U12045 (N_12045,N_7948,N_9397);
nor U12046 (N_12046,N_7039,N_7777);
or U12047 (N_12047,N_8868,N_11787);
or U12048 (N_12048,N_8541,N_6367);
nor U12049 (N_12049,N_8358,N_6349);
nand U12050 (N_12050,N_6637,N_9985);
xnor U12051 (N_12051,N_6505,N_11581);
or U12052 (N_12052,N_9912,N_9891);
xnor U12053 (N_12053,N_9225,N_8353);
or U12054 (N_12054,N_8314,N_9978);
nor U12055 (N_12055,N_6915,N_6409);
nand U12056 (N_12056,N_8458,N_10933);
and U12057 (N_12057,N_8230,N_7203);
nor U12058 (N_12058,N_8879,N_6115);
nand U12059 (N_12059,N_6213,N_6183);
nor U12060 (N_12060,N_9318,N_9164);
xnor U12061 (N_12061,N_6821,N_9109);
and U12062 (N_12062,N_9234,N_11739);
and U12063 (N_12063,N_6765,N_9915);
xnor U12064 (N_12064,N_8572,N_6736);
and U12065 (N_12065,N_10887,N_10818);
nand U12066 (N_12066,N_7093,N_11365);
or U12067 (N_12067,N_7989,N_11381);
or U12068 (N_12068,N_8133,N_6908);
nor U12069 (N_12069,N_7641,N_8481);
nor U12070 (N_12070,N_8131,N_6297);
nand U12071 (N_12071,N_6798,N_11022);
and U12072 (N_12072,N_8989,N_11570);
nand U12073 (N_12073,N_11460,N_7858);
nand U12074 (N_12074,N_11312,N_9106);
xnor U12075 (N_12075,N_11723,N_9884);
nand U12076 (N_12076,N_8226,N_8398);
nor U12077 (N_12077,N_7148,N_11767);
and U12078 (N_12078,N_8801,N_6599);
nand U12079 (N_12079,N_6655,N_7586);
xor U12080 (N_12080,N_6249,N_10066);
xnor U12081 (N_12081,N_11169,N_11736);
nor U12082 (N_12082,N_11572,N_10264);
xor U12083 (N_12083,N_8733,N_9677);
or U12084 (N_12084,N_9243,N_11404);
and U12085 (N_12085,N_7211,N_9472);
and U12086 (N_12086,N_11828,N_11768);
or U12087 (N_12087,N_8134,N_10061);
or U12088 (N_12088,N_8176,N_6627);
or U12089 (N_12089,N_6377,N_9195);
nand U12090 (N_12090,N_10875,N_6280);
or U12091 (N_12091,N_7192,N_11817);
xor U12092 (N_12092,N_10171,N_8023);
nor U12093 (N_12093,N_7978,N_11651);
or U12094 (N_12094,N_8403,N_8544);
or U12095 (N_12095,N_10244,N_7454);
and U12096 (N_12096,N_11658,N_7924);
nor U12097 (N_12097,N_11420,N_6139);
or U12098 (N_12098,N_9003,N_6714);
nand U12099 (N_12099,N_10402,N_8401);
or U12100 (N_12100,N_10869,N_10807);
nand U12101 (N_12101,N_6430,N_11152);
nand U12102 (N_12102,N_6177,N_10358);
nand U12103 (N_12103,N_6404,N_11471);
nand U12104 (N_12104,N_7418,N_7218);
xnor U12105 (N_12105,N_8662,N_7073);
or U12106 (N_12106,N_10148,N_7347);
nand U12107 (N_12107,N_9664,N_11503);
nand U12108 (N_12108,N_8787,N_8035);
nand U12109 (N_12109,N_9876,N_6023);
nand U12110 (N_12110,N_8119,N_10483);
nand U12111 (N_12111,N_8764,N_10243);
nand U12112 (N_12112,N_11631,N_6232);
nand U12113 (N_12113,N_11431,N_6082);
and U12114 (N_12114,N_9505,N_6577);
nand U12115 (N_12115,N_6410,N_9517);
or U12116 (N_12116,N_10528,N_11488);
nand U12117 (N_12117,N_10740,N_10461);
nor U12118 (N_12118,N_8416,N_10071);
nand U12119 (N_12119,N_10502,N_6257);
or U12120 (N_12120,N_10544,N_7838);
or U12121 (N_12121,N_10761,N_6193);
nand U12122 (N_12122,N_8056,N_9378);
nand U12123 (N_12123,N_11469,N_9189);
xor U12124 (N_12124,N_8823,N_10043);
and U12125 (N_12125,N_9804,N_10806);
nor U12126 (N_12126,N_9489,N_10749);
nor U12127 (N_12127,N_7444,N_11305);
nor U12128 (N_12128,N_11345,N_8737);
nor U12129 (N_12129,N_10586,N_10101);
or U12130 (N_12130,N_10877,N_11567);
nor U12131 (N_12131,N_9638,N_11178);
xnor U12132 (N_12132,N_10515,N_8021);
and U12133 (N_12133,N_9337,N_6310);
and U12134 (N_12134,N_7932,N_6966);
nor U12135 (N_12135,N_6805,N_11222);
xnor U12136 (N_12136,N_6358,N_9077);
xnor U12137 (N_12137,N_8108,N_8836);
nand U12138 (N_12138,N_9269,N_8978);
and U12139 (N_12139,N_8773,N_9137);
nor U12140 (N_12140,N_7084,N_7290);
nor U12141 (N_12141,N_9019,N_10460);
and U12142 (N_12142,N_11956,N_8804);
xnor U12143 (N_12143,N_11368,N_9083);
nand U12144 (N_12144,N_10636,N_8635);
nand U12145 (N_12145,N_10425,N_11843);
nand U12146 (N_12146,N_9706,N_9032);
xor U12147 (N_12147,N_10282,N_6034);
nor U12148 (N_12148,N_10283,N_7531);
and U12149 (N_12149,N_10065,N_8560);
nor U12150 (N_12150,N_11976,N_10334);
or U12151 (N_12151,N_9231,N_6776);
nand U12152 (N_12152,N_11924,N_11329);
or U12153 (N_12153,N_10119,N_7548);
nand U12154 (N_12154,N_9709,N_7200);
nand U12155 (N_12155,N_11207,N_7149);
nor U12156 (N_12156,N_7054,N_6842);
or U12157 (N_12157,N_6059,N_8686);
nor U12158 (N_12158,N_11673,N_11000);
xor U12159 (N_12159,N_11752,N_7107);
and U12160 (N_12160,N_10359,N_6981);
nand U12161 (N_12161,N_11332,N_10622);
nand U12162 (N_12162,N_7297,N_6439);
or U12163 (N_12163,N_6450,N_7905);
and U12164 (N_12164,N_11445,N_8622);
xnor U12165 (N_12165,N_11142,N_11480);
nand U12166 (N_12166,N_6418,N_8513);
and U12167 (N_12167,N_11136,N_10078);
nand U12168 (N_12168,N_9056,N_9042);
nor U12169 (N_12169,N_6595,N_10547);
and U12170 (N_12170,N_11882,N_6866);
or U12171 (N_12171,N_10023,N_8586);
nand U12172 (N_12172,N_9655,N_6406);
xor U12173 (N_12173,N_9238,N_11234);
or U12174 (N_12174,N_7806,N_9220);
or U12175 (N_12175,N_9085,N_8750);
nand U12176 (N_12176,N_7856,N_9832);
or U12177 (N_12177,N_11680,N_6964);
and U12178 (N_12178,N_8433,N_7996);
nor U12179 (N_12179,N_10340,N_7086);
nand U12180 (N_12180,N_11848,N_11521);
nand U12181 (N_12181,N_11929,N_11738);
nand U12182 (N_12182,N_7308,N_8359);
nor U12183 (N_12183,N_6062,N_8752);
nor U12184 (N_12184,N_9806,N_9658);
nor U12185 (N_12185,N_6181,N_9261);
nor U12186 (N_12186,N_10388,N_9108);
or U12187 (N_12187,N_7434,N_10414);
nand U12188 (N_12188,N_8191,N_6510);
or U12189 (N_12189,N_9073,N_9105);
xor U12190 (N_12190,N_11449,N_9939);
and U12191 (N_12191,N_10542,N_10769);
and U12192 (N_12192,N_11316,N_6042);
nand U12193 (N_12193,N_10293,N_9969);
or U12194 (N_12194,N_9590,N_10439);
nand U12195 (N_12195,N_7529,N_10493);
and U12196 (N_12196,N_8435,N_10919);
xor U12197 (N_12197,N_9565,N_9508);
nor U12198 (N_12198,N_8066,N_6835);
nor U12199 (N_12199,N_9089,N_8708);
xor U12200 (N_12200,N_7333,N_7357);
nor U12201 (N_12201,N_11026,N_11705);
and U12202 (N_12202,N_8294,N_9786);
xnor U12203 (N_12203,N_11347,N_10382);
nand U12204 (N_12204,N_8471,N_7736);
nor U12205 (N_12205,N_6899,N_10986);
nand U12206 (N_12206,N_10182,N_7078);
or U12207 (N_12207,N_6465,N_9482);
and U12208 (N_12208,N_7921,N_6998);
nand U12209 (N_12209,N_6486,N_7768);
or U12210 (N_12210,N_8179,N_9368);
nand U12211 (N_12211,N_9280,N_9249);
nand U12212 (N_12212,N_9130,N_9864);
or U12213 (N_12213,N_10781,N_10565);
nor U12214 (N_12214,N_9200,N_11193);
or U12215 (N_12215,N_10891,N_11112);
and U12216 (N_12216,N_11247,N_11394);
xor U12217 (N_12217,N_8499,N_9589);
nor U12218 (N_12218,N_6861,N_9058);
and U12219 (N_12219,N_11831,N_10640);
and U12220 (N_12220,N_8805,N_9650);
nand U12221 (N_12221,N_6277,N_8731);
or U12222 (N_12222,N_8952,N_10489);
and U12223 (N_12223,N_7998,N_8852);
xnor U12224 (N_12224,N_10741,N_6803);
or U12225 (N_12225,N_8813,N_8188);
xnor U12226 (N_12226,N_8778,N_10600);
and U12227 (N_12227,N_11444,N_6693);
and U12228 (N_12228,N_9409,N_8116);
nor U12229 (N_12229,N_10820,N_10085);
or U12230 (N_12230,N_10910,N_10407);
nand U12231 (N_12231,N_10580,N_11300);
and U12232 (N_12232,N_7942,N_9393);
nand U12233 (N_12233,N_8751,N_7461);
nand U12234 (N_12234,N_6996,N_7786);
nand U12235 (N_12235,N_8740,N_11496);
or U12236 (N_12236,N_10159,N_6609);
and U12237 (N_12237,N_6057,N_7617);
xor U12238 (N_12238,N_6125,N_10231);
nor U12239 (N_12239,N_11890,N_7300);
or U12240 (N_12240,N_8365,N_8436);
nand U12241 (N_12241,N_9445,N_10755);
and U12242 (N_12242,N_7275,N_9268);
and U12243 (N_12243,N_9413,N_7817);
nand U12244 (N_12244,N_10177,N_11288);
nand U12245 (N_12245,N_9099,N_11157);
or U12246 (N_12246,N_7344,N_10911);
or U12247 (N_12247,N_9711,N_9104);
nand U12248 (N_12248,N_9325,N_8380);
or U12249 (N_12249,N_6596,N_7289);
and U12250 (N_12250,N_9687,N_7734);
or U12251 (N_12251,N_9155,N_11641);
nand U12252 (N_12252,N_6878,N_10338);
or U12253 (N_12253,N_10226,N_11561);
nand U12254 (N_12254,N_11183,N_7636);
and U12255 (N_12255,N_10691,N_7059);
or U12256 (N_12256,N_8067,N_9293);
nand U12257 (N_12257,N_6823,N_11746);
and U12258 (N_12258,N_6894,N_9097);
and U12259 (N_12259,N_7901,N_6101);
nor U12260 (N_12260,N_9792,N_10527);
nand U12261 (N_12261,N_10537,N_9983);
nor U12262 (N_12262,N_10039,N_11771);
and U12263 (N_12263,N_9849,N_6470);
nor U12264 (N_12264,N_6110,N_11683);
or U12265 (N_12265,N_9470,N_6551);
xnor U12266 (N_12266,N_11172,N_6635);
nor U12267 (N_12267,N_11814,N_6667);
nor U12268 (N_12268,N_11185,N_6585);
nor U12269 (N_12269,N_6931,N_6837);
or U12270 (N_12270,N_9053,N_9604);
nand U12271 (N_12271,N_11074,N_9525);
and U12272 (N_12272,N_8977,N_6905);
and U12273 (N_12273,N_6830,N_11210);
nor U12274 (N_12274,N_10627,N_9921);
nor U12275 (N_12275,N_8389,N_10325);
nand U12276 (N_12276,N_10568,N_9006);
xor U12277 (N_12277,N_11727,N_9784);
or U12278 (N_12278,N_6412,N_9815);
nand U12279 (N_12279,N_8162,N_8966);
nor U12280 (N_12280,N_11903,N_11416);
and U12281 (N_12281,N_9437,N_11064);
or U12282 (N_12282,N_8853,N_8603);
and U12283 (N_12283,N_7670,N_10849);
nand U12284 (N_12284,N_6018,N_10558);
nand U12285 (N_12285,N_8819,N_10585);
nor U12286 (N_12286,N_11295,N_10735);
and U12287 (N_12287,N_11912,N_9734);
nand U12288 (N_12288,N_6248,N_10042);
and U12289 (N_12289,N_11344,N_6888);
nand U12290 (N_12290,N_11248,N_9430);
nor U12291 (N_12291,N_8707,N_7615);
nor U12292 (N_12292,N_11686,N_11836);
nand U12293 (N_12293,N_7076,N_11273);
xnor U12294 (N_12294,N_7654,N_9093);
or U12295 (N_12295,N_6834,N_10736);
nand U12296 (N_12296,N_9350,N_6227);
nand U12297 (N_12297,N_10190,N_11379);
nand U12298 (N_12298,N_8307,N_6334);
nor U12299 (N_12299,N_8717,N_11459);
or U12300 (N_12300,N_6093,N_8734);
nor U12301 (N_12301,N_7585,N_6777);
xor U12302 (N_12302,N_9123,N_11684);
nand U12303 (N_12303,N_8838,N_8136);
or U12304 (N_12304,N_8525,N_6930);
nand U12305 (N_12305,N_6833,N_6729);
xnor U12306 (N_12306,N_8337,N_7433);
nor U12307 (N_12307,N_6376,N_11292);
xor U12308 (N_12308,N_9509,N_8799);
and U12309 (N_12309,N_11881,N_6258);
nand U12310 (N_12310,N_6600,N_7431);
and U12311 (N_12311,N_10559,N_6532);
nand U12312 (N_12312,N_8316,N_9214);
and U12313 (N_12313,N_9674,N_8908);
nand U12314 (N_12314,N_10518,N_6702);
nor U12315 (N_12315,N_11710,N_9451);
or U12316 (N_12316,N_8935,N_11199);
nand U12317 (N_12317,N_9323,N_8017);
nor U12318 (N_12318,N_10017,N_11714);
or U12319 (N_12319,N_8795,N_7367);
or U12320 (N_12320,N_7842,N_10034);
and U12321 (N_12321,N_8317,N_6766);
nand U12322 (N_12322,N_8284,N_9802);
xor U12323 (N_12323,N_10831,N_10700);
or U12324 (N_12324,N_8379,N_9889);
and U12325 (N_12325,N_9575,N_7396);
nor U12326 (N_12326,N_9668,N_7462);
or U12327 (N_12327,N_10929,N_6529);
or U12328 (N_12328,N_10912,N_8864);
nor U12329 (N_12329,N_6346,N_11729);
and U12330 (N_12330,N_6009,N_10092);
nor U12331 (N_12331,N_10643,N_11776);
or U12332 (N_12332,N_7523,N_7197);
or U12333 (N_12333,N_8049,N_11517);
xor U12334 (N_12334,N_7945,N_6983);
nor U12335 (N_12335,N_8798,N_9467);
or U12336 (N_12336,N_10630,N_11871);
and U12337 (N_12337,N_10884,N_7646);
and U12338 (N_12338,N_10984,N_7019);
nor U12339 (N_12339,N_6441,N_11889);
nand U12340 (N_12340,N_8865,N_8537);
or U12341 (N_12341,N_8509,N_7280);
nor U12342 (N_12342,N_8076,N_6162);
nor U12343 (N_12343,N_6684,N_7943);
nand U12344 (N_12344,N_10152,N_8096);
nand U12345 (N_12345,N_9663,N_10242);
xnor U12346 (N_12346,N_8959,N_11334);
or U12347 (N_12347,N_7231,N_11050);
or U12348 (N_12348,N_8894,N_11845);
and U12349 (N_12349,N_11424,N_8817);
or U12350 (N_12350,N_9580,N_11255);
nand U12351 (N_12351,N_7887,N_8183);
or U12352 (N_12352,N_10900,N_9890);
nand U12353 (N_12353,N_7601,N_7730);
and U12354 (N_12354,N_11827,N_7279);
and U12355 (N_12355,N_7335,N_11901);
nor U12356 (N_12356,N_9582,N_9086);
nand U12357 (N_12357,N_10913,N_11410);
or U12358 (N_12358,N_10145,N_10713);
and U12359 (N_12359,N_10698,N_9041);
and U12360 (N_12360,N_10567,N_8759);
or U12361 (N_12361,N_9007,N_8271);
or U12362 (N_12362,N_10975,N_8539);
nand U12363 (N_12363,N_6174,N_10644);
nor U12364 (N_12364,N_8042,N_7398);
and U12365 (N_12365,N_11585,N_11914);
and U12366 (N_12366,N_8618,N_9158);
xor U12367 (N_12367,N_7649,N_9847);
and U12368 (N_12368,N_8334,N_11508);
or U12369 (N_12369,N_11280,N_8289);
nor U12370 (N_12370,N_11932,N_6301);
and U12371 (N_12371,N_7602,N_11626);
nor U12372 (N_12372,N_8788,N_7268);
nor U12373 (N_12373,N_10130,N_11540);
or U12374 (N_12374,N_8600,N_9899);
nor U12375 (N_12375,N_10982,N_7976);
nor U12376 (N_12376,N_9017,N_11134);
nor U12377 (N_12377,N_8336,N_11337);
or U12378 (N_12378,N_6116,N_7815);
and U12379 (N_12379,N_6975,N_9321);
xnor U12380 (N_12380,N_10363,N_11021);
nand U12381 (N_12381,N_6306,N_10943);
or U12382 (N_12382,N_7684,N_10339);
nor U12383 (N_12383,N_9645,N_11063);
nand U12384 (N_12384,N_6380,N_10941);
xor U12385 (N_12385,N_10253,N_10480);
nor U12386 (N_12386,N_11451,N_10328);
nand U12387 (N_12387,N_9630,N_8472);
nor U12388 (N_12388,N_6845,N_9216);
or U12389 (N_12389,N_11245,N_9702);
xor U12390 (N_12390,N_7725,N_6758);
or U12391 (N_12391,N_8834,N_6628);
nand U12392 (N_12392,N_9692,N_11395);
and U12393 (N_12393,N_11171,N_11635);
nand U12394 (N_12394,N_10020,N_8246);
or U12395 (N_12395,N_6157,N_6658);
or U12396 (N_12396,N_11933,N_6391);
nand U12397 (N_12397,N_6282,N_7871);
and U12398 (N_12398,N_10847,N_10670);
nand U12399 (N_12399,N_7714,N_11114);
nand U12400 (N_12400,N_11622,N_9453);
nor U12401 (N_12401,N_9532,N_6171);
and U12402 (N_12402,N_8848,N_8442);
or U12403 (N_12403,N_9892,N_11243);
nand U12404 (N_12404,N_10470,N_8610);
or U12405 (N_12405,N_6168,N_10230);
or U12406 (N_12406,N_9193,N_6158);
nand U12407 (N_12407,N_11423,N_11818);
or U12408 (N_12408,N_9913,N_10526);
and U12409 (N_12409,N_8828,N_9643);
and U12410 (N_12410,N_6080,N_6800);
or U12411 (N_12411,N_10709,N_9064);
nor U12412 (N_12412,N_8151,N_10812);
nor U12413 (N_12413,N_7666,N_9499);
nor U12414 (N_12414,N_7388,N_11040);
and U12415 (N_12415,N_6746,N_11490);
and U12416 (N_12416,N_9324,N_7277);
and U12417 (N_12417,N_9637,N_7517);
nand U12418 (N_12418,N_11809,N_9241);
nand U12419 (N_12419,N_11556,N_10021);
and U12420 (N_12420,N_6856,N_7611);
and U12421 (N_12421,N_9274,N_10311);
nor U12422 (N_12422,N_9365,N_6241);
xnor U12423 (N_12423,N_9015,N_7514);
xor U12424 (N_12424,N_7669,N_7413);
xor U12425 (N_12425,N_6535,N_8248);
xor U12426 (N_12426,N_6104,N_6369);
nor U12427 (N_12427,N_7321,N_11801);
nor U12428 (N_12428,N_9036,N_10216);
or U12429 (N_12429,N_9551,N_11601);
or U12430 (N_12430,N_6732,N_6896);
nor U12431 (N_12431,N_9361,N_6753);
or U12432 (N_12432,N_8362,N_6913);
or U12433 (N_12433,N_7955,N_10990);
and U12434 (N_12434,N_7475,N_7037);
and U12435 (N_12435,N_8555,N_6849);
nor U12436 (N_12436,N_8546,N_9861);
nand U12437 (N_12437,N_7898,N_6809);
nand U12438 (N_12438,N_6933,N_11085);
and U12439 (N_12439,N_7574,N_7949);
or U12440 (N_12440,N_9528,N_11493);
nor U12441 (N_12441,N_8950,N_8187);
nor U12442 (N_12442,N_10004,N_11078);
or U12443 (N_12443,N_11502,N_10851);
or U12444 (N_12444,N_6760,N_7020);
or U12445 (N_12445,N_7099,N_7236);
or U12446 (N_12446,N_9483,N_8014);
or U12447 (N_12447,N_9809,N_9290);
nand U12448 (N_12448,N_11239,N_10077);
xor U12449 (N_12449,N_11665,N_10275);
nand U12450 (N_12450,N_8643,N_6173);
nor U12451 (N_12451,N_10886,N_10661);
and U12452 (N_12452,N_7828,N_7809);
xor U12453 (N_12453,N_8910,N_9340);
nor U12454 (N_12454,N_10676,N_8477);
or U12455 (N_12455,N_9735,N_10706);
or U12456 (N_12456,N_11175,N_7448);
and U12457 (N_12457,N_6957,N_7881);
nor U12458 (N_12458,N_7991,N_11458);
nand U12459 (N_12459,N_9870,N_9427);
and U12460 (N_12460,N_7349,N_10179);
nor U12461 (N_12461,N_11065,N_8711);
nor U12462 (N_12462,N_6457,N_9573);
nor U12463 (N_12463,N_8354,N_10380);
and U12464 (N_12464,N_10836,N_6133);
or U12465 (N_12465,N_11120,N_10906);
or U12466 (N_12466,N_11150,N_9068);
nor U12467 (N_12467,N_7052,N_7582);
nor U12468 (N_12468,N_6515,N_6621);
or U12469 (N_12469,N_10817,N_8140);
or U12470 (N_12470,N_8885,N_10333);
and U12471 (N_12471,N_8496,N_7629);
xor U12472 (N_12472,N_8969,N_9403);
nand U12473 (N_12473,N_11462,N_8459);
nand U12474 (N_12474,N_10464,N_7605);
and U12475 (N_12475,N_11392,N_10609);
nand U12476 (N_12476,N_11125,N_11256);
nor U12477 (N_12477,N_10729,N_10809);
nor U12478 (N_12478,N_7456,N_7940);
nand U12479 (N_12479,N_7464,N_7334);
or U12480 (N_12480,N_6016,N_11220);
or U12481 (N_12481,N_10685,N_7371);
nor U12482 (N_12482,N_8086,N_9132);
nand U12483 (N_12483,N_11760,N_8529);
nand U12484 (N_12484,N_10045,N_7747);
or U12485 (N_12485,N_6858,N_6978);
nand U12486 (N_12486,N_7745,N_9511);
and U12487 (N_12487,N_7458,N_11740);
and U12488 (N_12488,N_7159,N_8909);
and U12489 (N_12489,N_11587,N_10347);
and U12490 (N_12490,N_11548,N_10276);
and U12491 (N_12491,N_7801,N_6008);
or U12492 (N_12492,N_7535,N_7346);
or U12493 (N_12493,N_6206,N_10327);
or U12494 (N_12494,N_11061,N_9446);
nor U12495 (N_12495,N_9619,N_10165);
nor U12496 (N_12496,N_9315,N_10496);
or U12497 (N_12497,N_11005,N_9139);
and U12498 (N_12498,N_11266,N_10569);
xnor U12499 (N_12499,N_10263,N_11492);
nor U12500 (N_12500,N_6708,N_7697);
or U12501 (N_12501,N_7144,N_7511);
and U12502 (N_12502,N_7127,N_11780);
and U12503 (N_12503,N_10861,N_9946);
and U12504 (N_12504,N_8128,N_9418);
nand U12505 (N_12505,N_8774,N_8400);
and U12506 (N_12506,N_9829,N_8225);
or U12507 (N_12507,N_11741,N_8732);
or U12508 (N_12508,N_11749,N_9078);
nand U12509 (N_12509,N_8890,N_9987);
xnor U12510 (N_12510,N_7643,N_7519);
nor U12511 (N_12511,N_9233,N_10787);
and U12512 (N_12512,N_10285,N_11250);
or U12513 (N_12513,N_8990,N_7359);
and U12514 (N_12514,N_10210,N_9369);
nor U12515 (N_12515,N_7550,N_8542);
and U12516 (N_12516,N_10999,N_6456);
and U12517 (N_12517,N_7783,N_7350);
and U12518 (N_12518,N_6759,N_6069);
or U12519 (N_12519,N_7270,N_11681);
nand U12520 (N_12520,N_8533,N_9475);
nand U12521 (N_12521,N_6815,N_11180);
and U12522 (N_12522,N_7443,N_8484);
and U12523 (N_12523,N_8986,N_8347);
or U12524 (N_12524,N_10108,N_6687);
or U12525 (N_12525,N_7634,N_7061);
nand U12526 (N_12526,N_9389,N_8038);
xor U12527 (N_12527,N_10049,N_8998);
nand U12528 (N_12528,N_7907,N_10281);
nor U12529 (N_12529,N_8951,N_7723);
and U12530 (N_12530,N_11869,N_8229);
or U12531 (N_12531,N_8518,N_7453);
xnor U12532 (N_12532,N_11161,N_11677);
and U12533 (N_12533,N_8001,N_6544);
xor U12534 (N_12534,N_7135,N_11838);
nand U12535 (N_12535,N_6343,N_6973);
nor U12536 (N_12536,N_9052,N_7030);
and U12537 (N_12537,N_6172,N_10098);
xor U12538 (N_12538,N_7420,N_10647);
nand U12539 (N_12539,N_8753,N_11667);
nor U12540 (N_12540,N_11269,N_8611);
or U12541 (N_12541,N_11198,N_9986);
nand U12542 (N_12542,N_9357,N_8884);
nand U12543 (N_12543,N_11426,N_8408);
nor U12544 (N_12544,N_9633,N_8666);
and U12545 (N_12545,N_10019,N_9351);
and U12546 (N_12546,N_8173,N_6741);
nand U12547 (N_12547,N_11115,N_11646);
and U12548 (N_12548,N_7285,N_10137);
xor U12549 (N_12549,N_11435,N_7259);
xnor U12550 (N_12550,N_8897,N_8816);
or U12551 (N_12551,N_8682,N_10225);
and U12552 (N_12552,N_9920,N_11274);
nor U12553 (N_12553,N_6492,N_6659);
and U12554 (N_12554,N_9857,N_6041);
nor U12555 (N_12555,N_11509,N_8861);
nand U12556 (N_12556,N_7911,N_6897);
nand U12557 (N_12557,N_9009,N_9289);
nand U12558 (N_12558,N_7589,N_6004);
nor U12559 (N_12559,N_7103,N_9039);
nand U12560 (N_12560,N_6304,N_10416);
and U12561 (N_12561,N_9562,N_9258);
or U12562 (N_12562,N_7305,N_9610);
or U12563 (N_12563,N_7351,N_9564);
and U12564 (N_12564,N_10058,N_10780);
nand U12565 (N_12565,N_7587,N_10563);
nand U12566 (N_12566,N_6509,N_6190);
and U12567 (N_12567,N_6147,N_9203);
and U12568 (N_12568,N_11013,N_6802);
nand U12569 (N_12569,N_8006,N_10974);
nand U12570 (N_12570,N_9501,N_9479);
nand U12571 (N_12571,N_10632,N_6909);
nand U12572 (N_12572,N_6196,N_6814);
and U12573 (N_12573,N_10641,N_9546);
xor U12574 (N_12574,N_8193,N_7628);
or U12575 (N_12575,N_8534,N_7554);
or U12576 (N_12576,N_8906,N_8287);
or U12577 (N_12577,N_9126,N_6408);
or U12578 (N_12578,N_6891,N_10203);
nand U12579 (N_12579,N_6499,N_7987);
nor U12580 (N_12580,N_6947,N_10154);
nor U12581 (N_12581,N_6201,N_6079);
nor U12582 (N_12582,N_10185,N_11413);
or U12583 (N_12583,N_9143,N_9270);
or U12584 (N_12584,N_11688,N_11533);
nor U12585 (N_12585,N_9634,N_7962);
nor U12586 (N_12586,N_6122,N_10629);
or U12587 (N_12587,N_7694,N_8079);
xor U12588 (N_12588,N_6290,N_8192);
nand U12589 (N_12589,N_9911,N_6968);
or U12590 (N_12590,N_10738,N_7408);
and U12591 (N_12591,N_7665,N_7411);
nand U12592 (N_12592,N_9218,N_8202);
nor U12593 (N_12593,N_7772,N_10922);
and U12594 (N_12594,N_8854,N_10595);
nor U12595 (N_12595,N_11879,N_11999);
nor U12596 (N_12596,N_11592,N_9764);
and U12597 (N_12597,N_11129,N_8974);
nor U12598 (N_12598,N_9918,N_11246);
nand U12599 (N_12599,N_9741,N_6792);
and U12600 (N_12600,N_7743,N_7119);
or U12601 (N_12601,N_9673,N_8743);
or U12602 (N_12602,N_11747,N_8434);
nand U12603 (N_12603,N_10675,N_9840);
and U12604 (N_12604,N_7399,N_11265);
or U12605 (N_12605,N_7819,N_9833);
or U12606 (N_12606,N_6649,N_7927);
and U12607 (N_12607,N_6914,N_10390);
and U12608 (N_12608,N_7198,N_8152);
nand U12609 (N_12609,N_9141,N_6530);
nor U12610 (N_12610,N_7538,N_11858);
or U12611 (N_12611,N_10573,N_6831);
xor U12612 (N_12612,N_7661,N_8397);
nor U12613 (N_12613,N_8843,N_6048);
nor U12614 (N_12614,N_8418,N_9502);
xnor U12615 (N_12615,N_10088,N_8887);
nand U12616 (N_12616,N_9147,N_11812);
nor U12617 (N_12617,N_10788,N_7352);
or U12618 (N_12618,N_7284,N_6960);
nor U12619 (N_12619,N_8658,N_8875);
or U12620 (N_12620,N_6399,N_6182);
nand U12621 (N_12621,N_9667,N_8280);
or U12622 (N_12622,N_7288,N_6132);
nand U12623 (N_12623,N_8955,N_7062);
and U12624 (N_12624,N_6817,N_7234);
nand U12625 (N_12625,N_11339,N_10794);
nand U12626 (N_12626,N_8517,N_11380);
or U12627 (N_12627,N_9776,N_11575);
and U12628 (N_12628,N_11270,N_6683);
and U12629 (N_12629,N_11685,N_9701);
and U12630 (N_12630,N_8943,N_10451);
nand U12631 (N_12631,N_8027,N_9682);
xnor U12632 (N_12632,N_9923,N_8968);
and U12633 (N_12633,N_7695,N_11948);
or U12634 (N_12634,N_9063,N_10160);
or U12635 (N_12635,N_8809,N_11870);
nor U12636 (N_12636,N_7720,N_9537);
and U12637 (N_12637,N_9720,N_10032);
nand U12638 (N_12638,N_8148,N_6325);
and U12639 (N_12639,N_10178,N_11930);
or U12640 (N_12640,N_6750,N_6612);
nor U12641 (N_12641,N_10279,N_6293);
nor U12642 (N_12642,N_6992,N_7317);
nor U12643 (N_12643,N_6061,N_7323);
xor U12644 (N_12644,N_8462,N_11957);
nand U12645 (N_12645,N_7118,N_11412);
and U12646 (N_12646,N_8143,N_11106);
nor U12647 (N_12647,N_6780,N_7925);
nand U12648 (N_12648,N_10010,N_8092);
nand U12649 (N_12649,N_9419,N_11963);
and U12650 (N_12650,N_11101,N_10883);
nand U12651 (N_12651,N_9563,N_10356);
and U12652 (N_12652,N_11562,N_11229);
nor U12653 (N_12653,N_11798,N_6045);
nor U12654 (N_12654,N_8929,N_10393);
and U12655 (N_12655,N_9254,N_10056);
and U12656 (N_12656,N_11484,N_6794);
nand U12657 (N_12657,N_9922,N_6389);
nand U12658 (N_12658,N_9358,N_7597);
and U12659 (N_12659,N_10619,N_6117);
nand U12660 (N_12660,N_11219,N_6917);
and U12661 (N_12661,N_7222,N_11102);
or U12662 (N_12662,N_10606,N_7506);
nand U12663 (N_12663,N_11209,N_10583);
or U12664 (N_12664,N_8013,N_7354);
nor U12665 (N_12665,N_11557,N_10187);
and U12666 (N_12666,N_10289,N_11039);
or U12667 (N_12667,N_10259,N_9173);
nor U12668 (N_12668,N_8322,N_9196);
xnor U12669 (N_12669,N_11539,N_10635);
and U12670 (N_12670,N_10625,N_10742);
and U12671 (N_12671,N_8178,N_9995);
nor U12672 (N_12672,N_6056,N_6284);
and U12673 (N_12673,N_8926,N_6782);
and U12674 (N_12674,N_10985,N_7132);
nand U12675 (N_12675,N_10557,N_9271);
nand U12676 (N_12676,N_10459,N_6885);
or U12677 (N_12677,N_8914,N_6836);
and U12678 (N_12678,N_11607,N_10987);
nor U12679 (N_12679,N_6077,N_11856);
and U12680 (N_12680,N_6690,N_8474);
and U12681 (N_12681,N_6451,N_11872);
or U12682 (N_12682,N_7545,N_9902);
nor U12683 (N_12683,N_9286,N_9577);
xnor U12684 (N_12684,N_6787,N_8832);
nand U12685 (N_12685,N_10651,N_9456);
or U12686 (N_12686,N_6027,N_9997);
xnor U12687 (N_12687,N_6706,N_8098);
or U12688 (N_12688,N_8830,N_10732);
and U12689 (N_12689,N_6186,N_6887);
nor U12690 (N_12690,N_8721,N_6747);
nor U12691 (N_12691,N_8084,N_7633);
and U12692 (N_12692,N_11762,N_11097);
nor U12693 (N_12693,N_9835,N_8480);
nor U12694 (N_12694,N_10455,N_7499);
nor U12695 (N_12695,N_11944,N_7698);
nor U12696 (N_12696,N_8840,N_6713);
or U12697 (N_12697,N_10446,N_8476);
or U12698 (N_12698,N_7110,N_10030);
nor U12699 (N_12699,N_6138,N_8939);
nor U12700 (N_12700,N_8520,N_6545);
nor U12701 (N_12701,N_8818,N_11455);
and U12702 (N_12702,N_9558,N_6982);
nand U12703 (N_12703,N_6176,N_9156);
and U12704 (N_12704,N_9824,N_9444);
nand U12705 (N_12705,N_7446,N_9008);
and U12706 (N_12706,N_9101,N_8438);
and U12707 (N_12707,N_10692,N_7364);
xnor U12708 (N_12708,N_8947,N_7724);
nand U12709 (N_12709,N_8161,N_10378);
nand U12710 (N_12710,N_10420,N_7737);
or U12711 (N_12711,N_11043,N_8429);
nand U12712 (N_12712,N_10006,N_7165);
nor U12713 (N_12713,N_7024,N_6020);
nand U12714 (N_12714,N_11725,N_9157);
and U12715 (N_12715,N_7656,N_6967);
nor U12716 (N_12716,N_9404,N_6972);
and U12717 (N_12717,N_8216,N_8790);
and U12718 (N_12718,N_9306,N_9928);
and U12719 (N_12719,N_8775,N_7792);
and U12720 (N_12720,N_11177,N_9457);
and U12721 (N_12721,N_8738,N_6216);
xor U12722 (N_12722,N_10474,N_8779);
nor U12723 (N_12723,N_9299,N_9842);
nand U12724 (N_12724,N_11790,N_6590);
nor U12725 (N_12725,N_11849,N_11144);
nand U12726 (N_12726,N_10837,N_9730);
nand U12727 (N_12727,N_10447,N_9311);
nand U12728 (N_12728,N_6865,N_6989);
xnor U12729 (N_12729,N_11168,N_9596);
nor U12730 (N_12730,N_10572,N_10733);
nand U12731 (N_12731,N_6639,N_6898);
nand U12732 (N_12732,N_11974,N_6266);
and U12733 (N_12733,N_10942,N_10718);
and U12734 (N_12734,N_9729,N_10048);
nor U12735 (N_12735,N_7315,N_11573);
and U12736 (N_12736,N_11737,N_7872);
and U12737 (N_12737,N_11893,N_6936);
and U12738 (N_12738,N_10613,N_9791);
nand U12739 (N_12739,N_9699,N_6673);
or U12740 (N_12740,N_9592,N_6594);
nor U12741 (N_12741,N_10050,N_10574);
nand U12742 (N_12742,N_11769,N_6215);
nand U12743 (N_12743,N_10172,N_9523);
nand U12744 (N_12744,N_10750,N_10902);
nand U12745 (N_12745,N_10989,N_7719);
nand U12746 (N_12746,N_7613,N_7298);
nor U12747 (N_12747,N_8547,N_7038);
or U12748 (N_12748,N_6854,N_9308);
nand U12749 (N_12749,N_8081,N_9414);
and U12750 (N_12750,N_10403,N_11487);
nand U12751 (N_12751,N_11024,N_10041);
nand U12752 (N_12752,N_6870,N_9134);
or U12753 (N_12753,N_11800,N_6087);
or U12754 (N_12754,N_11716,N_6068);
or U12755 (N_12755,N_9927,N_9961);
nand U12756 (N_12756,N_11197,N_7754);
and U12757 (N_12757,N_8166,N_11558);
nor U12758 (N_12758,N_6028,N_8387);
or U12759 (N_12759,N_8573,N_9405);
or U12760 (N_12760,N_6217,N_11886);
nand U12761 (N_12761,N_11206,N_7001);
nand U12762 (N_12762,N_9746,N_6819);
nand U12763 (N_12763,N_6956,N_7381);
xnor U12764 (N_12764,N_6223,N_8576);
xor U12765 (N_12765,N_6235,N_10091);
nor U12766 (N_12766,N_9512,N_9550);
or U12767 (N_12767,N_9989,N_7837);
and U12768 (N_12768,N_8127,N_7167);
and U12769 (N_12769,N_11119,N_7191);
and U12770 (N_12770,N_7383,N_6066);
and U12771 (N_12771,N_8409,N_7232);
nor U12772 (N_12772,N_11428,N_10070);
or U12773 (N_12773,N_8739,N_6512);
xor U12774 (N_12774,N_8366,N_7919);
nor U12775 (N_12775,N_6929,N_7023);
nor U12776 (N_12776,N_8210,N_6576);
or U12777 (N_12777,N_9893,N_7852);
nand U12778 (N_12778,N_10964,N_6626);
and U12779 (N_12779,N_7032,N_8402);
and U12780 (N_12780,N_11625,N_11713);
xor U12781 (N_12781,N_6630,N_8423);
nor U12782 (N_12782,N_9455,N_7455);
nor U12783 (N_12783,N_6489,N_10047);
xor U12784 (N_12784,N_7530,N_9338);
and U12785 (N_12785,N_6534,N_9209);
nor U12786 (N_12786,N_11373,N_7500);
nand U12787 (N_12787,N_6084,N_11140);
nor U12788 (N_12788,N_10795,N_11698);
or U12789 (N_12789,N_6466,N_10413);
and U12790 (N_12790,N_6519,N_6123);
or U12791 (N_12791,N_10500,N_10973);
or U12792 (N_12792,N_9492,N_9885);
xnor U12793 (N_12793,N_6414,N_7782);
and U12794 (N_12794,N_8363,N_6783);
xor U12795 (N_12795,N_10959,N_8735);
nand U12796 (N_12796,N_6503,N_6012);
xnor U12797 (N_12797,N_11732,N_7790);
and U12798 (N_12798,N_7920,N_8617);
nor U12799 (N_12799,N_7966,N_8340);
xor U12800 (N_12800,N_7063,N_9439);
nand U12801 (N_12801,N_6473,N_7722);
or U12802 (N_12802,N_10827,N_8608);
nor U12803 (N_12803,N_8141,N_8487);
and U12804 (N_12804,N_6476,N_11916);
and U12805 (N_12805,N_9309,N_6333);
nor U12806 (N_12806,N_10819,N_10428);
and U12807 (N_12807,N_6495,N_7518);
or U12808 (N_12808,N_9751,N_8281);
or U12809 (N_12809,N_10754,N_9778);
nor U12810 (N_12810,N_7760,N_9725);
xor U12811 (N_12811,N_8898,N_10801);
xnor U12812 (N_12812,N_6303,N_11995);
nand U12813 (N_12813,N_7577,N_10046);
or U12814 (N_12814,N_8508,N_11645);
nor U12815 (N_12815,N_6674,N_7082);
or U12816 (N_12816,N_7214,N_6986);
and U12817 (N_12817,N_10398,N_7498);
nor U12818 (N_12818,N_7992,N_8562);
nor U12819 (N_12819,N_6677,N_7796);
nor U12820 (N_12820,N_11935,N_9689);
nand U12821 (N_12821,N_6160,N_11285);
xnor U12822 (N_12822,N_8522,N_11497);
and U12823 (N_12823,N_11580,N_11482);
nor U12824 (N_12824,N_8437,N_11215);
or U12825 (N_12825,N_9230,N_9717);
or U12826 (N_12826,N_6360,N_10482);
and U12827 (N_12827,N_9654,N_7000);
nor U12828 (N_12828,N_9436,N_8053);
or U12829 (N_12829,N_10602,N_7048);
nand U12830 (N_12830,N_10590,N_10610);
and U12831 (N_12831,N_6632,N_9011);
nand U12832 (N_12832,N_9914,N_11343);
or U12833 (N_12833,N_6166,N_11975);
nand U12834 (N_12834,N_7158,N_10507);
nor U12835 (N_12835,N_6021,N_11402);
nor U12836 (N_12836,N_7136,N_10270);
nor U12837 (N_12837,N_9611,N_10215);
and U12838 (N_12838,N_10992,N_7508);
or U12839 (N_12839,N_6010,N_8614);
nand U12840 (N_12840,N_11795,N_6808);
nand U12841 (N_12841,N_6723,N_11253);
nor U12842 (N_12842,N_9518,N_6671);
xor U12843 (N_12843,N_7956,N_9334);
nor U12844 (N_12844,N_8500,N_8036);
and U12845 (N_12845,N_11690,N_8186);
or U12846 (N_12846,N_7816,N_9094);
xnor U12847 (N_12847,N_11654,N_8447);
or U12848 (N_12848,N_10370,N_7598);
or U12849 (N_12849,N_7671,N_11033);
nor U12850 (N_12850,N_6827,N_8681);
nand U12851 (N_12851,N_6295,N_6421);
and U12852 (N_12852,N_10157,N_7994);
or U12853 (N_12853,N_10599,N_9984);
and U12854 (N_12854,N_11240,N_6165);
xor U12855 (N_12855,N_9360,N_11603);
nor U12856 (N_12856,N_7864,N_6988);
and U12857 (N_12857,N_8454,N_6664);
nand U12858 (N_12858,N_10663,N_11510);
nor U12859 (N_12859,N_10371,N_6696);
nand U12860 (N_12860,N_8112,N_11574);
or U12861 (N_12861,N_7854,N_11734);
nand U12862 (N_12862,N_11466,N_11203);
xnor U12863 (N_12863,N_6584,N_6959);
and U12864 (N_12864,N_8842,N_11514);
nor U12865 (N_12865,N_8282,N_10885);
nor U12866 (N_12866,N_7094,N_10330);
nand U12867 (N_12867,N_10524,N_10848);
and U12868 (N_12868,N_6005,N_8695);
nand U12869 (N_12869,N_11073,N_9205);
and U12870 (N_12870,N_9965,N_6994);
and U12871 (N_12871,N_11807,N_9621);
and U12872 (N_12872,N_9826,N_11759);
and U12873 (N_12873,N_10064,N_8050);
nand U12874 (N_12874,N_7895,N_10173);
nor U12875 (N_12875,N_11606,N_7325);
and U12876 (N_12876,N_8198,N_8800);
and U12877 (N_12877,N_10681,N_10679);
xor U12878 (N_12878,N_10843,N_9644);
and U12879 (N_12879,N_6761,N_11452);
nor U12880 (N_12880,N_7502,N_10124);
nand U12881 (N_12881,N_6541,N_6778);
and U12882 (N_12882,N_7988,N_7291);
xnor U12883 (N_12883,N_10799,N_11195);
or U12884 (N_12884,N_9330,N_9858);
nor U12885 (N_12885,N_9001,N_9079);
or U12886 (N_12886,N_9872,N_8766);
or U12887 (N_12887,N_6771,N_11045);
nand U12888 (N_12888,N_6855,N_6807);
and U12889 (N_12889,N_9830,N_7293);
nand U12890 (N_12890,N_10410,N_10680);
xor U12891 (N_12891,N_7731,N_6863);
and U12892 (N_12892,N_9762,N_8057);
and U12893 (N_12893,N_11612,N_11081);
xnor U12894 (N_12894,N_8925,N_9754);
nand U12895 (N_12895,N_7440,N_10953);
or U12896 (N_12896,N_6262,N_6680);
and U12897 (N_12897,N_11341,N_10062);
nor U12898 (N_12898,N_9212,N_9026);
nand U12899 (N_12899,N_9329,N_6383);
and U12900 (N_12900,N_8088,N_8285);
and U12901 (N_12901,N_10471,N_9005);
xnor U12902 (N_12902,N_11438,N_6434);
and U12903 (N_12903,N_9744,N_11874);
nand U12904 (N_12904,N_7757,N_10813);
xnor U12905 (N_12905,N_10156,N_7184);
nor U12906 (N_12906,N_11283,N_11154);
xnor U12907 (N_12907,N_11188,N_8217);
nand U12908 (N_12908,N_11941,N_9670);
nor U12909 (N_12909,N_10011,N_11403);
and U12910 (N_12910,N_11122,N_7557);
nor U12911 (N_12911,N_6225,N_9181);
xnor U12912 (N_12912,N_6700,N_8903);
and U12913 (N_12913,N_11408,N_7522);
nand U12914 (N_12914,N_10903,N_9547);
or U12915 (N_12915,N_11089,N_7811);
nand U12916 (N_12916,N_11094,N_8961);
or U12917 (N_12917,N_6208,N_8306);
or U12918 (N_12918,N_8822,N_7328);
and U12919 (N_12919,N_11696,N_7944);
or U12920 (N_12920,N_9950,N_8299);
xor U12921 (N_12921,N_6214,N_10054);
nand U12922 (N_12922,N_11214,N_11868);
and U12923 (N_12923,N_6715,N_8478);
or U12924 (N_12924,N_8415,N_10810);
nor U12925 (N_12925,N_8000,N_6553);
nor U12926 (N_12926,N_6091,N_6339);
xor U12927 (N_12927,N_11495,N_7679);
or U12928 (N_12928,N_11997,N_6405);
and U12929 (N_12929,N_6429,N_10192);
nor U12930 (N_12930,N_10730,N_9608);
nand U12931 (N_12931,N_10707,N_10016);
xor U12932 (N_12932,N_10762,N_6498);
nand U12933 (N_12933,N_11006,N_11938);
and U12934 (N_12934,N_7703,N_11925);
and U12935 (N_12935,N_6211,N_8833);
or U12936 (N_12936,N_10737,N_7595);
and U12937 (N_12937,N_7739,N_8651);
nand U12938 (N_12938,N_11421,N_11057);
nand U12939 (N_12939,N_8005,N_10634);
or U12940 (N_12940,N_8058,N_11221);
nand U12941 (N_12941,N_10009,N_8763);
and U12942 (N_12942,N_10864,N_11885);
xor U12943 (N_12943,N_9726,N_10856);
nor U12944 (N_12944,N_6744,N_9916);
and U12945 (N_12945,N_10201,N_10826);
or U12946 (N_12946,N_6454,N_7533);
and U12947 (N_12947,N_7166,N_6876);
xor U12948 (N_12948,N_10852,N_9867);
xnor U12949 (N_12949,N_8277,N_8233);
or U12950 (N_12950,N_7763,N_11110);
nand U12951 (N_12951,N_8902,N_6011);
or U12952 (N_12952,N_10516,N_8305);
or U12953 (N_12953,N_11184,N_7467);
and U12954 (N_12954,N_6017,N_6490);
nand U12955 (N_12955,N_7573,N_10089);
or U12956 (N_12956,N_6390,N_8941);
nand U12957 (N_12957,N_8713,N_6675);
or U12958 (N_12958,N_7311,N_8062);
xor U12959 (N_12959,N_9490,N_7789);
and U12960 (N_12960,N_9304,N_6111);
nor U12961 (N_12961,N_9114,N_9162);
nand U12962 (N_12962,N_8504,N_9463);
nand U12963 (N_12963,N_9151,N_7196);
or U12964 (N_12964,N_11722,N_9713);
nor U12965 (N_12965,N_8642,N_11475);
nor U12966 (N_12966,N_9481,N_10596);
or U12967 (N_12967,N_8502,N_10899);
and U12968 (N_12968,N_9480,N_7157);
nand U12969 (N_12969,N_9707,N_10441);
xnor U12970 (N_12970,N_8376,N_6105);
nor U12971 (N_12971,N_9756,N_7985);
or U12972 (N_12972,N_11278,N_6163);
xor U12973 (N_12973,N_8670,N_8132);
xnor U12974 (N_12974,N_11030,N_11405);
xor U12975 (N_12975,N_11676,N_9851);
or U12976 (N_12976,N_6526,N_6646);
nand U12977 (N_12977,N_11720,N_8785);
nor U12978 (N_12978,N_6620,N_11786);
or U12979 (N_12979,N_9793,N_7343);
and U12980 (N_12980,N_6841,N_11586);
nor U12981 (N_12981,N_6812,N_11331);
nand U12982 (N_12982,N_10509,N_7668);
or U12983 (N_12983,N_10350,N_6135);
nand U12984 (N_12984,N_11648,N_9967);
or U12985 (N_12985,N_8074,N_11841);
nor U12986 (N_12986,N_7774,N_7990);
nand U12987 (N_12987,N_11080,N_11037);
or U12988 (N_12988,N_9051,N_11016);
and U12989 (N_12989,N_6507,N_11333);
nand U12990 (N_12990,N_10752,N_6514);
nor U12991 (N_12991,N_9594,N_9942);
or U12992 (N_12992,N_9047,N_10689);
nor U12993 (N_12993,N_10174,N_7607);
or U12994 (N_12994,N_9524,N_7894);
or U12995 (N_12995,N_6275,N_10722);
nor U12996 (N_12996,N_8566,N_7833);
and U12997 (N_12997,N_9990,N_9049);
or U12998 (N_12998,N_9055,N_6342);
and U12999 (N_12999,N_8197,N_9880);
nand U13000 (N_13000,N_11325,N_6446);
and U13001 (N_13001,N_10097,N_7829);
xnor U13002 (N_13002,N_10419,N_7863);
nand U13003 (N_13003,N_8850,N_9265);
nand U13004 (N_13004,N_7257,N_10519);
nand U13005 (N_13005,N_9057,N_9844);
nand U13006 (N_13006,N_7637,N_7603);
xnor U13007 (N_13007,N_11182,N_11551);
nand U13008 (N_13008,N_10564,N_10208);
nand U13009 (N_13009,N_9345,N_11289);
nor U13010 (N_13010,N_9579,N_8718);
nand U13011 (N_13011,N_6562,N_11643);
or U13012 (N_13012,N_11068,N_10086);
and U13013 (N_13013,N_9777,N_9605);
xnor U13014 (N_13014,N_9232,N_10829);
nand U13015 (N_13015,N_10063,N_7152);
nor U13016 (N_13016,N_8054,N_6222);
nor U13017 (N_13017,N_8946,N_11067);
nor U13018 (N_13018,N_8964,N_8020);
or U13019 (N_13019,N_8170,N_10529);
nand U13020 (N_13020,N_8758,N_10473);
xnor U13021 (N_13021,N_7896,N_10200);
and U13022 (N_13022,N_8856,N_6305);
nor U13023 (N_13023,N_8045,N_11390);
xor U13024 (N_13024,N_8182,N_9897);
and U13025 (N_13025,N_7248,N_9498);
and U13026 (N_13026,N_11058,N_9343);
nor U13027 (N_13027,N_9281,N_10318);
nor U13028 (N_13028,N_11877,N_9898);
nand U13029 (N_13029,N_8007,N_6799);
or U13030 (N_13030,N_9819,N_6950);
or U13031 (N_13031,N_7457,N_11212);
or U13032 (N_13032,N_7385,N_8443);
and U13033 (N_13033,N_10303,N_8310);
or U13034 (N_13034,N_9424,N_9705);
nor U13035 (N_13035,N_8552,N_7003);
and U13036 (N_13036,N_6431,N_9421);
nor U13037 (N_13037,N_8927,N_7830);
xor U13038 (N_13038,N_8252,N_10153);
nor U13039 (N_13039,N_7501,N_6652);
or U13040 (N_13040,N_7470,N_8526);
and U13041 (N_13041,N_8855,N_9874);
nand U13042 (N_13042,N_7664,N_8432);
or U13043 (N_13043,N_10533,N_7097);
and U13044 (N_13044,N_9120,N_6263);
nor U13045 (N_13045,N_9845,N_6720);
xor U13046 (N_13046,N_7631,N_6663);
and U13047 (N_13047,N_6574,N_11808);
or U13048 (N_13048,N_9906,N_6478);
nor U13049 (N_13049,N_9346,N_9585);
nor U13050 (N_13050,N_11719,N_8046);
or U13051 (N_13051,N_8742,N_6738);
nand U13052 (N_13052,N_9519,N_7145);
nor U13053 (N_13053,N_8630,N_10131);
xor U13054 (N_13054,N_10949,N_7855);
nand U13055 (N_13055,N_10404,N_11525);
or U13056 (N_13056,N_11430,N_11652);
nor U13057 (N_13057,N_10923,N_8507);
and U13058 (N_13058,N_7025,N_11702);
or U13059 (N_13059,N_10914,N_9383);
nor U13060 (N_13060,N_9970,N_9124);
or U13061 (N_13061,N_10081,N_11303);
and U13062 (N_13062,N_6337,N_9469);
and U13063 (N_13063,N_11745,N_11546);
and U13064 (N_13064,N_9179,N_11427);
or U13065 (N_13065,N_8761,N_8228);
or U13066 (N_13066,N_10716,N_11158);
nand U13067 (N_13067,N_8121,N_11824);
and U13068 (N_13068,N_9569,N_7116);
nor U13069 (N_13069,N_9917,N_10746);
or U13070 (N_13070,N_10701,N_7594);
nand U13071 (N_13071,N_6963,N_6583);
xnor U13072 (N_13072,N_10453,N_8172);
and U13073 (N_13073,N_11597,N_6309);
nand U13074 (N_13074,N_6872,N_11775);
nor U13075 (N_13075,N_11318,N_7012);
or U13076 (N_13076,N_7199,N_6392);
and U13077 (N_13077,N_11894,N_9013);
nor U13078 (N_13078,N_8494,N_7609);
nor U13079 (N_13079,N_10665,N_9302);
nor U13080 (N_13080,N_8385,N_11327);
nor U13081 (N_13081,N_10638,N_7618);
nor U13082 (N_13082,N_7208,N_8026);
and U13083 (N_13083,N_10823,N_7952);
nor U13084 (N_13084,N_7749,N_8694);
nor U13085 (N_13085,N_8558,N_6939);
xnor U13086 (N_13086,N_11348,N_8190);
xnor U13087 (N_13087,N_11384,N_6419);
or U13088 (N_13088,N_10368,N_9387);
xnor U13089 (N_13089,N_7541,N_6650);
nor U13090 (N_13090,N_11955,N_10120);
nor U13091 (N_13091,N_6734,N_10000);
or U13092 (N_13092,N_11750,N_9122);
or U13093 (N_13093,N_6032,N_7689);
and U13094 (N_13094,N_6088,N_9443);
nor U13095 (N_13095,N_7374,N_8424);
nor U13096 (N_13096,N_9262,N_6977);
and U13097 (N_13097,N_11252,N_6560);
or U13098 (N_13098,N_10274,N_9242);
or U13099 (N_13099,N_7642,N_6832);
nor U13100 (N_13100,N_10053,N_11620);
or U13101 (N_13101,N_8770,N_6238);
and U13102 (N_13102,N_10822,N_9442);
nand U13103 (N_13103,N_11287,N_10257);
or U13104 (N_13104,N_11660,N_8960);
nor U13105 (N_13105,N_9759,N_10682);
nor U13106 (N_13106,N_6167,N_7361);
and U13107 (N_13107,N_7339,N_9253);
or U13108 (N_13108,N_7672,N_9066);
nand U13109 (N_13109,N_6520,N_8936);
nor U13110 (N_13110,N_9133,N_10538);
nand U13111 (N_13111,N_10927,N_7449);
and U13112 (N_13112,N_11236,N_8649);
nor U13113 (N_13113,N_10804,N_8653);
or U13114 (N_13114,N_8803,N_9601);
nand U13115 (N_13115,N_11244,N_11116);
nand U13116 (N_13116,N_6298,N_6641);
nor U13117 (N_13117,N_8195,N_7108);
nor U13118 (N_13118,N_8196,N_11268);
or U13119 (N_13119,N_7036,N_6326);
or U13120 (N_13120,N_9295,N_11436);
nand U13121 (N_13121,N_9964,N_7391);
or U13122 (N_13122,N_9941,N_7282);
and U13123 (N_13123,N_10890,N_11383);
nand U13124 (N_13124,N_11241,N_10512);
or U13125 (N_13125,N_11920,N_6459);
and U13126 (N_13126,N_8699,N_6847);
and U13127 (N_13127,N_6816,N_7133);
or U13128 (N_13128,N_11568,N_7102);
nand U13129 (N_13129,N_7892,N_7401);
nand U13130 (N_13130,N_10146,N_7014);
nand U13131 (N_13131,N_8011,N_11793);
or U13132 (N_13132,N_8245,N_7572);
nand U13133 (N_13133,N_11731,N_10305);
nand U13134 (N_13134,N_9588,N_6387);
xor U13135 (N_13135,N_7130,N_6767);
and U13136 (N_13136,N_11072,N_10007);
nand U13137 (N_13137,N_8175,N_9237);
or U13138 (N_13138,N_7857,N_10026);
or U13139 (N_13139,N_9332,N_8019);
or U13140 (N_13140,N_11796,N_9398);
xnor U13141 (N_13141,N_6086,N_11946);
xnor U13142 (N_13142,N_7219,N_9300);
and U13143 (N_13143,N_11317,N_7580);
nor U13144 (N_13144,N_7341,N_6647);
xnor U13145 (N_13145,N_7848,N_8338);
and U13146 (N_13146,N_6935,N_8706);
and U13147 (N_13147,N_8238,N_6025);
and U13148 (N_13148,N_11985,N_6109);
nor U13149 (N_13149,N_10639,N_7755);
or U13150 (N_13150,N_9255,N_9510);
or U13151 (N_13151,N_7916,N_7709);
and U13152 (N_13152,N_6113,N_10697);
xnor U13153 (N_13153,N_11335,N_7154);
and U13154 (N_13154,N_11323,N_8293);
or U13155 (N_13155,N_10690,N_8802);
nand U13156 (N_13156,N_8748,N_10631);
and U13157 (N_13157,N_11489,N_10720);
nand U13158 (N_13158,N_9656,N_9722);
or U13159 (N_13159,N_11272,N_8381);
xnor U13160 (N_13160,N_6388,N_10317);
nor U13161 (N_13161,N_8792,N_11519);
nand U13162 (N_13162,N_9468,N_8538);
or U13163 (N_13163,N_9149,N_7667);
or U13164 (N_13164,N_7465,N_9372);
or U13165 (N_13165,N_7179,N_10603);
nor U13166 (N_13166,N_9721,N_7186);
nand U13167 (N_13167,N_11797,N_6140);
or U13168 (N_13168,N_7240,N_7326);
or U13169 (N_13169,N_8393,N_8725);
and U13170 (N_13170,N_10576,N_8032);
or U13171 (N_13171,N_9277,N_9349);
nor U13172 (N_13172,N_7778,N_9174);
or U13173 (N_13173,N_11637,N_11733);
nor U13174 (N_13174,N_8360,N_7027);
and U13175 (N_13175,N_8657,N_10597);
nand U13176 (N_13176,N_6323,N_11973);
xor U13177 (N_13177,N_7101,N_8623);
and U13178 (N_13178,N_9031,N_9553);
xnor U13179 (N_13179,N_6875,N_8339);
nand U13180 (N_13180,N_6152,N_6153);
nor U13181 (N_13181,N_9877,N_9727);
nand U13182 (N_13182,N_10109,N_6881);
or U13183 (N_13183,N_10379,N_8262);
xor U13184 (N_13184,N_10405,N_10374);
or U13185 (N_13185,N_7773,N_8628);
nor U13186 (N_13186,N_6941,N_7534);
or U13187 (N_13187,N_9117,N_7914);
nor U13188 (N_13188,N_9708,N_11754);
nand U13189 (N_13189,N_7226,N_11961);
nand U13190 (N_13190,N_8448,N_10025);
xor U13191 (N_13191,N_11128,N_10217);
nand U13192 (N_13192,N_10909,N_11494);
nand U13193 (N_13193,N_6824,N_8530);
nand U13194 (N_13194,N_7590,N_11151);
or U13195 (N_13195,N_6569,N_7161);
nand U13196 (N_13196,N_11830,N_8466);
nor U13197 (N_13197,N_10346,N_9747);
and U13198 (N_13198,N_8100,N_9127);
and U13199 (N_13199,N_11194,N_11829);
or U13200 (N_13200,N_8768,N_9869);
nand U13201 (N_13201,N_7918,N_7043);
nor U13202 (N_13202,N_9775,N_9247);
or U13203 (N_13203,N_9570,N_11422);
or U13204 (N_13204,N_9538,N_8568);
or U13205 (N_13205,N_11954,N_9211);
and U13206 (N_13206,N_8270,N_8283);
or U13207 (N_13207,N_7009,N_6202);
xor U13208 (N_13208,N_10467,N_11032);
or U13209 (N_13209,N_11216,N_7681);
or U13210 (N_13210,N_10227,N_6366);
nor U13211 (N_13211,N_8486,N_7933);
nand U13212 (N_13212,N_10412,N_6518);
nor U13213 (N_13213,N_11810,N_8625);
nand U13214 (N_13214,N_10844,N_9805);
and U13215 (N_13215,N_11774,N_6999);
nand U13216 (N_13216,N_10143,N_6396);
or U13217 (N_13217,N_10079,N_6588);
and U13218 (N_13218,N_11537,N_7400);
nand U13219 (N_13219,N_6175,N_6155);
nor U13220 (N_13220,N_9111,N_9037);
or U13221 (N_13221,N_9600,N_7393);
or U13222 (N_13222,N_10463,N_7382);
and U13223 (N_13223,N_7986,N_8420);
or U13224 (N_13224,N_11353,N_7878);
and U13225 (N_13225,N_10060,N_10628);
or U13226 (N_13226,N_6270,N_11748);
nand U13227 (N_13227,N_8377,N_7010);
or U13228 (N_13228,N_9425,N_7752);
or U13229 (N_13229,N_7929,N_11582);
nor U13230 (N_13230,N_10534,N_8988);
nand U13231 (N_13231,N_10617,N_9591);
nor U13232 (N_13232,N_6099,N_11861);
or U13233 (N_13233,N_7329,N_7960);
xor U13234 (N_13234,N_9159,N_9142);
and U13235 (N_13235,N_6395,N_11712);
nand U13236 (N_13236,N_10038,N_7375);
nand U13237 (N_13237,N_8218,N_10117);
nand U13238 (N_13238,N_7592,N_10814);
nand U13239 (N_13239,N_9796,N_11742);
nor U13240 (N_13240,N_9719,N_7369);
or U13241 (N_13241,N_9781,N_11069);
nand U13242 (N_13242,N_6703,N_10189);
nand U13243 (N_13243,N_6474,N_9059);
and U13244 (N_13244,N_8827,N_10193);
or U13245 (N_13245,N_6363,N_7194);
nand U13246 (N_13246,N_8123,N_11943);
or U13247 (N_13247,N_6923,N_9244);
nor U13248 (N_13248,N_11862,N_6050);
and U13249 (N_13249,N_10221,N_8068);
or U13250 (N_13250,N_9339,N_8326);
or U13251 (N_13251,N_8213,N_8917);
nor U13252 (N_13252,N_6546,N_11141);
nand U13253 (N_13253,N_8839,N_9381);
and U13254 (N_13254,N_7771,N_8286);
or U13255 (N_13255,N_11313,N_10448);
nor U13256 (N_13256,N_9178,N_9541);
or U13257 (N_13257,N_8335,N_11309);
nor U13258 (N_13258,N_8370,N_8386);
xnor U13259 (N_13259,N_7899,N_9229);
xnor U13260 (N_13260,N_9949,N_8321);
or U13261 (N_13261,N_7690,N_7775);
or U13262 (N_13262,N_10440,N_11307);
nor U13263 (N_13263,N_9925,N_6725);
or U13264 (N_13264,N_10386,N_7390);
nand U13265 (N_13265,N_9084,N_6022);
xor U13266 (N_13266,N_8811,N_10935);
nor U13267 (N_13267,N_6299,N_6469);
or U13268 (N_13268,N_6145,N_6335);
nor U13269 (N_13269,N_10677,N_8679);
nor U13270 (N_13270,N_6361,N_11564);
nor U13271 (N_13271,N_7844,N_11664);
or U13272 (N_13272,N_9336,N_9718);
nor U13273 (N_13273,N_7704,N_9640);
nand U13274 (N_13274,N_9102,N_9454);
or U13275 (N_13275,N_7098,N_8288);
nand U13276 (N_13276,N_7124,N_10743);
nand U13277 (N_13277,N_7302,N_8771);
nor U13278 (N_13278,N_9678,N_7733);
nor U13279 (N_13279,N_11299,N_7057);
and U13280 (N_13280,N_7313,N_7822);
and U13281 (N_13281,N_10005,N_10968);
and U13282 (N_13282,N_11541,N_7867);
nor U13283 (N_13283,N_11121,N_6910);
and U13284 (N_13284,N_10857,N_6024);
nor U13285 (N_13285,N_9929,N_6292);
nor U13286 (N_13286,N_6697,N_7378);
and U13287 (N_13287,N_8700,N_11009);
nor U13288 (N_13288,N_10162,N_9852);
nand U13289 (N_13289,N_11387,N_11689);
and U13290 (N_13290,N_8064,N_6940);
xnor U13291 (N_13291,N_6995,N_10366);
xnor U13292 (N_13292,N_8080,N_8523);
and U13293 (N_13293,N_7225,N_6364);
nand U13294 (N_13294,N_8512,N_8982);
nor U13295 (N_13295,N_7273,N_10611);
or U13296 (N_13296,N_6296,N_8578);
nand U13297 (N_13297,N_11905,N_6843);
nor U13298 (N_13298,N_7496,N_9215);
or U13299 (N_13299,N_7487,N_6869);
or U13300 (N_13300,N_7645,N_8345);
nand U13301 (N_13301,N_11155,N_6668);
nand U13302 (N_13302,N_7490,N_10678);
and U13303 (N_13303,N_8563,N_7627);
xor U13304 (N_13304,N_6279,N_11926);
and U13305 (N_13305,N_11358,N_11357);
and U13306 (N_13306,N_9938,N_10938);
or U13307 (N_13307,N_10186,N_7578);
or U13308 (N_13308,N_9417,N_6884);
nand U13309 (N_13309,N_8253,N_10868);
xor U13310 (N_13310,N_11019,N_8535);
and U13311 (N_13311,N_6159,N_11276);
and U13312 (N_13312,N_11008,N_8620);
and U13313 (N_13313,N_7294,N_10195);
or U13314 (N_13314,N_6351,N_10779);
nand U13315 (N_13315,N_7466,N_11003);
nand U13316 (N_13316,N_6136,N_8495);
and U13317 (N_13317,N_11321,N_7639);
nand U13318 (N_13318,N_8863,N_6874);
and U13319 (N_13319,N_9297,N_9477);
nand U13320 (N_13320,N_8259,N_10114);
nor U13321 (N_13321,N_8696,N_7392);
or U13322 (N_13322,N_11389,N_6848);
nor U13323 (N_13323,N_10981,N_10501);
xor U13324 (N_13324,N_9113,N_6608);
and U13325 (N_13325,N_9248,N_11695);
and U13326 (N_13326,N_9736,N_7520);
nor U13327 (N_13327,N_11978,N_10372);
and U13328 (N_13328,N_10342,N_8741);
or U13329 (N_13329,N_10816,N_8870);
nor U13330 (N_13330,N_10391,N_7151);
nand U13331 (N_13331,N_7687,N_10082);
nand U13332 (N_13332,N_8373,N_7223);
and U13333 (N_13333,N_8587,N_11044);
and U13334 (N_13334,N_7011,N_8652);
or U13335 (N_13335,N_11576,N_8412);
and U13336 (N_13336,N_9060,N_8155);
nand U13337 (N_13337,N_6864,N_6927);
xor U13338 (N_13338,N_7266,N_9566);
nor U13339 (N_13339,N_7202,N_6691);
nor U13340 (N_13340,N_11351,N_8120);
or U13341 (N_13341,N_7527,N_11306);
and U13342 (N_13342,N_9690,N_7360);
or U13343 (N_13343,N_10957,N_6593);
xnor U13344 (N_13344,N_11996,N_9680);
nor U13345 (N_13345,N_6327,N_7460);
and U13346 (N_13346,N_11228,N_6300);
and U13347 (N_13347,N_6161,N_6063);
xor U13348 (N_13348,N_11170,N_9834);
and U13349 (N_13349,N_6665,N_11230);
and U13350 (N_13350,N_9347,N_8675);
xnor U13351 (N_13351,N_8554,N_11298);
and U13352 (N_13352,N_6592,N_11528);
nor U13353 (N_13353,N_7246,N_9543);
or U13354 (N_13354,N_6991,N_7958);
xnor U13355 (N_13355,N_6007,N_6622);
or U13356 (N_13356,N_10768,N_6768);
xor U13357 (N_13357,N_11919,N_9320);
nor U13358 (N_13358,N_6370,N_8812);
nor U13359 (N_13359,N_11457,N_11979);
nor U13360 (N_13360,N_7068,N_11934);
nand U13361 (N_13361,N_10988,N_9187);
and U13362 (N_13362,N_7623,N_6484);
nor U13363 (N_13363,N_9935,N_8844);
nand U13364 (N_13364,N_11330,N_9048);
and U13365 (N_13365,N_6524,N_11811);
nand U13366 (N_13366,N_11486,N_9953);
or U13367 (N_13367,N_9940,N_9314);
nor U13368 (N_13368,N_6149,N_6523);
xor U13369 (N_13369,N_8461,N_8874);
xnor U13370 (N_13370,N_6857,N_11227);
nand U13371 (N_13371,N_9257,N_9973);
xnor U13372 (N_13372,N_6203,N_9100);
or U13373 (N_13373,N_8866,N_11258);
and U13374 (N_13374,N_8767,N_8047);
nand U13375 (N_13375,N_9839,N_11461);
and U13376 (N_13376,N_9493,N_6877);
nor U13377 (N_13377,N_9868,N_11018);
nand U13378 (N_13378,N_6212,N_10726);
nor U13379 (N_13379,N_7591,N_6347);
nor U13380 (N_13380,N_8010,N_6234);
or U13381 (N_13381,N_7342,N_7659);
nand U13382 (N_13382,N_9535,N_8967);
and U13383 (N_13383,N_9963,N_10326);
nor U13384 (N_13384,N_6393,N_10406);
or U13385 (N_13385,N_6078,N_11082);
and U13386 (N_13386,N_9098,N_8845);
nand U13387 (N_13387,N_9497,N_9710);
or U13388 (N_13388,N_10457,N_7791);
xor U13389 (N_13389,N_11534,N_6770);
xor U13390 (N_13390,N_6638,N_9688);
or U13391 (N_13391,N_8901,N_10969);
nor U13392 (N_13392,N_11031,N_10783);
and U13393 (N_13393,N_7072,N_7797);
nor U13394 (N_13394,N_6619,N_10704);
or U13395 (N_13395,N_8208,N_8515);
nand U13396 (N_13396,N_10702,N_8669);
nor U13397 (N_13397,N_7824,N_7770);
nor U13398 (N_13398,N_7053,N_8239);
or U13399 (N_13399,N_10424,N_8860);
nor U13400 (N_13400,N_6618,N_7081);
nor U13401 (N_13401,N_10669,N_10384);
nand U13402 (N_13402,N_8516,N_10921);
xor U13403 (N_13403,N_9639,N_11201);
and U13404 (N_13404,N_11569,N_7491);
nand U13405 (N_13405,N_7941,N_10917);
xor U13406 (N_13406,N_11315,N_6127);
and U13407 (N_13407,N_6948,N_9128);
or U13408 (N_13408,N_7193,N_10490);
nor U13409 (N_13409,N_11832,N_9797);
nor U13410 (N_13410,N_7488,N_11880);
nor U13411 (N_13411,N_11970,N_8944);
nand U13412 (N_13412,N_8728,N_9628);
and U13413 (N_13413,N_9034,N_10415);
and U13414 (N_13414,N_8956,N_8422);
and U13415 (N_13415,N_9112,N_7414);
and U13416 (N_13416,N_6660,N_7271);
nand U13417 (N_13417,N_8249,N_10551);
and U13418 (N_13418,N_11029,N_6312);
nor U13419 (N_13419,N_8791,N_11364);
or U13420 (N_13420,N_9448,N_7251);
nand U13421 (N_13421,N_9291,N_7891);
and U13422 (N_13422,N_10970,N_6245);
or U13423 (N_13423,N_7109,N_10434);
nand U13424 (N_13424,N_7345,N_10083);
or U13425 (N_13425,N_11609,N_6246);
xnor U13426 (N_13426,N_7486,N_10345);
nor U13427 (N_13427,N_11633,N_6437);
nor U13428 (N_13428,N_10930,N_11839);
nor U13429 (N_13429,N_7982,N_6426);
and U13430 (N_13430,N_8154,N_9450);
nor U13431 (N_13431,N_11023,N_10727);
and U13432 (N_13432,N_9954,N_9811);
nand U13433 (N_13433,N_7310,N_10614);
and U13434 (N_13434,N_10401,N_11511);
or U13435 (N_13435,N_6539,N_10841);
or U13436 (N_13436,N_9197,N_10247);
xnor U13437 (N_13437,N_11450,N_6784);
or U13438 (N_13438,N_10481,N_8886);
and U13439 (N_13439,N_9733,N_11991);
nand U13440 (N_13440,N_6435,N_11202);
nor U13441 (N_13441,N_8730,N_7087);
xnor U13442 (N_13442,N_10113,N_6355);
and U13443 (N_13443,N_7450,N_9681);
xnor U13444 (N_13444,N_7647,N_7377);
or U13445 (N_13445,N_11336,N_9522);
or U13446 (N_13446,N_7441,N_11505);
and U13447 (N_13447,N_7015,N_11231);
or U13448 (N_13448,N_8570,N_9161);
nand U13449 (N_13449,N_9279,N_6942);
nor U13450 (N_13450,N_8660,N_11578);
nor U13451 (N_13451,N_6549,N_8250);
nand U13452 (N_13452,N_7509,N_10202);
nand U13453 (N_13453,N_6642,N_8680);
nand U13454 (N_13454,N_7524,N_8346);
nor U13455 (N_13455,N_7373,N_6095);
and U13456 (N_13456,N_6124,N_10161);
nor U13457 (N_13457,N_8457,N_11233);
xnor U13458 (N_13458,N_10846,N_7803);
or U13459 (N_13459,N_10299,N_6883);
xor U13460 (N_13460,N_8702,N_6047);
and U13461 (N_13461,N_6890,N_7606);
xnor U13462 (N_13462,N_11238,N_6198);
or U13463 (N_13463,N_10948,N_11964);
and U13464 (N_13464,N_10712,N_10667);
xnor U13465 (N_13465,N_9303,N_9728);
or U13466 (N_13466,N_6142,N_11697);
nand U13467 (N_13467,N_10307,N_9571);
nand U13468 (N_13468,N_8189,N_10184);
or U13469 (N_13469,N_8672,N_8727);
or U13470 (N_13470,N_10438,N_9958);
xnor U13471 (N_13471,N_9411,N_11765);
and U13472 (N_13472,N_10905,N_9067);
and U13473 (N_13473,N_6043,N_9883);
or U13474 (N_13474,N_9294,N_8243);
or U13475 (N_13475,N_10331,N_10587);
nand U13476 (N_13476,N_6195,N_10966);
and U13477 (N_13477,N_8479,N_6141);
and U13478 (N_13478,N_11764,N_11936);
and U13479 (N_13479,N_6494,N_9549);
and U13480 (N_13480,N_6398,N_6316);
and U13481 (N_13481,N_10555,N_9000);
nand U13482 (N_13482,N_8814,N_9198);
and U13483 (N_13483,N_8468,N_9103);
or U13484 (N_13484,N_6980,N_10068);
nor U13485 (N_13485,N_9919,N_11123);
nor U13486 (N_13486,N_9952,N_8160);
nor U13487 (N_13487,N_6191,N_10396);
nor U13488 (N_13488,N_7946,N_7178);
xnor U13489 (N_13489,N_7700,N_8102);
or U13490 (N_13490,N_6144,N_11692);
and U13491 (N_13491,N_9947,N_8521);
or U13492 (N_13492,N_7515,N_7424);
and U13493 (N_13493,N_11666,N_8754);
and U13494 (N_13494,N_10655,N_7614);
nand U13495 (N_13495,N_10488,N_6460);
or U13496 (N_13496,N_8091,N_9014);
or U13497 (N_13497,N_11931,N_7923);
or U13498 (N_13498,N_10882,N_10094);
nor U13499 (N_13499,N_6769,N_7997);
nor U13500 (N_13500,N_8404,N_9661);
and U13501 (N_13501,N_8783,N_10525);
or U13502 (N_13502,N_7442,N_10290);
or U13503 (N_13503,N_8575,N_8724);
nor U13504 (N_13504,N_7540,N_7558);
nor U13505 (N_13505,N_10498,N_9384);
nor U13506 (N_13506,N_8545,N_10792);
nor U13507 (N_13507,N_7963,N_9460);
nand U13508 (N_13508,N_7741,N_10879);
nand U13509 (N_13509,N_9813,N_10874);
and U13510 (N_13510,N_6422,N_9578);
or U13511 (N_13511,N_7970,N_8030);
and U13512 (N_13512,N_10335,N_9887);
nand U13513 (N_13513,N_7563,N_7742);
and U13514 (N_13514,N_11382,N_9222);
and U13515 (N_13515,N_8569,N_9798);
and U13516 (N_13516,N_6332,N_7040);
nand U13517 (N_13517,N_6900,N_10170);
nor U13518 (N_13518,N_7612,N_10104);
or U13519 (N_13519,N_7576,N_10658);
and U13520 (N_13520,N_9556,N_11785);
and U13521 (N_13521,N_6984,N_7033);
or U13522 (N_13522,N_8206,N_7870);
nand U13523 (N_13523,N_11017,N_7295);
or U13524 (N_13524,N_7922,N_10674);
nand U13525 (N_13525,N_7213,N_9962);
xor U13526 (N_13526,N_11104,N_8413);
and U13527 (N_13527,N_6252,N_8073);
xnor U13528 (N_13528,N_7890,N_11324);
and U13529 (N_13529,N_10808,N_7394);
and U13530 (N_13530,N_7217,N_9135);
nand U13531 (N_13531,N_9937,N_10971);
nand U13532 (N_13532,N_11545,N_10321);
nor U13533 (N_13533,N_11501,N_9180);
or U13534 (N_13534,N_6352,N_7079);
or U13535 (N_13535,N_6606,N_10650);
nand U13536 (N_13536,N_8003,N_7045);
or U13537 (N_13537,N_8641,N_9183);
nor U13538 (N_13538,N_6051,N_6427);
nand U13539 (N_13539,N_8406,N_7939);
xnor U13540 (N_13540,N_9993,N_8881);
nor U13541 (N_13541,N_7847,N_11515);
nor U13542 (N_13542,N_10560,N_8150);
or U13543 (N_13543,N_9900,N_9422);
nor U13544 (N_13544,N_10751,N_7138);
and U13545 (N_13545,N_10872,N_9760);
nand U13546 (N_13546,N_6705,N_6485);
nand U13547 (N_13547,N_10417,N_11217);
nand U13548 (N_13548,N_8972,N_11011);
or U13549 (N_13549,N_8571,N_9154);
nand U13550 (N_13550,N_10188,N_7875);
nand U13551 (N_13551,N_8503,N_9629);
nor U13552 (N_13552,N_9459,N_6281);
and U13553 (N_13553,N_7556,N_11555);
or U13554 (N_13554,N_8157,N_6901);
nor U13555 (N_13555,N_10012,N_8796);
and U13556 (N_13556,N_7092,N_11366);
nand U13557 (N_13557,N_11873,N_9107);
and U13558 (N_13558,N_9624,N_7984);
and U13559 (N_13559,N_9471,N_11038);
nor U13560 (N_13560,N_7143,N_6458);
or U13561 (N_13561,N_10309,N_6774);
or U13562 (N_13562,N_8701,N_7568);
and U13563 (N_13563,N_9322,N_11983);
and U13564 (N_13564,N_6550,N_7160);
nand U13565 (N_13565,N_7233,N_9821);
nand U13566 (N_13566,N_10668,N_10520);
and U13567 (N_13567,N_7995,N_8388);
or U13568 (N_13568,N_11297,N_8931);
xnor U13569 (N_13569,N_8528,N_11614);
nor U13570 (N_13570,N_10604,N_9412);
nand U13571 (N_13571,N_9335,N_7077);
and U13572 (N_13572,N_8824,N_9366);
nand U13573 (N_13573,N_7583,N_11470);
and U13574 (N_13574,N_7562,N_10375);
nor U13575 (N_13575,N_10556,N_10492);
or U13576 (N_13576,N_6743,N_10418);
and U13577 (N_13577,N_11145,N_9267);
nand U13578 (N_13578,N_7447,N_9352);
nor U13579 (N_13579,N_8034,N_11007);
nand U13580 (N_13580,N_8780,N_7163);
or U13581 (N_13581,N_7428,N_6852);
or U13582 (N_13582,N_7676,N_7134);
nor U13583 (N_13583,N_8473,N_8527);
xnor U13584 (N_13584,N_8807,N_6688);
and U13585 (N_13585,N_9669,N_11524);
and U13586 (N_13586,N_6558,N_10462);
nand U13587 (N_13587,N_9886,N_8453);
nor U13588 (N_13588,N_11251,N_6313);
and U13589 (N_13589,N_9703,N_7439);
nor U13590 (N_13590,N_7055,N_10508);
or U13591 (N_13591,N_10472,N_11047);
and U13592 (N_13592,N_8938,N_11149);
xnor U13593 (N_13593,N_8597,N_11267);
nor U13594 (N_13594,N_9494,N_9371);
nor U13595 (N_13595,N_8664,N_6772);
xnor U13596 (N_13596,N_9184,N_7821);
nor U13597 (N_13597,N_8215,N_11682);
nor U13598 (N_13598,N_6423,N_10945);
or U13599 (N_13599,N_8557,N_9256);
nor U13600 (N_13600,N_10140,N_11772);
or U13601 (N_13601,N_6943,N_8240);
nor U13602 (N_13602,N_11917,N_9118);
and U13603 (N_13603,N_6682,N_9948);
and U13604 (N_13604,N_10980,N_7525);
nand U13605 (N_13605,N_9836,N_8221);
or U13606 (N_13606,N_11529,N_11895);
nand U13607 (N_13607,N_8979,N_7693);
nand U13608 (N_13608,N_10196,N_9903);
nand U13609 (N_13609,N_9691,N_11784);
nand U13610 (N_13610,N_9043,N_11913);
and U13611 (N_13611,N_10036,N_7254);
nor U13612 (N_13612,N_8016,N_7677);
nor U13613 (N_13613,N_11761,N_8722);
nor U13614 (N_13614,N_9693,N_11456);
or U13615 (N_13615,N_7204,N_8688);
or U13616 (N_13616,N_11051,N_8138);
nor U13617 (N_13617,N_11160,N_6810);
nand U13618 (N_13618,N_7793,N_10387);
or U13619 (N_13619,N_9823,N_7804);
nor U13620 (N_13620,N_9988,N_6517);
xor U13621 (N_13621,N_9843,N_9160);
nand U13622 (N_13622,N_9333,N_6804);
or U13623 (N_13623,N_9559,N_10616);
or U13624 (N_13624,N_9557,N_11516);
or U13625 (N_13625,N_6256,N_6107);
and U13626 (N_13626,N_9671,N_9980);
or U13627 (N_13627,N_9080,N_6072);
or U13628 (N_13628,N_8826,N_7320);
and U13629 (N_13629,N_8414,N_9850);
and U13630 (N_13630,N_7972,N_10593);
nand U13631 (N_13631,N_8212,N_10789);
nand U13632 (N_13632,N_7182,N_11662);
nand U13633 (N_13633,N_8087,N_10854);
nand U13634 (N_13634,N_9581,N_6779);
and U13635 (N_13635,N_8970,N_9081);
or U13636 (N_13636,N_8371,N_8697);
or U13637 (N_13637,N_7041,N_6944);
or U13638 (N_13638,N_8214,N_6286);
nand U13639 (N_13639,N_11535,N_8862);
or U13640 (N_13640,N_6073,N_7947);
xor U13641 (N_13641,N_8668,N_7363);
xor U13642 (N_13642,N_7879,N_8945);
and U13643 (N_13643,N_7650,N_9402);
and U13644 (N_13644,N_7493,N_9207);
and U13645 (N_13645,N_11196,N_7319);
and U13646 (N_13646,N_10554,N_6654);
and U13647 (N_13647,N_7372,N_11947);
and U13648 (N_13648,N_9686,N_7278);
nand U13649 (N_13649,N_10468,N_10958);
nor U13650 (N_13650,N_6764,N_10138);
nand U13651 (N_13651,N_7513,N_11049);
nor U13652 (N_13652,N_10978,N_11618);
or U13653 (N_13653,N_6384,N_8171);
xor U13654 (N_13654,N_9896,N_6556);
xor U13655 (N_13655,N_11743,N_10207);
nor U13656 (N_13656,N_10828,N_7604);
nor U13657 (N_13657,N_6228,N_7265);
or U13658 (N_13658,N_6581,N_10118);
or U13659 (N_13659,N_8247,N_7227);
and U13660 (N_13660,N_6952,N_8319);
or U13661 (N_13661,N_6694,N_9951);
nor U13662 (N_13662,N_6239,N_8663);
xor U13663 (N_13663,N_7494,N_11138);
or U13664 (N_13664,N_6751,N_9440);
xnor U13665 (N_13665,N_10147,N_6634);
or U13666 (N_13666,N_10776,N_10550);
or U13667 (N_13667,N_6644,N_8973);
or U13668 (N_13668,N_6271,N_11910);
nor U13669 (N_13669,N_6742,N_6610);
nand U13670 (N_13670,N_9296,N_11844);
nand U13671 (N_13671,N_9683,N_8789);
nand U13672 (N_13672,N_6651,N_6240);
nand U13673 (N_13673,N_10753,N_7915);
or U13674 (N_13674,N_10122,N_6749);
and U13675 (N_13675,N_9871,N_9185);
nand U13676 (N_13676,N_11711,N_11949);
nand U13677 (N_13677,N_10653,N_6112);
and U13678 (N_13678,N_11417,N_7410);
xor U13679 (N_13679,N_10830,N_8029);
nand U13680 (N_13680,N_8463,N_8580);
xor U13681 (N_13681,N_8278,N_10517);
nand U13682 (N_13682,N_11699,N_10234);
xnor U13683 (N_13683,N_9362,N_8255);
nand U13684 (N_13684,N_10336,N_11087);
nand U13685 (N_13685,N_11878,N_6924);
and U13686 (N_13686,N_7818,N_10880);
nor U13687 (N_13687,N_11986,N_10310);
or U13688 (N_13688,N_10932,N_9732);
nor U13689 (N_13689,N_10158,N_8320);
and U13690 (N_13690,N_9555,N_10705);
xor U13691 (N_13691,N_11579,N_8489);
nor U13692 (N_13692,N_7711,N_7579);
or U13693 (N_13693,N_7835,N_8344);
xnor U13694 (N_13694,N_8678,N_8342);
or U13695 (N_13695,N_7926,N_6797);
and U13696 (N_13696,N_7189,N_11708);
nand U13697 (N_13697,N_10277,N_6773);
nor U13698 (N_13698,N_11687,N_9420);
xor U13699 (N_13699,N_9095,N_6965);
nor U13700 (N_13700,N_9814,N_6903);
and U13701 (N_13701,N_7180,N_6657);
nor U13702 (N_13702,N_9593,N_8626);
and U13703 (N_13703,N_9527,N_10268);
nand U13704 (N_13704,N_11103,N_11595);
and U13705 (N_13705,N_10096,N_10747);
nor U13706 (N_13706,N_11060,N_11779);
nor U13707 (N_13707,N_6906,N_8634);
nand U13708 (N_13708,N_9545,N_7125);
and U13709 (N_13709,N_11543,N_11730);
and U13710 (N_13710,N_8328,N_6411);
or U13711 (N_13711,N_9812,N_8071);
nand U13712 (N_13712,N_8085,N_11994);
nor U13713 (N_13713,N_9273,N_10479);
and U13714 (N_13714,N_7977,N_9758);
nand U13715 (N_13715,N_8638,N_8349);
nor U13716 (N_13716,N_11623,N_6291);
nand U13717 (N_13717,N_11679,N_7368);
nor U13718 (N_13718,N_11433,N_7516);
nor U13719 (N_13719,N_11401,N_10435);
nor U13720 (N_13720,N_6733,N_6044);
or U13721 (N_13721,N_8242,N_11059);
or U13722 (N_13722,N_6571,N_11984);
or U13723 (N_13723,N_6513,N_10301);
or U13724 (N_13724,N_9194,N_6330);
and U13725 (N_13725,N_11782,N_6097);
nor U13726 (N_13726,N_7559,N_7337);
or U13727 (N_13727,N_11640,N_6826);
nand U13728 (N_13728,N_10908,N_11962);
xor U13729 (N_13729,N_8065,N_11211);
or U13730 (N_13730,N_6597,N_11463);
xnor U13731 (N_13731,N_7387,N_9319);
and U13732 (N_13732,N_10313,N_9790);
xnor U13733 (N_13733,N_6987,N_10764);
and U13734 (N_13734,N_11628,N_8806);
nor U13735 (N_13735,N_10955,N_9515);
and U13736 (N_13736,N_6579,N_9283);
and U13737 (N_13737,N_9263,N_11004);
xnor U13738 (N_13738,N_8040,N_9516);
nand U13739 (N_13739,N_8954,N_9028);
nand U13740 (N_13740,N_8089,N_6130);
nor U13741 (N_13741,N_7660,N_6178);
nand U13742 (N_13742,N_7126,N_6187);
nand U13743 (N_13743,N_7776,N_6911);
or U13744 (N_13744,N_11897,N_11131);
nor U13745 (N_13745,N_6090,N_10353);
nor U13746 (N_13746,N_9882,N_10561);
nand U13747 (N_13747,N_11518,N_8883);
xnor U13748 (N_13748,N_8729,N_7713);
nand U13749 (N_13749,N_10765,N_6269);
nor U13750 (N_13750,N_6307,N_8333);
nand U13751 (N_13751,N_8490,N_10436);
nand U13752 (N_13752,N_6645,N_10892);
nor U13753 (N_13753,N_11661,N_9012);
and U13754 (N_13754,N_11411,N_11781);
nand U13755 (N_13755,N_10367,N_11070);
or U13756 (N_13756,N_11139,N_7810);
and U13757 (N_13757,N_8237,N_8257);
nor U13758 (N_13758,N_7566,N_7066);
or U13759 (N_13759,N_10939,N_7307);
xnor U13760 (N_13760,N_6261,N_11636);
nand U13761 (N_13761,N_7799,N_9695);
and U13762 (N_13762,N_8934,N_8757);
nor U13763 (N_13763,N_6662,N_8810);
nand U13764 (N_13764,N_9392,N_8309);
or U13765 (N_13765,N_11473,N_8232);
and U13766 (N_13766,N_11566,N_11036);
and U13767 (N_13767,N_6516,N_8980);
or U13768 (N_13768,N_10167,N_7071);
xor U13769 (N_13769,N_11583,N_8492);
or U13770 (N_13770,N_7832,N_8142);
nor U13771 (N_13771,N_11375,N_7355);
nand U13772 (N_13772,N_6287,N_7865);
and U13773 (N_13773,N_10549,N_7505);
and U13774 (N_13774,N_7366,N_10745);
nor U13775 (N_13775,N_10672,N_11899);
xor U13776 (N_13776,N_10839,N_11133);
and U13777 (N_13777,N_11166,N_11399);
or U13778 (N_13778,N_6504,N_11164);
nor U13779 (N_13779,N_8209,N_8323);
and U13780 (N_13780,N_6049,N_8784);
and U13781 (N_13781,N_7258,N_10840);
nor U13782 (N_13782,N_10377,N_8331);
nand U13783 (N_13783,N_11604,N_7430);
or U13784 (N_13784,N_9395,N_6862);
nand U13785 (N_13785,N_9223,N_6374);
nor U13786 (N_13786,N_10123,N_11559);
nand U13787 (N_13787,N_7332,N_7861);
or U13788 (N_13788,N_10947,N_11167);
xnor U13789 (N_13789,N_11627,N_11084);
and U13790 (N_13790,N_10865,N_7253);
or U13791 (N_13791,N_9712,N_11418);
or U13792 (N_13792,N_6566,N_8015);
nor U13793 (N_13793,N_9033,N_9050);
or U13794 (N_13794,N_6443,N_9182);
nand U13795 (N_13795,N_7546,N_11361);
or U13796 (N_13796,N_11179,N_7338);
nand U13797 (N_13797,N_11237,N_7169);
nor U13798 (N_13798,N_9110,N_7060);
nand U13799 (N_13799,N_11577,N_8156);
nand U13800 (N_13800,N_7993,N_9071);
nand U13801 (N_13801,N_7304,N_8318);
or U13802 (N_13802,N_10002,N_10031);
and U13803 (N_13803,N_10150,N_7205);
xnor U13804 (N_13804,N_6712,N_7584);
and U13805 (N_13805,N_11359,N_10385);
and U13806 (N_13806,N_9441,N_6379);
nor U13807 (N_13807,N_6120,N_10577);
nand U13808 (N_13808,N_7692,N_11100);
and U13809 (N_13809,N_6064,N_11659);
nand U13810 (N_13810,N_8577,N_11835);
or U13811 (N_13811,N_9092,N_9434);
and U13812 (N_13812,N_8794,N_7244);
and U13813 (N_13813,N_6472,N_9895);
and U13814 (N_13814,N_6420,N_11904);
nor U13815 (N_13815,N_8002,N_6192);
nand U13816 (N_13816,N_9614,N_6381);
xor U13817 (N_13817,N_7171,N_7090);
nor U13818 (N_13818,N_9647,N_10237);
nand U13819 (N_13819,N_6179,N_6945);
or U13820 (N_13820,N_7859,N_9116);
nand U13821 (N_13821,N_11965,N_11624);
nor U13822 (N_13822,N_6265,N_6613);
nand U13823 (N_13823,N_10662,N_10811);
nor U13824 (N_13824,N_10197,N_8889);
and U13825 (N_13825,N_9761,N_7758);
and U13826 (N_13826,N_8896,N_11876);
or U13827 (N_13827,N_8295,N_11958);
and U13828 (N_13828,N_11400,N_9054);
and U13829 (N_13829,N_8975,N_6433);
nand U13830 (N_13830,N_6679,N_7303);
and U13831 (N_13831,N_10295,N_6321);
or U13832 (N_13832,N_9428,N_10087);
and U13833 (N_13833,N_10645,N_10562);
xor U13834 (N_13834,N_11056,N_10715);
and U13835 (N_13835,N_10426,N_7588);
or U13836 (N_13836,N_8786,N_9278);
and U13837 (N_13837,N_6200,N_11671);
and U13838 (N_13838,N_7686,N_8624);
and U13839 (N_13839,N_11286,N_9933);
xor U13840 (N_13840,N_11851,N_8920);
xor U13841 (N_13841,N_9224,N_8543);
nor U13842 (N_13842,N_8470,N_7903);
nand U13843 (N_13843,N_8912,N_10998);
and U13844 (N_13844,N_7630,N_6692);
nor U13845 (N_13845,N_7953,N_11884);
nor U13846 (N_13846,N_11888,N_11959);
or U13847 (N_13847,N_6547,N_10292);
and U13848 (N_13848,N_9374,N_6728);
nand U13849 (N_13849,N_10008,N_10169);
and U13850 (N_13850,N_8747,N_9944);
nand U13851 (N_13851,N_10223,N_10626);
nand U13852 (N_13852,N_7067,N_9410);
and U13853 (N_13853,N_11819,N_9342);
nor U13854 (N_13854,N_9924,N_6226);
nand U13855 (N_13855,N_10180,N_9091);
or U13856 (N_13856,N_6707,N_10513);
or U13857 (N_13857,N_6288,N_6143);
or U13858 (N_13858,N_8745,N_6294);
nand U13859 (N_13859,N_10389,N_8052);
nor U13860 (N_13860,N_9831,N_6154);
or U13861 (N_13861,N_8399,N_11213);
nand U13862 (N_13862,N_8654,N_8691);
nor U13863 (N_13863,N_8684,N_11655);
nand U13864 (N_13864,N_11191,N_11028);
nor U13865 (N_13865,N_9520,N_11553);
or U13866 (N_13866,N_10102,N_6479);
xor U13867 (N_13867,N_10411,N_10400);
and U13868 (N_13868,N_10466,N_11842);
and U13869 (N_13869,N_9617,N_11669);
and U13870 (N_13870,N_8139,N_8111);
nand U13871 (N_13871,N_11596,N_8716);
nor U13872 (N_13872,N_10214,N_7425);
nor U13873 (N_13873,N_8687,N_6464);
or U13874 (N_13874,N_7114,N_9770);
and U13875 (N_13875,N_7435,N_7174);
and U13876 (N_13876,N_9531,N_11825);
and U13877 (N_13877,N_10399,N_7735);
and U13878 (N_13878,N_11887,N_9206);
or U13879 (N_13879,N_7299,N_6631);
nor U13880 (N_13880,N_7477,N_10859);
nor U13881 (N_13881,N_7292,N_6954);
or U13882 (N_13882,N_10699,N_10454);
nand U13883 (N_13883,N_9163,N_10579);
nand U13884 (N_13884,N_10915,N_9662);
and U13885 (N_13885,N_7035,N_7769);
nor U13886 (N_13886,N_9246,N_9649);
nor U13887 (N_13887,N_10245,N_9974);
xnor U13888 (N_13888,N_11354,N_7699);
or U13889 (N_13889,N_10605,N_10027);
nand U13890 (N_13890,N_8090,N_10771);
nor U13891 (N_13891,N_7674,N_9875);
nor U13892 (N_13892,N_8061,N_10800);
nor U13893 (N_13893,N_11615,N_8378);
or U13894 (N_13894,N_6455,N_11109);
and U13895 (N_13895,N_6278,N_8899);
or U13896 (N_13896,N_6121,N_11249);
nand U13897 (N_13897,N_7860,N_10531);
xor U13898 (N_13898,N_9354,N_6365);
and U13899 (N_13899,N_11588,N_6268);
nor U13900 (N_13900,N_11854,N_6030);
nor U13901 (N_13901,N_8983,N_10241);
or U13902 (N_13902,N_6491,N_9506);
and U13903 (N_13903,N_10523,N_10151);
xnor U13904 (N_13904,N_9788,N_7973);
or U13905 (N_13905,N_8692,N_6250);
nor U13906 (N_13906,N_10514,N_6838);
and U13907 (N_13907,N_8312,N_7201);
xnor U13908 (N_13908,N_7176,N_6689);
or U13909 (N_13909,N_8113,N_10944);
and U13910 (N_13910,N_9190,N_10721);
and U13911 (N_13911,N_11554,N_10219);
and U13912 (N_13912,N_7471,N_6604);
or U13913 (N_13913,N_8550,N_6962);
and U13914 (N_13914,N_7190,N_6462);
or U13915 (N_13915,N_11770,N_11314);
or U13916 (N_13916,N_7570,N_11530);
and U13917 (N_13917,N_9062,N_8384);
nand U13918 (N_13918,N_10950,N_6730);
nor U13919 (N_13919,N_8451,N_11118);
nor U13920 (N_13920,N_7269,N_11002);
nor U13921 (N_13921,N_6251,N_9552);
nand U13922 (N_13922,N_7287,N_11701);
nand U13923 (N_13923,N_9972,N_6259);
or U13924 (N_13924,N_9023,N_10928);
or U13925 (N_13925,N_7029,N_9285);
and U13926 (N_13926,N_6669,N_10271);
nor U13927 (N_13927,N_8115,N_8464);
or U13928 (N_13928,N_6487,N_6083);
and U13929 (N_13929,N_8797,N_6126);
and U13930 (N_13930,N_11127,N_8772);
or U13931 (N_13931,N_10786,N_10422);
nand U13932 (N_13932,N_9004,N_6785);
or U13933 (N_13933,N_7340,N_8106);
or U13934 (N_13934,N_7406,N_8976);
nand U13935 (N_13935,N_6722,N_10308);
and U13936 (N_13936,N_6587,N_11728);
and U13937 (N_13937,N_6636,N_10951);
and U13938 (N_13938,N_7397,N_8300);
nor U13939 (N_13939,N_7085,N_8009);
and U13940 (N_13940,N_11644,N_7021);
nor U13941 (N_13941,N_11602,N_8223);
and U13942 (N_13942,N_8375,N_9979);
or U13943 (N_13943,N_6955,N_10266);
or U13944 (N_13944,N_9394,N_10570);
nand U13945 (N_13945,N_8683,N_7928);
and U13946 (N_13946,N_9866,N_11794);
or U13947 (N_13947,N_9863,N_10256);
or U13948 (N_13948,N_7478,N_6754);
and U13949 (N_13949,N_10983,N_9618);
and U13950 (N_13950,N_11223,N_11605);
and U13951 (N_13951,N_7532,N_8627);
or U13952 (N_13952,N_7096,N_10621);
nor U13953 (N_13953,N_9763,N_9276);
xnor U13954 (N_13954,N_6156,N_10588);
xnor U13955 (N_13955,N_11532,N_10784);
or U13956 (N_13956,N_10212,N_8093);
nand U13957 (N_13957,N_11981,N_8327);
and U13958 (N_13958,N_7261,N_9245);
and U13959 (N_13959,N_8129,N_8744);
nor U13960 (N_13960,N_8070,N_8352);
nand U13961 (N_13961,N_9328,N_9665);
and U13962 (N_13962,N_10235,N_11356);
and U13963 (N_13963,N_10895,N_11823);
or U13964 (N_13964,N_9433,N_11478);
or U13965 (N_13965,N_8723,N_9723);
or U13966 (N_13966,N_8655,N_11350);
nor U13967 (N_13967,N_7549,N_8837);
or U13968 (N_13968,N_10936,N_10878);
and U13969 (N_13969,N_7142,N_9679);
and U13970 (N_13970,N_7954,N_6070);
nand U13971 (N_13971,N_9176,N_9250);
xor U13972 (N_13972,N_6071,N_10862);
xor U13973 (N_13973,N_7407,N_9534);
xor U13974 (N_13974,N_10168,N_10615);
nor U13975 (N_13975,N_8911,N_11406);
nor U13976 (N_13976,N_7897,N_7567);
or U13977 (N_13977,N_6283,N_9461);
and U13978 (N_13978,N_7930,N_11670);
and U13979 (N_13979,N_10803,N_7091);
nand U13980 (N_13980,N_6974,N_6582);
xnor U13981 (N_13981,N_9478,N_11090);
nor U13982 (N_13982,N_9331,N_11834);
nor U13983 (N_13983,N_8589,N_10361);
nor U13984 (N_13984,N_7380,N_7419);
nor U13985 (N_13985,N_7140,N_8117);
or U13986 (N_13986,N_7437,N_8126);
nor U13987 (N_13987,N_6919,N_6572);
nor U13988 (N_13988,N_6055,N_10067);
nor U13989 (N_13989,N_8236,N_10487);
nor U13990 (N_13990,N_9474,N_11649);
nand U13991 (N_13991,N_9530,N_6320);
or U13992 (N_13992,N_8164,N_11657);
nand U13993 (N_13993,N_11066,N_10233);
and U13994 (N_13994,N_8673,N_9131);
or U13995 (N_13995,N_7422,N_8872);
nand U13996 (N_13996,N_8279,N_11111);
and U13997 (N_13997,N_10961,N_6314);
nand U13998 (N_13998,N_7224,N_7787);
xor U13999 (N_13999,N_6417,N_11077);
and U14000 (N_14000,N_6527,N_11259);
nor U14001 (N_14001,N_11906,N_11448);
nand U14002 (N_14002,N_11940,N_6790);
and U14003 (N_14003,N_11481,N_8124);
or U14004 (N_14004,N_6039,N_6453);
nand U14005 (N_14005,N_9449,N_10536);
nand U14006 (N_14006,N_8267,N_7331);
xnor U14007 (N_14007,N_7685,N_6436);
or U14008 (N_14008,N_7780,N_8203);
and U14009 (N_14009,N_9800,N_10601);
nor U14010 (N_14010,N_8469,N_11137);
or U14011 (N_14011,N_9859,N_9810);
and U14012 (N_14012,N_11866,N_9287);
and U14013 (N_14013,N_8762,N_11378);
nor U14014 (N_14014,N_9260,N_10254);
nand U14015 (N_14015,N_9363,N_8984);
nand U14016 (N_14016,N_9167,N_8356);
and U14017 (N_14017,N_6415,N_8177);
nand U14018 (N_14018,N_8392,N_11319);
or U14019 (N_14019,N_10802,N_10294);
nand U14020 (N_14020,N_8957,N_10322);
nand U14021 (N_14021,N_8372,N_7185);
nor U14022 (N_14022,N_9072,N_6726);
nor U14023 (N_14023,N_9239,N_6616);
nand U14024 (N_14024,N_6482,N_7705);
nand U14025 (N_14025,N_9635,N_7046);
nand U14026 (N_14026,N_8639,N_6788);
nand U14027 (N_14027,N_8907,N_10748);
xor U14028 (N_14028,N_9568,N_11055);
nor U14029 (N_14029,N_7504,N_11642);
or U14030 (N_14030,N_11506,N_9121);
or U14031 (N_14031,N_8777,N_8234);
and U14032 (N_14032,N_10267,N_6611);
and U14033 (N_14033,N_10324,N_9801);
or U14034 (N_14034,N_10918,N_8324);
nand U14035 (N_14035,N_9305,N_7389);
nand U14036 (N_14036,N_6656,N_10835);
and U14037 (N_14037,N_10723,N_6868);
nor U14038 (N_14038,N_11896,N_7005);
nor U14039 (N_14039,N_9145,N_9061);
or U14040 (N_14040,N_8606,N_11376);
nor U14041 (N_14041,N_10495,N_9996);
nand U14042 (N_14042,N_9208,N_7512);
and U14043 (N_14043,N_9992,N_9901);
or U14044 (N_14044,N_10076,N_7281);
nor U14045 (N_14045,N_7164,N_11130);
nor U14046 (N_14046,N_6828,N_9344);
or U14047 (N_14047,N_11176,N_11472);
or U14048 (N_14048,N_10204,N_9675);
nor U14049 (N_14049,N_10546,N_6014);
xnor U14050 (N_14050,N_10834,N_7013);
nor U14051 (N_14051,N_9934,N_7937);
nand U14052 (N_14052,N_9272,N_10369);
nor U14053 (N_14053,N_8311,N_9166);
nand U14054 (N_14054,N_9355,N_7904);
nor U14055 (N_14055,N_10960,N_7495);
nor U14056 (N_14056,N_10708,N_7906);
or U14057 (N_14057,N_10458,N_6748);
xnor U14058 (N_14058,N_7417,N_10867);
nor U14059 (N_14059,N_6811,N_9438);
and U14060 (N_14060,N_7766,N_6575);
and U14061 (N_14061,N_11621,N_10129);
nand U14062 (N_14062,N_10269,N_9795);
nor U14063 (N_14063,N_6442,N_10469);
xnor U14064 (N_14064,N_11439,N_11891);
and U14065 (N_14065,N_7416,N_9391);
or U14066 (N_14066,N_9435,N_10646);
and U14067 (N_14067,N_7552,N_9076);
nand U14068 (N_14068,N_9743,N_6114);
and U14069 (N_14069,N_9217,N_11096);
or U14070 (N_14070,N_6317,N_7748);
and U14071 (N_14071,N_8710,N_6207);
or U14072 (N_14072,N_10059,N_8871);
nor U14073 (N_14073,N_11218,N_9862);
and U14074 (N_14074,N_6169,N_7432);
nor U14075 (N_14075,N_7445,N_10894);
or U14076 (N_14076,N_9431,N_8599);
nand U14077 (N_14077,N_8291,N_7459);
and U14078 (N_14078,N_10889,N_9905);
nor U14079 (N_14079,N_7050,N_9651);
nand U14080 (N_14080,N_11552,N_6624);
or U14081 (N_14081,N_7551,N_11088);
nand U14082 (N_14082,N_7785,N_7910);
nand U14083 (N_14083,N_8169,N_10871);
or U14084 (N_14084,N_8519,N_11086);
or U14085 (N_14085,N_7620,N_6094);
xnor U14086 (N_14086,N_9606,N_9977);
and U14087 (N_14087,N_8425,N_7146);
nand U14088 (N_14088,N_11296,N_10757);
or U14089 (N_14089,N_11753,N_8043);
nand U14090 (N_14090,N_10373,N_11124);
nand U14091 (N_14091,N_6354,N_10693);
or U14092 (N_14092,N_10744,N_6289);
or U14093 (N_14093,N_11804,N_7175);
nand U14094 (N_14094,N_10592,N_7682);
nand U14095 (N_14095,N_9138,N_9808);
nand U14096 (N_14096,N_10125,N_6825);
or U14097 (N_14097,N_7120,N_8167);
nor U14098 (N_14098,N_6763,N_8260);
and U14099 (N_14099,N_7967,N_8857);
and U14100 (N_14100,N_7247,N_9779);
nor U14101 (N_14101,N_11547,N_6148);
and U14102 (N_14102,N_11001,N_10652);
nand U14103 (N_14103,N_7917,N_8094);
or U14104 (N_14104,N_7008,N_6829);
or U14105 (N_14105,N_6204,N_11998);
nand U14106 (N_14106,N_7651,N_11691);
nand U14107 (N_14107,N_9817,N_10881);
or U14108 (N_14108,N_6276,N_11454);
nand U14109 (N_14109,N_7625,N_7825);
nor U14110 (N_14110,N_6573,N_7542);
nor U14111 (N_14111,N_9219,N_7610);
xor U14112 (N_14112,N_11414,N_9930);
nand U14113 (N_14113,N_10688,N_10920);
nand U14114 (N_14114,N_8916,N_8583);
nor U14115 (N_14115,N_10778,N_6820);
nor U14116 (N_14116,N_6000,N_10449);
or U14117 (N_14117,N_7241,N_10954);
nor U14118 (N_14118,N_7230,N_9991);
nor U14119 (N_14119,N_7883,N_9574);
nand U14120 (N_14120,N_8867,N_10349);
nor U14121 (N_14121,N_11474,N_10543);
nor U14122 (N_14122,N_10607,N_11966);
or U14123 (N_14123,N_6357,N_6918);
xor U14124 (N_14124,N_7537,N_8493);
or U14125 (N_14125,N_8981,N_11027);
or U14126 (N_14126,N_11945,N_7128);
nor U14127 (N_14127,N_7426,N_11294);
xnor U14128 (N_14128,N_11853,N_10095);
nor U14129 (N_14129,N_9353,N_6990);
or U14130 (N_14130,N_7137,N_8677);
and U14131 (N_14131,N_10314,N_8135);
nor U14132 (N_14132,N_10255,N_8665);
nand U14133 (N_14133,N_9846,N_11953);
nand U14134 (N_14134,N_9773,N_8077);
nor U14135 (N_14135,N_11290,N_8647);
and U14136 (N_14136,N_7007,N_10452);
nor U14137 (N_14137,N_11113,N_11694);
or U14138 (N_14138,N_11989,N_7006);
xnor U14139 (N_14139,N_7873,N_8033);
and U14140 (N_14140,N_10842,N_8892);
nand U14141 (N_14141,N_8227,N_10815);
xor U14142 (N_14142,N_11593,N_7544);
and U14143 (N_14143,N_9168,N_8593);
nand U14144 (N_14144,N_6019,N_6731);
nand U14145 (N_14145,N_11591,N_8428);
nor U14146 (N_14146,N_7959,N_8078);
or U14147 (N_14147,N_7260,N_11189);
nand U14148 (N_14148,N_10142,N_10300);
nand U14149 (N_14149,N_7575,N_11663);
nor U14150 (N_14150,N_9228,N_11107);
nand U14151 (N_14151,N_10444,N_6907);
nor U14152 (N_14152,N_8958,N_10433);
nand U14153 (N_14153,N_10222,N_6035);
or U14154 (N_14154,N_11507,N_8004);
or U14155 (N_14155,N_7489,N_7327);
nor U14156 (N_14156,N_10996,N_8302);
nor U14157 (N_14157,N_8579,N_10409);
nor U14158 (N_14158,N_6860,N_10503);
nor U14159 (N_14159,N_10545,N_11326);
and U14160 (N_14160,N_7051,N_9632);
nand U14161 (N_14161,N_7468,N_10860);
nand U14162 (N_14162,N_9495,N_7421);
xnor U14163 (N_14163,N_8953,N_11766);
and U14164 (N_14164,N_10144,N_8268);
nand U14165 (N_14165,N_6100,N_6565);
nor U14166 (N_14166,N_6496,N_9316);
nor U14167 (N_14167,N_9266,N_8629);
or U14168 (N_14168,N_10121,N_11434);
and U14169 (N_14169,N_9065,N_11485);
or U14170 (N_14170,N_7764,N_8329);
and U14171 (N_14171,N_8357,N_8145);
nor U14172 (N_14172,N_7795,N_10084);
nor U14173 (N_14173,N_10111,N_7732);
nor U14174 (N_14174,N_8251,N_6629);
and U14175 (N_14175,N_6564,N_6356);
nor U14176 (N_14176,N_9521,N_8674);
or U14177 (N_14177,N_10110,N_7974);
or U14178 (N_14178,N_11260,N_9406);
or U14179 (N_14179,N_11538,N_11447);
and U14180 (N_14180,N_9542,N_6264);
xor U14181 (N_14181,N_6432,N_11304);
nand U14182 (N_14182,N_11650,N_7964);
nand U14183 (N_14183,N_9794,N_11902);
nor U14184 (N_14184,N_7348,N_10376);
nor U14185 (N_14185,N_6448,N_6716);
and U14186 (N_14186,N_10994,N_11988);
nand U14187 (N_14187,N_6735,N_9129);
nand U14188 (N_14188,N_8153,N_7100);
or U14189 (N_14189,N_8609,N_11328);
nor U14190 (N_14190,N_6013,N_9171);
nor U14191 (N_14191,N_7276,N_10475);
nor U14192 (N_14192,N_8181,N_8690);
or U14193 (N_14193,N_11783,N_7403);
or U14194 (N_14194,N_11187,N_7472);
xnor U14195 (N_14195,N_6331,N_10394);
nor U14196 (N_14196,N_10686,N_6372);
and U14197 (N_14197,N_7729,N_6993);
nand U14198 (N_14198,N_9998,N_6793);
and U14199 (N_14199,N_8782,N_7798);
or U14200 (N_14200,N_8846,N_10352);
nand U14201 (N_14201,N_9465,N_8417);
and U14202 (N_14202,N_10229,N_8895);
nand U14203 (N_14203,N_11826,N_6128);
or U14204 (N_14204,N_10103,N_9659);
and U14205 (N_14205,N_11108,N_9625);
nor U14206 (N_14206,N_8581,N_9745);
nand U14207 (N_14207,N_9548,N_10332);
xor U14208 (N_14208,N_7476,N_7049);
nand U14209 (N_14209,N_8012,N_6345);
nor U14210 (N_14210,N_11020,N_9881);
and U14211 (N_14211,N_8204,N_8419);
or U14212 (N_14212,N_9146,N_10141);
nand U14213 (N_14213,N_6851,N_11046);
nor U14214 (N_14214,N_7728,N_6089);
xnor U14215 (N_14215,N_8199,N_10408);
xnor U14216 (N_14216,N_11491,N_10898);
nand U14217 (N_14217,N_7653,N_10916);
nand U14218 (N_14218,N_8276,N_7106);
nor U14219 (N_14219,N_8965,N_9612);
or U14220 (N_14220,N_9603,N_7112);
and U14221 (N_14221,N_7423,N_11840);
nand U14222 (N_14222,N_10633,N_9087);
nor U14223 (N_14223,N_9313,N_9676);
or U14224 (N_14224,N_7187,N_7663);
and U14225 (N_14225,N_8607,N_8072);
nor U14226 (N_14226,N_6666,N_8869);
or U14227 (N_14227,N_9153,N_10649);
or U14228 (N_14228,N_8410,N_11707);
nor U14229 (N_14229,N_6806,N_9191);
or U14230 (N_14230,N_6979,N_7252);
and U14231 (N_14231,N_6709,N_11386);
or U14232 (N_14232,N_10485,N_8426);
nor U14233 (N_14233,N_9115,N_7961);
nand U14234 (N_14234,N_8254,N_6643);
and U14235 (N_14235,N_10581,N_9447);
or U14236 (N_14236,N_9865,N_10100);
and U14237 (N_14237,N_11520,N_7726);
nand U14238 (N_14238,N_9715,N_10725);
and U14239 (N_14239,N_10934,N_6893);
or U14240 (N_14240,N_6243,N_9769);
nand U14241 (N_14241,N_9382,N_8083);
xor U14242 (N_14242,N_8427,N_8350);
and U14243 (N_14243,N_8913,N_6681);
nand U14244 (N_14244,N_10684,N_6873);
and U14245 (N_14245,N_10756,N_11993);
and U14246 (N_14246,N_6461,N_9310);
or U14247 (N_14247,N_8137,N_8194);
and U14248 (N_14248,N_6795,N_11425);
or U14249 (N_14249,N_11159,N_6285);
or U14250 (N_14250,N_6985,N_8440);
or U14251 (N_14251,N_10946,N_10341);
nand U14252 (N_14252,N_7560,N_6129);
nor U14253 (N_14253,N_7058,N_10683);
nor U14254 (N_14254,N_8873,N_6502);
nor U14255 (N_14255,N_6699,N_6184);
or U14256 (N_14256,N_9737,N_11951);
nand U14257 (N_14257,N_11571,N_6137);
xnor U14258 (N_14258,N_6555,N_10128);
nand U14259 (N_14259,N_10760,N_6598);
nand U14260 (N_14260,N_11960,N_10465);
nor U14261 (N_14261,N_7836,N_6026);
and U14262 (N_14262,N_10383,N_9544);
and U14263 (N_14263,N_9491,N_11791);
nor U14264 (N_14264,N_6467,N_6633);
nand U14265 (N_14265,N_6640,N_10013);
nor U14266 (N_14266,N_10362,N_9202);
nand U14267 (N_14267,N_7016,N_10191);
xnor U14268 (N_14268,N_10003,N_8594);
nor U14269 (N_14269,N_11527,N_7662);
and U14270 (N_14270,N_10719,N_8900);
or U14271 (N_14271,N_6867,N_11668);
nand U14272 (N_14272,N_10302,N_11254);
nor U14273 (N_14273,N_10997,N_7767);
nand U14274 (N_14274,N_10796,N_8591);
nor U14275 (N_14275,N_9904,N_7017);
or U14276 (N_14276,N_6740,N_10116);
nand U14277 (N_14277,N_10798,N_7781);
nor U14278 (N_14278,N_9854,N_8631);
and U14279 (N_14279,N_9186,N_8567);
nor U14280 (N_14280,N_11226,N_6563);
and U14281 (N_14281,N_9646,N_6118);
nand U14282 (N_14282,N_6180,N_6698);
nor U14283 (N_14283,N_11143,N_10777);
and U14284 (N_14284,N_11261,N_8235);
or U14285 (N_14285,N_7362,N_6348);
and U14286 (N_14286,N_10055,N_8689);
nand U14287 (N_14287,N_7497,N_9022);
nand U14288 (N_14288,N_7571,N_11751);
or U14289 (N_14289,N_6511,N_8491);
and U14290 (N_14290,N_11147,N_6737);
and U14291 (N_14291,N_11908,N_11349);
xor U14292 (N_14292,N_10199,N_10236);
nand U14293 (N_14293,N_9910,N_10758);
nand U14294 (N_14294,N_7210,N_9750);
and U14295 (N_14295,N_11340,N_8024);
xor U14296 (N_14296,N_9125,N_11822);
nand U14297 (N_14297,N_11755,N_6951);
nor U14298 (N_14298,N_7155,N_7600);
nor U14299 (N_14299,N_10824,N_9700);
nand U14300 (N_14300,N_8878,N_7710);
nor U14301 (N_14301,N_8482,N_10731);
xor U14302 (N_14302,N_11190,N_7717);
nor U14303 (N_14303,N_6428,N_11360);
nor U14304 (N_14304,N_11805,N_10431);
and U14305 (N_14305,N_7675,N_9029);
and U14306 (N_14306,N_8149,N_11833);
or U14307 (N_14307,N_10136,N_11852);
nand U14308 (N_14308,N_7412,N_11098);
nor U14309 (N_14309,N_8661,N_6444);
nor U14310 (N_14310,N_11465,N_11362);
and U14311 (N_14311,N_6844,N_10540);
and U14312 (N_14312,N_11898,N_9386);
and U14313 (N_14313,N_6452,N_8831);
nor U14314 (N_14314,N_11977,N_7312);
nor U14315 (N_14315,N_11693,N_7028);
nand U14316 (N_14316,N_11629,N_7249);
nor U14317 (N_14317,N_7215,N_9742);
nand U14318 (N_14318,N_9878,N_10287);
or U14319 (N_14319,N_8646,N_8211);
xor U14320 (N_14320,N_10728,N_6926);
or U14321 (N_14321,N_7536,N_7652);
or U14322 (N_14322,N_8709,N_8439);
and U14323 (N_14323,N_9396,N_9312);
nand U14324 (N_14324,N_10724,N_10694);
nand U14325 (N_14325,N_7678,N_7718);
and U14326 (N_14326,N_7839,N_11653);
and U14327 (N_14327,N_10238,N_7968);
nor U14328 (N_14328,N_6997,N_7358);
nand U14329 (N_14329,N_9799,N_8585);
and U14330 (N_14330,N_7673,N_8656);
nor U14331 (N_14331,N_11443,N_9375);
xor U14332 (N_14332,N_9227,N_8069);
or U14333 (N_14333,N_9199,N_6046);
or U14334 (N_14334,N_6031,N_10505);
nor U14335 (N_14335,N_11135,N_9016);
or U14336 (N_14336,N_9599,N_11921);
nand U14337 (N_14337,N_11338,N_9822);
or U14338 (N_14338,N_10976,N_7843);
nor U14339 (N_14339,N_9748,N_11907);
nand U14340 (N_14340,N_8109,N_8815);
nor U14341 (N_14341,N_10249,N_9150);
nand U14342 (N_14342,N_11675,N_10734);
xor U14343 (N_14343,N_7122,N_10028);
or U14344 (N_14344,N_8456,N_7228);
nand U14345 (N_14345,N_8483,N_9040);
or U14346 (N_14346,N_9908,N_6971);
nand U14347 (N_14347,N_11062,N_8303);
or U14348 (N_14348,N_11918,N_10351);
nand U14349 (N_14349,N_9175,N_8595);
nor U14350 (N_14350,N_10364,N_8110);
and U14351 (N_14351,N_10209,N_8390);
and U14352 (N_14352,N_7619,N_11015);
xnor U14353 (N_14353,N_6536,N_9317);
and U14354 (N_14354,N_8374,N_9768);
nand U14355 (N_14355,N_7807,N_10952);
and U14356 (N_14356,N_10135,N_7188);
xnor U14357 (N_14357,N_11536,N_6853);
and U14358 (N_14358,N_11132,N_7156);
nor U14359 (N_14359,N_7884,N_9724);
and U14360 (N_14360,N_8367,N_11232);
nor U14361 (N_14361,N_9370,N_8698);
nor U14362 (N_14362,N_7365,N_11242);
and U14363 (N_14363,N_10897,N_6818);
nand U14364 (N_14364,N_11969,N_10711);
xnor U14365 (N_14365,N_11374,N_7593);
or U14366 (N_14366,N_10206,N_8996);
xnor U14367 (N_14367,N_8602,N_8765);
nand U14368 (N_14368,N_6449,N_8114);
or U14369 (N_14369,N_6580,N_8037);
nand U14370 (N_14370,N_9021,N_11367);
and U14371 (N_14371,N_8275,N_10589);
nand U14372 (N_14372,N_6685,N_10962);
or U14373 (N_14373,N_7283,N_6719);
and U14374 (N_14374,N_9560,N_8893);
and U14375 (N_14375,N_6932,N_9367);
nor U14376 (N_14376,N_9739,N_10642);
or U14377 (N_14377,N_6328,N_11656);
and U14378 (N_14378,N_6554,N_11616);
or U14379 (N_14379,N_6098,N_7004);
and U14380 (N_14380,N_9466,N_8633);
or U14381 (N_14381,N_11531,N_9731);
and U14382 (N_14382,N_7324,N_11721);
and U14383 (N_14383,N_10924,N_9848);
and U14384 (N_14384,N_9787,N_11863);
nand U14385 (N_14385,N_9020,N_7309);
or U14386 (N_14386,N_7042,N_7800);
and U14387 (N_14387,N_11611,N_7436);
nor U14388 (N_14388,N_10656,N_8501);
xor U14389 (N_14389,N_7528,N_10198);
nand U14390 (N_14390,N_7150,N_10870);
or U14391 (N_14391,N_7975,N_7473);
or U14392 (N_14392,N_10896,N_9416);
or U14393 (N_14393,N_8269,N_7170);
or U14394 (N_14394,N_10164,N_10163);
nand U14395 (N_14395,N_8348,N_7115);
nor U14396 (N_14396,N_6934,N_6561);
and U14397 (N_14397,N_11397,N_7296);
xnor U14398 (N_14398,N_10763,N_8582);
nor U14399 (N_14399,N_8055,N_7242);
or U14400 (N_14400,N_9044,N_7044);
or U14401 (N_14401,N_6194,N_10260);
or U14402 (N_14402,N_10001,N_6704);
nand U14403 (N_14403,N_6210,N_11479);
nand U14404 (N_14404,N_9192,N_6548);
or U14405 (N_14405,N_6085,N_8590);
or U14406 (N_14406,N_6488,N_8825);
nor U14407 (N_14407,N_7845,N_10033);
nor U14408 (N_14408,N_9572,N_10979);
nor U14409 (N_14409,N_9931,N_8146);
xor U14410 (N_14410,N_7846,N_7539);
nand U14411 (N_14411,N_7702,N_6359);
nor U14412 (N_14412,N_10323,N_8937);
nor U14413 (N_14413,N_6102,N_8411);
nor U14414 (N_14414,N_9088,N_9757);
nor U14415 (N_14415,N_8184,N_9526);
and U14416 (N_14416,N_8640,N_7802);
nor U14417 (N_14417,N_7336,N_7696);
nor U14418 (N_14418,N_10246,N_8099);
or U14419 (N_14419,N_9626,N_7479);
nor U14420 (N_14420,N_11277,N_8549);
nand U14421 (N_14421,N_9136,N_7827);
nor U14422 (N_14422,N_8756,N_8650);
nand U14423 (N_14423,N_10080,N_11560);
and U14424 (N_14424,N_8905,N_11715);
nor U14425 (N_14425,N_8613,N_9966);
xnor U14426 (N_14426,N_9554,N_7971);
nor U14427 (N_14427,N_7765,N_10044);
nor U14428 (N_14428,N_7794,N_7510);
nor U14429 (N_14429,N_10687,N_6591);
or U14430 (N_14430,N_7235,N_10273);
or U14431 (N_14431,N_8829,N_8693);
or U14432 (N_14432,N_9144,N_11264);
nand U14433 (N_14433,N_6272,N_9598);
or U14434 (N_14434,N_9423,N_6076);
nor U14435 (N_14435,N_7153,N_10069);
nand U14436 (N_14436,N_9458,N_11053);
nand U14437 (N_14437,N_10258,N_10497);
or U14438 (N_14438,N_6146,N_7526);
or U14439 (N_14439,N_6813,N_8712);
nor U14440 (N_14440,N_8498,N_7243);
xnor U14441 (N_14441,N_8343,N_8636);
nor U14442 (N_14442,N_9765,N_6497);
nand U14443 (N_14443,N_9373,N_8497);
nor U14444 (N_14444,N_11369,N_8540);
nor U14445 (N_14445,N_7306,N_11778);
and U14446 (N_14446,N_7484,N_11262);
and U14447 (N_14447,N_9879,N_10265);
nand U14448 (N_14448,N_9816,N_11922);
xor U14449 (N_14449,N_8430,N_9487);
nand U14450 (N_14450,N_11522,N_10456);
xor U14451 (N_14451,N_10541,N_11012);
nor U14452 (N_14452,N_10759,N_8736);
xnor U14453 (N_14453,N_11980,N_7485);
nand U14454 (N_14454,N_6791,N_7707);
nand U14455 (N_14455,N_10766,N_9752);
nor U14456 (N_14456,N_8407,N_9825);
nor U14457 (N_14457,N_6678,N_11281);
or U14458 (N_14458,N_11076,N_8103);
nor U14459 (N_14459,N_6721,N_8467);
nand U14460 (N_14460,N_9018,N_6617);
xor U14461 (N_14461,N_11610,N_7162);
nor U14462 (N_14462,N_9607,N_6373);
and U14463 (N_14463,N_10484,N_6711);
nor U14464 (N_14464,N_6483,N_8793);
or U14465 (N_14465,N_8308,N_7168);
nor U14466 (N_14466,N_6578,N_7262);
or U14467 (N_14467,N_9771,N_6067);
nand U14468 (N_14468,N_7834,N_6231);
nor U14469 (N_14469,N_8705,N_6344);
and U14470 (N_14470,N_8882,N_8118);
nor U14471 (N_14471,N_6775,N_8180);
nor U14472 (N_14472,N_6471,N_6522);
and U14473 (N_14473,N_9818,N_7263);
and U14474 (N_14474,N_11275,N_8301);
nand U14475 (N_14475,N_8369,N_9999);
or U14476 (N_14476,N_8851,N_7812);
xnor U14477 (N_14477,N_9586,N_11523);
or U14478 (N_14478,N_10024,N_6150);
nor U14479 (N_14479,N_8940,N_7882);
nand U14480 (N_14480,N_9660,N_10348);
and U14481 (N_14481,N_8018,N_8719);
and U14482 (N_14482,N_8383,N_11972);
nand U14483 (N_14483,N_11010,N_7877);
or U14484 (N_14484,N_9327,N_8452);
nand U14485 (N_14485,N_9976,N_6002);
or U14486 (N_14486,N_8330,N_10423);
nand U14487 (N_14487,N_6340,N_6724);
or U14488 (N_14488,N_7981,N_6438);
or U14489 (N_14489,N_7759,N_7750);
or U14490 (N_14490,N_8596,N_10995);
or U14491 (N_14491,N_8224,N_8531);
or U14492 (N_14492,N_7885,N_10343);
and U14493 (N_14493,N_11311,N_6407);
and U14494 (N_14494,N_10105,N_9288);
and U14495 (N_14495,N_6661,N_11706);
or U14496 (N_14496,N_9172,N_8703);
and U14497 (N_14497,N_6052,N_7469);
nor U14498 (N_14498,N_11773,N_8364);
nand U14499 (N_14499,N_11200,N_6567);
or U14500 (N_14500,N_11526,N_6481);
xor U14501 (N_14501,N_6756,N_6440);
nor U14502 (N_14502,N_8962,N_11915);
or U14503 (N_14503,N_6542,N_6528);
xor U14504 (N_14504,N_8720,N_10710);
nor U14505 (N_14505,N_10155,N_11371);
and U14506 (N_14506,N_8776,N_10838);
nand U14507 (N_14507,N_9348,N_10224);
nand U14508 (N_14508,N_10072,N_9838);
nand U14509 (N_14509,N_6846,N_7207);
or U14510 (N_14510,N_8125,N_9177);
or U14511 (N_14511,N_9464,N_11442);
nor U14512 (N_14512,N_11342,N_6324);
or U14513 (N_14513,N_10297,N_7869);
xor U14514 (N_14514,N_7386,N_11476);
nand U14515 (N_14515,N_11608,N_10491);
or U14516 (N_14516,N_9807,N_6015);
or U14517 (N_14517,N_10620,N_11724);
nor U14518 (N_14518,N_9069,N_6253);
and U14519 (N_14519,N_8031,N_7507);
nor U14520 (N_14520,N_6075,N_10907);
and U14521 (N_14521,N_7405,N_11717);
nor U14522 (N_14522,N_7056,N_11638);
nand U14523 (N_14523,N_8985,N_10093);
nand U14524 (N_14524,N_8632,N_8421);
or U14525 (N_14525,N_10664,N_8714);
or U14526 (N_14526,N_6614,N_6916);
and U14527 (N_14527,N_6922,N_10925);
nand U14528 (N_14528,N_6879,N_10315);
nor U14529 (N_14529,N_10316,N_6653);
or U14530 (N_14530,N_7999,N_6976);
xnor U14531 (N_14531,N_11173,N_8559);
nand U14532 (N_14532,N_6501,N_9341);
and U14533 (N_14533,N_6267,N_6054);
xnor U14534 (N_14534,N_10893,N_6969);
and U14535 (N_14535,N_10478,N_8514);
and U14536 (N_14536,N_10637,N_10967);
or U14537 (N_14537,N_7622,N_11672);
xnor U14538 (N_14538,N_6170,N_7123);
and U14539 (N_14539,N_6871,N_6859);
and U14540 (N_14540,N_7503,N_10977);
nand U14541 (N_14541,N_8769,N_7658);
and U14542 (N_14542,N_11208,N_8556);
nand U14543 (N_14543,N_7492,N_7888);
and U14544 (N_14544,N_10112,N_10858);
nand U14545 (N_14545,N_6003,N_8615);
and U14546 (N_14546,N_8220,N_7080);
and U14547 (N_14547,N_6500,N_7070);
and U14548 (N_14548,N_8948,N_10972);
and U14549 (N_14549,N_11911,N_9252);
or U14550 (N_14550,N_7239,N_9685);
or U14551 (N_14551,N_6850,N_6670);
nand U14552 (N_14552,N_7089,N_10511);
nand U14553 (N_14553,N_9828,N_10262);
nand U14554 (N_14554,N_11117,N_11363);
nand U14555 (N_14555,N_8685,N_11639);
nor U14556 (N_14556,N_8025,N_7596);
or U14557 (N_14557,N_9894,N_10430);
nand U14558 (N_14558,N_6378,N_6001);
and U14559 (N_14559,N_8097,N_8304);
and U14560 (N_14560,N_6375,N_9853);
nand U14561 (N_14561,N_7083,N_11165);
or U14562 (N_14562,N_6385,N_11042);
or U14563 (N_14563,N_7172,N_10074);
nor U14564 (N_14564,N_6413,N_7415);
or U14565 (N_14565,N_11735,N_6695);
and U14566 (N_14566,N_6092,N_8044);
or U14567 (N_14567,N_7902,N_6311);
or U14568 (N_14568,N_10770,N_8888);
nand U14569 (N_14569,N_10296,N_8265);
nor U14570 (N_14570,N_10090,N_8158);
and U14571 (N_14571,N_8313,N_6920);
nand U14572 (N_14572,N_7564,N_6254);
nor U14573 (N_14573,N_10149,N_10659);
or U14574 (N_14574,N_6318,N_11952);
nand U14575 (N_14575,N_7965,N_11432);
and U14576 (N_14576,N_8995,N_7480);
or U14577 (N_14577,N_10477,N_11105);
xor U14578 (N_14578,N_11619,N_9595);
or U14579 (N_14579,N_8315,N_9170);
xor U14580 (N_14580,N_6188,N_8241);
or U14581 (N_14581,N_9025,N_8441);
nor U14582 (N_14582,N_8405,N_7402);
xnor U14583 (N_14583,N_7640,N_6586);
or U14584 (N_14584,N_10018,N_6189);
and U14585 (N_14585,N_8039,N_10714);
or U14586 (N_14586,N_6463,N_8781);
and U14587 (N_14587,N_7245,N_8648);
nor U14588 (N_14588,N_8361,N_7147);
or U14589 (N_14589,N_8616,N_10075);
nand U14590 (N_14590,N_6247,N_6237);
and U14591 (N_14591,N_9971,N_9503);
nand U14592 (N_14592,N_8726,N_10251);
nand U14593 (N_14593,N_6796,N_10040);
and U14594 (N_14594,N_6538,N_10445);
or U14595 (N_14595,N_11153,N_9075);
or U14596 (N_14596,N_9221,N_7761);
or U14597 (N_14597,N_6882,N_11483);
nand U14598 (N_14598,N_10584,N_7983);
or U14599 (N_14599,N_10739,N_9694);
or U14600 (N_14600,N_6221,N_7565);
nor U14601 (N_14601,N_11971,N_9301);
or U14602 (N_14602,N_7547,N_7173);
and U14603 (N_14603,N_11820,N_9780);
and U14604 (N_14604,N_10791,N_11678);
nand U14605 (N_14605,N_7912,N_11813);
and U14606 (N_14606,N_8551,N_9981);
and U14607 (N_14607,N_6029,N_7635);
or U14608 (N_14608,N_10608,N_11393);
nor U14609 (N_14609,N_11950,N_9514);
nor U14610 (N_14610,N_6134,N_10298);
nor U14611 (N_14611,N_6540,N_7788);
or U14612 (N_14612,N_10790,N_6053);
nor U14613 (N_14613,N_9602,N_6185);
or U14614 (N_14614,N_6058,N_11803);
xnor U14615 (N_14615,N_7206,N_9377);
nand U14616 (N_14616,N_7316,N_8592);
or U14617 (N_14617,N_9356,N_10022);
nor U14618 (N_14618,N_9803,N_11181);
nor U14619 (N_14619,N_8168,N_11589);
nor U14620 (N_14620,N_6403,N_9583);
nand U14621 (N_14621,N_6236,N_6839);
nand U14622 (N_14622,N_10499,N_10365);
nand U14623 (N_14623,N_6065,N_11674);
and U14624 (N_14624,N_11467,N_7712);
and U14625 (N_14625,N_11744,N_7808);
nor U14626 (N_14626,N_11968,N_11513);
nor U14627 (N_14627,N_9380,N_11429);
xor U14628 (N_14628,N_11647,N_9070);
and U14629 (N_14629,N_8922,N_10286);
nor U14630 (N_14630,N_10888,N_7451);
and U14631 (N_14631,N_9500,N_11441);
or U14632 (N_14632,N_6033,N_7047);
and U14633 (N_14633,N_11939,N_7853);
and U14634 (N_14634,N_8821,N_11726);
nor U14635 (N_14635,N_7935,N_6131);
or U14636 (N_14636,N_7909,N_8915);
nand U14637 (N_14637,N_11320,N_8949);
nor U14638 (N_14638,N_8222,N_7463);
nor U14639 (N_14639,N_9968,N_7938);
nand U14640 (N_14640,N_7740,N_6416);
nor U14641 (N_14641,N_8584,N_9298);
and U14642 (N_14642,N_7691,N_8877);
or U14643 (N_14643,N_10772,N_6710);
nand U14644 (N_14644,N_9627,N_10357);
nand U14645 (N_14645,N_11718,N_9782);
or U14646 (N_14646,N_8511,N_9783);
nand U14647 (N_14647,N_11146,N_6400);
xnor U14648 (N_14648,N_10218,N_10552);
and U14649 (N_14649,N_6255,N_10126);
nor U14650 (N_14650,N_11990,N_8449);
nand U14651 (N_14651,N_6164,N_9657);
and U14652 (N_14652,N_11923,N_7322);
and U14653 (N_14653,N_8808,N_7075);
and U14654 (N_14654,N_9767,N_9698);
or U14655 (N_14655,N_8292,N_8147);
nand U14656 (N_14656,N_11512,N_11377);
nor U14657 (N_14657,N_11398,N_7762);
or U14658 (N_14658,N_11816,N_7840);
or U14659 (N_14659,N_8928,N_7621);
and U14660 (N_14660,N_6543,N_8933);
and U14661 (N_14661,N_8987,N_9772);
nand U14662 (N_14662,N_11263,N_11041);
nor U14663 (N_14663,N_7876,N_8849);
xor U14664 (N_14664,N_8536,N_7427);
nor U14665 (N_14665,N_6717,N_10504);
nor U14666 (N_14666,N_6244,N_8859);
or U14667 (N_14667,N_6603,N_9090);
nor U14668 (N_14668,N_9235,N_11850);
nor U14669 (N_14669,N_6568,N_6480);
and U14670 (N_14670,N_7022,N_10591);
nand U14671 (N_14671,N_10360,N_11052);
and U14672 (N_14672,N_6302,N_6686);
nand U14673 (N_14673,N_7105,N_11498);
and U14674 (N_14674,N_9956,N_11054);
nor U14675 (N_14675,N_10904,N_11099);
or U14676 (N_14676,N_10284,N_8075);
or U14677 (N_14677,N_10320,N_6625);
nor U14678 (N_14678,N_9432,N_11156);
or U14679 (N_14679,N_11370,N_8930);
and U14680 (N_14680,N_7267,N_7250);
nand U14681 (N_14681,N_7951,N_9616);
and U14682 (N_14682,N_8266,N_7908);
xnor U14683 (N_14683,N_7229,N_9539);
and U14684 (N_14684,N_6623,N_8715);
and U14685 (N_14685,N_11204,N_9452);
xnor U14686 (N_14686,N_9926,N_10450);
nor U14687 (N_14687,N_6038,N_6260);
and U14688 (N_14688,N_8574,N_11703);
and U14689 (N_14689,N_10767,N_11777);
nor U14690 (N_14690,N_9226,N_8256);
or U14691 (N_14691,N_11821,N_10035);
nand U14692 (N_14692,N_11909,N_7936);
nor U14693 (N_14693,N_10648,N_7979);
and U14694 (N_14694,N_6006,N_10354);
and U14695 (N_14695,N_10355,N_7934);
xor U14696 (N_14696,N_7626,N_8008);
nand U14697 (N_14697,N_7715,N_9484);
xnor U14698 (N_14698,N_7181,N_10194);
and U14699 (N_14699,N_7805,N_8891);
and U14700 (N_14700,N_9169,N_8051);
xnor U14701 (N_14701,N_9561,N_9388);
nor U14702 (N_14702,N_10775,N_10057);
xor U14703 (N_14703,N_7237,N_6880);
and U14704 (N_14704,N_6218,N_10873);
or U14705 (N_14705,N_6739,N_6424);
nor U14706 (N_14706,N_9429,N_10782);
nand U14707 (N_14707,N_6220,N_6273);
or U14708 (N_14708,N_8298,N_8601);
and U14709 (N_14709,N_6197,N_11763);
nor U14710 (N_14710,N_6970,N_6081);
nor U14711 (N_14711,N_9030,N_8841);
and U14712 (N_14712,N_11163,N_7648);
nand U14713 (N_14713,N_7301,N_11865);
or U14714 (N_14714,N_7141,N_8604);
nor U14715 (N_14715,N_10671,N_9140);
and U14716 (N_14716,N_6074,N_8637);
nor U14717 (N_14717,N_10863,N_7744);
xor U14718 (N_14718,N_9210,N_8847);
xor U14719 (N_14719,N_7751,N_7483);
and U14720 (N_14720,N_6937,N_9648);
nor U14721 (N_14721,N_7624,N_11279);
or U14722 (N_14722,N_10774,N_7238);
nor U14723 (N_14723,N_10051,N_9251);
nor U14724 (N_14724,N_11942,N_10623);
and U14725 (N_14725,N_8122,N_10228);
and U14726 (N_14726,N_9584,N_10312);
nor U14727 (N_14727,N_9401,N_11883);
and U14728 (N_14728,N_9587,N_7220);
or U14729 (N_14729,N_8082,N_9609);
nand U14730 (N_14730,N_11308,N_7543);
nand U14731 (N_14731,N_9955,N_10494);
nand U14732 (N_14732,N_10014,N_11322);
nor U14733 (N_14733,N_10421,N_9943);
nand U14734 (N_14734,N_8524,N_7779);
and U14735 (N_14735,N_8105,N_8382);
xor U14736 (N_14736,N_6904,N_6477);
nor U14737 (N_14737,N_11542,N_8992);
nand U14738 (N_14738,N_11446,N_7950);
xor U14739 (N_14739,N_9201,N_10598);
or U14740 (N_14740,N_6676,N_11867);
nor U14741 (N_14741,N_11837,N_7481);
nand U14742 (N_14742,N_8475,N_7286);
nor U14743 (N_14743,N_10304,N_8548);
nor U14744 (N_14744,N_10239,N_9035);
nor U14745 (N_14745,N_11271,N_11600);
and U14746 (N_14746,N_9841,N_11992);
and U14747 (N_14747,N_11391,N_6445);
nand U14748 (N_14748,N_7862,N_7608);
nor U14749 (N_14749,N_7680,N_7274);
or U14750 (N_14750,N_11477,N_10866);
nand U14751 (N_14751,N_8671,N_7034);
nor U14752 (N_14752,N_6953,N_11632);
nand U14753 (N_14753,N_8605,N_11385);
or U14754 (N_14754,N_6892,N_11704);
nand U14755 (N_14755,N_9010,N_9540);
and U14756 (N_14756,N_11504,N_8645);
nand U14757 (N_14757,N_6958,N_10037);
nand U14758 (N_14758,N_8060,N_7216);
or U14759 (N_14759,N_8028,N_10695);
nor U14760 (N_14760,N_10291,N_11855);
nand U14761 (N_14761,N_9504,N_6506);
nor U14762 (N_14762,N_6525,N_8104);
or U14763 (N_14763,N_7314,N_8130);
nor U14764 (N_14764,N_8621,N_7104);
xnor U14765 (N_14765,N_11372,N_11806);
nand U14766 (N_14766,N_6601,N_6447);
or U14767 (N_14767,N_9766,N_10486);
xnor U14768 (N_14768,N_11282,N_6589);
nor U14769 (N_14769,N_8174,N_10329);
or U14770 (N_14770,N_9860,N_7957);
and U14771 (N_14771,N_9641,N_10240);
nor U14772 (N_14772,N_11409,N_11927);
or U14773 (N_14773,N_6961,N_10539);
nor U14774 (N_14774,N_9188,N_10937);
or U14775 (N_14775,N_6949,N_9082);
and U14776 (N_14776,N_11346,N_6338);
nor U14777 (N_14777,N_10015,N_9284);
nor U14778 (N_14778,N_7117,N_10099);
nor U14779 (N_14779,N_10107,N_6468);
or U14780 (N_14780,N_11257,N_8022);
and U14781 (N_14781,N_8341,N_10717);
nand U14782 (N_14782,N_8485,N_6570);
and U14783 (N_14783,N_8165,N_7209);
and U14784 (N_14784,N_8200,N_6789);
nand U14785 (N_14785,N_7886,N_11415);
nand U14786 (N_14786,N_8561,N_10850);
or U14787 (N_14787,N_7851,N_10855);
or U14788 (N_14788,N_9046,N_8880);
nand U14789 (N_14789,N_8921,N_9496);
and U14790 (N_14790,N_6336,N_11419);
and U14791 (N_14791,N_9002,N_11550);
or U14792 (N_14792,N_11967,N_7889);
nand U14793 (N_14793,N_8351,N_8876);
and U14794 (N_14794,N_10821,N_10654);
nand U14795 (N_14795,N_8835,N_8924);
nor U14796 (N_14796,N_9148,N_8644);
nor U14797 (N_14797,N_11700,N_9307);
and U14798 (N_14798,N_7131,N_7738);
or U14799 (N_14799,N_7706,N_11291);
nor U14800 (N_14800,N_8455,N_9982);
nand U14801 (N_14801,N_9364,N_10532);
or U14802 (N_14802,N_11174,N_9024);
and U14803 (N_14803,N_9236,N_7831);
nor U14804 (N_14804,N_11613,N_8858);
xnor U14805 (N_14805,N_8095,N_6353);
nand U14806 (N_14806,N_11205,N_7823);
xnor U14807 (N_14807,N_7330,N_6938);
xor U14808 (N_14808,N_9613,N_8296);
and U14809 (N_14809,N_7069,N_7900);
and U14810 (N_14810,N_11544,N_11982);
or U14811 (N_14811,N_10392,N_10773);
nor U14812 (N_14812,N_11048,N_9390);
and U14813 (N_14813,N_10443,N_10548);
nand U14814 (N_14814,N_9820,N_8297);
or U14815 (N_14815,N_9213,N_11034);
and U14816 (N_14816,N_10530,N_11617);
nand U14817 (N_14817,N_6425,N_9960);
or U14818 (N_14818,N_10432,N_8460);
and U14819 (N_14819,N_6219,N_8059);
nor U14820 (N_14820,N_11148,N_6394);
nand U14821 (N_14821,N_6036,N_11310);
or U14822 (N_14822,N_6607,N_6308);
and U14823 (N_14823,N_11598,N_7599);
and U14824 (N_14824,N_11192,N_11630);
or U14825 (N_14825,N_8760,N_7376);
nand U14826 (N_14826,N_10166,N_11091);
nand U14827 (N_14827,N_11293,N_10427);
nor U14828 (N_14828,N_10582,N_10106);
or U14829 (N_14829,N_7183,N_9909);
xor U14830 (N_14830,N_7657,N_7874);
nor U14831 (N_14831,N_10506,N_11857);
nand U14832 (N_14832,N_11388,N_10278);
or U14833 (N_14833,N_6895,N_6602);
nand U14834 (N_14834,N_6386,N_9855);
or U14835 (N_14835,N_8205,N_6886);
or U14836 (N_14836,N_9704,N_10845);
nor U14837 (N_14837,N_9856,N_6475);
or U14838 (N_14838,N_6928,N_7555);
nand U14839 (N_14839,N_8444,N_11634);
nand U14840 (N_14840,N_6205,N_9755);
and U14841 (N_14841,N_9045,N_11928);
nor U14842 (N_14842,N_6745,N_9932);
and U14843 (N_14843,N_11792,N_11396);
and U14844 (N_14844,N_9888,N_9749);
or U14845 (N_14845,N_11355,N_6368);
nand U14846 (N_14846,N_6648,N_10853);
or U14847 (N_14847,N_8355,N_9486);
nor U14848 (N_14848,N_8391,N_6199);
nand U14849 (N_14849,N_11709,N_8971);
or U14850 (N_14850,N_11092,N_11847);
or U14851 (N_14851,N_7113,N_10134);
nor U14852 (N_14852,N_10797,N_10825);
and U14853 (N_14853,N_6533,N_11162);
and U14854 (N_14854,N_9873,N_8396);
nand U14855 (N_14855,N_6925,N_9379);
and U14856 (N_14856,N_11789,N_7814);
xor U14857 (N_14857,N_6762,N_10175);
nor U14858 (N_14858,N_6718,N_6402);
nor U14859 (N_14859,N_10963,N_10657);
and U14860 (N_14860,N_6060,N_10381);
nor U14861 (N_14861,N_6233,N_9259);
or U14862 (N_14862,N_6397,N_10578);
or U14863 (N_14863,N_8048,N_10127);
nand U14864 (N_14864,N_10306,N_6508);
xnor U14865 (N_14865,N_8942,N_11352);
or U14866 (N_14866,N_9642,N_9359);
or U14867 (N_14867,N_8263,N_6902);
nor U14868 (N_14868,N_7074,N_6362);
and U14869 (N_14869,N_11499,N_10926);
nor U14870 (N_14870,N_9326,N_7384);
nand U14871 (N_14871,N_7931,N_10220);
or U14872 (N_14872,N_6151,N_7452);
nand U14873 (N_14873,N_8994,N_10395);
nor U14874 (N_14874,N_7002,N_10176);
nor U14875 (N_14875,N_8261,N_7111);
or U14876 (N_14876,N_9399,N_9936);
xor U14877 (N_14877,N_8272,N_8290);
nor U14878 (N_14878,N_11846,N_9507);
nor U14879 (N_14879,N_6371,N_6315);
or U14880 (N_14880,N_9096,N_8553);
or U14881 (N_14881,N_8488,N_10252);
nor U14882 (N_14882,N_8163,N_11235);
nand U14883 (N_14883,N_11407,N_11224);
nand U14884 (N_14884,N_6605,N_7868);
nand U14885 (N_14885,N_9975,N_6224);
and U14886 (N_14886,N_8749,N_9753);
or U14887 (N_14887,N_6946,N_6921);
nor U14888 (N_14888,N_9027,N_10429);
nand U14889 (N_14889,N_7370,N_9615);
and U14890 (N_14890,N_10232,N_8904);
and U14891 (N_14891,N_9623,N_7756);
or U14892 (N_14892,N_10673,N_11859);
nor U14893 (N_14893,N_11815,N_9827);
or U14894 (N_14894,N_6230,N_7569);
nor U14895 (N_14895,N_10991,N_7727);
xnor U14896 (N_14896,N_6229,N_7482);
nand U14897 (N_14897,N_10029,N_8107);
nand U14898 (N_14898,N_9597,N_11464);
and U14899 (N_14899,N_11079,N_7638);
nor U14900 (N_14900,N_8932,N_7632);
xor U14901 (N_14901,N_11301,N_7913);
nand U14902 (N_14902,N_9696,N_7688);
and U14903 (N_14903,N_10397,N_6757);
nor U14904 (N_14904,N_11563,N_7644);
or U14905 (N_14905,N_10940,N_6531);
nor U14906 (N_14906,N_7018,N_8445);
nand U14907 (N_14907,N_11802,N_9789);
nand U14908 (N_14908,N_6521,N_11083);
nand U14909 (N_14909,N_7139,N_7064);
xnor U14910 (N_14910,N_7129,N_7813);
and U14911 (N_14911,N_10510,N_10666);
and U14912 (N_14912,N_8207,N_7716);
or U14913 (N_14913,N_7850,N_8244);
nor U14914 (N_14914,N_7820,N_11440);
nand U14915 (N_14915,N_7177,N_9407);
nand U14916 (N_14916,N_9785,N_8746);
or U14917 (N_14917,N_10133,N_6108);
nor U14918 (N_14918,N_6040,N_10785);
nor U14919 (N_14919,N_11799,N_10805);
nor U14920 (N_14920,N_9620,N_7753);
nand U14921 (N_14921,N_9165,N_6329);
nor U14922 (N_14922,N_7438,N_6552);
and U14923 (N_14923,N_7474,N_7980);
nand U14924 (N_14924,N_9738,N_9376);
xor U14925 (N_14925,N_8963,N_9837);
or U14926 (N_14926,N_11756,N_7065);
nor U14927 (N_14927,N_7581,N_6801);
and U14928 (N_14928,N_8755,N_10344);
nand U14929 (N_14929,N_10132,N_6727);
nor U14930 (N_14930,N_6537,N_10437);
and U14931 (N_14931,N_7701,N_9672);
and U14932 (N_14932,N_7255,N_11590);
nand U14933 (N_14933,N_11500,N_9684);
xor U14934 (N_14934,N_7841,N_6615);
nand U14935 (N_14935,N_9415,N_9994);
nand U14936 (N_14936,N_9204,N_11892);
nand U14937 (N_14937,N_8258,N_11864);
or U14938 (N_14938,N_11594,N_8659);
and U14939 (N_14939,N_10442,N_10476);
nand U14940 (N_14940,N_7893,N_10535);
nand U14941 (N_14941,N_9119,N_10052);
and U14942 (N_14942,N_8465,N_7866);
nand U14943 (N_14943,N_11900,N_10931);
nor U14944 (N_14944,N_6822,N_9400);
nor U14945 (N_14945,N_11599,N_9152);
or U14946 (N_14946,N_10319,N_9652);
or U14947 (N_14947,N_7031,N_10181);
or U14948 (N_14948,N_7256,N_8395);
or U14949 (N_14949,N_8564,N_6350);
nand U14950 (N_14950,N_11035,N_10965);
nand U14951 (N_14951,N_7318,N_6672);
nor U14952 (N_14952,N_9622,N_9907);
nor U14953 (N_14953,N_8506,N_8588);
or U14954 (N_14954,N_10571,N_6037);
nand U14955 (N_14955,N_6209,N_9666);
xnor U14956 (N_14956,N_8101,N_7826);
or U14957 (N_14957,N_8532,N_10624);
nor U14958 (N_14958,N_10793,N_11225);
nand U14959 (N_14959,N_7409,N_10213);
or U14960 (N_14960,N_8667,N_10956);
nand U14961 (N_14961,N_10211,N_8185);
nor U14962 (N_14962,N_6912,N_11584);
xnor U14963 (N_14963,N_11987,N_11186);
or U14964 (N_14964,N_9653,N_6755);
nand U14965 (N_14965,N_8394,N_9292);
nand U14966 (N_14966,N_6752,N_8565);
or U14967 (N_14967,N_8918,N_6319);
nand U14968 (N_14968,N_11071,N_6382);
xnor U14969 (N_14969,N_10833,N_6557);
or U14970 (N_14970,N_11126,N_9488);
nor U14971 (N_14971,N_10073,N_10660);
or U14972 (N_14972,N_9385,N_7353);
nor U14973 (N_14973,N_6781,N_9038);
nor U14974 (N_14974,N_8325,N_8041);
or U14975 (N_14975,N_8450,N_9636);
xor U14976 (N_14976,N_6103,N_7746);
and U14977 (N_14977,N_11875,N_7221);
or U14978 (N_14978,N_8332,N_9697);
nor U14979 (N_14979,N_9529,N_7395);
nor U14980 (N_14980,N_9533,N_7969);
nor U14981 (N_14981,N_9959,N_9740);
or U14982 (N_14982,N_11284,N_10272);
xor U14983 (N_14983,N_11075,N_9476);
xor U14984 (N_14984,N_9513,N_9275);
and U14985 (N_14985,N_6242,N_6096);
nor U14986 (N_14986,N_11025,N_9240);
or U14987 (N_14987,N_6322,N_8993);
or U14988 (N_14988,N_11453,N_8991);
and U14989 (N_14989,N_8368,N_11302);
nor U14990 (N_14990,N_6401,N_11757);
and U14991 (N_14991,N_6840,N_9631);
and U14992 (N_14992,N_10612,N_9714);
or U14993 (N_14993,N_9473,N_7212);
and U14994 (N_14994,N_8273,N_11758);
nand U14995 (N_14995,N_10337,N_10280);
and U14996 (N_14996,N_6889,N_8144);
nand U14997 (N_14997,N_11437,N_8619);
or U14998 (N_14998,N_7616,N_7655);
nand U14999 (N_14999,N_11093,N_10575);
nor U15000 (N_15000,N_11010,N_6503);
nand U15001 (N_15001,N_9480,N_10935);
or U15002 (N_15002,N_10151,N_9481);
xnor U15003 (N_15003,N_7133,N_6886);
nor U15004 (N_15004,N_6145,N_6911);
and U15005 (N_15005,N_9882,N_6917);
and U15006 (N_15006,N_9047,N_9945);
and U15007 (N_15007,N_6682,N_9640);
nor U15008 (N_15008,N_8409,N_6230);
and U15009 (N_15009,N_6991,N_6306);
and U15010 (N_15010,N_8356,N_7945);
nand U15011 (N_15011,N_7484,N_7213);
and U15012 (N_15012,N_7862,N_9545);
nor U15013 (N_15013,N_9838,N_7157);
and U15014 (N_15014,N_10221,N_7292);
and U15015 (N_15015,N_11919,N_8513);
nand U15016 (N_15016,N_9050,N_11432);
nand U15017 (N_15017,N_10835,N_7828);
nor U15018 (N_15018,N_9229,N_9717);
nor U15019 (N_15019,N_11712,N_9492);
xnor U15020 (N_15020,N_7868,N_8364);
and U15021 (N_15021,N_6346,N_8586);
nor U15022 (N_15022,N_7453,N_10120);
and U15023 (N_15023,N_9743,N_7289);
nor U15024 (N_15024,N_11540,N_6767);
and U15025 (N_15025,N_7362,N_8312);
xnor U15026 (N_15026,N_9923,N_6765);
nand U15027 (N_15027,N_6047,N_11980);
nand U15028 (N_15028,N_8882,N_10392);
and U15029 (N_15029,N_6385,N_6701);
xor U15030 (N_15030,N_6359,N_10206);
or U15031 (N_15031,N_9707,N_9329);
xor U15032 (N_15032,N_6014,N_9793);
nand U15033 (N_15033,N_8362,N_6744);
nor U15034 (N_15034,N_6247,N_11271);
or U15035 (N_15035,N_8757,N_11226);
nor U15036 (N_15036,N_7555,N_10849);
nor U15037 (N_15037,N_7613,N_7373);
xor U15038 (N_15038,N_11946,N_11175);
xnor U15039 (N_15039,N_7191,N_10448);
nand U15040 (N_15040,N_7338,N_11219);
xor U15041 (N_15041,N_7678,N_6327);
nand U15042 (N_15042,N_7771,N_10447);
nor U15043 (N_15043,N_11010,N_11005);
nor U15044 (N_15044,N_10067,N_11940);
xor U15045 (N_15045,N_8260,N_11614);
nor U15046 (N_15046,N_6848,N_6086);
nand U15047 (N_15047,N_7631,N_8800);
nand U15048 (N_15048,N_9603,N_6804);
or U15049 (N_15049,N_11448,N_11937);
and U15050 (N_15050,N_9675,N_6489);
or U15051 (N_15051,N_6464,N_7907);
and U15052 (N_15052,N_8685,N_10023);
nand U15053 (N_15053,N_9262,N_9878);
nor U15054 (N_15054,N_6517,N_6493);
nor U15055 (N_15055,N_7823,N_10078);
or U15056 (N_15056,N_9844,N_7307);
nand U15057 (N_15057,N_8569,N_10366);
and U15058 (N_15058,N_7010,N_9819);
nand U15059 (N_15059,N_9105,N_11649);
and U15060 (N_15060,N_10262,N_11839);
or U15061 (N_15061,N_6460,N_6575);
and U15062 (N_15062,N_10449,N_11105);
nor U15063 (N_15063,N_11025,N_10803);
nor U15064 (N_15064,N_6154,N_11245);
nand U15065 (N_15065,N_8362,N_7838);
and U15066 (N_15066,N_11696,N_10389);
xor U15067 (N_15067,N_7067,N_6182);
nand U15068 (N_15068,N_9196,N_8522);
or U15069 (N_15069,N_7601,N_10914);
or U15070 (N_15070,N_9743,N_11316);
nand U15071 (N_15071,N_7253,N_6603);
nand U15072 (N_15072,N_7606,N_8100);
or U15073 (N_15073,N_9323,N_10863);
nand U15074 (N_15074,N_10403,N_6675);
xnor U15075 (N_15075,N_10650,N_11900);
or U15076 (N_15076,N_8700,N_9956);
nor U15077 (N_15077,N_11392,N_11106);
and U15078 (N_15078,N_8505,N_7083);
nor U15079 (N_15079,N_7190,N_11284);
xnor U15080 (N_15080,N_8124,N_10391);
xor U15081 (N_15081,N_11908,N_11384);
xnor U15082 (N_15082,N_9454,N_8955);
and U15083 (N_15083,N_11172,N_7532);
and U15084 (N_15084,N_7798,N_11809);
and U15085 (N_15085,N_8193,N_6941);
and U15086 (N_15086,N_9645,N_9464);
or U15087 (N_15087,N_8596,N_6954);
xnor U15088 (N_15088,N_7657,N_11554);
nand U15089 (N_15089,N_9550,N_10607);
or U15090 (N_15090,N_8780,N_7379);
nor U15091 (N_15091,N_6191,N_8739);
nand U15092 (N_15092,N_9613,N_11026);
nor U15093 (N_15093,N_10163,N_6529);
and U15094 (N_15094,N_9617,N_10484);
or U15095 (N_15095,N_11601,N_7960);
nand U15096 (N_15096,N_8973,N_7126);
xor U15097 (N_15097,N_8766,N_10623);
nand U15098 (N_15098,N_10117,N_7619);
nor U15099 (N_15099,N_9906,N_11176);
nand U15100 (N_15100,N_6644,N_8022);
or U15101 (N_15101,N_9164,N_11964);
nor U15102 (N_15102,N_8820,N_11941);
and U15103 (N_15103,N_10503,N_6067);
and U15104 (N_15104,N_9628,N_6396);
nand U15105 (N_15105,N_11789,N_11091);
or U15106 (N_15106,N_11195,N_9584);
nand U15107 (N_15107,N_9419,N_6550);
or U15108 (N_15108,N_11263,N_8316);
or U15109 (N_15109,N_11631,N_7554);
nor U15110 (N_15110,N_9173,N_6923);
nand U15111 (N_15111,N_9466,N_10618);
nor U15112 (N_15112,N_7811,N_7193);
and U15113 (N_15113,N_11348,N_10437);
and U15114 (N_15114,N_7034,N_11750);
and U15115 (N_15115,N_7185,N_7163);
nor U15116 (N_15116,N_10633,N_8034);
or U15117 (N_15117,N_10938,N_7825);
nand U15118 (N_15118,N_11179,N_7491);
or U15119 (N_15119,N_7063,N_9329);
nand U15120 (N_15120,N_7321,N_7749);
or U15121 (N_15121,N_11329,N_11463);
nand U15122 (N_15122,N_6459,N_10428);
xnor U15123 (N_15123,N_11386,N_11931);
xor U15124 (N_15124,N_7985,N_6640);
or U15125 (N_15125,N_8902,N_11329);
nand U15126 (N_15126,N_8989,N_9297);
nand U15127 (N_15127,N_9144,N_11524);
or U15128 (N_15128,N_10546,N_8389);
nor U15129 (N_15129,N_9111,N_7077);
nor U15130 (N_15130,N_8183,N_8181);
nor U15131 (N_15131,N_6468,N_8891);
nand U15132 (N_15132,N_9680,N_11275);
and U15133 (N_15133,N_9740,N_9519);
and U15134 (N_15134,N_10121,N_11339);
and U15135 (N_15135,N_10883,N_9178);
nor U15136 (N_15136,N_9569,N_6555);
and U15137 (N_15137,N_10579,N_9282);
nor U15138 (N_15138,N_8501,N_11708);
nor U15139 (N_15139,N_8578,N_11805);
nand U15140 (N_15140,N_6600,N_9956);
and U15141 (N_15141,N_7673,N_11071);
and U15142 (N_15142,N_7606,N_9091);
nor U15143 (N_15143,N_7329,N_9107);
nor U15144 (N_15144,N_6550,N_9451);
and U15145 (N_15145,N_8968,N_6091);
or U15146 (N_15146,N_10168,N_8924);
or U15147 (N_15147,N_10679,N_11955);
or U15148 (N_15148,N_11095,N_7153);
or U15149 (N_15149,N_9978,N_9778);
nand U15150 (N_15150,N_9986,N_6127);
xor U15151 (N_15151,N_8364,N_10220);
nor U15152 (N_15152,N_9614,N_6870);
nor U15153 (N_15153,N_8693,N_8274);
or U15154 (N_15154,N_10117,N_8100);
nor U15155 (N_15155,N_11836,N_9346);
nor U15156 (N_15156,N_11807,N_9498);
or U15157 (N_15157,N_9699,N_7655);
nor U15158 (N_15158,N_7312,N_11737);
or U15159 (N_15159,N_8478,N_6653);
and U15160 (N_15160,N_11743,N_8110);
nor U15161 (N_15161,N_10898,N_9728);
or U15162 (N_15162,N_10462,N_8143);
nand U15163 (N_15163,N_11787,N_11663);
or U15164 (N_15164,N_8746,N_8353);
nand U15165 (N_15165,N_6926,N_6010);
or U15166 (N_15166,N_7681,N_6353);
nand U15167 (N_15167,N_9655,N_6765);
and U15168 (N_15168,N_7471,N_8712);
nand U15169 (N_15169,N_9650,N_11057);
nor U15170 (N_15170,N_11145,N_6918);
nand U15171 (N_15171,N_11275,N_7393);
and U15172 (N_15172,N_8021,N_6385);
or U15173 (N_15173,N_7173,N_9215);
nor U15174 (N_15174,N_8709,N_11189);
and U15175 (N_15175,N_11640,N_9738);
xor U15176 (N_15176,N_10274,N_6967);
nor U15177 (N_15177,N_8026,N_10520);
nand U15178 (N_15178,N_8660,N_10142);
xor U15179 (N_15179,N_7663,N_9734);
nor U15180 (N_15180,N_9122,N_10169);
and U15181 (N_15181,N_8520,N_7694);
nor U15182 (N_15182,N_6242,N_7547);
or U15183 (N_15183,N_11105,N_6468);
and U15184 (N_15184,N_7671,N_10607);
and U15185 (N_15185,N_10264,N_8164);
xor U15186 (N_15186,N_11781,N_9298);
nand U15187 (N_15187,N_10685,N_11350);
and U15188 (N_15188,N_9412,N_10959);
or U15189 (N_15189,N_10706,N_8015);
nand U15190 (N_15190,N_10150,N_9302);
nand U15191 (N_15191,N_9753,N_8644);
and U15192 (N_15192,N_9971,N_6940);
nor U15193 (N_15193,N_11700,N_10824);
or U15194 (N_15194,N_6114,N_10452);
and U15195 (N_15195,N_10785,N_10645);
or U15196 (N_15196,N_11540,N_6460);
xnor U15197 (N_15197,N_9852,N_10664);
nor U15198 (N_15198,N_9383,N_9899);
or U15199 (N_15199,N_6295,N_9571);
nor U15200 (N_15200,N_9910,N_8767);
and U15201 (N_15201,N_8245,N_6434);
nand U15202 (N_15202,N_8104,N_8253);
nor U15203 (N_15203,N_8954,N_8446);
and U15204 (N_15204,N_11808,N_8226);
nor U15205 (N_15205,N_6090,N_6210);
nor U15206 (N_15206,N_9292,N_8938);
and U15207 (N_15207,N_7291,N_10365);
nor U15208 (N_15208,N_9836,N_8117);
xor U15209 (N_15209,N_7871,N_8497);
xor U15210 (N_15210,N_9739,N_11122);
nand U15211 (N_15211,N_8701,N_7398);
or U15212 (N_15212,N_8550,N_11395);
and U15213 (N_15213,N_8308,N_9781);
nand U15214 (N_15214,N_11173,N_9453);
and U15215 (N_15215,N_10342,N_8925);
nand U15216 (N_15216,N_10729,N_6630);
or U15217 (N_15217,N_7893,N_7577);
and U15218 (N_15218,N_9188,N_10960);
and U15219 (N_15219,N_6189,N_9985);
nand U15220 (N_15220,N_9932,N_10632);
nand U15221 (N_15221,N_6643,N_11796);
nand U15222 (N_15222,N_9088,N_6805);
nor U15223 (N_15223,N_9632,N_6856);
or U15224 (N_15224,N_8090,N_11098);
and U15225 (N_15225,N_10642,N_10315);
nand U15226 (N_15226,N_6408,N_9519);
or U15227 (N_15227,N_8921,N_6823);
and U15228 (N_15228,N_8711,N_9158);
nand U15229 (N_15229,N_11748,N_10387);
and U15230 (N_15230,N_10040,N_6524);
nand U15231 (N_15231,N_6830,N_6423);
or U15232 (N_15232,N_10597,N_11401);
nand U15233 (N_15233,N_11848,N_7682);
nor U15234 (N_15234,N_9997,N_11444);
nor U15235 (N_15235,N_8168,N_6397);
and U15236 (N_15236,N_6971,N_6431);
nand U15237 (N_15237,N_6292,N_11806);
or U15238 (N_15238,N_8362,N_9771);
nor U15239 (N_15239,N_8001,N_11068);
nor U15240 (N_15240,N_11472,N_9736);
or U15241 (N_15241,N_7415,N_6714);
nor U15242 (N_15242,N_11190,N_8995);
xnor U15243 (N_15243,N_8989,N_6332);
or U15244 (N_15244,N_8180,N_8616);
or U15245 (N_15245,N_8929,N_7619);
xnor U15246 (N_15246,N_10383,N_7394);
xor U15247 (N_15247,N_9235,N_11201);
nor U15248 (N_15248,N_11215,N_9569);
or U15249 (N_15249,N_6291,N_9273);
and U15250 (N_15250,N_6723,N_9322);
or U15251 (N_15251,N_9453,N_8964);
or U15252 (N_15252,N_7374,N_11572);
xor U15253 (N_15253,N_9362,N_9506);
or U15254 (N_15254,N_9895,N_7870);
nand U15255 (N_15255,N_6497,N_10620);
or U15256 (N_15256,N_7903,N_6044);
and U15257 (N_15257,N_9336,N_10967);
xor U15258 (N_15258,N_6631,N_8279);
nand U15259 (N_15259,N_9165,N_9338);
or U15260 (N_15260,N_8919,N_11405);
and U15261 (N_15261,N_11447,N_10801);
nand U15262 (N_15262,N_10735,N_6553);
or U15263 (N_15263,N_6783,N_8373);
nand U15264 (N_15264,N_6804,N_10554);
xnor U15265 (N_15265,N_6546,N_10755);
nor U15266 (N_15266,N_10254,N_9351);
and U15267 (N_15267,N_8713,N_8699);
xnor U15268 (N_15268,N_6116,N_11778);
and U15269 (N_15269,N_11532,N_7215);
nor U15270 (N_15270,N_11778,N_6987);
nor U15271 (N_15271,N_9821,N_10623);
nor U15272 (N_15272,N_10270,N_10527);
nand U15273 (N_15273,N_10359,N_11165);
xor U15274 (N_15274,N_11485,N_6042);
nand U15275 (N_15275,N_7928,N_8399);
and U15276 (N_15276,N_9140,N_7264);
or U15277 (N_15277,N_11517,N_8560);
and U15278 (N_15278,N_11406,N_6807);
or U15279 (N_15279,N_7604,N_11321);
nor U15280 (N_15280,N_6144,N_10210);
nor U15281 (N_15281,N_7244,N_8791);
and U15282 (N_15282,N_9642,N_10051);
and U15283 (N_15283,N_7066,N_7902);
nand U15284 (N_15284,N_6152,N_11243);
or U15285 (N_15285,N_9870,N_10325);
and U15286 (N_15286,N_9189,N_9875);
or U15287 (N_15287,N_9221,N_6880);
and U15288 (N_15288,N_6984,N_7421);
nor U15289 (N_15289,N_7933,N_6920);
or U15290 (N_15290,N_10467,N_9468);
nor U15291 (N_15291,N_9837,N_10939);
and U15292 (N_15292,N_8621,N_10970);
nand U15293 (N_15293,N_11602,N_7820);
nor U15294 (N_15294,N_9210,N_9014);
nand U15295 (N_15295,N_9696,N_7950);
xor U15296 (N_15296,N_10685,N_10300);
or U15297 (N_15297,N_8141,N_11285);
nand U15298 (N_15298,N_9123,N_6041);
or U15299 (N_15299,N_8905,N_9366);
or U15300 (N_15300,N_10380,N_6526);
xnor U15301 (N_15301,N_10304,N_6499);
nor U15302 (N_15302,N_6374,N_10117);
and U15303 (N_15303,N_6651,N_6129);
xnor U15304 (N_15304,N_6231,N_11054);
or U15305 (N_15305,N_11952,N_8388);
and U15306 (N_15306,N_8273,N_11425);
and U15307 (N_15307,N_6471,N_7518);
and U15308 (N_15308,N_9312,N_10921);
nand U15309 (N_15309,N_8855,N_10619);
and U15310 (N_15310,N_8569,N_10920);
and U15311 (N_15311,N_8619,N_10932);
and U15312 (N_15312,N_8298,N_9295);
or U15313 (N_15313,N_10616,N_8090);
nand U15314 (N_15314,N_6842,N_11415);
and U15315 (N_15315,N_11431,N_6999);
and U15316 (N_15316,N_9577,N_9235);
and U15317 (N_15317,N_9772,N_9037);
or U15318 (N_15318,N_8589,N_10444);
nor U15319 (N_15319,N_9033,N_9566);
nand U15320 (N_15320,N_6154,N_11834);
and U15321 (N_15321,N_11597,N_10846);
or U15322 (N_15322,N_8987,N_11891);
nor U15323 (N_15323,N_8811,N_9269);
nor U15324 (N_15324,N_8127,N_11999);
or U15325 (N_15325,N_7778,N_9741);
nand U15326 (N_15326,N_11447,N_6893);
or U15327 (N_15327,N_6567,N_6179);
and U15328 (N_15328,N_11048,N_6275);
and U15329 (N_15329,N_7987,N_8538);
xor U15330 (N_15330,N_7079,N_7944);
and U15331 (N_15331,N_7842,N_10711);
or U15332 (N_15332,N_9468,N_6806);
and U15333 (N_15333,N_8132,N_7365);
nor U15334 (N_15334,N_10958,N_8955);
or U15335 (N_15335,N_7796,N_8080);
or U15336 (N_15336,N_8139,N_7628);
nor U15337 (N_15337,N_9163,N_9002);
or U15338 (N_15338,N_6767,N_10310);
or U15339 (N_15339,N_10122,N_6513);
or U15340 (N_15340,N_7011,N_10315);
or U15341 (N_15341,N_8092,N_9965);
and U15342 (N_15342,N_8008,N_7064);
and U15343 (N_15343,N_10042,N_6553);
and U15344 (N_15344,N_10688,N_10170);
nor U15345 (N_15345,N_10244,N_8784);
xor U15346 (N_15346,N_9802,N_11338);
nand U15347 (N_15347,N_10152,N_9683);
and U15348 (N_15348,N_7433,N_7956);
nor U15349 (N_15349,N_11917,N_9115);
nor U15350 (N_15350,N_6247,N_9430);
nor U15351 (N_15351,N_6287,N_6990);
nor U15352 (N_15352,N_8064,N_11826);
nor U15353 (N_15353,N_6480,N_7771);
or U15354 (N_15354,N_11704,N_10327);
nand U15355 (N_15355,N_8705,N_6770);
nand U15356 (N_15356,N_9458,N_6909);
nand U15357 (N_15357,N_6268,N_6185);
nor U15358 (N_15358,N_6360,N_6237);
nand U15359 (N_15359,N_11314,N_8886);
nand U15360 (N_15360,N_8511,N_6602);
and U15361 (N_15361,N_7042,N_10230);
or U15362 (N_15362,N_7218,N_11547);
or U15363 (N_15363,N_9163,N_10688);
nand U15364 (N_15364,N_9176,N_10639);
nand U15365 (N_15365,N_8279,N_11550);
or U15366 (N_15366,N_11270,N_8286);
nor U15367 (N_15367,N_8530,N_10013);
nor U15368 (N_15368,N_9452,N_11569);
nor U15369 (N_15369,N_9160,N_11828);
and U15370 (N_15370,N_7507,N_11837);
or U15371 (N_15371,N_7929,N_8441);
or U15372 (N_15372,N_7954,N_8799);
or U15373 (N_15373,N_10712,N_9753);
nor U15374 (N_15374,N_10920,N_8224);
xor U15375 (N_15375,N_6918,N_9069);
and U15376 (N_15376,N_8529,N_10342);
nand U15377 (N_15377,N_6842,N_11958);
nor U15378 (N_15378,N_9393,N_10853);
nand U15379 (N_15379,N_7628,N_10478);
xnor U15380 (N_15380,N_10205,N_8612);
xnor U15381 (N_15381,N_6810,N_7908);
and U15382 (N_15382,N_11764,N_6737);
nor U15383 (N_15383,N_6142,N_7034);
and U15384 (N_15384,N_9398,N_6838);
and U15385 (N_15385,N_8893,N_7349);
nor U15386 (N_15386,N_7993,N_7001);
or U15387 (N_15387,N_7475,N_8707);
nor U15388 (N_15388,N_7708,N_11614);
and U15389 (N_15389,N_8894,N_7376);
xor U15390 (N_15390,N_9981,N_8339);
nand U15391 (N_15391,N_11629,N_7403);
or U15392 (N_15392,N_10065,N_6762);
and U15393 (N_15393,N_6947,N_7151);
or U15394 (N_15394,N_7979,N_11704);
xnor U15395 (N_15395,N_9999,N_6563);
nor U15396 (N_15396,N_11805,N_7333);
nand U15397 (N_15397,N_11711,N_7246);
nor U15398 (N_15398,N_11823,N_9862);
nor U15399 (N_15399,N_9688,N_11382);
or U15400 (N_15400,N_6000,N_8466);
or U15401 (N_15401,N_10982,N_11695);
or U15402 (N_15402,N_9449,N_11952);
and U15403 (N_15403,N_10247,N_9103);
or U15404 (N_15404,N_10702,N_7778);
nor U15405 (N_15405,N_10285,N_8016);
xnor U15406 (N_15406,N_10044,N_10496);
or U15407 (N_15407,N_6999,N_11272);
nor U15408 (N_15408,N_10200,N_10575);
nor U15409 (N_15409,N_8853,N_6423);
nor U15410 (N_15410,N_8058,N_9703);
xnor U15411 (N_15411,N_9136,N_8394);
nand U15412 (N_15412,N_11503,N_11530);
or U15413 (N_15413,N_10026,N_7228);
xnor U15414 (N_15414,N_8061,N_11979);
or U15415 (N_15415,N_6321,N_9681);
or U15416 (N_15416,N_6366,N_11710);
and U15417 (N_15417,N_6167,N_7761);
and U15418 (N_15418,N_9662,N_6696);
or U15419 (N_15419,N_9867,N_6910);
and U15420 (N_15420,N_9800,N_7734);
nor U15421 (N_15421,N_6513,N_6326);
xor U15422 (N_15422,N_6530,N_9531);
nor U15423 (N_15423,N_9961,N_10604);
or U15424 (N_15424,N_6766,N_9501);
xor U15425 (N_15425,N_10490,N_11345);
or U15426 (N_15426,N_8479,N_11597);
nand U15427 (N_15427,N_10226,N_6627);
or U15428 (N_15428,N_6467,N_11424);
or U15429 (N_15429,N_11433,N_11818);
nand U15430 (N_15430,N_11248,N_7266);
and U15431 (N_15431,N_11653,N_10055);
and U15432 (N_15432,N_8439,N_10950);
and U15433 (N_15433,N_11756,N_7852);
or U15434 (N_15434,N_9153,N_10199);
nor U15435 (N_15435,N_7290,N_7338);
or U15436 (N_15436,N_10897,N_10606);
nor U15437 (N_15437,N_10411,N_11486);
nand U15438 (N_15438,N_6980,N_6637);
or U15439 (N_15439,N_7912,N_10178);
and U15440 (N_15440,N_7161,N_6699);
nand U15441 (N_15441,N_9901,N_6792);
nor U15442 (N_15442,N_11665,N_7876);
and U15443 (N_15443,N_8489,N_10363);
and U15444 (N_15444,N_6602,N_11152);
nand U15445 (N_15445,N_9346,N_8497);
and U15446 (N_15446,N_7872,N_6581);
and U15447 (N_15447,N_9427,N_7686);
nand U15448 (N_15448,N_9314,N_8437);
nand U15449 (N_15449,N_10976,N_7937);
nor U15450 (N_15450,N_6084,N_11631);
or U15451 (N_15451,N_11835,N_6475);
xnor U15452 (N_15452,N_10796,N_9023);
nor U15453 (N_15453,N_7281,N_8455);
xor U15454 (N_15454,N_10348,N_11995);
nor U15455 (N_15455,N_6496,N_9744);
or U15456 (N_15456,N_10544,N_10070);
xor U15457 (N_15457,N_10947,N_11937);
xnor U15458 (N_15458,N_11959,N_9078);
nor U15459 (N_15459,N_6814,N_8726);
xor U15460 (N_15460,N_10684,N_9303);
nor U15461 (N_15461,N_10321,N_7104);
xor U15462 (N_15462,N_9933,N_10055);
or U15463 (N_15463,N_7844,N_8528);
nand U15464 (N_15464,N_7030,N_10045);
nand U15465 (N_15465,N_6789,N_11351);
and U15466 (N_15466,N_10736,N_6129);
or U15467 (N_15467,N_6118,N_8935);
xnor U15468 (N_15468,N_6465,N_7068);
and U15469 (N_15469,N_11056,N_7010);
nor U15470 (N_15470,N_11739,N_8458);
and U15471 (N_15471,N_6862,N_10160);
nand U15472 (N_15472,N_9855,N_8640);
nor U15473 (N_15473,N_11614,N_7434);
nor U15474 (N_15474,N_6399,N_10025);
and U15475 (N_15475,N_10851,N_8652);
or U15476 (N_15476,N_10698,N_10417);
nor U15477 (N_15477,N_11213,N_9489);
or U15478 (N_15478,N_8619,N_6604);
or U15479 (N_15479,N_10671,N_9461);
and U15480 (N_15480,N_11168,N_8823);
or U15481 (N_15481,N_7210,N_7112);
nand U15482 (N_15482,N_7672,N_7429);
or U15483 (N_15483,N_6287,N_11659);
and U15484 (N_15484,N_7268,N_10555);
or U15485 (N_15485,N_8319,N_11204);
nand U15486 (N_15486,N_7023,N_10976);
nor U15487 (N_15487,N_10734,N_9912);
and U15488 (N_15488,N_9965,N_11339);
xnor U15489 (N_15489,N_9571,N_10644);
or U15490 (N_15490,N_10730,N_11265);
or U15491 (N_15491,N_9741,N_9771);
and U15492 (N_15492,N_9004,N_10813);
or U15493 (N_15493,N_7106,N_6807);
or U15494 (N_15494,N_8781,N_11535);
nand U15495 (N_15495,N_10288,N_10979);
nor U15496 (N_15496,N_6934,N_9064);
or U15497 (N_15497,N_9459,N_6015);
or U15498 (N_15498,N_9504,N_9666);
xnor U15499 (N_15499,N_7737,N_8034);
or U15500 (N_15500,N_7797,N_6611);
and U15501 (N_15501,N_6782,N_8722);
nor U15502 (N_15502,N_11170,N_8682);
nor U15503 (N_15503,N_8682,N_9875);
nand U15504 (N_15504,N_6494,N_10364);
or U15505 (N_15505,N_6664,N_6342);
nor U15506 (N_15506,N_10985,N_9943);
xor U15507 (N_15507,N_9410,N_10836);
nand U15508 (N_15508,N_8052,N_7821);
xor U15509 (N_15509,N_10873,N_8954);
and U15510 (N_15510,N_8175,N_7636);
xor U15511 (N_15511,N_11797,N_7894);
nand U15512 (N_15512,N_9681,N_10013);
and U15513 (N_15513,N_10786,N_9021);
or U15514 (N_15514,N_8046,N_8501);
or U15515 (N_15515,N_9707,N_11139);
and U15516 (N_15516,N_10634,N_7659);
nor U15517 (N_15517,N_11295,N_9949);
nand U15518 (N_15518,N_7557,N_9934);
nor U15519 (N_15519,N_6999,N_8066);
nand U15520 (N_15520,N_9242,N_8351);
nand U15521 (N_15521,N_10201,N_7303);
or U15522 (N_15522,N_9520,N_8434);
nand U15523 (N_15523,N_8966,N_11846);
nand U15524 (N_15524,N_10219,N_9206);
nor U15525 (N_15525,N_7258,N_6992);
or U15526 (N_15526,N_9959,N_9923);
and U15527 (N_15527,N_11181,N_8973);
and U15528 (N_15528,N_9322,N_7172);
nor U15529 (N_15529,N_9256,N_9613);
or U15530 (N_15530,N_7745,N_8713);
nor U15531 (N_15531,N_8509,N_9133);
nor U15532 (N_15532,N_9849,N_11902);
and U15533 (N_15533,N_9310,N_6800);
or U15534 (N_15534,N_10722,N_8190);
and U15535 (N_15535,N_8266,N_7547);
nand U15536 (N_15536,N_8187,N_8354);
or U15537 (N_15537,N_11415,N_8791);
nor U15538 (N_15538,N_7189,N_7126);
xnor U15539 (N_15539,N_6634,N_11745);
or U15540 (N_15540,N_8160,N_10529);
nor U15541 (N_15541,N_6797,N_8982);
and U15542 (N_15542,N_8157,N_7364);
or U15543 (N_15543,N_6022,N_8162);
xor U15544 (N_15544,N_10891,N_11631);
xor U15545 (N_15545,N_10581,N_7619);
or U15546 (N_15546,N_6537,N_6168);
nand U15547 (N_15547,N_8201,N_11150);
nand U15548 (N_15548,N_10548,N_10425);
and U15549 (N_15549,N_10041,N_8036);
nor U15550 (N_15550,N_10663,N_9336);
xor U15551 (N_15551,N_7157,N_10357);
nor U15552 (N_15552,N_11765,N_7943);
nor U15553 (N_15553,N_7083,N_6613);
or U15554 (N_15554,N_10968,N_6445);
nand U15555 (N_15555,N_11748,N_10090);
nor U15556 (N_15556,N_8441,N_7162);
xor U15557 (N_15557,N_8809,N_9549);
xnor U15558 (N_15558,N_10202,N_8258);
or U15559 (N_15559,N_11370,N_10336);
and U15560 (N_15560,N_9253,N_10649);
and U15561 (N_15561,N_7253,N_11181);
xnor U15562 (N_15562,N_6726,N_10200);
nor U15563 (N_15563,N_9811,N_7777);
and U15564 (N_15564,N_10794,N_10547);
and U15565 (N_15565,N_11568,N_6192);
nor U15566 (N_15566,N_9275,N_8554);
and U15567 (N_15567,N_7253,N_8951);
nand U15568 (N_15568,N_6652,N_6794);
nor U15569 (N_15569,N_8398,N_9690);
and U15570 (N_15570,N_10123,N_11604);
xor U15571 (N_15571,N_8350,N_6854);
and U15572 (N_15572,N_6968,N_6430);
and U15573 (N_15573,N_6794,N_11175);
xnor U15574 (N_15574,N_10418,N_7197);
nor U15575 (N_15575,N_6884,N_8888);
and U15576 (N_15576,N_6890,N_9180);
and U15577 (N_15577,N_8545,N_10061);
or U15578 (N_15578,N_7385,N_10734);
nor U15579 (N_15579,N_6767,N_10143);
nand U15580 (N_15580,N_11670,N_7708);
xor U15581 (N_15581,N_10124,N_11792);
xnor U15582 (N_15582,N_11803,N_6974);
nand U15583 (N_15583,N_10191,N_6542);
or U15584 (N_15584,N_9985,N_6964);
nand U15585 (N_15585,N_7370,N_6820);
and U15586 (N_15586,N_10045,N_7867);
nor U15587 (N_15587,N_9317,N_8574);
or U15588 (N_15588,N_11745,N_9083);
or U15589 (N_15589,N_10691,N_10793);
nand U15590 (N_15590,N_6751,N_11112);
and U15591 (N_15591,N_7731,N_7619);
or U15592 (N_15592,N_7175,N_11818);
and U15593 (N_15593,N_7749,N_8255);
xor U15594 (N_15594,N_9889,N_7130);
or U15595 (N_15595,N_8510,N_7156);
nor U15596 (N_15596,N_10771,N_8849);
xnor U15597 (N_15597,N_7161,N_6613);
nand U15598 (N_15598,N_11695,N_9229);
xnor U15599 (N_15599,N_7871,N_6740);
and U15600 (N_15600,N_6923,N_10574);
or U15601 (N_15601,N_10716,N_6444);
or U15602 (N_15602,N_9318,N_11743);
nor U15603 (N_15603,N_10272,N_7702);
and U15604 (N_15604,N_8820,N_8287);
xnor U15605 (N_15605,N_6071,N_8029);
nor U15606 (N_15606,N_10077,N_9117);
or U15607 (N_15607,N_10188,N_10530);
nor U15608 (N_15608,N_8229,N_10528);
nand U15609 (N_15609,N_11019,N_6791);
or U15610 (N_15610,N_9864,N_9853);
nor U15611 (N_15611,N_6035,N_9039);
nand U15612 (N_15612,N_6058,N_9164);
nand U15613 (N_15613,N_6658,N_11942);
nor U15614 (N_15614,N_8805,N_6056);
xnor U15615 (N_15615,N_9914,N_11418);
nor U15616 (N_15616,N_6134,N_8031);
nand U15617 (N_15617,N_8122,N_7689);
nor U15618 (N_15618,N_6338,N_7296);
nand U15619 (N_15619,N_10080,N_6736);
and U15620 (N_15620,N_8080,N_9211);
nor U15621 (N_15621,N_10777,N_6288);
nand U15622 (N_15622,N_10943,N_9740);
or U15623 (N_15623,N_6511,N_8688);
and U15624 (N_15624,N_8885,N_10012);
xnor U15625 (N_15625,N_7743,N_6241);
nor U15626 (N_15626,N_9665,N_11363);
or U15627 (N_15627,N_6049,N_11833);
and U15628 (N_15628,N_8027,N_10095);
or U15629 (N_15629,N_10525,N_11447);
and U15630 (N_15630,N_11792,N_9634);
xor U15631 (N_15631,N_9880,N_8923);
nand U15632 (N_15632,N_11525,N_10187);
or U15633 (N_15633,N_10072,N_6482);
nor U15634 (N_15634,N_10667,N_10549);
nand U15635 (N_15635,N_8508,N_6040);
and U15636 (N_15636,N_10017,N_9525);
and U15637 (N_15637,N_9135,N_7235);
nor U15638 (N_15638,N_8370,N_6229);
or U15639 (N_15639,N_10743,N_9286);
nand U15640 (N_15640,N_6238,N_8968);
and U15641 (N_15641,N_6290,N_6789);
nor U15642 (N_15642,N_11737,N_6038);
and U15643 (N_15643,N_7793,N_6381);
or U15644 (N_15644,N_9046,N_6434);
nand U15645 (N_15645,N_7275,N_10830);
and U15646 (N_15646,N_8446,N_6088);
nand U15647 (N_15647,N_7771,N_8687);
and U15648 (N_15648,N_7881,N_10456);
nand U15649 (N_15649,N_9249,N_8299);
or U15650 (N_15650,N_11405,N_6827);
nor U15651 (N_15651,N_9874,N_7749);
nor U15652 (N_15652,N_8550,N_9992);
nand U15653 (N_15653,N_9363,N_7892);
and U15654 (N_15654,N_7986,N_7648);
nor U15655 (N_15655,N_8247,N_7488);
and U15656 (N_15656,N_11296,N_8181);
nand U15657 (N_15657,N_11281,N_10532);
or U15658 (N_15658,N_6448,N_7239);
nor U15659 (N_15659,N_11287,N_6208);
nor U15660 (N_15660,N_11771,N_7916);
nand U15661 (N_15661,N_10815,N_9933);
nand U15662 (N_15662,N_7325,N_8277);
nand U15663 (N_15663,N_10625,N_7430);
and U15664 (N_15664,N_7543,N_8881);
or U15665 (N_15665,N_8848,N_10388);
nand U15666 (N_15666,N_11230,N_8691);
nand U15667 (N_15667,N_11533,N_9172);
nor U15668 (N_15668,N_8121,N_11270);
or U15669 (N_15669,N_7081,N_9171);
and U15670 (N_15670,N_7267,N_8053);
xor U15671 (N_15671,N_10884,N_7928);
and U15672 (N_15672,N_11104,N_6668);
or U15673 (N_15673,N_7635,N_11962);
and U15674 (N_15674,N_10151,N_10519);
nor U15675 (N_15675,N_7623,N_8915);
nand U15676 (N_15676,N_11918,N_7514);
and U15677 (N_15677,N_7032,N_10500);
nor U15678 (N_15678,N_10091,N_6492);
nor U15679 (N_15679,N_11910,N_8582);
and U15680 (N_15680,N_8972,N_8148);
nand U15681 (N_15681,N_7260,N_11067);
or U15682 (N_15682,N_10492,N_7456);
nor U15683 (N_15683,N_9025,N_6065);
nor U15684 (N_15684,N_10859,N_8320);
and U15685 (N_15685,N_6249,N_7314);
and U15686 (N_15686,N_7766,N_6502);
nand U15687 (N_15687,N_8755,N_6658);
nor U15688 (N_15688,N_11303,N_7500);
nor U15689 (N_15689,N_9718,N_8590);
and U15690 (N_15690,N_10878,N_10007);
xnor U15691 (N_15691,N_6789,N_7026);
or U15692 (N_15692,N_7692,N_10654);
or U15693 (N_15693,N_11096,N_9740);
nand U15694 (N_15694,N_11805,N_7954);
and U15695 (N_15695,N_10923,N_7442);
nor U15696 (N_15696,N_8968,N_11678);
nor U15697 (N_15697,N_6940,N_11235);
nand U15698 (N_15698,N_11728,N_6329);
nor U15699 (N_15699,N_10822,N_8229);
nand U15700 (N_15700,N_7548,N_7665);
or U15701 (N_15701,N_7784,N_10386);
and U15702 (N_15702,N_8382,N_6859);
or U15703 (N_15703,N_7016,N_10213);
nor U15704 (N_15704,N_7562,N_7056);
and U15705 (N_15705,N_9173,N_9199);
xnor U15706 (N_15706,N_6385,N_11471);
and U15707 (N_15707,N_7022,N_9977);
or U15708 (N_15708,N_11522,N_11616);
nand U15709 (N_15709,N_10378,N_7195);
nand U15710 (N_15710,N_8519,N_7638);
or U15711 (N_15711,N_9877,N_8373);
nand U15712 (N_15712,N_8823,N_11905);
nor U15713 (N_15713,N_7817,N_6475);
nor U15714 (N_15714,N_10796,N_7975);
nand U15715 (N_15715,N_6441,N_9257);
or U15716 (N_15716,N_10664,N_6973);
and U15717 (N_15717,N_7019,N_8402);
nand U15718 (N_15718,N_6596,N_8945);
nand U15719 (N_15719,N_6197,N_8342);
or U15720 (N_15720,N_8748,N_7103);
and U15721 (N_15721,N_11155,N_6951);
or U15722 (N_15722,N_9474,N_9687);
and U15723 (N_15723,N_6235,N_10386);
and U15724 (N_15724,N_10398,N_8752);
and U15725 (N_15725,N_7658,N_7225);
nand U15726 (N_15726,N_8183,N_6363);
nand U15727 (N_15727,N_7874,N_11980);
nand U15728 (N_15728,N_6354,N_8243);
nand U15729 (N_15729,N_11726,N_9360);
nor U15730 (N_15730,N_6644,N_6325);
and U15731 (N_15731,N_11818,N_10931);
or U15732 (N_15732,N_8614,N_10553);
xor U15733 (N_15733,N_11698,N_11664);
xnor U15734 (N_15734,N_9863,N_9174);
nor U15735 (N_15735,N_11344,N_11449);
and U15736 (N_15736,N_11018,N_6062);
or U15737 (N_15737,N_8701,N_9219);
or U15738 (N_15738,N_10427,N_9896);
xor U15739 (N_15739,N_11953,N_7805);
or U15740 (N_15740,N_6130,N_7139);
nor U15741 (N_15741,N_6798,N_10128);
nand U15742 (N_15742,N_8260,N_7707);
or U15743 (N_15743,N_11094,N_10182);
nand U15744 (N_15744,N_9094,N_7652);
and U15745 (N_15745,N_11135,N_7308);
nand U15746 (N_15746,N_7311,N_6224);
nand U15747 (N_15747,N_6132,N_6368);
and U15748 (N_15748,N_9244,N_11934);
and U15749 (N_15749,N_10298,N_6210);
and U15750 (N_15750,N_10227,N_7222);
or U15751 (N_15751,N_9926,N_7883);
nand U15752 (N_15752,N_8718,N_6278);
nand U15753 (N_15753,N_11842,N_8040);
xnor U15754 (N_15754,N_9441,N_6083);
or U15755 (N_15755,N_11846,N_8786);
nor U15756 (N_15756,N_11043,N_9642);
nand U15757 (N_15757,N_7075,N_7648);
and U15758 (N_15758,N_11262,N_9209);
or U15759 (N_15759,N_6010,N_9316);
or U15760 (N_15760,N_7587,N_7070);
nand U15761 (N_15761,N_8990,N_11583);
nor U15762 (N_15762,N_6371,N_11706);
nand U15763 (N_15763,N_11726,N_9687);
nand U15764 (N_15764,N_7616,N_7364);
nand U15765 (N_15765,N_11330,N_9852);
nor U15766 (N_15766,N_8654,N_11012);
nor U15767 (N_15767,N_10083,N_6944);
nor U15768 (N_15768,N_6044,N_9168);
nor U15769 (N_15769,N_8271,N_11057);
nand U15770 (N_15770,N_6288,N_7044);
xor U15771 (N_15771,N_10642,N_7217);
and U15772 (N_15772,N_11106,N_8060);
or U15773 (N_15773,N_11243,N_6692);
nor U15774 (N_15774,N_9828,N_8185);
or U15775 (N_15775,N_9295,N_10457);
nor U15776 (N_15776,N_9980,N_10692);
or U15777 (N_15777,N_6801,N_9458);
nor U15778 (N_15778,N_10355,N_11307);
xnor U15779 (N_15779,N_8524,N_7136);
nand U15780 (N_15780,N_8358,N_8382);
nand U15781 (N_15781,N_11421,N_11792);
nor U15782 (N_15782,N_6485,N_8692);
nand U15783 (N_15783,N_6360,N_7582);
and U15784 (N_15784,N_7273,N_6149);
nand U15785 (N_15785,N_6953,N_11668);
and U15786 (N_15786,N_6241,N_10210);
or U15787 (N_15787,N_7995,N_10169);
nand U15788 (N_15788,N_11914,N_11594);
and U15789 (N_15789,N_7333,N_7309);
nand U15790 (N_15790,N_7765,N_9019);
or U15791 (N_15791,N_11676,N_8227);
nand U15792 (N_15792,N_11941,N_6408);
nor U15793 (N_15793,N_10007,N_10947);
and U15794 (N_15794,N_7978,N_7806);
nor U15795 (N_15795,N_10085,N_9696);
nand U15796 (N_15796,N_8558,N_6971);
and U15797 (N_15797,N_11673,N_7645);
nand U15798 (N_15798,N_11249,N_10977);
nand U15799 (N_15799,N_10497,N_8809);
nand U15800 (N_15800,N_6844,N_9748);
or U15801 (N_15801,N_7103,N_9326);
nor U15802 (N_15802,N_8830,N_11641);
or U15803 (N_15803,N_9359,N_7644);
or U15804 (N_15804,N_11589,N_8633);
nand U15805 (N_15805,N_9460,N_6415);
and U15806 (N_15806,N_11935,N_10665);
xor U15807 (N_15807,N_9291,N_8426);
nor U15808 (N_15808,N_9137,N_9825);
or U15809 (N_15809,N_6080,N_9211);
nor U15810 (N_15810,N_10181,N_9730);
nand U15811 (N_15811,N_9828,N_9219);
and U15812 (N_15812,N_8904,N_6327);
or U15813 (N_15813,N_10157,N_8203);
nor U15814 (N_15814,N_9063,N_11832);
nor U15815 (N_15815,N_7335,N_11743);
and U15816 (N_15816,N_6308,N_10437);
and U15817 (N_15817,N_8778,N_7759);
nand U15818 (N_15818,N_10116,N_9723);
and U15819 (N_15819,N_8456,N_8716);
and U15820 (N_15820,N_10541,N_11630);
and U15821 (N_15821,N_8357,N_11317);
and U15822 (N_15822,N_11366,N_9993);
nor U15823 (N_15823,N_9712,N_7357);
or U15824 (N_15824,N_6959,N_9618);
nor U15825 (N_15825,N_10544,N_8606);
nand U15826 (N_15826,N_7947,N_11869);
xnor U15827 (N_15827,N_9018,N_8014);
nand U15828 (N_15828,N_6557,N_9539);
or U15829 (N_15829,N_11821,N_6000);
nand U15830 (N_15830,N_9321,N_6251);
nor U15831 (N_15831,N_9831,N_10836);
or U15832 (N_15832,N_11737,N_11218);
and U15833 (N_15833,N_8542,N_6381);
or U15834 (N_15834,N_8982,N_9993);
nand U15835 (N_15835,N_8186,N_9027);
nor U15836 (N_15836,N_11711,N_6920);
nor U15837 (N_15837,N_7677,N_11790);
or U15838 (N_15838,N_6362,N_9714);
nand U15839 (N_15839,N_10605,N_8023);
nor U15840 (N_15840,N_6943,N_6173);
and U15841 (N_15841,N_7628,N_7099);
nand U15842 (N_15842,N_7661,N_10501);
and U15843 (N_15843,N_7090,N_11587);
nor U15844 (N_15844,N_11531,N_8027);
nor U15845 (N_15845,N_7185,N_9478);
nand U15846 (N_15846,N_10524,N_6894);
and U15847 (N_15847,N_7465,N_11026);
or U15848 (N_15848,N_6321,N_6770);
or U15849 (N_15849,N_8826,N_6372);
nor U15850 (N_15850,N_8650,N_6753);
nor U15851 (N_15851,N_6281,N_7303);
nand U15852 (N_15852,N_8544,N_9705);
nor U15853 (N_15853,N_8677,N_9504);
nor U15854 (N_15854,N_6051,N_8698);
nor U15855 (N_15855,N_9786,N_7675);
nor U15856 (N_15856,N_9086,N_8341);
nor U15857 (N_15857,N_10188,N_9039);
nor U15858 (N_15858,N_9064,N_10973);
nor U15859 (N_15859,N_7093,N_9831);
nand U15860 (N_15860,N_6049,N_6293);
or U15861 (N_15861,N_10408,N_6447);
nand U15862 (N_15862,N_6207,N_10451);
and U15863 (N_15863,N_7130,N_7465);
or U15864 (N_15864,N_7003,N_11974);
and U15865 (N_15865,N_8712,N_8163);
nor U15866 (N_15866,N_10516,N_9065);
nand U15867 (N_15867,N_10009,N_7919);
nand U15868 (N_15868,N_9473,N_8059);
nor U15869 (N_15869,N_8548,N_10144);
or U15870 (N_15870,N_8728,N_9474);
nand U15871 (N_15871,N_8222,N_9925);
or U15872 (N_15872,N_6556,N_9160);
nand U15873 (N_15873,N_9320,N_10334);
nand U15874 (N_15874,N_10362,N_7888);
nor U15875 (N_15875,N_9313,N_8649);
and U15876 (N_15876,N_6502,N_10455);
nor U15877 (N_15877,N_9687,N_11441);
or U15878 (N_15878,N_7997,N_7495);
or U15879 (N_15879,N_6663,N_6987);
or U15880 (N_15880,N_6900,N_11951);
nor U15881 (N_15881,N_8874,N_9544);
xor U15882 (N_15882,N_9776,N_10820);
or U15883 (N_15883,N_11906,N_7117);
or U15884 (N_15884,N_11532,N_7925);
and U15885 (N_15885,N_9101,N_10000);
nand U15886 (N_15886,N_11794,N_6763);
nor U15887 (N_15887,N_8285,N_6171);
nand U15888 (N_15888,N_10650,N_7834);
and U15889 (N_15889,N_10068,N_9258);
nor U15890 (N_15890,N_10018,N_10708);
and U15891 (N_15891,N_10760,N_11694);
or U15892 (N_15892,N_9382,N_10863);
or U15893 (N_15893,N_8079,N_7191);
or U15894 (N_15894,N_11614,N_10793);
nand U15895 (N_15895,N_8872,N_10323);
xnor U15896 (N_15896,N_9270,N_7737);
nor U15897 (N_15897,N_11566,N_6625);
and U15898 (N_15898,N_10758,N_11251);
and U15899 (N_15899,N_7783,N_10548);
nand U15900 (N_15900,N_10050,N_9404);
nand U15901 (N_15901,N_10520,N_11295);
and U15902 (N_15902,N_10125,N_9427);
and U15903 (N_15903,N_10260,N_8673);
or U15904 (N_15904,N_7757,N_10768);
nand U15905 (N_15905,N_6121,N_6947);
nor U15906 (N_15906,N_7619,N_10649);
nor U15907 (N_15907,N_9210,N_7644);
nand U15908 (N_15908,N_11252,N_11686);
nor U15909 (N_15909,N_10963,N_7024);
nor U15910 (N_15910,N_10984,N_8519);
nor U15911 (N_15911,N_8247,N_11419);
xor U15912 (N_15912,N_9025,N_11511);
or U15913 (N_15913,N_7459,N_7484);
nand U15914 (N_15914,N_6350,N_7171);
xnor U15915 (N_15915,N_6811,N_10201);
nand U15916 (N_15916,N_7414,N_10281);
nor U15917 (N_15917,N_6338,N_7560);
or U15918 (N_15918,N_8496,N_11771);
nand U15919 (N_15919,N_8659,N_8358);
or U15920 (N_15920,N_8266,N_9408);
nor U15921 (N_15921,N_10654,N_7191);
or U15922 (N_15922,N_11051,N_11467);
nor U15923 (N_15923,N_10619,N_9336);
or U15924 (N_15924,N_7631,N_11209);
nor U15925 (N_15925,N_10677,N_9983);
xor U15926 (N_15926,N_9333,N_9832);
nand U15927 (N_15927,N_10660,N_8453);
and U15928 (N_15928,N_6582,N_6446);
nand U15929 (N_15929,N_11088,N_8845);
or U15930 (N_15930,N_9515,N_7212);
nor U15931 (N_15931,N_8660,N_7882);
and U15932 (N_15932,N_10845,N_10057);
or U15933 (N_15933,N_9347,N_11749);
and U15934 (N_15934,N_9824,N_6810);
nor U15935 (N_15935,N_10462,N_8161);
and U15936 (N_15936,N_8996,N_8736);
nand U15937 (N_15937,N_9379,N_7469);
or U15938 (N_15938,N_10583,N_11249);
xnor U15939 (N_15939,N_6456,N_9552);
nor U15940 (N_15940,N_10653,N_8315);
nor U15941 (N_15941,N_6903,N_9186);
xor U15942 (N_15942,N_10707,N_11855);
nor U15943 (N_15943,N_6133,N_9825);
or U15944 (N_15944,N_10246,N_8338);
nand U15945 (N_15945,N_9076,N_9218);
nand U15946 (N_15946,N_11437,N_8003);
nand U15947 (N_15947,N_8421,N_6055);
or U15948 (N_15948,N_9601,N_9505);
nor U15949 (N_15949,N_9351,N_6495);
nand U15950 (N_15950,N_7980,N_10813);
xor U15951 (N_15951,N_8603,N_6992);
and U15952 (N_15952,N_6299,N_8607);
nor U15953 (N_15953,N_9131,N_7134);
nand U15954 (N_15954,N_9291,N_7005);
nand U15955 (N_15955,N_10558,N_10453);
nor U15956 (N_15956,N_11137,N_7230);
nand U15957 (N_15957,N_6685,N_7459);
nand U15958 (N_15958,N_10300,N_7136);
and U15959 (N_15959,N_10758,N_6298);
or U15960 (N_15960,N_6598,N_9290);
xor U15961 (N_15961,N_11799,N_6930);
or U15962 (N_15962,N_7597,N_10628);
nand U15963 (N_15963,N_9816,N_7562);
or U15964 (N_15964,N_8869,N_10091);
and U15965 (N_15965,N_6549,N_11958);
or U15966 (N_15966,N_6109,N_6657);
xnor U15967 (N_15967,N_9311,N_10863);
or U15968 (N_15968,N_6044,N_6884);
or U15969 (N_15969,N_10177,N_8153);
or U15970 (N_15970,N_7165,N_11504);
and U15971 (N_15971,N_11551,N_10596);
and U15972 (N_15972,N_8011,N_11599);
or U15973 (N_15973,N_9903,N_7891);
nor U15974 (N_15974,N_6588,N_6374);
nand U15975 (N_15975,N_7878,N_8837);
xnor U15976 (N_15976,N_8804,N_10653);
or U15977 (N_15977,N_9830,N_10338);
nand U15978 (N_15978,N_7682,N_11612);
and U15979 (N_15979,N_6093,N_11741);
or U15980 (N_15980,N_11071,N_11290);
nand U15981 (N_15981,N_6980,N_9109);
and U15982 (N_15982,N_7719,N_6947);
or U15983 (N_15983,N_9261,N_10219);
or U15984 (N_15984,N_9408,N_10725);
or U15985 (N_15985,N_9829,N_8389);
and U15986 (N_15986,N_9140,N_7136);
nand U15987 (N_15987,N_11279,N_9203);
nor U15988 (N_15988,N_10649,N_8179);
nor U15989 (N_15989,N_8992,N_8913);
and U15990 (N_15990,N_11268,N_8950);
or U15991 (N_15991,N_6889,N_9688);
and U15992 (N_15992,N_11802,N_9500);
nor U15993 (N_15993,N_9566,N_10374);
nor U15994 (N_15994,N_10315,N_9896);
nor U15995 (N_15995,N_11479,N_6280);
nand U15996 (N_15996,N_6077,N_11208);
nor U15997 (N_15997,N_7641,N_10862);
and U15998 (N_15998,N_8317,N_8658);
nand U15999 (N_15999,N_6823,N_9655);
xor U16000 (N_16000,N_11336,N_9842);
nor U16001 (N_16001,N_11859,N_7509);
and U16002 (N_16002,N_8829,N_10607);
nand U16003 (N_16003,N_9734,N_8181);
and U16004 (N_16004,N_11452,N_6170);
or U16005 (N_16005,N_7938,N_8521);
xor U16006 (N_16006,N_6893,N_6501);
and U16007 (N_16007,N_6054,N_8876);
and U16008 (N_16008,N_10476,N_7363);
or U16009 (N_16009,N_6027,N_10053);
or U16010 (N_16010,N_11854,N_11796);
nor U16011 (N_16011,N_10512,N_10497);
or U16012 (N_16012,N_6235,N_8648);
nand U16013 (N_16013,N_6250,N_10311);
and U16014 (N_16014,N_10415,N_8095);
nor U16015 (N_16015,N_6085,N_6469);
nor U16016 (N_16016,N_7236,N_7175);
nor U16017 (N_16017,N_7764,N_6850);
nor U16018 (N_16018,N_8074,N_8384);
nor U16019 (N_16019,N_9138,N_10951);
and U16020 (N_16020,N_7097,N_7557);
or U16021 (N_16021,N_6624,N_8030);
nor U16022 (N_16022,N_10495,N_10561);
nand U16023 (N_16023,N_7502,N_7090);
xnor U16024 (N_16024,N_7677,N_9668);
xor U16025 (N_16025,N_7212,N_6506);
nor U16026 (N_16026,N_11770,N_8768);
nor U16027 (N_16027,N_9427,N_6701);
nor U16028 (N_16028,N_7337,N_10628);
nand U16029 (N_16029,N_8575,N_7478);
and U16030 (N_16030,N_9769,N_10094);
or U16031 (N_16031,N_9315,N_11840);
and U16032 (N_16032,N_7789,N_8438);
nand U16033 (N_16033,N_9665,N_11903);
nor U16034 (N_16034,N_10925,N_6744);
nor U16035 (N_16035,N_7542,N_6887);
nor U16036 (N_16036,N_8309,N_7888);
and U16037 (N_16037,N_11785,N_8837);
nand U16038 (N_16038,N_10037,N_11227);
or U16039 (N_16039,N_11651,N_10865);
or U16040 (N_16040,N_8445,N_10152);
or U16041 (N_16041,N_7430,N_8495);
and U16042 (N_16042,N_10506,N_7628);
and U16043 (N_16043,N_6439,N_6371);
xor U16044 (N_16044,N_6412,N_11824);
nand U16045 (N_16045,N_11388,N_10206);
nand U16046 (N_16046,N_8120,N_7153);
or U16047 (N_16047,N_8000,N_11584);
or U16048 (N_16048,N_6544,N_9014);
nor U16049 (N_16049,N_11073,N_9480);
nor U16050 (N_16050,N_6638,N_6274);
xor U16051 (N_16051,N_10784,N_11598);
and U16052 (N_16052,N_6922,N_7085);
nor U16053 (N_16053,N_10140,N_11458);
nand U16054 (N_16054,N_10902,N_11301);
nor U16055 (N_16055,N_6867,N_6780);
nand U16056 (N_16056,N_6587,N_10070);
nor U16057 (N_16057,N_6650,N_10038);
or U16058 (N_16058,N_7304,N_11899);
nand U16059 (N_16059,N_10913,N_6364);
nand U16060 (N_16060,N_10934,N_7079);
xnor U16061 (N_16061,N_11451,N_6635);
or U16062 (N_16062,N_8126,N_11091);
nor U16063 (N_16063,N_9855,N_6529);
or U16064 (N_16064,N_9189,N_9707);
or U16065 (N_16065,N_10980,N_9904);
and U16066 (N_16066,N_11407,N_7357);
nor U16067 (N_16067,N_6403,N_7727);
or U16068 (N_16068,N_8437,N_7629);
nand U16069 (N_16069,N_6988,N_11767);
or U16070 (N_16070,N_9024,N_7165);
and U16071 (N_16071,N_6095,N_8305);
or U16072 (N_16072,N_11327,N_7213);
or U16073 (N_16073,N_9491,N_6364);
nor U16074 (N_16074,N_6012,N_8569);
and U16075 (N_16075,N_8773,N_6359);
or U16076 (N_16076,N_7609,N_7667);
or U16077 (N_16077,N_6972,N_10420);
nor U16078 (N_16078,N_8130,N_8501);
nand U16079 (N_16079,N_10840,N_9693);
nor U16080 (N_16080,N_8386,N_11580);
nand U16081 (N_16081,N_7632,N_8376);
nor U16082 (N_16082,N_7935,N_7688);
nor U16083 (N_16083,N_9838,N_7099);
nand U16084 (N_16084,N_6195,N_11427);
or U16085 (N_16085,N_10663,N_9949);
and U16086 (N_16086,N_6383,N_8751);
or U16087 (N_16087,N_6637,N_10276);
nor U16088 (N_16088,N_11267,N_10587);
nor U16089 (N_16089,N_11126,N_8436);
nand U16090 (N_16090,N_6282,N_11567);
or U16091 (N_16091,N_11959,N_7864);
nor U16092 (N_16092,N_6733,N_11304);
or U16093 (N_16093,N_9776,N_9252);
nor U16094 (N_16094,N_6906,N_10009);
or U16095 (N_16095,N_11634,N_6032);
nor U16096 (N_16096,N_11432,N_9341);
or U16097 (N_16097,N_7752,N_8530);
nand U16098 (N_16098,N_6703,N_11587);
nand U16099 (N_16099,N_10458,N_9836);
xnor U16100 (N_16100,N_11583,N_6979);
nor U16101 (N_16101,N_11366,N_10845);
or U16102 (N_16102,N_9326,N_8124);
and U16103 (N_16103,N_8134,N_11771);
and U16104 (N_16104,N_9788,N_8003);
nand U16105 (N_16105,N_6815,N_10127);
or U16106 (N_16106,N_9642,N_6797);
nor U16107 (N_16107,N_9299,N_9758);
nand U16108 (N_16108,N_9007,N_6740);
nor U16109 (N_16109,N_8040,N_10597);
nor U16110 (N_16110,N_7168,N_7270);
nor U16111 (N_16111,N_7005,N_7313);
nor U16112 (N_16112,N_10676,N_11835);
and U16113 (N_16113,N_10818,N_10077);
and U16114 (N_16114,N_11898,N_7285);
nand U16115 (N_16115,N_9773,N_6872);
or U16116 (N_16116,N_9731,N_7493);
and U16117 (N_16117,N_9829,N_7847);
nor U16118 (N_16118,N_11745,N_8219);
or U16119 (N_16119,N_7793,N_8047);
nand U16120 (N_16120,N_10174,N_8291);
nand U16121 (N_16121,N_9455,N_6057);
nor U16122 (N_16122,N_7566,N_10663);
nand U16123 (N_16123,N_10434,N_6437);
nor U16124 (N_16124,N_11258,N_7177);
and U16125 (N_16125,N_11791,N_10578);
nand U16126 (N_16126,N_11449,N_9597);
xnor U16127 (N_16127,N_7189,N_9944);
or U16128 (N_16128,N_7278,N_11771);
nand U16129 (N_16129,N_11681,N_8998);
and U16130 (N_16130,N_6960,N_11271);
nand U16131 (N_16131,N_7741,N_6171);
nor U16132 (N_16132,N_8411,N_9724);
nand U16133 (N_16133,N_11418,N_8550);
nor U16134 (N_16134,N_11235,N_6450);
nand U16135 (N_16135,N_7845,N_11811);
nand U16136 (N_16136,N_11892,N_11147);
xnor U16137 (N_16137,N_11594,N_8050);
nand U16138 (N_16138,N_10142,N_7430);
nor U16139 (N_16139,N_9240,N_11023);
or U16140 (N_16140,N_7212,N_7339);
or U16141 (N_16141,N_10074,N_8920);
and U16142 (N_16142,N_6691,N_8574);
and U16143 (N_16143,N_7775,N_6175);
nor U16144 (N_16144,N_6751,N_7244);
nor U16145 (N_16145,N_11135,N_11811);
or U16146 (N_16146,N_9626,N_6665);
and U16147 (N_16147,N_8313,N_6874);
xnor U16148 (N_16148,N_6605,N_9649);
nand U16149 (N_16149,N_11036,N_11155);
or U16150 (N_16150,N_9369,N_10497);
and U16151 (N_16151,N_11468,N_6974);
and U16152 (N_16152,N_8808,N_9538);
nor U16153 (N_16153,N_8354,N_10739);
or U16154 (N_16154,N_6998,N_9513);
or U16155 (N_16155,N_10843,N_9083);
or U16156 (N_16156,N_8941,N_6466);
or U16157 (N_16157,N_7792,N_7962);
and U16158 (N_16158,N_11548,N_11764);
nand U16159 (N_16159,N_6332,N_8693);
nand U16160 (N_16160,N_7917,N_11010);
nor U16161 (N_16161,N_10941,N_11388);
nor U16162 (N_16162,N_11732,N_7649);
xnor U16163 (N_16163,N_10458,N_10442);
nor U16164 (N_16164,N_6027,N_7032);
or U16165 (N_16165,N_10134,N_11645);
nor U16166 (N_16166,N_6758,N_9502);
nand U16167 (N_16167,N_9521,N_8462);
xnor U16168 (N_16168,N_8049,N_11871);
or U16169 (N_16169,N_7018,N_11110);
or U16170 (N_16170,N_7465,N_8886);
nor U16171 (N_16171,N_7058,N_9018);
nand U16172 (N_16172,N_6135,N_8392);
and U16173 (N_16173,N_7336,N_9830);
nand U16174 (N_16174,N_6254,N_10994);
nand U16175 (N_16175,N_7846,N_7270);
nand U16176 (N_16176,N_9319,N_10923);
and U16177 (N_16177,N_6139,N_6316);
nor U16178 (N_16178,N_6270,N_8476);
and U16179 (N_16179,N_9909,N_8458);
or U16180 (N_16180,N_9169,N_9902);
nor U16181 (N_16181,N_8718,N_7829);
nand U16182 (N_16182,N_11422,N_9828);
nor U16183 (N_16183,N_6339,N_7725);
and U16184 (N_16184,N_11888,N_8046);
nor U16185 (N_16185,N_6688,N_11287);
nand U16186 (N_16186,N_8004,N_7308);
nor U16187 (N_16187,N_11152,N_9591);
and U16188 (N_16188,N_11618,N_6349);
and U16189 (N_16189,N_7627,N_11188);
and U16190 (N_16190,N_7793,N_11130);
nand U16191 (N_16191,N_9380,N_7113);
nand U16192 (N_16192,N_9493,N_8713);
and U16193 (N_16193,N_10158,N_11232);
or U16194 (N_16194,N_9545,N_9131);
nand U16195 (N_16195,N_9732,N_9385);
nor U16196 (N_16196,N_11218,N_7878);
nor U16197 (N_16197,N_7352,N_7215);
nand U16198 (N_16198,N_8236,N_6082);
xnor U16199 (N_16199,N_10202,N_6048);
and U16200 (N_16200,N_9121,N_10057);
and U16201 (N_16201,N_10165,N_9830);
nand U16202 (N_16202,N_7522,N_11107);
nor U16203 (N_16203,N_11270,N_8218);
nor U16204 (N_16204,N_7415,N_8245);
xnor U16205 (N_16205,N_8657,N_8213);
or U16206 (N_16206,N_7999,N_6595);
nand U16207 (N_16207,N_9614,N_8175);
or U16208 (N_16208,N_10949,N_11995);
xnor U16209 (N_16209,N_10211,N_6475);
xnor U16210 (N_16210,N_6569,N_9098);
and U16211 (N_16211,N_10198,N_7948);
and U16212 (N_16212,N_9341,N_6670);
nor U16213 (N_16213,N_8924,N_9787);
or U16214 (N_16214,N_11700,N_8019);
nand U16215 (N_16215,N_9692,N_10354);
and U16216 (N_16216,N_10445,N_9132);
nand U16217 (N_16217,N_8205,N_10141);
or U16218 (N_16218,N_11104,N_9917);
nand U16219 (N_16219,N_10873,N_11841);
and U16220 (N_16220,N_11979,N_8005);
and U16221 (N_16221,N_9841,N_11167);
and U16222 (N_16222,N_10296,N_11574);
or U16223 (N_16223,N_10999,N_11389);
nand U16224 (N_16224,N_7580,N_11781);
and U16225 (N_16225,N_6007,N_6759);
or U16226 (N_16226,N_11322,N_9544);
nor U16227 (N_16227,N_8264,N_6876);
nor U16228 (N_16228,N_6765,N_6947);
or U16229 (N_16229,N_7057,N_9341);
and U16230 (N_16230,N_10545,N_10407);
nor U16231 (N_16231,N_9857,N_8261);
xnor U16232 (N_16232,N_11822,N_9964);
nand U16233 (N_16233,N_6673,N_9881);
and U16234 (N_16234,N_6598,N_8810);
nand U16235 (N_16235,N_6092,N_6255);
nor U16236 (N_16236,N_9136,N_6536);
and U16237 (N_16237,N_9477,N_8075);
or U16238 (N_16238,N_10399,N_9764);
and U16239 (N_16239,N_9891,N_7988);
nor U16240 (N_16240,N_9005,N_11222);
nand U16241 (N_16241,N_7204,N_9995);
nand U16242 (N_16242,N_7414,N_10534);
or U16243 (N_16243,N_6892,N_11462);
or U16244 (N_16244,N_8116,N_7454);
or U16245 (N_16245,N_11423,N_10552);
and U16246 (N_16246,N_7989,N_7075);
xor U16247 (N_16247,N_6238,N_9429);
and U16248 (N_16248,N_6288,N_11227);
or U16249 (N_16249,N_10759,N_11006);
and U16250 (N_16250,N_7708,N_6549);
nand U16251 (N_16251,N_7209,N_6928);
and U16252 (N_16252,N_8603,N_7667);
or U16253 (N_16253,N_8805,N_6610);
nand U16254 (N_16254,N_10299,N_8846);
nand U16255 (N_16255,N_11252,N_11984);
nor U16256 (N_16256,N_11991,N_10754);
xnor U16257 (N_16257,N_10495,N_9102);
xor U16258 (N_16258,N_11552,N_7743);
or U16259 (N_16259,N_11138,N_8498);
nor U16260 (N_16260,N_9308,N_6260);
and U16261 (N_16261,N_11860,N_10715);
and U16262 (N_16262,N_10740,N_9174);
nor U16263 (N_16263,N_11029,N_11614);
and U16264 (N_16264,N_11274,N_9769);
and U16265 (N_16265,N_10953,N_10622);
nand U16266 (N_16266,N_7060,N_11203);
xor U16267 (N_16267,N_7861,N_10786);
nand U16268 (N_16268,N_7616,N_10825);
or U16269 (N_16269,N_10059,N_7151);
or U16270 (N_16270,N_7607,N_9365);
or U16271 (N_16271,N_6610,N_10085);
or U16272 (N_16272,N_11971,N_10964);
or U16273 (N_16273,N_7435,N_8538);
nor U16274 (N_16274,N_9758,N_6067);
or U16275 (N_16275,N_11844,N_8835);
and U16276 (N_16276,N_9388,N_11721);
nor U16277 (N_16277,N_10364,N_7867);
or U16278 (N_16278,N_9457,N_6404);
or U16279 (N_16279,N_7309,N_8868);
nor U16280 (N_16280,N_11053,N_9207);
xor U16281 (N_16281,N_6495,N_11352);
nor U16282 (N_16282,N_9926,N_8808);
nor U16283 (N_16283,N_9634,N_8576);
and U16284 (N_16284,N_6710,N_6222);
or U16285 (N_16285,N_6714,N_11111);
or U16286 (N_16286,N_7557,N_11639);
or U16287 (N_16287,N_9151,N_11850);
or U16288 (N_16288,N_10816,N_11708);
or U16289 (N_16289,N_11471,N_7259);
nand U16290 (N_16290,N_11183,N_10468);
nand U16291 (N_16291,N_8828,N_7294);
and U16292 (N_16292,N_8712,N_10538);
nor U16293 (N_16293,N_8227,N_8983);
or U16294 (N_16294,N_8558,N_8918);
and U16295 (N_16295,N_10064,N_7024);
and U16296 (N_16296,N_7029,N_6662);
nand U16297 (N_16297,N_11857,N_11357);
nor U16298 (N_16298,N_7972,N_7674);
or U16299 (N_16299,N_6152,N_8022);
nor U16300 (N_16300,N_6400,N_8951);
and U16301 (N_16301,N_11659,N_11084);
and U16302 (N_16302,N_10189,N_9702);
and U16303 (N_16303,N_6366,N_11829);
nor U16304 (N_16304,N_11611,N_8302);
nor U16305 (N_16305,N_10102,N_10088);
nor U16306 (N_16306,N_9028,N_6001);
and U16307 (N_16307,N_7852,N_8547);
and U16308 (N_16308,N_9683,N_6990);
nor U16309 (N_16309,N_8062,N_10416);
nor U16310 (N_16310,N_11671,N_7433);
and U16311 (N_16311,N_9244,N_7098);
and U16312 (N_16312,N_8339,N_9296);
or U16313 (N_16313,N_7339,N_11918);
and U16314 (N_16314,N_6117,N_10569);
or U16315 (N_16315,N_9442,N_10500);
or U16316 (N_16316,N_10234,N_10984);
or U16317 (N_16317,N_11350,N_11787);
and U16318 (N_16318,N_7719,N_8409);
nand U16319 (N_16319,N_8284,N_9110);
or U16320 (N_16320,N_11497,N_9484);
nor U16321 (N_16321,N_10167,N_9112);
nand U16322 (N_16322,N_11867,N_6304);
nor U16323 (N_16323,N_10483,N_11230);
nor U16324 (N_16324,N_11432,N_8125);
or U16325 (N_16325,N_6007,N_11433);
nor U16326 (N_16326,N_11228,N_10130);
nand U16327 (N_16327,N_10362,N_9014);
or U16328 (N_16328,N_11688,N_6449);
or U16329 (N_16329,N_10072,N_6008);
and U16330 (N_16330,N_10864,N_9399);
or U16331 (N_16331,N_7159,N_10445);
nand U16332 (N_16332,N_9374,N_7327);
and U16333 (N_16333,N_6024,N_10488);
nand U16334 (N_16334,N_7005,N_8728);
or U16335 (N_16335,N_6092,N_6238);
and U16336 (N_16336,N_7647,N_9588);
or U16337 (N_16337,N_9721,N_6686);
nand U16338 (N_16338,N_7117,N_11361);
nor U16339 (N_16339,N_6971,N_6407);
xnor U16340 (N_16340,N_8587,N_8728);
and U16341 (N_16341,N_7091,N_8657);
or U16342 (N_16342,N_7767,N_11699);
or U16343 (N_16343,N_9560,N_11461);
nand U16344 (N_16344,N_6974,N_6916);
and U16345 (N_16345,N_11051,N_7148);
xor U16346 (N_16346,N_7020,N_7431);
and U16347 (N_16347,N_6951,N_10479);
and U16348 (N_16348,N_11629,N_11439);
and U16349 (N_16349,N_7859,N_11698);
and U16350 (N_16350,N_9841,N_11425);
and U16351 (N_16351,N_7732,N_8918);
nor U16352 (N_16352,N_11533,N_6169);
or U16353 (N_16353,N_10148,N_9996);
and U16354 (N_16354,N_7044,N_9082);
nand U16355 (N_16355,N_9207,N_8249);
and U16356 (N_16356,N_11815,N_10117);
or U16357 (N_16357,N_11918,N_11244);
nor U16358 (N_16358,N_11687,N_8406);
nor U16359 (N_16359,N_6315,N_7413);
nor U16360 (N_16360,N_6749,N_11159);
and U16361 (N_16361,N_8788,N_8217);
and U16362 (N_16362,N_8791,N_10652);
and U16363 (N_16363,N_8289,N_9481);
nor U16364 (N_16364,N_6555,N_11701);
nor U16365 (N_16365,N_11357,N_8754);
nand U16366 (N_16366,N_7023,N_8064);
nand U16367 (N_16367,N_7597,N_11108);
or U16368 (N_16368,N_10442,N_8753);
xor U16369 (N_16369,N_11456,N_6222);
and U16370 (N_16370,N_7282,N_7196);
or U16371 (N_16371,N_10930,N_10371);
nand U16372 (N_16372,N_7526,N_11448);
nand U16373 (N_16373,N_7916,N_11027);
or U16374 (N_16374,N_7915,N_10094);
and U16375 (N_16375,N_11403,N_6268);
nand U16376 (N_16376,N_11017,N_11897);
nand U16377 (N_16377,N_10035,N_10285);
nand U16378 (N_16378,N_10359,N_9376);
xor U16379 (N_16379,N_11062,N_9751);
or U16380 (N_16380,N_10438,N_6740);
nor U16381 (N_16381,N_10708,N_11839);
nand U16382 (N_16382,N_6364,N_7676);
xnor U16383 (N_16383,N_9647,N_8784);
nand U16384 (N_16384,N_6145,N_9630);
nand U16385 (N_16385,N_10573,N_9931);
and U16386 (N_16386,N_9223,N_9153);
nand U16387 (N_16387,N_8157,N_7594);
nand U16388 (N_16388,N_9800,N_6317);
nand U16389 (N_16389,N_11194,N_6470);
and U16390 (N_16390,N_8627,N_9420);
or U16391 (N_16391,N_9003,N_11605);
nand U16392 (N_16392,N_6203,N_6683);
nor U16393 (N_16393,N_11102,N_9501);
or U16394 (N_16394,N_6265,N_7022);
nand U16395 (N_16395,N_9043,N_8935);
and U16396 (N_16396,N_7963,N_7292);
or U16397 (N_16397,N_9007,N_9209);
xnor U16398 (N_16398,N_8802,N_9115);
nor U16399 (N_16399,N_11866,N_11131);
xor U16400 (N_16400,N_11508,N_7353);
and U16401 (N_16401,N_10821,N_10723);
or U16402 (N_16402,N_9509,N_8063);
or U16403 (N_16403,N_11330,N_7002);
nand U16404 (N_16404,N_6030,N_10204);
xor U16405 (N_16405,N_8543,N_6395);
nand U16406 (N_16406,N_6574,N_10007);
and U16407 (N_16407,N_7814,N_11442);
and U16408 (N_16408,N_7561,N_8997);
nor U16409 (N_16409,N_11263,N_10250);
nand U16410 (N_16410,N_9387,N_11863);
nor U16411 (N_16411,N_9207,N_9500);
or U16412 (N_16412,N_9419,N_6289);
nand U16413 (N_16413,N_11167,N_8768);
or U16414 (N_16414,N_7345,N_10923);
xnor U16415 (N_16415,N_10594,N_9344);
nor U16416 (N_16416,N_10036,N_11923);
and U16417 (N_16417,N_6226,N_8582);
and U16418 (N_16418,N_9173,N_7680);
and U16419 (N_16419,N_10965,N_8623);
nand U16420 (N_16420,N_11118,N_7485);
xor U16421 (N_16421,N_6466,N_6876);
nor U16422 (N_16422,N_10414,N_7428);
or U16423 (N_16423,N_7846,N_6709);
and U16424 (N_16424,N_8276,N_10828);
nand U16425 (N_16425,N_9031,N_8445);
nor U16426 (N_16426,N_8955,N_7384);
nor U16427 (N_16427,N_6687,N_9969);
nor U16428 (N_16428,N_8814,N_6024);
nor U16429 (N_16429,N_7475,N_8992);
and U16430 (N_16430,N_6401,N_8030);
and U16431 (N_16431,N_7836,N_10533);
nor U16432 (N_16432,N_8815,N_6258);
or U16433 (N_16433,N_8127,N_11388);
and U16434 (N_16434,N_7094,N_8646);
or U16435 (N_16435,N_10700,N_6793);
nand U16436 (N_16436,N_6679,N_11312);
nand U16437 (N_16437,N_10779,N_7755);
and U16438 (N_16438,N_9504,N_8870);
nand U16439 (N_16439,N_6726,N_6087);
nor U16440 (N_16440,N_10565,N_11412);
nor U16441 (N_16441,N_11440,N_6353);
nor U16442 (N_16442,N_11046,N_9079);
or U16443 (N_16443,N_11718,N_6386);
and U16444 (N_16444,N_8701,N_11919);
or U16445 (N_16445,N_10328,N_11373);
nor U16446 (N_16446,N_9200,N_10693);
and U16447 (N_16447,N_9834,N_11495);
nor U16448 (N_16448,N_6676,N_7939);
nand U16449 (N_16449,N_11433,N_6973);
nor U16450 (N_16450,N_7808,N_7113);
nor U16451 (N_16451,N_6240,N_10647);
and U16452 (N_16452,N_10325,N_6146);
or U16453 (N_16453,N_6834,N_6166);
nand U16454 (N_16454,N_6686,N_10688);
or U16455 (N_16455,N_6597,N_11769);
and U16456 (N_16456,N_6035,N_6431);
or U16457 (N_16457,N_6704,N_9515);
xnor U16458 (N_16458,N_11791,N_7076);
and U16459 (N_16459,N_8784,N_6817);
nor U16460 (N_16460,N_10385,N_7969);
nor U16461 (N_16461,N_6788,N_10218);
and U16462 (N_16462,N_6254,N_6604);
nor U16463 (N_16463,N_11235,N_10575);
or U16464 (N_16464,N_11190,N_8172);
nand U16465 (N_16465,N_7684,N_11744);
nor U16466 (N_16466,N_8587,N_6792);
or U16467 (N_16467,N_10167,N_9707);
nor U16468 (N_16468,N_7056,N_7553);
and U16469 (N_16469,N_8244,N_9996);
and U16470 (N_16470,N_9131,N_7805);
or U16471 (N_16471,N_8909,N_10746);
xor U16472 (N_16472,N_10910,N_9584);
or U16473 (N_16473,N_6599,N_7870);
and U16474 (N_16474,N_6878,N_9745);
and U16475 (N_16475,N_9234,N_7513);
nand U16476 (N_16476,N_7787,N_10598);
or U16477 (N_16477,N_7967,N_7853);
or U16478 (N_16478,N_7739,N_9805);
xor U16479 (N_16479,N_11956,N_6369);
xor U16480 (N_16480,N_9023,N_10203);
or U16481 (N_16481,N_10103,N_11731);
xnor U16482 (N_16482,N_6090,N_6062);
or U16483 (N_16483,N_11039,N_11166);
nand U16484 (N_16484,N_7218,N_8267);
or U16485 (N_16485,N_8152,N_10862);
xnor U16486 (N_16486,N_9897,N_7402);
xnor U16487 (N_16487,N_7750,N_6993);
nor U16488 (N_16488,N_7129,N_9859);
nand U16489 (N_16489,N_9278,N_10938);
nor U16490 (N_16490,N_8001,N_11413);
nand U16491 (N_16491,N_7878,N_8474);
or U16492 (N_16492,N_8439,N_10307);
or U16493 (N_16493,N_7537,N_9728);
nand U16494 (N_16494,N_6849,N_6244);
xnor U16495 (N_16495,N_9678,N_9046);
nand U16496 (N_16496,N_9605,N_7462);
nand U16497 (N_16497,N_7814,N_9388);
xor U16498 (N_16498,N_8323,N_7140);
or U16499 (N_16499,N_10324,N_9472);
nand U16500 (N_16500,N_11425,N_6145);
and U16501 (N_16501,N_10868,N_9176);
nand U16502 (N_16502,N_9231,N_6644);
and U16503 (N_16503,N_8498,N_11611);
and U16504 (N_16504,N_7720,N_8741);
and U16505 (N_16505,N_9471,N_7296);
and U16506 (N_16506,N_11189,N_10955);
or U16507 (N_16507,N_9161,N_9259);
nor U16508 (N_16508,N_7016,N_10580);
or U16509 (N_16509,N_8224,N_10724);
or U16510 (N_16510,N_8879,N_9683);
nand U16511 (N_16511,N_6053,N_9990);
or U16512 (N_16512,N_7534,N_6808);
nor U16513 (N_16513,N_10616,N_10215);
and U16514 (N_16514,N_9987,N_6284);
or U16515 (N_16515,N_7631,N_6579);
nand U16516 (N_16516,N_9139,N_7323);
nor U16517 (N_16517,N_11192,N_10818);
or U16518 (N_16518,N_7109,N_8983);
or U16519 (N_16519,N_9683,N_9869);
xnor U16520 (N_16520,N_9429,N_11609);
nand U16521 (N_16521,N_9288,N_10220);
nand U16522 (N_16522,N_10732,N_10484);
and U16523 (N_16523,N_11185,N_10230);
nor U16524 (N_16524,N_11925,N_7154);
nor U16525 (N_16525,N_11600,N_11611);
xor U16526 (N_16526,N_6132,N_7107);
nand U16527 (N_16527,N_6351,N_6691);
or U16528 (N_16528,N_11883,N_6682);
nand U16529 (N_16529,N_9417,N_10310);
nor U16530 (N_16530,N_7664,N_8816);
nor U16531 (N_16531,N_9564,N_7129);
nor U16532 (N_16532,N_7108,N_6440);
and U16533 (N_16533,N_11165,N_6038);
nand U16534 (N_16534,N_6277,N_10039);
nand U16535 (N_16535,N_8715,N_11861);
or U16536 (N_16536,N_9704,N_6562);
nor U16537 (N_16537,N_9921,N_10941);
or U16538 (N_16538,N_9639,N_7310);
nor U16539 (N_16539,N_9627,N_9819);
nor U16540 (N_16540,N_8139,N_11322);
and U16541 (N_16541,N_6414,N_11709);
or U16542 (N_16542,N_11654,N_8459);
nor U16543 (N_16543,N_6017,N_9140);
nand U16544 (N_16544,N_11918,N_7510);
nand U16545 (N_16545,N_8141,N_9028);
or U16546 (N_16546,N_8868,N_7123);
nand U16547 (N_16547,N_10869,N_8338);
nor U16548 (N_16548,N_6062,N_9461);
or U16549 (N_16549,N_10244,N_6189);
or U16550 (N_16550,N_7164,N_10664);
or U16551 (N_16551,N_8334,N_6788);
nand U16552 (N_16552,N_9175,N_7314);
and U16553 (N_16553,N_6190,N_8561);
and U16554 (N_16554,N_8680,N_8291);
and U16555 (N_16555,N_7331,N_7459);
and U16556 (N_16556,N_8747,N_7414);
nand U16557 (N_16557,N_7128,N_8308);
nand U16558 (N_16558,N_8089,N_7678);
and U16559 (N_16559,N_6024,N_10302);
xor U16560 (N_16560,N_7836,N_7944);
nor U16561 (N_16561,N_6356,N_11096);
nand U16562 (N_16562,N_9138,N_8445);
xor U16563 (N_16563,N_10301,N_6079);
nand U16564 (N_16564,N_6764,N_8586);
nor U16565 (N_16565,N_7422,N_11684);
xor U16566 (N_16566,N_11893,N_6469);
nor U16567 (N_16567,N_7539,N_6731);
and U16568 (N_16568,N_6398,N_10913);
nor U16569 (N_16569,N_8862,N_7624);
or U16570 (N_16570,N_6917,N_8931);
or U16571 (N_16571,N_6950,N_8968);
and U16572 (N_16572,N_8523,N_9346);
nand U16573 (N_16573,N_11854,N_6257);
xor U16574 (N_16574,N_11090,N_11257);
or U16575 (N_16575,N_7357,N_9607);
nand U16576 (N_16576,N_7611,N_6188);
or U16577 (N_16577,N_10947,N_8319);
or U16578 (N_16578,N_10230,N_6468);
nand U16579 (N_16579,N_11075,N_6459);
nor U16580 (N_16580,N_7161,N_11707);
nor U16581 (N_16581,N_10573,N_6832);
and U16582 (N_16582,N_10274,N_11548);
or U16583 (N_16583,N_9666,N_10635);
xnor U16584 (N_16584,N_10313,N_11109);
and U16585 (N_16585,N_9008,N_7625);
or U16586 (N_16586,N_6090,N_8645);
xor U16587 (N_16587,N_9126,N_9042);
and U16588 (N_16588,N_6943,N_8057);
or U16589 (N_16589,N_7070,N_11909);
and U16590 (N_16590,N_9936,N_6716);
nor U16591 (N_16591,N_8897,N_10496);
and U16592 (N_16592,N_10075,N_7903);
xnor U16593 (N_16593,N_10175,N_6806);
nor U16594 (N_16594,N_10098,N_9245);
nor U16595 (N_16595,N_7070,N_9590);
or U16596 (N_16596,N_9297,N_10901);
nor U16597 (N_16597,N_9843,N_9406);
and U16598 (N_16598,N_9474,N_11929);
xor U16599 (N_16599,N_11127,N_7894);
or U16600 (N_16600,N_8363,N_6593);
nor U16601 (N_16601,N_8234,N_9106);
nand U16602 (N_16602,N_6715,N_8543);
or U16603 (N_16603,N_8149,N_11972);
nor U16604 (N_16604,N_7035,N_7269);
nor U16605 (N_16605,N_8449,N_10032);
xnor U16606 (N_16606,N_7991,N_9998);
and U16607 (N_16607,N_10970,N_9684);
or U16608 (N_16608,N_11047,N_9481);
and U16609 (N_16609,N_9471,N_9405);
nand U16610 (N_16610,N_10666,N_6993);
and U16611 (N_16611,N_8322,N_8166);
nor U16612 (N_16612,N_10572,N_7004);
and U16613 (N_16613,N_10476,N_9515);
nand U16614 (N_16614,N_6333,N_6824);
or U16615 (N_16615,N_6169,N_11289);
nor U16616 (N_16616,N_8195,N_7489);
nand U16617 (N_16617,N_9351,N_7716);
and U16618 (N_16618,N_8764,N_8242);
nor U16619 (N_16619,N_6800,N_11805);
nor U16620 (N_16620,N_7964,N_9868);
xnor U16621 (N_16621,N_6565,N_11914);
nor U16622 (N_16622,N_9938,N_11851);
or U16623 (N_16623,N_10049,N_8797);
and U16624 (N_16624,N_6142,N_11021);
nand U16625 (N_16625,N_7957,N_7308);
or U16626 (N_16626,N_10775,N_10755);
or U16627 (N_16627,N_11072,N_10535);
and U16628 (N_16628,N_6589,N_6357);
and U16629 (N_16629,N_11374,N_10502);
nand U16630 (N_16630,N_8916,N_11309);
or U16631 (N_16631,N_9989,N_7087);
and U16632 (N_16632,N_9450,N_6559);
or U16633 (N_16633,N_6602,N_11141);
and U16634 (N_16634,N_6086,N_6417);
and U16635 (N_16635,N_8419,N_11137);
nor U16636 (N_16636,N_9381,N_6683);
or U16637 (N_16637,N_10285,N_8583);
and U16638 (N_16638,N_10113,N_6736);
nor U16639 (N_16639,N_7691,N_10787);
nand U16640 (N_16640,N_11342,N_8641);
or U16641 (N_16641,N_10416,N_10400);
nand U16642 (N_16642,N_7690,N_6631);
or U16643 (N_16643,N_10572,N_7777);
nor U16644 (N_16644,N_7118,N_7443);
nand U16645 (N_16645,N_8323,N_9510);
nor U16646 (N_16646,N_9814,N_6720);
or U16647 (N_16647,N_9390,N_6794);
nor U16648 (N_16648,N_6419,N_11661);
or U16649 (N_16649,N_7281,N_10585);
xnor U16650 (N_16650,N_9762,N_10864);
nor U16651 (N_16651,N_9925,N_7091);
nand U16652 (N_16652,N_7167,N_7942);
and U16653 (N_16653,N_6844,N_9780);
nor U16654 (N_16654,N_8392,N_11343);
nand U16655 (N_16655,N_10897,N_9027);
nor U16656 (N_16656,N_11810,N_7570);
or U16657 (N_16657,N_10356,N_9251);
nor U16658 (N_16658,N_10406,N_11353);
and U16659 (N_16659,N_9826,N_6320);
or U16660 (N_16660,N_7878,N_10095);
and U16661 (N_16661,N_8044,N_10005);
nor U16662 (N_16662,N_8294,N_9205);
or U16663 (N_16663,N_8080,N_11754);
and U16664 (N_16664,N_7326,N_7399);
nor U16665 (N_16665,N_8156,N_11887);
or U16666 (N_16666,N_10143,N_9179);
nor U16667 (N_16667,N_8412,N_9070);
and U16668 (N_16668,N_8805,N_8184);
nor U16669 (N_16669,N_10548,N_9164);
or U16670 (N_16670,N_9177,N_6461);
nand U16671 (N_16671,N_11663,N_7174);
nor U16672 (N_16672,N_11107,N_9338);
xnor U16673 (N_16673,N_7476,N_6424);
nor U16674 (N_16674,N_8015,N_7927);
and U16675 (N_16675,N_7880,N_8952);
nor U16676 (N_16676,N_11403,N_9586);
nand U16677 (N_16677,N_9343,N_7602);
nand U16678 (N_16678,N_11841,N_10511);
or U16679 (N_16679,N_9407,N_8764);
and U16680 (N_16680,N_7389,N_9438);
nor U16681 (N_16681,N_10376,N_6542);
xor U16682 (N_16682,N_6190,N_11780);
nor U16683 (N_16683,N_8082,N_9539);
nand U16684 (N_16684,N_6202,N_8620);
nor U16685 (N_16685,N_10486,N_7822);
or U16686 (N_16686,N_6117,N_9989);
nand U16687 (N_16687,N_11492,N_7230);
xor U16688 (N_16688,N_11811,N_11873);
xor U16689 (N_16689,N_10941,N_8667);
or U16690 (N_16690,N_6418,N_9804);
and U16691 (N_16691,N_9228,N_10602);
nor U16692 (N_16692,N_8023,N_7102);
nor U16693 (N_16693,N_9082,N_7547);
and U16694 (N_16694,N_7329,N_6218);
nor U16695 (N_16695,N_11717,N_9354);
nand U16696 (N_16696,N_9105,N_9433);
and U16697 (N_16697,N_8014,N_7111);
or U16698 (N_16698,N_9569,N_10311);
nor U16699 (N_16699,N_9342,N_7392);
nand U16700 (N_16700,N_9458,N_7127);
nor U16701 (N_16701,N_10624,N_7115);
xor U16702 (N_16702,N_11480,N_9503);
nor U16703 (N_16703,N_11863,N_8691);
or U16704 (N_16704,N_6248,N_9910);
nor U16705 (N_16705,N_7140,N_6383);
or U16706 (N_16706,N_6416,N_10350);
and U16707 (N_16707,N_9503,N_10701);
and U16708 (N_16708,N_6892,N_6320);
and U16709 (N_16709,N_10224,N_6025);
and U16710 (N_16710,N_7109,N_10286);
nor U16711 (N_16711,N_11128,N_6195);
and U16712 (N_16712,N_11163,N_8278);
nand U16713 (N_16713,N_8597,N_7501);
nor U16714 (N_16714,N_11153,N_11845);
nor U16715 (N_16715,N_11694,N_11476);
nor U16716 (N_16716,N_6176,N_11321);
nor U16717 (N_16717,N_8543,N_10639);
nand U16718 (N_16718,N_6823,N_6028);
nor U16719 (N_16719,N_7632,N_7788);
nand U16720 (N_16720,N_6907,N_10281);
nand U16721 (N_16721,N_10840,N_6273);
nor U16722 (N_16722,N_7433,N_7890);
and U16723 (N_16723,N_6876,N_9741);
nor U16724 (N_16724,N_9052,N_6875);
nor U16725 (N_16725,N_7211,N_8294);
nand U16726 (N_16726,N_11799,N_9307);
nor U16727 (N_16727,N_6133,N_6096);
and U16728 (N_16728,N_8447,N_6124);
and U16729 (N_16729,N_7965,N_7981);
xor U16730 (N_16730,N_8682,N_10292);
nand U16731 (N_16731,N_6945,N_6284);
nor U16732 (N_16732,N_8111,N_9277);
nand U16733 (N_16733,N_10819,N_8910);
nor U16734 (N_16734,N_10306,N_11084);
and U16735 (N_16735,N_9974,N_6508);
nand U16736 (N_16736,N_6019,N_6742);
and U16737 (N_16737,N_9693,N_9567);
nand U16738 (N_16738,N_9141,N_11187);
nand U16739 (N_16739,N_6714,N_6358);
nor U16740 (N_16740,N_9970,N_11379);
nor U16741 (N_16741,N_7008,N_6054);
nor U16742 (N_16742,N_7954,N_10306);
or U16743 (N_16743,N_8585,N_11824);
or U16744 (N_16744,N_8010,N_11039);
nor U16745 (N_16745,N_8929,N_7718);
or U16746 (N_16746,N_10706,N_11413);
xor U16747 (N_16747,N_7526,N_9554);
or U16748 (N_16748,N_11022,N_8345);
and U16749 (N_16749,N_10100,N_11774);
nor U16750 (N_16750,N_6138,N_6915);
nand U16751 (N_16751,N_10771,N_10919);
nor U16752 (N_16752,N_11885,N_6162);
or U16753 (N_16753,N_8880,N_9969);
nand U16754 (N_16754,N_6299,N_11071);
nand U16755 (N_16755,N_11281,N_8452);
nor U16756 (N_16756,N_10399,N_7106);
nand U16757 (N_16757,N_9361,N_11993);
nor U16758 (N_16758,N_11693,N_7912);
nand U16759 (N_16759,N_7781,N_8425);
nor U16760 (N_16760,N_9178,N_8168);
nand U16761 (N_16761,N_7337,N_9458);
nand U16762 (N_16762,N_9152,N_9218);
nand U16763 (N_16763,N_7487,N_11464);
xnor U16764 (N_16764,N_9313,N_9262);
and U16765 (N_16765,N_6228,N_10720);
nor U16766 (N_16766,N_7329,N_11932);
and U16767 (N_16767,N_10517,N_9315);
nor U16768 (N_16768,N_8164,N_6758);
or U16769 (N_16769,N_7627,N_8334);
nand U16770 (N_16770,N_6630,N_7831);
and U16771 (N_16771,N_9482,N_10210);
xnor U16772 (N_16772,N_9164,N_10639);
or U16773 (N_16773,N_6190,N_10277);
nand U16774 (N_16774,N_7529,N_7930);
and U16775 (N_16775,N_7826,N_6085);
xor U16776 (N_16776,N_6878,N_11209);
nor U16777 (N_16777,N_6875,N_10230);
xor U16778 (N_16778,N_7524,N_7884);
and U16779 (N_16779,N_7531,N_7183);
nor U16780 (N_16780,N_11646,N_9067);
nor U16781 (N_16781,N_11562,N_9263);
or U16782 (N_16782,N_7110,N_9097);
nand U16783 (N_16783,N_9929,N_10680);
or U16784 (N_16784,N_9381,N_10191);
and U16785 (N_16785,N_10489,N_8489);
xnor U16786 (N_16786,N_9137,N_10675);
xor U16787 (N_16787,N_7488,N_9789);
nor U16788 (N_16788,N_7843,N_9189);
nand U16789 (N_16789,N_7074,N_6807);
and U16790 (N_16790,N_6698,N_7198);
nor U16791 (N_16791,N_8594,N_10479);
nor U16792 (N_16792,N_11081,N_11793);
nor U16793 (N_16793,N_8916,N_7598);
xnor U16794 (N_16794,N_6944,N_9853);
nor U16795 (N_16795,N_10434,N_8692);
or U16796 (N_16796,N_11316,N_8823);
nand U16797 (N_16797,N_11783,N_10074);
and U16798 (N_16798,N_8039,N_9727);
xnor U16799 (N_16799,N_9437,N_9662);
nor U16800 (N_16800,N_9896,N_7376);
or U16801 (N_16801,N_9289,N_11453);
nor U16802 (N_16802,N_11906,N_9317);
nor U16803 (N_16803,N_9133,N_9345);
nor U16804 (N_16804,N_7243,N_8518);
nand U16805 (N_16805,N_11662,N_9957);
and U16806 (N_16806,N_8736,N_8011);
xnor U16807 (N_16807,N_10346,N_11865);
nand U16808 (N_16808,N_10250,N_6816);
nand U16809 (N_16809,N_10314,N_10031);
xor U16810 (N_16810,N_10517,N_11964);
nor U16811 (N_16811,N_7974,N_9100);
or U16812 (N_16812,N_11607,N_7525);
and U16813 (N_16813,N_10357,N_8774);
nand U16814 (N_16814,N_6805,N_7800);
nor U16815 (N_16815,N_11012,N_6516);
nand U16816 (N_16816,N_11037,N_9416);
nand U16817 (N_16817,N_8964,N_9371);
or U16818 (N_16818,N_6520,N_7145);
xor U16819 (N_16819,N_9127,N_7622);
xnor U16820 (N_16820,N_7809,N_7527);
nor U16821 (N_16821,N_6905,N_11958);
nor U16822 (N_16822,N_11947,N_11754);
nand U16823 (N_16823,N_8173,N_11176);
and U16824 (N_16824,N_11871,N_9852);
nor U16825 (N_16825,N_8191,N_8024);
nor U16826 (N_16826,N_7851,N_7999);
nor U16827 (N_16827,N_7268,N_11821);
nor U16828 (N_16828,N_7719,N_6279);
nor U16829 (N_16829,N_7259,N_11813);
nor U16830 (N_16830,N_11053,N_10905);
and U16831 (N_16831,N_7928,N_9337);
or U16832 (N_16832,N_10320,N_9614);
or U16833 (N_16833,N_10547,N_11141);
nand U16834 (N_16834,N_7702,N_11476);
or U16835 (N_16835,N_10373,N_9038);
nand U16836 (N_16836,N_6456,N_6632);
nor U16837 (N_16837,N_8754,N_10566);
or U16838 (N_16838,N_6887,N_10906);
nand U16839 (N_16839,N_9728,N_6438);
nor U16840 (N_16840,N_10066,N_6116);
and U16841 (N_16841,N_10506,N_10787);
nor U16842 (N_16842,N_10865,N_7156);
or U16843 (N_16843,N_7215,N_7207);
nor U16844 (N_16844,N_8123,N_11138);
and U16845 (N_16845,N_7339,N_11318);
nand U16846 (N_16846,N_6821,N_7615);
nand U16847 (N_16847,N_10832,N_6709);
nor U16848 (N_16848,N_9190,N_11709);
xor U16849 (N_16849,N_11530,N_8732);
nor U16850 (N_16850,N_7967,N_6225);
or U16851 (N_16851,N_11261,N_11664);
or U16852 (N_16852,N_7383,N_7617);
nor U16853 (N_16853,N_8793,N_6629);
or U16854 (N_16854,N_10769,N_6215);
nand U16855 (N_16855,N_10683,N_8886);
nand U16856 (N_16856,N_8944,N_8985);
nor U16857 (N_16857,N_11714,N_8285);
and U16858 (N_16858,N_11086,N_8745);
nor U16859 (N_16859,N_9055,N_6069);
or U16860 (N_16860,N_7381,N_6524);
nand U16861 (N_16861,N_10887,N_7427);
nand U16862 (N_16862,N_11227,N_6291);
or U16863 (N_16863,N_9848,N_7417);
or U16864 (N_16864,N_8995,N_6914);
xor U16865 (N_16865,N_6665,N_10905);
nor U16866 (N_16866,N_9916,N_11999);
and U16867 (N_16867,N_7747,N_6903);
nor U16868 (N_16868,N_9203,N_10703);
xor U16869 (N_16869,N_9605,N_10482);
or U16870 (N_16870,N_9054,N_7712);
xor U16871 (N_16871,N_9124,N_8820);
nor U16872 (N_16872,N_10133,N_11806);
nor U16873 (N_16873,N_11602,N_7492);
nor U16874 (N_16874,N_11501,N_9271);
nor U16875 (N_16875,N_9838,N_6028);
nor U16876 (N_16876,N_6778,N_9589);
nand U16877 (N_16877,N_11123,N_9384);
nor U16878 (N_16878,N_7346,N_7331);
and U16879 (N_16879,N_11289,N_10541);
nor U16880 (N_16880,N_11105,N_8777);
nand U16881 (N_16881,N_10018,N_8715);
nand U16882 (N_16882,N_6310,N_6816);
xnor U16883 (N_16883,N_10403,N_7449);
and U16884 (N_16884,N_10424,N_6829);
and U16885 (N_16885,N_10955,N_7355);
nor U16886 (N_16886,N_7515,N_6225);
or U16887 (N_16887,N_11943,N_11251);
and U16888 (N_16888,N_9736,N_11951);
or U16889 (N_16889,N_7720,N_7747);
or U16890 (N_16890,N_7971,N_9943);
or U16891 (N_16891,N_10988,N_7062);
xor U16892 (N_16892,N_6586,N_6019);
and U16893 (N_16893,N_7701,N_11349);
nor U16894 (N_16894,N_7978,N_8666);
or U16895 (N_16895,N_6784,N_10946);
and U16896 (N_16896,N_11243,N_10582);
or U16897 (N_16897,N_11203,N_11595);
or U16898 (N_16898,N_6091,N_10799);
or U16899 (N_16899,N_6115,N_6001);
or U16900 (N_16900,N_8928,N_7529);
nand U16901 (N_16901,N_10027,N_10966);
nand U16902 (N_16902,N_11382,N_9077);
nand U16903 (N_16903,N_8113,N_8213);
nor U16904 (N_16904,N_9851,N_10211);
nor U16905 (N_16905,N_8493,N_11922);
and U16906 (N_16906,N_6592,N_7674);
nand U16907 (N_16907,N_10531,N_6034);
nand U16908 (N_16908,N_8553,N_8734);
nand U16909 (N_16909,N_11336,N_8859);
xnor U16910 (N_16910,N_10185,N_9457);
nand U16911 (N_16911,N_8640,N_6691);
or U16912 (N_16912,N_11325,N_6286);
nor U16913 (N_16913,N_9267,N_9874);
nand U16914 (N_16914,N_6535,N_7088);
xnor U16915 (N_16915,N_7615,N_9092);
nor U16916 (N_16916,N_10261,N_10737);
and U16917 (N_16917,N_7843,N_7101);
nand U16918 (N_16918,N_6523,N_11130);
and U16919 (N_16919,N_10172,N_6421);
xnor U16920 (N_16920,N_10222,N_10509);
nand U16921 (N_16921,N_6762,N_10539);
xor U16922 (N_16922,N_9461,N_8653);
nand U16923 (N_16923,N_10123,N_9683);
and U16924 (N_16924,N_7869,N_7451);
nand U16925 (N_16925,N_9115,N_11670);
or U16926 (N_16926,N_9995,N_8546);
nor U16927 (N_16927,N_9967,N_8760);
or U16928 (N_16928,N_10705,N_11009);
nor U16929 (N_16929,N_10350,N_11235);
nand U16930 (N_16930,N_9654,N_8151);
nor U16931 (N_16931,N_9379,N_8226);
nand U16932 (N_16932,N_6114,N_7056);
or U16933 (N_16933,N_8417,N_11413);
nor U16934 (N_16934,N_7848,N_9075);
and U16935 (N_16935,N_11216,N_10123);
xnor U16936 (N_16936,N_6811,N_10003);
nor U16937 (N_16937,N_10005,N_9343);
nor U16938 (N_16938,N_10915,N_6187);
nand U16939 (N_16939,N_8402,N_10646);
or U16940 (N_16940,N_11940,N_10352);
nor U16941 (N_16941,N_10864,N_9562);
xnor U16942 (N_16942,N_7551,N_7602);
nor U16943 (N_16943,N_7839,N_11742);
and U16944 (N_16944,N_7038,N_9708);
nand U16945 (N_16945,N_8998,N_6050);
or U16946 (N_16946,N_9216,N_11626);
nor U16947 (N_16947,N_11095,N_10035);
nand U16948 (N_16948,N_7249,N_7305);
or U16949 (N_16949,N_9822,N_7042);
or U16950 (N_16950,N_6400,N_6410);
or U16951 (N_16951,N_11787,N_9040);
nor U16952 (N_16952,N_9908,N_11011);
nor U16953 (N_16953,N_6124,N_8589);
nand U16954 (N_16954,N_9287,N_6216);
or U16955 (N_16955,N_6895,N_11319);
and U16956 (N_16956,N_7275,N_8210);
or U16957 (N_16957,N_10773,N_7063);
xor U16958 (N_16958,N_7341,N_9408);
nand U16959 (N_16959,N_8569,N_10918);
and U16960 (N_16960,N_10254,N_8456);
nand U16961 (N_16961,N_10628,N_6748);
and U16962 (N_16962,N_8974,N_10805);
or U16963 (N_16963,N_9716,N_11552);
nand U16964 (N_16964,N_10733,N_9376);
nand U16965 (N_16965,N_7153,N_10295);
xnor U16966 (N_16966,N_10924,N_10699);
or U16967 (N_16967,N_11725,N_11560);
or U16968 (N_16968,N_9597,N_11832);
and U16969 (N_16969,N_9937,N_11713);
nand U16970 (N_16970,N_11792,N_7348);
or U16971 (N_16971,N_9931,N_6402);
nor U16972 (N_16972,N_9334,N_10842);
or U16973 (N_16973,N_7865,N_7193);
or U16974 (N_16974,N_9024,N_8460);
or U16975 (N_16975,N_9210,N_9726);
nand U16976 (N_16976,N_7463,N_6761);
nand U16977 (N_16977,N_9561,N_9081);
and U16978 (N_16978,N_7955,N_6806);
and U16979 (N_16979,N_11200,N_6894);
nand U16980 (N_16980,N_8949,N_10932);
nand U16981 (N_16981,N_8379,N_7263);
or U16982 (N_16982,N_9185,N_7407);
and U16983 (N_16983,N_10431,N_11332);
and U16984 (N_16984,N_6418,N_9036);
xnor U16985 (N_16985,N_9439,N_10980);
or U16986 (N_16986,N_7465,N_9005);
or U16987 (N_16987,N_9301,N_6659);
nand U16988 (N_16988,N_9734,N_10623);
nor U16989 (N_16989,N_7959,N_11990);
or U16990 (N_16990,N_6432,N_10775);
nor U16991 (N_16991,N_10152,N_10784);
or U16992 (N_16992,N_10934,N_7417);
and U16993 (N_16993,N_10388,N_8849);
xor U16994 (N_16994,N_8288,N_11435);
nand U16995 (N_16995,N_7811,N_10679);
and U16996 (N_16996,N_11222,N_11777);
nor U16997 (N_16997,N_9557,N_6787);
nor U16998 (N_16998,N_8593,N_6549);
and U16999 (N_16999,N_8023,N_9479);
or U17000 (N_17000,N_10003,N_11371);
or U17001 (N_17001,N_9187,N_9338);
and U17002 (N_17002,N_10407,N_6349);
or U17003 (N_17003,N_7137,N_9795);
nor U17004 (N_17004,N_10326,N_11194);
nor U17005 (N_17005,N_8908,N_8826);
nand U17006 (N_17006,N_8964,N_9355);
or U17007 (N_17007,N_10888,N_7458);
nand U17008 (N_17008,N_6363,N_8718);
nand U17009 (N_17009,N_9164,N_9791);
or U17010 (N_17010,N_9093,N_8295);
nor U17011 (N_17011,N_7753,N_10907);
nand U17012 (N_17012,N_8179,N_9359);
or U17013 (N_17013,N_11377,N_10107);
nand U17014 (N_17014,N_7382,N_9767);
nor U17015 (N_17015,N_7891,N_9018);
or U17016 (N_17016,N_6823,N_10714);
nor U17017 (N_17017,N_6026,N_11355);
nor U17018 (N_17018,N_11286,N_8673);
nor U17019 (N_17019,N_10373,N_6260);
nor U17020 (N_17020,N_8808,N_8513);
and U17021 (N_17021,N_11130,N_11661);
nor U17022 (N_17022,N_7883,N_8766);
nor U17023 (N_17023,N_7776,N_7473);
xnor U17024 (N_17024,N_9403,N_6379);
and U17025 (N_17025,N_6619,N_8791);
nand U17026 (N_17026,N_10997,N_7175);
xor U17027 (N_17027,N_9437,N_11174);
and U17028 (N_17028,N_11885,N_8349);
xor U17029 (N_17029,N_8393,N_10531);
nor U17030 (N_17030,N_6825,N_8342);
nand U17031 (N_17031,N_11198,N_11253);
or U17032 (N_17032,N_10538,N_8094);
xnor U17033 (N_17033,N_7468,N_7492);
xor U17034 (N_17034,N_6421,N_10017);
nor U17035 (N_17035,N_11455,N_7228);
nand U17036 (N_17036,N_8358,N_8196);
or U17037 (N_17037,N_11274,N_7289);
nor U17038 (N_17038,N_11170,N_8515);
nor U17039 (N_17039,N_10111,N_6801);
or U17040 (N_17040,N_11232,N_9152);
nand U17041 (N_17041,N_8307,N_10777);
and U17042 (N_17042,N_11705,N_8183);
nor U17043 (N_17043,N_6151,N_10826);
nand U17044 (N_17044,N_7008,N_9136);
or U17045 (N_17045,N_11669,N_6728);
or U17046 (N_17046,N_11746,N_8951);
and U17047 (N_17047,N_10494,N_7704);
nand U17048 (N_17048,N_7872,N_11162);
or U17049 (N_17049,N_7433,N_6288);
nor U17050 (N_17050,N_11243,N_8880);
nor U17051 (N_17051,N_10427,N_9443);
nor U17052 (N_17052,N_8894,N_11002);
and U17053 (N_17053,N_9302,N_6068);
or U17054 (N_17054,N_9320,N_11217);
or U17055 (N_17055,N_7170,N_9517);
or U17056 (N_17056,N_10358,N_11044);
nand U17057 (N_17057,N_10001,N_8035);
xor U17058 (N_17058,N_10520,N_7551);
nand U17059 (N_17059,N_7780,N_6457);
or U17060 (N_17060,N_7402,N_10527);
and U17061 (N_17061,N_6076,N_8212);
and U17062 (N_17062,N_8998,N_11797);
nor U17063 (N_17063,N_7612,N_6596);
nor U17064 (N_17064,N_7632,N_7027);
and U17065 (N_17065,N_6294,N_8397);
and U17066 (N_17066,N_6447,N_10271);
nand U17067 (N_17067,N_6019,N_6061);
or U17068 (N_17068,N_6099,N_11404);
and U17069 (N_17069,N_9094,N_8458);
or U17070 (N_17070,N_6239,N_10992);
xor U17071 (N_17071,N_6908,N_6635);
and U17072 (N_17072,N_10202,N_6189);
or U17073 (N_17073,N_6618,N_10349);
or U17074 (N_17074,N_11085,N_8292);
and U17075 (N_17075,N_11847,N_10255);
nand U17076 (N_17076,N_7218,N_8518);
xnor U17077 (N_17077,N_7918,N_10516);
nor U17078 (N_17078,N_9270,N_6275);
and U17079 (N_17079,N_6301,N_6296);
nor U17080 (N_17080,N_6281,N_8652);
nand U17081 (N_17081,N_11561,N_7545);
nand U17082 (N_17082,N_10541,N_8508);
or U17083 (N_17083,N_10105,N_6152);
nand U17084 (N_17084,N_6337,N_9031);
nor U17085 (N_17085,N_10423,N_7211);
and U17086 (N_17086,N_11898,N_6257);
xnor U17087 (N_17087,N_10673,N_6645);
nor U17088 (N_17088,N_8146,N_9872);
nand U17089 (N_17089,N_10040,N_7329);
xnor U17090 (N_17090,N_8709,N_10811);
xor U17091 (N_17091,N_10370,N_10569);
or U17092 (N_17092,N_7166,N_11987);
and U17093 (N_17093,N_6176,N_8337);
or U17094 (N_17094,N_9915,N_10577);
and U17095 (N_17095,N_10785,N_9963);
or U17096 (N_17096,N_7314,N_9017);
nand U17097 (N_17097,N_8773,N_8866);
and U17098 (N_17098,N_11175,N_8496);
or U17099 (N_17099,N_7701,N_8219);
nor U17100 (N_17100,N_6988,N_10236);
nor U17101 (N_17101,N_6672,N_8332);
nor U17102 (N_17102,N_10255,N_9396);
and U17103 (N_17103,N_6034,N_9813);
or U17104 (N_17104,N_6391,N_8577);
nand U17105 (N_17105,N_10628,N_8537);
xor U17106 (N_17106,N_9943,N_9270);
and U17107 (N_17107,N_9040,N_10793);
nand U17108 (N_17108,N_11706,N_11910);
nand U17109 (N_17109,N_8892,N_6080);
nor U17110 (N_17110,N_7831,N_9206);
and U17111 (N_17111,N_6302,N_6257);
nor U17112 (N_17112,N_8355,N_6482);
nor U17113 (N_17113,N_7449,N_10245);
nand U17114 (N_17114,N_9309,N_10790);
nand U17115 (N_17115,N_11328,N_7259);
or U17116 (N_17116,N_9345,N_7927);
or U17117 (N_17117,N_7827,N_10796);
and U17118 (N_17118,N_6857,N_8487);
nand U17119 (N_17119,N_10930,N_8492);
xor U17120 (N_17120,N_9929,N_11737);
and U17121 (N_17121,N_7592,N_8907);
nor U17122 (N_17122,N_11820,N_11984);
nor U17123 (N_17123,N_10426,N_7859);
nand U17124 (N_17124,N_6040,N_11138);
nand U17125 (N_17125,N_10607,N_11901);
or U17126 (N_17126,N_10337,N_8738);
nor U17127 (N_17127,N_11250,N_7388);
or U17128 (N_17128,N_10962,N_9289);
and U17129 (N_17129,N_10306,N_7437);
nor U17130 (N_17130,N_6200,N_9532);
or U17131 (N_17131,N_10240,N_10659);
or U17132 (N_17132,N_10305,N_10096);
and U17133 (N_17133,N_8191,N_10463);
and U17134 (N_17134,N_6080,N_10675);
nor U17135 (N_17135,N_7253,N_9426);
nor U17136 (N_17136,N_11348,N_6379);
nand U17137 (N_17137,N_11839,N_9860);
or U17138 (N_17138,N_10456,N_6699);
nand U17139 (N_17139,N_6634,N_11194);
nor U17140 (N_17140,N_9725,N_8770);
and U17141 (N_17141,N_7908,N_11109);
nor U17142 (N_17142,N_8821,N_9768);
or U17143 (N_17143,N_11269,N_10946);
or U17144 (N_17144,N_8464,N_10281);
or U17145 (N_17145,N_9585,N_6990);
and U17146 (N_17146,N_7636,N_9525);
and U17147 (N_17147,N_11651,N_6327);
nand U17148 (N_17148,N_9773,N_10265);
and U17149 (N_17149,N_9126,N_9798);
nand U17150 (N_17150,N_7650,N_10440);
xor U17151 (N_17151,N_9092,N_10053);
xor U17152 (N_17152,N_9381,N_6022);
nand U17153 (N_17153,N_8880,N_11319);
nand U17154 (N_17154,N_8297,N_9223);
and U17155 (N_17155,N_10037,N_6045);
or U17156 (N_17156,N_7067,N_7450);
nand U17157 (N_17157,N_8368,N_11914);
nor U17158 (N_17158,N_8186,N_9150);
and U17159 (N_17159,N_10013,N_10781);
or U17160 (N_17160,N_7499,N_11457);
nor U17161 (N_17161,N_11374,N_7807);
and U17162 (N_17162,N_9736,N_6230);
or U17163 (N_17163,N_10543,N_11523);
and U17164 (N_17164,N_10639,N_11282);
and U17165 (N_17165,N_6085,N_11966);
or U17166 (N_17166,N_6385,N_9121);
or U17167 (N_17167,N_8453,N_7821);
and U17168 (N_17168,N_9328,N_9104);
nand U17169 (N_17169,N_9514,N_7689);
nor U17170 (N_17170,N_10030,N_9472);
nor U17171 (N_17171,N_11000,N_11733);
or U17172 (N_17172,N_11584,N_11544);
nand U17173 (N_17173,N_6157,N_11775);
nor U17174 (N_17174,N_7358,N_11859);
nor U17175 (N_17175,N_7441,N_9556);
nor U17176 (N_17176,N_6929,N_8525);
and U17177 (N_17177,N_8941,N_7671);
or U17178 (N_17178,N_6442,N_7775);
nor U17179 (N_17179,N_9660,N_9784);
nand U17180 (N_17180,N_6479,N_8124);
nand U17181 (N_17181,N_11021,N_7807);
nand U17182 (N_17182,N_11241,N_10641);
xor U17183 (N_17183,N_9213,N_8892);
nand U17184 (N_17184,N_11718,N_8499);
and U17185 (N_17185,N_7075,N_9690);
nor U17186 (N_17186,N_6389,N_10115);
and U17187 (N_17187,N_10423,N_10020);
nand U17188 (N_17188,N_9717,N_11215);
nand U17189 (N_17189,N_8251,N_7644);
nand U17190 (N_17190,N_8168,N_8579);
nor U17191 (N_17191,N_7693,N_11209);
or U17192 (N_17192,N_11361,N_7034);
or U17193 (N_17193,N_8967,N_9878);
or U17194 (N_17194,N_7575,N_9522);
or U17195 (N_17195,N_9329,N_9486);
or U17196 (N_17196,N_8724,N_9497);
and U17197 (N_17197,N_11427,N_7014);
or U17198 (N_17198,N_7378,N_6927);
nor U17199 (N_17199,N_9164,N_7610);
nor U17200 (N_17200,N_10375,N_6814);
and U17201 (N_17201,N_9031,N_7544);
xor U17202 (N_17202,N_10653,N_11192);
or U17203 (N_17203,N_8281,N_6343);
nor U17204 (N_17204,N_7019,N_8457);
or U17205 (N_17205,N_6404,N_11563);
nor U17206 (N_17206,N_10276,N_7061);
or U17207 (N_17207,N_7483,N_8209);
and U17208 (N_17208,N_9492,N_11485);
nand U17209 (N_17209,N_11502,N_10408);
nor U17210 (N_17210,N_7467,N_8767);
nor U17211 (N_17211,N_7078,N_10429);
and U17212 (N_17212,N_6529,N_11072);
or U17213 (N_17213,N_8212,N_6105);
nand U17214 (N_17214,N_10252,N_9204);
or U17215 (N_17215,N_7379,N_11309);
or U17216 (N_17216,N_10407,N_10003);
and U17217 (N_17217,N_6679,N_8706);
and U17218 (N_17218,N_9330,N_9090);
or U17219 (N_17219,N_6229,N_9737);
and U17220 (N_17220,N_9303,N_10798);
or U17221 (N_17221,N_6059,N_9679);
and U17222 (N_17222,N_6108,N_11806);
nor U17223 (N_17223,N_10275,N_7275);
or U17224 (N_17224,N_7397,N_7351);
and U17225 (N_17225,N_6418,N_10765);
nand U17226 (N_17226,N_9203,N_9838);
nand U17227 (N_17227,N_7318,N_7915);
nand U17228 (N_17228,N_11292,N_6503);
or U17229 (N_17229,N_6643,N_7629);
nand U17230 (N_17230,N_6456,N_11053);
nor U17231 (N_17231,N_6142,N_7874);
nor U17232 (N_17232,N_6568,N_7757);
nor U17233 (N_17233,N_9545,N_9093);
nand U17234 (N_17234,N_9985,N_7332);
xnor U17235 (N_17235,N_6664,N_10893);
and U17236 (N_17236,N_7501,N_6963);
nor U17237 (N_17237,N_7296,N_6585);
nor U17238 (N_17238,N_11784,N_9384);
nand U17239 (N_17239,N_9344,N_11826);
and U17240 (N_17240,N_6820,N_6524);
nand U17241 (N_17241,N_6274,N_11602);
nand U17242 (N_17242,N_8238,N_11158);
xnor U17243 (N_17243,N_8051,N_11231);
nand U17244 (N_17244,N_11850,N_9813);
nand U17245 (N_17245,N_7882,N_8584);
or U17246 (N_17246,N_8468,N_7462);
nand U17247 (N_17247,N_8171,N_9985);
or U17248 (N_17248,N_7736,N_8929);
xnor U17249 (N_17249,N_9577,N_6825);
nor U17250 (N_17250,N_6692,N_10045);
or U17251 (N_17251,N_8759,N_10406);
or U17252 (N_17252,N_8998,N_11057);
or U17253 (N_17253,N_6485,N_8687);
or U17254 (N_17254,N_11729,N_8085);
nand U17255 (N_17255,N_8448,N_10638);
or U17256 (N_17256,N_11828,N_9818);
nand U17257 (N_17257,N_7777,N_11474);
xor U17258 (N_17258,N_6745,N_6617);
xnor U17259 (N_17259,N_7761,N_8102);
xnor U17260 (N_17260,N_9477,N_6480);
and U17261 (N_17261,N_7581,N_9898);
or U17262 (N_17262,N_11516,N_10860);
nand U17263 (N_17263,N_7889,N_7820);
nor U17264 (N_17264,N_11314,N_10335);
or U17265 (N_17265,N_10484,N_9903);
nand U17266 (N_17266,N_7910,N_8149);
xor U17267 (N_17267,N_8944,N_9723);
and U17268 (N_17268,N_10258,N_9686);
nand U17269 (N_17269,N_7648,N_8355);
nand U17270 (N_17270,N_7564,N_6354);
or U17271 (N_17271,N_7899,N_6142);
nor U17272 (N_17272,N_6264,N_7050);
xnor U17273 (N_17273,N_11614,N_9145);
and U17274 (N_17274,N_10301,N_8305);
nand U17275 (N_17275,N_9436,N_8985);
and U17276 (N_17276,N_9100,N_11649);
nor U17277 (N_17277,N_11568,N_11862);
or U17278 (N_17278,N_11283,N_11323);
nand U17279 (N_17279,N_6807,N_9910);
or U17280 (N_17280,N_7068,N_8740);
nand U17281 (N_17281,N_7081,N_8097);
xnor U17282 (N_17282,N_11420,N_6929);
nand U17283 (N_17283,N_10650,N_8519);
or U17284 (N_17284,N_8506,N_6121);
and U17285 (N_17285,N_10700,N_10485);
nor U17286 (N_17286,N_10570,N_7483);
and U17287 (N_17287,N_11837,N_6476);
and U17288 (N_17288,N_6276,N_9997);
nor U17289 (N_17289,N_11299,N_7969);
nor U17290 (N_17290,N_9802,N_9189);
and U17291 (N_17291,N_10309,N_7373);
nand U17292 (N_17292,N_11385,N_10721);
xnor U17293 (N_17293,N_10612,N_7614);
nor U17294 (N_17294,N_11421,N_9433);
and U17295 (N_17295,N_6977,N_10202);
nor U17296 (N_17296,N_8780,N_10599);
or U17297 (N_17297,N_7540,N_9006);
or U17298 (N_17298,N_8151,N_8985);
nand U17299 (N_17299,N_9129,N_11867);
nor U17300 (N_17300,N_6743,N_7379);
nor U17301 (N_17301,N_8952,N_10033);
or U17302 (N_17302,N_7796,N_6439);
nor U17303 (N_17303,N_9073,N_9394);
xnor U17304 (N_17304,N_6479,N_6198);
and U17305 (N_17305,N_9590,N_9436);
or U17306 (N_17306,N_11468,N_11783);
nand U17307 (N_17307,N_6674,N_8988);
nor U17308 (N_17308,N_10980,N_9136);
nand U17309 (N_17309,N_7555,N_7017);
nand U17310 (N_17310,N_10090,N_9913);
nor U17311 (N_17311,N_10209,N_7382);
or U17312 (N_17312,N_6411,N_8887);
xor U17313 (N_17313,N_6116,N_6702);
and U17314 (N_17314,N_7056,N_6835);
nand U17315 (N_17315,N_7150,N_9458);
nand U17316 (N_17316,N_8236,N_7039);
nand U17317 (N_17317,N_6859,N_7771);
or U17318 (N_17318,N_11899,N_11873);
nand U17319 (N_17319,N_9054,N_8298);
nor U17320 (N_17320,N_8795,N_8721);
nand U17321 (N_17321,N_7323,N_10236);
nand U17322 (N_17322,N_7453,N_9122);
nor U17323 (N_17323,N_9176,N_7682);
nor U17324 (N_17324,N_6349,N_10801);
nand U17325 (N_17325,N_6745,N_6297);
nor U17326 (N_17326,N_7163,N_10522);
nor U17327 (N_17327,N_10067,N_10748);
and U17328 (N_17328,N_7307,N_9371);
and U17329 (N_17329,N_6345,N_7570);
and U17330 (N_17330,N_7924,N_7339);
or U17331 (N_17331,N_8605,N_7268);
or U17332 (N_17332,N_9921,N_8633);
xnor U17333 (N_17333,N_8224,N_7275);
or U17334 (N_17334,N_8803,N_10673);
nand U17335 (N_17335,N_8697,N_6546);
or U17336 (N_17336,N_8631,N_6202);
or U17337 (N_17337,N_7156,N_8087);
and U17338 (N_17338,N_6838,N_8035);
or U17339 (N_17339,N_10352,N_8626);
nor U17340 (N_17340,N_7905,N_7077);
nor U17341 (N_17341,N_11660,N_10712);
nand U17342 (N_17342,N_8684,N_7417);
xnor U17343 (N_17343,N_6323,N_6760);
nor U17344 (N_17344,N_11912,N_9939);
nand U17345 (N_17345,N_10020,N_6355);
and U17346 (N_17346,N_11973,N_7979);
nor U17347 (N_17347,N_10834,N_10751);
nor U17348 (N_17348,N_10890,N_8232);
xnor U17349 (N_17349,N_7882,N_6606);
nor U17350 (N_17350,N_10312,N_6269);
or U17351 (N_17351,N_10067,N_9686);
nand U17352 (N_17352,N_8059,N_8276);
nor U17353 (N_17353,N_7443,N_7608);
nand U17354 (N_17354,N_11133,N_10754);
nor U17355 (N_17355,N_11842,N_11229);
and U17356 (N_17356,N_10924,N_11698);
and U17357 (N_17357,N_6926,N_7104);
xnor U17358 (N_17358,N_8489,N_6691);
or U17359 (N_17359,N_11229,N_6979);
nor U17360 (N_17360,N_6961,N_11347);
and U17361 (N_17361,N_11663,N_9832);
and U17362 (N_17362,N_9726,N_9395);
and U17363 (N_17363,N_7527,N_8195);
and U17364 (N_17364,N_7766,N_7032);
and U17365 (N_17365,N_7614,N_6337);
nand U17366 (N_17366,N_7780,N_6640);
or U17367 (N_17367,N_7289,N_11240);
and U17368 (N_17368,N_11559,N_9424);
xnor U17369 (N_17369,N_10189,N_11519);
nor U17370 (N_17370,N_11740,N_10045);
and U17371 (N_17371,N_11720,N_10434);
or U17372 (N_17372,N_8085,N_11061);
or U17373 (N_17373,N_7685,N_9708);
and U17374 (N_17374,N_9775,N_8662);
nor U17375 (N_17375,N_11813,N_8695);
nand U17376 (N_17376,N_9498,N_10869);
nor U17377 (N_17377,N_7874,N_11771);
nor U17378 (N_17378,N_9459,N_6935);
or U17379 (N_17379,N_9883,N_8513);
xor U17380 (N_17380,N_11459,N_7293);
nand U17381 (N_17381,N_7716,N_7111);
nand U17382 (N_17382,N_10343,N_10552);
nand U17383 (N_17383,N_8531,N_6212);
and U17384 (N_17384,N_7443,N_6170);
nor U17385 (N_17385,N_10761,N_10420);
and U17386 (N_17386,N_10555,N_6068);
nor U17387 (N_17387,N_7740,N_11134);
nand U17388 (N_17388,N_9030,N_11840);
nand U17389 (N_17389,N_6270,N_8887);
and U17390 (N_17390,N_11519,N_6413);
nand U17391 (N_17391,N_11157,N_7853);
and U17392 (N_17392,N_11544,N_6899);
or U17393 (N_17393,N_9595,N_10065);
nand U17394 (N_17394,N_7313,N_7791);
and U17395 (N_17395,N_8408,N_8391);
and U17396 (N_17396,N_11344,N_10964);
and U17397 (N_17397,N_8436,N_9491);
nor U17398 (N_17398,N_6350,N_9597);
nand U17399 (N_17399,N_6785,N_10486);
and U17400 (N_17400,N_10001,N_7305);
and U17401 (N_17401,N_9230,N_8346);
xnor U17402 (N_17402,N_7506,N_6139);
nor U17403 (N_17403,N_7913,N_6912);
and U17404 (N_17404,N_7657,N_10413);
xnor U17405 (N_17405,N_6433,N_11541);
nand U17406 (N_17406,N_10824,N_7321);
nand U17407 (N_17407,N_7068,N_11292);
nor U17408 (N_17408,N_9486,N_7630);
and U17409 (N_17409,N_9032,N_8123);
nand U17410 (N_17410,N_8412,N_7276);
nor U17411 (N_17411,N_11825,N_7501);
xnor U17412 (N_17412,N_11213,N_7544);
nand U17413 (N_17413,N_8715,N_11165);
nor U17414 (N_17414,N_10529,N_11949);
nor U17415 (N_17415,N_6659,N_6636);
or U17416 (N_17416,N_11086,N_6740);
and U17417 (N_17417,N_10743,N_9437);
nor U17418 (N_17418,N_10544,N_8492);
and U17419 (N_17419,N_11525,N_7381);
and U17420 (N_17420,N_9842,N_7255);
nand U17421 (N_17421,N_10560,N_10811);
and U17422 (N_17422,N_11519,N_11265);
and U17423 (N_17423,N_9246,N_11045);
and U17424 (N_17424,N_9171,N_6358);
nor U17425 (N_17425,N_11633,N_8451);
nand U17426 (N_17426,N_7520,N_10286);
xnor U17427 (N_17427,N_6925,N_8570);
and U17428 (N_17428,N_8042,N_8174);
and U17429 (N_17429,N_10927,N_8849);
nor U17430 (N_17430,N_10564,N_7506);
or U17431 (N_17431,N_7636,N_10770);
and U17432 (N_17432,N_11197,N_8682);
nor U17433 (N_17433,N_7520,N_7907);
or U17434 (N_17434,N_10443,N_9793);
and U17435 (N_17435,N_11800,N_6744);
nand U17436 (N_17436,N_8850,N_8934);
or U17437 (N_17437,N_7879,N_7957);
xnor U17438 (N_17438,N_6651,N_9089);
nand U17439 (N_17439,N_8570,N_10913);
or U17440 (N_17440,N_8313,N_6985);
xnor U17441 (N_17441,N_8310,N_8202);
or U17442 (N_17442,N_7048,N_11381);
xor U17443 (N_17443,N_7893,N_11884);
nor U17444 (N_17444,N_8684,N_7895);
nand U17445 (N_17445,N_7341,N_8451);
and U17446 (N_17446,N_9169,N_10559);
nand U17447 (N_17447,N_9620,N_10145);
or U17448 (N_17448,N_6978,N_11169);
nor U17449 (N_17449,N_8883,N_7165);
nand U17450 (N_17450,N_10051,N_8938);
nand U17451 (N_17451,N_10484,N_8373);
nor U17452 (N_17452,N_10594,N_8649);
and U17453 (N_17453,N_6452,N_10539);
or U17454 (N_17454,N_9186,N_11132);
or U17455 (N_17455,N_8117,N_10409);
nand U17456 (N_17456,N_11555,N_6996);
nor U17457 (N_17457,N_8906,N_10357);
xor U17458 (N_17458,N_9678,N_8146);
or U17459 (N_17459,N_7162,N_7033);
nand U17460 (N_17460,N_10484,N_6226);
nand U17461 (N_17461,N_9572,N_9356);
or U17462 (N_17462,N_11745,N_10514);
nand U17463 (N_17463,N_8829,N_10303);
or U17464 (N_17464,N_6797,N_11391);
nand U17465 (N_17465,N_11510,N_6559);
or U17466 (N_17466,N_7308,N_9095);
or U17467 (N_17467,N_11265,N_10556);
or U17468 (N_17468,N_10117,N_10460);
nand U17469 (N_17469,N_6091,N_8300);
xor U17470 (N_17470,N_7494,N_8616);
nor U17471 (N_17471,N_7098,N_8138);
or U17472 (N_17472,N_7424,N_9753);
nor U17473 (N_17473,N_10860,N_6171);
nand U17474 (N_17474,N_6954,N_8515);
nor U17475 (N_17475,N_7464,N_8601);
xor U17476 (N_17476,N_8404,N_11437);
and U17477 (N_17477,N_9978,N_10916);
and U17478 (N_17478,N_6470,N_8499);
xor U17479 (N_17479,N_11363,N_11414);
xor U17480 (N_17480,N_11961,N_9788);
nor U17481 (N_17481,N_11870,N_7491);
or U17482 (N_17482,N_11396,N_11146);
nand U17483 (N_17483,N_6401,N_11901);
and U17484 (N_17484,N_7491,N_11720);
nor U17485 (N_17485,N_11044,N_10168);
and U17486 (N_17486,N_9750,N_10347);
and U17487 (N_17487,N_10742,N_7298);
nor U17488 (N_17488,N_9475,N_9000);
nor U17489 (N_17489,N_6992,N_9425);
nor U17490 (N_17490,N_9769,N_6064);
or U17491 (N_17491,N_8078,N_6482);
nor U17492 (N_17492,N_11911,N_7518);
nor U17493 (N_17493,N_7398,N_10037);
nand U17494 (N_17494,N_8988,N_7527);
nor U17495 (N_17495,N_7742,N_7555);
or U17496 (N_17496,N_9165,N_9070);
and U17497 (N_17497,N_10837,N_10567);
nor U17498 (N_17498,N_10233,N_6204);
or U17499 (N_17499,N_6324,N_6400);
and U17500 (N_17500,N_8060,N_6675);
or U17501 (N_17501,N_6232,N_7000);
or U17502 (N_17502,N_7976,N_8880);
nand U17503 (N_17503,N_10210,N_6565);
nand U17504 (N_17504,N_7918,N_11548);
or U17505 (N_17505,N_10353,N_9847);
nand U17506 (N_17506,N_9357,N_11627);
nand U17507 (N_17507,N_8059,N_10565);
nor U17508 (N_17508,N_7910,N_11416);
nand U17509 (N_17509,N_10803,N_7035);
and U17510 (N_17510,N_8099,N_8403);
xor U17511 (N_17511,N_11942,N_9912);
xnor U17512 (N_17512,N_11940,N_10720);
or U17513 (N_17513,N_9081,N_6422);
or U17514 (N_17514,N_6313,N_7020);
and U17515 (N_17515,N_10308,N_8901);
and U17516 (N_17516,N_10885,N_7759);
nor U17517 (N_17517,N_8641,N_7475);
or U17518 (N_17518,N_10020,N_11793);
nor U17519 (N_17519,N_7601,N_10115);
and U17520 (N_17520,N_9106,N_10894);
xnor U17521 (N_17521,N_7618,N_8644);
and U17522 (N_17522,N_11666,N_10708);
nor U17523 (N_17523,N_11821,N_6174);
nor U17524 (N_17524,N_8656,N_11423);
nor U17525 (N_17525,N_11391,N_9595);
nand U17526 (N_17526,N_11344,N_8571);
nand U17527 (N_17527,N_10317,N_10879);
or U17528 (N_17528,N_9691,N_7595);
nor U17529 (N_17529,N_6462,N_11893);
and U17530 (N_17530,N_7996,N_6540);
nand U17531 (N_17531,N_9832,N_11849);
or U17532 (N_17532,N_6588,N_10590);
and U17533 (N_17533,N_6678,N_8275);
or U17534 (N_17534,N_10334,N_7464);
or U17535 (N_17535,N_8327,N_10467);
nand U17536 (N_17536,N_10669,N_10802);
nor U17537 (N_17537,N_9942,N_6955);
nor U17538 (N_17538,N_9340,N_8132);
nand U17539 (N_17539,N_6263,N_8676);
or U17540 (N_17540,N_8288,N_6901);
and U17541 (N_17541,N_7003,N_6176);
or U17542 (N_17542,N_10870,N_10133);
nor U17543 (N_17543,N_8318,N_8386);
and U17544 (N_17544,N_6661,N_10531);
and U17545 (N_17545,N_8278,N_11692);
xnor U17546 (N_17546,N_10719,N_11521);
or U17547 (N_17547,N_7096,N_10155);
xor U17548 (N_17548,N_6670,N_7821);
nor U17549 (N_17549,N_8776,N_10867);
nor U17550 (N_17550,N_11737,N_7150);
nor U17551 (N_17551,N_10283,N_6554);
xor U17552 (N_17552,N_6397,N_9910);
and U17553 (N_17553,N_9796,N_7195);
and U17554 (N_17554,N_9169,N_8275);
or U17555 (N_17555,N_10812,N_6243);
nor U17556 (N_17556,N_10040,N_11876);
or U17557 (N_17557,N_10063,N_10841);
nor U17558 (N_17558,N_9099,N_8351);
or U17559 (N_17559,N_7391,N_10720);
nand U17560 (N_17560,N_6898,N_7905);
nor U17561 (N_17561,N_7769,N_7804);
nor U17562 (N_17562,N_11470,N_10868);
or U17563 (N_17563,N_10838,N_11546);
and U17564 (N_17564,N_9067,N_10376);
xnor U17565 (N_17565,N_11824,N_11761);
nor U17566 (N_17566,N_7966,N_10603);
or U17567 (N_17567,N_6699,N_9728);
nor U17568 (N_17568,N_10888,N_11117);
and U17569 (N_17569,N_7848,N_7611);
nor U17570 (N_17570,N_10980,N_6832);
nor U17571 (N_17571,N_9553,N_11039);
and U17572 (N_17572,N_7317,N_11514);
nor U17573 (N_17573,N_9751,N_9781);
xor U17574 (N_17574,N_9229,N_8247);
nor U17575 (N_17575,N_10695,N_7816);
or U17576 (N_17576,N_11981,N_11132);
nand U17577 (N_17577,N_10015,N_8928);
and U17578 (N_17578,N_8806,N_9273);
and U17579 (N_17579,N_7421,N_9298);
and U17580 (N_17580,N_8278,N_6531);
or U17581 (N_17581,N_10825,N_10983);
and U17582 (N_17582,N_8190,N_9411);
nor U17583 (N_17583,N_10778,N_10885);
nand U17584 (N_17584,N_8373,N_8826);
nand U17585 (N_17585,N_9338,N_8704);
or U17586 (N_17586,N_10188,N_11124);
nand U17587 (N_17587,N_7207,N_10898);
nand U17588 (N_17588,N_7223,N_10252);
nor U17589 (N_17589,N_7836,N_11070);
nand U17590 (N_17590,N_7140,N_10617);
or U17591 (N_17591,N_6459,N_9505);
nor U17592 (N_17592,N_10515,N_10113);
nand U17593 (N_17593,N_11466,N_6616);
nand U17594 (N_17594,N_9369,N_10434);
or U17595 (N_17595,N_8518,N_7332);
or U17596 (N_17596,N_7515,N_11116);
nand U17597 (N_17597,N_10490,N_9739);
or U17598 (N_17598,N_8028,N_9189);
nor U17599 (N_17599,N_9577,N_8292);
or U17600 (N_17600,N_10100,N_6947);
nor U17601 (N_17601,N_8669,N_6568);
or U17602 (N_17602,N_7438,N_10054);
nor U17603 (N_17603,N_8000,N_7963);
nand U17604 (N_17604,N_11707,N_10961);
nand U17605 (N_17605,N_7142,N_6127);
nor U17606 (N_17606,N_8900,N_8758);
or U17607 (N_17607,N_10803,N_8791);
nand U17608 (N_17608,N_7866,N_6701);
nor U17609 (N_17609,N_9876,N_11034);
or U17610 (N_17610,N_11755,N_6985);
nand U17611 (N_17611,N_9767,N_11836);
nor U17612 (N_17612,N_8656,N_10145);
and U17613 (N_17613,N_11638,N_9684);
or U17614 (N_17614,N_7805,N_10429);
nor U17615 (N_17615,N_6851,N_10864);
and U17616 (N_17616,N_8428,N_9888);
nor U17617 (N_17617,N_6808,N_7583);
and U17618 (N_17618,N_9778,N_11724);
and U17619 (N_17619,N_11295,N_7010);
and U17620 (N_17620,N_6196,N_7789);
or U17621 (N_17621,N_11381,N_9116);
and U17622 (N_17622,N_8678,N_9681);
or U17623 (N_17623,N_9224,N_9263);
nor U17624 (N_17624,N_7033,N_6535);
nor U17625 (N_17625,N_8651,N_6426);
or U17626 (N_17626,N_7532,N_8498);
nor U17627 (N_17627,N_8834,N_8384);
and U17628 (N_17628,N_8838,N_9044);
and U17629 (N_17629,N_7147,N_7293);
nand U17630 (N_17630,N_11160,N_6718);
nor U17631 (N_17631,N_7891,N_7326);
and U17632 (N_17632,N_7244,N_6348);
or U17633 (N_17633,N_8212,N_6322);
nor U17634 (N_17634,N_9758,N_9242);
or U17635 (N_17635,N_11441,N_7784);
nand U17636 (N_17636,N_7502,N_10290);
and U17637 (N_17637,N_6385,N_11442);
nor U17638 (N_17638,N_10320,N_11959);
nand U17639 (N_17639,N_9261,N_11986);
nor U17640 (N_17640,N_10179,N_11904);
or U17641 (N_17641,N_10728,N_10108);
and U17642 (N_17642,N_6244,N_11691);
or U17643 (N_17643,N_9225,N_8799);
and U17644 (N_17644,N_9403,N_7431);
nand U17645 (N_17645,N_9264,N_9549);
or U17646 (N_17646,N_9922,N_6717);
nor U17647 (N_17647,N_8148,N_9531);
and U17648 (N_17648,N_6693,N_8157);
or U17649 (N_17649,N_11002,N_6303);
or U17650 (N_17650,N_10574,N_9633);
nand U17651 (N_17651,N_11341,N_9470);
nand U17652 (N_17652,N_9418,N_7108);
nor U17653 (N_17653,N_7342,N_11223);
or U17654 (N_17654,N_6882,N_11846);
nand U17655 (N_17655,N_10793,N_9321);
nor U17656 (N_17656,N_6014,N_8830);
or U17657 (N_17657,N_11311,N_8520);
nor U17658 (N_17658,N_9632,N_10369);
nor U17659 (N_17659,N_8253,N_9357);
nor U17660 (N_17660,N_6499,N_8061);
and U17661 (N_17661,N_10315,N_11192);
nor U17662 (N_17662,N_11504,N_7396);
nand U17663 (N_17663,N_9938,N_11860);
and U17664 (N_17664,N_9149,N_10050);
and U17665 (N_17665,N_10748,N_8056);
xor U17666 (N_17666,N_8106,N_8964);
and U17667 (N_17667,N_8632,N_8797);
and U17668 (N_17668,N_11562,N_7389);
or U17669 (N_17669,N_11126,N_9635);
nand U17670 (N_17670,N_9527,N_6842);
and U17671 (N_17671,N_8810,N_10909);
nor U17672 (N_17672,N_11147,N_7304);
nor U17673 (N_17673,N_6266,N_6064);
or U17674 (N_17674,N_10957,N_10247);
nor U17675 (N_17675,N_8329,N_8964);
and U17676 (N_17676,N_9609,N_9161);
and U17677 (N_17677,N_9461,N_7584);
and U17678 (N_17678,N_9622,N_11046);
nor U17679 (N_17679,N_7471,N_9043);
nand U17680 (N_17680,N_7674,N_7258);
and U17681 (N_17681,N_11688,N_9826);
nand U17682 (N_17682,N_6907,N_10932);
or U17683 (N_17683,N_10577,N_8127);
and U17684 (N_17684,N_8829,N_9398);
or U17685 (N_17685,N_11684,N_11346);
nand U17686 (N_17686,N_11134,N_11450);
nand U17687 (N_17687,N_6608,N_10099);
nand U17688 (N_17688,N_6592,N_7795);
nor U17689 (N_17689,N_7443,N_10207);
and U17690 (N_17690,N_8572,N_9367);
and U17691 (N_17691,N_7657,N_11727);
nand U17692 (N_17692,N_9963,N_7471);
and U17693 (N_17693,N_11038,N_7234);
or U17694 (N_17694,N_7532,N_9620);
nor U17695 (N_17695,N_9174,N_7336);
and U17696 (N_17696,N_9585,N_10220);
nor U17697 (N_17697,N_8928,N_11208);
or U17698 (N_17698,N_7786,N_9883);
or U17699 (N_17699,N_6109,N_7316);
nor U17700 (N_17700,N_8923,N_9259);
and U17701 (N_17701,N_8330,N_11030);
nand U17702 (N_17702,N_10867,N_8888);
nand U17703 (N_17703,N_8937,N_6067);
nor U17704 (N_17704,N_7548,N_8840);
nand U17705 (N_17705,N_7212,N_11006);
or U17706 (N_17706,N_8507,N_7545);
and U17707 (N_17707,N_7514,N_9844);
nand U17708 (N_17708,N_6551,N_6615);
and U17709 (N_17709,N_11144,N_7818);
nand U17710 (N_17710,N_7855,N_6186);
xnor U17711 (N_17711,N_11678,N_10961);
nor U17712 (N_17712,N_7447,N_9790);
nor U17713 (N_17713,N_6500,N_9612);
nand U17714 (N_17714,N_7744,N_7222);
nand U17715 (N_17715,N_6743,N_11612);
nand U17716 (N_17716,N_6427,N_8081);
xnor U17717 (N_17717,N_8657,N_9348);
and U17718 (N_17718,N_11645,N_10791);
or U17719 (N_17719,N_10603,N_7178);
and U17720 (N_17720,N_7716,N_10467);
and U17721 (N_17721,N_9987,N_11756);
or U17722 (N_17722,N_9028,N_6506);
nor U17723 (N_17723,N_11148,N_8876);
nand U17724 (N_17724,N_11484,N_9734);
or U17725 (N_17725,N_10965,N_11550);
nor U17726 (N_17726,N_7314,N_6256);
and U17727 (N_17727,N_7682,N_9837);
xor U17728 (N_17728,N_9309,N_8397);
and U17729 (N_17729,N_11221,N_11656);
or U17730 (N_17730,N_9028,N_11210);
and U17731 (N_17731,N_11342,N_11024);
nand U17732 (N_17732,N_11082,N_7750);
xnor U17733 (N_17733,N_10426,N_11687);
and U17734 (N_17734,N_7333,N_8287);
nand U17735 (N_17735,N_11419,N_8150);
or U17736 (N_17736,N_7390,N_8516);
or U17737 (N_17737,N_11157,N_6428);
xor U17738 (N_17738,N_6719,N_6004);
nor U17739 (N_17739,N_6832,N_10998);
nand U17740 (N_17740,N_10240,N_7984);
nor U17741 (N_17741,N_10809,N_8521);
or U17742 (N_17742,N_8324,N_6104);
and U17743 (N_17743,N_11297,N_11487);
nand U17744 (N_17744,N_6082,N_10043);
and U17745 (N_17745,N_9201,N_7830);
and U17746 (N_17746,N_8805,N_8757);
or U17747 (N_17747,N_8793,N_9467);
nor U17748 (N_17748,N_9497,N_7212);
and U17749 (N_17749,N_6756,N_7363);
xor U17750 (N_17750,N_7775,N_10673);
and U17751 (N_17751,N_6545,N_9603);
nor U17752 (N_17752,N_6809,N_6847);
xor U17753 (N_17753,N_10849,N_11848);
nor U17754 (N_17754,N_8796,N_9171);
and U17755 (N_17755,N_10426,N_8014);
xnor U17756 (N_17756,N_8074,N_8973);
nor U17757 (N_17757,N_10934,N_6758);
nor U17758 (N_17758,N_10075,N_7554);
xnor U17759 (N_17759,N_11995,N_7193);
nand U17760 (N_17760,N_7440,N_6093);
and U17761 (N_17761,N_10017,N_6034);
nand U17762 (N_17762,N_8852,N_8760);
nand U17763 (N_17763,N_9916,N_10177);
nor U17764 (N_17764,N_9472,N_6734);
nand U17765 (N_17765,N_7575,N_6820);
nand U17766 (N_17766,N_9919,N_9163);
or U17767 (N_17767,N_9321,N_7507);
nor U17768 (N_17768,N_8549,N_8512);
or U17769 (N_17769,N_9650,N_9663);
or U17770 (N_17770,N_6172,N_7186);
nor U17771 (N_17771,N_10813,N_10893);
nor U17772 (N_17772,N_7433,N_8830);
nor U17773 (N_17773,N_7369,N_6921);
and U17774 (N_17774,N_7508,N_11248);
and U17775 (N_17775,N_9983,N_7779);
nand U17776 (N_17776,N_7595,N_6863);
nor U17777 (N_17777,N_11028,N_7093);
and U17778 (N_17778,N_7827,N_11280);
xnor U17779 (N_17779,N_8392,N_8972);
or U17780 (N_17780,N_11880,N_11186);
nor U17781 (N_17781,N_11580,N_9253);
nand U17782 (N_17782,N_6396,N_7122);
and U17783 (N_17783,N_6791,N_9744);
or U17784 (N_17784,N_11934,N_9693);
nand U17785 (N_17785,N_8590,N_8774);
and U17786 (N_17786,N_6654,N_7601);
nor U17787 (N_17787,N_9231,N_10721);
and U17788 (N_17788,N_6528,N_6861);
and U17789 (N_17789,N_10122,N_9581);
or U17790 (N_17790,N_6718,N_7819);
and U17791 (N_17791,N_11447,N_7180);
nor U17792 (N_17792,N_10502,N_7128);
xor U17793 (N_17793,N_7004,N_7703);
nand U17794 (N_17794,N_8739,N_6394);
nor U17795 (N_17795,N_6916,N_9832);
xor U17796 (N_17796,N_10479,N_9963);
nand U17797 (N_17797,N_6023,N_6754);
and U17798 (N_17798,N_8315,N_8358);
or U17799 (N_17799,N_9626,N_10163);
nor U17800 (N_17800,N_7797,N_7822);
and U17801 (N_17801,N_6586,N_6478);
and U17802 (N_17802,N_11858,N_7140);
and U17803 (N_17803,N_6903,N_7328);
nor U17804 (N_17804,N_10705,N_9029);
nor U17805 (N_17805,N_6413,N_10669);
nand U17806 (N_17806,N_7643,N_11183);
or U17807 (N_17807,N_8475,N_9370);
xor U17808 (N_17808,N_10993,N_6558);
or U17809 (N_17809,N_6441,N_6657);
or U17810 (N_17810,N_9215,N_10489);
nand U17811 (N_17811,N_7550,N_7166);
or U17812 (N_17812,N_7297,N_9545);
nand U17813 (N_17813,N_11606,N_7414);
nor U17814 (N_17814,N_6657,N_7635);
nand U17815 (N_17815,N_11957,N_11603);
nor U17816 (N_17816,N_7720,N_11358);
nor U17817 (N_17817,N_10670,N_7758);
xnor U17818 (N_17818,N_11033,N_7587);
nand U17819 (N_17819,N_6924,N_8621);
nor U17820 (N_17820,N_7986,N_7251);
and U17821 (N_17821,N_8047,N_7140);
nor U17822 (N_17822,N_8825,N_8139);
or U17823 (N_17823,N_11933,N_10675);
nor U17824 (N_17824,N_7226,N_8734);
or U17825 (N_17825,N_8283,N_6341);
or U17826 (N_17826,N_8999,N_6695);
nor U17827 (N_17827,N_6169,N_10002);
and U17828 (N_17828,N_6310,N_11540);
nor U17829 (N_17829,N_6019,N_9601);
and U17830 (N_17830,N_8450,N_9961);
nor U17831 (N_17831,N_10327,N_11781);
nor U17832 (N_17832,N_7815,N_7024);
or U17833 (N_17833,N_6641,N_7860);
nand U17834 (N_17834,N_9198,N_11751);
nor U17835 (N_17835,N_7999,N_8002);
and U17836 (N_17836,N_10499,N_7045);
nor U17837 (N_17837,N_7281,N_11760);
or U17838 (N_17838,N_6014,N_6502);
and U17839 (N_17839,N_8857,N_7877);
nand U17840 (N_17840,N_7756,N_7470);
and U17841 (N_17841,N_9431,N_6043);
nor U17842 (N_17842,N_8902,N_6527);
nand U17843 (N_17843,N_10558,N_6904);
nor U17844 (N_17844,N_9262,N_8950);
nor U17845 (N_17845,N_10154,N_11263);
xnor U17846 (N_17846,N_11478,N_10240);
and U17847 (N_17847,N_6382,N_10403);
and U17848 (N_17848,N_11065,N_11594);
nor U17849 (N_17849,N_7691,N_10631);
and U17850 (N_17850,N_10734,N_8325);
and U17851 (N_17851,N_11513,N_10328);
xor U17852 (N_17852,N_11612,N_6677);
nand U17853 (N_17853,N_6230,N_11940);
nand U17854 (N_17854,N_9987,N_11904);
or U17855 (N_17855,N_10958,N_9829);
nand U17856 (N_17856,N_7294,N_8235);
nand U17857 (N_17857,N_10272,N_9413);
and U17858 (N_17858,N_6414,N_10819);
or U17859 (N_17859,N_10962,N_9063);
xnor U17860 (N_17860,N_7021,N_6351);
nand U17861 (N_17861,N_10544,N_10069);
nand U17862 (N_17862,N_9836,N_6695);
or U17863 (N_17863,N_11395,N_11799);
xnor U17864 (N_17864,N_10313,N_10773);
nand U17865 (N_17865,N_6983,N_11120);
and U17866 (N_17866,N_11508,N_10026);
and U17867 (N_17867,N_11933,N_8583);
or U17868 (N_17868,N_6283,N_6798);
nand U17869 (N_17869,N_11244,N_7174);
nor U17870 (N_17870,N_6753,N_6061);
or U17871 (N_17871,N_10392,N_9872);
and U17872 (N_17872,N_7403,N_11588);
and U17873 (N_17873,N_11820,N_7967);
nand U17874 (N_17874,N_7443,N_6645);
nand U17875 (N_17875,N_7919,N_9702);
and U17876 (N_17876,N_8292,N_9912);
nor U17877 (N_17877,N_11637,N_8388);
nand U17878 (N_17878,N_8699,N_9016);
xor U17879 (N_17879,N_6150,N_10113);
nor U17880 (N_17880,N_10912,N_10804);
or U17881 (N_17881,N_11226,N_10735);
nor U17882 (N_17882,N_6391,N_11947);
nand U17883 (N_17883,N_8054,N_8642);
xnor U17884 (N_17884,N_8540,N_9793);
or U17885 (N_17885,N_8241,N_10852);
nand U17886 (N_17886,N_6094,N_8226);
or U17887 (N_17887,N_6296,N_8341);
nor U17888 (N_17888,N_8233,N_11201);
nand U17889 (N_17889,N_6384,N_8768);
and U17890 (N_17890,N_10974,N_8395);
xnor U17891 (N_17891,N_6128,N_9922);
or U17892 (N_17892,N_9662,N_9541);
xor U17893 (N_17893,N_6695,N_7058);
or U17894 (N_17894,N_10026,N_8860);
nand U17895 (N_17895,N_6203,N_8686);
or U17896 (N_17896,N_7050,N_10095);
or U17897 (N_17897,N_10275,N_9583);
nand U17898 (N_17898,N_7472,N_6602);
nand U17899 (N_17899,N_10335,N_7231);
and U17900 (N_17900,N_7977,N_10883);
and U17901 (N_17901,N_7977,N_10927);
nand U17902 (N_17902,N_9092,N_10918);
xor U17903 (N_17903,N_10321,N_6849);
and U17904 (N_17904,N_10892,N_10354);
nor U17905 (N_17905,N_7801,N_6941);
nor U17906 (N_17906,N_11924,N_6651);
nand U17907 (N_17907,N_8039,N_7880);
nor U17908 (N_17908,N_10179,N_11010);
and U17909 (N_17909,N_7792,N_11048);
nand U17910 (N_17910,N_6303,N_6945);
and U17911 (N_17911,N_11982,N_9432);
or U17912 (N_17912,N_10752,N_6671);
nand U17913 (N_17913,N_10207,N_6869);
and U17914 (N_17914,N_9423,N_10466);
nand U17915 (N_17915,N_10931,N_11449);
nor U17916 (N_17916,N_10839,N_11809);
or U17917 (N_17917,N_10043,N_7230);
nand U17918 (N_17918,N_7040,N_7850);
nand U17919 (N_17919,N_10748,N_9477);
or U17920 (N_17920,N_9866,N_11967);
nor U17921 (N_17921,N_9162,N_8156);
xor U17922 (N_17922,N_8335,N_11301);
nand U17923 (N_17923,N_7719,N_11478);
nor U17924 (N_17924,N_7802,N_9122);
and U17925 (N_17925,N_9324,N_8392);
and U17926 (N_17926,N_8418,N_8505);
xor U17927 (N_17927,N_10676,N_8418);
xor U17928 (N_17928,N_10994,N_6758);
nand U17929 (N_17929,N_9295,N_6957);
nor U17930 (N_17930,N_6338,N_7902);
or U17931 (N_17931,N_6341,N_9656);
nor U17932 (N_17932,N_11366,N_7728);
and U17933 (N_17933,N_11426,N_11572);
xnor U17934 (N_17934,N_8341,N_6033);
nor U17935 (N_17935,N_6030,N_11296);
nand U17936 (N_17936,N_7330,N_6619);
or U17937 (N_17937,N_8569,N_10686);
or U17938 (N_17938,N_7161,N_9082);
or U17939 (N_17939,N_7608,N_7129);
and U17940 (N_17940,N_7911,N_10158);
and U17941 (N_17941,N_10320,N_7225);
and U17942 (N_17942,N_8688,N_6820);
and U17943 (N_17943,N_11586,N_9488);
nor U17944 (N_17944,N_8635,N_7590);
nand U17945 (N_17945,N_10379,N_7894);
or U17946 (N_17946,N_10286,N_9551);
nor U17947 (N_17947,N_8549,N_9213);
and U17948 (N_17948,N_11077,N_11627);
and U17949 (N_17949,N_8241,N_9861);
nand U17950 (N_17950,N_9910,N_7875);
nor U17951 (N_17951,N_8163,N_6605);
nor U17952 (N_17952,N_7837,N_9994);
or U17953 (N_17953,N_9453,N_11757);
or U17954 (N_17954,N_10229,N_9737);
or U17955 (N_17955,N_9899,N_8834);
xor U17956 (N_17956,N_8011,N_7955);
or U17957 (N_17957,N_11806,N_7823);
or U17958 (N_17958,N_6858,N_6837);
nor U17959 (N_17959,N_11747,N_8374);
nand U17960 (N_17960,N_9031,N_9398);
and U17961 (N_17961,N_11145,N_8284);
and U17962 (N_17962,N_10370,N_10199);
xnor U17963 (N_17963,N_11117,N_11692);
nand U17964 (N_17964,N_11984,N_11840);
and U17965 (N_17965,N_10912,N_8942);
or U17966 (N_17966,N_8196,N_10832);
nor U17967 (N_17967,N_7257,N_7627);
or U17968 (N_17968,N_7564,N_9632);
nand U17969 (N_17969,N_8040,N_6397);
nor U17970 (N_17970,N_11551,N_11972);
xor U17971 (N_17971,N_6528,N_8073);
nand U17972 (N_17972,N_6607,N_10123);
or U17973 (N_17973,N_11834,N_9555);
or U17974 (N_17974,N_9736,N_7081);
and U17975 (N_17975,N_11179,N_8873);
or U17976 (N_17976,N_11728,N_8360);
nand U17977 (N_17977,N_7918,N_6069);
nand U17978 (N_17978,N_7709,N_8508);
nor U17979 (N_17979,N_7929,N_6100);
or U17980 (N_17980,N_11074,N_10037);
nand U17981 (N_17981,N_9745,N_7615);
nor U17982 (N_17982,N_10294,N_8344);
and U17983 (N_17983,N_9520,N_9396);
and U17984 (N_17984,N_9918,N_6572);
and U17985 (N_17985,N_11387,N_7404);
nor U17986 (N_17986,N_10608,N_11821);
nor U17987 (N_17987,N_10871,N_9210);
xnor U17988 (N_17988,N_9982,N_9389);
and U17989 (N_17989,N_6173,N_11683);
xnor U17990 (N_17990,N_9851,N_8594);
and U17991 (N_17991,N_8967,N_8370);
and U17992 (N_17992,N_9440,N_9826);
nand U17993 (N_17993,N_10655,N_7757);
or U17994 (N_17994,N_9951,N_7226);
and U17995 (N_17995,N_11487,N_6560);
or U17996 (N_17996,N_10811,N_6243);
or U17997 (N_17997,N_8141,N_8680);
or U17998 (N_17998,N_6015,N_7448);
or U17999 (N_17999,N_9817,N_7606);
nand U18000 (N_18000,N_16626,N_17017);
and U18001 (N_18001,N_17871,N_12903);
nor U18002 (N_18002,N_15427,N_14387);
nor U18003 (N_18003,N_14209,N_16591);
or U18004 (N_18004,N_15585,N_17409);
or U18005 (N_18005,N_12058,N_14747);
nand U18006 (N_18006,N_14970,N_15798);
nand U18007 (N_18007,N_14153,N_16069);
nand U18008 (N_18008,N_17684,N_13755);
and U18009 (N_18009,N_14896,N_14127);
and U18010 (N_18010,N_15945,N_13411);
or U18011 (N_18011,N_16924,N_12392);
nor U18012 (N_18012,N_12296,N_17220);
or U18013 (N_18013,N_14635,N_14894);
or U18014 (N_18014,N_16759,N_15528);
nand U18015 (N_18015,N_15034,N_12937);
or U18016 (N_18016,N_13703,N_16129);
and U18017 (N_18017,N_13350,N_17571);
nor U18018 (N_18018,N_14562,N_12872);
xnor U18019 (N_18019,N_14689,N_14913);
nor U18020 (N_18020,N_15865,N_13460);
and U18021 (N_18021,N_15363,N_14015);
nor U18022 (N_18022,N_13534,N_17381);
xnor U18023 (N_18023,N_14488,N_16170);
and U18024 (N_18024,N_15048,N_15820);
nand U18025 (N_18025,N_15184,N_14274);
nand U18026 (N_18026,N_12482,N_15937);
xor U18027 (N_18027,N_16314,N_15221);
xor U18028 (N_18028,N_17654,N_16784);
and U18029 (N_18029,N_13255,N_13836);
or U18030 (N_18030,N_16427,N_17345);
nor U18031 (N_18031,N_14502,N_13256);
nand U18032 (N_18032,N_14926,N_13257);
or U18033 (N_18033,N_17576,N_15892);
nor U18034 (N_18034,N_12632,N_17940);
nor U18035 (N_18035,N_16773,N_15115);
nor U18036 (N_18036,N_17064,N_13389);
and U18037 (N_18037,N_13502,N_12253);
nor U18038 (N_18038,N_13833,N_16143);
nand U18039 (N_18039,N_16823,N_14371);
nor U18040 (N_18040,N_12424,N_16769);
and U18041 (N_18041,N_17330,N_13192);
or U18042 (N_18042,N_16414,N_14220);
and U18043 (N_18043,N_14390,N_17873);
xnor U18044 (N_18044,N_15842,N_13537);
nand U18045 (N_18045,N_15959,N_15822);
or U18046 (N_18046,N_13203,N_13393);
or U18047 (N_18047,N_14658,N_17586);
nand U18048 (N_18048,N_13417,N_12250);
and U18049 (N_18049,N_16426,N_17605);
xnor U18050 (N_18050,N_15011,N_12785);
nand U18051 (N_18051,N_17096,N_15452);
nand U18052 (N_18052,N_12023,N_15101);
nand U18053 (N_18053,N_13967,N_15881);
and U18054 (N_18054,N_15387,N_14656);
nor U18055 (N_18055,N_15744,N_17322);
and U18056 (N_18056,N_12752,N_12748);
nand U18057 (N_18057,N_15480,N_13916);
nor U18058 (N_18058,N_17513,N_14580);
and U18059 (N_18059,N_14565,N_17315);
nand U18060 (N_18060,N_17868,N_15830);
nand U18061 (N_18061,N_17420,N_14255);
nand U18062 (N_18062,N_17189,N_17646);
xor U18063 (N_18063,N_17151,N_16188);
nand U18064 (N_18064,N_13463,N_14944);
nand U18065 (N_18065,N_13337,N_12866);
or U18066 (N_18066,N_14461,N_13218);
nand U18067 (N_18067,N_15500,N_14105);
or U18068 (N_18068,N_13541,N_13959);
or U18069 (N_18069,N_14285,N_16517);
or U18070 (N_18070,N_16142,N_15467);
and U18071 (N_18071,N_15326,N_12894);
nor U18072 (N_18072,N_14150,N_14763);
nor U18073 (N_18073,N_14422,N_13662);
and U18074 (N_18074,N_15025,N_17369);
and U18075 (N_18075,N_12484,N_15149);
or U18076 (N_18076,N_13615,N_17737);
or U18077 (N_18077,N_12323,N_14912);
or U18078 (N_18078,N_17145,N_17668);
and U18079 (N_18079,N_17792,N_15927);
or U18080 (N_18080,N_15251,N_13569);
and U18081 (N_18081,N_16471,N_12462);
and U18082 (N_18082,N_14138,N_14732);
nand U18083 (N_18083,N_12855,N_14536);
nand U18084 (N_18084,N_16052,N_14631);
and U18085 (N_18085,N_13596,N_15999);
or U18086 (N_18086,N_16841,N_12776);
nand U18087 (N_18087,N_15590,N_16323);
or U18088 (N_18088,N_12681,N_13905);
xnor U18089 (N_18089,N_13206,N_13428);
xnor U18090 (N_18090,N_15209,N_13369);
xnor U18091 (N_18091,N_15155,N_13957);
xor U18092 (N_18092,N_13397,N_15236);
xnor U18093 (N_18093,N_12832,N_15206);
or U18094 (N_18094,N_16801,N_17262);
and U18095 (N_18095,N_16435,N_16293);
nand U18096 (N_18096,N_15402,N_12810);
nor U18097 (N_18097,N_13012,N_12616);
nand U18098 (N_18098,N_16523,N_13374);
or U18099 (N_18099,N_13189,N_17698);
nor U18100 (N_18100,N_13077,N_16086);
and U18101 (N_18101,N_12517,N_14554);
nand U18102 (N_18102,N_14675,N_17298);
or U18103 (N_18103,N_14762,N_16429);
and U18104 (N_18104,N_12339,N_15435);
nor U18105 (N_18105,N_12581,N_17713);
nand U18106 (N_18106,N_12825,N_15022);
or U18107 (N_18107,N_13222,N_12699);
and U18108 (N_18108,N_16265,N_14979);
nand U18109 (N_18109,N_14314,N_17986);
or U18110 (N_18110,N_17647,N_17196);
nor U18111 (N_18111,N_13367,N_15990);
or U18112 (N_18112,N_17612,N_17689);
or U18113 (N_18113,N_12527,N_16346);
nand U18114 (N_18114,N_15385,N_14780);
nand U18115 (N_18115,N_15168,N_12508);
nand U18116 (N_18116,N_14609,N_16957);
nor U18117 (N_18117,N_13447,N_12700);
nand U18118 (N_18118,N_12698,N_14339);
and U18119 (N_18119,N_16425,N_16187);
and U18120 (N_18120,N_12818,N_16623);
nand U18121 (N_18121,N_13119,N_16139);
and U18122 (N_18122,N_12547,N_13053);
and U18123 (N_18123,N_12912,N_14513);
nand U18124 (N_18124,N_16900,N_13507);
nand U18125 (N_18125,N_14578,N_17523);
nor U18126 (N_18126,N_14409,N_14813);
xnor U18127 (N_18127,N_16544,N_14332);
or U18128 (N_18128,N_13995,N_17815);
nor U18129 (N_18129,N_14289,N_12704);
or U18130 (N_18130,N_16621,N_14741);
nor U18131 (N_18131,N_16467,N_17499);
and U18132 (N_18132,N_15083,N_14602);
or U18133 (N_18133,N_13472,N_16761);
or U18134 (N_18134,N_15190,N_16412);
and U18135 (N_18135,N_17246,N_16787);
or U18136 (N_18136,N_15028,N_15694);
nand U18137 (N_18137,N_13558,N_14610);
nand U18138 (N_18138,N_12230,N_15741);
nand U18139 (N_18139,N_13835,N_15476);
or U18140 (N_18140,N_15026,N_15068);
xor U18141 (N_18141,N_15245,N_15051);
or U18142 (N_18142,N_13830,N_14987);
xor U18143 (N_18143,N_14383,N_17733);
nor U18144 (N_18144,N_12823,N_16961);
nand U18145 (N_18145,N_17888,N_17492);
or U18146 (N_18146,N_17990,N_14948);
nor U18147 (N_18147,N_14052,N_15644);
or U18148 (N_18148,N_12404,N_13184);
nor U18149 (N_18149,N_17756,N_15244);
nand U18150 (N_18150,N_13887,N_12329);
nand U18151 (N_18151,N_12430,N_16689);
and U18152 (N_18152,N_16887,N_13055);
nand U18153 (N_18153,N_13458,N_14393);
nand U18154 (N_18154,N_16655,N_12728);
nand U18155 (N_18155,N_16227,N_15040);
and U18156 (N_18156,N_12348,N_15570);
xnor U18157 (N_18157,N_17263,N_12035);
nand U18158 (N_18158,N_13088,N_16388);
nor U18159 (N_18159,N_15648,N_16844);
and U18160 (N_18160,N_14438,N_12958);
nor U18161 (N_18161,N_16356,N_16449);
nand U18162 (N_18162,N_12809,N_13542);
nor U18163 (N_18163,N_17944,N_16145);
or U18164 (N_18164,N_12051,N_13092);
xor U18165 (N_18165,N_17349,N_15786);
or U18166 (N_18166,N_16124,N_12934);
or U18167 (N_18167,N_17179,N_15855);
nor U18168 (N_18168,N_17811,N_13038);
and U18169 (N_18169,N_12350,N_14096);
xor U18170 (N_18170,N_13820,N_13545);
or U18171 (N_18171,N_16690,N_13501);
nor U18172 (N_18172,N_12237,N_12852);
or U18173 (N_18173,N_16223,N_16861);
or U18174 (N_18174,N_15611,N_15941);
or U18175 (N_18175,N_14938,N_14873);
nor U18176 (N_18176,N_17209,N_16409);
nor U18177 (N_18177,N_16751,N_13348);
nor U18178 (N_18178,N_13332,N_17639);
nand U18179 (N_18179,N_15397,N_14687);
nand U18180 (N_18180,N_12873,N_14801);
and U18181 (N_18181,N_12732,N_12883);
nand U18182 (N_18182,N_15535,N_17242);
or U18183 (N_18183,N_16664,N_13150);
nor U18184 (N_18184,N_17249,N_12477);
or U18185 (N_18185,N_17665,N_13111);
or U18186 (N_18186,N_16274,N_16110);
nand U18187 (N_18187,N_15507,N_15984);
nor U18188 (N_18188,N_14297,N_13095);
nor U18189 (N_18189,N_17552,N_16553);
or U18190 (N_18190,N_14647,N_12762);
nand U18191 (N_18191,N_14047,N_14521);
and U18192 (N_18192,N_16081,N_14112);
or U18193 (N_18193,N_15808,N_16629);
or U18194 (N_18194,N_13765,N_15204);
or U18195 (N_18195,N_13052,N_17254);
and U18196 (N_18196,N_17769,N_12111);
and U18197 (N_18197,N_14241,N_12099);
or U18198 (N_18198,N_13028,N_15376);
or U18199 (N_18199,N_15750,N_12869);
or U18200 (N_18200,N_14910,N_13990);
nor U18201 (N_18201,N_12901,N_17282);
and U18202 (N_18202,N_17454,N_17204);
nand U18203 (N_18203,N_14778,N_14365);
nand U18204 (N_18204,N_17724,N_16648);
or U18205 (N_18205,N_13778,N_15112);
xor U18206 (N_18206,N_13375,N_15021);
nand U18207 (N_18207,N_15304,N_16041);
or U18208 (N_18208,N_12624,N_17182);
and U18209 (N_18209,N_15958,N_12672);
and U18210 (N_18210,N_14625,N_17116);
and U18211 (N_18211,N_13193,N_17915);
nor U18212 (N_18212,N_12980,N_12805);
nor U18213 (N_18213,N_14092,N_13847);
nor U18214 (N_18214,N_12360,N_15605);
nand U18215 (N_18215,N_15854,N_13964);
and U18216 (N_18216,N_15488,N_15131);
or U18217 (N_18217,N_14564,N_17983);
nor U18218 (N_18218,N_15567,N_12028);
and U18219 (N_18219,N_16739,N_13180);
nand U18220 (N_18220,N_14142,N_12629);
nand U18221 (N_18221,N_17895,N_15721);
nand U18222 (N_18222,N_14341,N_13761);
nand U18223 (N_18223,N_16277,N_13041);
nor U18224 (N_18224,N_12463,N_13285);
xnor U18225 (N_18225,N_17533,N_15866);
or U18226 (N_18226,N_14522,N_13479);
and U18227 (N_18227,N_14799,N_14369);
nand U18228 (N_18228,N_14348,N_13081);
nor U18229 (N_18229,N_12145,N_12812);
or U18230 (N_18230,N_15166,N_14198);
xor U18231 (N_18231,N_17408,N_16272);
and U18232 (N_18232,N_15041,N_16260);
or U18233 (N_18233,N_17743,N_15635);
nand U18234 (N_18234,N_15268,N_16300);
nand U18235 (N_18235,N_17098,N_15875);
nand U18236 (N_18236,N_16952,N_17467);
nor U18237 (N_18237,N_15153,N_16093);
xnor U18238 (N_18238,N_16672,N_15401);
or U18239 (N_18239,N_15270,N_15829);
nor U18240 (N_18240,N_17723,N_16509);
or U18241 (N_18241,N_12643,N_14247);
or U18242 (N_18242,N_14306,N_12718);
nor U18243 (N_18243,N_13171,N_13293);
nor U18244 (N_18244,N_12181,N_17522);
and U18245 (N_18245,N_13554,N_16804);
or U18246 (N_18246,N_13614,N_15896);
or U18247 (N_18247,N_16497,N_12514);
and U18248 (N_18248,N_17329,N_17909);
or U18249 (N_18249,N_16975,N_14161);
nor U18250 (N_18250,N_15754,N_13767);
or U18251 (N_18251,N_13823,N_13717);
xor U18252 (N_18252,N_13602,N_13186);
and U18253 (N_18253,N_16571,N_13704);
and U18254 (N_18254,N_13110,N_14388);
and U18255 (N_18255,N_14962,N_17540);
and U18256 (N_18256,N_16458,N_14943);
and U18257 (N_18257,N_12995,N_15349);
nand U18258 (N_18258,N_13327,N_12331);
nor U18259 (N_18259,N_12496,N_16728);
and U18260 (N_18260,N_17122,N_14680);
nand U18261 (N_18261,N_17328,N_15019);
or U18262 (N_18262,N_17334,N_17047);
nor U18263 (N_18263,N_12357,N_15092);
nor U18264 (N_18264,N_13581,N_13082);
or U18265 (N_18265,N_13888,N_15716);
and U18266 (N_18266,N_12723,N_14405);
or U18267 (N_18267,N_16935,N_15237);
xor U18268 (N_18268,N_14002,N_17163);
and U18269 (N_18269,N_15793,N_16051);
or U18270 (N_18270,N_17350,N_17885);
nor U18271 (N_18271,N_12612,N_14166);
or U18272 (N_18272,N_12533,N_14355);
or U18273 (N_18273,N_12131,N_14623);
or U18274 (N_18274,N_16053,N_16813);
nor U18275 (N_18275,N_13023,N_15502);
nand U18276 (N_18276,N_15096,N_12876);
nand U18277 (N_18277,N_14908,N_12395);
nand U18278 (N_18278,N_13484,N_15046);
nand U18279 (N_18279,N_15422,N_12436);
nor U18280 (N_18280,N_16546,N_12166);
nor U18281 (N_18281,N_12095,N_13474);
and U18282 (N_18282,N_13850,N_15626);
nor U18283 (N_18283,N_15711,N_14619);
nor U18284 (N_18284,N_14109,N_16874);
and U18285 (N_18285,N_12011,N_13059);
xnor U18286 (N_18286,N_15620,N_12641);
and U18287 (N_18287,N_12158,N_15652);
xnor U18288 (N_18288,N_15969,N_17186);
xor U18289 (N_18289,N_15418,N_16456);
nand U18290 (N_18290,N_15185,N_16014);
nor U18291 (N_18291,N_12308,N_12300);
and U18292 (N_18292,N_12639,N_16049);
and U18293 (N_18293,N_17553,N_16491);
nor U18294 (N_18294,N_12662,N_13438);
nor U18295 (N_18295,N_16944,N_14673);
nor U18296 (N_18296,N_15224,N_15802);
or U18297 (N_18297,N_12362,N_15767);
nor U18298 (N_18298,N_13779,N_13656);
or U18299 (N_18299,N_15459,N_15998);
and U18300 (N_18300,N_12566,N_13920);
nand U18301 (N_18301,N_13176,N_13577);
nor U18302 (N_18302,N_15643,N_13245);
nor U18303 (N_18303,N_14328,N_16383);
nand U18304 (N_18304,N_15010,N_13191);
nor U18305 (N_18305,N_13152,N_14050);
nand U18306 (N_18306,N_12685,N_16270);
nor U18307 (N_18307,N_14666,N_15729);
or U18308 (N_18308,N_13525,N_16616);
nand U18309 (N_18309,N_15409,N_17391);
nand U18310 (N_18310,N_16422,N_14088);
xor U18311 (N_18311,N_15858,N_17011);
nand U18312 (N_18312,N_17863,N_14524);
nand U18313 (N_18313,N_17133,N_15734);
nand U18314 (N_18314,N_16815,N_13031);
nor U18315 (N_18315,N_17355,N_12645);
and U18316 (N_18316,N_15053,N_15072);
or U18317 (N_18317,N_17837,N_14641);
or U18318 (N_18318,N_13776,N_15306);
nand U18319 (N_18319,N_13935,N_12528);
xor U18320 (N_18320,N_16074,N_13793);
nand U18321 (N_18321,N_13324,N_16357);
nor U18322 (N_18322,N_15317,N_13410);
xnor U18323 (N_18323,N_15226,N_17216);
nor U18324 (N_18324,N_12144,N_14091);
and U18325 (N_18325,N_14221,N_15904);
nand U18326 (N_18326,N_17487,N_12214);
or U18327 (N_18327,N_15549,N_15692);
or U18328 (N_18328,N_12147,N_17864);
nand U18329 (N_18329,N_15017,N_15141);
nor U18330 (N_18330,N_12261,N_16249);
or U18331 (N_18331,N_16583,N_15843);
nand U18332 (N_18332,N_15443,N_12212);
and U18333 (N_18333,N_17070,N_15521);
nor U18334 (N_18334,N_14428,N_16879);
nor U18335 (N_18335,N_12758,N_17542);
nor U18336 (N_18336,N_14304,N_15546);
or U18337 (N_18337,N_13377,N_15806);
or U18338 (N_18338,N_17604,N_16811);
nand U18339 (N_18339,N_14612,N_12476);
xor U18340 (N_18340,N_13208,N_17643);
and U18341 (N_18341,N_13925,N_16355);
nand U18342 (N_18342,N_15302,N_14756);
or U18343 (N_18343,N_14914,N_16710);
or U18344 (N_18344,N_13570,N_16130);
and U18345 (N_18345,N_17911,N_17388);
and U18346 (N_18346,N_14389,N_17292);
or U18347 (N_18347,N_16466,N_15908);
or U18348 (N_18348,N_15523,N_13802);
nor U18349 (N_18349,N_12282,N_14668);
and U18350 (N_18350,N_17949,N_16624);
nand U18351 (N_18351,N_16561,N_12013);
nor U18352 (N_18352,N_17968,N_17482);
nor U18353 (N_18353,N_14063,N_13163);
nor U18354 (N_18354,N_12063,N_17306);
or U18355 (N_18355,N_14646,N_12289);
xor U18356 (N_18356,N_15145,N_13643);
xor U18357 (N_18357,N_15559,N_14642);
nand U18358 (N_18358,N_16920,N_16488);
nand U18359 (N_18359,N_15389,N_17072);
nor U18360 (N_18360,N_16108,N_16237);
or U18361 (N_18361,N_14421,N_13113);
nand U18362 (N_18362,N_16097,N_14185);
xor U18363 (N_18363,N_14116,N_15484);
nand U18364 (N_18364,N_15837,N_15577);
nand U18365 (N_18365,N_16882,N_14725);
or U18366 (N_18366,N_12717,N_15686);
nor U18367 (N_18367,N_13017,N_12456);
or U18368 (N_18368,N_12152,N_16613);
or U18369 (N_18369,N_13403,N_12500);
nor U18370 (N_18370,N_16235,N_15726);
and U18371 (N_18371,N_13344,N_16638);
nand U18372 (N_18372,N_13866,N_17117);
and U18373 (N_18373,N_12659,N_15923);
and U18374 (N_18374,N_12295,N_17853);
or U18375 (N_18375,N_14147,N_12139);
nand U18376 (N_18376,N_15200,N_17879);
nor U18377 (N_18377,N_15928,N_17916);
nand U18378 (N_18378,N_14437,N_15586);
or U18379 (N_18379,N_14346,N_12516);
or U18380 (N_18380,N_17446,N_16415);
and U18381 (N_18381,N_15170,N_17929);
and U18382 (N_18382,N_17061,N_12303);
and U18383 (N_18383,N_15685,N_16642);
and U18384 (N_18384,N_17595,N_16895);
nand U18385 (N_18385,N_13628,N_15981);
nand U18386 (N_18386,N_16927,N_17875);
nand U18387 (N_18387,N_15449,N_14386);
and U18388 (N_18388,N_13302,N_14354);
nand U18389 (N_18389,N_16596,N_12724);
or U18390 (N_18390,N_16791,N_12322);
nand U18391 (N_18391,N_16390,N_16670);
nand U18392 (N_18392,N_13215,N_13966);
xor U18393 (N_18393,N_17180,N_13625);
nand U18394 (N_18394,N_17283,N_16993);
xor U18395 (N_18395,N_12077,N_14575);
and U18396 (N_18396,N_16540,N_16408);
nor U18397 (N_18397,N_17183,N_17285);
nor U18398 (N_18398,N_14089,N_14001);
or U18399 (N_18399,N_14552,N_15225);
or U18400 (N_18400,N_12067,N_16551);
nor U18401 (N_18401,N_16726,N_14923);
or U18402 (N_18402,N_17430,N_15047);
and U18403 (N_18403,N_16119,N_15247);
or U18404 (N_18404,N_14989,N_15616);
or U18405 (N_18405,N_17237,N_12783);
nor U18406 (N_18406,N_14830,N_15093);
and U18407 (N_18407,N_12870,N_14459);
xnor U18408 (N_18408,N_15606,N_16389);
or U18409 (N_18409,N_13013,N_15633);
and U18410 (N_18410,N_17049,N_15656);
nand U18411 (N_18411,N_13477,N_13797);
nand U18412 (N_18412,N_17662,N_12976);
and U18413 (N_18413,N_12799,N_14076);
nor U18414 (N_18414,N_12179,N_14541);
nor U18415 (N_18415,N_16280,N_12149);
and U18416 (N_18416,N_13198,N_13864);
nor U18417 (N_18417,N_14519,N_14560);
nand U18418 (N_18418,N_12843,N_13018);
nor U18419 (N_18419,N_16406,N_14082);
nor U18420 (N_18420,N_16457,N_12966);
nand U18421 (N_18421,N_16822,N_17611);
and U18422 (N_18422,N_16196,N_14413);
or U18423 (N_18423,N_16515,N_17690);
and U18424 (N_18424,N_16537,N_12079);
nor U18425 (N_18425,N_15780,N_16434);
xnor U18426 (N_18426,N_17042,N_14456);
nand U18427 (N_18427,N_15207,N_17019);
or U18428 (N_18428,N_17829,N_13977);
and U18429 (N_18429,N_15634,N_17067);
nor U18430 (N_18430,N_13241,N_15006);
nor U18431 (N_18431,N_16331,N_16891);
nand U18432 (N_18432,N_12816,N_13346);
and U18433 (N_18433,N_14471,N_13370);
and U18434 (N_18434,N_12688,N_12156);
nor U18435 (N_18435,N_14173,N_12199);
or U18436 (N_18436,N_16794,N_13739);
xnor U18437 (N_18437,N_12834,N_12352);
and U18438 (N_18438,N_16369,N_13843);
nand U18439 (N_18439,N_16122,N_14985);
nor U18440 (N_18440,N_14998,N_17955);
and U18441 (N_18441,N_12693,N_12651);
and U18442 (N_18442,N_15036,N_14904);
or U18443 (N_18443,N_12907,N_14286);
nor U18444 (N_18444,N_16547,N_12066);
nand U18445 (N_18445,N_15698,N_13406);
or U18446 (N_18446,N_17100,N_16582);
nor U18447 (N_18447,N_14293,N_12803);
nor U18448 (N_18448,N_16386,N_17245);
nand U18449 (N_18449,N_13732,N_16632);
nand U18450 (N_18450,N_15084,N_17036);
and U18451 (N_18451,N_12005,N_17531);
xnor U18452 (N_18452,N_12429,N_15105);
nor U18453 (N_18453,N_14754,N_15794);
nand U18454 (N_18454,N_17372,N_15610);
nor U18455 (N_18455,N_14994,N_13854);
and U18456 (N_18456,N_12371,N_15974);
nor U18457 (N_18457,N_17975,N_15763);
nand U18458 (N_18458,N_15540,N_12080);
and U18459 (N_18459,N_15550,N_17481);
nand U18460 (N_18460,N_16605,N_13243);
nand U18461 (N_18461,N_15862,N_17597);
nand U18462 (N_18462,N_12102,N_12828);
nor U18463 (N_18463,N_16486,N_13865);
and U18464 (N_18464,N_17749,N_16166);
nand U18465 (N_18465,N_13358,N_14125);
nand U18466 (N_18466,N_14555,N_15396);
nand U18467 (N_18467,N_17834,N_13046);
or U18468 (N_18468,N_12634,N_12737);
and U18469 (N_18469,N_14489,N_15677);
and U18470 (N_18470,N_13550,N_13499);
or U18471 (N_18471,N_16203,N_12222);
nor U18472 (N_18472,N_17860,N_12773);
and U18473 (N_18473,N_17993,N_13659);
and U18474 (N_18474,N_14796,N_14534);
and U18475 (N_18475,N_12757,N_12284);
nand U18476 (N_18476,N_15779,N_13899);
nand U18477 (N_18477,N_12374,N_13647);
xnor U18478 (N_18478,N_16233,N_16001);
nor U18479 (N_18479,N_14561,N_13666);
or U18480 (N_18480,N_12251,N_17987);
or U18481 (N_18481,N_17203,N_14336);
nor U18482 (N_18482,N_13679,N_12422);
or U18483 (N_18483,N_16795,N_17704);
or U18484 (N_18484,N_12633,N_13952);
and U18485 (N_18485,N_13291,N_12435);
nor U18486 (N_18486,N_12187,N_15433);
nand U18487 (N_18487,N_13840,N_14996);
and U18488 (N_18488,N_16185,N_12246);
nor U18489 (N_18489,N_17020,N_12782);
or U18490 (N_18490,N_17271,N_13003);
and U18491 (N_18491,N_12990,N_15529);
or U18492 (N_18492,N_14679,N_13881);
or U18493 (N_18493,N_12689,N_16911);
nor U18494 (N_18494,N_14073,N_14556);
or U18495 (N_18495,N_12085,N_13387);
nor U18496 (N_18496,N_17805,N_17405);
and U18497 (N_18497,N_13837,N_14533);
nor U18498 (N_18498,N_17976,N_12649);
nor U18499 (N_18499,N_14827,N_17802);
or U18500 (N_18500,N_15107,N_12298);
and U18501 (N_18501,N_12155,N_13391);
nor U18502 (N_18502,N_14810,N_13872);
and U18503 (N_18503,N_14497,N_12536);
nor U18504 (N_18504,N_16612,N_16169);
and U18505 (N_18505,N_13494,N_13109);
nand U18506 (N_18506,N_17187,N_17686);
nand U18507 (N_18507,N_12751,N_12086);
nor U18508 (N_18508,N_17700,N_15882);
and U18509 (N_18509,N_13224,N_12091);
nand U18510 (N_18510,N_17979,N_14041);
nand U18511 (N_18511,N_14742,N_13708);
xnor U18512 (N_18512,N_13815,N_17716);
xor U18513 (N_18513,N_16716,N_13211);
nor U18514 (N_18514,N_15323,N_16027);
or U18515 (N_18515,N_16692,N_15076);
xnor U18516 (N_18516,N_13268,N_12210);
xor U18517 (N_18517,N_12550,N_13062);
nor U18518 (N_18518,N_14457,N_14981);
or U18519 (N_18519,N_13347,N_17599);
and U18520 (N_18520,N_12969,N_17053);
xor U18521 (N_18521,N_17074,N_15514);
nor U18522 (N_18522,N_12857,N_14394);
xnor U18523 (N_18523,N_14430,N_16304);
nand U18524 (N_18524,N_12411,N_17087);
nand U18525 (N_18525,N_15768,N_16857);
nand U18526 (N_18526,N_13076,N_17732);
xor U18527 (N_18527,N_17620,N_17688);
or U18528 (N_18528,N_15004,N_16478);
nand U18529 (N_18529,N_16697,N_15778);
nand U18530 (N_18530,N_17554,N_14915);
and U18531 (N_18531,N_15408,N_14512);
and U18532 (N_18532,N_17429,N_17939);
or U18533 (N_18533,N_14593,N_17343);
and U18534 (N_18534,N_16824,N_16392);
and U18535 (N_18535,N_12389,N_15087);
nand U18536 (N_18536,N_14767,N_14023);
nand U18537 (N_18537,N_12485,N_15678);
nand U18538 (N_18538,N_17326,N_12548);
and U18539 (N_18539,N_16352,N_14771);
xor U18540 (N_18540,N_12355,N_12442);
or U18541 (N_18541,N_12878,N_16089);
nand U18542 (N_18542,N_14490,N_13832);
and U18543 (N_18543,N_13437,N_14284);
xor U18544 (N_18544,N_12075,N_13829);
nor U18545 (N_18545,N_13326,N_15576);
or U18546 (N_18546,N_14862,N_15863);
and U18547 (N_18547,N_17985,N_13632);
and U18548 (N_18548,N_15018,N_15903);
or U18549 (N_18549,N_14053,N_16136);
or U18550 (N_18550,N_14093,N_16133);
or U18551 (N_18551,N_16229,N_13890);
nand U18552 (N_18552,N_12697,N_16572);
nor U18553 (N_18553,N_13650,N_16943);
nor U18554 (N_18554,N_14925,N_14898);
nand U18555 (N_18555,N_12960,N_16776);
nand U18556 (N_18556,N_13449,N_17105);
xor U18557 (N_18557,N_15841,N_12819);
or U18558 (N_18558,N_13261,N_14786);
and U18559 (N_18559,N_15483,N_14329);
xnor U18560 (N_18560,N_14320,N_12291);
xor U18561 (N_18561,N_13945,N_15447);
nand U18562 (N_18562,N_17764,N_16306);
or U18563 (N_18563,N_17622,N_16214);
nor U18564 (N_18564,N_12087,N_16854);
and U18565 (N_18565,N_17274,N_17443);
nor U18566 (N_18566,N_13953,N_15759);
and U18567 (N_18567,N_16036,N_14854);
nand U18568 (N_18568,N_13758,N_13857);
and U18569 (N_18569,N_13757,N_14058);
or U18570 (N_18570,N_13773,N_14880);
xor U18571 (N_18571,N_16526,N_17135);
nand U18572 (N_18572,N_17498,N_14710);
nand U18573 (N_18573,N_16645,N_16184);
and U18574 (N_18574,N_15872,N_16370);
nor U18575 (N_18575,N_16319,N_14258);
and U18576 (N_18576,N_17473,N_14918);
and U18577 (N_18577,N_16153,N_15809);
nand U18578 (N_18578,N_14482,N_16539);
and U18579 (N_18579,N_14038,N_12807);
and U18580 (N_18580,N_13670,N_17653);
and U18581 (N_18581,N_16731,N_12307);
nand U18582 (N_18582,N_15313,N_13587);
nor U18583 (N_18583,N_13595,N_17027);
nand U18584 (N_18584,N_16361,N_14470);
nand U18585 (N_18585,N_13690,N_14966);
nand U18586 (N_18586,N_17401,N_13338);
or U18587 (N_18587,N_12423,N_16992);
or U18588 (N_18588,N_17610,N_13523);
and U18589 (N_18589,N_17472,N_16711);
or U18590 (N_18590,N_15614,N_16808);
and U18591 (N_18591,N_15687,N_14779);
and U18592 (N_18592,N_17337,N_16030);
or U18593 (N_18593,N_13819,N_12660);
and U18594 (N_18594,N_17891,N_14648);
xor U18595 (N_18595,N_13482,N_13196);
or U18596 (N_18596,N_14866,N_14037);
nor U18597 (N_18597,N_15844,N_16251);
and U18598 (N_18598,N_17305,N_13547);
and U18599 (N_18599,N_17856,N_13296);
nand U18600 (N_18600,N_13914,N_12440);
nor U18601 (N_18601,N_17568,N_13902);
xor U18602 (N_18602,N_17735,N_13166);
nand U18603 (N_18603,N_14877,N_15617);
and U18604 (N_18604,N_14223,N_16707);
nand U18605 (N_18605,N_12761,N_14620);
nand U18606 (N_18606,N_12126,N_17219);
or U18607 (N_18607,N_12949,N_15619);
nor U18608 (N_18608,N_15063,N_15353);
and U18609 (N_18609,N_15789,N_13727);
nand U18610 (N_18610,N_14323,N_14714);
or U18611 (N_18611,N_14148,N_14036);
and U18612 (N_18612,N_16472,N_14585);
nand U18613 (N_18613,N_15542,N_12302);
nor U18614 (N_18614,N_14034,N_13488);
nor U18615 (N_18615,N_12759,N_16064);
nand U18616 (N_18616,N_14179,N_17458);
nand U18617 (N_18617,N_17692,N_16267);
and U18618 (N_18618,N_15562,N_12044);
or U18619 (N_18619,N_12571,N_13427);
xor U18620 (N_18620,N_14468,N_16865);
nand U18621 (N_18621,N_12998,N_16528);
nor U18622 (N_18622,N_14683,N_13022);
and U18623 (N_18623,N_13042,N_14347);
or U18624 (N_18624,N_17747,N_13000);
and U18625 (N_18625,N_14883,N_17176);
nor U18626 (N_18626,N_14057,N_15384);
nor U18627 (N_18627,N_13939,N_13320);
or U18628 (N_18628,N_16241,N_14257);
nor U18629 (N_18629,N_12554,N_14043);
or U18630 (N_18630,N_13630,N_17232);
nor U18631 (N_18631,N_15828,N_13390);
or U18632 (N_18632,N_13972,N_17782);
or U18633 (N_18633,N_13520,N_15320);
or U18634 (N_18634,N_14922,N_16312);
or U18635 (N_18635,N_12716,N_13195);
nand U18636 (N_18636,N_16285,N_17957);
or U18637 (N_18637,N_16827,N_16598);
nand U18638 (N_18638,N_12804,N_16079);
nor U18639 (N_18639,N_17589,N_16483);
nor U18640 (N_18640,N_12078,N_13172);
nor U18641 (N_18641,N_14713,N_16482);
nand U18642 (N_18642,N_16418,N_16398);
or U18643 (N_18643,N_16842,N_16929);
nor U18644 (N_18644,N_15378,N_14791);
or U18645 (N_18645,N_12262,N_15522);
nand U18646 (N_18646,N_12268,N_14124);
nor U18647 (N_18647,N_14491,N_17852);
nor U18648 (N_18648,N_13784,N_14418);
nor U18649 (N_18649,N_12082,N_16378);
xor U18650 (N_18650,N_16164,N_15563);
nand U18651 (N_18651,N_15274,N_14162);
and U18652 (N_18652,N_16615,N_14643);
nand U18653 (N_18653,N_12963,N_12908);
and U18654 (N_18654,N_13069,N_17028);
and U18655 (N_18655,N_15720,N_14792);
nor U18656 (N_18656,N_14755,N_12658);
nand U18657 (N_18657,N_14398,N_15039);
nor U18658 (N_18658,N_15412,N_15582);
or U18659 (N_18659,N_15653,N_16946);
and U18660 (N_18660,N_14460,N_17193);
nand U18661 (N_18661,N_16178,N_12902);
or U18662 (N_18662,N_12206,N_15089);
or U18663 (N_18663,N_14950,N_15503);
or U18664 (N_18664,N_15106,N_15428);
xnor U18665 (N_18665,N_12356,N_15737);
and U18666 (N_18666,N_15910,N_15061);
nand U18667 (N_18667,N_12271,N_13325);
and U18668 (N_18668,N_13589,N_15211);
xor U18669 (N_18669,N_17632,N_12984);
xnor U18670 (N_18670,N_13409,N_17880);
nor U18671 (N_18671,N_14267,N_12970);
nor U18672 (N_18672,N_17761,N_12183);
or U18673 (N_18673,N_14480,N_12572);
nand U18674 (N_18674,N_14858,N_15324);
and U18675 (N_18675,N_12987,N_17517);
xnor U18676 (N_18676,N_16444,N_13824);
and U18677 (N_18677,N_12345,N_13394);
nand U18678 (N_18678,N_12584,N_13859);
nor U18679 (N_18679,N_17363,N_12630);
or U18680 (N_18680,N_15929,N_12709);
xnor U18681 (N_18681,N_16450,N_13713);
and U18682 (N_18682,N_13143,N_13894);
nor U18683 (N_18683,N_16843,N_15719);
or U18684 (N_18684,N_12655,N_13551);
and U18685 (N_18685,N_16758,N_12197);
and U18686 (N_18686,N_15801,N_13168);
or U18687 (N_18687,N_16661,N_13617);
nor U18688 (N_18688,N_12218,N_16128);
or U18689 (N_18689,N_17808,N_16004);
or U18690 (N_18690,N_14795,N_14357);
nand U18691 (N_18691,N_16755,N_12927);
nor U18692 (N_18692,N_13600,N_15395);
or U18693 (N_18693,N_12292,N_12933);
or U18694 (N_18694,N_14448,N_17395);
or U18695 (N_18695,N_14392,N_13909);
and U18696 (N_18696,N_16330,N_12244);
nor U18697 (N_18697,N_14263,N_15826);
xor U18698 (N_18698,N_15917,N_14711);
nor U18699 (N_18699,N_17780,N_17967);
nand U18700 (N_18700,N_13559,N_14201);
nand U18701 (N_18701,N_17172,N_12712);
nor U18702 (N_18702,N_16573,N_14213);
nor U18703 (N_18703,N_17511,N_14404);
nor U18704 (N_18704,N_15758,N_17421);
xor U18705 (N_18705,N_17131,N_12238);
and U18706 (N_18706,N_13631,N_13724);
nand U18707 (N_18707,N_16363,N_14743);
nand U18708 (N_18708,N_12388,N_14651);
or U18709 (N_18709,N_13099,N_12668);
nor U18710 (N_18710,N_16407,N_12019);
or U18711 (N_18711,N_16362,N_15623);
nand U18712 (N_18712,N_16496,N_12314);
and U18713 (N_18713,N_13469,N_17198);
nor U18714 (N_18714,N_17640,N_17269);
nand U18715 (N_18715,N_13980,N_15136);
nand U18716 (N_18716,N_14352,N_17406);
nand U18717 (N_18717,N_13074,N_14044);
or U18718 (N_18718,N_12979,N_12454);
nor U18719 (N_18719,N_14407,N_13738);
or U18720 (N_18720,N_13505,N_14537);
or U18721 (N_18721,N_15078,N_17898);
and U18722 (N_18722,N_17339,N_16402);
nor U18723 (N_18723,N_16225,N_17286);
nor U18724 (N_18724,N_13436,N_14272);
or U18725 (N_18725,N_16949,N_12638);
nor U18726 (N_18726,N_13816,N_14403);
nor U18727 (N_18727,N_16956,N_12130);
nor U18728 (N_18728,N_17845,N_12701);
xor U18729 (N_18729,N_17787,N_14054);
nand U18730 (N_18730,N_17712,N_15899);
or U18731 (N_18731,N_15194,N_15769);
nand U18732 (N_18732,N_14824,N_16078);
nor U18733 (N_18733,N_12499,N_13392);
nor U18734 (N_18734,N_13800,N_13927);
and U18735 (N_18735,N_15424,N_17857);
nor U18736 (N_18736,N_17687,N_17008);
nor U18737 (N_18737,N_17365,N_12943);
nand U18738 (N_18738,N_15962,N_13297);
nand U18739 (N_18739,N_14262,N_14543);
nor U18740 (N_18740,N_15173,N_16618);
nor U18741 (N_18741,N_14205,N_14587);
and U18742 (N_18742,N_12209,N_14960);
nand U18743 (N_18743,N_14061,N_13274);
nor U18744 (N_18744,N_17442,N_13491);
and U18745 (N_18745,N_16563,N_14180);
or U18746 (N_18746,N_17223,N_15888);
nand U18747 (N_18747,N_17159,N_15399);
or U18748 (N_18748,N_12480,N_14074);
and U18749 (N_18749,N_12860,N_16550);
and U18750 (N_18750,N_14530,N_15895);
and U18751 (N_18751,N_15961,N_13340);
xor U18752 (N_18752,N_12363,N_17928);
and U18753 (N_18753,N_17119,N_14123);
and U18754 (N_18754,N_17084,N_13424);
nand U18755 (N_18755,N_12400,N_14065);
nand U18756 (N_18756,N_16562,N_16190);
and U18757 (N_18757,N_12620,N_16947);
and U18758 (N_18758,N_12243,N_17024);
or U18759 (N_18759,N_15539,N_14532);
nand U18760 (N_18760,N_13267,N_13244);
or U18761 (N_18761,N_16889,N_12004);
nand U18762 (N_18762,N_16151,N_13153);
or U18763 (N_18763,N_16866,N_13956);
nand U18764 (N_18764,N_15642,N_14464);
and U18765 (N_18765,N_13810,N_12211);
or U18766 (N_18766,N_15884,N_16852);
and U18767 (N_18767,N_14505,N_13246);
and U18768 (N_18768,N_17076,N_12189);
nand U18769 (N_18769,N_14029,N_16982);
nand U18770 (N_18770,N_12378,N_12273);
xor U18771 (N_18771,N_17806,N_12530);
nand U18772 (N_18772,N_16168,N_14280);
nand U18773 (N_18773,N_16595,N_17630);
or U18774 (N_18774,N_14798,N_17660);
nand U18775 (N_18775,N_15544,N_17476);
xor U18776 (N_18776,N_13950,N_15516);
nand U18777 (N_18777,N_12171,N_13983);
nand U18778 (N_18778,N_17428,N_16431);
nand U18779 (N_18779,N_15897,N_15533);
or U18780 (N_18780,N_17798,N_14245);
nor U18781 (N_18781,N_15868,N_13286);
xnor U18782 (N_18782,N_15257,N_15597);
nor U18783 (N_18783,N_16643,N_16120);
nand U18784 (N_18784,N_15989,N_12252);
nor U18785 (N_18785,N_12039,N_16181);
and U18786 (N_18786,N_16328,N_16264);
and U18787 (N_18787,N_15552,N_15358);
and U18788 (N_18788,N_17394,N_15281);
and U18789 (N_18789,N_12993,N_13272);
or U18790 (N_18790,N_17515,N_17433);
xnor U18791 (N_18791,N_16193,N_14746);
nand U18792 (N_18792,N_12236,N_16096);
nor U18793 (N_18793,N_15016,N_13728);
nand U18794 (N_18794,N_12967,N_17386);
nand U18795 (N_18795,N_16845,N_13140);
nor U18796 (N_18796,N_16729,N_14697);
xor U18797 (N_18797,N_16673,N_12811);
nand U18798 (N_18798,N_15596,N_14976);
nor U18799 (N_18799,N_14298,N_16340);
and U18800 (N_18800,N_15310,N_17547);
nand U18801 (N_18801,N_17991,N_13202);
and U18802 (N_18802,N_14892,N_16910);
xnor U18803 (N_18803,N_14544,N_12009);
nand U18804 (N_18804,N_12887,N_15290);
xor U18805 (N_18805,N_16082,N_13592);
nand U18806 (N_18806,N_12790,N_12753);
or U18807 (N_18807,N_13665,N_15287);
nor U18808 (N_18808,N_17543,N_14443);
and U18809 (N_18809,N_13989,N_15612);
nand U18810 (N_18810,N_16704,N_16724);
nand U18811 (N_18811,N_14622,N_17007);
and U18812 (N_18812,N_14846,N_13309);
nor U18813 (N_18813,N_13054,N_16644);
and U18814 (N_18814,N_12945,N_16353);
or U18815 (N_18815,N_17021,N_12695);
or U18816 (N_18816,N_16375,N_14232);
xnor U18817 (N_18817,N_13306,N_14548);
or U18818 (N_18818,N_12168,N_13342);
xnor U18819 (N_18819,N_16259,N_12100);
nor U18820 (N_18820,N_16380,N_13811);
xnor U18821 (N_18821,N_17488,N_16611);
xor U18822 (N_18822,N_12768,N_13642);
or U18823 (N_18823,N_16584,N_13487);
nand U18824 (N_18824,N_15792,N_12714);
and U18825 (N_18825,N_16625,N_17912);
xnor U18826 (N_18826,N_13591,N_15383);
or U18827 (N_18827,N_16394,N_13503);
xor U18828 (N_18828,N_17423,N_12789);
nand U18829 (N_18829,N_13451,N_15337);
nor U18830 (N_18830,N_15023,N_16525);
nor U18831 (N_18831,N_12607,N_14106);
and U18832 (N_18832,N_12275,N_15942);
xnor U18833 (N_18833,N_14069,N_15641);
and U18834 (N_18834,N_12784,N_14579);
and U18835 (N_18835,N_14715,N_17821);
nor U18836 (N_18836,N_17086,N_17085);
nand U18837 (N_18837,N_15398,N_12827);
nor U18838 (N_18838,N_16928,N_17057);
nor U18839 (N_18839,N_17419,N_13770);
nor U18840 (N_18840,N_12178,N_14856);
nor U18841 (N_18841,N_12376,N_15595);
xor U18842 (N_18842,N_17147,N_13001);
and U18843 (N_18843,N_12959,N_15867);
nand U18844 (N_18844,N_13748,N_17437);
xnor U18845 (N_18845,N_16480,N_14144);
nand U18846 (N_18846,N_13608,N_14446);
and U18847 (N_18847,N_13601,N_13043);
nor U18848 (N_18848,N_16016,N_14252);
and U18849 (N_18849,N_14420,N_12367);
nand U18850 (N_18850,N_15976,N_13958);
and U18851 (N_18851,N_15456,N_13480);
or U18852 (N_18852,N_15289,N_12049);
nor U18853 (N_18853,N_16485,N_14844);
and U18854 (N_18854,N_15952,N_13968);
xnor U18855 (N_18855,N_16713,N_13682);
and U18856 (N_18856,N_14338,N_17616);
nand U18857 (N_18857,N_13855,N_17126);
or U18858 (N_18858,N_12366,N_17907);
nand U18859 (N_18859,N_12003,N_12956);
xor U18860 (N_18860,N_16391,N_12491);
xor U18861 (N_18861,N_15104,N_12327);
nand U18862 (N_18862,N_17789,N_14935);
nor U18863 (N_18863,N_14014,N_17346);
nor U18864 (N_18864,N_15057,N_14465);
nor U18865 (N_18865,N_17973,N_12397);
and U18866 (N_18866,N_12092,N_14385);
nor U18867 (N_18867,N_14805,N_12176);
and U18868 (N_18868,N_16860,N_16656);
xnor U18869 (N_18869,N_15163,N_15508);
nor U18870 (N_18870,N_14492,N_13723);
and U18871 (N_18871,N_13557,N_17158);
and U18872 (N_18872,N_13217,N_14748);
nor U18873 (N_18873,N_12889,N_12793);
nor U18874 (N_18874,N_14559,N_13135);
or U18875 (N_18875,N_16043,N_14817);
or U18876 (N_18876,N_15752,N_12200);
and U18877 (N_18877,N_17521,N_13237);
nor U18878 (N_18878,N_14822,N_16735);
or U18879 (N_18879,N_17956,N_15538);
and U18880 (N_18880,N_16696,N_16103);
nor U18881 (N_18881,N_15133,N_15406);
xor U18882 (N_18882,N_15773,N_13334);
and U18883 (N_18883,N_17279,N_13313);
nand U18884 (N_18884,N_15102,N_16737);
nand U18885 (N_18885,N_16913,N_12495);
nor U18886 (N_18886,N_14160,N_16989);
or U18887 (N_18887,N_17954,N_15501);
or U18888 (N_18888,N_16112,N_16440);
and U18889 (N_18889,N_12950,N_14807);
and U18890 (N_18890,N_13906,N_17483);
nand U18891 (N_18891,N_14849,N_14882);
or U18892 (N_18892,N_12022,N_12637);
nor U18893 (N_18893,N_17265,N_14449);
nor U18894 (N_18894,N_14301,N_16207);
or U18895 (N_18895,N_14563,N_12774);
xnor U18896 (N_18896,N_17900,N_12233);
and U18897 (N_18897,N_17592,N_14939);
nand U18898 (N_18898,N_16796,N_16627);
and U18899 (N_18899,N_17567,N_12276);
or U18900 (N_18900,N_17862,N_17023);
xor U18901 (N_18901,N_15787,N_17095);
nor U18902 (N_18902,N_12646,N_16347);
and U18903 (N_18903,N_14583,N_17445);
nand U18904 (N_18904,N_14538,N_12871);
nand U18905 (N_18905,N_13740,N_17001);
nand U18906 (N_18906,N_17697,N_17508);
and U18907 (N_18907,N_13579,N_15697);
or U18908 (N_18908,N_14677,N_12923);
nor U18909 (N_18909,N_15253,N_12564);
xnor U18910 (N_18910,N_13814,N_12110);
and U18911 (N_18911,N_15264,N_13842);
or U18912 (N_18912,N_16455,N_15944);
and U18913 (N_18913,N_15548,N_15745);
or U18914 (N_18914,N_16607,N_13010);
nor U18915 (N_18915,N_16519,N_13429);
or U18916 (N_18916,N_13689,N_14937);
and U18917 (N_18917,N_12690,N_16806);
xnor U18918 (N_18918,N_13283,N_14721);
nor U18919 (N_18919,N_15382,N_14961);
nand U18920 (N_18920,N_16970,N_17083);
nor U18921 (N_18921,N_12242,N_12557);
xnor U18922 (N_18922,N_14953,N_17783);
and U18923 (N_18923,N_14876,N_15113);
nor U18924 (N_18924,N_14984,N_17464);
or U18925 (N_18925,N_16248,N_17146);
and U18926 (N_18926,N_13035,N_14569);
and U18927 (N_18927,N_12502,N_13122);
or U18928 (N_18928,N_14291,N_14749);
nand U18929 (N_18929,N_12301,N_14433);
and U18930 (N_18930,N_16084,N_15419);
nand U18931 (N_18931,N_14956,N_13709);
nor U18932 (N_18932,N_13919,N_15182);
nand U18933 (N_18933,N_16687,N_14655);
xnor U18934 (N_18934,N_12123,N_14706);
and U18935 (N_18935,N_16532,N_12361);
xor U18936 (N_18936,N_13834,N_15015);
xor U18937 (N_18937,N_13075,N_17951);
and U18938 (N_18938,N_17148,N_14042);
xor U18939 (N_18939,N_14726,N_14134);
nor U18940 (N_18940,N_12228,N_16890);
nand U18941 (N_18941,N_16684,N_12452);
or U18942 (N_18942,N_16760,N_16152);
or U18943 (N_18943,N_15551,N_15286);
nand U18944 (N_18944,N_17545,N_14294);
nand U18945 (N_18945,N_13351,N_14776);
or U18946 (N_18946,N_16442,N_17776);
nor U18947 (N_18947,N_16177,N_16792);
nor U18948 (N_18948,N_17489,N_14207);
or U18949 (N_18949,N_16599,N_12103);
nor U18950 (N_18950,N_15360,N_13024);
xnor U18951 (N_18951,N_16065,N_13025);
nor U18952 (N_18952,N_12839,N_15118);
nor U18953 (N_18953,N_14122,N_15080);
nand U18954 (N_18954,N_16470,N_15602);
and U18955 (N_18955,N_16162,N_15589);
nor U18956 (N_18956,N_15811,N_12002);
nor U18957 (N_18957,N_17277,N_13521);
nor U18958 (N_18958,N_12734,N_16017);
or U18959 (N_18959,N_17613,N_15584);
nor U18960 (N_18960,N_13142,N_15982);
nor U18961 (N_18961,N_16100,N_15050);
or U18962 (N_18962,N_13856,N_13470);
nand U18963 (N_18963,N_16848,N_12278);
and U18964 (N_18964,N_12119,N_15122);
and U18965 (N_18965,N_15519,N_12297);
nor U18966 (N_18966,N_17519,N_13073);
or U18967 (N_18967,N_13457,N_15407);
nand U18968 (N_18968,N_12906,N_14071);
and U18969 (N_18969,N_15322,N_17417);
nor U18970 (N_18970,N_13675,N_12140);
and U18971 (N_18971,N_14924,N_15355);
nand U18972 (N_18972,N_15713,N_17373);
xor U18973 (N_18973,N_16454,N_16853);
and U18974 (N_18974,N_16230,N_12593);
nand U18975 (N_18975,N_15201,N_12647);
nor U18976 (N_18976,N_13008,N_13485);
xnor U18977 (N_18977,N_16554,N_12328);
and U18978 (N_18978,N_13948,N_17636);
xor U18979 (N_18979,N_12657,N_17859);
nand U18980 (N_18980,N_15886,N_13991);
nand U18981 (N_18981,N_13677,N_13156);
nor U18982 (N_18982,N_14075,N_17318);
or U18983 (N_18983,N_15696,N_13988);
or U18984 (N_18984,N_12190,N_13846);
nor U18985 (N_18985,N_14194,N_12160);
or U18986 (N_18986,N_14777,N_17002);
nor U18987 (N_18987,N_13301,N_14540);
nand U18988 (N_18988,N_15128,N_17034);
or U18989 (N_18989,N_14349,N_13721);
or U18990 (N_18990,N_14977,N_17969);
and U18991 (N_18991,N_16753,N_16850);
nor U18992 (N_18992,N_13085,N_17721);
and U18993 (N_18993,N_15968,N_14429);
or U18994 (N_18994,N_14903,N_13165);
and U18995 (N_18995,N_14900,N_14744);
nand U18996 (N_18996,N_16295,N_16182);
nand U18997 (N_18997,N_13048,N_14064);
or U18998 (N_18998,N_16183,N_14604);
or U18999 (N_18999,N_14803,N_14508);
and U19000 (N_19000,N_17257,N_13125);
and U19001 (N_19001,N_15444,N_13498);
and U19002 (N_19002,N_15977,N_14751);
nor U19003 (N_19003,N_16305,N_16453);
and U19004 (N_19004,N_12749,N_17803);
and U19005 (N_19005,N_12503,N_16500);
and U19006 (N_19006,N_14319,N_12574);
nor U19007 (N_19007,N_15151,N_14476);
nand U19008 (N_19008,N_16080,N_13671);
nor U19009 (N_19009,N_15666,N_14159);
nor U19010 (N_19010,N_14797,N_16066);
xor U19011 (N_19011,N_13335,N_13225);
and U19012 (N_19012,N_13715,N_12915);
xor U19013 (N_19013,N_17762,N_17781);
and U19014 (N_19014,N_12433,N_17921);
or U19015 (N_19015,N_16793,N_15366);
or U19016 (N_19016,N_14672,N_16817);
and U19017 (N_19017,N_17235,N_14982);
and U19018 (N_19018,N_12673,N_13380);
nand U19019 (N_19019,N_14375,N_17865);
nor U19020 (N_19020,N_13290,N_13040);
xnor U19021 (N_19021,N_15915,N_15035);
nand U19022 (N_19022,N_14539,N_12465);
xor U19023 (N_19023,N_13384,N_13839);
xor U19024 (N_19024,N_13164,N_15618);
or U19025 (N_19025,N_14499,N_13414);
and U19026 (N_19026,N_12879,N_16732);
or U19027 (N_19027,N_13431,N_14172);
nor U19028 (N_19028,N_15943,N_13588);
or U19029 (N_19029,N_16050,N_12249);
or U19030 (N_19030,N_15935,N_13571);
or U19031 (N_19031,N_12027,N_15291);
xor U19032 (N_19032,N_12105,N_13475);
nand U19033 (N_19033,N_12490,N_17828);
and U19034 (N_19034,N_16003,N_13039);
nand U19035 (N_19035,N_14078,N_14577);
nor U19036 (N_19036,N_16810,N_12794);
and U19037 (N_19037,N_15566,N_15262);
xor U19038 (N_19038,N_17556,N_16015);
nor U19039 (N_19039,N_16494,N_17451);
or U19040 (N_19040,N_12216,N_17258);
xor U19041 (N_19041,N_17252,N_16658);
xnor U19042 (N_19042,N_13102,N_17858);
nand U19043 (N_19043,N_13913,N_15810);
nand U19044 (N_19044,N_16105,N_12854);
xnor U19045 (N_19045,N_14660,N_12010);
xnor U19046 (N_19046,N_14764,N_16837);
nand U19047 (N_19047,N_17593,N_12569);
or U19048 (N_19048,N_16002,N_14649);
xor U19049 (N_19049,N_16531,N_17233);
and U19050 (N_19050,N_15161,N_13227);
nand U19051 (N_19051,N_16364,N_16620);
nor U19052 (N_19052,N_14259,N_14253);
nand U19053 (N_19053,N_14445,N_17656);
or U19054 (N_19054,N_16146,N_12154);
nand U19055 (N_19055,N_17861,N_17243);
and U19056 (N_19056,N_15624,N_12408);
nor U19057 (N_19057,N_15804,N_16068);
nor U19058 (N_19058,N_15771,N_13500);
xnor U19059 (N_19059,N_14588,N_14974);
nor U19060 (N_19060,N_15511,N_16154);
and U19061 (N_19061,N_15835,N_15718);
nor U19062 (N_19062,N_12245,N_17013);
and U19063 (N_19063,N_14397,N_16764);
or U19064 (N_19064,N_12663,N_17127);
xor U19065 (N_19065,N_16464,N_12996);
nor U19066 (N_19066,N_17585,N_13897);
xnor U19067 (N_19067,N_12116,N_16349);
nor U19068 (N_19068,N_14959,N_12815);
nand U19069 (N_19069,N_14952,N_15933);
xor U19070 (N_19070,N_16819,N_17755);
nor U19071 (N_19071,N_17727,N_16971);
or U19072 (N_19072,N_16452,N_17661);
nor U19073 (N_19073,N_12065,N_12259);
and U19074 (N_19074,N_17195,N_13214);
and U19075 (N_19075,N_12285,N_15282);
and U19076 (N_19076,N_12159,N_14178);
xnor U19077 (N_19077,N_16351,N_14834);
and U19078 (N_19078,N_14440,N_17710);
nor U19079 (N_19079,N_15423,N_12319);
nor U19080 (N_19080,N_15911,N_16802);
nand U19081 (N_19081,N_15203,N_12175);
nor U19082 (N_19082,N_17770,N_15898);
and U19083 (N_19083,N_14969,N_12304);
nor U19084 (N_19084,N_17043,N_17397);
nand U19085 (N_19085,N_13860,N_17794);
or U19086 (N_19086,N_13036,N_15757);
and U19087 (N_19087,N_17479,N_15143);
xnor U19088 (N_19088,N_13756,N_15860);
or U19089 (N_19089,N_15189,N_15919);
and U19090 (N_19090,N_17069,N_15478);
and U19091 (N_19091,N_17125,N_16662);
nand U19092 (N_19092,N_17649,N_12334);
or U19093 (N_19093,N_15833,N_12260);
nor U19094 (N_19094,N_12587,N_12801);
and U19095 (N_19095,N_12330,N_14444);
and U19096 (N_19096,N_15055,N_14236);
nor U19097 (N_19097,N_12665,N_13827);
nand U19098 (N_19098,N_17140,N_15058);
xnor U19099 (N_19099,N_14372,N_16055);
xor U19100 (N_19100,N_15486,N_14200);
and U19101 (N_19101,N_15239,N_15196);
nor U19102 (N_19102,N_16213,N_16106);
and U19103 (N_19103,N_17801,N_12676);
nand U19104 (N_19104,N_12098,N_12399);
and U19105 (N_19105,N_14728,N_13769);
and U19106 (N_19106,N_15655,N_15913);
and U19107 (N_19107,N_16299,N_16985);
nor U19108 (N_19108,N_16736,N_12895);
or U19109 (N_19109,N_17325,N_13308);
nand U19110 (N_19110,N_15228,N_15679);
xor U19111 (N_19111,N_12320,N_12177);
nor U19112 (N_19112,N_13654,N_13786);
and U19113 (N_19113,N_14145,N_12470);
and U19114 (N_19114,N_15150,N_16567);
nand U19115 (N_19115,N_15367,N_13467);
nor U19116 (N_19116,N_14670,N_12652);
or U19117 (N_19117,N_15254,N_14833);
xnor U19118 (N_19118,N_13107,N_17598);
nand U19119 (N_19119,N_13373,N_16557);
or U19120 (N_19120,N_13714,N_12121);
and U19121 (N_19121,N_17234,N_17240);
nor U19122 (N_19122,N_14911,N_13687);
nor U19123 (N_19123,N_14237,N_15840);
xor U19124 (N_19124,N_13928,N_16006);
and U19125 (N_19125,N_15846,N_13145);
and U19126 (N_19126,N_14012,N_12929);
xor U19127 (N_19127,N_14832,N_12611);
or U19128 (N_19128,N_15859,N_16683);
or U19129 (N_19129,N_14736,N_12669);
or U19130 (N_19130,N_17486,N_13987);
or U19131 (N_19131,N_16118,N_13402);
nand U19132 (N_19132,N_16789,N_16291);
nor U19133 (N_19133,N_12401,N_12867);
nor U19134 (N_19134,N_17778,N_17165);
nor U19135 (N_19135,N_16067,N_15580);
and U19136 (N_19136,N_15178,N_17296);
or U19137 (N_19137,N_16159,N_12985);
nand U19138 (N_19138,N_12396,N_14218);
nor U19139 (N_19139,N_13007,N_13955);
xor U19140 (N_19140,N_16396,N_16385);
nor U19141 (N_19141,N_16807,N_13707);
or U19142 (N_19142,N_15749,N_17830);
xor U19143 (N_19143,N_16438,N_13926);
or U19144 (N_19144,N_14171,N_16950);
nor U19145 (N_19145,N_15066,N_14527);
nor U19146 (N_19146,N_13486,N_12510);
and U19147 (N_19147,N_12309,N_17910);
nand U19148 (N_19148,N_12565,N_15246);
or U19149 (N_19149,N_12975,N_12626);
and U19150 (N_19150,N_17218,N_16757);
and U19151 (N_19151,N_17694,N_17530);
or U19152 (N_19152,N_14692,N_16511);
xor U19153 (N_19153,N_14889,N_12340);
xnor U19154 (N_19154,N_16657,N_15531);
nand U19155 (N_19155,N_16520,N_15649);
and U19156 (N_19156,N_16877,N_13408);
nand U19157 (N_19157,N_14967,N_16176);
or U19158 (N_19158,N_15564,N_17438);
or U19159 (N_19159,N_14473,N_16897);
nand U19160 (N_19160,N_14999,N_13456);
nand U19161 (N_19161,N_12730,N_17188);
nand U19162 (N_19162,N_17431,N_12324);
xnor U19163 (N_19163,N_16610,N_16965);
or U19164 (N_19164,N_16722,N_13322);
nor U19165 (N_19165,N_12137,N_16033);
nor U19166 (N_19166,N_15940,N_15142);
nor U19167 (N_19167,N_15466,N_14163);
and U19168 (N_19168,N_14231,N_15077);
and U19169 (N_19169,N_16436,N_14067);
or U19170 (N_19170,N_15064,N_12431);
or U19171 (N_19171,N_15847,N_14202);
nor U19172 (N_19172,N_12654,N_12493);
and U19173 (N_19173,N_12153,N_14990);
nand U19174 (N_19174,N_17672,N_15972);
nand U19175 (N_19175,N_16038,N_16564);
nand U19176 (N_19176,N_12443,N_15183);
and U19177 (N_19177,N_12599,N_12057);
nand U19178 (N_19178,N_15790,N_17938);
xnor U19179 (N_19179,N_16413,N_16192);
or U19180 (N_19180,N_15593,N_17063);
nand U19181 (N_19181,N_12413,N_13371);
nand U19182 (N_19182,N_17619,N_17974);
nand U19183 (N_19183,N_17923,N_17629);
nor U19184 (N_19184,N_14968,N_13978);
xnor U19185 (N_19185,N_17705,N_17617);
and U19186 (N_19186,N_12851,N_13357);
nand U19187 (N_19187,N_16013,N_16847);
or U19188 (N_19188,N_17799,N_14021);
and U19189 (N_19189,N_13777,N_15127);
nand U19190 (N_19190,N_14695,N_15465);
nand U19191 (N_19191,N_14701,N_15164);
nand U19192 (N_19192,N_14864,N_14028);
and U19193 (N_19193,N_12188,N_14196);
xnor U19194 (N_19194,N_17826,N_12434);
nor U19195 (N_19195,N_12263,N_12494);
nor U19196 (N_19196,N_12733,N_12511);
xor U19197 (N_19197,N_16292,N_15878);
nand U19198 (N_19198,N_13121,N_16785);
or U19199 (N_19199,N_17748,N_13032);
nor U19200 (N_19200,N_17925,N_16986);
and U19201 (N_19201,N_14290,N_16126);
nand U19202 (N_19202,N_15431,N_17230);
or U19203 (N_19203,N_15116,N_16109);
and U19204 (N_19204,N_12708,N_16031);
nor U19205 (N_19205,N_16983,N_14917);
nand U19206 (N_19206,N_14279,N_17952);
and U19207 (N_19207,N_16307,N_16980);
nor U19208 (N_19208,N_14062,N_14240);
and U19209 (N_19209,N_17758,N_16150);
or U19210 (N_19210,N_15905,N_12754);
nor U19211 (N_19211,N_17740,N_16712);
nor U19212 (N_19212,N_14599,N_14342);
xnor U19213 (N_19213,N_14667,N_12104);
nor U19214 (N_19214,N_14973,N_14855);
nor U19215 (N_19215,N_14550,N_12012);
or U19216 (N_19216,N_16144,N_14895);
and U19217 (N_19217,N_17924,N_12164);
or U19218 (N_19218,N_14316,N_15248);
nor U19219 (N_19219,N_16377,N_14208);
nand U19220 (N_19220,N_17358,N_15265);
nor U19221 (N_19221,N_15174,N_12964);
nor U19222 (N_19222,N_14860,N_12769);
xor U19223 (N_19223,N_14553,N_12526);
xnor U19224 (N_19224,N_17500,N_17657);
xor U19225 (N_19225,N_12445,N_14885);
nand U19226 (N_19226,N_13067,N_13328);
xnor U19227 (N_19227,N_17272,N_16695);
or U19228 (N_19228,N_15646,N_13459);
and U19229 (N_19229,N_17261,N_16075);
nor U19230 (N_19230,N_12661,N_15400);
and U19231 (N_19231,N_13789,N_14551);
or U19232 (N_19232,N_16941,N_13667);
or U19233 (N_19233,N_14676,N_15494);
nor U19234 (N_19234,N_17637,N_17784);
and U19235 (N_19235,N_15760,N_13086);
and U19236 (N_19236,N_13134,N_12940);
nand U19237 (N_19237,N_12580,N_17302);
xnor U19238 (N_19238,N_13068,N_17963);
or U19239 (N_19239,N_13790,N_16600);
and U19240 (N_19240,N_14453,N_16102);
xnor U19241 (N_19241,N_15572,N_14376);
or U19242 (N_19242,N_16790,N_17908);
and U19243 (N_19243,N_17332,N_12897);
nor U19244 (N_19244,N_15901,N_15329);
and U19245 (N_19245,N_15995,N_17785);
or U19246 (N_19246,N_12394,N_12583);
nor U19247 (N_19247,N_12097,N_17981);
nand U19248 (N_19248,N_12900,N_13087);
nand U19249 (N_19249,N_13576,N_13782);
and U19250 (N_19250,N_16297,N_16262);
and U19251 (N_19251,N_17922,N_13562);
nand U19252 (N_19252,N_14203,N_15825);
or U19253 (N_19253,N_17767,N_17132);
or U19254 (N_19254,N_15838,N_13598);
nand U19255 (N_19255,N_15125,N_12916);
or U19256 (N_19256,N_17854,N_15027);
and U19257 (N_19257,N_12725,N_12847);
nand U19258 (N_19258,N_17503,N_16559);
and U19259 (N_19259,N_13175,N_14432);
nand U19260 (N_19260,N_17060,N_12138);
and U19261 (N_19261,N_13141,N_12899);
or U19262 (N_19262,N_12921,N_13548);
or U19263 (N_19263,N_16421,N_13162);
nand U19264 (N_19264,N_16933,N_12142);
or U19265 (N_19265,N_16886,N_16308);
xor U19266 (N_19266,N_16475,N_12914);
and U19267 (N_19267,N_16289,N_12603);
or U19268 (N_19268,N_16701,N_15764);
or U19269 (N_19269,N_13657,N_12489);
nor U19270 (N_19270,N_15060,N_13892);
xnor U19271 (N_19271,N_13321,N_14921);
or U19272 (N_19272,N_16926,N_13020);
nor U19273 (N_19273,N_16238,N_16451);
nand U19274 (N_19274,N_12896,N_13079);
and U19275 (N_19275,N_17671,N_14377);
nor U19276 (N_19276,N_13300,N_12042);
or U19277 (N_19277,N_17143,N_13812);
or U19278 (N_19278,N_14455,N_17777);
and U19279 (N_19279,N_17614,N_16721);
nand U19280 (N_19280,N_17791,N_17795);
nor U19281 (N_19281,N_17960,N_14017);
or U19282 (N_19282,N_14839,N_13744);
nor U19283 (N_19283,N_17441,N_13645);
xnor U19284 (N_19284,N_12055,N_12888);
nand U19285 (N_19285,N_12602,N_14224);
xor U19286 (N_19286,N_14835,N_15714);
nand U19287 (N_19287,N_12519,N_14566);
or U19288 (N_19288,N_17528,N_15588);
nor U19289 (N_19289,N_17818,N_12258);
or U19290 (N_19290,N_17478,N_14753);
and U19291 (N_19291,N_14315,N_16738);
and U19292 (N_19292,N_15930,N_16411);
and U19293 (N_19293,N_15137,N_16009);
nor U19294 (N_19294,N_12315,N_13177);
and U19295 (N_19295,N_17775,N_12196);
nor U19296 (N_19296,N_17664,N_15223);
or U19297 (N_19297,N_13047,N_15413);
xor U19298 (N_19298,N_17579,N_13269);
nand U19299 (N_19299,N_15232,N_15573);
nand U19300 (N_19300,N_17768,N_16581);
or U19301 (N_19301,N_14308,N_12405);
and U19302 (N_19302,N_13005,N_17178);
xnor U19303 (N_19303,N_13364,N_12604);
and U19304 (N_19304,N_13681,N_17754);
or U19305 (N_19305,N_15031,N_13658);
nor U19306 (N_19306,N_15658,N_13240);
nand U19307 (N_19307,N_12472,N_12846);
nand U19308 (N_19308,N_13841,N_16171);
nand U19309 (N_19309,N_16826,N_16247);
and U19310 (N_19310,N_13629,N_17120);
nor U19311 (N_19311,N_14942,N_16978);
xor U19312 (N_19312,N_17822,N_13618);
or U19313 (N_19313,N_13536,N_17501);
nor U19314 (N_19314,N_12136,N_13011);
nor U19315 (N_19315,N_14009,N_13004);
or U19316 (N_19316,N_12589,N_15086);
xor U19317 (N_19317,N_14644,N_15800);
or U19318 (N_19318,N_13903,N_15179);
nor U19319 (N_19319,N_12542,N_12313);
or U19320 (N_19320,N_13807,N_13197);
nand U19321 (N_19321,N_16499,N_17870);
and U19322 (N_19322,N_17699,N_13597);
nand U19323 (N_19323,N_16665,N_14802);
and U19324 (N_19324,N_14531,N_12992);
or U19325 (N_19325,N_16253,N_17744);
xnor U19326 (N_19326,N_12625,N_12191);
or U19327 (N_19327,N_12359,N_14479);
or U19328 (N_19328,N_12692,N_13910);
and U19329 (N_19329,N_15088,N_14111);
nor U19330 (N_19330,N_14210,N_14056);
nor U19331 (N_19331,N_13924,N_16228);
and U19332 (N_19332,N_13676,N_12439);
or U19333 (N_19333,N_17934,N_15348);
nor U19334 (N_19334,N_12438,N_16622);
or U19335 (N_19335,N_14826,N_17299);
nand U19336 (N_19336,N_15165,N_13311);
nand U19337 (N_19337,N_12062,N_17725);
nand U19338 (N_19338,N_13578,N_15005);
nand U19339 (N_19339,N_12539,N_16040);
or U19340 (N_19340,N_17236,N_15992);
or U19341 (N_19341,N_14545,N_14638);
nor U19342 (N_19342,N_15258,N_13084);
or U19343 (N_19343,N_12890,N_13307);
or U19344 (N_19344,N_12596,N_15560);
nor U19345 (N_19345,N_13907,N_16777);
or U19346 (N_19346,N_13729,N_15948);
xor U19347 (N_19347,N_17384,N_14268);
or U19348 (N_19348,N_14809,N_13098);
nand U19349 (N_19349,N_17452,N_12525);
xor U19350 (N_19350,N_17192,N_14188);
or U19351 (N_19351,N_14963,N_15279);
or U19352 (N_19352,N_14843,N_16771);
or U19353 (N_19353,N_17114,N_14800);
xnor U19354 (N_19354,N_14299,N_12466);
nor U19355 (N_19355,N_15267,N_16538);
nor U19356 (N_19356,N_12333,N_17793);
and U19357 (N_19357,N_15305,N_16750);
and U19358 (N_19358,N_15717,N_12427);
or U19359 (N_19359,N_15604,N_17065);
or U19360 (N_19360,N_14246,N_15342);
nand U19361 (N_19361,N_13889,N_15630);
and U19362 (N_19362,N_17844,N_13181);
or U19363 (N_19363,N_16816,N_17945);
and U19364 (N_19364,N_12488,N_17720);
or U19365 (N_19365,N_17558,N_16923);
nor U19366 (N_19366,N_16430,N_15079);
or U19367 (N_19367,N_14165,N_14149);
xor U19368 (N_19368,N_14717,N_15834);
and U19369 (N_19369,N_14463,N_12225);
nand U19370 (N_19370,N_15997,N_12858);
and U19371 (N_19371,N_17199,N_16894);
nor U19372 (N_19372,N_17313,N_13673);
nor U19373 (N_19373,N_12983,N_16745);
and U19374 (N_19374,N_12069,N_17290);
and U19375 (N_19375,N_13584,N_12391);
xor U19376 (N_19376,N_13083,N_12577);
nor U19377 (N_19377,N_17745,N_14136);
or U19378 (N_19378,N_16514,N_17760);
nor U19379 (N_19379,N_13057,N_14382);
nor U19380 (N_19380,N_17942,N_12635);
and U19381 (N_19381,N_12845,N_16536);
and U19382 (N_19382,N_17104,N_16437);
nand U19383 (N_19383,N_15925,N_13080);
nor U19384 (N_19384,N_16173,N_14738);
nor U19385 (N_19385,N_17634,N_15162);
or U19386 (N_19386,N_16973,N_15205);
xor U19387 (N_19387,N_17266,N_14639);
nand U19388 (N_19388,N_13984,N_15269);
or U19389 (N_19389,N_14624,N_15392);
and U19390 (N_19390,N_14110,N_15782);
or U19391 (N_19391,N_16393,N_16668);
xnor U19392 (N_19392,N_16694,N_16315);
nor U19393 (N_19393,N_15429,N_15960);
and U19394 (N_19394,N_14789,N_17016);
xnor U19395 (N_19395,N_12379,N_16577);
nor U19396 (N_19396,N_12694,N_15297);
and U19397 (N_19397,N_12132,N_14708);
and U19398 (N_19398,N_15216,N_16132);
nor U19399 (N_19399,N_15334,N_14735);
nand U19400 (N_19400,N_13509,N_17615);
nor U19401 (N_19401,N_12619,N_14310);
nor U19402 (N_19402,N_13105,N_15463);
nor U19403 (N_19403,N_14400,N_16688);
or U19404 (N_19404,N_17819,N_14662);
and U19405 (N_19405,N_14436,N_17368);
and U19406 (N_19406,N_14381,N_17840);
or U19407 (N_19407,N_17197,N_16762);
and U19408 (N_19408,N_14645,N_17129);
nor U19409 (N_19409,N_14439,N_16510);
or U19410 (N_19410,N_13030,N_16379);
or U19411 (N_19411,N_13844,N_15381);
or U19412 (N_19412,N_15134,N_15495);
xor U19413 (N_19413,N_15707,N_16158);
nor U19414 (N_19414,N_13400,N_14360);
xnor U19415 (N_19415,N_12739,N_12792);
or U19416 (N_19416,N_12458,N_16835);
or U19417 (N_19417,N_16749,N_17398);
nor U19418 (N_19418,N_12269,N_17809);
and U19419 (N_19419,N_16994,N_16720);
nor U19420 (N_19420,N_17030,N_13440);
and U19421 (N_19421,N_13235,N_17904);
nand U19422 (N_19422,N_13071,N_14191);
nor U19423 (N_19423,N_12918,N_13318);
and U19424 (N_19424,N_14669,N_12016);
and U19425 (N_19425,N_14727,N_15215);
and U19426 (N_19426,N_13639,N_17603);
and U19427 (N_19427,N_13620,N_13759);
and U19428 (N_19428,N_17812,N_14235);
nor U19429 (N_19429,N_14243,N_14603);
and U19430 (N_19430,N_17920,N_14696);
nor U19431 (N_19431,N_12377,N_12585);
xnor U19432 (N_19432,N_15894,N_12412);
nor U19433 (N_19433,N_12817,N_12108);
nand U19434 (N_19434,N_17138,N_16180);
nor U19435 (N_19435,N_16549,N_17574);
nand U19436 (N_19436,N_14661,N_17562);
or U19437 (N_19437,N_12338,N_17389);
and U19438 (N_19438,N_15242,N_12974);
nor U19439 (N_19439,N_16502,N_14472);
and U19440 (N_19440,N_16579,N_14087);
and U19441 (N_19441,N_12567,N_13763);
and U19442 (N_19442,N_13139,N_12460);
or U19443 (N_19443,N_15651,N_15702);
nand U19444 (N_19444,N_14337,N_12173);
nor U19445 (N_19445,N_17590,N_16653);
and U19446 (N_19446,N_13468,N_16239);
or U19447 (N_19447,N_12856,N_16748);
nor U19448 (N_19448,N_14462,N_16321);
nand U19449 (N_19449,N_15957,N_13213);
nor U19450 (N_19450,N_17040,N_12886);
and U19451 (N_19451,N_17738,N_12201);
and U19452 (N_19452,N_12650,N_15796);
and U19453 (N_19453,N_17006,N_17091);
or U19454 (N_19454,N_15766,N_15553);
nor U19455 (N_19455,N_14814,N_16542);
nor U19456 (N_19456,N_17659,N_15471);
nand U19457 (N_19457,N_16703,N_17485);
nand U19458 (N_19458,N_17677,N_15001);
nor U19459 (N_19459,N_14107,N_13170);
or U19460 (N_19460,N_14192,N_15728);
nor U19461 (N_19461,N_17202,N_17474);
nor U19462 (N_19462,N_12540,N_12426);
xnor U19463 (N_19463,N_14094,N_12337);
nor U19464 (N_19464,N_16400,N_13582);
nand U19465 (N_19465,N_12820,N_16805);
nor U19466 (N_19466,N_13641,N_14128);
and U19467 (N_19467,N_17324,N_13026);
nand U19468 (N_19468,N_17168,N_13161);
and U19469 (N_19469,N_14511,N_15090);
nand U19470 (N_19470,N_15436,N_17009);
nand U19471 (N_19471,N_12594,N_14759);
nor U19472 (N_19472,N_13852,N_16878);
nand U19473 (N_19473,N_17514,N_17827);
nor U19474 (N_19474,N_12129,N_12101);
nor U19475 (N_19475,N_14326,N_17383);
and U19476 (N_19476,N_17177,N_13445);
or U19477 (N_19477,N_14836,N_17471);
nand U19478 (N_19478,N_16032,N_15922);
xor U19479 (N_19479,N_17056,N_17626);
or U19480 (N_19480,N_12448,N_17774);
nor U19481 (N_19481,N_15235,N_15126);
nand U19482 (N_19482,N_14700,N_16076);
nor U19483 (N_19483,N_17435,N_12671);
nand U19484 (N_19484,N_13603,N_15454);
or U19485 (N_19485,N_17238,N_15375);
or U19486 (N_19486,N_14525,N_12957);
and U19487 (N_19487,N_15372,N_16772);
or U19488 (N_19488,N_13954,N_17899);
and U19489 (N_19489,N_13712,N_15365);
nor U19490 (N_19490,N_17866,N_15158);
or U19491 (N_19491,N_12184,N_13194);
and U19492 (N_19492,N_13239,N_15601);
nor U19493 (N_19493,N_13090,N_15420);
nand U19494 (N_19494,N_15704,N_13287);
nand U19495 (N_19495,N_15672,N_12913);
or U19496 (N_19496,N_12621,N_15273);
or U19497 (N_19497,N_14295,N_14607);
or U19498 (N_19498,N_14636,N_17225);
and U19499 (N_19499,N_16883,N_13573);
nand U19500 (N_19500,N_13441,N_15712);
or U19501 (N_19501,N_17088,N_16374);
xnor U19502 (N_19502,N_16809,N_15762);
or U19503 (N_19503,N_15455,N_17608);
or U19504 (N_19504,N_16107,N_13731);
nor U19505 (N_19505,N_15280,N_17393);
nor U19506 (N_19506,N_16083,N_14340);
xor U19507 (N_19507,N_15336,N_17892);
or U19508 (N_19508,N_14248,N_12636);
nor U19509 (N_19509,N_13787,N_17800);
or U19510 (N_19510,N_15748,N_15338);
nor U19511 (N_19511,N_13533,N_16218);
and U19512 (N_19512,N_14510,N_16873);
nand U19513 (N_19513,N_17638,N_16432);
and U19514 (N_19514,N_13606,N_14331);
and U19515 (N_19515,N_12898,N_14275);
nand U19516 (N_19516,N_13771,N_16635);
nand U19517 (N_19517,N_17004,N_12615);
nand U19518 (N_19518,N_14427,N_16232);
and U19519 (N_19519,N_14888,N_14719);
nand U19520 (N_19520,N_15873,N_12691);
or U19521 (N_19521,N_14175,N_14431);
nand U19522 (N_19522,N_13319,N_14077);
nor U19523 (N_19523,N_17439,N_16675);
nand U19524 (N_19524,N_12288,N_14019);
nand U19525 (N_19525,N_13289,N_16803);
xor U19526 (N_19526,N_13637,N_15380);
nor U19527 (N_19527,N_16219,N_16602);
nand U19528 (N_19528,N_14131,N_13691);
and U19529 (N_19529,N_13644,N_17031);
or U19530 (N_19530,N_12981,N_15791);
or U19531 (N_19531,N_16189,N_17882);
nand U19532 (N_19532,N_13136,N_17703);
or U19533 (N_19533,N_15675,N_14557);
or U19534 (N_19534,N_13694,N_16282);
or U19535 (N_19535,N_12750,N_17101);
nor U19536 (N_19536,N_15416,N_16195);
xor U19537 (N_19537,N_14705,N_14401);
nand U19538 (N_19538,N_13940,N_16023);
nand U19539 (N_19539,N_16324,N_15345);
nor U19540 (N_19540,N_15243,N_12425);
nand U19541 (N_19541,N_12501,N_17935);
nor U19542 (N_19542,N_14251,N_13063);
xor U19543 (N_19543,N_16667,N_13719);
xnor U19544 (N_19544,N_15354,N_17427);
nor U19545 (N_19545,N_12598,N_14788);
nand U19546 (N_19546,N_15231,N_15037);
and U19547 (N_19547,N_17412,N_17550);
or U19548 (N_19548,N_17150,N_17336);
nand U19549 (N_19549,N_15893,N_13312);
nor U19550 (N_19550,N_17352,N_12205);
or U19551 (N_19551,N_15473,N_17025);
or U19552 (N_19552,N_15132,N_12204);
xor U19553 (N_19553,N_12628,N_17118);
xor U19554 (N_19554,N_15956,N_14234);
nand U19555 (N_19555,N_16575,N_14718);
nand U19556 (N_19556,N_17843,N_15936);
nand U19557 (N_19557,N_12713,N_15283);
or U19558 (N_19558,N_17144,N_13813);
or U19559 (N_19559,N_14143,N_13271);
nand U19560 (N_19560,N_13443,N_13066);
xor U19561 (N_19561,N_17206,N_12351);
xnor U19562 (N_19562,N_15924,N_15665);
and U19563 (N_19563,N_16825,N_15472);
nand U19564 (N_19564,N_17718,N_15003);
nand U19565 (N_19565,N_12518,N_16681);
nand U19566 (N_19566,N_12736,N_17440);
or U19567 (N_19567,N_14722,N_15973);
and U19568 (N_19568,N_13454,N_15219);
nor U19569 (N_19569,N_14614,N_16966);
or U19570 (N_19570,N_17077,N_15775);
nand U19571 (N_19571,N_17816,N_12578);
and U19572 (N_19572,N_15938,N_17893);
or U19573 (N_19573,N_13775,N_13733);
nor U19574 (N_19574,N_12219,N_12904);
nand U19575 (N_19575,N_17157,N_14154);
and U19576 (N_19576,N_13749,N_15784);
nor U19577 (N_19577,N_16301,N_15774);
and U19578 (N_19578,N_17759,N_17426);
nand U19579 (N_19579,N_13413,N_17572);
or U19580 (N_19580,N_15191,N_16350);
and U19581 (N_19581,N_13360,N_15195);
xnor U19582 (N_19582,N_15208,N_13568);
nand U19583 (N_19583,N_13382,N_12954);
nor U19584 (N_19584,N_12862,N_14378);
nand U19585 (N_19585,N_13174,N_16888);
nor U19586 (N_19586,N_12317,N_13640);
nand U19587 (N_19587,N_12588,N_15978);
xnor U19588 (N_19588,N_12088,N_12372);
nand U19589 (N_19589,N_15008,N_16641);
xor U19590 (N_19590,N_17139,N_14723);
xnor U19591 (N_19591,N_12763,N_12125);
xnor U19592 (N_19592,N_12948,N_16958);
or U19593 (N_19593,N_12254,N_13065);
nor U19594 (N_19594,N_17903,N_15374);
nand U19595 (N_19595,N_16798,N_17267);
nand U19596 (N_19596,N_17855,N_13730);
nand U19597 (N_19597,N_17497,N_14737);
xnor U19598 (N_19598,N_16095,N_14567);
nor U19599 (N_19599,N_14542,N_12522);
nor U19600 (N_19600,N_14628,N_13961);
or U19601 (N_19601,N_12255,N_13726);
and U19602 (N_19602,N_12513,N_15715);
nor U19603 (N_19603,N_16636,N_15877);
and U19604 (N_19604,N_15812,N_16336);
xnor U19605 (N_19605,N_12562,N_17790);
or U19606 (N_19606,N_14212,N_15172);
nand U19607 (N_19607,N_15879,N_12342);
nand U19608 (N_19608,N_13893,N_13613);
nand U19609 (N_19609,N_17570,N_13508);
nor U19610 (N_19610,N_14066,N_15415);
and U19611 (N_19611,N_12194,N_15645);
or U19612 (N_19612,N_13522,N_17817);
and U19613 (N_19613,N_12383,N_13664);
nor U19614 (N_19614,N_16179,N_16677);
nor U19615 (N_19615,N_13696,N_16960);
nand U19616 (N_19616,N_13388,N_13982);
nor U19617 (N_19617,N_13693,N_13292);
or U19618 (N_19618,N_12025,N_13273);
or U19619 (N_19619,N_13452,N_12046);
nor U19620 (N_19620,N_15699,N_12756);
or U19621 (N_19621,N_13242,N_15130);
nand U19622 (N_19622,N_17280,N_15032);
nor U19623 (N_19623,N_15625,N_14214);
xor U19624 (N_19624,N_12073,N_14417);
and U19625 (N_19625,N_16044,N_17532);
nand U19626 (N_19626,N_16298,N_16812);
nor U19627 (N_19627,N_13117,N_16503);
nand U19628 (N_19628,N_15524,N_14114);
nand U19629 (N_19629,N_15676,N_17999);
and U19630 (N_19630,N_12486,N_17936);
nand U19631 (N_19631,N_12537,N_16868);
nand U19632 (N_19632,N_12605,N_14177);
and U19633 (N_19633,N_13574,N_17275);
nor U19634 (N_19634,N_17469,N_15663);
xor U19635 (N_19635,N_13298,N_17018);
and U19636 (N_19636,N_12932,N_17099);
nand U19637 (N_19637,N_12332,N_15167);
nor U19638 (N_19638,N_14995,N_17162);
nand U19639 (N_19639,N_16273,N_15052);
or U19640 (N_19640,N_15033,N_13801);
or U19641 (N_19641,N_17820,N_12040);
or U19642 (N_19642,N_16818,N_15909);
nand U19643 (N_19643,N_12017,N_14051);
nor U19644 (N_19644,N_15256,N_17906);
nor U19645 (N_19645,N_15598,N_12217);
xnor U19646 (N_19646,N_14370,N_12165);
xnor U19647 (N_19647,N_14615,N_15332);
nand U19648 (N_19648,N_12107,N_17897);
and U19649 (N_19649,N_15498,N_13943);
nand U19650 (N_19650,N_14195,N_13339);
or U19651 (N_19651,N_15341,N_14702);
or U19652 (N_19652,N_15659,N_13442);
nor U19653 (N_19653,N_12720,N_15751);
nor U19654 (N_19654,N_15857,N_14884);
nand U19655 (N_19655,N_16423,N_16633);
and U19656 (N_19656,N_17174,N_14366);
nor U19657 (N_19657,N_16085,N_17200);
or U19658 (N_19658,N_12703,N_17462);
nand U19659 (N_19659,N_17958,N_12457);
or U19660 (N_19660,N_16025,N_12545);
nand U19661 (N_19661,N_13646,N_13669);
and U19662 (N_19662,N_16022,N_13232);
nand U19663 (N_19663,N_13478,N_14592);
nor U19664 (N_19664,N_15014,N_17340);
nand U19665 (N_19665,N_15603,N_13050);
nand U19666 (N_19666,N_15111,N_12481);
nor U19667 (N_19667,N_16395,N_15044);
xnor U19668 (N_19668,N_12745,N_17779);
nand U19669 (N_19669,N_17080,N_14745);
and U19670 (N_19670,N_12955,N_13229);
nor U19671 (N_19671,N_13120,N_14794);
or U19672 (N_19672,N_14452,N_12133);
and U19673 (N_19673,N_12808,N_13560);
nand U19674 (N_19674,N_14469,N_16508);
nand U19675 (N_19675,N_16217,N_17103);
nor U19676 (N_19676,N_15870,N_16367);
nor U19677 (N_19677,N_16589,N_16316);
nor U19678 (N_19678,N_17217,N_14343);
xor U19679 (N_19679,N_14475,N_12962);
xor U19680 (N_19680,N_13216,N_12344);
and U19681 (N_19681,N_17701,N_16498);
or U19682 (N_19682,N_17037,N_17251);
or U19683 (N_19683,N_12910,N_17839);
nand U19684 (N_19684,N_13209,N_17977);
and U19685 (N_19685,N_15074,N_17317);
nor U19686 (N_19686,N_16020,N_14359);
and U19687 (N_19687,N_12721,N_15029);
nor U19688 (N_19688,N_13751,N_17377);
and U19689 (N_19689,N_13448,N_17152);
and U19690 (N_19690,N_13612,N_12965);
or U19691 (N_19691,N_17092,N_16922);
nand U19692 (N_19692,N_16855,N_17396);
xor U19693 (N_19693,N_16317,N_15299);
or U19694 (N_19694,N_13663,N_17652);
nor U19695 (N_19695,N_12760,N_14571);
and U19696 (N_19696,N_17757,N_15327);
or U19697 (N_19697,N_12521,N_17509);
or U19698 (N_19698,N_13376,N_14940);
nand U19699 (N_19699,N_17931,N_14219);
nor U19700 (N_19700,N_12410,N_13648);
nor U19701 (N_19701,N_13481,N_17107);
nor U19702 (N_19702,N_13878,N_17538);
and U19703 (N_19703,N_16505,N_15403);
and U19704 (N_19704,N_14600,N_17149);
nand U19705 (N_19705,N_12727,N_17890);
nor U19706 (N_19706,N_16936,N_17311);
or U19707 (N_19707,N_17175,N_17773);
or U19708 (N_19708,N_16047,N_14688);
or U19709 (N_19709,N_13412,N_14632);
nor U19710 (N_19710,N_16024,N_14334);
nor U19711 (N_19711,N_13750,N_15330);
nand U19712 (N_19712,N_17493,N_17066);
nor U19713 (N_19713,N_16261,N_15621);
or U19714 (N_19714,N_15229,N_13493);
or U19715 (N_19715,N_13190,N_12863);
nor U19716 (N_19716,N_15373,N_16556);
nor U19717 (N_19717,N_15296,N_14811);
xor U19718 (N_19718,N_14083,N_15579);
nand U19719 (N_19719,N_13329,N_13946);
or U19720 (N_19720,N_12568,N_12034);
and U19721 (N_19721,N_16258,N_14322);
nor U19722 (N_19722,N_12841,N_13668);
and U19723 (N_19723,N_17035,N_14481);
and U19724 (N_19724,N_15964,N_15670);
xor U19725 (N_19725,N_15309,N_16329);
nand U19726 (N_19726,N_14256,N_15410);
nand U19727 (N_19727,N_13126,N_14520);
and U19728 (N_19728,N_16410,N_13148);
and U19729 (N_19729,N_13262,N_12505);
nor U19730 (N_19730,N_17601,N_13530);
nor U19731 (N_19731,N_13515,N_12556);
nor U19732 (N_19732,N_16884,N_14281);
and U19733 (N_19733,N_16898,N_16628);
and U19734 (N_19734,N_13716,N_14227);
or U19735 (N_19735,N_17213,N_14164);
and U19736 (N_19736,N_15198,N_17055);
and U19737 (N_19737,N_16902,N_14033);
and U19738 (N_19738,N_14168,N_17526);
and U19739 (N_19739,N_13281,N_13333);
nand U19740 (N_19740,N_13276,N_13674);
or U19741 (N_19741,N_16870,N_14007);
nor U19742 (N_19742,N_13260,N_12606);
or U19743 (N_19743,N_16288,N_16904);
and U19744 (N_19744,N_13882,N_13516);
and U19745 (N_19745,N_16250,N_14426);
nor U19746 (N_19746,N_17587,N_13886);
and U19747 (N_19747,N_12248,N_13710);
or U19748 (N_19748,N_15776,N_13270);
nor U19749 (N_19749,N_15818,N_15914);
and U19750 (N_19750,N_13942,N_17181);
nand U19751 (N_19751,N_17333,N_17335);
nand U19752 (N_19752,N_16240,N_14139);
and U19753 (N_19753,N_17212,N_16569);
or U19754 (N_19754,N_15394,N_12930);
or U19755 (N_19755,N_15045,N_16543);
or U19756 (N_19756,N_15012,N_13610);
and U19757 (N_19757,N_15261,N_12112);
or U19758 (N_19758,N_14691,N_17264);
or U19759 (N_19759,N_14072,N_12507);
nor U19760 (N_19760,N_13254,N_14983);
nand U19761 (N_19761,N_15100,N_12555);
or U19762 (N_19762,N_12354,N_15390);
nor U19763 (N_19763,N_13407,N_16465);
or U19764 (N_19764,N_17354,N_14850);
and U19765 (N_19765,N_12081,N_14955);
xor U19766 (N_19766,N_14928,N_16348);
or U19767 (N_19767,N_17124,N_14606);
and U19768 (N_19768,N_14988,N_16931);
nand U19769 (N_19769,N_14774,N_14769);
and U19770 (N_19770,N_13908,N_12265);
nor U19771 (N_19771,N_14434,N_17506);
nand U19772 (N_19772,N_12775,N_17772);
xor U19773 (N_19773,N_14494,N_13097);
nand U19774 (N_19774,N_13904,N_13686);
or U19775 (N_19775,N_12679,N_12702);
or U19776 (N_19776,N_16208,N_14155);
or U19777 (N_19777,N_15627,N_13826);
nor U19778 (N_19778,N_16660,N_14419);
and U19779 (N_19779,N_12601,N_13185);
and U19780 (N_19780,N_14699,N_16649);
nor U19781 (N_19781,N_15622,N_17932);
nor U19782 (N_19782,N_13207,N_12207);
nand U19783 (N_19783,N_15996,N_14972);
nor U19784 (N_19784,N_16962,N_16046);
nand U19785 (N_19785,N_15187,N_14187);
and U19786 (N_19786,N_14874,N_17425);
nor U19787 (N_19787,N_17387,N_15085);
or U19788 (N_19788,N_12432,N_15657);
and U19789 (N_19789,N_14863,N_15856);
nand U19790 (N_19790,N_15722,N_14773);
nor U19791 (N_19791,N_14363,N_15993);
or U19792 (N_19792,N_15723,N_13146);
or U19793 (N_19793,N_17997,N_14515);
or U19794 (N_19794,N_12056,N_15742);
or U19795 (N_19795,N_12041,N_17222);
nor U19796 (N_19796,N_14412,N_13330);
and U19797 (N_19797,N_12909,N_14547);
xnor U19798 (N_19798,N_15683,N_14206);
and U19799 (N_19799,N_13653,N_13781);
nand U19800 (N_19800,N_16548,N_17804);
nor U19801 (N_19801,N_17607,N_12279);
and U19802 (N_19802,N_15525,N_14992);
xor U19803 (N_19803,N_13234,N_13938);
or U19804 (N_19804,N_12939,N_15543);
and U19805 (N_19805,N_13626,N_12364);
and U19806 (N_19806,N_16659,N_13743);
or U19807 (N_19807,N_16156,N_14229);
or U19808 (N_19808,N_17561,N_12227);
nor U19809 (N_19809,N_17402,N_16029);
nand U19810 (N_19810,N_17627,N_14934);
nor U19811 (N_19811,N_16072,N_17847);
and U19812 (N_19812,N_12549,N_17327);
nand U19813 (N_19813,N_12892,N_14941);
nor U19814 (N_19814,N_16037,N_17667);
or U19815 (N_19815,N_13621,N_16647);
nand U19816 (N_19816,N_13266,N_13929);
or U19817 (N_19817,N_13435,N_14570);
nand U19818 (N_19818,N_14772,N_16278);
nor U19819 (N_19819,N_17484,N_16198);
or U19820 (N_19820,N_13649,N_12582);
nor U19821 (N_19821,N_13627,N_17404);
nor U19822 (N_19822,N_16344,N_13058);
nand U19823 (N_19823,N_15054,N_16504);
nor U19824 (N_19824,N_16114,N_14020);
nand U19825 (N_19825,N_15135,N_16372);
or U19826 (N_19826,N_12560,N_16617);
xnor U19827 (N_19827,N_12203,N_13426);
nor U19828 (N_19828,N_14682,N_16972);
nand U19829 (N_19829,N_14517,N_13089);
nor U19830 (N_19830,N_17134,N_15460);
and U19831 (N_19831,N_15271,N_13825);
or U19832 (N_19832,N_14358,N_12109);
nor U19833 (N_19833,N_13401,N_12235);
nand U19834 (N_19834,N_16310,N_16991);
nor U19835 (N_19835,N_13519,N_16460);
nor U19836 (N_19836,N_17546,N_16224);
and U19837 (N_19837,N_16194,N_12561);
or U19838 (N_19838,N_15705,N_14055);
nor U19839 (N_19839,N_15755,N_13792);
or U19840 (N_19840,N_12127,N_13796);
nand U19841 (N_19841,N_13029,N_13985);
and U19842 (N_19842,N_15836,N_13200);
nor U19843 (N_19843,N_16558,N_16246);
or U19844 (N_19844,N_17374,N_16981);
and U19845 (N_19845,N_12172,N_14841);
and U19846 (N_19846,N_14313,N_14831);
or U19847 (N_19847,N_13853,N_17039);
nor U19848 (N_19848,N_17073,N_17378);
nor U19849 (N_19849,N_13798,N_17872);
nor U19850 (N_19850,N_16885,N_14783);
nand U19851 (N_19851,N_15441,N_14085);
nand U19852 (N_19852,N_16997,N_14906);
nand U19853 (N_19853,N_15110,N_14853);
nor U19854 (N_19854,N_16257,N_16593);
nor U19855 (N_19855,N_16365,N_14523);
and U19856 (N_19856,N_15321,N_15532);
nor U19857 (N_19857,N_12666,N_15554);
or U19858 (N_19858,N_13464,N_12349);
or U19859 (N_19859,N_15907,N_17022);
nand U19860 (N_19860,N_16359,N_12777);
and U19861 (N_19861,N_15181,N_17044);
nand U19862 (N_19862,N_16786,N_17537);
and U19863 (N_19863,N_15654,N_12670);
or U19864 (N_19864,N_16294,N_14596);
nor U19865 (N_19865,N_14048,N_17341);
or U19866 (N_19866,N_13315,N_14410);
and U19867 (N_19867,N_17309,N_12822);
xor U19868 (N_19868,N_13752,N_14008);
and U19869 (N_19869,N_15700,N_14484);
nor U19870 (N_19870,N_13705,N_17623);
or U19871 (N_19871,N_17648,N_16639);
and U19872 (N_19872,N_16706,N_15637);
and U19873 (N_19873,N_13253,N_14681);
nor U19874 (N_19874,N_14361,N_16405);
or U19875 (N_19875,N_13877,N_12813);
and U19876 (N_19876,N_12592,N_16266);
nor U19877 (N_19877,N_13015,N_17366);
and U19878 (N_19878,N_12523,N_17399);
and U19879 (N_19879,N_14302,N_14467);
nor U19880 (N_19880,N_17108,N_13511);
nor U19881 (N_19881,N_12731,N_16358);
and U19882 (N_19882,N_12015,N_14630);
or U19883 (N_19883,N_14356,N_17214);
and U19884 (N_19884,N_14828,N_15148);
or U19885 (N_19885,N_12982,N_16215);
nor U19886 (N_19886,N_15545,N_14311);
nor U19887 (N_19887,N_17869,N_15727);
or U19888 (N_19888,N_15991,N_13323);
and U19889 (N_19889,N_14277,N_13524);
nor U19890 (N_19890,N_15095,N_13720);
or U19891 (N_19891,N_17221,N_17005);
and U19892 (N_19892,N_14782,N_16404);
nand U19893 (N_19893,N_12373,N_13037);
nand U19894 (N_19894,N_12617,N_15743);
nor U19895 (N_19895,N_16134,N_13951);
and U19896 (N_19896,N_16676,N_13736);
nor U19897 (N_19897,N_17293,N_15470);
or U19898 (N_19898,N_17207,N_15462);
nor U19899 (N_19899,N_12570,N_17943);
and U19900 (N_19900,N_14233,N_12835);
nand U19901 (N_19901,N_17674,N_16901);
xor U19902 (N_19902,N_16867,N_13116);
or U19903 (N_19903,N_16384,N_13803);
or U19904 (N_19904,N_17651,N_14024);
xor U19905 (N_19905,N_15370,N_14287);
nor U19906 (N_19906,N_12270,N_16286);
nand U19907 (N_19907,N_14416,N_12781);
xnor U19908 (N_19908,N_15351,N_15710);
nand U19909 (N_19909,N_17848,N_15263);
xnor U19910 (N_19910,N_14215,N_13794);
nor U19911 (N_19911,N_14156,N_14046);
or U19912 (N_19912,N_17447,N_17961);
nand U19913 (N_19913,N_13735,N_15411);
and U19914 (N_19914,N_13804,N_17173);
and U19915 (N_19915,N_12471,N_14842);
nor U19916 (N_19916,N_15359,N_17914);
and U19917 (N_19917,N_12318,N_14820);
xnor U19918 (N_19918,N_14514,N_17555);
nor U19919 (N_19919,N_12492,N_15278);
or U19920 (N_19920,N_16522,N_17227);
nor U19921 (N_19921,N_17171,N_14932);
or U19922 (N_19922,N_12779,N_13518);
xor U19923 (N_19923,N_14787,N_16533);
nor U19924 (N_19924,N_12951,N_12614);
and U19925 (N_19925,N_15852,N_12687);
nand U19926 (N_19926,N_13737,N_15512);
or U19927 (N_19927,N_12280,N_14425);
nand U19928 (N_19928,N_14045,N_15217);
nor U19929 (N_19929,N_15325,N_16463);
nand U19930 (N_19930,N_13868,N_12535);
nor U19931 (N_19931,N_14765,N_16303);
or U19932 (N_19932,N_13531,N_12664);
or U19933 (N_19933,N_15193,N_15120);
nand U19934 (N_19934,N_16121,N_16042);
or U19935 (N_19935,N_13123,N_13258);
and U19936 (N_19936,N_13495,N_17972);
or U19937 (N_19937,N_12719,N_17320);
nand U19938 (N_19938,N_14598,N_16601);
or U19939 (N_19939,N_12838,N_12865);
or U19940 (N_19940,N_15939,N_15154);
nand U19941 (N_19941,N_17824,N_17457);
nor U19942 (N_19942,N_17416,N_17786);
or U19943 (N_19943,N_16832,N_13167);
and U19944 (N_19944,N_13419,N_13975);
nor U19945 (N_19945,N_17211,N_12795);
and U19946 (N_19946,N_14591,N_13986);
or U19947 (N_19947,N_15631,N_17062);
or U19948 (N_19948,N_12767,N_12045);
nand U19949 (N_19949,N_15091,N_15983);
nor U19950 (N_19950,N_13130,N_16428);
nand U19951 (N_19951,N_12007,N_12551);
nand U19952 (N_19952,N_13974,N_16197);
or U19953 (N_19953,N_12836,N_12415);
or U19954 (N_19954,N_14130,N_16780);
nand U19955 (N_19955,N_12848,N_13418);
nor U19956 (N_19956,N_14411,N_14010);
nand U19957 (N_19957,N_15513,N_15587);
nand U19958 (N_19958,N_12859,N_14823);
nor U19959 (N_19959,N_13937,N_16045);
nor U19960 (N_19960,N_16468,N_15690);
nor U19961 (N_19961,N_14451,N_15608);
and U19962 (N_19962,N_16640,N_14657);
nor U19963 (N_19963,N_12771,N_16148);
and U19964 (N_19964,N_13504,N_14027);
and U19965 (N_19965,N_17728,N_17752);
nor U19966 (N_19966,N_13154,N_13949);
xor U19967 (N_19967,N_14549,N_17194);
nand U19968 (N_19968,N_16111,N_17215);
nor U19969 (N_19969,N_12935,N_17544);
and U19970 (N_19970,N_14283,N_12911);
or U19971 (N_19971,N_15357,N_15821);
nand U19972 (N_19972,N_14650,N_16131);
and U19973 (N_19973,N_15578,N_13378);
nor U19974 (N_19974,N_17535,N_14936);
nand U19975 (N_19975,N_12198,N_17966);
nor U19976 (N_19976,N_15509,N_12640);
nor U19977 (N_19977,N_13132,N_12312);
nand U19978 (N_19978,N_13310,N_12504);
or U19979 (N_19979,N_13399,N_15988);
or U19980 (N_19980,N_17256,N_14030);
nor U19981 (N_19981,N_16765,N_17516);
nand U19982 (N_19982,N_17765,N_13655);
or U19983 (N_19983,N_14881,N_15547);
and U19984 (N_19984,N_13182,N_15926);
or U19985 (N_19985,N_16568,N_15307);
nand U19986 (N_19986,N_12124,N_14379);
nand U19987 (N_19987,N_12978,N_17633);
and U19988 (N_19988,N_13151,N_15530);
or U19989 (N_19989,N_17507,N_13483);
and U19990 (N_19990,N_13556,N_15947);
nand U19991 (N_19991,N_16513,N_15662);
nor U19992 (N_19992,N_17319,N_16495);
or U19993 (N_19993,N_16976,N_17741);
nor U19994 (N_19994,N_15318,N_15199);
nand U19995 (N_19995,N_12325,N_17270);
nand U19996 (N_19996,N_13760,N_17121);
nor U19997 (N_19997,N_13848,N_13944);
or U19998 (N_19998,N_14887,N_12973);
and U19999 (N_19999,N_13917,N_15293);
nor U20000 (N_20000,N_12226,N_17512);
nor U20001 (N_20001,N_12743,N_14704);
or U20002 (N_20002,N_16828,N_17717);
nand U20003 (N_20003,N_14276,N_13462);
nand U20004 (N_20004,N_16104,N_17155);
and U20005 (N_20005,N_13279,N_16094);
nand U20006 (N_20006,N_14006,N_17551);
nor U20007 (N_20007,N_14292,N_15124);
or U20008 (N_20008,N_14126,N_15889);
and U20009 (N_20009,N_13862,N_14617);
and U20010 (N_20010,N_12128,N_14222);
nand U20011 (N_20011,N_12498,N_17367);
nor U20012 (N_20012,N_15157,N_17709);
or U20013 (N_20013,N_12240,N_16708);
and U20014 (N_20014,N_14273,N_16839);
nor U20015 (N_20015,N_15650,N_16587);
nand U20016 (N_20016,N_16529,N_17344);
and U20017 (N_20017,N_17415,N_17504);
or U20018 (N_20018,N_12524,N_16007);
nand U20019 (N_20019,N_16269,N_14729);
nand U20020 (N_20020,N_12798,N_15638);
nor U20021 (N_20021,N_14478,N_13680);
nor U20022 (N_20022,N_17362,N_15361);
nor U20023 (N_20023,N_12487,N_12114);
nand U20024 (N_20024,N_14652,N_17106);
nand U20025 (N_20025,N_15558,N_17407);
nor U20026 (N_20026,N_14097,N_16469);
xnor U20027 (N_20027,N_15266,N_17303);
or U20028 (N_20028,N_15887,N_16876);
or U20029 (N_20029,N_17371,N_14957);
and U20030 (N_20030,N_16054,N_13965);
nor U20031 (N_20031,N_15918,N_12849);
or U20032 (N_20032,N_13398,N_16332);
nor U20033 (N_20033,N_14506,N_17831);
or U20034 (N_20034,N_13034,N_14893);
nor U20035 (N_20035,N_16326,N_14760);
or U20036 (N_20036,N_13561,N_16010);
or U20037 (N_20037,N_14458,N_14825);
nor U20038 (N_20038,N_15285,N_16671);
nor U20039 (N_20039,N_16254,N_15788);
and U20040 (N_20040,N_13305,N_16283);
and U20041 (N_20041,N_15541,N_15294);
nand U20042 (N_20042,N_13513,N_12844);
nor U20043 (N_20043,N_13692,N_16039);
nor U20044 (N_20044,N_15038,N_12534);
nand U20045 (N_20045,N_17696,N_17867);
and U20046 (N_20046,N_15056,N_13231);
nor U20047 (N_20047,N_12346,N_13564);
nor U20048 (N_20048,N_12014,N_15276);
nor U20049 (N_20049,N_17878,N_13249);
nor U20050 (N_20050,N_14364,N_16963);
nor U20051 (N_20051,N_16846,N_13799);
and U20052 (N_20052,N_12675,N_16091);
nand U20053 (N_20053,N_12917,N_13996);
and U20054 (N_20054,N_16334,N_14946);
nand U20055 (N_20055,N_15414,N_13187);
or U20056 (N_20056,N_17905,N_16998);
and U20057 (N_20057,N_15437,N_15496);
nor U20058 (N_20058,N_13446,N_14947);
and U20059 (N_20059,N_13818,N_13918);
nand U20060 (N_20060,N_17370,N_13875);
nand U20061 (N_20061,N_13870,N_17580);
nor U20062 (N_20062,N_13808,N_17418);
nor U20063 (N_20063,N_12294,N_16381);
nand U20064 (N_20064,N_16746,N_14847);
or U20065 (N_20065,N_12387,N_14851);
nand U20066 (N_20066,N_16524,N_14690);
nor U20067 (N_20067,N_15260,N_16945);
and U20068 (N_20068,N_14707,N_16155);
nor U20069 (N_20069,N_15438,N_17926);
nor U20070 (N_20070,N_12048,N_15218);
nand U20071 (N_20071,N_16527,N_16341);
and U20072 (N_20072,N_13652,N_14288);
or U20073 (N_20073,N_17094,N_17090);
nand U20074 (N_20074,N_15377,N_16774);
and U20075 (N_20075,N_15951,N_14454);
nand U20076 (N_20076,N_17141,N_17490);
nor U20077 (N_20077,N_17226,N_12467);
or U20078 (N_20078,N_15364,N_12024);
nor U20079 (N_20079,N_14784,N_14608);
nor U20080 (N_20080,N_14626,N_14486);
or U20081 (N_20081,N_15681,N_14678);
or U20082 (N_20082,N_13867,N_13147);
and U20083 (N_20083,N_15975,N_12390);
nand U20084 (N_20084,N_15740,N_15814);
or U20085 (N_20085,N_16905,N_17136);
nand U20086 (N_20086,N_17625,N_14758);
and U20087 (N_20087,N_16814,N_15152);
or U20088 (N_20088,N_17502,N_16709);
or U20089 (N_20089,N_17814,N_15772);
nor U20090 (N_20090,N_13725,N_14344);
or U20091 (N_20091,N_17123,N_12150);
and U20092 (N_20092,N_17413,N_12446);
nor U20093 (N_20093,N_14325,N_12232);
and U20094 (N_20094,N_14060,N_13546);
nor U20095 (N_20095,N_14733,N_16318);
and U20096 (N_20096,N_13072,N_13128);
and U20097 (N_20097,N_17045,N_14685);
and U20098 (N_20098,N_14775,N_17505);
and U20099 (N_20099,N_13745,N_16256);
or U20100 (N_20100,N_15468,N_14664);
and U20101 (N_20101,N_16763,N_14035);
and U20102 (N_20102,N_15439,N_14157);
and U20103 (N_20103,N_17838,N_16420);
or U20104 (N_20104,N_17436,N_12461);
or U20105 (N_20105,N_14264,N_17596);
and U20106 (N_20106,N_13575,N_13821);
nand U20107 (N_20107,N_14730,N_15432);
xor U20108 (N_20108,N_16275,N_14000);
nor U20109 (N_20109,N_15042,N_15575);
or U20110 (N_20110,N_15469,N_13248);
and U20111 (N_20111,N_12090,N_14193);
or U20112 (N_20112,N_15761,N_16281);
nand U20113 (N_20113,N_17284,N_16019);
nand U20114 (N_20114,N_14901,N_13496);
nand U20115 (N_20115,N_15950,N_12994);
and U20116 (N_20116,N_16788,N_17466);
nor U20117 (N_20117,N_15049,N_13831);
xnor U20118 (N_20118,N_15446,N_14597);
or U20119 (N_20119,N_15451,N_15007);
nand U20120 (N_20120,N_14584,N_15458);
and U20121 (N_20121,N_17573,N_13471);
or U20122 (N_20122,N_13619,N_13544);
or U20123 (N_20123,N_14930,N_12479);
nor U20124 (N_20124,N_16163,N_17033);
nand U20125 (N_20125,N_12997,N_15839);
or U20126 (N_20126,N_15831,N_14117);
nand U20127 (N_20127,N_12840,N_15295);
nor U20128 (N_20128,N_14815,N_13355);
or U20129 (N_20129,N_15284,N_17650);
or U20130 (N_20130,N_12305,N_16098);
or U20131 (N_20131,N_12157,N_17161);
nor U20132 (N_20132,N_15489,N_12084);
xor U20133 (N_20133,N_12683,N_17456);
and U20134 (N_20134,N_16325,N_14099);
xnor U20135 (N_20135,N_15062,N_16937);
or U20136 (N_20136,N_12316,N_17565);
nand U20137 (N_20137,N_17000,N_14684);
and U20138 (N_20138,N_12417,N_17691);
xor U20139 (N_20139,N_12072,N_17536);
or U20140 (N_20140,N_13275,N_12746);
nand U20141 (N_20141,N_13915,N_13764);
nand U20142 (N_20142,N_15607,N_15510);
xor U20143 (N_20143,N_12512,N_16734);
or U20144 (N_20144,N_14261,N_17321);
and U20145 (N_20145,N_13609,N_14151);
nand U20146 (N_20146,N_17154,N_12118);
nor U20147 (N_20147,N_17359,N_13506);
or U20148 (N_20148,N_17012,N_15371);
nand U20149 (N_20149,N_13672,N_17376);
nor U20150 (N_20150,N_14890,N_16940);
nor U20151 (N_20151,N_13633,N_16252);
nand U20152 (N_20152,N_16342,N_13352);
or U20153 (N_20153,N_15583,N_16903);
nor U20154 (N_20154,N_15000,N_15594);
xor U20155 (N_20155,N_12038,N_14621);
or U20156 (N_20156,N_15146,N_17896);
and U20157 (N_20157,N_17250,N_12797);
and U20158 (N_20158,N_13490,N_16376);
nand U20159 (N_20159,N_13294,N_12622);
or U20160 (N_20160,N_17841,N_15536);
or U20161 (N_20161,N_14101,N_14916);
nand U20162 (N_20162,N_17032,N_13078);
and U20163 (N_20163,N_13129,N_12115);
nor U20164 (N_20164,N_13226,N_17702);
xor U20165 (N_20165,N_17635,N_12420);
or U20166 (N_20166,N_15356,N_14931);
nor U20167 (N_20167,N_12464,N_17312);
nor U20168 (N_20168,N_17539,N_15615);
or U20169 (N_20169,N_15340,N_17591);
xor U20170 (N_20170,N_15043,N_17751);
and U20171 (N_20171,N_17719,N_17937);
or U20172 (N_20172,N_13103,N_13051);
and U20173 (N_20173,N_12008,N_15212);
and U20174 (N_20174,N_16631,N_14875);
or U20175 (N_20175,N_17998,N_17953);
xor U20176 (N_20176,N_13199,N_13895);
nand U20177 (N_20177,N_15849,N_12546);
or U20178 (N_20178,N_16211,N_12398);
and U20179 (N_20179,N_12036,N_12368);
or U20180 (N_20180,N_16244,N_17534);
or U20181 (N_20181,N_15156,N_14103);
nor U20182 (N_20182,N_17248,N_15169);
nor U20183 (N_20183,N_17079,N_15474);
and U20184 (N_20184,N_12403,N_14640);
and U20185 (N_20185,N_13439,N_13622);
and U20186 (N_20186,N_14011,N_12627);
and U20187 (N_20187,N_15971,N_13947);
nor U20188 (N_20188,N_13963,N_13616);
nand U20189 (N_20189,N_16691,N_14829);
nor U20190 (N_20190,N_14951,N_12293);
xor U20191 (N_20191,N_15736,N_14447);
and U20192 (N_20192,N_14663,N_12744);
nor U20193 (N_20193,N_17170,N_14487);
or U20194 (N_20194,N_15900,N_12215);
or U20195 (N_20195,N_13205,N_17128);
nor U20196 (N_20196,N_15669,N_14576);
nor U20197 (N_20197,N_16212,N_15319);
and U20198 (N_20198,N_16535,N_17813);
nand U20199 (N_20199,N_12707,N_17052);
and U20200 (N_20200,N_12283,N_15192);
nand U20201 (N_20201,N_16781,N_12538);
nor U20202 (N_20202,N_17380,N_16948);
xnor U20203 (N_20203,N_12882,N_12674);
nand U20204 (N_20204,N_17231,N_13754);
and U20205 (N_20205,N_17679,N_15506);
nand U20206 (N_20206,N_17807,N_13204);
xor U20207 (N_20207,N_12881,N_13006);
and U20208 (N_20208,N_12586,N_17201);
nor U20209 (N_20209,N_17477,N_12257);
nor U20210 (N_20210,N_12272,N_12182);
nor U20211 (N_20211,N_13766,N_15569);
and U20212 (N_20212,N_14573,N_12162);
and U20213 (N_20213,N_16714,N_15568);
or U20214 (N_20214,N_16541,N_12868);
xor U20215 (N_20215,N_15098,N_15065);
xnor U20216 (N_20216,N_15912,N_16302);
and U20217 (N_20217,N_16829,N_15640);
and U20218 (N_20218,N_14399,N_15555);
or U20219 (N_20219,N_14886,N_17734);
or U20220 (N_20220,N_15739,N_17902);
nor U20221 (N_20221,N_15222,N_17097);
nor U20222 (N_20222,N_14654,N_16160);
nand U20223 (N_20223,N_17295,N_17965);
nand U20224 (N_20224,N_15475,N_13210);
nand U20225 (N_20225,N_15565,N_14694);
xnor U20226 (N_20226,N_17297,N_14740);
nor U20227 (N_20227,N_15316,N_16766);
nand U20228 (N_20228,N_15689,N_15537);
and U20229 (N_20229,N_14230,N_15632);
nand U20230 (N_20230,N_12613,N_16778);
nand U20231 (N_20231,N_15534,N_13421);
or U20232 (N_20232,N_17746,N_13565);
or U20233 (N_20233,N_13461,N_15186);
nor U20234 (N_20234,N_12310,N_14590);
xnor U20235 (N_20235,N_14167,N_13492);
xnor U20236 (N_20236,N_14674,N_13316);
nor U20237 (N_20237,N_12193,N_12922);
or U20238 (N_20238,N_12029,N_14040);
and U20239 (N_20239,N_17304,N_14945);
nand U20240 (N_20240,N_12989,N_14059);
or U20241 (N_20241,N_13220,N_15140);
and U20242 (N_20242,N_15667,N_16279);
or U20243 (N_20243,N_12202,N_14905);
xnor U20244 (N_20244,N_15249,N_15103);
or U20245 (N_20245,N_14368,N_16831);
nor U20246 (N_20246,N_16919,N_16115);
and U20247 (N_20247,N_15591,N_16730);
or U20248 (N_20248,N_13381,N_15430);
nor U20249 (N_20249,N_16864,N_16311);
and U20250 (N_20250,N_17832,N_16800);
or U20251 (N_20251,N_13809,N_12563);
nor U20252 (N_20252,N_16880,N_12497);
nand U20253 (N_20253,N_17444,N_14080);
and U20254 (N_20254,N_16967,N_17753);
and U20255 (N_20255,N_16951,N_12185);
and U20256 (N_20256,N_17058,N_16062);
nand U20257 (N_20257,N_14818,N_12030);
or U20258 (N_20258,N_13131,N_15119);
or U20259 (N_20259,N_12961,N_14975);
nor U20260 (N_20260,N_16566,N_15703);
and U20261 (N_20261,N_16744,N_14734);
or U20262 (N_20262,N_17289,N_15682);
nand U20263 (N_20263,N_15159,N_14249);
nor U20264 (N_20264,N_17950,N_16057);
and U20265 (N_20265,N_17314,N_14837);
nor U20266 (N_20266,N_13623,N_13973);
and U20267 (N_20267,N_14594,N_16727);
and U20268 (N_20268,N_13361,N_12358);
nor U20269 (N_20269,N_13538,N_16725);
or U20270 (N_20270,N_16231,N_17153);
nand U20271 (N_20271,N_13992,N_12071);
nand U20272 (N_20272,N_12266,N_17810);
and U20273 (N_20273,N_17287,N_15493);
and U20274 (N_20274,N_16872,N_12000);
or U20275 (N_20275,N_17575,N_12076);
or U20276 (N_20276,N_14653,N_15664);
nor U20277 (N_20277,N_16939,N_17169);
nor U20278 (N_20278,N_17185,N_12247);
and U20279 (N_20279,N_12469,N_13762);
or U20280 (N_20280,N_17351,N_12826);
nor U20281 (N_20281,N_13178,N_17894);
nand U20282 (N_20282,N_13343,N_14949);
and U20283 (N_20283,N_12644,N_13061);
nand U20284 (N_20284,N_17331,N_14804);
and U20285 (N_20285,N_17948,N_16236);
nand U20286 (N_20286,N_16608,N_14790);
nor U20287 (N_20287,N_16863,N_15177);
nand U20288 (N_20288,N_14119,N_16907);
and U20289 (N_20289,N_16088,N_16360);
or U20290 (N_20290,N_16205,N_16339);
nand U20291 (N_20291,N_14307,N_14204);
or U20292 (N_20292,N_13108,N_12788);
nor U20293 (N_20293,N_13933,N_12381);
or U20294 (N_20294,N_17642,N_15175);
nand U20295 (N_20295,N_12299,N_16366);
xnor U20296 (N_20296,N_12686,N_16775);
nand U20297 (N_20297,N_15497,N_14997);
nand U20298 (N_20298,N_13016,N_14605);
nand U20299 (N_20299,N_13049,N_14211);
xor U20300 (N_20300,N_13753,N_13405);
nor U20301 (N_20301,N_16101,N_12677);
and U20302 (N_20302,N_12648,N_13282);
nor U20303 (N_20303,N_12925,N_12971);
nand U20304 (N_20304,N_14978,N_17941);
or U20305 (N_20305,N_13891,N_13230);
and U20306 (N_20306,N_17142,N_17239);
xnor U20307 (N_20307,N_12952,N_15869);
nand U20308 (N_20308,N_13742,N_16116);
or U20309 (N_20309,N_17917,N_14500);
nor U20310 (N_20310,N_17609,N_14104);
nand U20311 (N_20311,N_13783,N_14980);
and U20312 (N_20312,N_17455,N_14242);
nand U20313 (N_20313,N_17276,N_16186);
nor U20314 (N_20314,N_15725,N_14121);
nor U20315 (N_20315,N_13572,N_13863);
and U20316 (N_20316,N_13785,N_14958);
and U20317 (N_20317,N_16552,N_14518);
and U20318 (N_20318,N_15823,N_15328);
nand U20319 (N_20319,N_13149,N_16172);
and U20320 (N_20320,N_13611,N_12977);
or U20321 (N_20321,N_15883,N_13354);
nand U20322 (N_20322,N_13685,N_16849);
nor U20323 (N_20323,N_15735,N_12120);
and U20324 (N_20324,N_16165,N_13304);
and U20325 (N_20325,N_16767,N_16743);
nor U20326 (N_20326,N_16942,N_17461);
and U20327 (N_20327,N_14296,N_12234);
and U20328 (N_20328,N_15404,N_17846);
nand U20329 (N_20329,N_15214,N_13114);
nor U20330 (N_20330,N_13941,N_13911);
and U20331 (N_20331,N_12321,N_15816);
nor U20332 (N_20332,N_12167,N_12141);
or U20333 (N_20333,N_15561,N_17849);
or U20334 (N_20334,N_15890,N_17947);
or U20335 (N_20335,N_13236,N_14031);
nor U20336 (N_20336,N_16290,N_14574);
nand U20337 (N_20337,N_13636,N_14879);
nand U20338 (N_20338,N_12738,N_14350);
nand U20339 (N_20339,N_13450,N_14781);
nand U20340 (N_20340,N_16719,N_14335);
nand U20341 (N_20341,N_12880,N_12094);
nor U20342 (N_20342,N_14158,N_12473);
nand U20343 (N_20343,N_17581,N_17459);
and U20344 (N_20344,N_13683,N_13923);
and U20345 (N_20345,N_17763,N_17089);
nor U20346 (N_20346,N_12064,N_12772);
and U20347 (N_20347,N_13345,N_16484);
nand U20348 (N_20348,N_17569,N_16487);
nand U20349 (N_20349,N_14300,N_17414);
and U20350 (N_20350,N_15114,N_13527);
xor U20351 (N_20351,N_14414,N_15706);
and U20352 (N_20352,N_17964,N_17050);
nor U20353 (N_20353,N_17673,N_17160);
and U20354 (N_20354,N_12428,N_13838);
nand U20355 (N_20355,N_13706,N_13594);
or U20356 (N_20356,N_15445,N_15144);
nand U20357 (N_20357,N_13353,N_14137);
or U20358 (N_20358,N_14816,N_17480);
nand U20359 (N_20359,N_12558,N_16996);
and U20360 (N_20360,N_16797,N_13383);
or U20361 (N_20361,N_17992,N_12113);
and U20362 (N_20362,N_14629,N_17606);
xor U20363 (N_20363,N_15346,N_17392);
and U20364 (N_20364,N_14317,N_16461);
or U20365 (N_20365,N_14266,N_13455);
or U20366 (N_20366,N_12336,N_17884);
nand U20367 (N_20367,N_14330,N_12710);
nand U20368 (N_20368,N_17410,N_14186);
or U20369 (N_20369,N_16705,N_15803);
or U20370 (N_20370,N_13466,N_16401);
or U20371 (N_20371,N_12083,N_15520);
xnor U20372 (N_20372,N_17750,N_17288);
and U20373 (N_20373,N_13660,N_12478);
nand U20374 (N_20374,N_14582,N_17449);
nand U20375 (N_20375,N_17766,N_16912);
nor U20376 (N_20376,N_16570,N_17361);
and U20377 (N_20377,N_14493,N_16741);
nand U20378 (N_20378,N_12174,N_13385);
nor U20379 (N_20379,N_16479,N_17883);
and U20380 (N_20380,N_15906,N_15075);
nand U20381 (N_20381,N_14070,N_13979);
nand U20382 (N_20382,N_17190,N_15527);
or U20383 (N_20383,N_13774,N_14859);
and U20384 (N_20384,N_16216,N_17887);
or U20385 (N_20385,N_17988,N_12928);
or U20386 (N_20386,N_14731,N_17137);
nand U20387 (N_20387,N_13932,N_16397);
or U20388 (N_20388,N_15123,N_14507);
xor U20389 (N_20389,N_16201,N_13543);
or U20390 (N_20390,N_17048,N_14374);
and U20391 (N_20391,N_17041,N_12747);
nand U20392 (N_20392,N_13934,N_13684);
nand U20393 (N_20393,N_16448,N_16011);
nand U20394 (N_20394,N_17113,N_16222);
xnor U20395 (N_20395,N_12696,N_16399);
nor U20396 (N_20396,N_14870,N_16371);
or U20397 (N_20397,N_14872,N_12787);
nor U20398 (N_20398,N_14395,N_13444);
nand U20399 (N_20399,N_17984,N_12459);
nand U20400 (N_20400,N_12437,N_12060);
and U20401 (N_20401,N_17495,N_16799);
and U20402 (N_20402,N_13971,N_13583);
or U20403 (N_20403,N_14485,N_17156);
nor U20404 (N_20404,N_14239,N_12053);
or U20405 (N_20405,N_17628,N_12931);
xnor U20406 (N_20406,N_15067,N_14929);
or U20407 (N_20407,N_16893,N_15448);
xnor U20408 (N_20408,N_14637,N_16686);
nand U20409 (N_20409,N_13936,N_12070);
nand U20410 (N_20410,N_12711,N_17015);
nor U20411 (N_20411,N_17247,N_17093);
or U20412 (N_20412,N_16578,N_17268);
and U20413 (N_20413,N_16090,N_13998);
or U20414 (N_20414,N_12653,N_15963);
nand U20415 (N_20415,N_16862,N_17682);
nor U20416 (N_20416,N_12553,N_14867);
nand U20417 (N_20417,N_16209,N_14384);
or U20418 (N_20418,N_15986,N_15362);
or U20419 (N_20419,N_15574,N_14362);
and U20420 (N_20420,N_12375,N_15747);
nand U20421 (N_20421,N_14954,N_17675);
nand U20422 (N_20422,N_14353,N_13179);
xor U20423 (N_20423,N_17253,N_14244);
nand U20424 (N_20424,N_17618,N_12290);
and U20425 (N_20425,N_12093,N_13711);
or U20426 (N_20426,N_12618,N_17051);
nor U20427 (N_20427,N_15629,N_13212);
nand U20428 (N_20428,N_17959,N_12096);
nor U20429 (N_20429,N_14819,N_17886);
and U20430 (N_20430,N_15233,N_16507);
or U20431 (N_20431,N_13851,N_13879);
nor U20432 (N_20432,N_15252,N_16590);
nor U20433 (N_20433,N_12061,N_13822);
and U20434 (N_20434,N_16609,N_12220);
or U20435 (N_20435,N_15505,N_14589);
or U20436 (N_20436,N_13921,N_14546);
or U20437 (N_20437,N_16200,N_16925);
and U20438 (N_20438,N_12802,N_13489);
or U20439 (N_20439,N_13590,N_16881);
nand U20440 (N_20440,N_16840,N_12402);
xor U20441 (N_20441,N_15331,N_13372);
nor U20442 (N_20442,N_14450,N_13303);
or U20443 (N_20443,N_12919,N_17736);
xnor U20444 (N_20444,N_16368,N_17520);
nand U20445 (N_20445,N_15081,N_12037);
xnor U20446 (N_20446,N_15671,N_13651);
nor U20447 (N_20447,N_15129,N_14659);
or U20448 (N_20448,N_15819,N_17836);
nand U20449 (N_20449,N_16875,N_16892);
and U20450 (N_20450,N_13423,N_12715);
xor U20451 (N_20451,N_12552,N_15202);
nor U20452 (N_20452,N_14367,N_12287);
and U20453 (N_20453,N_14032,N_14477);
and U20454 (N_20454,N_13027,N_12419);
xnor U20455 (N_20455,N_13096,N_17655);
or U20456 (N_20456,N_16969,N_17010);
or U20457 (N_20457,N_12947,N_15701);
and U20458 (N_20458,N_17102,N_16953);
nand U20459 (N_20459,N_13284,N_12353);
nor U20460 (N_20460,N_17068,N_12409);
and U20461 (N_20461,N_12068,N_17003);
and U20462 (N_20462,N_14113,N_16987);
nor U20463 (N_20463,N_17919,N_13510);
nor U20464 (N_20464,N_17578,N_17946);
or U20465 (N_20465,N_16276,N_14423);
and U20466 (N_20466,N_14496,N_15934);
nand U20467 (N_20467,N_14709,N_14498);
nor U20468 (N_20468,N_12941,N_15970);
nand U20469 (N_20469,N_15777,N_15227);
or U20470 (N_20470,N_16606,N_12800);
or U20471 (N_20471,N_12369,N_13425);
nand U20472 (N_20472,N_13173,N_12451);
or U20473 (N_20473,N_16018,N_12842);
nand U20474 (N_20474,N_16373,N_15490);
or U20475 (N_20475,N_13395,N_16836);
nor U20476 (N_20476,N_14118,N_14986);
nand U20477 (N_20477,N_13101,N_13526);
nand U20478 (N_20478,N_15312,N_16008);
or U20479 (N_20479,N_12163,N_14611);
nor U20480 (N_20480,N_17930,N_13264);
nor U20481 (N_20481,N_13019,N_13422);
nor U20482 (N_20482,N_12382,N_15891);
nor U20483 (N_20483,N_14183,N_14869);
nand U20484 (N_20484,N_17584,N_16335);
and U20485 (N_20485,N_13014,N_12778);
nor U20486 (N_20486,N_12742,N_15421);
nand U20487 (N_20487,N_14228,N_12755);
xnor U20488 (N_20488,N_16056,N_16070);
nor U20489 (N_20489,N_12050,N_12735);
nand U20490 (N_20490,N_12837,N_16117);
or U20491 (N_20491,N_16512,N_17851);
nor U20492 (N_20492,N_14840,N_13884);
xnor U20493 (N_20493,N_17294,N_15369);
nand U20494 (N_20494,N_13535,N_16059);
nor U20495 (N_20495,N_13605,N_16592);
and U20496 (N_20496,N_14309,N_16382);
nor U20497 (N_20497,N_17833,N_13060);
nor U20498 (N_20498,N_13259,N_16127);
and U20499 (N_20499,N_15880,N_16702);
and U20500 (N_20500,N_14005,N_12134);
and U20501 (N_20501,N_13365,N_17109);
xnor U20502 (N_20502,N_13415,N_16322);
nand U20503 (N_20503,N_16700,N_13638);
nand U20504 (N_20504,N_17889,N_12610);
nor U20505 (N_20505,N_16021,N_17681);
nor U20506 (N_20506,N_13702,N_16666);
xor U20507 (N_20507,N_15300,N_15315);
xor U20508 (N_20508,N_17208,N_12520);
nor U20509 (N_20509,N_15386,N_16245);
or U20510 (N_20510,N_12264,N_17557);
and U20511 (N_20511,N_17527,N_17644);
or U20512 (N_20512,N_16220,N_15388);
nor U20513 (N_20513,N_14965,N_15824);
nand U20514 (N_20514,N_13858,N_16296);
nor U20515 (N_20515,N_12764,N_12223);
xor U20516 (N_20516,N_14049,N_14686);
or U20517 (N_20517,N_14808,N_17307);
nand U20518 (N_20518,N_12018,N_15238);
or U20519 (N_20519,N_15417,N_17496);
or U20520 (N_20520,N_15709,N_16663);
nand U20521 (N_20521,N_15817,N_15733);
nand U20522 (N_20522,N_14891,N_12043);
nor U20523 (N_20523,N_14004,N_12286);
or U20524 (N_20524,N_13661,N_16914);
or U20525 (N_20525,N_13849,N_14724);
nor U20526 (N_20526,N_12509,N_16048);
xor U20527 (N_20527,N_13869,N_12416);
nor U20528 (N_20528,N_16545,N_17448);
nor U20529 (N_20529,N_13688,N_13805);
nor U20530 (N_20530,N_16768,N_12729);
nand U20531 (N_20531,N_12421,N_14189);
nand U20532 (N_20532,N_16138,N_14132);
and U20533 (N_20533,N_16263,N_13791);
nor U20534 (N_20534,N_13607,N_12740);
nand U20535 (N_20535,N_14305,N_15303);
xor U20536 (N_20536,N_13552,N_14003);
and U20537 (N_20537,N_17670,N_13416);
xnor U20538 (N_20538,N_15347,N_15259);
nor U20539 (N_20539,N_14250,N_13634);
and U20540 (N_20540,N_16964,N_16012);
and U20541 (N_20541,N_14396,N_15668);
nor U20542 (N_20542,N_13999,N_12765);
nand U20543 (N_20543,N_13133,N_13188);
nor U20544 (N_20544,N_17432,N_12418);
and U20545 (N_20545,N_17594,N_16934);
nand U20546 (N_20546,N_15213,N_14086);
or U20547 (N_20547,N_12924,N_15661);
nor U20548 (N_20548,N_17494,N_14081);
nor U20549 (N_20549,N_12441,N_13201);
and U20550 (N_20550,N_12864,N_17424);
or U20551 (N_20551,N_12893,N_14269);
and U20552 (N_20552,N_16147,N_15965);
nor U20553 (N_20553,N_16652,N_14483);
nand U20554 (N_20554,N_17164,N_12195);
nand U20555 (N_20555,N_13962,N_12089);
nor U20556 (N_20556,N_17881,N_16242);
xnor U20557 (N_20557,N_12833,N_13263);
nor U20558 (N_20558,N_13434,N_15250);
and U20559 (N_20559,N_15864,N_17014);
nor U20560 (N_20560,N_13453,N_16838);
nor U20561 (N_20561,N_16035,N_17111);
or U20562 (N_20562,N_13157,N_17739);
nor U20563 (N_20563,N_14408,N_16343);
or U20564 (N_20564,N_15171,N_14529);
or U20565 (N_20565,N_15954,N_13599);
nor U20566 (N_20566,N_12450,N_14586);
or U20567 (N_20567,N_13473,N_17788);
or U20568 (N_20568,N_15861,N_12609);
and U20569 (N_20569,N_15693,N_13359);
and U20570 (N_20570,N_12033,N_16073);
nand U20571 (N_20571,N_14278,N_13768);
nor U20572 (N_20572,N_14120,N_16859);
and U20573 (N_20573,N_17382,N_13160);
xor U20574 (N_20574,N_17641,N_15639);
nor U20575 (N_20575,N_16167,N_16918);
nor U20576 (N_20576,N_13567,N_17678);
and U20577 (N_20577,N_16834,N_16403);
and U20578 (N_20578,N_16521,N_17524);
nand U20579 (N_20579,N_15379,N_12274);
nand U20580 (N_20580,N_14793,N_12680);
or U20581 (N_20581,N_16740,N_13093);
or U20582 (N_20582,N_15885,N_13876);
xnor U20583 (N_20583,N_15674,N_14282);
and U20584 (N_20584,N_17112,N_12335);
or U20585 (N_20585,N_15746,N_12306);
nor U20586 (N_20586,N_13356,N_13233);
and U20587 (N_20587,N_16682,N_12926);
xor U20588 (N_20588,N_14345,N_15073);
nand U20589 (N_20589,N_13871,N_17167);
and U20590 (N_20590,N_14509,N_13970);
and U20591 (N_20591,N_16477,N_17360);
and U20592 (N_20592,N_16433,N_12722);
nor U20593 (N_20593,N_12796,N_17205);
nand U20594 (N_20594,N_15160,N_13278);
nand U20595 (N_20595,N_14504,N_17730);
xor U20596 (N_20596,N_14535,N_15853);
nor U20597 (N_20597,N_15765,N_15275);
or U20598 (N_20598,N_15724,N_12559);
and U20599 (N_20599,N_13104,N_13228);
xnor U20600 (N_20600,N_14402,N_16646);
or U20601 (N_20601,N_15009,N_17191);
or U20602 (N_20602,N_12705,N_13532);
nand U20603 (N_20603,N_12885,N_14927);
xor U20604 (N_20604,N_12020,N_17255);
or U20605 (N_20605,N_17933,N_13420);
or U20606 (N_20606,N_14785,N_15314);
nand U20607 (N_20607,N_12180,N_13795);
nand U20608 (N_20608,N_15921,N_14391);
and U20609 (N_20609,N_12824,N_12146);
and U20610 (N_20610,N_17075,N_16445);
nand U20611 (N_20611,N_16680,N_12341);
nor U20612 (N_20612,N_12151,N_16830);
and U20613 (N_20613,N_15108,N_16492);
or U20614 (N_20614,N_13277,N_16820);
nor U20615 (N_20615,N_14665,N_15932);
nor U20616 (N_20616,N_16871,N_15592);
and U20617 (N_20617,N_16327,N_17082);
nand U20618 (N_20618,N_13922,N_17722);
nor U20619 (N_20619,N_15916,N_17970);
nor U20620 (N_20620,N_13299,N_13528);
and U20621 (N_20621,N_15485,N_14495);
nor U20622 (N_20622,N_12786,N_13363);
nor U20623 (N_20623,N_14018,N_16921);
or U20624 (N_20624,N_15425,N_14199);
xnor U20625 (N_20625,N_15071,N_15139);
or U20626 (N_20626,N_13349,N_12861);
nand U20627 (N_20627,N_15691,N_17564);
nand U20628 (N_20628,N_15030,N_17796);
nand U20629 (N_20629,N_12455,N_14899);
nor U20630 (N_20630,N_14750,N_16782);
and U20631 (N_20631,N_17680,N_16604);
nand U20632 (N_20632,N_14920,N_17130);
or U20633 (N_20633,N_14568,N_13695);
nor U20634 (N_20634,N_12944,N_17228);
and U20635 (N_20635,N_15094,N_16005);
or U20636 (N_20636,N_13553,N_15967);
nand U20637 (N_20637,N_15850,N_13930);
and U20638 (N_20638,N_16135,N_16099);
or U20639 (N_20639,N_13465,N_16685);
or U20640 (N_20640,N_14068,N_16202);
nand U20641 (N_20641,N_16968,N_17621);
nor U20642 (N_20642,N_15434,N_12239);
nand U20643 (N_20643,N_17281,N_13368);
nand U20644 (N_20644,N_12682,N_17300);
nor U20645 (N_20645,N_14897,N_17422);
nand U20646 (N_20646,N_12814,N_17029);
nand U20647 (N_20647,N_13788,N_15980);
or U20648 (N_20648,N_12942,N_15180);
nor U20649 (N_20649,N_15255,N_16742);
and U20650 (N_20650,N_13699,N_13874);
nor U20651 (N_20651,N_13094,N_13873);
nand U20652 (N_20652,N_14254,N_13137);
nand U20653 (N_20653,N_17876,N_15994);
or U20654 (N_20654,N_15797,N_16534);
nand U20655 (N_20655,N_12821,N_12386);
nand U20656 (N_20656,N_13091,N_15479);
and U20657 (N_20657,N_14260,N_16899);
nand U20658 (N_20658,N_15333,N_13432);
nand U20659 (N_20659,N_16752,N_16462);
nor U20660 (N_20660,N_17342,N_13144);
xnor U20661 (N_20661,N_16619,N_14435);
xor U20662 (N_20662,N_15461,N_15393);
xnor U20663 (N_20663,N_15680,N_17470);
nand U20664 (N_20664,N_12224,N_12531);
nor U20665 (N_20665,N_16959,N_13517);
or U20666 (N_20666,N_16255,N_16756);
nor U20667 (N_20667,N_12231,N_14141);
or U20668 (N_20668,N_12059,N_12468);
and U20669 (N_20669,N_13772,N_16481);
nand U20670 (N_20670,N_17560,N_16338);
nand U20671 (N_20671,N_14878,N_16473);
nor U20672 (N_20672,N_14993,N_13336);
and U20673 (N_20673,N_14321,N_14441);
nand U20674 (N_20674,N_16990,N_17078);
and U20675 (N_20675,N_12281,N_17874);
xnor U20676 (N_20676,N_13247,N_13314);
or U20677 (N_20677,N_16137,N_13295);
nor U20678 (N_20678,N_12326,N_12831);
nor U20679 (N_20679,N_15176,N_14739);
or U20680 (N_20680,N_15277,N_15311);
nand U20681 (N_20681,N_17658,N_15464);
nor U20682 (N_20682,N_13100,N_15756);
nand U20683 (N_20683,N_13604,N_13806);
or U20684 (N_20684,N_17244,N_12026);
and U20685 (N_20685,N_12277,N_14752);
and U20686 (N_20686,N_16446,N_15082);
xnor U20687 (N_20687,N_14720,N_12208);
nand U20688 (N_20688,N_17645,N_16650);
nand U20689 (N_20689,N_17996,N_13540);
nor U20690 (N_20690,N_14558,N_16175);
or U20691 (N_20691,N_12021,N_16674);
or U20692 (N_20692,N_13331,N_15556);
nand U20693 (N_20693,N_13433,N_17038);
nor U20694 (N_20694,N_13746,N_16490);
nor U20695 (N_20695,N_16416,N_14265);
xor U20696 (N_20696,N_15813,N_16988);
and U20697 (N_20697,N_14146,N_17241);
and U20698 (N_20698,N_12741,N_15599);
xor U20699 (N_20699,N_12543,N_14270);
nand U20700 (N_20700,N_16087,N_17463);
nand U20701 (N_20701,N_13219,N_16506);
and U20702 (N_20702,N_16614,N_17559);
and U20703 (N_20703,N_12444,N_14380);
nor U20704 (N_20704,N_12474,N_12631);
xor U20705 (N_20705,N_12726,N_17683);
and U20706 (N_20706,N_15121,N_13780);
nor U20707 (N_20707,N_15526,N_13566);
xor U20708 (N_20708,N_17115,N_15210);
nand U20709 (N_20709,N_17460,N_16979);
nand U20710 (N_20710,N_13021,N_16058);
nor U20711 (N_20711,N_14933,N_15117);
nor U20712 (N_20712,N_17797,N_14140);
nor U20713 (N_20713,N_13563,N_15799);
or U20714 (N_20714,N_14821,N_13379);
nor U20715 (N_20715,N_17729,N_17913);
nand U20716 (N_20716,N_16113,N_13969);
and U20717 (N_20717,N_12074,N_14991);
xor U20718 (N_20718,N_12874,N_15613);
or U20719 (N_20719,N_16699,N_16574);
nand U20720 (N_20720,N_15805,N_16597);
nor U20721 (N_20721,N_15230,N_17356);
nor U20722 (N_20722,N_15871,N_17706);
or U20723 (N_20723,N_13396,N_13585);
nor U20724 (N_20724,N_15985,N_13845);
nor U20725 (N_20725,N_15557,N_13238);
nand U20726 (N_20726,N_12600,N_16932);
nor U20727 (N_20727,N_12347,N_13896);
and U20728 (N_20728,N_14595,N_17994);
xor U20729 (N_20729,N_13221,N_17624);
or U20730 (N_20730,N_12143,N_14768);
and U20731 (N_20731,N_14633,N_12780);
or U20732 (N_20732,N_14226,N_13009);
nand U20733 (N_20733,N_16896,N_13138);
or U20734 (N_20734,N_17491,N_13861);
and U20735 (N_20735,N_16555,N_15059);
or U20736 (N_20736,N_14351,N_16234);
or U20737 (N_20737,N_17663,N_13734);
or U20738 (N_20738,N_16443,N_16493);
nor U20739 (N_20739,N_13701,N_15848);
xor U20740 (N_20740,N_16459,N_15581);
or U20741 (N_20741,N_16125,N_12054);
or U20742 (N_20742,N_15795,N_12850);
nor U20743 (N_20743,N_16206,N_15827);
or U20744 (N_20744,N_16586,N_16955);
xor U20745 (N_20745,N_14501,N_12001);
or U20746 (N_20746,N_14528,N_14373);
nor U20747 (N_20747,N_17566,N_12256);
nand U20748 (N_20748,N_17685,N_17995);
or U20749 (N_20749,N_16271,N_14098);
or U20750 (N_20750,N_15240,N_13976);
and U20751 (N_20751,N_15949,N_17989);
and U20752 (N_20752,N_14170,N_17707);
or U20753 (N_20753,N_15753,N_16284);
xor U20754 (N_20754,N_17259,N_13118);
and U20755 (N_20755,N_17877,N_15147);
or U20756 (N_20756,N_13127,N_15688);
and U20757 (N_20757,N_17548,N_15344);
nor U20758 (N_20758,N_14424,N_13280);
nand U20759 (N_20759,N_16123,N_17475);
nor U20760 (N_20760,N_16909,N_12186);
nand U20761 (N_20761,N_12393,N_15684);
nor U20762 (N_20762,N_15946,N_12891);
and U20763 (N_20763,N_14766,N_16354);
nor U20764 (N_20764,N_14216,N_16077);
and U20765 (N_20765,N_12311,N_17054);
and U20766 (N_20766,N_14238,N_15628);
nor U20767 (N_20767,N_12169,N_12384);
or U20768 (N_20768,N_14133,N_16779);
and U20769 (N_20769,N_16210,N_15902);
or U20770 (N_20770,N_17434,N_14770);
or U20771 (N_20771,N_12576,N_13931);
nor U20772 (N_20772,N_14190,N_16821);
nand U20773 (N_20773,N_15874,N_13362);
and U20774 (N_20774,N_13635,N_17825);
nand U20775 (N_20775,N_16723,N_12031);
or U20776 (N_20776,N_13045,N_12999);
or U20777 (N_20777,N_17400,N_16930);
nor U20778 (N_20778,N_16157,N_14671);
nand U20779 (N_20779,N_17403,N_17726);
nand U20780 (N_20780,N_15350,N_12579);
and U20781 (N_20781,N_17714,N_14812);
nor U20782 (N_20782,N_12453,N_17541);
nor U20783 (N_20783,N_14716,N_14871);
xor U20784 (N_20784,N_17166,N_15492);
or U20785 (N_20785,N_16747,N_17353);
or U20786 (N_20786,N_12905,N_12988);
nand U20787 (N_20787,N_15832,N_14333);
nand U20788 (N_20788,N_16833,N_17771);
nor U20789 (N_20789,N_15636,N_13593);
nor U20790 (N_20790,N_16476,N_12667);
nor U20791 (N_20791,N_12623,N_12229);
nor U20792 (N_20792,N_17563,N_13341);
xnor U20793 (N_20793,N_15339,N_13828);
nand U20794 (N_20794,N_13994,N_15920);
nand U20795 (N_20795,N_13497,N_13033);
or U20796 (N_20796,N_12267,N_13404);
or U20797 (N_20797,N_16733,N_17850);
xnor U20798 (N_20798,N_14152,N_13900);
xor U20799 (N_20799,N_15298,N_12642);
or U20800 (N_20800,N_12573,N_13981);
nor U20801 (N_20801,N_16908,N_14627);
nand U20802 (N_20802,N_14613,N_16149);
or U20803 (N_20803,N_16938,N_15851);
nand U20804 (N_20804,N_16447,N_16560);
xnor U20805 (N_20805,N_16199,N_16174);
nand U20806 (N_20806,N_16439,N_12541);
and U20807 (N_20807,N_16518,N_12946);
nand U20808 (N_20808,N_15487,N_17842);
nand U20809 (N_20809,N_14095,N_14909);
nor U20810 (N_20810,N_16419,N_13251);
xnor U20811 (N_20811,N_13317,N_17323);
xor U20812 (N_20812,N_14634,N_12591);
nor U20813 (N_20813,N_13718,N_16770);
and U20814 (N_20814,N_14090,N_15517);
nor U20815 (N_20815,N_16268,N_14857);
or U20816 (N_20816,N_16140,N_14217);
nor U20817 (N_20817,N_13115,N_15292);
nand U20818 (N_20818,N_14852,N_17453);
xnor U20819 (N_20819,N_14327,N_13722);
and U20820 (N_20820,N_17348,N_17529);
nor U20821 (N_20821,N_15097,N_13885);
or U20822 (N_20822,N_16585,N_13366);
xnor U20823 (N_20823,N_17390,N_16851);
and U20824 (N_20824,N_13159,N_12449);
nor U20825 (N_20825,N_12192,N_13250);
nor U20826 (N_20826,N_12170,N_14225);
or U20827 (N_20827,N_16576,N_17210);
nand U20828 (N_20828,N_13539,N_17549);
nor U20829 (N_20829,N_12117,N_15481);
or U20830 (N_20830,N_15220,N_17600);
nand U20831 (N_20831,N_13002,N_16915);
and U20832 (N_20832,N_12529,N_16580);
xnor U20833 (N_20833,N_15405,N_16424);
nand U20834 (N_20834,N_12122,N_16869);
or U20835 (N_20835,N_15352,N_17364);
xor U20836 (N_20836,N_12968,N_16669);
xor U20837 (N_20837,N_16333,N_16783);
nor U20838 (N_20838,N_17026,N_16034);
xnor U20839 (N_20839,N_17588,N_13549);
and U20840 (N_20840,N_17385,N_13064);
nand U20841 (N_20841,N_12407,N_12953);
nand U20842 (N_20842,N_17059,N_16226);
and U20843 (N_20843,N_17110,N_16698);
nand U20844 (N_20844,N_15070,N_16906);
and U20845 (N_20845,N_17375,N_14838);
or U20846 (N_20846,N_14100,N_14466);
or U20847 (N_20847,N_16754,N_15673);
and U20848 (N_20848,N_15440,N_13056);
nand U20849 (N_20849,N_12575,N_16654);
and U20850 (N_20850,N_12385,N_15069);
nand U20851 (N_20851,N_14516,N_15966);
or U20852 (N_20852,N_17273,N_15845);
and U20853 (N_20853,N_16717,N_16977);
nor U20854 (N_20854,N_14022,N_13880);
nand U20855 (N_20855,N_12936,N_16516);
and U20856 (N_20856,N_12532,N_17577);
nand U20857 (N_20857,N_13817,N_14135);
nor U20858 (N_20858,N_16221,N_17525);
nor U20859 (N_20859,N_13586,N_17669);
nor U20860 (N_20860,N_17835,N_15482);
and U20861 (N_20861,N_14324,N_13580);
nor U20862 (N_20862,N_17291,N_12830);
nor U20863 (N_20863,N_15013,N_14848);
or U20864 (N_20864,N_17411,N_13747);
or U20865 (N_20865,N_17583,N_12447);
or U20866 (N_20866,N_12544,N_14197);
nand U20867 (N_20867,N_14108,N_16387);
and U20868 (N_20868,N_13529,N_15343);
xnor U20869 (N_20869,N_12343,N_12706);
or U20870 (N_20870,N_13476,N_14703);
and U20871 (N_20871,N_17742,N_17278);
nor U20872 (N_20872,N_12938,N_14026);
and U20873 (N_20873,N_15099,N_12365);
and U20874 (N_20874,N_15571,N_13993);
or U20875 (N_20875,N_15024,N_17918);
and U20876 (N_20876,N_15785,N_12991);
nand U20877 (N_20877,N_16060,N_17071);
or U20878 (N_20878,N_13158,N_14757);
nor U20879 (N_20879,N_13430,N_14907);
and U20880 (N_20880,N_13106,N_16999);
xnor U20881 (N_20881,N_16337,N_14861);
and U20882 (N_20882,N_14526,N_16026);
and U20883 (N_20883,N_15426,N_14503);
and U20884 (N_20884,N_16634,N_17602);
and U20885 (N_20885,N_16594,N_12213);
nor U20886 (N_20886,N_14271,N_12972);
and U20887 (N_20887,N_15301,N_13169);
nand U20888 (N_20888,N_12380,N_16856);
and U20889 (N_20889,N_12791,N_15953);
or U20890 (N_20890,N_12806,N_15732);
nor U20891 (N_20891,N_15499,N_15955);
nor U20892 (N_20892,N_15368,N_14601);
nand U20893 (N_20893,N_14902,N_13960);
nand U20894 (N_20894,N_12884,N_14572);
or U20895 (N_20895,N_17962,N_15197);
nand U20896 (N_20896,N_14698,N_14318);
nor U20897 (N_20897,N_12106,N_17184);
nor U20898 (N_20898,N_15504,N_17347);
nand U20899 (N_20899,N_15987,N_14971);
and U20900 (N_20900,N_15979,N_12684);
nand U20901 (N_20901,N_17316,N_17450);
or U20902 (N_20902,N_15738,N_15647);
and U20903 (N_20903,N_15781,N_14079);
nand U20904 (N_20904,N_13912,N_15450);
nor U20905 (N_20905,N_14415,N_12770);
nand U20906 (N_20906,N_17338,N_14964);
and U20907 (N_20907,N_17465,N_13678);
nand U20908 (N_20908,N_16441,N_14474);
nand U20909 (N_20909,N_16000,N_16028);
nand U20910 (N_20910,N_15931,N_12877);
nand U20911 (N_20911,N_15002,N_14845);
nand U20912 (N_20912,N_17693,N_15783);
xnor U20913 (N_20913,N_14039,N_17695);
nor U20914 (N_20914,N_16630,N_16061);
nor U20915 (N_20915,N_12148,N_15491);
and U20916 (N_20916,N_15188,N_17357);
or U20917 (N_20917,N_12608,N_17260);
and U20918 (N_20918,N_13288,N_15730);
and U20919 (N_20919,N_12135,N_15477);
and U20920 (N_20920,N_17823,N_16063);
and U20921 (N_20921,N_14618,N_12656);
and U20922 (N_20922,N_17715,N_16530);
and U20923 (N_20923,N_15391,N_14025);
and U20924 (N_20924,N_16489,N_16718);
nand U20925 (N_20925,N_13223,N_13741);
and U20926 (N_20926,N_14169,N_16474);
or U20927 (N_20927,N_14013,N_17468);
and U20928 (N_20928,N_14176,N_15515);
xor U20929 (N_20929,N_17901,N_14806);
and U20930 (N_20930,N_17582,N_13044);
nand U20931 (N_20931,N_13898,N_13512);
nor U20932 (N_20932,N_17301,N_15138);
and U20933 (N_20933,N_16637,N_15770);
or U20934 (N_20934,N_13112,N_12161);
nand U20935 (N_20935,N_14865,N_15457);
nor U20936 (N_20936,N_15442,N_13386);
and U20937 (N_20937,N_17229,N_17518);
nand U20938 (N_20938,N_17927,N_13155);
and U20939 (N_20939,N_14115,N_16092);
and U20940 (N_20940,N_15815,N_12506);
or U20941 (N_20941,N_15609,N_14919);
and U20942 (N_20942,N_16678,N_13883);
nand U20943 (N_20943,N_17308,N_17631);
or U20944 (N_20944,N_12920,N_15731);
nand U20945 (N_20945,N_16603,N_17971);
nor U20946 (N_20946,N_15695,N_16693);
nand U20947 (N_20947,N_16071,N_17310);
or U20948 (N_20948,N_13901,N_13514);
nand U20949 (N_20949,N_17379,N_15708);
nor U20950 (N_20950,N_16345,N_16916);
and U20951 (N_20951,N_12414,N_17980);
nor U20952 (N_20952,N_14084,N_16161);
nand U20953 (N_20953,N_14761,N_12406);
nor U20954 (N_20954,N_13700,N_12221);
and U20955 (N_20955,N_17666,N_16243);
and U20956 (N_20956,N_14102,N_12853);
nand U20957 (N_20957,N_15453,N_14182);
or U20958 (N_20958,N_16974,N_14312);
or U20959 (N_20959,N_14181,N_15807);
and U20960 (N_20960,N_15876,N_12829);
or U20961 (N_20961,N_17224,N_14442);
or U20962 (N_20962,N_12052,N_12047);
and U20963 (N_20963,N_12032,N_17978);
and U20964 (N_20964,N_14184,N_17982);
xnor U20965 (N_20965,N_12766,N_12678);
and U20966 (N_20966,N_15109,N_13070);
nand U20967 (N_20967,N_16995,N_17081);
nand U20968 (N_20968,N_13124,N_12483);
or U20969 (N_20969,N_15272,N_16204);
nand U20970 (N_20970,N_17708,N_17731);
nand U20971 (N_20971,N_15518,N_12006);
xnor U20972 (N_20972,N_13698,N_16313);
or U20973 (N_20973,N_15308,N_13624);
xnor U20974 (N_20974,N_14616,N_13183);
xnor U20975 (N_20975,N_16715,N_16651);
xor U20976 (N_20976,N_12595,N_14129);
nor U20977 (N_20977,N_13555,N_13252);
nor U20978 (N_20978,N_16287,N_14174);
nand U20979 (N_20979,N_15234,N_16565);
or U20980 (N_20980,N_17046,N_16309);
nor U20981 (N_20981,N_17510,N_15020);
or U20982 (N_20982,N_17711,N_12370);
or U20983 (N_20983,N_16141,N_16588);
or U20984 (N_20984,N_14581,N_12875);
nor U20985 (N_20985,N_13697,N_16417);
and U20986 (N_20986,N_12475,N_15335);
or U20987 (N_20987,N_14712,N_15600);
nor U20988 (N_20988,N_12590,N_13997);
nor U20989 (N_20989,N_15241,N_12515);
nor U20990 (N_20990,N_16954,N_15660);
nand U20991 (N_20991,N_14868,N_14406);
nand U20992 (N_20992,N_15288,N_14693);
xnor U20993 (N_20993,N_12241,N_16320);
nor U20994 (N_20994,N_16501,N_16191);
and U20995 (N_20995,N_12597,N_16858);
nand U20996 (N_20996,N_14303,N_16917);
nor U20997 (N_20997,N_14016,N_16679);
nand U20998 (N_20998,N_17676,N_12986);
nor U20999 (N_20999,N_16984,N_13265);
nor U21000 (N_21000,N_13971,N_16155);
nor U21001 (N_21001,N_14764,N_17275);
nand U21002 (N_21002,N_13015,N_12357);
or U21003 (N_21003,N_17337,N_16534);
and U21004 (N_21004,N_14370,N_14426);
and U21005 (N_21005,N_13383,N_14990);
or U21006 (N_21006,N_16440,N_16616);
and U21007 (N_21007,N_12444,N_14249);
xor U21008 (N_21008,N_16433,N_16643);
nand U21009 (N_21009,N_17086,N_13957);
or U21010 (N_21010,N_16493,N_12225);
and U21011 (N_21011,N_16440,N_12103);
and U21012 (N_21012,N_15323,N_12064);
nand U21013 (N_21013,N_14139,N_16860);
nor U21014 (N_21014,N_17188,N_13308);
nor U21015 (N_21015,N_16100,N_15743);
and U21016 (N_21016,N_17982,N_14875);
nor U21017 (N_21017,N_14947,N_15737);
nand U21018 (N_21018,N_16257,N_12991);
xnor U21019 (N_21019,N_17463,N_14524);
nand U21020 (N_21020,N_17652,N_16669);
xnor U21021 (N_21021,N_12690,N_12763);
nor U21022 (N_21022,N_14921,N_13231);
or U21023 (N_21023,N_16070,N_16216);
nor U21024 (N_21024,N_16582,N_17998);
nor U21025 (N_21025,N_13089,N_17545);
and U21026 (N_21026,N_15723,N_17660);
and U21027 (N_21027,N_13080,N_16084);
and U21028 (N_21028,N_14580,N_16422);
xnor U21029 (N_21029,N_16285,N_13300);
nand U21030 (N_21030,N_17322,N_17966);
or U21031 (N_21031,N_12857,N_16215);
and U21032 (N_21032,N_15822,N_17296);
or U21033 (N_21033,N_13854,N_12162);
and U21034 (N_21034,N_17462,N_14086);
or U21035 (N_21035,N_15726,N_16281);
and U21036 (N_21036,N_14827,N_13312);
xor U21037 (N_21037,N_12650,N_13715);
and U21038 (N_21038,N_14319,N_15135);
nor U21039 (N_21039,N_14902,N_15410);
nor U21040 (N_21040,N_16394,N_15057);
or U21041 (N_21041,N_16780,N_14583);
nand U21042 (N_21042,N_17905,N_15285);
or U21043 (N_21043,N_13418,N_15185);
and U21044 (N_21044,N_15962,N_13661);
nor U21045 (N_21045,N_16692,N_14469);
nor U21046 (N_21046,N_15197,N_17224);
or U21047 (N_21047,N_16503,N_16702);
nand U21048 (N_21048,N_17352,N_12131);
or U21049 (N_21049,N_12662,N_17027);
nand U21050 (N_21050,N_14157,N_17606);
or U21051 (N_21051,N_14669,N_13382);
nand U21052 (N_21052,N_12773,N_15547);
or U21053 (N_21053,N_17563,N_17802);
or U21054 (N_21054,N_17472,N_14479);
nand U21055 (N_21055,N_12455,N_17692);
or U21056 (N_21056,N_14607,N_17456);
or U21057 (N_21057,N_17991,N_12932);
and U21058 (N_21058,N_16888,N_12303);
and U21059 (N_21059,N_15922,N_17197);
and U21060 (N_21060,N_15771,N_16088);
or U21061 (N_21061,N_13355,N_15887);
and U21062 (N_21062,N_15039,N_12625);
nor U21063 (N_21063,N_17665,N_14776);
xnor U21064 (N_21064,N_14007,N_12753);
xnor U21065 (N_21065,N_17483,N_17142);
or U21066 (N_21066,N_13378,N_16059);
nor U21067 (N_21067,N_17762,N_13660);
nor U21068 (N_21068,N_12619,N_12503);
and U21069 (N_21069,N_13226,N_14208);
or U21070 (N_21070,N_16011,N_14438);
xor U21071 (N_21071,N_17161,N_16499);
xor U21072 (N_21072,N_14273,N_16224);
nand U21073 (N_21073,N_14026,N_15538);
and U21074 (N_21074,N_13479,N_16223);
nor U21075 (N_21075,N_17157,N_14283);
or U21076 (N_21076,N_15824,N_17514);
nor U21077 (N_21077,N_13863,N_16777);
or U21078 (N_21078,N_12639,N_12732);
and U21079 (N_21079,N_14904,N_17210);
xnor U21080 (N_21080,N_16877,N_15487);
or U21081 (N_21081,N_13036,N_12201);
xnor U21082 (N_21082,N_14801,N_12036);
xor U21083 (N_21083,N_16025,N_13253);
nand U21084 (N_21084,N_17996,N_17522);
xnor U21085 (N_21085,N_16739,N_15389);
nor U21086 (N_21086,N_17860,N_15003);
nand U21087 (N_21087,N_16796,N_15024);
nor U21088 (N_21088,N_12204,N_12146);
xor U21089 (N_21089,N_12351,N_14257);
nor U21090 (N_21090,N_15284,N_17203);
or U21091 (N_21091,N_14950,N_12411);
nand U21092 (N_21092,N_15921,N_15602);
nand U21093 (N_21093,N_17591,N_14498);
nor U21094 (N_21094,N_15756,N_13028);
nor U21095 (N_21095,N_13966,N_14148);
nand U21096 (N_21096,N_12481,N_12944);
xnor U21097 (N_21097,N_12688,N_12221);
nand U21098 (N_21098,N_13846,N_12149);
nand U21099 (N_21099,N_13956,N_12979);
and U21100 (N_21100,N_14137,N_17766);
or U21101 (N_21101,N_13069,N_14548);
and U21102 (N_21102,N_17042,N_15835);
nor U21103 (N_21103,N_14567,N_12102);
or U21104 (N_21104,N_15089,N_15632);
or U21105 (N_21105,N_12016,N_16490);
nand U21106 (N_21106,N_14292,N_12934);
or U21107 (N_21107,N_14411,N_12897);
nor U21108 (N_21108,N_12622,N_17260);
nor U21109 (N_21109,N_15939,N_17274);
and U21110 (N_21110,N_14647,N_13327);
or U21111 (N_21111,N_15991,N_15020);
xor U21112 (N_21112,N_13381,N_17535);
nand U21113 (N_21113,N_13565,N_15575);
and U21114 (N_21114,N_15762,N_16095);
or U21115 (N_21115,N_13071,N_13288);
nor U21116 (N_21116,N_14556,N_12869);
nand U21117 (N_21117,N_14223,N_12031);
nor U21118 (N_21118,N_13326,N_12739);
or U21119 (N_21119,N_14284,N_12193);
and U21120 (N_21120,N_16511,N_12796);
or U21121 (N_21121,N_12135,N_16851);
xor U21122 (N_21122,N_14992,N_13516);
or U21123 (N_21123,N_16335,N_16768);
or U21124 (N_21124,N_17528,N_13741);
and U21125 (N_21125,N_12609,N_16599);
xnor U21126 (N_21126,N_12734,N_17285);
and U21127 (N_21127,N_16517,N_12174);
nor U21128 (N_21128,N_15370,N_12414);
and U21129 (N_21129,N_16129,N_16114);
nor U21130 (N_21130,N_14277,N_14600);
and U21131 (N_21131,N_15797,N_16436);
nand U21132 (N_21132,N_14908,N_15425);
or U21133 (N_21133,N_12404,N_13305);
and U21134 (N_21134,N_12671,N_13093);
nor U21135 (N_21135,N_14025,N_12716);
nand U21136 (N_21136,N_15635,N_17122);
nor U21137 (N_21137,N_12747,N_13921);
or U21138 (N_21138,N_13379,N_13089);
nand U21139 (N_21139,N_15312,N_13919);
xor U21140 (N_21140,N_12029,N_12812);
nand U21141 (N_21141,N_17897,N_15759);
nand U21142 (N_21142,N_16834,N_15127);
and U21143 (N_21143,N_15825,N_16297);
xnor U21144 (N_21144,N_17046,N_13175);
nor U21145 (N_21145,N_13578,N_12614);
or U21146 (N_21146,N_16577,N_14524);
or U21147 (N_21147,N_16398,N_17247);
nand U21148 (N_21148,N_17851,N_14724);
nor U21149 (N_21149,N_14100,N_15753);
nor U21150 (N_21150,N_14518,N_12323);
or U21151 (N_21151,N_14312,N_12337);
nor U21152 (N_21152,N_13179,N_16530);
nor U21153 (N_21153,N_12802,N_13448);
or U21154 (N_21154,N_13397,N_15267);
nor U21155 (N_21155,N_14920,N_16294);
and U21156 (N_21156,N_17954,N_14980);
nor U21157 (N_21157,N_14451,N_13620);
or U21158 (N_21158,N_12534,N_16794);
nand U21159 (N_21159,N_15335,N_14430);
or U21160 (N_21160,N_15297,N_12789);
and U21161 (N_21161,N_15590,N_16286);
nor U21162 (N_21162,N_13093,N_17427);
xnor U21163 (N_21163,N_15542,N_14384);
nor U21164 (N_21164,N_17954,N_15479);
nor U21165 (N_21165,N_17082,N_15948);
and U21166 (N_21166,N_12193,N_16964);
nor U21167 (N_21167,N_15139,N_15798);
or U21168 (N_21168,N_13103,N_15253);
nand U21169 (N_21169,N_17871,N_13646);
nor U21170 (N_21170,N_14887,N_16956);
nor U21171 (N_21171,N_16573,N_13052);
or U21172 (N_21172,N_12778,N_17365);
nor U21173 (N_21173,N_16557,N_13611);
and U21174 (N_21174,N_12750,N_14077);
xor U21175 (N_21175,N_14491,N_12886);
xor U21176 (N_21176,N_17959,N_12575);
xnor U21177 (N_21177,N_17030,N_17458);
xnor U21178 (N_21178,N_17110,N_14537);
nand U21179 (N_21179,N_15845,N_13847);
nor U21180 (N_21180,N_17662,N_12195);
or U21181 (N_21181,N_13208,N_12562);
and U21182 (N_21182,N_16968,N_13028);
nand U21183 (N_21183,N_14889,N_13207);
or U21184 (N_21184,N_13061,N_13720);
nor U21185 (N_21185,N_15955,N_17766);
nor U21186 (N_21186,N_16466,N_17837);
xnor U21187 (N_21187,N_13022,N_16260);
nand U21188 (N_21188,N_15441,N_15018);
nor U21189 (N_21189,N_13351,N_12990);
or U21190 (N_21190,N_12987,N_12490);
nand U21191 (N_21191,N_16539,N_12801);
or U21192 (N_21192,N_13069,N_12402);
or U21193 (N_21193,N_12063,N_17115);
nor U21194 (N_21194,N_17225,N_16434);
nand U21195 (N_21195,N_17546,N_17049);
or U21196 (N_21196,N_13590,N_16894);
and U21197 (N_21197,N_13798,N_12668);
and U21198 (N_21198,N_13070,N_15020);
and U21199 (N_21199,N_17366,N_14874);
nand U21200 (N_21200,N_13860,N_17480);
xnor U21201 (N_21201,N_16344,N_13708);
nand U21202 (N_21202,N_16864,N_15032);
nor U21203 (N_21203,N_17290,N_12705);
or U21204 (N_21204,N_15739,N_12406);
or U21205 (N_21205,N_16076,N_17830);
nor U21206 (N_21206,N_16300,N_14372);
or U21207 (N_21207,N_17213,N_17084);
nand U21208 (N_21208,N_17023,N_13380);
and U21209 (N_21209,N_14348,N_13431);
nor U21210 (N_21210,N_17195,N_17247);
and U21211 (N_21211,N_16936,N_12978);
and U21212 (N_21212,N_14350,N_16262);
and U21213 (N_21213,N_12466,N_13142);
or U21214 (N_21214,N_15155,N_17512);
and U21215 (N_21215,N_13500,N_14845);
nand U21216 (N_21216,N_17539,N_12109);
xor U21217 (N_21217,N_13866,N_13587);
or U21218 (N_21218,N_12241,N_13363);
nand U21219 (N_21219,N_16125,N_12052);
nor U21220 (N_21220,N_17545,N_14224);
nand U21221 (N_21221,N_13617,N_14275);
nand U21222 (N_21222,N_16185,N_13946);
nand U21223 (N_21223,N_14877,N_16033);
and U21224 (N_21224,N_16964,N_15416);
nor U21225 (N_21225,N_15762,N_17062);
or U21226 (N_21226,N_14298,N_12882);
or U21227 (N_21227,N_14702,N_13763);
or U21228 (N_21228,N_17806,N_16980);
and U21229 (N_21229,N_13574,N_14827);
nand U21230 (N_21230,N_14404,N_17619);
nand U21231 (N_21231,N_17031,N_17697);
xnor U21232 (N_21232,N_17361,N_17772);
nand U21233 (N_21233,N_15425,N_14139);
nor U21234 (N_21234,N_16402,N_14488);
or U21235 (N_21235,N_12467,N_12236);
nor U21236 (N_21236,N_14955,N_15877);
and U21237 (N_21237,N_16319,N_12235);
nand U21238 (N_21238,N_16517,N_12077);
and U21239 (N_21239,N_14652,N_15141);
and U21240 (N_21240,N_13801,N_17755);
or U21241 (N_21241,N_12774,N_17610);
or U21242 (N_21242,N_12936,N_14371);
and U21243 (N_21243,N_17224,N_12465);
nand U21244 (N_21244,N_12559,N_12804);
nand U21245 (N_21245,N_16968,N_17747);
xnor U21246 (N_21246,N_14085,N_14799);
or U21247 (N_21247,N_14093,N_15119);
nand U21248 (N_21248,N_13265,N_15505);
nor U21249 (N_21249,N_15512,N_16342);
nand U21250 (N_21250,N_13549,N_15308);
and U21251 (N_21251,N_14246,N_15423);
and U21252 (N_21252,N_15605,N_15435);
nand U21253 (N_21253,N_13684,N_16847);
nand U21254 (N_21254,N_17160,N_15134);
nor U21255 (N_21255,N_12413,N_15643);
or U21256 (N_21256,N_13027,N_16023);
and U21257 (N_21257,N_13506,N_16224);
nor U21258 (N_21258,N_15545,N_15153);
nand U21259 (N_21259,N_13141,N_14058);
or U21260 (N_21260,N_16545,N_13405);
nand U21261 (N_21261,N_12968,N_13940);
nand U21262 (N_21262,N_17215,N_14884);
and U21263 (N_21263,N_14174,N_15467);
or U21264 (N_21264,N_12798,N_16832);
nand U21265 (N_21265,N_12231,N_13102);
nand U21266 (N_21266,N_16017,N_14231);
or U21267 (N_21267,N_14436,N_15482);
nor U21268 (N_21268,N_17500,N_16341);
and U21269 (N_21269,N_14693,N_15075);
or U21270 (N_21270,N_13111,N_13429);
and U21271 (N_21271,N_16334,N_17374);
nor U21272 (N_21272,N_12482,N_17818);
xor U21273 (N_21273,N_12169,N_14620);
xnor U21274 (N_21274,N_14472,N_15531);
nor U21275 (N_21275,N_15926,N_15594);
and U21276 (N_21276,N_16607,N_17440);
or U21277 (N_21277,N_14360,N_15015);
and U21278 (N_21278,N_17862,N_13105);
and U21279 (N_21279,N_16529,N_12050);
xnor U21280 (N_21280,N_16990,N_13633);
and U21281 (N_21281,N_17010,N_14885);
and U21282 (N_21282,N_16253,N_16789);
nor U21283 (N_21283,N_16383,N_16964);
xor U21284 (N_21284,N_17615,N_12903);
nand U21285 (N_21285,N_15558,N_15318);
or U21286 (N_21286,N_16393,N_12420);
nor U21287 (N_21287,N_12854,N_15401);
or U21288 (N_21288,N_13270,N_14860);
nor U21289 (N_21289,N_14338,N_12203);
or U21290 (N_21290,N_12714,N_15482);
and U21291 (N_21291,N_17662,N_15248);
xnor U21292 (N_21292,N_17681,N_16566);
nand U21293 (N_21293,N_12521,N_17470);
nand U21294 (N_21294,N_16648,N_16307);
nand U21295 (N_21295,N_13216,N_17213);
or U21296 (N_21296,N_13208,N_15556);
xnor U21297 (N_21297,N_15936,N_13048);
nor U21298 (N_21298,N_14674,N_12628);
or U21299 (N_21299,N_14728,N_15705);
nand U21300 (N_21300,N_17298,N_17532);
nand U21301 (N_21301,N_17178,N_17670);
or U21302 (N_21302,N_16703,N_12385);
nand U21303 (N_21303,N_12098,N_17930);
or U21304 (N_21304,N_17694,N_13253);
xor U21305 (N_21305,N_14043,N_16615);
and U21306 (N_21306,N_15170,N_16651);
nand U21307 (N_21307,N_14708,N_12398);
nand U21308 (N_21308,N_16533,N_17616);
nand U21309 (N_21309,N_14959,N_12521);
xor U21310 (N_21310,N_17348,N_17301);
and U21311 (N_21311,N_14776,N_14989);
xor U21312 (N_21312,N_16169,N_16268);
and U21313 (N_21313,N_15374,N_17672);
and U21314 (N_21314,N_14187,N_12042);
nor U21315 (N_21315,N_13410,N_12339);
or U21316 (N_21316,N_13700,N_16251);
xnor U21317 (N_21317,N_15775,N_13204);
nand U21318 (N_21318,N_14736,N_17885);
nand U21319 (N_21319,N_14727,N_17998);
and U21320 (N_21320,N_17776,N_15235);
nor U21321 (N_21321,N_17222,N_12908);
and U21322 (N_21322,N_16688,N_16672);
nor U21323 (N_21323,N_15477,N_16060);
and U21324 (N_21324,N_14049,N_15552);
nor U21325 (N_21325,N_16529,N_16611);
or U21326 (N_21326,N_14531,N_14997);
and U21327 (N_21327,N_13865,N_12108);
or U21328 (N_21328,N_12758,N_12465);
or U21329 (N_21329,N_12432,N_13105);
and U21330 (N_21330,N_17008,N_17713);
or U21331 (N_21331,N_14547,N_16301);
and U21332 (N_21332,N_13139,N_15198);
nand U21333 (N_21333,N_13859,N_15678);
and U21334 (N_21334,N_16417,N_12254);
or U21335 (N_21335,N_17761,N_12293);
nor U21336 (N_21336,N_12367,N_13213);
nor U21337 (N_21337,N_16654,N_15463);
xnor U21338 (N_21338,N_13611,N_12829);
or U21339 (N_21339,N_12393,N_17384);
or U21340 (N_21340,N_12467,N_16640);
nor U21341 (N_21341,N_13746,N_12869);
nor U21342 (N_21342,N_14456,N_12178);
nand U21343 (N_21343,N_13396,N_15227);
nor U21344 (N_21344,N_17060,N_13352);
xor U21345 (N_21345,N_14496,N_14706);
nor U21346 (N_21346,N_16358,N_13015);
and U21347 (N_21347,N_13323,N_14255);
and U21348 (N_21348,N_17815,N_12415);
and U21349 (N_21349,N_17043,N_12367);
and U21350 (N_21350,N_12225,N_15079);
and U21351 (N_21351,N_12470,N_13033);
nor U21352 (N_21352,N_12024,N_17885);
and U21353 (N_21353,N_14611,N_17764);
and U21354 (N_21354,N_14013,N_17711);
nand U21355 (N_21355,N_15736,N_12233);
nor U21356 (N_21356,N_12976,N_16688);
xor U21357 (N_21357,N_14519,N_17643);
or U21358 (N_21358,N_14938,N_13952);
and U21359 (N_21359,N_14292,N_17264);
and U21360 (N_21360,N_16936,N_14583);
xnor U21361 (N_21361,N_15703,N_12820);
nand U21362 (N_21362,N_13978,N_17530);
and U21363 (N_21363,N_16600,N_12419);
or U21364 (N_21364,N_17784,N_14342);
and U21365 (N_21365,N_15584,N_13001);
nand U21366 (N_21366,N_17571,N_17603);
and U21367 (N_21367,N_12034,N_16390);
nand U21368 (N_21368,N_15472,N_12668);
nor U21369 (N_21369,N_12403,N_17499);
xnor U21370 (N_21370,N_15080,N_13844);
nand U21371 (N_21371,N_13902,N_12116);
and U21372 (N_21372,N_14646,N_12959);
or U21373 (N_21373,N_15707,N_14145);
and U21374 (N_21374,N_15387,N_15560);
and U21375 (N_21375,N_17839,N_14104);
and U21376 (N_21376,N_16495,N_17329);
or U21377 (N_21377,N_13767,N_12205);
and U21378 (N_21378,N_14764,N_15209);
nand U21379 (N_21379,N_13232,N_15188);
and U21380 (N_21380,N_15402,N_13266);
nand U21381 (N_21381,N_12663,N_13768);
or U21382 (N_21382,N_12275,N_15599);
xor U21383 (N_21383,N_17004,N_12823);
nor U21384 (N_21384,N_15565,N_17718);
or U21385 (N_21385,N_17183,N_16464);
nor U21386 (N_21386,N_14693,N_14113);
nor U21387 (N_21387,N_15650,N_17433);
nand U21388 (N_21388,N_13507,N_17949);
or U21389 (N_21389,N_13391,N_14470);
or U21390 (N_21390,N_16610,N_14940);
or U21391 (N_21391,N_14173,N_15401);
nor U21392 (N_21392,N_15653,N_14056);
nand U21393 (N_21393,N_16292,N_13262);
nor U21394 (N_21394,N_16412,N_15413);
or U21395 (N_21395,N_12102,N_12399);
nand U21396 (N_21396,N_14676,N_12052);
and U21397 (N_21397,N_12670,N_14883);
nor U21398 (N_21398,N_14680,N_13308);
nand U21399 (N_21399,N_17273,N_12789);
or U21400 (N_21400,N_15480,N_16409);
nor U21401 (N_21401,N_12660,N_15394);
nor U21402 (N_21402,N_17965,N_15385);
nand U21403 (N_21403,N_12400,N_16200);
nor U21404 (N_21404,N_12075,N_15006);
and U21405 (N_21405,N_13084,N_14555);
nand U21406 (N_21406,N_14961,N_17443);
or U21407 (N_21407,N_15415,N_12586);
nand U21408 (N_21408,N_13093,N_14855);
or U21409 (N_21409,N_17044,N_17346);
and U21410 (N_21410,N_14080,N_12682);
or U21411 (N_21411,N_17261,N_12322);
nor U21412 (N_21412,N_12447,N_16037);
or U21413 (N_21413,N_15363,N_13308);
nand U21414 (N_21414,N_12175,N_17931);
and U21415 (N_21415,N_16844,N_17668);
and U21416 (N_21416,N_17797,N_17924);
nor U21417 (N_21417,N_13508,N_16730);
and U21418 (N_21418,N_12164,N_15704);
xor U21419 (N_21419,N_13589,N_14149);
nor U21420 (N_21420,N_14355,N_15669);
or U21421 (N_21421,N_17653,N_14495);
and U21422 (N_21422,N_14952,N_13077);
nand U21423 (N_21423,N_17756,N_13400);
nand U21424 (N_21424,N_14381,N_13403);
and U21425 (N_21425,N_12394,N_12598);
nand U21426 (N_21426,N_17644,N_17647);
nand U21427 (N_21427,N_16854,N_13498);
and U21428 (N_21428,N_12330,N_13270);
nor U21429 (N_21429,N_17669,N_13429);
and U21430 (N_21430,N_16806,N_14576);
nor U21431 (N_21431,N_16079,N_16168);
nand U21432 (N_21432,N_17943,N_13491);
nand U21433 (N_21433,N_12317,N_14134);
nor U21434 (N_21434,N_13364,N_12642);
or U21435 (N_21435,N_12770,N_12411);
or U21436 (N_21436,N_12952,N_16670);
and U21437 (N_21437,N_12109,N_15698);
nor U21438 (N_21438,N_15449,N_12023);
and U21439 (N_21439,N_16332,N_16231);
xnor U21440 (N_21440,N_14546,N_17988);
and U21441 (N_21441,N_17578,N_15262);
nor U21442 (N_21442,N_13254,N_17701);
or U21443 (N_21443,N_15015,N_16038);
xnor U21444 (N_21444,N_17238,N_12244);
nor U21445 (N_21445,N_13653,N_17313);
nor U21446 (N_21446,N_15490,N_17185);
or U21447 (N_21447,N_12049,N_16301);
nand U21448 (N_21448,N_14328,N_15972);
nor U21449 (N_21449,N_13419,N_12321);
and U21450 (N_21450,N_13383,N_12069);
nand U21451 (N_21451,N_16352,N_15808);
nand U21452 (N_21452,N_17952,N_14260);
or U21453 (N_21453,N_17095,N_13291);
nor U21454 (N_21454,N_14212,N_16932);
nor U21455 (N_21455,N_15966,N_16404);
nor U21456 (N_21456,N_15247,N_14934);
and U21457 (N_21457,N_14300,N_12475);
nand U21458 (N_21458,N_15477,N_14629);
nand U21459 (N_21459,N_16394,N_15779);
xor U21460 (N_21460,N_14172,N_17486);
and U21461 (N_21461,N_16207,N_12648);
nor U21462 (N_21462,N_17954,N_16200);
nor U21463 (N_21463,N_12778,N_17102);
nand U21464 (N_21464,N_16701,N_12339);
or U21465 (N_21465,N_13991,N_13601);
and U21466 (N_21466,N_16721,N_15490);
nand U21467 (N_21467,N_15590,N_14284);
nand U21468 (N_21468,N_16262,N_17769);
nand U21469 (N_21469,N_15929,N_15928);
nor U21470 (N_21470,N_15073,N_17989);
nand U21471 (N_21471,N_16767,N_13581);
or U21472 (N_21472,N_13517,N_12959);
nor U21473 (N_21473,N_14625,N_15879);
or U21474 (N_21474,N_17857,N_13476);
nand U21475 (N_21475,N_12260,N_16654);
xor U21476 (N_21476,N_14291,N_12416);
nor U21477 (N_21477,N_16669,N_17508);
or U21478 (N_21478,N_15423,N_16820);
nor U21479 (N_21479,N_14385,N_15250);
nand U21480 (N_21480,N_16524,N_16512);
nand U21481 (N_21481,N_14628,N_14579);
and U21482 (N_21482,N_16903,N_13672);
xor U21483 (N_21483,N_14424,N_17245);
or U21484 (N_21484,N_14108,N_15364);
nor U21485 (N_21485,N_16705,N_12973);
and U21486 (N_21486,N_17402,N_14931);
and U21487 (N_21487,N_15408,N_15601);
xnor U21488 (N_21488,N_14893,N_16067);
and U21489 (N_21489,N_14452,N_12157);
nand U21490 (N_21490,N_16767,N_15684);
nand U21491 (N_21491,N_14912,N_12949);
or U21492 (N_21492,N_14904,N_17435);
nand U21493 (N_21493,N_17715,N_14116);
nor U21494 (N_21494,N_15061,N_15676);
nand U21495 (N_21495,N_17630,N_12649);
and U21496 (N_21496,N_16664,N_15119);
or U21497 (N_21497,N_14330,N_15749);
nand U21498 (N_21498,N_15651,N_15705);
and U21499 (N_21499,N_15450,N_17314);
and U21500 (N_21500,N_17641,N_17944);
or U21501 (N_21501,N_13635,N_17486);
and U21502 (N_21502,N_16211,N_17009);
nand U21503 (N_21503,N_14477,N_14969);
nand U21504 (N_21504,N_14141,N_15342);
nand U21505 (N_21505,N_16217,N_12215);
xnor U21506 (N_21506,N_15823,N_17270);
xnor U21507 (N_21507,N_12142,N_13699);
nand U21508 (N_21508,N_16141,N_15713);
nor U21509 (N_21509,N_13702,N_16712);
nor U21510 (N_21510,N_16311,N_14569);
xor U21511 (N_21511,N_16402,N_13713);
nor U21512 (N_21512,N_14358,N_16904);
nand U21513 (N_21513,N_16394,N_15150);
nand U21514 (N_21514,N_14066,N_16356);
nand U21515 (N_21515,N_15831,N_12249);
nor U21516 (N_21516,N_16026,N_12995);
nand U21517 (N_21517,N_15159,N_16585);
or U21518 (N_21518,N_15107,N_17765);
or U21519 (N_21519,N_13185,N_14469);
and U21520 (N_21520,N_13304,N_14387);
nor U21521 (N_21521,N_12948,N_15930);
or U21522 (N_21522,N_13353,N_14837);
and U21523 (N_21523,N_15410,N_16612);
xor U21524 (N_21524,N_16508,N_16445);
and U21525 (N_21525,N_15155,N_16249);
nand U21526 (N_21526,N_12758,N_13341);
xor U21527 (N_21527,N_16399,N_16579);
nor U21528 (N_21528,N_12579,N_12975);
nor U21529 (N_21529,N_16351,N_15148);
nand U21530 (N_21530,N_13461,N_14478);
and U21531 (N_21531,N_13576,N_16697);
nand U21532 (N_21532,N_12474,N_16723);
and U21533 (N_21533,N_16914,N_13429);
and U21534 (N_21534,N_16703,N_12929);
or U21535 (N_21535,N_13250,N_17193);
and U21536 (N_21536,N_12567,N_12989);
xor U21537 (N_21537,N_15224,N_12923);
nand U21538 (N_21538,N_14855,N_12742);
and U21539 (N_21539,N_13729,N_12926);
nor U21540 (N_21540,N_12437,N_17549);
xor U21541 (N_21541,N_12756,N_12154);
nand U21542 (N_21542,N_14213,N_16902);
nor U21543 (N_21543,N_12133,N_16936);
and U21544 (N_21544,N_17726,N_14504);
nor U21545 (N_21545,N_16797,N_14653);
nand U21546 (N_21546,N_17657,N_17512);
xnor U21547 (N_21547,N_17625,N_15640);
and U21548 (N_21548,N_13774,N_13787);
nor U21549 (N_21549,N_15965,N_13482);
nand U21550 (N_21550,N_15362,N_16463);
or U21551 (N_21551,N_16968,N_16992);
nor U21552 (N_21552,N_14093,N_12839);
or U21553 (N_21553,N_17685,N_15207);
nor U21554 (N_21554,N_12032,N_15944);
nor U21555 (N_21555,N_17934,N_13422);
nand U21556 (N_21556,N_16302,N_12365);
nor U21557 (N_21557,N_17635,N_16917);
nor U21558 (N_21558,N_14081,N_13883);
nand U21559 (N_21559,N_14803,N_17827);
nand U21560 (N_21560,N_14798,N_13665);
or U21561 (N_21561,N_16162,N_15299);
and U21562 (N_21562,N_15887,N_13275);
nor U21563 (N_21563,N_13416,N_15532);
and U21564 (N_21564,N_17892,N_16733);
nor U21565 (N_21565,N_12285,N_17640);
nor U21566 (N_21566,N_14656,N_15139);
and U21567 (N_21567,N_13498,N_14294);
nand U21568 (N_21568,N_16320,N_14942);
and U21569 (N_21569,N_15368,N_14196);
nor U21570 (N_21570,N_15280,N_16380);
nand U21571 (N_21571,N_12505,N_17485);
and U21572 (N_21572,N_14307,N_17060);
or U21573 (N_21573,N_13980,N_17582);
nand U21574 (N_21574,N_13150,N_13821);
and U21575 (N_21575,N_13660,N_16082);
nand U21576 (N_21576,N_12377,N_16852);
nor U21577 (N_21577,N_13278,N_13536);
nand U21578 (N_21578,N_13050,N_14631);
nor U21579 (N_21579,N_12910,N_15842);
nor U21580 (N_21580,N_17055,N_16029);
nor U21581 (N_21581,N_17072,N_14651);
nor U21582 (N_21582,N_15752,N_17980);
nor U21583 (N_21583,N_12708,N_12354);
nor U21584 (N_21584,N_12934,N_17447);
or U21585 (N_21585,N_14928,N_17608);
nor U21586 (N_21586,N_13415,N_14930);
or U21587 (N_21587,N_15200,N_17258);
nor U21588 (N_21588,N_13121,N_16028);
xnor U21589 (N_21589,N_16555,N_17165);
and U21590 (N_21590,N_12351,N_12718);
and U21591 (N_21591,N_14677,N_16822);
nor U21592 (N_21592,N_12853,N_17367);
nor U21593 (N_21593,N_12018,N_17319);
and U21594 (N_21594,N_12638,N_14386);
xnor U21595 (N_21595,N_14756,N_14761);
or U21596 (N_21596,N_14060,N_16640);
or U21597 (N_21597,N_12708,N_17608);
and U21598 (N_21598,N_13858,N_12120);
nor U21599 (N_21599,N_15217,N_15210);
nand U21600 (N_21600,N_15187,N_12987);
nor U21601 (N_21601,N_16421,N_17875);
and U21602 (N_21602,N_15663,N_14632);
nor U21603 (N_21603,N_13611,N_13647);
and U21604 (N_21604,N_16535,N_16837);
and U21605 (N_21605,N_15415,N_14513);
or U21606 (N_21606,N_12191,N_16434);
or U21607 (N_21607,N_16222,N_17240);
xor U21608 (N_21608,N_14111,N_13006);
nor U21609 (N_21609,N_12142,N_13891);
nand U21610 (N_21610,N_13525,N_13844);
nor U21611 (N_21611,N_16689,N_17662);
and U21612 (N_21612,N_16897,N_13642);
nand U21613 (N_21613,N_13155,N_17230);
nor U21614 (N_21614,N_17218,N_17207);
xor U21615 (N_21615,N_15694,N_15778);
or U21616 (N_21616,N_12353,N_17896);
nor U21617 (N_21617,N_17002,N_12588);
nor U21618 (N_21618,N_16640,N_12194);
or U21619 (N_21619,N_16107,N_14684);
or U21620 (N_21620,N_17459,N_17265);
and U21621 (N_21621,N_12187,N_13228);
or U21622 (N_21622,N_16187,N_14101);
nand U21623 (N_21623,N_13527,N_13352);
nor U21624 (N_21624,N_17016,N_17707);
and U21625 (N_21625,N_15949,N_16367);
and U21626 (N_21626,N_17837,N_13767);
nor U21627 (N_21627,N_12319,N_15491);
xnor U21628 (N_21628,N_15716,N_15484);
or U21629 (N_21629,N_15041,N_14914);
nor U21630 (N_21630,N_14732,N_15825);
xnor U21631 (N_21631,N_12153,N_17598);
nor U21632 (N_21632,N_15426,N_16566);
and U21633 (N_21633,N_14918,N_15332);
nor U21634 (N_21634,N_13652,N_13975);
and U21635 (N_21635,N_14595,N_15320);
and U21636 (N_21636,N_17656,N_17655);
nor U21637 (N_21637,N_12711,N_14089);
nor U21638 (N_21638,N_16166,N_13618);
or U21639 (N_21639,N_15796,N_12839);
or U21640 (N_21640,N_16168,N_13949);
and U21641 (N_21641,N_17909,N_12719);
nand U21642 (N_21642,N_14370,N_12746);
nor U21643 (N_21643,N_14025,N_16991);
and U21644 (N_21644,N_17889,N_13112);
nand U21645 (N_21645,N_14239,N_14699);
nand U21646 (N_21646,N_17650,N_14772);
nor U21647 (N_21647,N_13589,N_17110);
or U21648 (N_21648,N_15919,N_16162);
and U21649 (N_21649,N_12018,N_17784);
nand U21650 (N_21650,N_15559,N_13475);
nand U21651 (N_21651,N_17852,N_13715);
xor U21652 (N_21652,N_13219,N_14425);
or U21653 (N_21653,N_15343,N_13972);
nand U21654 (N_21654,N_16066,N_14759);
and U21655 (N_21655,N_12730,N_17149);
and U21656 (N_21656,N_14627,N_17535);
and U21657 (N_21657,N_13786,N_16385);
or U21658 (N_21658,N_12616,N_15749);
or U21659 (N_21659,N_12977,N_17157);
xor U21660 (N_21660,N_16746,N_16650);
and U21661 (N_21661,N_12775,N_12472);
nand U21662 (N_21662,N_17221,N_16684);
nor U21663 (N_21663,N_12156,N_14181);
nand U21664 (N_21664,N_15042,N_15838);
nor U21665 (N_21665,N_12741,N_16197);
or U21666 (N_21666,N_15395,N_13721);
or U21667 (N_21667,N_17447,N_15936);
nor U21668 (N_21668,N_13747,N_13378);
nand U21669 (N_21669,N_17427,N_15536);
xnor U21670 (N_21670,N_12062,N_15737);
nor U21671 (N_21671,N_14853,N_15105);
nand U21672 (N_21672,N_15365,N_13962);
and U21673 (N_21673,N_12025,N_15637);
and U21674 (N_21674,N_13998,N_12258);
nand U21675 (N_21675,N_14715,N_13403);
xor U21676 (N_21676,N_12765,N_17894);
and U21677 (N_21677,N_12649,N_17575);
nor U21678 (N_21678,N_14459,N_17828);
and U21679 (N_21679,N_15122,N_15493);
or U21680 (N_21680,N_17529,N_13767);
xor U21681 (N_21681,N_13760,N_13432);
or U21682 (N_21682,N_13222,N_15608);
and U21683 (N_21683,N_17013,N_15051);
nor U21684 (N_21684,N_14405,N_12975);
and U21685 (N_21685,N_17383,N_12807);
nand U21686 (N_21686,N_13428,N_14538);
nand U21687 (N_21687,N_13729,N_17553);
and U21688 (N_21688,N_14979,N_13507);
and U21689 (N_21689,N_14887,N_14397);
nor U21690 (N_21690,N_14141,N_12740);
and U21691 (N_21691,N_17276,N_17828);
and U21692 (N_21692,N_16489,N_15332);
or U21693 (N_21693,N_16189,N_12521);
xor U21694 (N_21694,N_16737,N_17532);
or U21695 (N_21695,N_17359,N_14453);
or U21696 (N_21696,N_15393,N_17370);
and U21697 (N_21697,N_15437,N_14163);
nor U21698 (N_21698,N_17266,N_16783);
nand U21699 (N_21699,N_12809,N_15944);
nor U21700 (N_21700,N_13476,N_12700);
nand U21701 (N_21701,N_17550,N_12457);
and U21702 (N_21702,N_15176,N_15220);
nor U21703 (N_21703,N_15240,N_13990);
nor U21704 (N_21704,N_17293,N_17790);
and U21705 (N_21705,N_14141,N_15860);
nand U21706 (N_21706,N_15591,N_13100);
and U21707 (N_21707,N_13723,N_16436);
nand U21708 (N_21708,N_13026,N_17700);
nand U21709 (N_21709,N_13770,N_13288);
xor U21710 (N_21710,N_12554,N_16805);
nand U21711 (N_21711,N_12074,N_17744);
nor U21712 (N_21712,N_16336,N_15196);
nand U21713 (N_21713,N_13942,N_16065);
xnor U21714 (N_21714,N_12420,N_16409);
or U21715 (N_21715,N_15532,N_16826);
nand U21716 (N_21716,N_15842,N_17391);
nand U21717 (N_21717,N_13159,N_14555);
or U21718 (N_21718,N_12086,N_13817);
xnor U21719 (N_21719,N_12595,N_12743);
and U21720 (N_21720,N_14564,N_13955);
or U21721 (N_21721,N_16274,N_13004);
or U21722 (N_21722,N_16186,N_14105);
and U21723 (N_21723,N_13465,N_13951);
and U21724 (N_21724,N_16699,N_15498);
nor U21725 (N_21725,N_17273,N_13002);
nor U21726 (N_21726,N_12951,N_14328);
xor U21727 (N_21727,N_12537,N_14056);
or U21728 (N_21728,N_13819,N_15669);
nand U21729 (N_21729,N_14723,N_14300);
nor U21730 (N_21730,N_12915,N_12418);
nand U21731 (N_21731,N_13579,N_13448);
and U21732 (N_21732,N_17284,N_13742);
nand U21733 (N_21733,N_12603,N_15537);
or U21734 (N_21734,N_14052,N_15954);
nor U21735 (N_21735,N_12592,N_16828);
or U21736 (N_21736,N_16606,N_17959);
xnor U21737 (N_21737,N_16243,N_16221);
nand U21738 (N_21738,N_14564,N_17750);
or U21739 (N_21739,N_15831,N_16558);
nor U21740 (N_21740,N_13207,N_16200);
and U21741 (N_21741,N_12954,N_15862);
and U21742 (N_21742,N_17191,N_14834);
nand U21743 (N_21743,N_17645,N_17592);
and U21744 (N_21744,N_13665,N_13980);
or U21745 (N_21745,N_13060,N_17005);
nand U21746 (N_21746,N_17020,N_17323);
nor U21747 (N_21747,N_16263,N_16265);
or U21748 (N_21748,N_12864,N_13080);
nor U21749 (N_21749,N_17045,N_16715);
nand U21750 (N_21750,N_12181,N_14511);
nand U21751 (N_21751,N_17550,N_13214);
or U21752 (N_21752,N_12581,N_15820);
nand U21753 (N_21753,N_14517,N_13175);
and U21754 (N_21754,N_16398,N_12936);
xor U21755 (N_21755,N_17497,N_13069);
and U21756 (N_21756,N_14280,N_13091);
and U21757 (N_21757,N_15765,N_16781);
and U21758 (N_21758,N_14356,N_15936);
and U21759 (N_21759,N_12629,N_12719);
nor U21760 (N_21760,N_15133,N_14981);
and U21761 (N_21761,N_17803,N_16222);
and U21762 (N_21762,N_13576,N_14080);
nand U21763 (N_21763,N_12202,N_15911);
and U21764 (N_21764,N_14061,N_14617);
nor U21765 (N_21765,N_15347,N_15833);
nor U21766 (N_21766,N_12933,N_13303);
nor U21767 (N_21767,N_16162,N_16223);
xor U21768 (N_21768,N_17251,N_16958);
nor U21769 (N_21769,N_16971,N_12310);
and U21770 (N_21770,N_15414,N_15834);
nand U21771 (N_21771,N_13040,N_15202);
and U21772 (N_21772,N_12563,N_12987);
nor U21773 (N_21773,N_16918,N_14975);
nand U21774 (N_21774,N_17153,N_12820);
or U21775 (N_21775,N_17265,N_17009);
and U21776 (N_21776,N_12874,N_17683);
and U21777 (N_21777,N_14784,N_15570);
xor U21778 (N_21778,N_12650,N_16011);
nand U21779 (N_21779,N_12533,N_12547);
nor U21780 (N_21780,N_16977,N_13548);
nand U21781 (N_21781,N_12158,N_12820);
xnor U21782 (N_21782,N_13033,N_13221);
and U21783 (N_21783,N_17300,N_14702);
xor U21784 (N_21784,N_12909,N_15594);
nor U21785 (N_21785,N_16094,N_12817);
xnor U21786 (N_21786,N_13550,N_12915);
or U21787 (N_21787,N_17789,N_17124);
or U21788 (N_21788,N_15296,N_12412);
xor U21789 (N_21789,N_13362,N_13097);
xnor U21790 (N_21790,N_13597,N_16749);
nor U21791 (N_21791,N_12407,N_17162);
or U21792 (N_21792,N_16148,N_17085);
nor U21793 (N_21793,N_14442,N_15468);
and U21794 (N_21794,N_16813,N_16719);
nand U21795 (N_21795,N_14849,N_12835);
nand U21796 (N_21796,N_15540,N_14699);
and U21797 (N_21797,N_13476,N_15464);
and U21798 (N_21798,N_14809,N_17569);
and U21799 (N_21799,N_14047,N_17753);
nand U21800 (N_21800,N_14797,N_16934);
and U21801 (N_21801,N_12458,N_14884);
or U21802 (N_21802,N_17983,N_15817);
nor U21803 (N_21803,N_12423,N_16977);
xnor U21804 (N_21804,N_12645,N_15573);
nor U21805 (N_21805,N_14099,N_17758);
or U21806 (N_21806,N_16787,N_16074);
and U21807 (N_21807,N_13909,N_16463);
and U21808 (N_21808,N_16741,N_17791);
nor U21809 (N_21809,N_14761,N_13727);
or U21810 (N_21810,N_16928,N_17696);
nand U21811 (N_21811,N_17956,N_13579);
or U21812 (N_21812,N_17567,N_13795);
or U21813 (N_21813,N_14876,N_13188);
xor U21814 (N_21814,N_17184,N_14883);
and U21815 (N_21815,N_15763,N_13715);
or U21816 (N_21816,N_12674,N_13568);
or U21817 (N_21817,N_15267,N_13603);
or U21818 (N_21818,N_15040,N_13007);
and U21819 (N_21819,N_15171,N_13625);
nor U21820 (N_21820,N_15370,N_16294);
or U21821 (N_21821,N_15994,N_15175);
nand U21822 (N_21822,N_12269,N_17923);
and U21823 (N_21823,N_16686,N_15491);
and U21824 (N_21824,N_17685,N_17519);
nor U21825 (N_21825,N_17186,N_12742);
nor U21826 (N_21826,N_14743,N_13264);
or U21827 (N_21827,N_12368,N_17028);
xor U21828 (N_21828,N_12567,N_12196);
and U21829 (N_21829,N_17865,N_16369);
xor U21830 (N_21830,N_12226,N_15987);
or U21831 (N_21831,N_13747,N_12622);
nand U21832 (N_21832,N_14863,N_12560);
nor U21833 (N_21833,N_14793,N_13079);
and U21834 (N_21834,N_12505,N_15758);
nand U21835 (N_21835,N_12320,N_12038);
and U21836 (N_21836,N_16220,N_17871);
nand U21837 (N_21837,N_14274,N_13230);
nor U21838 (N_21838,N_13915,N_17617);
or U21839 (N_21839,N_13174,N_15667);
and U21840 (N_21840,N_14060,N_16563);
nor U21841 (N_21841,N_17471,N_16667);
nor U21842 (N_21842,N_14492,N_14537);
and U21843 (N_21843,N_17068,N_13597);
nand U21844 (N_21844,N_12841,N_16219);
and U21845 (N_21845,N_13155,N_12686);
or U21846 (N_21846,N_14122,N_12085);
or U21847 (N_21847,N_13410,N_14994);
xnor U21848 (N_21848,N_12622,N_15007);
nand U21849 (N_21849,N_12606,N_13377);
and U21850 (N_21850,N_13005,N_14737);
and U21851 (N_21851,N_14436,N_16793);
or U21852 (N_21852,N_14664,N_17143);
nand U21853 (N_21853,N_17136,N_17615);
nand U21854 (N_21854,N_15858,N_17155);
nor U21855 (N_21855,N_12695,N_14751);
or U21856 (N_21856,N_13420,N_12063);
nor U21857 (N_21857,N_13466,N_15473);
nand U21858 (N_21858,N_17382,N_14304);
or U21859 (N_21859,N_14521,N_14066);
xor U21860 (N_21860,N_14362,N_16894);
or U21861 (N_21861,N_15115,N_16656);
and U21862 (N_21862,N_13265,N_15185);
nand U21863 (N_21863,N_16418,N_12021);
nand U21864 (N_21864,N_16349,N_12338);
or U21865 (N_21865,N_13103,N_13448);
xnor U21866 (N_21866,N_16082,N_13118);
or U21867 (N_21867,N_14727,N_17170);
nand U21868 (N_21868,N_17830,N_12548);
xnor U21869 (N_21869,N_17593,N_16167);
and U21870 (N_21870,N_15386,N_13150);
or U21871 (N_21871,N_16219,N_15816);
or U21872 (N_21872,N_14029,N_12813);
nor U21873 (N_21873,N_16112,N_13620);
nor U21874 (N_21874,N_12733,N_14775);
nor U21875 (N_21875,N_15588,N_14846);
xnor U21876 (N_21876,N_17523,N_13336);
and U21877 (N_21877,N_16900,N_13850);
nand U21878 (N_21878,N_13782,N_14784);
nor U21879 (N_21879,N_15073,N_14237);
nor U21880 (N_21880,N_15869,N_17656);
xor U21881 (N_21881,N_15916,N_16916);
and U21882 (N_21882,N_17622,N_15640);
nand U21883 (N_21883,N_15117,N_17291);
or U21884 (N_21884,N_16894,N_13569);
nand U21885 (N_21885,N_17643,N_13665);
nand U21886 (N_21886,N_15415,N_17476);
nor U21887 (N_21887,N_12470,N_17038);
or U21888 (N_21888,N_17298,N_15969);
nand U21889 (N_21889,N_12379,N_14180);
xor U21890 (N_21890,N_15683,N_15325);
or U21891 (N_21891,N_14668,N_12591);
and U21892 (N_21892,N_16326,N_17359);
and U21893 (N_21893,N_15864,N_12697);
nor U21894 (N_21894,N_12917,N_13454);
or U21895 (N_21895,N_13492,N_14752);
or U21896 (N_21896,N_13117,N_16357);
or U21897 (N_21897,N_17192,N_16978);
or U21898 (N_21898,N_16114,N_13346);
nor U21899 (N_21899,N_13204,N_13643);
and U21900 (N_21900,N_13876,N_15740);
nand U21901 (N_21901,N_12200,N_12787);
or U21902 (N_21902,N_13430,N_14821);
and U21903 (N_21903,N_14103,N_16605);
and U21904 (N_21904,N_14547,N_16951);
nand U21905 (N_21905,N_12695,N_12592);
or U21906 (N_21906,N_17103,N_15999);
or U21907 (N_21907,N_15495,N_15187);
nor U21908 (N_21908,N_12643,N_13134);
nor U21909 (N_21909,N_14328,N_15440);
nor U21910 (N_21910,N_14073,N_15666);
xnor U21911 (N_21911,N_13173,N_14390);
nor U21912 (N_21912,N_13780,N_17111);
nand U21913 (N_21913,N_14976,N_12487);
and U21914 (N_21914,N_12266,N_14577);
or U21915 (N_21915,N_15462,N_16784);
and U21916 (N_21916,N_12072,N_15979);
xor U21917 (N_21917,N_17433,N_15933);
nor U21918 (N_21918,N_12618,N_16505);
nor U21919 (N_21919,N_14510,N_12698);
or U21920 (N_21920,N_17877,N_14925);
nor U21921 (N_21921,N_17573,N_16627);
nor U21922 (N_21922,N_14761,N_13457);
and U21923 (N_21923,N_12877,N_17940);
or U21924 (N_21924,N_14182,N_14541);
nor U21925 (N_21925,N_14645,N_13501);
nor U21926 (N_21926,N_14259,N_16544);
and U21927 (N_21927,N_17545,N_15624);
or U21928 (N_21928,N_16999,N_13958);
or U21929 (N_21929,N_14654,N_13722);
or U21930 (N_21930,N_16367,N_12634);
or U21931 (N_21931,N_15241,N_13775);
nor U21932 (N_21932,N_12109,N_13808);
or U21933 (N_21933,N_14946,N_13208);
nand U21934 (N_21934,N_12328,N_12842);
nand U21935 (N_21935,N_13316,N_15711);
nand U21936 (N_21936,N_16637,N_13036);
nand U21937 (N_21937,N_14376,N_12693);
and U21938 (N_21938,N_16651,N_14844);
and U21939 (N_21939,N_15709,N_16772);
or U21940 (N_21940,N_14409,N_14589);
xor U21941 (N_21941,N_14366,N_16265);
and U21942 (N_21942,N_14175,N_17363);
nor U21943 (N_21943,N_16496,N_12334);
nand U21944 (N_21944,N_15926,N_15680);
and U21945 (N_21945,N_16752,N_12920);
xor U21946 (N_21946,N_14125,N_16910);
and U21947 (N_21947,N_13990,N_12026);
or U21948 (N_21948,N_12288,N_15669);
or U21949 (N_21949,N_15489,N_12525);
and U21950 (N_21950,N_15632,N_16700);
or U21951 (N_21951,N_16608,N_17975);
nor U21952 (N_21952,N_15913,N_17493);
and U21953 (N_21953,N_14612,N_14037);
and U21954 (N_21954,N_12343,N_13951);
xor U21955 (N_21955,N_13926,N_16072);
nand U21956 (N_21956,N_14440,N_15713);
or U21957 (N_21957,N_13864,N_12901);
nand U21958 (N_21958,N_14590,N_16568);
nand U21959 (N_21959,N_17776,N_12824);
nor U21960 (N_21960,N_17872,N_17836);
xor U21961 (N_21961,N_17064,N_16153);
xor U21962 (N_21962,N_13482,N_13944);
or U21963 (N_21963,N_12761,N_15210);
or U21964 (N_21964,N_14136,N_14798);
nand U21965 (N_21965,N_13400,N_17437);
xnor U21966 (N_21966,N_15896,N_14726);
xnor U21967 (N_21967,N_15033,N_17512);
and U21968 (N_21968,N_13869,N_14558);
xor U21969 (N_21969,N_13288,N_17307);
nor U21970 (N_21970,N_17921,N_15420);
and U21971 (N_21971,N_12761,N_12993);
nand U21972 (N_21972,N_13025,N_16110);
or U21973 (N_21973,N_12136,N_14626);
xor U21974 (N_21974,N_14866,N_14126);
nand U21975 (N_21975,N_15244,N_12996);
or U21976 (N_21976,N_12936,N_13031);
or U21977 (N_21977,N_15668,N_16431);
nand U21978 (N_21978,N_12266,N_17635);
xnor U21979 (N_21979,N_16617,N_17514);
xor U21980 (N_21980,N_12872,N_13076);
or U21981 (N_21981,N_13553,N_17554);
and U21982 (N_21982,N_16255,N_16939);
nand U21983 (N_21983,N_14789,N_13164);
nor U21984 (N_21984,N_14502,N_17336);
or U21985 (N_21985,N_17336,N_15026);
and U21986 (N_21986,N_16935,N_14758);
nor U21987 (N_21987,N_12881,N_15309);
and U21988 (N_21988,N_15146,N_12486);
nor U21989 (N_21989,N_16170,N_12294);
nand U21990 (N_21990,N_15795,N_15110);
and U21991 (N_21991,N_12393,N_13260);
and U21992 (N_21992,N_13163,N_17074);
and U21993 (N_21993,N_14665,N_16658);
and U21994 (N_21994,N_12234,N_12834);
nand U21995 (N_21995,N_12499,N_13876);
and U21996 (N_21996,N_12996,N_16566);
and U21997 (N_21997,N_12645,N_13983);
nand U21998 (N_21998,N_12849,N_13541);
nand U21999 (N_21999,N_15267,N_15989);
nor U22000 (N_22000,N_17186,N_12695);
nor U22001 (N_22001,N_16998,N_16063);
nor U22002 (N_22002,N_15804,N_13344);
xor U22003 (N_22003,N_16878,N_15987);
nand U22004 (N_22004,N_13708,N_15838);
or U22005 (N_22005,N_14890,N_15759);
nand U22006 (N_22006,N_15793,N_16548);
and U22007 (N_22007,N_14370,N_14181);
or U22008 (N_22008,N_14061,N_17325);
and U22009 (N_22009,N_16705,N_17889);
or U22010 (N_22010,N_15263,N_13065);
nand U22011 (N_22011,N_15354,N_13664);
nor U22012 (N_22012,N_17163,N_16933);
and U22013 (N_22013,N_13091,N_16739);
and U22014 (N_22014,N_15231,N_12581);
or U22015 (N_22015,N_15967,N_16157);
nand U22016 (N_22016,N_15362,N_12041);
nand U22017 (N_22017,N_13910,N_15675);
or U22018 (N_22018,N_14680,N_16306);
nor U22019 (N_22019,N_16278,N_12643);
nand U22020 (N_22020,N_16815,N_12375);
and U22021 (N_22021,N_14955,N_12027);
nand U22022 (N_22022,N_12856,N_14633);
nand U22023 (N_22023,N_13810,N_13702);
nand U22024 (N_22024,N_14418,N_16700);
nand U22025 (N_22025,N_12909,N_13750);
nor U22026 (N_22026,N_12363,N_17810);
xnor U22027 (N_22027,N_12802,N_12512);
and U22028 (N_22028,N_13684,N_16199);
nand U22029 (N_22029,N_12353,N_17334);
nor U22030 (N_22030,N_16851,N_16352);
xor U22031 (N_22031,N_12913,N_14245);
and U22032 (N_22032,N_12470,N_14126);
nand U22033 (N_22033,N_14471,N_14053);
and U22034 (N_22034,N_13616,N_14079);
or U22035 (N_22035,N_17587,N_15523);
and U22036 (N_22036,N_13084,N_14896);
nand U22037 (N_22037,N_17410,N_12909);
or U22038 (N_22038,N_15073,N_16038);
and U22039 (N_22039,N_17043,N_12634);
xnor U22040 (N_22040,N_12294,N_17555);
nand U22041 (N_22041,N_15664,N_14027);
or U22042 (N_22042,N_14465,N_13736);
and U22043 (N_22043,N_16334,N_15621);
nand U22044 (N_22044,N_17403,N_12120);
nor U22045 (N_22045,N_14067,N_16308);
nor U22046 (N_22046,N_16716,N_13304);
nor U22047 (N_22047,N_15214,N_13872);
nor U22048 (N_22048,N_15983,N_14562);
or U22049 (N_22049,N_13150,N_15903);
nand U22050 (N_22050,N_12072,N_14611);
nor U22051 (N_22051,N_16955,N_17799);
or U22052 (N_22052,N_14583,N_17498);
or U22053 (N_22053,N_13171,N_15706);
and U22054 (N_22054,N_13660,N_16635);
and U22055 (N_22055,N_14777,N_13216);
nor U22056 (N_22056,N_17833,N_13176);
and U22057 (N_22057,N_14886,N_16521);
or U22058 (N_22058,N_15102,N_12404);
xnor U22059 (N_22059,N_14008,N_14180);
nor U22060 (N_22060,N_12993,N_12846);
xnor U22061 (N_22061,N_16772,N_15219);
or U22062 (N_22062,N_12234,N_15123);
nand U22063 (N_22063,N_17989,N_13636);
xnor U22064 (N_22064,N_15332,N_15164);
nand U22065 (N_22065,N_17750,N_12384);
nand U22066 (N_22066,N_14296,N_16514);
and U22067 (N_22067,N_14871,N_13323);
or U22068 (N_22068,N_12783,N_16439);
or U22069 (N_22069,N_12293,N_12848);
nand U22070 (N_22070,N_15444,N_14811);
nor U22071 (N_22071,N_15110,N_17482);
nor U22072 (N_22072,N_15217,N_15935);
and U22073 (N_22073,N_14053,N_17299);
nand U22074 (N_22074,N_17942,N_15585);
nor U22075 (N_22075,N_15053,N_16489);
and U22076 (N_22076,N_13192,N_12561);
xor U22077 (N_22077,N_14656,N_16791);
nand U22078 (N_22078,N_16117,N_17868);
and U22079 (N_22079,N_13172,N_13611);
or U22080 (N_22080,N_12471,N_12039);
nor U22081 (N_22081,N_15480,N_12575);
or U22082 (N_22082,N_13041,N_14422);
or U22083 (N_22083,N_17070,N_15302);
or U22084 (N_22084,N_16171,N_15477);
xnor U22085 (N_22085,N_16439,N_15919);
xor U22086 (N_22086,N_16121,N_12321);
nor U22087 (N_22087,N_15436,N_14423);
or U22088 (N_22088,N_13981,N_17596);
and U22089 (N_22089,N_13203,N_13953);
or U22090 (N_22090,N_12080,N_14942);
or U22091 (N_22091,N_17012,N_17488);
and U22092 (N_22092,N_12652,N_17236);
or U22093 (N_22093,N_13275,N_12368);
nand U22094 (N_22094,N_12515,N_15462);
xor U22095 (N_22095,N_16088,N_15663);
and U22096 (N_22096,N_12469,N_15461);
nor U22097 (N_22097,N_12845,N_16136);
xor U22098 (N_22098,N_14023,N_12466);
and U22099 (N_22099,N_14339,N_13678);
xor U22100 (N_22100,N_15881,N_16350);
nor U22101 (N_22101,N_16244,N_14619);
and U22102 (N_22102,N_15655,N_17156);
and U22103 (N_22103,N_15708,N_17558);
nor U22104 (N_22104,N_14162,N_15109);
and U22105 (N_22105,N_12142,N_12564);
nor U22106 (N_22106,N_13661,N_13059);
nor U22107 (N_22107,N_12191,N_14841);
nor U22108 (N_22108,N_17256,N_12479);
nor U22109 (N_22109,N_12283,N_16812);
nand U22110 (N_22110,N_16146,N_13477);
nor U22111 (N_22111,N_17613,N_15943);
nor U22112 (N_22112,N_12464,N_15760);
or U22113 (N_22113,N_17956,N_16889);
and U22114 (N_22114,N_15672,N_12923);
nor U22115 (N_22115,N_15362,N_13276);
nand U22116 (N_22116,N_13629,N_15168);
and U22117 (N_22117,N_13546,N_13045);
nor U22118 (N_22118,N_16627,N_16836);
and U22119 (N_22119,N_13854,N_14047);
nand U22120 (N_22120,N_17480,N_16866);
nand U22121 (N_22121,N_12353,N_12837);
or U22122 (N_22122,N_17990,N_17565);
and U22123 (N_22123,N_13941,N_16940);
nand U22124 (N_22124,N_16083,N_14134);
nor U22125 (N_22125,N_16070,N_13830);
xnor U22126 (N_22126,N_17457,N_16117);
and U22127 (N_22127,N_15353,N_17998);
nor U22128 (N_22128,N_16285,N_14018);
or U22129 (N_22129,N_15865,N_12405);
nand U22130 (N_22130,N_12982,N_12111);
or U22131 (N_22131,N_15300,N_15350);
or U22132 (N_22132,N_15884,N_16284);
nor U22133 (N_22133,N_15295,N_15788);
xnor U22134 (N_22134,N_17412,N_14547);
and U22135 (N_22135,N_14268,N_12148);
or U22136 (N_22136,N_14276,N_12117);
or U22137 (N_22137,N_12735,N_12076);
nand U22138 (N_22138,N_14786,N_14010);
and U22139 (N_22139,N_14829,N_15883);
nor U22140 (N_22140,N_14560,N_14631);
or U22141 (N_22141,N_13691,N_13374);
nand U22142 (N_22142,N_12574,N_15341);
and U22143 (N_22143,N_12400,N_16512);
nor U22144 (N_22144,N_12285,N_14225);
and U22145 (N_22145,N_12426,N_13494);
nand U22146 (N_22146,N_13849,N_15743);
nor U22147 (N_22147,N_13709,N_14625);
nor U22148 (N_22148,N_14932,N_12856);
nand U22149 (N_22149,N_16804,N_15039);
xor U22150 (N_22150,N_13807,N_13565);
and U22151 (N_22151,N_14357,N_14733);
or U22152 (N_22152,N_16257,N_15498);
nor U22153 (N_22153,N_13588,N_16087);
and U22154 (N_22154,N_14551,N_17314);
nor U22155 (N_22155,N_14139,N_14027);
xnor U22156 (N_22156,N_15314,N_17090);
nand U22157 (N_22157,N_17292,N_17125);
or U22158 (N_22158,N_12287,N_12860);
and U22159 (N_22159,N_14545,N_16284);
nor U22160 (N_22160,N_15486,N_17021);
and U22161 (N_22161,N_16376,N_16218);
and U22162 (N_22162,N_14721,N_12115);
nor U22163 (N_22163,N_14544,N_15716);
nor U22164 (N_22164,N_14985,N_13106);
nand U22165 (N_22165,N_16523,N_14189);
and U22166 (N_22166,N_15171,N_16796);
nor U22167 (N_22167,N_17725,N_17240);
and U22168 (N_22168,N_13261,N_16224);
and U22169 (N_22169,N_17832,N_15265);
nand U22170 (N_22170,N_13449,N_12908);
nand U22171 (N_22171,N_13420,N_16339);
nand U22172 (N_22172,N_12616,N_15802);
xor U22173 (N_22173,N_15680,N_14046);
nand U22174 (N_22174,N_14018,N_17656);
nand U22175 (N_22175,N_13317,N_12640);
nand U22176 (N_22176,N_12346,N_16538);
nor U22177 (N_22177,N_12265,N_12792);
or U22178 (N_22178,N_12241,N_13913);
and U22179 (N_22179,N_12263,N_16690);
xor U22180 (N_22180,N_17741,N_13177);
nor U22181 (N_22181,N_13497,N_16288);
nor U22182 (N_22182,N_13151,N_16115);
nand U22183 (N_22183,N_13284,N_13892);
nand U22184 (N_22184,N_14742,N_16143);
and U22185 (N_22185,N_14065,N_15262);
nor U22186 (N_22186,N_13834,N_14874);
nor U22187 (N_22187,N_15917,N_14542);
nand U22188 (N_22188,N_15188,N_16231);
nand U22189 (N_22189,N_16207,N_12141);
nor U22190 (N_22190,N_16920,N_17455);
nor U22191 (N_22191,N_14884,N_13208);
and U22192 (N_22192,N_13920,N_15439);
or U22193 (N_22193,N_14620,N_16839);
xnor U22194 (N_22194,N_13059,N_14432);
and U22195 (N_22195,N_15780,N_12222);
nor U22196 (N_22196,N_13715,N_13247);
nand U22197 (N_22197,N_12808,N_14041);
or U22198 (N_22198,N_13559,N_14822);
nor U22199 (N_22199,N_13064,N_13578);
or U22200 (N_22200,N_15958,N_15943);
xnor U22201 (N_22201,N_14568,N_13333);
nand U22202 (N_22202,N_16389,N_17592);
or U22203 (N_22203,N_12826,N_12763);
and U22204 (N_22204,N_13138,N_12937);
nor U22205 (N_22205,N_13165,N_16534);
nor U22206 (N_22206,N_17538,N_16238);
xor U22207 (N_22207,N_15488,N_17004);
or U22208 (N_22208,N_14426,N_15533);
nor U22209 (N_22209,N_12234,N_13505);
nand U22210 (N_22210,N_16004,N_14512);
xor U22211 (N_22211,N_13869,N_17851);
xnor U22212 (N_22212,N_13137,N_16767);
nand U22213 (N_22213,N_12653,N_13425);
and U22214 (N_22214,N_17822,N_15450);
nor U22215 (N_22215,N_12755,N_16861);
and U22216 (N_22216,N_17662,N_16890);
or U22217 (N_22217,N_15505,N_13235);
nand U22218 (N_22218,N_13390,N_17745);
nor U22219 (N_22219,N_13869,N_17328);
nand U22220 (N_22220,N_16867,N_14469);
nor U22221 (N_22221,N_12421,N_17097);
nand U22222 (N_22222,N_13403,N_17734);
nor U22223 (N_22223,N_13935,N_13823);
or U22224 (N_22224,N_15142,N_13526);
or U22225 (N_22225,N_14241,N_13426);
nor U22226 (N_22226,N_15749,N_13359);
nand U22227 (N_22227,N_16236,N_12449);
nand U22228 (N_22228,N_14933,N_15055);
nor U22229 (N_22229,N_17920,N_17341);
nor U22230 (N_22230,N_17893,N_16208);
nand U22231 (N_22231,N_17971,N_14658);
and U22232 (N_22232,N_15870,N_12158);
and U22233 (N_22233,N_16116,N_17593);
nand U22234 (N_22234,N_14751,N_14188);
nor U22235 (N_22235,N_13538,N_15138);
or U22236 (N_22236,N_12033,N_17141);
and U22237 (N_22237,N_13414,N_13312);
nand U22238 (N_22238,N_15285,N_16246);
nand U22239 (N_22239,N_17958,N_17283);
nor U22240 (N_22240,N_14568,N_13526);
nand U22241 (N_22241,N_17232,N_13951);
nand U22242 (N_22242,N_16627,N_16748);
and U22243 (N_22243,N_15375,N_15627);
nor U22244 (N_22244,N_14742,N_12335);
and U22245 (N_22245,N_17309,N_13227);
nor U22246 (N_22246,N_14651,N_14286);
nand U22247 (N_22247,N_16434,N_16052);
xor U22248 (N_22248,N_12169,N_17245);
nand U22249 (N_22249,N_12055,N_13926);
nor U22250 (N_22250,N_17506,N_12851);
or U22251 (N_22251,N_13483,N_13489);
and U22252 (N_22252,N_14369,N_12424);
nand U22253 (N_22253,N_13576,N_12203);
and U22254 (N_22254,N_15656,N_15136);
nand U22255 (N_22255,N_12837,N_16830);
nand U22256 (N_22256,N_16731,N_13671);
and U22257 (N_22257,N_16968,N_14630);
or U22258 (N_22258,N_12649,N_15492);
nor U22259 (N_22259,N_15589,N_14369);
and U22260 (N_22260,N_16913,N_14781);
xnor U22261 (N_22261,N_16902,N_14189);
nand U22262 (N_22262,N_15440,N_13940);
and U22263 (N_22263,N_17905,N_16454);
nand U22264 (N_22264,N_17803,N_13806);
and U22265 (N_22265,N_12270,N_17943);
or U22266 (N_22266,N_16733,N_16100);
nor U22267 (N_22267,N_12699,N_12294);
nor U22268 (N_22268,N_13461,N_16415);
nor U22269 (N_22269,N_16613,N_13650);
nand U22270 (N_22270,N_17865,N_14105);
nand U22271 (N_22271,N_14098,N_12294);
or U22272 (N_22272,N_12738,N_17421);
nand U22273 (N_22273,N_15187,N_13433);
xnor U22274 (N_22274,N_12566,N_12406);
or U22275 (N_22275,N_16540,N_13460);
and U22276 (N_22276,N_13025,N_17035);
nor U22277 (N_22277,N_14269,N_12422);
or U22278 (N_22278,N_15949,N_12034);
and U22279 (N_22279,N_17435,N_12268);
nand U22280 (N_22280,N_16553,N_17047);
xnor U22281 (N_22281,N_16072,N_16708);
and U22282 (N_22282,N_14857,N_17296);
nor U22283 (N_22283,N_12092,N_16346);
or U22284 (N_22284,N_12272,N_13091);
nand U22285 (N_22285,N_13704,N_16793);
nand U22286 (N_22286,N_13633,N_17473);
nand U22287 (N_22287,N_14387,N_14088);
xnor U22288 (N_22288,N_15826,N_15785);
nand U22289 (N_22289,N_14865,N_13720);
or U22290 (N_22290,N_15386,N_13190);
xor U22291 (N_22291,N_12339,N_15741);
nor U22292 (N_22292,N_17284,N_13981);
or U22293 (N_22293,N_17998,N_12174);
or U22294 (N_22294,N_17659,N_14792);
nand U22295 (N_22295,N_12481,N_12060);
or U22296 (N_22296,N_15183,N_14782);
nor U22297 (N_22297,N_15383,N_12911);
nand U22298 (N_22298,N_14607,N_15693);
nand U22299 (N_22299,N_12323,N_14101);
nor U22300 (N_22300,N_14793,N_16360);
or U22301 (N_22301,N_14082,N_15029);
and U22302 (N_22302,N_12295,N_17414);
nand U22303 (N_22303,N_12758,N_13081);
and U22304 (N_22304,N_13171,N_13078);
or U22305 (N_22305,N_12079,N_13939);
nand U22306 (N_22306,N_15846,N_12499);
and U22307 (N_22307,N_16786,N_17593);
nand U22308 (N_22308,N_15408,N_14594);
or U22309 (N_22309,N_14628,N_17758);
or U22310 (N_22310,N_12115,N_12952);
nor U22311 (N_22311,N_14129,N_16057);
nand U22312 (N_22312,N_12970,N_16311);
nor U22313 (N_22313,N_16993,N_14198);
or U22314 (N_22314,N_14357,N_12780);
or U22315 (N_22315,N_17542,N_17372);
and U22316 (N_22316,N_14290,N_16984);
nor U22317 (N_22317,N_12768,N_16070);
xnor U22318 (N_22318,N_14386,N_17297);
nand U22319 (N_22319,N_12111,N_13537);
and U22320 (N_22320,N_17285,N_17674);
nor U22321 (N_22321,N_13686,N_16600);
xor U22322 (N_22322,N_13997,N_13306);
and U22323 (N_22323,N_17044,N_17408);
nand U22324 (N_22324,N_12277,N_16784);
nand U22325 (N_22325,N_17532,N_15823);
nand U22326 (N_22326,N_14531,N_16005);
nor U22327 (N_22327,N_16845,N_16534);
nor U22328 (N_22328,N_14706,N_15113);
and U22329 (N_22329,N_14950,N_17684);
nand U22330 (N_22330,N_13082,N_17574);
nor U22331 (N_22331,N_14910,N_16301);
or U22332 (N_22332,N_12974,N_17393);
or U22333 (N_22333,N_14759,N_16544);
or U22334 (N_22334,N_12243,N_12752);
xor U22335 (N_22335,N_12333,N_17633);
nand U22336 (N_22336,N_13459,N_14758);
and U22337 (N_22337,N_13995,N_14473);
nand U22338 (N_22338,N_17026,N_12285);
xor U22339 (N_22339,N_15345,N_14660);
nor U22340 (N_22340,N_12295,N_15792);
and U22341 (N_22341,N_16935,N_13342);
and U22342 (N_22342,N_15277,N_16303);
nand U22343 (N_22343,N_14560,N_13562);
nand U22344 (N_22344,N_12221,N_16434);
and U22345 (N_22345,N_12765,N_15382);
nor U22346 (N_22346,N_15312,N_12666);
and U22347 (N_22347,N_17846,N_16313);
xnor U22348 (N_22348,N_14190,N_17107);
xor U22349 (N_22349,N_12329,N_16491);
and U22350 (N_22350,N_12258,N_13003);
xor U22351 (N_22351,N_12895,N_16086);
nand U22352 (N_22352,N_17000,N_12242);
or U22353 (N_22353,N_17408,N_15166);
nor U22354 (N_22354,N_14537,N_14160);
nor U22355 (N_22355,N_16015,N_12451);
and U22356 (N_22356,N_14577,N_16538);
and U22357 (N_22357,N_16759,N_13762);
or U22358 (N_22358,N_16795,N_17961);
nor U22359 (N_22359,N_17383,N_12886);
or U22360 (N_22360,N_12268,N_16117);
and U22361 (N_22361,N_16635,N_13522);
or U22362 (N_22362,N_14524,N_17650);
or U22363 (N_22363,N_15276,N_14572);
or U22364 (N_22364,N_16164,N_16512);
or U22365 (N_22365,N_15008,N_13607);
nor U22366 (N_22366,N_15435,N_15186);
or U22367 (N_22367,N_13179,N_13146);
nor U22368 (N_22368,N_17478,N_13481);
nor U22369 (N_22369,N_17884,N_12117);
xnor U22370 (N_22370,N_16731,N_15244);
xor U22371 (N_22371,N_14089,N_13492);
nor U22372 (N_22372,N_17265,N_14791);
or U22373 (N_22373,N_12848,N_15900);
or U22374 (N_22374,N_15018,N_17570);
nand U22375 (N_22375,N_13640,N_13419);
or U22376 (N_22376,N_17495,N_12552);
or U22377 (N_22377,N_14538,N_16747);
nor U22378 (N_22378,N_14408,N_13992);
or U22379 (N_22379,N_12432,N_14455);
nor U22380 (N_22380,N_16648,N_12312);
nand U22381 (N_22381,N_12094,N_12172);
nand U22382 (N_22382,N_12504,N_17407);
nor U22383 (N_22383,N_13749,N_17436);
xor U22384 (N_22384,N_14116,N_15028);
or U22385 (N_22385,N_16675,N_15665);
nor U22386 (N_22386,N_16850,N_12409);
xnor U22387 (N_22387,N_14463,N_17879);
or U22388 (N_22388,N_16194,N_15708);
nand U22389 (N_22389,N_14377,N_13797);
nor U22390 (N_22390,N_14167,N_17345);
nand U22391 (N_22391,N_13106,N_14348);
nor U22392 (N_22392,N_17552,N_17772);
and U22393 (N_22393,N_14286,N_15514);
or U22394 (N_22394,N_14643,N_12349);
or U22395 (N_22395,N_14410,N_16966);
and U22396 (N_22396,N_12116,N_14588);
nor U22397 (N_22397,N_16183,N_12073);
nand U22398 (N_22398,N_15472,N_14015);
nor U22399 (N_22399,N_16304,N_14853);
nor U22400 (N_22400,N_17246,N_15085);
xor U22401 (N_22401,N_15124,N_15295);
nand U22402 (N_22402,N_12724,N_15054);
or U22403 (N_22403,N_15283,N_15550);
and U22404 (N_22404,N_15655,N_15588);
nor U22405 (N_22405,N_13349,N_12037);
xor U22406 (N_22406,N_15472,N_12663);
or U22407 (N_22407,N_14777,N_16168);
nand U22408 (N_22408,N_15326,N_13608);
nor U22409 (N_22409,N_15466,N_13598);
and U22410 (N_22410,N_15766,N_15590);
nor U22411 (N_22411,N_13904,N_17010);
and U22412 (N_22412,N_17206,N_14858);
or U22413 (N_22413,N_16615,N_15523);
xnor U22414 (N_22414,N_16395,N_12874);
or U22415 (N_22415,N_17644,N_15120);
xor U22416 (N_22416,N_13529,N_15520);
nor U22417 (N_22417,N_14182,N_13297);
nor U22418 (N_22418,N_17986,N_15693);
nand U22419 (N_22419,N_16901,N_14148);
and U22420 (N_22420,N_13085,N_15795);
and U22421 (N_22421,N_15078,N_17107);
and U22422 (N_22422,N_14889,N_15780);
nor U22423 (N_22423,N_15655,N_16161);
or U22424 (N_22424,N_14400,N_17613);
or U22425 (N_22425,N_13261,N_13800);
nand U22426 (N_22426,N_15711,N_14731);
nor U22427 (N_22427,N_16753,N_16637);
nand U22428 (N_22428,N_17265,N_12218);
nand U22429 (N_22429,N_17435,N_17357);
and U22430 (N_22430,N_12242,N_15534);
or U22431 (N_22431,N_12022,N_15391);
nand U22432 (N_22432,N_13693,N_17156);
and U22433 (N_22433,N_13469,N_17410);
nand U22434 (N_22434,N_14167,N_12313);
nand U22435 (N_22435,N_12646,N_16487);
nand U22436 (N_22436,N_15996,N_12626);
nor U22437 (N_22437,N_15233,N_17168);
and U22438 (N_22438,N_12837,N_17819);
and U22439 (N_22439,N_13738,N_14132);
or U22440 (N_22440,N_17325,N_16192);
or U22441 (N_22441,N_17298,N_12152);
and U22442 (N_22442,N_16968,N_17441);
or U22443 (N_22443,N_14752,N_12914);
nand U22444 (N_22444,N_14165,N_16182);
and U22445 (N_22445,N_16444,N_12872);
or U22446 (N_22446,N_16155,N_13836);
and U22447 (N_22447,N_12117,N_14156);
and U22448 (N_22448,N_17549,N_14005);
nand U22449 (N_22449,N_15740,N_15546);
xnor U22450 (N_22450,N_15832,N_15799);
nor U22451 (N_22451,N_12653,N_12248);
and U22452 (N_22452,N_13953,N_13139);
nand U22453 (N_22453,N_15320,N_13321);
nand U22454 (N_22454,N_15691,N_16163);
nand U22455 (N_22455,N_13252,N_14460);
nand U22456 (N_22456,N_15630,N_14624);
nand U22457 (N_22457,N_14021,N_12170);
nand U22458 (N_22458,N_13570,N_15195);
or U22459 (N_22459,N_14931,N_16145);
and U22460 (N_22460,N_15922,N_15775);
and U22461 (N_22461,N_14204,N_16500);
nor U22462 (N_22462,N_16811,N_15027);
or U22463 (N_22463,N_15948,N_13388);
or U22464 (N_22464,N_17986,N_16316);
and U22465 (N_22465,N_15308,N_17763);
or U22466 (N_22466,N_13523,N_13499);
or U22467 (N_22467,N_14080,N_15005);
nand U22468 (N_22468,N_17954,N_15503);
nand U22469 (N_22469,N_13934,N_15212);
nor U22470 (N_22470,N_12511,N_12063);
nor U22471 (N_22471,N_16968,N_14716);
xnor U22472 (N_22472,N_16376,N_15528);
and U22473 (N_22473,N_17917,N_16325);
nand U22474 (N_22474,N_13285,N_17003);
nand U22475 (N_22475,N_15016,N_12316);
nand U22476 (N_22476,N_17696,N_15022);
nor U22477 (N_22477,N_16575,N_12702);
nor U22478 (N_22478,N_12908,N_15824);
or U22479 (N_22479,N_14578,N_12487);
xnor U22480 (N_22480,N_13797,N_13212);
and U22481 (N_22481,N_15614,N_12121);
or U22482 (N_22482,N_15249,N_13870);
nand U22483 (N_22483,N_16407,N_15831);
or U22484 (N_22484,N_13393,N_17488);
or U22485 (N_22485,N_17573,N_16562);
and U22486 (N_22486,N_14955,N_15149);
nor U22487 (N_22487,N_15458,N_15082);
xor U22488 (N_22488,N_17726,N_17281);
nor U22489 (N_22489,N_17213,N_14076);
and U22490 (N_22490,N_15202,N_13310);
nand U22491 (N_22491,N_16269,N_14035);
and U22492 (N_22492,N_14459,N_12584);
nand U22493 (N_22493,N_17695,N_17754);
xnor U22494 (N_22494,N_17953,N_17729);
nor U22495 (N_22495,N_16347,N_15671);
nor U22496 (N_22496,N_13173,N_13782);
nor U22497 (N_22497,N_17897,N_13450);
or U22498 (N_22498,N_13899,N_17544);
nor U22499 (N_22499,N_12676,N_14908);
nand U22500 (N_22500,N_13678,N_14831);
and U22501 (N_22501,N_15000,N_14242);
and U22502 (N_22502,N_16460,N_13435);
or U22503 (N_22503,N_12352,N_16952);
nor U22504 (N_22504,N_17077,N_13873);
nor U22505 (N_22505,N_16119,N_13134);
nand U22506 (N_22506,N_13377,N_17331);
or U22507 (N_22507,N_14098,N_12602);
or U22508 (N_22508,N_13621,N_17672);
nand U22509 (N_22509,N_17175,N_12273);
nand U22510 (N_22510,N_17227,N_17068);
nor U22511 (N_22511,N_16066,N_16447);
and U22512 (N_22512,N_17590,N_14986);
nor U22513 (N_22513,N_15815,N_15880);
or U22514 (N_22514,N_16929,N_12502);
nand U22515 (N_22515,N_15931,N_13071);
and U22516 (N_22516,N_14173,N_17003);
and U22517 (N_22517,N_13994,N_17773);
and U22518 (N_22518,N_16644,N_13926);
or U22519 (N_22519,N_17806,N_12249);
or U22520 (N_22520,N_16842,N_14554);
nor U22521 (N_22521,N_12223,N_14348);
and U22522 (N_22522,N_13146,N_15719);
or U22523 (N_22523,N_12882,N_13948);
nand U22524 (N_22524,N_16050,N_16393);
nor U22525 (N_22525,N_16699,N_13659);
or U22526 (N_22526,N_16234,N_15458);
or U22527 (N_22527,N_13290,N_16121);
nand U22528 (N_22528,N_16821,N_15785);
or U22529 (N_22529,N_13129,N_12996);
nor U22530 (N_22530,N_15533,N_14357);
nor U22531 (N_22531,N_12372,N_12198);
nand U22532 (N_22532,N_15149,N_12471);
nand U22533 (N_22533,N_12912,N_15412);
nor U22534 (N_22534,N_16406,N_16699);
nand U22535 (N_22535,N_16944,N_12351);
nor U22536 (N_22536,N_15538,N_14820);
or U22537 (N_22537,N_16355,N_13440);
nor U22538 (N_22538,N_13669,N_13519);
and U22539 (N_22539,N_12503,N_17431);
nor U22540 (N_22540,N_15835,N_15144);
nand U22541 (N_22541,N_16440,N_17828);
and U22542 (N_22542,N_16005,N_16802);
and U22543 (N_22543,N_16258,N_14163);
and U22544 (N_22544,N_14350,N_17784);
nand U22545 (N_22545,N_16101,N_17924);
or U22546 (N_22546,N_16436,N_17243);
nand U22547 (N_22547,N_17372,N_17640);
xor U22548 (N_22548,N_16994,N_14407);
xnor U22549 (N_22549,N_12712,N_12357);
and U22550 (N_22550,N_15761,N_15831);
nand U22551 (N_22551,N_12717,N_13149);
xnor U22552 (N_22552,N_14072,N_16872);
and U22553 (N_22553,N_13101,N_13007);
nor U22554 (N_22554,N_12859,N_17555);
and U22555 (N_22555,N_17435,N_15614);
and U22556 (N_22556,N_17254,N_14046);
nand U22557 (N_22557,N_15577,N_16124);
or U22558 (N_22558,N_17049,N_16295);
nor U22559 (N_22559,N_14414,N_17161);
xnor U22560 (N_22560,N_14966,N_14040);
nand U22561 (N_22561,N_13350,N_17007);
and U22562 (N_22562,N_17520,N_14863);
nor U22563 (N_22563,N_13224,N_13532);
nand U22564 (N_22564,N_14053,N_17274);
nor U22565 (N_22565,N_17766,N_13412);
or U22566 (N_22566,N_12663,N_15105);
or U22567 (N_22567,N_17815,N_15333);
nand U22568 (N_22568,N_12100,N_14963);
and U22569 (N_22569,N_15600,N_12397);
nand U22570 (N_22570,N_13716,N_16197);
nor U22571 (N_22571,N_16743,N_12533);
or U22572 (N_22572,N_15019,N_17639);
nand U22573 (N_22573,N_17375,N_14030);
and U22574 (N_22574,N_17203,N_14033);
xnor U22575 (N_22575,N_12636,N_17108);
and U22576 (N_22576,N_16367,N_14079);
and U22577 (N_22577,N_17026,N_13124);
nand U22578 (N_22578,N_13298,N_13549);
nand U22579 (N_22579,N_15977,N_14648);
and U22580 (N_22580,N_12391,N_16646);
nor U22581 (N_22581,N_15296,N_17652);
and U22582 (N_22582,N_15913,N_14036);
xor U22583 (N_22583,N_14146,N_12514);
nor U22584 (N_22584,N_15298,N_12772);
and U22585 (N_22585,N_16631,N_13281);
nor U22586 (N_22586,N_12989,N_15673);
or U22587 (N_22587,N_16338,N_15649);
or U22588 (N_22588,N_17972,N_12024);
xor U22589 (N_22589,N_13439,N_12659);
nand U22590 (N_22590,N_15307,N_17865);
nor U22591 (N_22591,N_13902,N_14896);
nor U22592 (N_22592,N_13181,N_15185);
nor U22593 (N_22593,N_16850,N_16534);
nand U22594 (N_22594,N_17247,N_12619);
and U22595 (N_22595,N_12766,N_13244);
or U22596 (N_22596,N_15917,N_17381);
and U22597 (N_22597,N_15203,N_13369);
nor U22598 (N_22598,N_15836,N_12486);
or U22599 (N_22599,N_15179,N_16119);
nor U22600 (N_22600,N_12377,N_14744);
nor U22601 (N_22601,N_14454,N_16858);
or U22602 (N_22602,N_15692,N_12320);
nor U22603 (N_22603,N_14109,N_15746);
nor U22604 (N_22604,N_14117,N_16072);
nor U22605 (N_22605,N_14358,N_14326);
nor U22606 (N_22606,N_12235,N_12776);
nor U22607 (N_22607,N_12657,N_17360);
or U22608 (N_22608,N_16782,N_16850);
and U22609 (N_22609,N_12446,N_16599);
nand U22610 (N_22610,N_17363,N_17080);
nand U22611 (N_22611,N_14983,N_13252);
xor U22612 (N_22612,N_15360,N_14001);
and U22613 (N_22613,N_17051,N_12064);
nor U22614 (N_22614,N_13576,N_17083);
nor U22615 (N_22615,N_14716,N_16242);
nand U22616 (N_22616,N_17499,N_17171);
nor U22617 (N_22617,N_16143,N_12994);
nand U22618 (N_22618,N_13167,N_13823);
and U22619 (N_22619,N_17921,N_15953);
nor U22620 (N_22620,N_17382,N_13501);
nand U22621 (N_22621,N_12819,N_13650);
nand U22622 (N_22622,N_16034,N_12230);
or U22623 (N_22623,N_16919,N_15564);
nor U22624 (N_22624,N_12716,N_17176);
nand U22625 (N_22625,N_17298,N_13705);
nor U22626 (N_22626,N_12378,N_12421);
nor U22627 (N_22627,N_12032,N_16541);
or U22628 (N_22628,N_13801,N_16993);
and U22629 (N_22629,N_17534,N_14427);
and U22630 (N_22630,N_12557,N_14589);
nand U22631 (N_22631,N_16558,N_17721);
or U22632 (N_22632,N_17532,N_12409);
nor U22633 (N_22633,N_14071,N_16472);
and U22634 (N_22634,N_14310,N_14348);
nor U22635 (N_22635,N_15765,N_12095);
nand U22636 (N_22636,N_16927,N_17706);
nor U22637 (N_22637,N_13908,N_15887);
or U22638 (N_22638,N_16253,N_13604);
or U22639 (N_22639,N_15551,N_12473);
and U22640 (N_22640,N_17599,N_12405);
nor U22641 (N_22641,N_14348,N_13924);
nor U22642 (N_22642,N_15849,N_17277);
or U22643 (N_22643,N_14654,N_17727);
nand U22644 (N_22644,N_14690,N_17128);
xnor U22645 (N_22645,N_15074,N_14909);
and U22646 (N_22646,N_15575,N_12738);
nor U22647 (N_22647,N_12817,N_12549);
nand U22648 (N_22648,N_13583,N_12880);
nor U22649 (N_22649,N_17102,N_12042);
and U22650 (N_22650,N_14361,N_14715);
nand U22651 (N_22651,N_15913,N_16644);
or U22652 (N_22652,N_12809,N_14213);
nand U22653 (N_22653,N_12570,N_16128);
xor U22654 (N_22654,N_15223,N_13628);
nand U22655 (N_22655,N_16561,N_16607);
nand U22656 (N_22656,N_17054,N_16728);
nand U22657 (N_22657,N_17805,N_14906);
and U22658 (N_22658,N_14539,N_15504);
and U22659 (N_22659,N_16862,N_17653);
and U22660 (N_22660,N_14683,N_14682);
nand U22661 (N_22661,N_12113,N_16572);
or U22662 (N_22662,N_15003,N_15071);
nor U22663 (N_22663,N_14500,N_15793);
nand U22664 (N_22664,N_16712,N_12961);
nor U22665 (N_22665,N_17583,N_16225);
or U22666 (N_22666,N_17868,N_15352);
nor U22667 (N_22667,N_16094,N_15128);
nor U22668 (N_22668,N_17017,N_16868);
nor U22669 (N_22669,N_14828,N_16108);
or U22670 (N_22670,N_14692,N_15705);
nand U22671 (N_22671,N_16953,N_14223);
or U22672 (N_22672,N_16903,N_13719);
or U22673 (N_22673,N_17571,N_16306);
nor U22674 (N_22674,N_12370,N_17303);
or U22675 (N_22675,N_16426,N_17710);
nor U22676 (N_22676,N_15538,N_16723);
nand U22677 (N_22677,N_14737,N_14936);
nand U22678 (N_22678,N_13146,N_15433);
or U22679 (N_22679,N_16187,N_14069);
and U22680 (N_22680,N_15259,N_15486);
nand U22681 (N_22681,N_13512,N_14194);
nand U22682 (N_22682,N_17071,N_15104);
nand U22683 (N_22683,N_17894,N_17887);
nand U22684 (N_22684,N_13484,N_15185);
nor U22685 (N_22685,N_12906,N_17003);
nor U22686 (N_22686,N_16926,N_12199);
nor U22687 (N_22687,N_12767,N_14474);
and U22688 (N_22688,N_16007,N_17173);
and U22689 (N_22689,N_13228,N_12604);
nor U22690 (N_22690,N_17217,N_16561);
and U22691 (N_22691,N_13268,N_13260);
xor U22692 (N_22692,N_14135,N_16769);
and U22693 (N_22693,N_14048,N_13555);
and U22694 (N_22694,N_16881,N_12796);
and U22695 (N_22695,N_13841,N_17038);
xor U22696 (N_22696,N_12585,N_17309);
or U22697 (N_22697,N_15628,N_17085);
or U22698 (N_22698,N_17938,N_12204);
or U22699 (N_22699,N_15323,N_13220);
xnor U22700 (N_22700,N_15251,N_13291);
nor U22701 (N_22701,N_12929,N_15272);
nor U22702 (N_22702,N_12093,N_15672);
nand U22703 (N_22703,N_16437,N_17714);
and U22704 (N_22704,N_15093,N_12328);
nor U22705 (N_22705,N_13370,N_16057);
nor U22706 (N_22706,N_16709,N_12142);
and U22707 (N_22707,N_17578,N_15127);
and U22708 (N_22708,N_16229,N_13367);
and U22709 (N_22709,N_12270,N_13868);
or U22710 (N_22710,N_15174,N_12077);
nor U22711 (N_22711,N_15075,N_17678);
or U22712 (N_22712,N_15924,N_13140);
or U22713 (N_22713,N_13287,N_14244);
and U22714 (N_22714,N_13615,N_13585);
nand U22715 (N_22715,N_13070,N_14600);
and U22716 (N_22716,N_17252,N_13241);
nand U22717 (N_22717,N_15903,N_16161);
nand U22718 (N_22718,N_15479,N_14327);
nor U22719 (N_22719,N_12480,N_17097);
and U22720 (N_22720,N_17400,N_15253);
and U22721 (N_22721,N_15427,N_16564);
and U22722 (N_22722,N_14789,N_17809);
nand U22723 (N_22723,N_14252,N_17819);
or U22724 (N_22724,N_14373,N_17534);
or U22725 (N_22725,N_16234,N_16487);
xnor U22726 (N_22726,N_16569,N_15937);
nand U22727 (N_22727,N_12684,N_13887);
or U22728 (N_22728,N_16551,N_16591);
nor U22729 (N_22729,N_16460,N_14103);
nor U22730 (N_22730,N_13945,N_15489);
or U22731 (N_22731,N_15557,N_16743);
nand U22732 (N_22732,N_17558,N_17581);
and U22733 (N_22733,N_14788,N_15887);
or U22734 (N_22734,N_17360,N_13423);
nand U22735 (N_22735,N_14174,N_17800);
nor U22736 (N_22736,N_13292,N_16292);
or U22737 (N_22737,N_14900,N_12392);
and U22738 (N_22738,N_13390,N_12034);
nand U22739 (N_22739,N_15744,N_15511);
and U22740 (N_22740,N_14514,N_12424);
nand U22741 (N_22741,N_13506,N_15937);
and U22742 (N_22742,N_13938,N_14961);
nor U22743 (N_22743,N_12700,N_15676);
nor U22744 (N_22744,N_15457,N_14018);
and U22745 (N_22745,N_15795,N_13060);
nor U22746 (N_22746,N_13234,N_13995);
nand U22747 (N_22747,N_14455,N_15008);
nor U22748 (N_22748,N_15120,N_12758);
or U22749 (N_22749,N_16948,N_12223);
nor U22750 (N_22750,N_12571,N_13529);
or U22751 (N_22751,N_17453,N_13608);
nor U22752 (N_22752,N_13165,N_15943);
nor U22753 (N_22753,N_16468,N_14246);
and U22754 (N_22754,N_16524,N_17893);
and U22755 (N_22755,N_17688,N_13754);
nand U22756 (N_22756,N_17001,N_12965);
or U22757 (N_22757,N_15264,N_14696);
nand U22758 (N_22758,N_13067,N_12138);
nor U22759 (N_22759,N_14830,N_15182);
nand U22760 (N_22760,N_14454,N_13283);
nor U22761 (N_22761,N_15353,N_14420);
nand U22762 (N_22762,N_17605,N_17562);
or U22763 (N_22763,N_15035,N_15169);
xor U22764 (N_22764,N_12898,N_13987);
nand U22765 (N_22765,N_15014,N_15412);
or U22766 (N_22766,N_13702,N_17828);
nor U22767 (N_22767,N_14611,N_14018);
or U22768 (N_22768,N_16195,N_14191);
nand U22769 (N_22769,N_14724,N_16958);
nand U22770 (N_22770,N_16563,N_12071);
nor U22771 (N_22771,N_13386,N_12737);
nand U22772 (N_22772,N_16328,N_13030);
and U22773 (N_22773,N_14263,N_14166);
and U22774 (N_22774,N_16960,N_15048);
or U22775 (N_22775,N_12569,N_17460);
nor U22776 (N_22776,N_17882,N_17002);
or U22777 (N_22777,N_12051,N_12083);
nor U22778 (N_22778,N_16602,N_14762);
nor U22779 (N_22779,N_13321,N_16345);
xnor U22780 (N_22780,N_14089,N_14797);
nand U22781 (N_22781,N_16481,N_14291);
and U22782 (N_22782,N_15284,N_12916);
nor U22783 (N_22783,N_16314,N_16125);
nor U22784 (N_22784,N_15287,N_12330);
or U22785 (N_22785,N_16006,N_12728);
nand U22786 (N_22786,N_14226,N_13125);
nor U22787 (N_22787,N_17640,N_16877);
nor U22788 (N_22788,N_12723,N_13492);
nor U22789 (N_22789,N_15413,N_13500);
and U22790 (N_22790,N_16610,N_16664);
nand U22791 (N_22791,N_16493,N_15501);
and U22792 (N_22792,N_12517,N_12397);
xor U22793 (N_22793,N_17791,N_14252);
xnor U22794 (N_22794,N_12163,N_15776);
and U22795 (N_22795,N_17885,N_13990);
nand U22796 (N_22796,N_16708,N_13882);
xnor U22797 (N_22797,N_15877,N_14106);
nand U22798 (N_22798,N_12489,N_12525);
nor U22799 (N_22799,N_12212,N_16496);
nand U22800 (N_22800,N_16847,N_15954);
and U22801 (N_22801,N_16776,N_17679);
and U22802 (N_22802,N_15163,N_12131);
nand U22803 (N_22803,N_12069,N_16730);
nand U22804 (N_22804,N_13091,N_15404);
or U22805 (N_22805,N_17337,N_16752);
xor U22806 (N_22806,N_16217,N_14163);
or U22807 (N_22807,N_17502,N_16589);
xor U22808 (N_22808,N_16269,N_17457);
or U22809 (N_22809,N_14421,N_12022);
or U22810 (N_22810,N_14593,N_14354);
nand U22811 (N_22811,N_12993,N_12448);
or U22812 (N_22812,N_14924,N_12458);
or U22813 (N_22813,N_16420,N_13789);
nor U22814 (N_22814,N_13717,N_17659);
nor U22815 (N_22815,N_15985,N_17700);
or U22816 (N_22816,N_12320,N_14393);
nand U22817 (N_22817,N_14294,N_17362);
nand U22818 (N_22818,N_16105,N_16878);
and U22819 (N_22819,N_13850,N_16156);
nand U22820 (N_22820,N_14893,N_17286);
xor U22821 (N_22821,N_16338,N_16332);
nor U22822 (N_22822,N_13015,N_13792);
or U22823 (N_22823,N_15270,N_12014);
and U22824 (N_22824,N_17325,N_15370);
nor U22825 (N_22825,N_16609,N_13968);
and U22826 (N_22826,N_12959,N_16589);
nand U22827 (N_22827,N_14701,N_16666);
nor U22828 (N_22828,N_12444,N_15172);
nor U22829 (N_22829,N_12002,N_16052);
and U22830 (N_22830,N_17411,N_14686);
and U22831 (N_22831,N_14877,N_13563);
nand U22832 (N_22832,N_13680,N_16831);
or U22833 (N_22833,N_13045,N_14908);
or U22834 (N_22834,N_16929,N_12612);
or U22835 (N_22835,N_14629,N_17825);
xor U22836 (N_22836,N_15580,N_16508);
and U22837 (N_22837,N_13130,N_16919);
nand U22838 (N_22838,N_16203,N_15122);
and U22839 (N_22839,N_12789,N_12766);
and U22840 (N_22840,N_16409,N_15987);
nor U22841 (N_22841,N_15532,N_14566);
nor U22842 (N_22842,N_13503,N_15982);
and U22843 (N_22843,N_16496,N_17492);
nand U22844 (N_22844,N_13772,N_17560);
nand U22845 (N_22845,N_14287,N_12143);
nand U22846 (N_22846,N_13043,N_14502);
nand U22847 (N_22847,N_17485,N_13510);
nand U22848 (N_22848,N_12294,N_13215);
nand U22849 (N_22849,N_16832,N_15946);
nand U22850 (N_22850,N_16663,N_16129);
and U22851 (N_22851,N_13117,N_16444);
xnor U22852 (N_22852,N_13807,N_16754);
nor U22853 (N_22853,N_12872,N_12190);
or U22854 (N_22854,N_16952,N_14032);
xor U22855 (N_22855,N_17635,N_12515);
or U22856 (N_22856,N_14021,N_15675);
xor U22857 (N_22857,N_13086,N_14785);
or U22858 (N_22858,N_14661,N_14165);
nor U22859 (N_22859,N_15808,N_12278);
nand U22860 (N_22860,N_15383,N_17911);
or U22861 (N_22861,N_13947,N_13676);
nand U22862 (N_22862,N_12332,N_17987);
xor U22863 (N_22863,N_17567,N_15393);
or U22864 (N_22864,N_15990,N_16863);
nand U22865 (N_22865,N_15263,N_16404);
nor U22866 (N_22866,N_13197,N_13118);
nand U22867 (N_22867,N_14999,N_12222);
nor U22868 (N_22868,N_17100,N_13076);
or U22869 (N_22869,N_13125,N_14463);
and U22870 (N_22870,N_17071,N_12158);
and U22871 (N_22871,N_17657,N_12696);
xor U22872 (N_22872,N_16400,N_16609);
and U22873 (N_22873,N_17058,N_15674);
and U22874 (N_22874,N_14452,N_13521);
nand U22875 (N_22875,N_12580,N_12321);
or U22876 (N_22876,N_14549,N_16303);
and U22877 (N_22877,N_13470,N_16024);
nand U22878 (N_22878,N_16237,N_13290);
xor U22879 (N_22879,N_15129,N_12063);
nand U22880 (N_22880,N_16877,N_12170);
nor U22881 (N_22881,N_12682,N_15680);
nand U22882 (N_22882,N_15912,N_13290);
nor U22883 (N_22883,N_14991,N_17687);
nand U22884 (N_22884,N_12959,N_14750);
nand U22885 (N_22885,N_16733,N_16749);
or U22886 (N_22886,N_16320,N_16999);
or U22887 (N_22887,N_17510,N_13231);
nor U22888 (N_22888,N_17469,N_14091);
and U22889 (N_22889,N_14882,N_16126);
and U22890 (N_22890,N_13334,N_17311);
nor U22891 (N_22891,N_13594,N_13626);
or U22892 (N_22892,N_14278,N_17358);
nand U22893 (N_22893,N_13561,N_13540);
nand U22894 (N_22894,N_14204,N_15803);
nand U22895 (N_22895,N_15235,N_17486);
and U22896 (N_22896,N_17529,N_17035);
nor U22897 (N_22897,N_17240,N_13118);
nand U22898 (N_22898,N_13874,N_16738);
and U22899 (N_22899,N_14255,N_16567);
or U22900 (N_22900,N_14320,N_15885);
and U22901 (N_22901,N_17876,N_16777);
nand U22902 (N_22902,N_14724,N_15943);
nand U22903 (N_22903,N_17501,N_14254);
nor U22904 (N_22904,N_17495,N_13794);
nand U22905 (N_22905,N_12103,N_17607);
nand U22906 (N_22906,N_15640,N_17878);
and U22907 (N_22907,N_14091,N_12589);
and U22908 (N_22908,N_12672,N_16520);
nand U22909 (N_22909,N_16433,N_17759);
nand U22910 (N_22910,N_16871,N_15777);
nor U22911 (N_22911,N_14891,N_15416);
nor U22912 (N_22912,N_13740,N_15607);
or U22913 (N_22913,N_12690,N_12167);
and U22914 (N_22914,N_13042,N_15709);
and U22915 (N_22915,N_13500,N_14027);
nand U22916 (N_22916,N_14624,N_15950);
xor U22917 (N_22917,N_16528,N_15273);
or U22918 (N_22918,N_13130,N_12113);
nor U22919 (N_22919,N_16064,N_13130);
or U22920 (N_22920,N_16511,N_15359);
nor U22921 (N_22921,N_15478,N_15538);
or U22922 (N_22922,N_14197,N_17422);
and U22923 (N_22923,N_12081,N_14352);
nand U22924 (N_22924,N_12214,N_12442);
or U22925 (N_22925,N_17854,N_16341);
and U22926 (N_22926,N_14332,N_17464);
or U22927 (N_22927,N_13176,N_13085);
or U22928 (N_22928,N_12975,N_15325);
nor U22929 (N_22929,N_17047,N_12344);
nand U22930 (N_22930,N_17462,N_14967);
or U22931 (N_22931,N_17208,N_13821);
or U22932 (N_22932,N_16280,N_15153);
nand U22933 (N_22933,N_17523,N_15810);
nand U22934 (N_22934,N_12822,N_12617);
and U22935 (N_22935,N_17710,N_15304);
xnor U22936 (N_22936,N_12771,N_16711);
or U22937 (N_22937,N_12419,N_14587);
nand U22938 (N_22938,N_12812,N_16464);
and U22939 (N_22939,N_17626,N_12343);
nand U22940 (N_22940,N_14568,N_16426);
nand U22941 (N_22941,N_14579,N_16276);
nand U22942 (N_22942,N_13588,N_17091);
nor U22943 (N_22943,N_14203,N_17660);
nand U22944 (N_22944,N_15251,N_13815);
nand U22945 (N_22945,N_12507,N_14632);
nor U22946 (N_22946,N_17011,N_14011);
nor U22947 (N_22947,N_13808,N_13333);
and U22948 (N_22948,N_13036,N_17548);
nand U22949 (N_22949,N_12064,N_12414);
nor U22950 (N_22950,N_13729,N_15504);
nor U22951 (N_22951,N_15584,N_12971);
and U22952 (N_22952,N_14910,N_15446);
xnor U22953 (N_22953,N_15741,N_15893);
and U22954 (N_22954,N_13561,N_13222);
nor U22955 (N_22955,N_13087,N_16681);
and U22956 (N_22956,N_17117,N_17492);
or U22957 (N_22957,N_16621,N_15376);
nor U22958 (N_22958,N_15391,N_12674);
nor U22959 (N_22959,N_17760,N_13720);
nor U22960 (N_22960,N_12727,N_15202);
or U22961 (N_22961,N_16072,N_13727);
or U22962 (N_22962,N_13229,N_14946);
and U22963 (N_22963,N_14297,N_13428);
nand U22964 (N_22964,N_14245,N_14839);
xnor U22965 (N_22965,N_16804,N_12065);
and U22966 (N_22966,N_12634,N_14227);
nor U22967 (N_22967,N_15129,N_13442);
and U22968 (N_22968,N_12679,N_15408);
xor U22969 (N_22969,N_13196,N_15938);
and U22970 (N_22970,N_14680,N_16519);
or U22971 (N_22971,N_16143,N_14754);
or U22972 (N_22972,N_16566,N_17899);
nor U22973 (N_22973,N_13247,N_17988);
xnor U22974 (N_22974,N_15452,N_17995);
nand U22975 (N_22975,N_16863,N_15299);
and U22976 (N_22976,N_12022,N_13399);
nor U22977 (N_22977,N_16902,N_13033);
nor U22978 (N_22978,N_12612,N_14704);
nand U22979 (N_22979,N_14669,N_14309);
nand U22980 (N_22980,N_12704,N_15299);
xnor U22981 (N_22981,N_17722,N_17877);
and U22982 (N_22982,N_17800,N_12077);
nand U22983 (N_22983,N_13157,N_13257);
nand U22984 (N_22984,N_17791,N_15713);
nand U22985 (N_22985,N_12952,N_16696);
or U22986 (N_22986,N_16038,N_12846);
nor U22987 (N_22987,N_17197,N_16113);
nand U22988 (N_22988,N_14198,N_14318);
and U22989 (N_22989,N_14094,N_13328);
nor U22990 (N_22990,N_15343,N_13790);
nand U22991 (N_22991,N_13765,N_13263);
and U22992 (N_22992,N_15537,N_14435);
xnor U22993 (N_22993,N_16923,N_15824);
nor U22994 (N_22994,N_16610,N_13825);
nor U22995 (N_22995,N_17175,N_13825);
and U22996 (N_22996,N_14623,N_17747);
and U22997 (N_22997,N_17060,N_16204);
nor U22998 (N_22998,N_15643,N_12955);
or U22999 (N_22999,N_14247,N_16640);
nor U23000 (N_23000,N_17530,N_15362);
nor U23001 (N_23001,N_13999,N_15206);
or U23002 (N_23002,N_13690,N_14200);
nand U23003 (N_23003,N_16203,N_13239);
nand U23004 (N_23004,N_13062,N_12442);
and U23005 (N_23005,N_13348,N_12509);
xor U23006 (N_23006,N_13877,N_14508);
nor U23007 (N_23007,N_14371,N_12278);
or U23008 (N_23008,N_17365,N_15537);
xnor U23009 (N_23009,N_16370,N_15233);
nand U23010 (N_23010,N_14013,N_12387);
and U23011 (N_23011,N_14206,N_12583);
nor U23012 (N_23012,N_17017,N_13574);
nand U23013 (N_23013,N_13704,N_12745);
or U23014 (N_23014,N_14142,N_15274);
nand U23015 (N_23015,N_15275,N_13600);
and U23016 (N_23016,N_12676,N_15725);
nor U23017 (N_23017,N_14496,N_15566);
and U23018 (N_23018,N_13160,N_13174);
nor U23019 (N_23019,N_15955,N_14425);
or U23020 (N_23020,N_16469,N_16743);
nor U23021 (N_23021,N_15610,N_15701);
nand U23022 (N_23022,N_12959,N_12398);
nand U23023 (N_23023,N_17423,N_15357);
or U23024 (N_23024,N_16968,N_16864);
and U23025 (N_23025,N_14631,N_16037);
xnor U23026 (N_23026,N_15506,N_16996);
or U23027 (N_23027,N_13648,N_17328);
or U23028 (N_23028,N_12591,N_15789);
xor U23029 (N_23029,N_14916,N_15021);
or U23030 (N_23030,N_14686,N_16788);
and U23031 (N_23031,N_15057,N_12081);
xnor U23032 (N_23032,N_14320,N_14844);
nand U23033 (N_23033,N_17431,N_17166);
or U23034 (N_23034,N_17744,N_15197);
nor U23035 (N_23035,N_14551,N_14163);
and U23036 (N_23036,N_15798,N_15435);
nor U23037 (N_23037,N_14344,N_17724);
nor U23038 (N_23038,N_17201,N_13006);
and U23039 (N_23039,N_16973,N_16108);
nand U23040 (N_23040,N_14192,N_14627);
or U23041 (N_23041,N_13875,N_17901);
or U23042 (N_23042,N_13757,N_14966);
nand U23043 (N_23043,N_16222,N_15239);
nor U23044 (N_23044,N_15108,N_15491);
xor U23045 (N_23045,N_16854,N_14553);
or U23046 (N_23046,N_17228,N_16185);
or U23047 (N_23047,N_15126,N_12360);
nor U23048 (N_23048,N_13022,N_14192);
or U23049 (N_23049,N_14618,N_15459);
nand U23050 (N_23050,N_16179,N_16478);
or U23051 (N_23051,N_16643,N_16362);
nor U23052 (N_23052,N_17478,N_17961);
nand U23053 (N_23053,N_12170,N_17036);
xnor U23054 (N_23054,N_16136,N_12015);
or U23055 (N_23055,N_12180,N_16533);
and U23056 (N_23056,N_16992,N_12216);
or U23057 (N_23057,N_14046,N_15898);
or U23058 (N_23058,N_17231,N_16616);
and U23059 (N_23059,N_12148,N_13363);
nor U23060 (N_23060,N_13308,N_14584);
nand U23061 (N_23061,N_13351,N_16222);
or U23062 (N_23062,N_16469,N_17529);
nand U23063 (N_23063,N_16438,N_15195);
xor U23064 (N_23064,N_16897,N_16657);
nand U23065 (N_23065,N_14231,N_14412);
nor U23066 (N_23066,N_13679,N_17856);
or U23067 (N_23067,N_13080,N_14957);
or U23068 (N_23068,N_16315,N_15843);
xnor U23069 (N_23069,N_14605,N_12344);
nor U23070 (N_23070,N_17323,N_13669);
and U23071 (N_23071,N_16297,N_14745);
or U23072 (N_23072,N_16100,N_16103);
nor U23073 (N_23073,N_16827,N_15171);
and U23074 (N_23074,N_12605,N_17874);
nand U23075 (N_23075,N_13933,N_17917);
nor U23076 (N_23076,N_16183,N_16576);
xnor U23077 (N_23077,N_14962,N_15964);
and U23078 (N_23078,N_17193,N_14616);
xor U23079 (N_23079,N_13396,N_15552);
or U23080 (N_23080,N_12738,N_15669);
and U23081 (N_23081,N_13334,N_16338);
nor U23082 (N_23082,N_13238,N_17081);
or U23083 (N_23083,N_17884,N_17536);
nand U23084 (N_23084,N_15670,N_14796);
nor U23085 (N_23085,N_15908,N_12019);
or U23086 (N_23086,N_12204,N_17267);
and U23087 (N_23087,N_17501,N_15723);
nand U23088 (N_23088,N_15831,N_14182);
or U23089 (N_23089,N_14198,N_12930);
or U23090 (N_23090,N_12104,N_16028);
or U23091 (N_23091,N_14566,N_12627);
xor U23092 (N_23092,N_12079,N_16230);
nor U23093 (N_23093,N_15671,N_13858);
xor U23094 (N_23094,N_12570,N_12232);
and U23095 (N_23095,N_14888,N_14773);
nor U23096 (N_23096,N_17556,N_13744);
or U23097 (N_23097,N_17202,N_12340);
nor U23098 (N_23098,N_15825,N_14621);
nor U23099 (N_23099,N_15034,N_13436);
nand U23100 (N_23100,N_12797,N_17453);
or U23101 (N_23101,N_16990,N_16456);
nor U23102 (N_23102,N_17575,N_17602);
or U23103 (N_23103,N_15000,N_16016);
nor U23104 (N_23104,N_13900,N_12269);
and U23105 (N_23105,N_17289,N_12522);
and U23106 (N_23106,N_17871,N_14477);
nand U23107 (N_23107,N_15088,N_14496);
and U23108 (N_23108,N_14838,N_17570);
and U23109 (N_23109,N_15758,N_17316);
xor U23110 (N_23110,N_12168,N_12568);
nand U23111 (N_23111,N_13750,N_13385);
nand U23112 (N_23112,N_15908,N_15366);
nor U23113 (N_23113,N_16864,N_12114);
nor U23114 (N_23114,N_15954,N_15551);
nand U23115 (N_23115,N_13534,N_14327);
and U23116 (N_23116,N_12510,N_14742);
or U23117 (N_23117,N_12173,N_15796);
or U23118 (N_23118,N_15885,N_12003);
nor U23119 (N_23119,N_15406,N_14275);
nand U23120 (N_23120,N_16192,N_14180);
xnor U23121 (N_23121,N_14818,N_14944);
and U23122 (N_23122,N_13829,N_17478);
and U23123 (N_23123,N_15707,N_16615);
or U23124 (N_23124,N_15706,N_12200);
and U23125 (N_23125,N_15592,N_16711);
and U23126 (N_23126,N_12013,N_16377);
nand U23127 (N_23127,N_13001,N_14340);
and U23128 (N_23128,N_12999,N_16161);
or U23129 (N_23129,N_17104,N_15045);
nor U23130 (N_23130,N_15457,N_15014);
or U23131 (N_23131,N_12941,N_14038);
xor U23132 (N_23132,N_13272,N_17954);
or U23133 (N_23133,N_12452,N_16291);
nand U23134 (N_23134,N_17737,N_12364);
and U23135 (N_23135,N_14316,N_16360);
nand U23136 (N_23136,N_13502,N_16996);
nand U23137 (N_23137,N_12694,N_15243);
xor U23138 (N_23138,N_14787,N_16200);
and U23139 (N_23139,N_15229,N_13448);
nand U23140 (N_23140,N_16151,N_14630);
nor U23141 (N_23141,N_15514,N_14386);
nand U23142 (N_23142,N_14078,N_16455);
or U23143 (N_23143,N_14216,N_16592);
and U23144 (N_23144,N_15554,N_13449);
xor U23145 (N_23145,N_16045,N_14220);
and U23146 (N_23146,N_17559,N_15531);
xor U23147 (N_23147,N_12002,N_16726);
and U23148 (N_23148,N_16167,N_15790);
or U23149 (N_23149,N_13081,N_13360);
nor U23150 (N_23150,N_14092,N_17518);
and U23151 (N_23151,N_14344,N_12564);
xnor U23152 (N_23152,N_15211,N_13055);
nand U23153 (N_23153,N_12411,N_15121);
xor U23154 (N_23154,N_16032,N_14671);
and U23155 (N_23155,N_15724,N_14459);
and U23156 (N_23156,N_17778,N_17767);
nor U23157 (N_23157,N_14091,N_14191);
or U23158 (N_23158,N_15891,N_15312);
or U23159 (N_23159,N_13785,N_12876);
xnor U23160 (N_23160,N_12120,N_14544);
xnor U23161 (N_23161,N_15886,N_15485);
nor U23162 (N_23162,N_15611,N_14812);
and U23163 (N_23163,N_14872,N_12544);
nand U23164 (N_23164,N_17418,N_13329);
nor U23165 (N_23165,N_15426,N_12876);
and U23166 (N_23166,N_13487,N_15426);
nor U23167 (N_23167,N_12505,N_14127);
nand U23168 (N_23168,N_13865,N_12728);
or U23169 (N_23169,N_14036,N_13299);
and U23170 (N_23170,N_12656,N_12690);
or U23171 (N_23171,N_12054,N_15230);
nor U23172 (N_23172,N_15176,N_12157);
nor U23173 (N_23173,N_15290,N_16291);
or U23174 (N_23174,N_15728,N_14005);
and U23175 (N_23175,N_13649,N_17535);
or U23176 (N_23176,N_17228,N_12532);
and U23177 (N_23177,N_13863,N_14387);
and U23178 (N_23178,N_16647,N_17413);
nor U23179 (N_23179,N_17590,N_17606);
and U23180 (N_23180,N_16379,N_17110);
nand U23181 (N_23181,N_14599,N_17761);
nor U23182 (N_23182,N_14200,N_12357);
and U23183 (N_23183,N_13025,N_15615);
and U23184 (N_23184,N_14017,N_13155);
or U23185 (N_23185,N_14617,N_12083);
nor U23186 (N_23186,N_14034,N_12667);
nand U23187 (N_23187,N_16367,N_12424);
nor U23188 (N_23188,N_12056,N_16953);
nand U23189 (N_23189,N_15999,N_14889);
nor U23190 (N_23190,N_15887,N_14776);
or U23191 (N_23191,N_17128,N_15102);
nor U23192 (N_23192,N_12304,N_14774);
or U23193 (N_23193,N_13725,N_14631);
xnor U23194 (N_23194,N_15617,N_12868);
xor U23195 (N_23195,N_16055,N_16667);
nand U23196 (N_23196,N_17878,N_13081);
or U23197 (N_23197,N_12041,N_17065);
or U23198 (N_23198,N_17453,N_13537);
xnor U23199 (N_23199,N_12912,N_16604);
or U23200 (N_23200,N_15735,N_16687);
nand U23201 (N_23201,N_14812,N_16630);
nand U23202 (N_23202,N_16199,N_13055);
and U23203 (N_23203,N_12757,N_15024);
and U23204 (N_23204,N_12036,N_17871);
or U23205 (N_23205,N_13397,N_16494);
nand U23206 (N_23206,N_15475,N_15397);
and U23207 (N_23207,N_12100,N_13799);
nand U23208 (N_23208,N_13852,N_13585);
or U23209 (N_23209,N_15120,N_12570);
nor U23210 (N_23210,N_13737,N_16523);
or U23211 (N_23211,N_14139,N_12560);
nor U23212 (N_23212,N_14921,N_17294);
xnor U23213 (N_23213,N_13584,N_13659);
and U23214 (N_23214,N_16464,N_14128);
and U23215 (N_23215,N_15004,N_14779);
nand U23216 (N_23216,N_16011,N_13166);
and U23217 (N_23217,N_14707,N_12261);
nor U23218 (N_23218,N_13265,N_16389);
nand U23219 (N_23219,N_16283,N_16430);
nand U23220 (N_23220,N_13298,N_13864);
nand U23221 (N_23221,N_12770,N_15388);
and U23222 (N_23222,N_12520,N_12603);
nand U23223 (N_23223,N_13489,N_13011);
and U23224 (N_23224,N_15708,N_16584);
nand U23225 (N_23225,N_16967,N_12108);
or U23226 (N_23226,N_16429,N_13118);
and U23227 (N_23227,N_13444,N_15578);
xor U23228 (N_23228,N_13622,N_15202);
or U23229 (N_23229,N_14268,N_16283);
and U23230 (N_23230,N_16337,N_12301);
and U23231 (N_23231,N_13237,N_14809);
xor U23232 (N_23232,N_14164,N_14428);
and U23233 (N_23233,N_17244,N_16978);
nor U23234 (N_23234,N_14875,N_17363);
or U23235 (N_23235,N_15357,N_17759);
nor U23236 (N_23236,N_13479,N_15093);
and U23237 (N_23237,N_12667,N_13607);
or U23238 (N_23238,N_14490,N_13231);
and U23239 (N_23239,N_15079,N_17214);
nor U23240 (N_23240,N_15752,N_15161);
and U23241 (N_23241,N_17092,N_12909);
nand U23242 (N_23242,N_12554,N_15668);
xor U23243 (N_23243,N_16883,N_16014);
nand U23244 (N_23244,N_14257,N_12241);
or U23245 (N_23245,N_12141,N_17185);
or U23246 (N_23246,N_13659,N_13376);
and U23247 (N_23247,N_17724,N_15796);
or U23248 (N_23248,N_14718,N_12884);
xor U23249 (N_23249,N_12168,N_13012);
and U23250 (N_23250,N_13879,N_17166);
or U23251 (N_23251,N_13235,N_12639);
nand U23252 (N_23252,N_14459,N_17202);
and U23253 (N_23253,N_13278,N_13368);
and U23254 (N_23254,N_16941,N_15455);
and U23255 (N_23255,N_17737,N_17428);
xor U23256 (N_23256,N_15071,N_13443);
nand U23257 (N_23257,N_13039,N_16027);
nor U23258 (N_23258,N_16821,N_17349);
nand U23259 (N_23259,N_14324,N_15857);
nand U23260 (N_23260,N_14846,N_16671);
and U23261 (N_23261,N_17750,N_12127);
nor U23262 (N_23262,N_13825,N_14048);
nor U23263 (N_23263,N_12182,N_15676);
nand U23264 (N_23264,N_12778,N_14298);
and U23265 (N_23265,N_14747,N_16706);
or U23266 (N_23266,N_13822,N_14125);
or U23267 (N_23267,N_14784,N_12033);
or U23268 (N_23268,N_15225,N_16155);
or U23269 (N_23269,N_17061,N_17786);
xor U23270 (N_23270,N_12485,N_14906);
nand U23271 (N_23271,N_17738,N_15012);
nor U23272 (N_23272,N_17707,N_14528);
and U23273 (N_23273,N_14025,N_13880);
or U23274 (N_23274,N_15967,N_17728);
or U23275 (N_23275,N_13106,N_16682);
nor U23276 (N_23276,N_12918,N_16597);
nor U23277 (N_23277,N_14387,N_13582);
or U23278 (N_23278,N_14943,N_13889);
nor U23279 (N_23279,N_16046,N_17588);
nor U23280 (N_23280,N_12742,N_16677);
and U23281 (N_23281,N_14016,N_13191);
nand U23282 (N_23282,N_15640,N_17262);
nand U23283 (N_23283,N_16007,N_15468);
and U23284 (N_23284,N_13165,N_15474);
and U23285 (N_23285,N_16773,N_13158);
and U23286 (N_23286,N_16004,N_15184);
and U23287 (N_23287,N_15397,N_17837);
or U23288 (N_23288,N_16825,N_17643);
or U23289 (N_23289,N_13547,N_16280);
nand U23290 (N_23290,N_16713,N_16611);
nor U23291 (N_23291,N_13882,N_15923);
and U23292 (N_23292,N_14159,N_15862);
or U23293 (N_23293,N_12078,N_12937);
or U23294 (N_23294,N_12261,N_17423);
xor U23295 (N_23295,N_17720,N_16769);
or U23296 (N_23296,N_17205,N_17887);
nor U23297 (N_23297,N_15875,N_17733);
and U23298 (N_23298,N_12891,N_13503);
xnor U23299 (N_23299,N_13603,N_13335);
nor U23300 (N_23300,N_17982,N_16539);
nand U23301 (N_23301,N_13131,N_13888);
xor U23302 (N_23302,N_12884,N_13737);
and U23303 (N_23303,N_17984,N_17085);
or U23304 (N_23304,N_14350,N_16702);
nor U23305 (N_23305,N_14455,N_15457);
xnor U23306 (N_23306,N_17626,N_17816);
nor U23307 (N_23307,N_12661,N_13255);
or U23308 (N_23308,N_17601,N_12113);
and U23309 (N_23309,N_13864,N_16934);
nor U23310 (N_23310,N_15212,N_17672);
and U23311 (N_23311,N_12549,N_16862);
nand U23312 (N_23312,N_17496,N_14553);
or U23313 (N_23313,N_16610,N_17275);
or U23314 (N_23314,N_13279,N_15983);
nor U23315 (N_23315,N_16633,N_12403);
nor U23316 (N_23316,N_13418,N_15109);
nand U23317 (N_23317,N_14588,N_14698);
nor U23318 (N_23318,N_16452,N_12942);
and U23319 (N_23319,N_12458,N_13147);
nor U23320 (N_23320,N_14708,N_14868);
nor U23321 (N_23321,N_12401,N_13252);
xor U23322 (N_23322,N_14408,N_13700);
nor U23323 (N_23323,N_12693,N_13309);
or U23324 (N_23324,N_12142,N_13321);
and U23325 (N_23325,N_17167,N_14500);
xnor U23326 (N_23326,N_15074,N_13639);
or U23327 (N_23327,N_17985,N_15321);
xnor U23328 (N_23328,N_12392,N_16953);
and U23329 (N_23329,N_15763,N_16373);
and U23330 (N_23330,N_17520,N_16397);
and U23331 (N_23331,N_13065,N_17529);
nor U23332 (N_23332,N_12014,N_17769);
nand U23333 (N_23333,N_14421,N_17180);
xor U23334 (N_23334,N_16023,N_17371);
or U23335 (N_23335,N_13767,N_12007);
and U23336 (N_23336,N_13874,N_13789);
and U23337 (N_23337,N_15513,N_13251);
nor U23338 (N_23338,N_14588,N_16756);
nand U23339 (N_23339,N_14082,N_17691);
or U23340 (N_23340,N_17546,N_16816);
nand U23341 (N_23341,N_14694,N_17067);
nand U23342 (N_23342,N_12441,N_15236);
or U23343 (N_23343,N_14925,N_13174);
nor U23344 (N_23344,N_15422,N_16099);
nor U23345 (N_23345,N_14826,N_12101);
or U23346 (N_23346,N_12234,N_14390);
nor U23347 (N_23347,N_16228,N_13752);
nor U23348 (N_23348,N_16892,N_15064);
and U23349 (N_23349,N_16039,N_16291);
and U23350 (N_23350,N_13800,N_15785);
nor U23351 (N_23351,N_15657,N_15208);
nor U23352 (N_23352,N_16194,N_17530);
or U23353 (N_23353,N_14878,N_15228);
nand U23354 (N_23354,N_17026,N_17743);
nor U23355 (N_23355,N_17339,N_16615);
or U23356 (N_23356,N_14623,N_13334);
nor U23357 (N_23357,N_12423,N_16702);
or U23358 (N_23358,N_12911,N_13611);
nor U23359 (N_23359,N_16404,N_14334);
or U23360 (N_23360,N_13266,N_17348);
and U23361 (N_23361,N_14802,N_17196);
nand U23362 (N_23362,N_14175,N_14283);
xor U23363 (N_23363,N_17830,N_16771);
or U23364 (N_23364,N_14188,N_13130);
xor U23365 (N_23365,N_13741,N_14410);
or U23366 (N_23366,N_13121,N_12089);
nor U23367 (N_23367,N_15793,N_15382);
nand U23368 (N_23368,N_16074,N_13178);
nand U23369 (N_23369,N_16863,N_17896);
nand U23370 (N_23370,N_12972,N_12360);
nor U23371 (N_23371,N_17575,N_12665);
nor U23372 (N_23372,N_13111,N_15383);
or U23373 (N_23373,N_17771,N_16929);
nor U23374 (N_23374,N_12632,N_14524);
nor U23375 (N_23375,N_13040,N_16571);
and U23376 (N_23376,N_16567,N_12652);
nor U23377 (N_23377,N_12518,N_12052);
nand U23378 (N_23378,N_13441,N_14850);
xor U23379 (N_23379,N_14978,N_16398);
nor U23380 (N_23380,N_16900,N_17390);
or U23381 (N_23381,N_12483,N_15322);
nor U23382 (N_23382,N_15604,N_16187);
nor U23383 (N_23383,N_17438,N_17535);
or U23384 (N_23384,N_16881,N_13049);
nor U23385 (N_23385,N_12058,N_14301);
nand U23386 (N_23386,N_12197,N_14861);
or U23387 (N_23387,N_16893,N_15118);
nand U23388 (N_23388,N_15855,N_13805);
or U23389 (N_23389,N_15618,N_14568);
nor U23390 (N_23390,N_13717,N_12055);
nor U23391 (N_23391,N_12960,N_15437);
or U23392 (N_23392,N_14497,N_15227);
and U23393 (N_23393,N_13025,N_16045);
nand U23394 (N_23394,N_14366,N_14959);
or U23395 (N_23395,N_14646,N_12743);
or U23396 (N_23396,N_16677,N_14652);
xnor U23397 (N_23397,N_15978,N_16400);
and U23398 (N_23398,N_15592,N_16431);
and U23399 (N_23399,N_17710,N_14313);
and U23400 (N_23400,N_14450,N_13861);
nor U23401 (N_23401,N_16291,N_15973);
nor U23402 (N_23402,N_14206,N_15556);
nand U23403 (N_23403,N_17818,N_16987);
or U23404 (N_23404,N_14455,N_14365);
or U23405 (N_23405,N_12722,N_16687);
and U23406 (N_23406,N_13507,N_14123);
and U23407 (N_23407,N_14167,N_14820);
xnor U23408 (N_23408,N_14634,N_14560);
nand U23409 (N_23409,N_13928,N_14165);
nand U23410 (N_23410,N_14959,N_14659);
xnor U23411 (N_23411,N_12149,N_12266);
and U23412 (N_23412,N_17851,N_16429);
nor U23413 (N_23413,N_12110,N_14416);
or U23414 (N_23414,N_17095,N_16186);
nor U23415 (N_23415,N_13101,N_12824);
xnor U23416 (N_23416,N_13303,N_16917);
nor U23417 (N_23417,N_17794,N_17322);
and U23418 (N_23418,N_12685,N_13835);
nand U23419 (N_23419,N_17839,N_14012);
nand U23420 (N_23420,N_12597,N_12418);
or U23421 (N_23421,N_13962,N_12594);
and U23422 (N_23422,N_15796,N_13264);
and U23423 (N_23423,N_16246,N_15901);
nor U23424 (N_23424,N_15487,N_17610);
or U23425 (N_23425,N_15542,N_16189);
and U23426 (N_23426,N_14283,N_13917);
nand U23427 (N_23427,N_14835,N_14885);
and U23428 (N_23428,N_13147,N_17153);
and U23429 (N_23429,N_16532,N_16981);
nand U23430 (N_23430,N_14966,N_17114);
nand U23431 (N_23431,N_14706,N_17472);
or U23432 (N_23432,N_16870,N_16487);
xnor U23433 (N_23433,N_16301,N_13973);
and U23434 (N_23434,N_13358,N_13227);
and U23435 (N_23435,N_15482,N_14134);
nor U23436 (N_23436,N_17229,N_12743);
and U23437 (N_23437,N_13029,N_17812);
xor U23438 (N_23438,N_13139,N_14171);
and U23439 (N_23439,N_12238,N_13531);
or U23440 (N_23440,N_14188,N_17095);
nor U23441 (N_23441,N_14884,N_13938);
nand U23442 (N_23442,N_15863,N_16181);
and U23443 (N_23443,N_12200,N_12192);
or U23444 (N_23444,N_12890,N_13819);
and U23445 (N_23445,N_12914,N_12508);
or U23446 (N_23446,N_13833,N_12840);
or U23447 (N_23447,N_12495,N_15187);
and U23448 (N_23448,N_15409,N_13729);
and U23449 (N_23449,N_15927,N_17171);
or U23450 (N_23450,N_14689,N_13527);
xnor U23451 (N_23451,N_17679,N_14251);
nor U23452 (N_23452,N_15820,N_16999);
nor U23453 (N_23453,N_12681,N_14718);
xor U23454 (N_23454,N_16457,N_14116);
nor U23455 (N_23455,N_13945,N_14785);
and U23456 (N_23456,N_17413,N_13685);
and U23457 (N_23457,N_17653,N_13817);
nand U23458 (N_23458,N_17531,N_12198);
or U23459 (N_23459,N_14174,N_12873);
nor U23460 (N_23460,N_17502,N_14653);
nand U23461 (N_23461,N_14757,N_14514);
and U23462 (N_23462,N_16499,N_16665);
and U23463 (N_23463,N_12706,N_12917);
nand U23464 (N_23464,N_16905,N_16535);
and U23465 (N_23465,N_12429,N_16591);
or U23466 (N_23466,N_16921,N_15949);
and U23467 (N_23467,N_15076,N_14295);
xor U23468 (N_23468,N_16462,N_14576);
nand U23469 (N_23469,N_15820,N_15548);
nand U23470 (N_23470,N_16709,N_13025);
or U23471 (N_23471,N_14940,N_17796);
nor U23472 (N_23472,N_17800,N_16882);
xor U23473 (N_23473,N_16116,N_16676);
and U23474 (N_23474,N_16773,N_13916);
nand U23475 (N_23475,N_13001,N_13569);
or U23476 (N_23476,N_13129,N_16509);
and U23477 (N_23477,N_16327,N_14780);
and U23478 (N_23478,N_13775,N_17485);
and U23479 (N_23479,N_13674,N_16324);
or U23480 (N_23480,N_17760,N_14607);
and U23481 (N_23481,N_17577,N_17804);
nand U23482 (N_23482,N_15568,N_15719);
xor U23483 (N_23483,N_15068,N_14725);
and U23484 (N_23484,N_14636,N_15503);
or U23485 (N_23485,N_17987,N_17650);
xor U23486 (N_23486,N_12014,N_12135);
nand U23487 (N_23487,N_17571,N_12915);
or U23488 (N_23488,N_12439,N_12476);
or U23489 (N_23489,N_15847,N_17832);
nand U23490 (N_23490,N_17526,N_16733);
nor U23491 (N_23491,N_12181,N_16868);
or U23492 (N_23492,N_14245,N_14756);
nor U23493 (N_23493,N_16635,N_14718);
nor U23494 (N_23494,N_13131,N_13756);
nand U23495 (N_23495,N_17991,N_17875);
nor U23496 (N_23496,N_15095,N_16296);
and U23497 (N_23497,N_12850,N_17158);
and U23498 (N_23498,N_15555,N_15406);
nand U23499 (N_23499,N_13228,N_15987);
nor U23500 (N_23500,N_13972,N_14053);
nand U23501 (N_23501,N_16840,N_12040);
or U23502 (N_23502,N_12440,N_17920);
or U23503 (N_23503,N_17710,N_12444);
nand U23504 (N_23504,N_14436,N_13893);
and U23505 (N_23505,N_14131,N_16909);
or U23506 (N_23506,N_17830,N_15638);
and U23507 (N_23507,N_15513,N_14007);
nand U23508 (N_23508,N_17338,N_14459);
nand U23509 (N_23509,N_14359,N_16996);
and U23510 (N_23510,N_15540,N_15369);
xnor U23511 (N_23511,N_13696,N_13776);
nor U23512 (N_23512,N_12997,N_14590);
or U23513 (N_23513,N_15108,N_16092);
and U23514 (N_23514,N_17719,N_14205);
and U23515 (N_23515,N_17118,N_17614);
or U23516 (N_23516,N_15068,N_14218);
and U23517 (N_23517,N_15476,N_15715);
nand U23518 (N_23518,N_14295,N_13871);
and U23519 (N_23519,N_17639,N_17193);
nor U23520 (N_23520,N_13937,N_17152);
nor U23521 (N_23521,N_17167,N_14645);
and U23522 (N_23522,N_16123,N_16768);
or U23523 (N_23523,N_14729,N_12221);
nor U23524 (N_23524,N_15152,N_13508);
nor U23525 (N_23525,N_13651,N_13326);
nand U23526 (N_23526,N_14885,N_14061);
nor U23527 (N_23527,N_12282,N_13597);
or U23528 (N_23528,N_16126,N_14819);
and U23529 (N_23529,N_15773,N_17822);
xnor U23530 (N_23530,N_12867,N_16227);
and U23531 (N_23531,N_12587,N_15502);
and U23532 (N_23532,N_17683,N_15717);
nand U23533 (N_23533,N_12300,N_16367);
nor U23534 (N_23534,N_14430,N_12157);
nor U23535 (N_23535,N_12501,N_13488);
or U23536 (N_23536,N_16313,N_17706);
xnor U23537 (N_23537,N_15715,N_16064);
nor U23538 (N_23538,N_12300,N_17581);
nand U23539 (N_23539,N_17456,N_12440);
or U23540 (N_23540,N_13688,N_12090);
nor U23541 (N_23541,N_15886,N_16482);
nand U23542 (N_23542,N_15601,N_13935);
nor U23543 (N_23543,N_13709,N_17448);
nor U23544 (N_23544,N_12958,N_17927);
nand U23545 (N_23545,N_12435,N_13575);
xor U23546 (N_23546,N_12444,N_14007);
and U23547 (N_23547,N_14093,N_16625);
and U23548 (N_23548,N_12874,N_15114);
and U23549 (N_23549,N_16048,N_16110);
nand U23550 (N_23550,N_15211,N_15180);
and U23551 (N_23551,N_17419,N_14812);
nand U23552 (N_23552,N_12976,N_16223);
nor U23553 (N_23553,N_16056,N_15848);
nand U23554 (N_23554,N_14410,N_15150);
and U23555 (N_23555,N_17719,N_16365);
and U23556 (N_23556,N_15144,N_17483);
nand U23557 (N_23557,N_16807,N_16865);
nor U23558 (N_23558,N_12104,N_15503);
nor U23559 (N_23559,N_12839,N_15013);
or U23560 (N_23560,N_14035,N_13426);
and U23561 (N_23561,N_15405,N_16371);
and U23562 (N_23562,N_13429,N_13009);
and U23563 (N_23563,N_16669,N_14843);
and U23564 (N_23564,N_14922,N_16839);
nor U23565 (N_23565,N_12947,N_16912);
and U23566 (N_23566,N_15175,N_16327);
nand U23567 (N_23567,N_15333,N_12548);
nor U23568 (N_23568,N_17140,N_15518);
nor U23569 (N_23569,N_14332,N_17236);
nor U23570 (N_23570,N_14845,N_15891);
and U23571 (N_23571,N_16133,N_16763);
nand U23572 (N_23572,N_12295,N_14560);
nand U23573 (N_23573,N_16818,N_16028);
nor U23574 (N_23574,N_12610,N_12240);
and U23575 (N_23575,N_12532,N_14313);
or U23576 (N_23576,N_14887,N_16457);
nand U23577 (N_23577,N_15082,N_16926);
and U23578 (N_23578,N_16658,N_12885);
and U23579 (N_23579,N_13487,N_15016);
nand U23580 (N_23580,N_12176,N_13376);
or U23581 (N_23581,N_17840,N_14447);
nor U23582 (N_23582,N_17543,N_13571);
or U23583 (N_23583,N_14294,N_16266);
nor U23584 (N_23584,N_16891,N_13553);
nand U23585 (N_23585,N_13911,N_16352);
or U23586 (N_23586,N_14401,N_16149);
or U23587 (N_23587,N_14220,N_17155);
and U23588 (N_23588,N_17751,N_13858);
nand U23589 (N_23589,N_15252,N_17411);
or U23590 (N_23590,N_12496,N_15573);
nand U23591 (N_23591,N_17758,N_16038);
or U23592 (N_23592,N_13078,N_14633);
or U23593 (N_23593,N_17546,N_16949);
or U23594 (N_23594,N_16284,N_12884);
or U23595 (N_23595,N_14536,N_16161);
and U23596 (N_23596,N_14131,N_16378);
nand U23597 (N_23597,N_14808,N_14316);
xnor U23598 (N_23598,N_13285,N_16207);
and U23599 (N_23599,N_14760,N_12281);
or U23600 (N_23600,N_15343,N_14716);
or U23601 (N_23601,N_17638,N_13698);
nand U23602 (N_23602,N_12246,N_13792);
xor U23603 (N_23603,N_17857,N_13354);
nand U23604 (N_23604,N_17153,N_13128);
xor U23605 (N_23605,N_15979,N_16890);
and U23606 (N_23606,N_17571,N_14354);
nor U23607 (N_23607,N_16684,N_12867);
or U23608 (N_23608,N_14460,N_17985);
and U23609 (N_23609,N_12164,N_14562);
and U23610 (N_23610,N_17580,N_14855);
nor U23611 (N_23611,N_17293,N_15963);
or U23612 (N_23612,N_16872,N_16315);
nand U23613 (N_23613,N_13497,N_14197);
nor U23614 (N_23614,N_16096,N_17948);
xnor U23615 (N_23615,N_14588,N_15962);
and U23616 (N_23616,N_12635,N_15337);
nand U23617 (N_23617,N_14582,N_12963);
and U23618 (N_23618,N_12294,N_12385);
nand U23619 (N_23619,N_14604,N_17876);
nor U23620 (N_23620,N_14515,N_13704);
nor U23621 (N_23621,N_16304,N_14789);
nand U23622 (N_23622,N_13711,N_17825);
or U23623 (N_23623,N_17226,N_17720);
or U23624 (N_23624,N_15914,N_13817);
nand U23625 (N_23625,N_13358,N_13657);
nand U23626 (N_23626,N_12407,N_16387);
nor U23627 (N_23627,N_14489,N_15267);
or U23628 (N_23628,N_17693,N_16453);
nor U23629 (N_23629,N_12750,N_13238);
or U23630 (N_23630,N_15780,N_16750);
or U23631 (N_23631,N_12153,N_14698);
or U23632 (N_23632,N_16161,N_14517);
or U23633 (N_23633,N_12221,N_14194);
and U23634 (N_23634,N_15512,N_14315);
and U23635 (N_23635,N_15895,N_14495);
nor U23636 (N_23636,N_12540,N_12139);
nor U23637 (N_23637,N_17095,N_12044);
and U23638 (N_23638,N_15329,N_17631);
or U23639 (N_23639,N_15682,N_16181);
nand U23640 (N_23640,N_14183,N_15350);
and U23641 (N_23641,N_14847,N_16181);
and U23642 (N_23642,N_14162,N_14981);
or U23643 (N_23643,N_16188,N_16775);
nor U23644 (N_23644,N_12197,N_13858);
or U23645 (N_23645,N_14003,N_16172);
nand U23646 (N_23646,N_12726,N_13697);
or U23647 (N_23647,N_13138,N_15243);
nand U23648 (N_23648,N_16442,N_12387);
nor U23649 (N_23649,N_13597,N_15774);
and U23650 (N_23650,N_15370,N_14985);
or U23651 (N_23651,N_13198,N_13834);
and U23652 (N_23652,N_12933,N_16849);
or U23653 (N_23653,N_17580,N_16993);
nor U23654 (N_23654,N_13309,N_16775);
nand U23655 (N_23655,N_16633,N_16281);
nor U23656 (N_23656,N_12960,N_13677);
and U23657 (N_23657,N_16361,N_12101);
and U23658 (N_23658,N_17199,N_17106);
nand U23659 (N_23659,N_12325,N_17089);
nand U23660 (N_23660,N_14231,N_14415);
nor U23661 (N_23661,N_16844,N_14771);
xor U23662 (N_23662,N_12135,N_16646);
nand U23663 (N_23663,N_13569,N_12707);
nor U23664 (N_23664,N_14639,N_17050);
xor U23665 (N_23665,N_17081,N_15511);
or U23666 (N_23666,N_16243,N_17464);
and U23667 (N_23667,N_14488,N_14934);
or U23668 (N_23668,N_15253,N_12946);
nand U23669 (N_23669,N_12026,N_13116);
nor U23670 (N_23670,N_16937,N_14127);
and U23671 (N_23671,N_16549,N_16509);
or U23672 (N_23672,N_12820,N_14768);
and U23673 (N_23673,N_17197,N_16816);
xnor U23674 (N_23674,N_12199,N_13063);
xor U23675 (N_23675,N_13436,N_14247);
or U23676 (N_23676,N_16778,N_13409);
and U23677 (N_23677,N_14328,N_14613);
nor U23678 (N_23678,N_17122,N_13112);
nand U23679 (N_23679,N_15219,N_16023);
nor U23680 (N_23680,N_14751,N_15207);
nand U23681 (N_23681,N_13488,N_14405);
and U23682 (N_23682,N_12523,N_16790);
xnor U23683 (N_23683,N_14059,N_12564);
or U23684 (N_23684,N_14149,N_13486);
and U23685 (N_23685,N_16293,N_13634);
nor U23686 (N_23686,N_16761,N_15621);
or U23687 (N_23687,N_14800,N_17258);
xor U23688 (N_23688,N_17268,N_15938);
and U23689 (N_23689,N_12727,N_13129);
nor U23690 (N_23690,N_13615,N_16470);
nor U23691 (N_23691,N_15399,N_14600);
nor U23692 (N_23692,N_13935,N_16432);
and U23693 (N_23693,N_14464,N_16062);
nor U23694 (N_23694,N_12048,N_15652);
and U23695 (N_23695,N_16321,N_14610);
nor U23696 (N_23696,N_12481,N_14096);
nand U23697 (N_23697,N_14363,N_12604);
or U23698 (N_23698,N_16179,N_14640);
nor U23699 (N_23699,N_15024,N_12327);
and U23700 (N_23700,N_15143,N_14604);
and U23701 (N_23701,N_17032,N_17600);
nand U23702 (N_23702,N_12099,N_12149);
nor U23703 (N_23703,N_17903,N_12247);
xor U23704 (N_23704,N_14418,N_13842);
nand U23705 (N_23705,N_12222,N_14742);
and U23706 (N_23706,N_15172,N_16621);
or U23707 (N_23707,N_17917,N_13364);
or U23708 (N_23708,N_17412,N_12816);
or U23709 (N_23709,N_17826,N_13838);
xor U23710 (N_23710,N_14720,N_15291);
and U23711 (N_23711,N_17542,N_15591);
or U23712 (N_23712,N_17463,N_13606);
nand U23713 (N_23713,N_13295,N_12013);
and U23714 (N_23714,N_15501,N_16059);
nand U23715 (N_23715,N_15300,N_17007);
or U23716 (N_23716,N_12005,N_15801);
and U23717 (N_23717,N_15724,N_13669);
or U23718 (N_23718,N_17202,N_13799);
nor U23719 (N_23719,N_15034,N_12175);
nand U23720 (N_23720,N_16716,N_17485);
xnor U23721 (N_23721,N_12757,N_15858);
nand U23722 (N_23722,N_13390,N_17160);
nor U23723 (N_23723,N_13045,N_13766);
and U23724 (N_23724,N_13770,N_15449);
and U23725 (N_23725,N_15849,N_17238);
xor U23726 (N_23726,N_12000,N_17217);
and U23727 (N_23727,N_17377,N_13937);
nor U23728 (N_23728,N_15387,N_17713);
nand U23729 (N_23729,N_17011,N_16165);
xor U23730 (N_23730,N_14333,N_17234);
and U23731 (N_23731,N_13045,N_14278);
xor U23732 (N_23732,N_12377,N_14353);
or U23733 (N_23733,N_17312,N_16696);
nand U23734 (N_23734,N_16444,N_16350);
or U23735 (N_23735,N_16153,N_14080);
nor U23736 (N_23736,N_17699,N_15195);
nand U23737 (N_23737,N_17381,N_16491);
nor U23738 (N_23738,N_14616,N_13681);
or U23739 (N_23739,N_14067,N_15861);
nor U23740 (N_23740,N_16224,N_13012);
xor U23741 (N_23741,N_16743,N_15727);
or U23742 (N_23742,N_13128,N_17434);
and U23743 (N_23743,N_12395,N_16289);
or U23744 (N_23744,N_17231,N_12683);
nor U23745 (N_23745,N_12015,N_12918);
xnor U23746 (N_23746,N_13574,N_17744);
xor U23747 (N_23747,N_12171,N_16030);
or U23748 (N_23748,N_14259,N_15253);
and U23749 (N_23749,N_12080,N_14757);
or U23750 (N_23750,N_16211,N_12533);
nor U23751 (N_23751,N_17870,N_16982);
nand U23752 (N_23752,N_16830,N_12467);
nor U23753 (N_23753,N_15759,N_17497);
or U23754 (N_23754,N_12657,N_17679);
or U23755 (N_23755,N_12363,N_17408);
nand U23756 (N_23756,N_13452,N_13216);
or U23757 (N_23757,N_12572,N_16415);
or U23758 (N_23758,N_15038,N_13187);
nand U23759 (N_23759,N_17456,N_12352);
nor U23760 (N_23760,N_17872,N_13288);
nor U23761 (N_23761,N_13945,N_17606);
nor U23762 (N_23762,N_14852,N_14790);
or U23763 (N_23763,N_17148,N_16398);
xor U23764 (N_23764,N_15287,N_16839);
and U23765 (N_23765,N_17129,N_12493);
and U23766 (N_23766,N_13342,N_16810);
xor U23767 (N_23767,N_15091,N_16225);
nand U23768 (N_23768,N_14698,N_15669);
or U23769 (N_23769,N_17191,N_15955);
nor U23770 (N_23770,N_16307,N_14500);
nand U23771 (N_23771,N_17253,N_16052);
nor U23772 (N_23772,N_16217,N_14838);
or U23773 (N_23773,N_17917,N_17673);
and U23774 (N_23774,N_16794,N_14624);
and U23775 (N_23775,N_13033,N_14126);
nand U23776 (N_23776,N_13207,N_17337);
nor U23777 (N_23777,N_14820,N_14150);
and U23778 (N_23778,N_14044,N_12518);
or U23779 (N_23779,N_13169,N_12313);
xnor U23780 (N_23780,N_15755,N_13092);
nand U23781 (N_23781,N_16320,N_13404);
or U23782 (N_23782,N_15343,N_13418);
nand U23783 (N_23783,N_14445,N_15042);
and U23784 (N_23784,N_16325,N_13420);
nor U23785 (N_23785,N_14875,N_12908);
nor U23786 (N_23786,N_14013,N_16190);
or U23787 (N_23787,N_17811,N_15124);
xnor U23788 (N_23788,N_17392,N_16960);
nand U23789 (N_23789,N_16910,N_12412);
nor U23790 (N_23790,N_14498,N_14805);
xor U23791 (N_23791,N_17861,N_12031);
and U23792 (N_23792,N_14127,N_16785);
nand U23793 (N_23793,N_15342,N_14949);
and U23794 (N_23794,N_12823,N_13430);
or U23795 (N_23795,N_13813,N_14766);
nor U23796 (N_23796,N_17712,N_13874);
nor U23797 (N_23797,N_13291,N_17403);
and U23798 (N_23798,N_16486,N_13069);
nand U23799 (N_23799,N_17735,N_17759);
and U23800 (N_23800,N_16180,N_15318);
nor U23801 (N_23801,N_16951,N_16709);
nand U23802 (N_23802,N_15093,N_16781);
and U23803 (N_23803,N_14950,N_16688);
or U23804 (N_23804,N_15764,N_16925);
xor U23805 (N_23805,N_16282,N_17203);
nor U23806 (N_23806,N_15954,N_16653);
nor U23807 (N_23807,N_16831,N_16241);
xnor U23808 (N_23808,N_15119,N_17308);
xor U23809 (N_23809,N_14850,N_12773);
or U23810 (N_23810,N_15984,N_17631);
or U23811 (N_23811,N_12036,N_13633);
or U23812 (N_23812,N_17707,N_12055);
or U23813 (N_23813,N_14474,N_17597);
xnor U23814 (N_23814,N_13616,N_15313);
and U23815 (N_23815,N_14946,N_12602);
nand U23816 (N_23816,N_13818,N_14545);
or U23817 (N_23817,N_17531,N_14596);
and U23818 (N_23818,N_13413,N_14457);
nor U23819 (N_23819,N_16164,N_16720);
and U23820 (N_23820,N_15426,N_15364);
and U23821 (N_23821,N_13809,N_16463);
and U23822 (N_23822,N_13040,N_14686);
and U23823 (N_23823,N_16548,N_15288);
nand U23824 (N_23824,N_15130,N_12638);
nand U23825 (N_23825,N_14543,N_17676);
nor U23826 (N_23826,N_14594,N_12224);
nor U23827 (N_23827,N_14739,N_17158);
xnor U23828 (N_23828,N_15146,N_13577);
nand U23829 (N_23829,N_12542,N_17935);
xnor U23830 (N_23830,N_17322,N_16993);
nor U23831 (N_23831,N_16117,N_16128);
xnor U23832 (N_23832,N_12267,N_16116);
nor U23833 (N_23833,N_17893,N_16282);
nand U23834 (N_23834,N_12178,N_15668);
nor U23835 (N_23835,N_14661,N_14354);
or U23836 (N_23836,N_17108,N_17420);
nand U23837 (N_23837,N_16885,N_16010);
xor U23838 (N_23838,N_14511,N_14272);
nand U23839 (N_23839,N_16357,N_14310);
or U23840 (N_23840,N_13909,N_16605);
nand U23841 (N_23841,N_13141,N_13861);
nand U23842 (N_23842,N_15388,N_15722);
nand U23843 (N_23843,N_12993,N_16532);
or U23844 (N_23844,N_14736,N_14318);
or U23845 (N_23845,N_13275,N_15870);
nand U23846 (N_23846,N_17884,N_16493);
and U23847 (N_23847,N_17908,N_17995);
or U23848 (N_23848,N_15324,N_13486);
or U23849 (N_23849,N_17972,N_13741);
xor U23850 (N_23850,N_14384,N_13532);
or U23851 (N_23851,N_15915,N_14133);
nand U23852 (N_23852,N_15461,N_12199);
or U23853 (N_23853,N_12399,N_13677);
nand U23854 (N_23854,N_13697,N_14372);
nor U23855 (N_23855,N_12472,N_14319);
xnor U23856 (N_23856,N_15616,N_12965);
or U23857 (N_23857,N_16310,N_14484);
and U23858 (N_23858,N_15017,N_17303);
nand U23859 (N_23859,N_16626,N_15922);
or U23860 (N_23860,N_16974,N_13704);
nor U23861 (N_23861,N_12392,N_12643);
nor U23862 (N_23862,N_15768,N_15905);
or U23863 (N_23863,N_15363,N_17569);
xor U23864 (N_23864,N_17919,N_12683);
nand U23865 (N_23865,N_12350,N_16383);
or U23866 (N_23866,N_15028,N_14531);
nor U23867 (N_23867,N_17619,N_16485);
or U23868 (N_23868,N_12707,N_14341);
nor U23869 (N_23869,N_16140,N_12150);
nor U23870 (N_23870,N_15621,N_12563);
nor U23871 (N_23871,N_15796,N_12834);
and U23872 (N_23872,N_13019,N_16719);
nor U23873 (N_23873,N_16827,N_12917);
xnor U23874 (N_23874,N_16536,N_15713);
nor U23875 (N_23875,N_12438,N_12060);
and U23876 (N_23876,N_15825,N_16928);
and U23877 (N_23877,N_17300,N_14932);
and U23878 (N_23878,N_13129,N_15036);
nand U23879 (N_23879,N_14234,N_15703);
nand U23880 (N_23880,N_14022,N_15010);
and U23881 (N_23881,N_12914,N_17076);
xnor U23882 (N_23882,N_12473,N_13190);
or U23883 (N_23883,N_14880,N_16904);
nand U23884 (N_23884,N_13583,N_14928);
or U23885 (N_23885,N_13119,N_12976);
or U23886 (N_23886,N_17666,N_14283);
nor U23887 (N_23887,N_17999,N_14958);
nor U23888 (N_23888,N_15282,N_13359);
nand U23889 (N_23889,N_12298,N_12759);
and U23890 (N_23890,N_16321,N_12994);
or U23891 (N_23891,N_16209,N_12028);
and U23892 (N_23892,N_15649,N_13894);
and U23893 (N_23893,N_17680,N_12421);
or U23894 (N_23894,N_13903,N_17697);
and U23895 (N_23895,N_12077,N_12597);
nand U23896 (N_23896,N_17915,N_16106);
or U23897 (N_23897,N_16768,N_13387);
and U23898 (N_23898,N_13468,N_17054);
nor U23899 (N_23899,N_14609,N_14674);
and U23900 (N_23900,N_13154,N_15701);
or U23901 (N_23901,N_13081,N_15039);
nand U23902 (N_23902,N_14082,N_15067);
nor U23903 (N_23903,N_16573,N_16150);
xor U23904 (N_23904,N_13550,N_15479);
nand U23905 (N_23905,N_12550,N_16118);
or U23906 (N_23906,N_14436,N_12302);
nand U23907 (N_23907,N_14994,N_17849);
or U23908 (N_23908,N_15837,N_13982);
nand U23909 (N_23909,N_13616,N_13730);
xor U23910 (N_23910,N_14378,N_12888);
or U23911 (N_23911,N_16948,N_15732);
nand U23912 (N_23912,N_17524,N_12693);
and U23913 (N_23913,N_13944,N_13023);
nand U23914 (N_23914,N_12236,N_17507);
xor U23915 (N_23915,N_14365,N_17121);
and U23916 (N_23916,N_17622,N_16068);
xnor U23917 (N_23917,N_12209,N_17599);
nor U23918 (N_23918,N_14154,N_15485);
and U23919 (N_23919,N_13105,N_15427);
nor U23920 (N_23920,N_15799,N_16520);
xnor U23921 (N_23921,N_14763,N_14870);
xnor U23922 (N_23922,N_17370,N_12791);
and U23923 (N_23923,N_17660,N_14873);
and U23924 (N_23924,N_14422,N_13159);
or U23925 (N_23925,N_16848,N_12583);
xnor U23926 (N_23926,N_13502,N_17561);
or U23927 (N_23927,N_16631,N_12769);
or U23928 (N_23928,N_14946,N_12863);
nand U23929 (N_23929,N_16305,N_13074);
nor U23930 (N_23930,N_12877,N_16884);
nor U23931 (N_23931,N_14949,N_13611);
or U23932 (N_23932,N_14506,N_14413);
nand U23933 (N_23933,N_12090,N_16681);
nand U23934 (N_23934,N_14742,N_14223);
xnor U23935 (N_23935,N_16847,N_12268);
nor U23936 (N_23936,N_17751,N_17412);
or U23937 (N_23937,N_13134,N_13477);
or U23938 (N_23938,N_15232,N_16844);
or U23939 (N_23939,N_17989,N_17660);
nor U23940 (N_23940,N_15898,N_13917);
nor U23941 (N_23941,N_16870,N_16108);
nor U23942 (N_23942,N_12274,N_12542);
or U23943 (N_23943,N_14676,N_12405);
nand U23944 (N_23944,N_16049,N_15792);
nor U23945 (N_23945,N_16922,N_13616);
and U23946 (N_23946,N_12723,N_15296);
nor U23947 (N_23947,N_17806,N_13991);
or U23948 (N_23948,N_13288,N_14083);
nor U23949 (N_23949,N_13194,N_12058);
nand U23950 (N_23950,N_13959,N_15082);
nand U23951 (N_23951,N_15297,N_17369);
nand U23952 (N_23952,N_17307,N_13535);
nor U23953 (N_23953,N_13641,N_16858);
or U23954 (N_23954,N_17167,N_17373);
and U23955 (N_23955,N_17729,N_17676);
xnor U23956 (N_23956,N_16408,N_12099);
or U23957 (N_23957,N_12344,N_14780);
or U23958 (N_23958,N_12540,N_15244);
nand U23959 (N_23959,N_12660,N_17759);
nand U23960 (N_23960,N_14888,N_13538);
or U23961 (N_23961,N_17859,N_15782);
nand U23962 (N_23962,N_14361,N_17428);
nor U23963 (N_23963,N_14244,N_14093);
or U23964 (N_23964,N_15021,N_16466);
nand U23965 (N_23965,N_17827,N_15257);
and U23966 (N_23966,N_12625,N_13643);
xnor U23967 (N_23967,N_12981,N_17834);
or U23968 (N_23968,N_16575,N_12662);
or U23969 (N_23969,N_14830,N_17285);
or U23970 (N_23970,N_14094,N_17179);
nand U23971 (N_23971,N_16169,N_16523);
nand U23972 (N_23972,N_16660,N_16152);
nand U23973 (N_23973,N_15170,N_16857);
and U23974 (N_23974,N_12182,N_16040);
nand U23975 (N_23975,N_12130,N_17664);
and U23976 (N_23976,N_17148,N_16069);
and U23977 (N_23977,N_15158,N_14408);
or U23978 (N_23978,N_17329,N_16879);
and U23979 (N_23979,N_13479,N_12476);
nor U23980 (N_23980,N_12332,N_14971);
xnor U23981 (N_23981,N_16629,N_15289);
nor U23982 (N_23982,N_13908,N_12330);
or U23983 (N_23983,N_13192,N_14101);
nand U23984 (N_23984,N_16204,N_15742);
nor U23985 (N_23985,N_12257,N_13948);
and U23986 (N_23986,N_15427,N_13006);
or U23987 (N_23987,N_17452,N_12900);
xnor U23988 (N_23988,N_15065,N_14485);
nand U23989 (N_23989,N_13722,N_12580);
nand U23990 (N_23990,N_13327,N_13868);
or U23991 (N_23991,N_17341,N_16225);
or U23992 (N_23992,N_15068,N_12338);
nand U23993 (N_23993,N_12498,N_16274);
nor U23994 (N_23994,N_17488,N_15371);
nand U23995 (N_23995,N_13484,N_15403);
nand U23996 (N_23996,N_15276,N_12493);
xnor U23997 (N_23997,N_17484,N_13832);
nand U23998 (N_23998,N_13284,N_15305);
xnor U23999 (N_23999,N_15347,N_14694);
or U24000 (N_24000,N_18591,N_22793);
nor U24001 (N_24001,N_22060,N_20544);
nand U24002 (N_24002,N_18742,N_19159);
nor U24003 (N_24003,N_23486,N_19796);
or U24004 (N_24004,N_20978,N_20687);
xor U24005 (N_24005,N_21825,N_21553);
nand U24006 (N_24006,N_23415,N_23037);
and U24007 (N_24007,N_20854,N_20578);
or U24008 (N_24008,N_20394,N_21709);
nand U24009 (N_24009,N_22298,N_23418);
nand U24010 (N_24010,N_21640,N_20074);
nor U24011 (N_24011,N_18348,N_19279);
nand U24012 (N_24012,N_23665,N_21969);
and U24013 (N_24013,N_23188,N_21592);
xnor U24014 (N_24014,N_20789,N_21841);
and U24015 (N_24015,N_21998,N_21874);
and U24016 (N_24016,N_23688,N_22147);
xor U24017 (N_24017,N_19287,N_21059);
or U24018 (N_24018,N_21144,N_19415);
nand U24019 (N_24019,N_18273,N_22500);
or U24020 (N_24020,N_22324,N_23777);
and U24021 (N_24021,N_20735,N_22317);
nand U24022 (N_24022,N_20292,N_20467);
nand U24023 (N_24023,N_21922,N_21618);
and U24024 (N_24024,N_22747,N_19151);
xnor U24025 (N_24025,N_20016,N_20300);
and U24026 (N_24026,N_23750,N_18843);
nand U24027 (N_24027,N_23247,N_21426);
nand U24028 (N_24028,N_20482,N_20895);
nand U24029 (N_24029,N_23467,N_18907);
and U24030 (N_24030,N_18604,N_18326);
and U24031 (N_24031,N_21780,N_22307);
or U24032 (N_24032,N_20620,N_20543);
and U24033 (N_24033,N_20521,N_21485);
or U24034 (N_24034,N_21529,N_22670);
xor U24035 (N_24035,N_18147,N_23899);
xor U24036 (N_24036,N_22337,N_20659);
nor U24037 (N_24037,N_22780,N_23321);
nor U24038 (N_24038,N_21774,N_21082);
and U24039 (N_24039,N_22020,N_20489);
and U24040 (N_24040,N_20990,N_18140);
nand U24041 (N_24041,N_20776,N_21562);
nor U24042 (N_24042,N_18322,N_19449);
nand U24043 (N_24043,N_18915,N_21542);
nand U24044 (N_24044,N_21465,N_21727);
nor U24045 (N_24045,N_23354,N_23838);
and U24046 (N_24046,N_18427,N_22244);
and U24047 (N_24047,N_22438,N_19184);
nor U24048 (N_24048,N_18357,N_20294);
nor U24049 (N_24049,N_22975,N_19305);
nand U24050 (N_24050,N_18696,N_21768);
nand U24051 (N_24051,N_20162,N_23618);
or U24052 (N_24052,N_19810,N_22136);
xor U24053 (N_24053,N_20275,N_23323);
nor U24054 (N_24054,N_18799,N_18557);
and U24055 (N_24055,N_22518,N_21717);
and U24056 (N_24056,N_19791,N_20425);
nor U24057 (N_24057,N_18004,N_18220);
nor U24058 (N_24058,N_21526,N_23461);
nor U24059 (N_24059,N_20032,N_18613);
or U24060 (N_24060,N_21375,N_18947);
nor U24061 (N_24061,N_20962,N_21677);
nor U24062 (N_24062,N_21633,N_23197);
nor U24063 (N_24063,N_18049,N_23196);
nand U24064 (N_24064,N_23042,N_20062);
or U24065 (N_24065,N_20638,N_19747);
and U24066 (N_24066,N_19120,N_20837);
and U24067 (N_24067,N_22185,N_19511);
or U24068 (N_24068,N_20167,N_23525);
nand U24069 (N_24069,N_21731,N_18761);
and U24070 (N_24070,N_19646,N_21885);
and U24071 (N_24071,N_23515,N_22669);
or U24072 (N_24072,N_21901,N_20959);
and U24073 (N_24073,N_22730,N_22375);
xor U24074 (N_24074,N_22373,N_22570);
or U24075 (N_24075,N_23979,N_22727);
and U24076 (N_24076,N_18228,N_21133);
nor U24077 (N_24077,N_22674,N_20897);
xnor U24078 (N_24078,N_18683,N_21718);
nor U24079 (N_24079,N_20081,N_20720);
nor U24080 (N_24080,N_21879,N_19825);
nand U24081 (N_24081,N_20546,N_20192);
nand U24082 (N_24082,N_21395,N_23768);
nand U24083 (N_24083,N_21685,N_19492);
and U24084 (N_24084,N_19008,N_20739);
nand U24085 (N_24085,N_22546,N_21594);
or U24086 (N_24086,N_23306,N_20665);
nor U24087 (N_24087,N_23405,N_22403);
and U24088 (N_24088,N_22251,N_19975);
nor U24089 (N_24089,N_23842,N_20039);
xnor U24090 (N_24090,N_18318,N_19389);
nor U24091 (N_24091,N_23945,N_23076);
and U24092 (N_24092,N_21971,N_20295);
or U24093 (N_24093,N_20820,N_19317);
or U24094 (N_24094,N_23684,N_21566);
nand U24095 (N_24095,N_19600,N_18744);
nand U24096 (N_24096,N_21453,N_21489);
nand U24097 (N_24097,N_21948,N_18405);
xnor U24098 (N_24098,N_18050,N_23474);
and U24099 (N_24099,N_20014,N_23767);
nor U24100 (N_24100,N_21050,N_19863);
nand U24101 (N_24101,N_19461,N_23692);
nand U24102 (N_24102,N_18837,N_21076);
and U24103 (N_24103,N_22031,N_21211);
nor U24104 (N_24104,N_20847,N_23381);
and U24105 (N_24105,N_20130,N_22114);
nand U24106 (N_24106,N_23783,N_23529);
nor U24107 (N_24107,N_23299,N_22914);
nand U24108 (N_24108,N_23335,N_19233);
and U24109 (N_24109,N_20148,N_21365);
xnor U24110 (N_24110,N_21800,N_22301);
nand U24111 (N_24111,N_19813,N_22666);
or U24112 (N_24112,N_18467,N_21267);
nor U24113 (N_24113,N_18292,N_19181);
or U24114 (N_24114,N_21330,N_21600);
nand U24115 (N_24115,N_21860,N_18756);
and U24116 (N_24116,N_19903,N_21246);
nor U24117 (N_24117,N_18227,N_21419);
nor U24118 (N_24118,N_18990,N_18370);
and U24119 (N_24119,N_20313,N_18387);
and U24120 (N_24120,N_18266,N_18710);
and U24121 (N_24121,N_20883,N_22163);
and U24122 (N_24122,N_23148,N_23357);
nand U24123 (N_24123,N_18859,N_20540);
and U24124 (N_24124,N_23911,N_18008);
nor U24125 (N_24125,N_18233,N_19998);
and U24126 (N_24126,N_22755,N_23030);
nor U24127 (N_24127,N_23186,N_20538);
or U24128 (N_24128,N_23159,N_21673);
or U24129 (N_24129,N_18075,N_22376);
xor U24130 (N_24130,N_23809,N_23730);
nor U24131 (N_24131,N_20189,N_20395);
or U24132 (N_24132,N_18983,N_19471);
xnor U24133 (N_24133,N_21507,N_21480);
nor U24134 (N_24134,N_21366,N_18987);
or U24135 (N_24135,N_23413,N_23457);
nor U24136 (N_24136,N_21493,N_23780);
and U24137 (N_24137,N_20670,N_21567);
nor U24138 (N_24138,N_23845,N_21397);
nand U24139 (N_24139,N_22109,N_22004);
and U24140 (N_24140,N_18412,N_18719);
or U24141 (N_24141,N_20663,N_23661);
nor U24142 (N_24142,N_22717,N_20184);
nor U24143 (N_24143,N_21369,N_19856);
nor U24144 (N_24144,N_20612,N_18299);
or U24145 (N_24145,N_20226,N_20080);
or U24146 (N_24146,N_20825,N_18737);
or U24147 (N_24147,N_20349,N_23640);
nand U24148 (N_24148,N_23479,N_20590);
and U24149 (N_24149,N_22140,N_18964);
nand U24150 (N_24150,N_18995,N_22826);
nor U24151 (N_24151,N_21137,N_19585);
xnor U24152 (N_24152,N_23353,N_19862);
xnor U24153 (N_24153,N_21354,N_19333);
and U24154 (N_24154,N_20332,N_22841);
nor U24155 (N_24155,N_21649,N_21794);
nor U24156 (N_24156,N_20966,N_18091);
and U24157 (N_24157,N_20449,N_23861);
or U24158 (N_24158,N_19841,N_20417);
or U24159 (N_24159,N_19092,N_19239);
and U24160 (N_24160,N_21376,N_20055);
nor U24161 (N_24161,N_19493,N_23904);
nor U24162 (N_24162,N_22724,N_20928);
or U24163 (N_24163,N_19078,N_22702);
nor U24164 (N_24164,N_19774,N_20823);
and U24165 (N_24165,N_21411,N_23850);
nor U24166 (N_24166,N_19743,N_20364);
xor U24167 (N_24167,N_21067,N_19827);
or U24168 (N_24168,N_18530,N_21071);
nor U24169 (N_24169,N_20605,N_18500);
and U24170 (N_24170,N_22206,N_21044);
or U24171 (N_24171,N_20899,N_18388);
nor U24172 (N_24172,N_18477,N_23227);
xor U24173 (N_24173,N_21864,N_18222);
or U24174 (N_24174,N_21103,N_21534);
or U24175 (N_24175,N_18338,N_20264);
and U24176 (N_24176,N_20678,N_20064);
nor U24177 (N_24177,N_22773,N_23012);
nor U24178 (N_24178,N_23604,N_23967);
or U24179 (N_24179,N_21997,N_23960);
nor U24180 (N_24180,N_21243,N_18706);
nor U24181 (N_24181,N_18209,N_23582);
and U24182 (N_24182,N_19028,N_23341);
nand U24183 (N_24183,N_22582,N_19327);
nand U24184 (N_24184,N_18638,N_18930);
xor U24185 (N_24185,N_22794,N_19535);
and U24186 (N_24186,N_21944,N_22475);
nor U24187 (N_24187,N_22810,N_22271);
nor U24188 (N_24188,N_22385,N_21152);
xor U24189 (N_24189,N_21325,N_21593);
xnor U24190 (N_24190,N_21266,N_19529);
or U24191 (N_24191,N_22377,N_19665);
and U24192 (N_24192,N_21464,N_21272);
nand U24193 (N_24193,N_18923,N_21737);
nand U24194 (N_24194,N_20229,N_20542);
xor U24195 (N_24195,N_18077,N_20366);
and U24196 (N_24196,N_20481,N_22563);
and U24197 (N_24197,N_23478,N_21916);
nor U24198 (N_24198,N_21488,N_20602);
and U24199 (N_24199,N_19296,N_23900);
nor U24200 (N_24200,N_21976,N_22188);
or U24201 (N_24201,N_20796,N_22953);
xor U24202 (N_24202,N_18496,N_22557);
nor U24203 (N_24203,N_21565,N_21006);
nor U24204 (N_24204,N_21691,N_20179);
or U24205 (N_24205,N_20375,N_22866);
nor U24206 (N_24206,N_18251,N_19572);
nand U24207 (N_24207,N_20971,N_22587);
and U24208 (N_24208,N_22692,N_19270);
xnor U24209 (N_24209,N_22567,N_20925);
xor U24210 (N_24210,N_19926,N_20180);
nor U24211 (N_24211,N_22941,N_19023);
and U24212 (N_24212,N_19524,N_22925);
nor U24213 (N_24213,N_21017,N_21966);
xor U24214 (N_24214,N_21106,N_20286);
nand U24215 (N_24215,N_23603,N_19635);
nor U24216 (N_24216,N_19306,N_18373);
xnor U24217 (N_24217,N_22121,N_19262);
or U24218 (N_24218,N_19976,N_19067);
and U24219 (N_24219,N_20894,N_18047);
and U24220 (N_24220,N_20611,N_19417);
nor U24221 (N_24221,N_21300,N_23984);
nand U24222 (N_24222,N_21757,N_19912);
nand U24223 (N_24223,N_18836,N_18079);
or U24224 (N_24224,N_18404,N_22857);
xor U24225 (N_24225,N_22005,N_21883);
or U24226 (N_24226,N_19961,N_20463);
nand U24227 (N_24227,N_23416,N_20912);
and U24228 (N_24228,N_21172,N_18128);
nand U24229 (N_24229,N_18991,N_21900);
nand U24230 (N_24230,N_22085,N_19872);
nand U24231 (N_24231,N_19176,N_21695);
or U24232 (N_24232,N_21316,N_20083);
nand U24233 (N_24233,N_19753,N_18498);
or U24234 (N_24234,N_18752,N_21753);
xnor U24235 (N_24235,N_20779,N_22365);
nor U24236 (N_24236,N_19993,N_19195);
nor U24237 (N_24237,N_18081,N_19981);
or U24238 (N_24238,N_20276,N_18482);
or U24239 (N_24239,N_21165,N_18682);
and U24240 (N_24240,N_18337,N_19057);
and U24241 (N_24241,N_21240,N_21089);
xor U24242 (N_24242,N_21867,N_21560);
or U24243 (N_24243,N_19016,N_19678);
and U24244 (N_24244,N_23107,N_20690);
and U24245 (N_24245,N_21229,N_22346);
nand U24246 (N_24246,N_19102,N_21742);
nor U24247 (N_24247,N_18774,N_19478);
nor U24248 (N_24248,N_23224,N_19125);
nand U24249 (N_24249,N_20245,N_23395);
or U24250 (N_24250,N_22710,N_18522);
nand U24251 (N_24251,N_18331,N_20545);
nor U24252 (N_24252,N_23814,N_20304);
and U24253 (N_24253,N_20501,N_20821);
and U24254 (N_24254,N_20655,N_20673);
or U24255 (N_24255,N_18981,N_18631);
and U24256 (N_24256,N_23480,N_23262);
or U24257 (N_24257,N_22167,N_19574);
and U24258 (N_24258,N_20900,N_20480);
nand U24259 (N_24259,N_18898,N_18224);
nor U24260 (N_24260,N_21555,N_18720);
or U24261 (N_24261,N_18608,N_22023);
or U24262 (N_24262,N_23837,N_22135);
xor U24263 (N_24263,N_19990,N_22082);
nand U24264 (N_24264,N_19359,N_20686);
nor U24265 (N_24265,N_19628,N_18254);
xnor U24266 (N_24266,N_22069,N_19174);
or U24267 (N_24267,N_21644,N_23512);
nor U24268 (N_24268,N_23709,N_22994);
and U24269 (N_24269,N_22433,N_20236);
and U24270 (N_24270,N_21228,N_20839);
or U24271 (N_24271,N_18126,N_21256);
nand U24272 (N_24272,N_21060,N_20432);
nor U24273 (N_24273,N_22656,N_19656);
and U24274 (N_24274,N_20944,N_18784);
nand U24275 (N_24275,N_18708,N_19439);
nand U24276 (N_24276,N_23174,N_20806);
and U24277 (N_24277,N_19892,N_20051);
nand U24278 (N_24278,N_21607,N_23446);
xor U24279 (N_24279,N_20293,N_20740);
nand U24280 (N_24280,N_21161,N_19475);
and U24281 (N_24281,N_23150,N_23071);
and U24282 (N_24282,N_18447,N_22574);
and U24283 (N_24283,N_23101,N_18377);
or U24284 (N_24284,N_23060,N_18645);
nor U24285 (N_24285,N_19653,N_20552);
xnor U24286 (N_24286,N_18432,N_19323);
nand U24287 (N_24287,N_21866,N_19851);
nand U24288 (N_24288,N_21798,N_22480);
or U24289 (N_24289,N_22673,N_21662);
nor U24290 (N_24290,N_21439,N_22164);
xor U24291 (N_24291,N_21745,N_21470);
nand U24292 (N_24292,N_19889,N_20694);
nand U24293 (N_24293,N_20154,N_23541);
and U24294 (N_24294,N_21062,N_21982);
xnor U24295 (N_24295,N_23737,N_19787);
nand U24296 (N_24296,N_20078,N_21069);
or U24297 (N_24297,N_20352,N_20774);
and U24298 (N_24298,N_22254,N_18911);
or U24299 (N_24299,N_20911,N_19559);
nor U24300 (N_24300,N_19380,N_22162);
xor U24301 (N_24301,N_18562,N_23172);
and U24302 (N_24302,N_18842,N_19466);
xor U24303 (N_24303,N_21833,N_23517);
nor U24304 (N_24304,N_22573,N_18693);
or U24305 (N_24305,N_22221,N_19060);
nand U24306 (N_24306,N_18421,N_23587);
or U24307 (N_24307,N_21838,N_19698);
nand U24308 (N_24308,N_23275,N_21206);
nand U24309 (N_24309,N_22002,N_22906);
xor U24310 (N_24310,N_23766,N_19875);
and U24311 (N_24311,N_21769,N_22840);
and U24312 (N_24312,N_18570,N_21094);
or U24313 (N_24313,N_21919,N_23173);
or U24314 (N_24314,N_19071,N_23852);
or U24315 (N_24315,N_22583,N_18466);
nand U24316 (N_24316,N_23986,N_19285);
and U24317 (N_24317,N_19697,N_18435);
nand U24318 (N_24318,N_19189,N_21558);
nor U24319 (N_24319,N_18606,N_19798);
and U24320 (N_24320,N_20407,N_22217);
and U24321 (N_24321,N_19596,N_19477);
nand U24322 (N_24322,N_19293,N_21019);
nor U24323 (N_24323,N_19036,N_21804);
nor U24324 (N_24324,N_23053,N_19281);
nor U24325 (N_24325,N_21574,N_19379);
nand U24326 (N_24326,N_22058,N_21937);
nor U24327 (N_24327,N_18345,N_18506);
nor U24328 (N_24328,N_22985,N_23181);
nor U24329 (N_24329,N_20608,N_21265);
nand U24330 (N_24330,N_19055,N_22675);
nor U24331 (N_24331,N_18476,N_22350);
nand U24332 (N_24332,N_23119,N_23505);
and U24333 (N_24333,N_22203,N_18669);
or U24334 (N_24334,N_18136,N_19548);
nor U24335 (N_24335,N_19828,N_22942);
or U24336 (N_24336,N_21079,N_20135);
and U24337 (N_24337,N_21713,N_19232);
and U24338 (N_24338,N_19474,N_19134);
xor U24339 (N_24339,N_21672,N_20539);
nand U24340 (N_24340,N_18650,N_23230);
nand U24341 (N_24341,N_18581,N_20744);
or U24342 (N_24342,N_18440,N_21886);
and U24343 (N_24343,N_21538,N_23261);
nand U24344 (N_24344,N_22243,N_18402);
and U24345 (N_24345,N_22202,N_19291);
or U24346 (N_24346,N_18367,N_23612);
and U24347 (N_24347,N_20792,N_19623);
nor U24348 (N_24348,N_19256,N_20798);
nand U24349 (N_24349,N_21182,N_18505);
or U24350 (N_24350,N_22105,N_23294);
nand U24351 (N_24351,N_20824,N_21875);
and U24352 (N_24352,N_21087,N_18146);
or U24353 (N_24353,N_21167,N_18112);
nand U24354 (N_24354,N_22699,N_22455);
or U24355 (N_24355,N_23745,N_18609);
or U24356 (N_24356,N_22310,N_20136);
and U24357 (N_24357,N_22124,N_21648);
and U24358 (N_24358,N_20222,N_21471);
and U24359 (N_24359,N_19240,N_22939);
nor U24360 (N_24360,N_19594,N_18463);
nand U24361 (N_24361,N_19541,N_18879);
or U24362 (N_24362,N_22623,N_19950);
xnor U24363 (N_24363,N_19497,N_23317);
xor U24364 (N_24364,N_22288,N_23207);
and U24365 (N_24365,N_18763,N_19978);
nor U24366 (N_24366,N_22600,N_23589);
nand U24367 (N_24367,N_21975,N_21651);
nor U24368 (N_24368,N_20337,N_19179);
xnor U24369 (N_24369,N_21850,N_23220);
nand U24370 (N_24370,N_18445,N_18518);
nor U24371 (N_24371,N_21616,N_19703);
or U24372 (N_24372,N_21950,N_23198);
or U24373 (N_24373,N_22458,N_19680);
and U24374 (N_24374,N_21043,N_19599);
and U24375 (N_24375,N_20931,N_20593);
xor U24376 (N_24376,N_18335,N_18150);
and U24377 (N_24377,N_19545,N_23371);
nand U24378 (N_24378,N_22149,N_23811);
nor U24379 (N_24379,N_19878,N_23470);
or U24380 (N_24380,N_18940,N_19253);
and U24381 (N_24381,N_18688,N_21350);
nand U24382 (N_24382,N_18198,N_19140);
nand U24383 (N_24383,N_19393,N_19971);
nor U24384 (N_24384,N_23564,N_18226);
and U24385 (N_24385,N_22395,N_20240);
and U24386 (N_24386,N_21571,N_22595);
or U24387 (N_24387,N_21097,N_21809);
nor U24388 (N_24388,N_18044,N_21360);
nand U24389 (N_24389,N_19946,N_20408);
nor U24390 (N_24390,N_18712,N_19068);
or U24391 (N_24391,N_21583,N_21924);
xnor U24392 (N_24392,N_23794,N_21889);
xnor U24393 (N_24393,N_21456,N_23919);
xor U24394 (N_24394,N_21552,N_22534);
and U24395 (N_24395,N_23453,N_21048);
nand U24396 (N_24396,N_20946,N_20564);
xor U24397 (N_24397,N_19898,N_23365);
xor U24398 (N_24398,N_18231,N_18828);
xor U24399 (N_24399,N_20471,N_21793);
and U24400 (N_24400,N_20008,N_23514);
and U24401 (N_24401,N_21314,N_23014);
nor U24402 (N_24402,N_23376,N_18384);
and U24403 (N_24403,N_19652,N_18071);
and U24404 (N_24404,N_23477,N_19962);
or U24405 (N_24405,N_22415,N_23624);
or U24406 (N_24406,N_18538,N_23905);
nor U24407 (N_24407,N_21258,N_23350);
and U24408 (N_24408,N_22388,N_21118);
or U24409 (N_24409,N_20967,N_23260);
nor U24410 (N_24410,N_22222,N_21675);
nor U24411 (N_24411,N_20802,N_21099);
nand U24412 (N_24412,N_22401,N_21641);
nor U24413 (N_24413,N_22503,N_23072);
nand U24414 (N_24414,N_23382,N_18428);
nor U24415 (N_24415,N_18814,N_19713);
or U24416 (N_24416,N_20152,N_20983);
nand U24417 (N_24417,N_22033,N_23191);
and U24418 (N_24418,N_21778,N_21911);
nor U24419 (N_24419,N_19601,N_23568);
nand U24420 (N_24420,N_20139,N_19900);
or U24421 (N_24421,N_20807,N_20217);
or U24422 (N_24422,N_22653,N_21789);
and U24423 (N_24423,N_21665,N_19761);
nand U24424 (N_24424,N_23211,N_23932);
nor U24425 (N_24425,N_18362,N_21289);
nand U24426 (N_24426,N_18301,N_23913);
and U24427 (N_24427,N_18003,N_18169);
nor U24428 (N_24428,N_22501,N_22099);
nand U24429 (N_24429,N_18212,N_21497);
or U24430 (N_24430,N_21792,N_18648);
or U24431 (N_24431,N_23848,N_23423);
nor U24432 (N_24432,N_20140,N_22348);
or U24433 (N_24433,N_22540,N_20428);
nand U24434 (N_24434,N_18309,N_18932);
and U24435 (N_24435,N_18130,N_18230);
xnor U24436 (N_24436,N_23310,N_21773);
nand U24437 (N_24437,N_20903,N_22657);
nor U24438 (N_24438,N_20936,N_18565);
nand U24439 (N_24439,N_19170,N_23417);
or U24440 (N_24440,N_18769,N_18257);
nand U24441 (N_24441,N_20566,N_22111);
nand U24442 (N_24442,N_19457,N_18268);
nand U24443 (N_24443,N_20705,N_19927);
nand U24444 (N_24444,N_19522,N_23548);
nor U24445 (N_24445,N_18630,N_23366);
nor U24446 (N_24446,N_21352,N_21026);
nand U24447 (N_24447,N_20650,N_18457);
nand U24448 (N_24448,N_18728,N_21909);
nor U24449 (N_24449,N_20289,N_20943);
nor U24450 (N_24450,N_18415,N_22431);
nand U24451 (N_24451,N_18647,N_18705);
nand U24452 (N_24452,N_19781,N_19476);
or U24453 (N_24453,N_18839,N_21634);
nand U24454 (N_24454,N_20872,N_22476);
and U24455 (N_24455,N_23798,N_20447);
nor U24456 (N_24456,N_21810,N_22787);
nor U24457 (N_24457,N_23106,N_22523);
nand U24458 (N_24458,N_20737,N_18078);
or U24459 (N_24459,N_22413,N_18471);
xor U24460 (N_24460,N_23146,N_22482);
nand U24461 (N_24461,N_18778,N_19375);
or U24462 (N_24462,N_22648,N_19918);
nor U24463 (N_24463,N_19320,N_23721);
nand U24464 (N_24464,N_20353,N_20299);
or U24465 (N_24465,N_20508,N_20851);
and U24466 (N_24466,N_23853,N_21361);
nand U24467 (N_24467,N_22853,N_22817);
and U24468 (N_24468,N_18238,N_19789);
and U24469 (N_24469,N_22402,N_22021);
and U24470 (N_24470,N_21199,N_20041);
nor U24471 (N_24471,N_20019,N_21827);
and U24472 (N_24472,N_18278,N_19326);
nor U24473 (N_24473,N_22224,N_20994);
xnor U24474 (N_24474,N_22616,N_18858);
and U24475 (N_24475,N_20347,N_22483);
nor U24476 (N_24476,N_20159,N_20923);
or U24477 (N_24477,N_23677,N_23723);
nand U24478 (N_24478,N_22931,N_23944);
nand U24479 (N_24479,N_18247,N_19182);
xnor U24480 (N_24480,N_23094,N_22586);
or U24481 (N_24481,N_21142,N_19696);
nor U24482 (N_24482,N_23574,N_18028);
and U24483 (N_24483,N_20054,N_22040);
xor U24484 (N_24484,N_19007,N_18759);
nor U24485 (N_24485,N_18588,N_19839);
or U24486 (N_24486,N_23637,N_22988);
nand U24487 (N_24487,N_23167,N_18066);
nor U24488 (N_24488,N_21157,N_18797);
nor U24489 (N_24489,N_19741,N_21363);
xor U24490 (N_24490,N_21054,N_20216);
nand U24491 (N_24491,N_20077,N_22446);
nor U24492 (N_24492,N_18640,N_20992);
nand U24493 (N_24493,N_22642,N_20384);
or U24494 (N_24494,N_20336,N_21057);
nand U24495 (N_24495,N_20919,N_20183);
and U24496 (N_24496,N_20360,N_22016);
or U24497 (N_24497,N_22678,N_21812);
nor U24498 (N_24498,N_22326,N_18743);
or U24499 (N_24499,N_23133,N_19592);
or U24500 (N_24500,N_20646,N_21214);
nor U24501 (N_24501,N_21338,N_21891);
nor U24502 (N_24502,N_22788,N_20142);
or U24503 (N_24503,N_23623,N_22977);
nor U24504 (N_24504,N_18142,N_23879);
nor U24505 (N_24505,N_18152,N_19913);
and U24506 (N_24506,N_23336,N_20531);
xor U24507 (N_24507,N_23866,N_21307);
nor U24508 (N_24508,N_22323,N_18276);
and U24509 (N_24509,N_18757,N_19226);
or U24510 (N_24510,N_19470,N_21910);
and U24511 (N_24511,N_20338,N_22132);
and U24512 (N_24512,N_18926,N_18969);
or U24513 (N_24513,N_19304,N_18244);
nand U24514 (N_24514,N_21158,N_22913);
and U24515 (N_24515,N_23595,N_20688);
or U24516 (N_24516,N_19777,N_23266);
or U24517 (N_24517,N_23531,N_22112);
or U24518 (N_24518,N_20389,N_20574);
and U24519 (N_24519,N_20208,N_21110);
nor U24520 (N_24520,N_21473,N_21114);
nand U24521 (N_24521,N_22339,N_20722);
nor U24522 (N_24522,N_19101,N_19609);
nor U24523 (N_24523,N_23482,N_21368);
or U24524 (N_24524,N_20233,N_19843);
and U24525 (N_24525,N_18989,N_19443);
nor U24526 (N_24526,N_18596,N_22974);
and U24527 (N_24527,N_18794,N_22877);
and U24528 (N_24528,N_18011,N_19832);
nand U24529 (N_24529,N_18820,N_18030);
and U24530 (N_24530,N_22426,N_21382);
nor U24531 (N_24531,N_21877,N_20422);
and U24532 (N_24532,N_18250,N_21126);
or U24533 (N_24533,N_21954,N_22095);
nand U24534 (N_24534,N_19308,N_23152);
nand U24535 (N_24535,N_23717,N_19723);
and U24536 (N_24536,N_20131,N_20121);
or U24537 (N_24537,N_21588,N_23057);
nor U24538 (N_24538,N_21457,N_23473);
or U24539 (N_24539,N_22605,N_22883);
and U24540 (N_24540,N_23871,N_18176);
nor U24541 (N_24541,N_23494,N_18881);
or U24542 (N_24542,N_20558,N_19146);
and U24543 (N_24543,N_19669,N_23755);
nor U24544 (N_24544,N_18074,N_20708);
nand U24545 (N_24545,N_21055,N_21579);
nand U24546 (N_24546,N_23887,N_20017);
and U24547 (N_24547,N_20549,N_23751);
xor U24548 (N_24548,N_23931,N_21221);
and U24549 (N_24549,N_21676,N_19177);
and U24550 (N_24550,N_20043,N_20072);
or U24551 (N_24551,N_19165,N_20814);
nor U24552 (N_24552,N_23458,N_19852);
nor U24553 (N_24553,N_23825,N_21010);
or U24554 (N_24554,N_20742,N_21706);
xor U24555 (N_24555,N_22516,N_19752);
nand U24556 (N_24556,N_18489,N_20397);
and U24557 (N_24557,N_18670,N_23171);
xnor U24558 (N_24558,N_23386,N_19505);
nand U24559 (N_24559,N_21117,N_20986);
and U24560 (N_24560,N_23539,N_21831);
xor U24561 (N_24561,N_21400,N_20654);
nor U24562 (N_24562,N_22749,N_23285);
or U24563 (N_24563,N_18114,N_22151);
xor U24564 (N_24564,N_21687,N_18904);
nand U24565 (N_24565,N_21232,N_18022);
or U24566 (N_24566,N_21430,N_21801);
or U24567 (N_24567,N_22044,N_22218);
and U24568 (N_24568,N_22220,N_23450);
and U24569 (N_24569,N_22525,N_21596);
nand U24570 (N_24570,N_20835,N_21708);
nand U24571 (N_24571,N_20734,N_23540);
nand U24572 (N_24572,N_18521,N_22828);
and U24573 (N_24573,N_21249,N_21164);
or U24574 (N_24574,N_23560,N_19412);
and U24575 (N_24575,N_21740,N_20383);
nand U24576 (N_24576,N_20497,N_22039);
nor U24577 (N_24577,N_22406,N_20253);
and U24578 (N_24578,N_19197,N_22541);
or U24579 (N_24579,N_23973,N_23346);
and U24580 (N_24580,N_22357,N_19506);
or U24581 (N_24581,N_22432,N_18403);
nor U24582 (N_24582,N_20382,N_20312);
or U24583 (N_24583,N_18097,N_22437);
nor U24584 (N_24584,N_22133,N_19691);
nand U24585 (N_24585,N_22978,N_20656);
nand U24586 (N_24586,N_21598,N_18636);
or U24587 (N_24587,N_21449,N_21970);
or U24588 (N_24588,N_22463,N_20682);
xnor U24589 (N_24589,N_20857,N_21720);
nor U24590 (N_24590,N_21904,N_18013);
nor U24591 (N_24591,N_21009,N_22989);
nand U24592 (N_24592,N_19538,N_19830);
nand U24593 (N_24593,N_19933,N_19649);
nor U24594 (N_24594,N_21065,N_21839);
nor U24595 (N_24595,N_18830,N_19807);
nand U24596 (N_24596,N_20704,N_20917);
nor U24597 (N_24597,N_20913,N_22728);
nor U24598 (N_24598,N_21432,N_20581);
or U24599 (N_24599,N_20767,N_22113);
or U24600 (N_24600,N_21930,N_21188);
nand U24601 (N_24601,N_18724,N_23597);
nand U24602 (N_24602,N_18829,N_20230);
nor U24603 (N_24603,N_23284,N_22533);
or U24604 (N_24604,N_23046,N_21113);
and U24605 (N_24605,N_22396,N_18555);
and U24606 (N_24606,N_21250,N_20033);
nand U24607 (N_24607,N_21724,N_18453);
and U24608 (N_24608,N_19214,N_21659);
xor U24609 (N_24609,N_23736,N_23351);
or U24610 (N_24610,N_23696,N_19893);
nand U24611 (N_24611,N_22923,N_20049);
or U24612 (N_24612,N_20004,N_21402);
nor U24613 (N_24613,N_21931,N_22638);
nand U24614 (N_24614,N_21549,N_19370);
nand U24615 (N_24615,N_23602,N_18064);
nand U24616 (N_24616,N_23025,N_18137);
nand U24617 (N_24617,N_19717,N_22076);
nand U24618 (N_24618,N_19654,N_18838);
or U24619 (N_24619,N_18986,N_22349);
nand U24620 (N_24620,N_23551,N_19560);
or U24621 (N_24621,N_21722,N_22238);
nand U24622 (N_24622,N_21101,N_23398);
nor U24623 (N_24623,N_20034,N_21239);
or U24624 (N_24624,N_23311,N_19923);
and U24625 (N_24625,N_20341,N_18484);
nor U24626 (N_24626,N_22854,N_20805);
nand U24627 (N_24627,N_19801,N_22952);
or U24628 (N_24628,N_23889,N_23139);
nand U24629 (N_24629,N_23448,N_18871);
and U24630 (N_24630,N_23629,N_20727);
nor U24631 (N_24631,N_21947,N_21888);
nor U24632 (N_24632,N_19881,N_19468);
or U24633 (N_24633,N_20562,N_21508);
nor U24634 (N_24634,N_19939,N_21514);
xor U24635 (N_24635,N_21528,N_21056);
nand U24636 (N_24636,N_22867,N_23915);
or U24637 (N_24637,N_20624,N_21111);
nor U24638 (N_24638,N_23318,N_18869);
or U24639 (N_24639,N_20904,N_18817);
and U24640 (N_24640,N_18184,N_23647);
and U24641 (N_24641,N_18572,N_22617);
nand U24642 (N_24642,N_23135,N_20866);
or U24643 (N_24643,N_20797,N_22495);
or U24644 (N_24644,N_23980,N_18856);
nor U24645 (N_24645,N_23731,N_21674);
and U24646 (N_24646,N_19530,N_22972);
nand U24647 (N_24647,N_20567,N_19965);
nor U24648 (N_24648,N_20093,N_22834);
and U24649 (N_24649,N_20537,N_23993);
and U24650 (N_24650,N_20648,N_23909);
or U24651 (N_24651,N_21186,N_19376);
and U24652 (N_24652,N_19034,N_23572);
or U24653 (N_24653,N_22709,N_22962);
nand U24654 (N_24654,N_20662,N_23527);
nor U24655 (N_24655,N_20743,N_19113);
nand U24656 (N_24656,N_22522,N_21550);
nor U24657 (N_24657,N_21237,N_19344);
or U24658 (N_24658,N_22812,N_19451);
nand U24659 (N_24659,N_21296,N_19073);
nor U24660 (N_24660,N_21999,N_19194);
xnor U24661 (N_24661,N_19797,N_20875);
nand U24662 (N_24662,N_20199,N_21295);
xor U24663 (N_24663,N_19952,N_20935);
xnor U24664 (N_24664,N_23655,N_23728);
nand U24665 (N_24665,N_18192,N_20933);
nand U24666 (N_24666,N_18548,N_18512);
or U24667 (N_24667,N_22226,N_19352);
nor U24668 (N_24668,N_20320,N_18143);
or U24669 (N_24669,N_22228,N_22682);
nand U24670 (N_24670,N_18840,N_18525);
or U24671 (N_24671,N_21617,N_21513);
nand U24672 (N_24672,N_18618,N_18722);
and U24673 (N_24673,N_21725,N_20715);
nor U24674 (N_24674,N_19751,N_18589);
xnor U24675 (N_24675,N_22367,N_23841);
or U24676 (N_24676,N_18741,N_23123);
or U24677 (N_24677,N_19683,N_23823);
and U24678 (N_24678,N_23545,N_19249);
and U24679 (N_24679,N_23881,N_23638);
nand U24680 (N_24680,N_20444,N_20021);
or U24681 (N_24681,N_20371,N_23265);
nand U24682 (N_24682,N_18746,N_18956);
nand U24683 (N_24683,N_21092,N_19702);
and U24684 (N_24684,N_18536,N_21816);
and U24685 (N_24685,N_21626,N_21466);
or U24686 (N_24686,N_22646,N_20791);
or U24687 (N_24687,N_21842,N_20887);
nor U24688 (N_24688,N_21213,N_22469);
xor U24689 (N_24689,N_22829,N_22832);
and U24690 (N_24690,N_23652,N_21476);
nand U24691 (N_24691,N_23017,N_19193);
or U24692 (N_24692,N_21615,N_23345);
and U24693 (N_24693,N_20050,N_18041);
xor U24694 (N_24694,N_23929,N_21291);
and U24695 (N_24695,N_21431,N_22698);
nand U24696 (N_24696,N_22405,N_18943);
nand U24697 (N_24697,N_18383,N_23201);
nor U24698 (N_24698,N_18861,N_23594);
and U24699 (N_24699,N_21765,N_23240);
and U24700 (N_24700,N_23164,N_19142);
nor U24701 (N_24701,N_18264,N_22097);
and U24702 (N_24702,N_19482,N_23437);
xor U24703 (N_24703,N_18024,N_22691);
and U24704 (N_24704,N_19131,N_22650);
nand U24705 (N_24705,N_19561,N_18654);
nand U24706 (N_24706,N_20773,N_23070);
nor U24707 (N_24707,N_21988,N_21960);
and U24708 (N_24708,N_20305,N_22886);
nand U24709 (N_24709,N_18715,N_22144);
nand U24710 (N_24710,N_21504,N_23048);
and U24711 (N_24711,N_22034,N_18936);
or U24712 (N_24712,N_18944,N_18617);
nand U24713 (N_24713,N_20469,N_23117);
or U24714 (N_24714,N_23633,N_19097);
or U24715 (N_24715,N_21436,N_19957);
nor U24716 (N_24716,N_19553,N_20405);
nor U24717 (N_24717,N_22369,N_18374);
nor U24718 (N_24718,N_20808,N_19063);
nor U24719 (N_24719,N_23826,N_21346);
nor U24720 (N_24720,N_21412,N_23689);
and U24721 (N_24721,N_19986,N_22798);
nand U24722 (N_24722,N_20751,N_21156);
xor U24723 (N_24723,N_22690,N_19896);
nor U24724 (N_24724,N_20197,N_19888);
or U24725 (N_24725,N_23643,N_23192);
nor U24726 (N_24726,N_23400,N_22491);
xnor U24727 (N_24727,N_23116,N_22783);
or U24728 (N_24728,N_22035,N_22499);
and U24729 (N_24729,N_20415,N_18849);
or U24730 (N_24730,N_22013,N_22393);
and U24731 (N_24731,N_21848,N_19576);
and U24732 (N_24732,N_18316,N_21479);
and U24733 (N_24733,N_19966,N_19328);
or U24734 (N_24734,N_20613,N_20801);
nor U24735 (N_24735,N_19335,N_21564);
and U24736 (N_24736,N_18270,N_19977);
and U24737 (N_24737,N_23293,N_23137);
nor U24738 (N_24738,N_21643,N_21772);
nand U24739 (N_24739,N_19616,N_22335);
nor U24740 (N_24740,N_18208,N_22799);
xnor U24741 (N_24741,N_21692,N_21120);
or U24742 (N_24742,N_20625,N_20309);
nor U24743 (N_24743,N_20117,N_19583);
and U24744 (N_24744,N_21183,N_19850);
or U24745 (N_24745,N_20982,N_18110);
nand U24746 (N_24746,N_21034,N_23077);
xnor U24747 (N_24747,N_23125,N_20830);
nor U24748 (N_24748,N_19901,N_19462);
and U24749 (N_24749,N_20161,N_19794);
nor U24750 (N_24750,N_19618,N_19109);
xnor U24751 (N_24751,N_19357,N_19202);
and U24752 (N_24752,N_20365,N_22391);
nand U24753 (N_24753,N_18379,N_20843);
and U24754 (N_24754,N_23752,N_22264);
xnor U24755 (N_24755,N_18914,N_23010);
nor U24756 (N_24756,N_19568,N_22568);
and U24757 (N_24757,N_18745,N_19634);
nand U24758 (N_24758,N_19107,N_21053);
nand U24759 (N_24759,N_19431,N_20479);
xor U24760 (N_24760,N_19217,N_21847);
nor U24761 (N_24761,N_20869,N_23108);
or U24762 (N_24762,N_19463,N_18779);
or U24763 (N_24763,N_19427,N_18812);
and U24764 (N_24764,N_18454,N_23223);
or U24765 (N_24765,N_20885,N_23639);
or U24766 (N_24766,N_18325,N_23775);
nor U24767 (N_24767,N_21189,N_20369);
nor U24768 (N_24768,N_22492,N_21173);
and U24769 (N_24769,N_22418,N_22776);
or U24770 (N_24770,N_19043,N_20858);
nand U24771 (N_24771,N_22937,N_22148);
and U24772 (N_24772,N_23064,N_22212);
or U24773 (N_24773,N_21920,N_19620);
nand U24774 (N_24774,N_18001,N_22256);
or U24775 (N_24775,N_20193,N_18768);
nand U24776 (N_24776,N_18319,N_22559);
nor U24777 (N_24777,N_18033,N_18411);
nor U24778 (N_24778,N_21000,N_19075);
or U24779 (N_24779,N_23156,N_21908);
and U24780 (N_24780,N_19989,N_21268);
or U24781 (N_24781,N_18520,N_18423);
nor U24782 (N_24782,N_20714,N_23951);
nor U24783 (N_24783,N_20958,N_19198);
or U24784 (N_24784,N_23343,N_22571);
xnor U24785 (N_24785,N_20999,N_22294);
or U24786 (N_24786,N_20582,N_23563);
nand U24787 (N_24787,N_20528,N_19087);
nand U24788 (N_24788,N_18725,N_18356);
nor U24789 (N_24789,N_23279,N_20126);
nor U24790 (N_24790,N_22624,N_18622);
and U24791 (N_24791,N_22982,N_22079);
or U24792 (N_24792,N_22126,N_23675);
nor U24793 (N_24793,N_19106,N_19746);
nor U24794 (N_24794,N_21462,N_21556);
nand U24795 (N_24795,N_23785,N_19115);
or U24796 (N_24796,N_18782,N_23297);
or U24797 (N_24797,N_19607,N_21201);
or U24798 (N_24798,N_18366,N_18834);
nand U24799 (N_24799,N_23475,N_23628);
and U24800 (N_24800,N_22419,N_22589);
nand U24801 (N_24801,N_20435,N_19156);
or U24802 (N_24802,N_22811,N_19274);
xor U24803 (N_24803,N_22608,N_22868);
nand U24804 (N_24804,N_20674,N_21073);
nor U24805 (N_24805,N_23658,N_21191);
or U24806 (N_24806,N_21638,N_18069);
nor U24807 (N_24807,N_22980,N_20856);
or U24808 (N_24808,N_20768,N_21169);
nor U24809 (N_24809,N_18473,N_23998);
nand U24810 (N_24810,N_23358,N_22277);
and U24811 (N_24811,N_18801,N_19410);
and U24812 (N_24812,N_21869,N_19502);
or U24813 (N_24813,N_20373,N_20533);
nor U24814 (N_24814,N_21741,N_21689);
and U24815 (N_24815,N_22056,N_22383);
nor U24816 (N_24816,N_21302,N_20870);
nand U24817 (N_24817,N_20243,N_23690);
xnor U24818 (N_24818,N_18900,N_18738);
or U24819 (N_24819,N_21844,N_22117);
nor U24820 (N_24820,N_23136,N_19598);
xor U24821 (N_24821,N_23710,N_20277);
nand U24822 (N_24822,N_22194,N_21478);
and U24823 (N_24823,N_22959,N_20587);
or U24824 (N_24824,N_20569,N_20211);
and U24825 (N_24825,N_21683,N_23055);
nor U24826 (N_24826,N_23695,N_20114);
or U24827 (N_24827,N_20242,N_18891);
or U24828 (N_24828,N_21575,N_19782);
nor U24829 (N_24829,N_23550,N_20109);
xnor U24830 (N_24830,N_20274,N_19569);
or U24831 (N_24831,N_23283,N_23003);
xnor U24832 (N_24832,N_21813,N_19577);
nor U24833 (N_24833,N_23249,N_23935);
or U24834 (N_24834,N_19991,N_21656);
nand U24835 (N_24835,N_20333,N_21629);
and U24836 (N_24836,N_21251,N_21559);
and U24837 (N_24837,N_18236,N_22354);
nor U24838 (N_24838,N_19460,N_21535);
and U24839 (N_24839,N_22880,N_18154);
and U24840 (N_24840,N_22477,N_21882);
and U24841 (N_24841,N_22042,N_19091);
nor U24842 (N_24842,N_22110,N_18409);
nor U24843 (N_24843,N_23649,N_22882);
nand U24844 (N_24844,N_19371,N_20433);
nor U24845 (N_24845,N_20572,N_18918);
xnor U24846 (N_24846,N_23606,N_18196);
xor U24847 (N_24847,N_23253,N_20120);
xor U24848 (N_24848,N_18002,N_23756);
nand U24849 (N_24849,N_19187,N_18877);
nor U24850 (N_24850,N_19894,N_19392);
nand U24851 (N_24851,N_20575,N_22029);
nor U24852 (N_24852,N_18850,N_19495);
nand U24853 (N_24853,N_19447,N_22146);
and U24854 (N_24854,N_18189,N_21965);
or U24855 (N_24855,N_21236,N_19928);
and U24856 (N_24856,N_20643,N_18702);
or U24857 (N_24857,N_21652,N_21102);
xor U24858 (N_24858,N_21627,N_22037);
or U24859 (N_24859,N_19615,N_21748);
and U24860 (N_24860,N_23654,N_19562);
or U24861 (N_24861,N_19996,N_19235);
xnor U24862 (N_24862,N_23847,N_21194);
nor U24863 (N_24863,N_20698,N_18162);
nand U24864 (N_24864,N_23501,N_20037);
nor U24865 (N_24865,N_21604,N_19563);
or U24866 (N_24866,N_18730,N_23080);
xor U24867 (N_24867,N_21499,N_23500);
or U24868 (N_24868,N_20716,N_21162);
nand U24869 (N_24869,N_18059,N_19228);
or U24870 (N_24870,N_20846,N_20213);
xor U24871 (N_24871,N_23454,N_23290);
nand U24872 (N_24872,N_23158,N_23210);
and U24873 (N_24873,N_21836,N_21989);
or U24874 (N_24874,N_22933,N_19870);
nand U24875 (N_24875,N_21786,N_19625);
and U24876 (N_24876,N_20692,N_20412);
and U24877 (N_24877,N_22819,N_23701);
nor U24878 (N_24878,N_20343,N_20416);
nand U24879 (N_24879,N_21818,N_22898);
and U24880 (N_24880,N_18601,N_23307);
and U24881 (N_24881,N_23367,N_23368);
nor U24882 (N_24882,N_18038,N_21846);
nor U24883 (N_24883,N_20256,N_19045);
and U24884 (N_24884,N_18684,N_23313);
nor U24885 (N_24885,N_21890,N_19910);
nand U24886 (N_24886,N_20493,N_21423);
nand U24887 (N_24887,N_19542,N_18372);
nand U24888 (N_24888,N_22729,N_20729);
nand U24889 (N_24889,N_23049,N_19776);
nor U24890 (N_24890,N_22551,N_20660);
nor U24891 (N_24891,N_20356,N_21668);
nand U24892 (N_24892,N_19744,N_19224);
nor U24893 (N_24893,N_19490,N_22313);
and U24894 (N_24894,N_19612,N_18042);
and U24895 (N_24895,N_23575,N_20046);
nand U24896 (N_24896,N_23584,N_22827);
or U24897 (N_24897,N_19582,N_23856);
nor U24898 (N_24898,N_21896,N_19373);
nor U24899 (N_24899,N_21837,N_20631);
and U24900 (N_24900,N_21303,N_19318);
or U24901 (N_24901,N_23271,N_19236);
nor U24902 (N_24902,N_19081,N_19085);
nand U24903 (N_24903,N_18553,N_23243);
or U24904 (N_24904,N_20173,N_18677);
nor U24905 (N_24905,N_18056,N_22242);
nor U24906 (N_24906,N_19488,N_23024);
or U24907 (N_24907,N_22900,N_23241);
or U24908 (N_24908,N_21322,N_22932);
or U24909 (N_24909,N_19136,N_18701);
and U24910 (N_24910,N_20495,N_18736);
nand U24911 (N_24911,N_18942,N_21418);
and U24912 (N_24912,N_20981,N_18785);
nor U24913 (N_24913,N_23791,N_18972);
and U24914 (N_24914,N_22731,N_20634);
and U24915 (N_24915,N_21320,N_19438);
xnor U24916 (N_24916,N_22316,N_18183);
or U24917 (N_24917,N_22790,N_20606);
or U24918 (N_24918,N_18896,N_18364);
or U24919 (N_24919,N_21525,N_18644);
and U24920 (N_24920,N_20442,N_21587);
nor U24921 (N_24921,N_18460,N_20893);
and U24922 (N_24922,N_19557,N_19510);
and U24923 (N_24923,N_23169,N_22627);
and U24924 (N_24924,N_21353,N_21016);
and U24925 (N_24925,N_20261,N_21404);
nor U24926 (N_24926,N_21516,N_21091);
nor U24927 (N_24927,N_18339,N_19390);
and U24928 (N_24928,N_19672,N_22633);
xnor U24929 (N_24929,N_21147,N_23965);
nor U24930 (N_24930,N_23537,N_20056);
or U24931 (N_24931,N_20576,N_19859);
and U24932 (N_24932,N_19824,N_23100);
and U24933 (N_24933,N_22759,N_19322);
or U24934 (N_24934,N_21586,N_19418);
nand U24935 (N_24935,N_23182,N_19099);
nor U24936 (N_24936,N_19029,N_23212);
nand U24937 (N_24937,N_20515,N_20073);
or U24938 (N_24938,N_21150,N_18641);
nor U24939 (N_24939,N_23406,N_21437);
or U24940 (N_24940,N_19079,N_18286);
nand U24941 (N_24941,N_21159,N_20234);
or U24942 (N_24942,N_23085,N_19489);
nand U24943 (N_24943,N_19547,N_23187);
xnor U24944 (N_24944,N_21690,N_23344);
or U24945 (N_24945,N_22411,N_18704);
or U24946 (N_24946,N_20151,N_23886);
or U24947 (N_24947,N_19757,N_23043);
nand U24948 (N_24948,N_19818,N_18234);
and U24949 (N_24949,N_20206,N_21756);
and U24950 (N_24950,N_21367,N_21510);
and U24951 (N_24951,N_18633,N_18663);
xnor U24952 (N_24952,N_22995,N_19611);
nand U24953 (N_24953,N_22028,N_18656);
and U24954 (N_24954,N_22363,N_20446);
nand U24955 (N_24955,N_20376,N_21870);
nor U24956 (N_24956,N_19434,N_18461);
xor U24957 (N_24957,N_22093,N_18999);
nor U24958 (N_24958,N_22046,N_19983);
nor U24959 (N_24959,N_19025,N_19907);
nor U24960 (N_24960,N_19760,N_21131);
xor U24961 (N_24961,N_20726,N_18789);
or U24962 (N_24962,N_19716,N_23997);
nand U24963 (N_24963,N_18998,N_20571);
nand U24964 (N_24964,N_18171,N_23822);
and U24965 (N_24965,N_21336,N_23773);
nor U24966 (N_24966,N_19342,N_22553);
or U24967 (N_24967,N_22874,N_22084);
and U24968 (N_24968,N_21166,N_20880);
and U24969 (N_24969,N_18138,N_20902);
and U24970 (N_24970,N_20118,N_20834);
and U24971 (N_24971,N_22156,N_23961);
and U24972 (N_24972,N_21608,N_22890);
and U24973 (N_24973,N_21035,N_18934);
or U24974 (N_24974,N_20926,N_23008);
and U24975 (N_24975,N_21107,N_21151);
xor U24976 (N_24976,N_22452,N_18474);
and U24977 (N_24977,N_23157,N_18875);
xor U24978 (N_24978,N_18905,N_22054);
and U24979 (N_24979,N_20028,N_19398);
or U24980 (N_24980,N_19756,N_23704);
xnor U24981 (N_24981,N_21109,N_19349);
and U24982 (N_24982,N_19640,N_20816);
or U24983 (N_24983,N_22245,N_20265);
and U24984 (N_24984,N_23533,N_23390);
xor U24985 (N_24985,N_19190,N_19944);
nor U24986 (N_24986,N_18659,N_21490);
xor U24987 (N_24987,N_21021,N_18971);
nor U24988 (N_24988,N_20833,N_20316);
and U24989 (N_24989,N_23747,N_23019);
nor U24990 (N_24990,N_21163,N_23748);
and U24991 (N_24991,N_22057,N_19103);
and U24992 (N_24992,N_19154,N_22636);
and U24993 (N_24993,N_19411,N_21548);
or U24994 (N_24994,N_23554,N_23384);
nand U24995 (N_24995,N_18163,N_18470);
or U24996 (N_24996,N_23463,N_21075);
nand U24997 (N_24997,N_19070,N_22216);
or U24998 (N_24998,N_18927,N_20732);
nand U24999 (N_24999,N_21362,N_19766);
and U25000 (N_25000,N_18458,N_22851);
or U25001 (N_25001,N_19246,N_19316);
nor U25002 (N_25002,N_20168,N_20809);
nand U25003 (N_25003,N_18452,N_22530);
nor U25004 (N_25004,N_21108,N_22104);
nand U25005 (N_25005,N_18786,N_22090);
nand U25006 (N_25006,N_18151,N_20584);
nand U25007 (N_25007,N_23121,N_18966);
or U25008 (N_25008,N_23672,N_22644);
and U25009 (N_25009,N_18805,N_19668);
nand U25010 (N_25010,N_23110,N_22761);
and U25011 (N_25011,N_19207,N_22448);
and U25012 (N_25012,N_22814,N_19404);
and U25013 (N_25013,N_23938,N_19943);
and U25014 (N_25014,N_22061,N_18735);
nand U25015 (N_25015,N_22733,N_19365);
nand U25016 (N_25016,N_21754,N_22319);
or U25017 (N_25017,N_19694,N_19916);
nor U25018 (N_25018,N_23707,N_18324);
or U25019 (N_25019,N_23421,N_21468);
and U25020 (N_25020,N_22922,N_23733);
or U25021 (N_25021,N_18919,N_18917);
and U25022 (N_25022,N_19074,N_19064);
or U25023 (N_25023,N_18508,N_20344);
nand U25024 (N_25024,N_21498,N_20239);
nor U25025 (N_25025,N_19720,N_18673);
and U25026 (N_25026,N_22380,N_20165);
xor U25027 (N_25027,N_19149,N_20328);
nand U25028 (N_25028,N_18913,N_20649);
and U25029 (N_25029,N_21759,N_19105);
and U25030 (N_25030,N_20505,N_22318);
or U25031 (N_25031,N_19730,N_21807);
or U25032 (N_25032,N_20456,N_19980);
xnor U25033 (N_25033,N_18394,N_22791);
and U25034 (N_25034,N_19402,N_22219);
nand U25035 (N_25035,N_23882,N_22744);
nor U25036 (N_25036,N_19039,N_21824);
or U25037 (N_25037,N_22329,N_20398);
nand U25038 (N_25038,N_19792,N_19909);
or U25039 (N_25039,N_18085,N_18436);
or U25040 (N_25040,N_19920,N_18675);
or U25041 (N_25041,N_18614,N_22763);
nor U25042 (N_25042,N_18197,N_18703);
and U25043 (N_25043,N_19963,N_18714);
or U25044 (N_25044,N_20214,N_18935);
or U25045 (N_25045,N_22342,N_19948);
nor U25046 (N_25046,N_21527,N_21345);
xor U25047 (N_25047,N_23259,N_20176);
or U25048 (N_25048,N_18368,N_21939);
and U25049 (N_25049,N_18734,N_21095);
nand U25050 (N_25050,N_18185,N_18798);
nand U25051 (N_25051,N_18982,N_21459);
xor U25052 (N_25052,N_23656,N_21622);
and U25053 (N_25053,N_20671,N_21198);
and U25054 (N_25054,N_21820,N_18841);
nor U25055 (N_25055,N_19126,N_21849);
nand U25056 (N_25056,N_18139,N_21313);
nor U25057 (N_25057,N_20626,N_18026);
or U25058 (N_25058,N_18502,N_20098);
or U25059 (N_25059,N_18920,N_18229);
or U25060 (N_25060,N_22610,N_23204);
nor U25061 (N_25061,N_19486,N_21078);
and U25062 (N_25062,N_23807,N_22374);
nor U25063 (N_25063,N_22153,N_18413);
or U25064 (N_25064,N_21275,N_22598);
or U25065 (N_25065,N_18773,N_22009);
nor U25066 (N_25066,N_23659,N_18916);
nand U25067 (N_25067,N_18263,N_18602);
or U25068 (N_25068,N_18170,N_22059);
and U25069 (N_25069,N_23536,N_18354);
or U25070 (N_25070,N_18890,N_22236);
and U25071 (N_25071,N_20380,N_23907);
or U25072 (N_25072,N_19339,N_23333);
nand U25073 (N_25073,N_20196,N_19367);
nor U25074 (N_25074,N_18410,N_19869);
and U25075 (N_25075,N_21958,N_22740);
nand U25076 (N_25076,N_18186,N_20813);
nand U25077 (N_25077,N_18243,N_23374);
nand U25078 (N_25078,N_20036,N_22174);
nor U25079 (N_25079,N_22987,N_22098);
or U25080 (N_25080,N_21088,N_19284);
nand U25081 (N_25081,N_23128,N_19877);
or U25082 (N_25082,N_20677,N_18131);
nand U25083 (N_25083,N_23426,N_18571);
and U25084 (N_25084,N_21898,N_22241);
nand U25085 (N_25085,N_20297,N_19773);
nor U25086 (N_25086,N_20718,N_19347);
nor U25087 (N_25087,N_23627,N_22864);
nor U25088 (N_25088,N_18950,N_21184);
nor U25089 (N_25089,N_19886,N_18545);
and U25090 (N_25090,N_19258,N_19163);
nand U25091 (N_25091,N_19942,N_22992);
and U25092 (N_25092,N_19251,N_23122);
nand U25093 (N_25093,N_20003,N_19230);
or U25094 (N_25094,N_18343,N_19769);
nand U25095 (N_25095,N_21925,N_22652);
or U25096 (N_25096,N_21012,N_22066);
nand U25097 (N_25097,N_20436,N_18621);
nor U25098 (N_25098,N_21417,N_23180);
nand U25099 (N_25099,N_19319,N_19821);
nor U25100 (N_25100,N_19846,N_20177);
nor U25101 (N_25101,N_19590,N_22229);
and U25102 (N_25102,N_19377,N_20326);
and U25103 (N_25103,N_22182,N_18122);
or U25104 (N_25104,N_21210,N_21334);
and U25105 (N_25105,N_22588,N_18054);
and U25106 (N_25106,N_22410,N_18671);
nand U25107 (N_25107,N_19780,N_21887);
or U25108 (N_25108,N_23255,N_18153);
xor U25109 (N_25109,N_20324,N_22460);
nor U25110 (N_25110,N_18627,N_19690);
nand U25111 (N_25111,N_18465,N_22253);
nor U25112 (N_25112,N_20031,N_22071);
nand U25113 (N_25113,N_21830,N_19440);
nand U25114 (N_25114,N_21463,N_19208);
nand U25115 (N_25115,N_23516,N_21628);
or U25116 (N_25116,N_21872,N_20012);
and U25117 (N_25117,N_19303,N_21802);
and U25118 (N_25118,N_19736,N_22808);
and U25119 (N_25119,N_21881,N_20681);
nor U25120 (N_25120,N_19687,N_22758);
nand U25121 (N_25121,N_19255,N_19812);
nand U25122 (N_25122,N_19867,N_18108);
xnor U25123 (N_25123,N_19995,N_23099);
xnor U25124 (N_25124,N_19264,N_21204);
and U25125 (N_25125,N_22409,N_23565);
and U25126 (N_25126,N_19020,N_20144);
nand U25127 (N_25127,N_23616,N_22924);
nand U25128 (N_25128,N_18980,N_19803);
and U25129 (N_25129,N_23660,N_19771);
and U25130 (N_25130,N_23000,N_22130);
and U25131 (N_25131,N_18246,N_23526);
nand U25132 (N_25132,N_19800,N_23925);
nor U25133 (N_25133,N_23700,N_21127);
nor U25134 (N_25134,N_23732,N_18957);
and U25135 (N_25135,N_19309,N_21856);
nor U25136 (N_25136,N_22576,N_21582);
or U25137 (N_25137,N_18178,N_21467);
or U25138 (N_25138,N_21980,N_20724);
xor U25139 (N_25139,N_19833,N_18358);
and U25140 (N_25140,N_18961,N_22429);
xnor U25141 (N_25141,N_23674,N_22197);
or U25142 (N_25142,N_19906,N_20555);
or U25143 (N_25143,N_23983,N_22341);
nand U25144 (N_25144,N_20684,N_22359);
and U25145 (N_25145,N_18516,N_19951);
nand U25146 (N_25146,N_23209,N_22843);
nand U25147 (N_25147,N_18297,N_19679);
nor U25148 (N_25148,N_21851,N_23926);
nand U25149 (N_25149,N_23218,N_19353);
and U25150 (N_25150,N_20956,N_20262);
or U25151 (N_25151,N_19416,N_18660);
and U25152 (N_25152,N_19168,N_19127);
nor U25153 (N_25153,N_21294,N_23803);
or U25154 (N_25154,N_20393,N_22180);
nand U25155 (N_25155,N_19465,N_20491);
xnor U25156 (N_25156,N_23890,N_22527);
or U25157 (N_25157,N_21693,N_22281);
nand U25158 (N_25158,N_18282,N_20335);
nand U25159 (N_25159,N_18723,N_21068);
or U25160 (N_25160,N_23120,N_19047);
and U25161 (N_25161,N_21934,N_20156);
and U25162 (N_25162,N_18057,N_19314);
and U25163 (N_25163,N_23287,N_18578);
and U25164 (N_25164,N_20831,N_21845);
and U25165 (N_25165,N_21262,N_21568);
xor U25166 (N_25166,N_22663,N_20873);
nor U25167 (N_25167,N_20879,N_22003);
xor U25168 (N_25168,N_23795,N_21271);
or U25169 (N_25169,N_18889,N_20878);
or U25170 (N_25170,N_23954,N_22478);
and U25171 (N_25171,N_21734,N_18866);
and U25172 (N_25172,N_21530,N_20296);
xor U25173 (N_25173,N_21735,N_19387);
nor U25174 (N_25174,N_22032,N_19002);
and U25175 (N_25175,N_21192,N_20058);
nor U25176 (N_25176,N_20372,N_21926);
or U25177 (N_25177,N_23738,N_18296);
nand U25178 (N_25178,N_21387,N_19518);
and U25179 (N_25179,N_23901,N_22205);
nor U25180 (N_25180,N_22145,N_23050);
nor U25181 (N_25181,N_22719,N_20788);
nor U25182 (N_25182,N_22486,N_19469);
and U25183 (N_25183,N_22231,N_19860);
nor U25184 (N_25184,N_21913,N_20146);
and U25185 (N_25185,N_19759,N_23836);
nor U25186 (N_25186,N_21434,N_22842);
or U25187 (N_25187,N_20832,N_22664);
nor U25188 (N_25188,N_23990,N_19396);
and U25189 (N_25189,N_23485,N_23644);
or U25190 (N_25190,N_20615,N_19570);
nand U25191 (N_25191,N_20201,N_20228);
or U25192 (N_25192,N_18365,N_20018);
nand U25193 (N_25193,N_18241,N_19959);
nand U25194 (N_25194,N_23078,N_21790);
nand U25195 (N_25195,N_18191,N_23481);
nand U25196 (N_25196,N_19879,N_19221);
or U25197 (N_25197,N_20589,N_22122);
and U25198 (N_25198,N_23232,N_20484);
or U25199 (N_25199,N_23394,N_18549);
nand U25200 (N_25200,N_23702,N_20710);
or U25201 (N_25201,N_18637,N_23566);
or U25202 (N_25202,N_22248,N_20178);
xnor U25203 (N_25203,N_22528,N_22063);
or U25204 (N_25204,N_20849,N_22961);
and U25205 (N_25205,N_23724,N_19408);
and U25206 (N_25206,N_21301,N_19033);
xor U25207 (N_25207,N_20220,N_23557);
nand U25208 (N_25208,N_20107,N_20134);
or U25209 (N_25209,N_20514,N_20128);
and U25210 (N_25210,N_19096,N_18347);
nand U25211 (N_25211,N_22166,N_22078);
xor U25212 (N_25212,N_19500,N_19086);
or U25213 (N_25213,N_19786,N_23815);
or U25214 (N_25214,N_23719,N_21795);
nor U25215 (N_25215,N_21744,N_19330);
nor U25216 (N_25216,N_22240,N_18806);
nand U25217 (N_25217,N_18430,N_21160);
nand U25218 (N_25218,N_23877,N_21446);
nand U25219 (N_25219,N_21020,N_23968);
nor U25220 (N_25220,N_23793,N_23023);
nand U25221 (N_25221,N_20527,N_23635);
xor U25222 (N_25222,N_20133,N_19076);
and U25223 (N_25223,N_20995,N_23903);
and U25224 (N_25224,N_20263,N_19137);
or U25225 (N_25225,N_23141,N_19595);
or U25226 (N_25226,N_21506,N_20439);
nor U25227 (N_25227,N_21337,N_19960);
and U25228 (N_25228,N_20160,N_19733);
or U25229 (N_25229,N_22545,N_22768);
or U25230 (N_25230,N_19622,N_18783);
nor U25231 (N_25231,N_18967,N_20970);
nor U25232 (N_25232,N_18992,N_20614);
or U25233 (N_25233,N_23897,N_21895);
nor U25234 (N_25234,N_23484,N_22661);
nor U25235 (N_25235,N_21688,N_21918);
nor U25236 (N_25236,N_19052,N_21180);
and U25237 (N_25237,N_23867,N_23974);
or U25238 (N_25238,N_18795,N_20084);
and U25239 (N_25239,N_23084,N_21269);
nor U25240 (N_25240,N_20357,N_19883);
nor U25241 (N_25241,N_22537,N_22971);
nand U25242 (N_25242,N_20221,N_19586);
nor U25243 (N_25243,N_21821,N_22322);
nand U25244 (N_25244,N_22628,N_23607);
nor U25245 (N_25245,N_22746,N_23599);
or U25246 (N_25246,N_21650,N_21755);
xnor U25247 (N_25247,N_22547,N_23503);
nor U25248 (N_25248,N_21746,N_18023);
and U25249 (N_25249,N_22927,N_22258);
nand U25250 (N_25250,N_20647,N_23631);
nand U25251 (N_25251,N_19820,N_23651);
nand U25252 (N_25252,N_19712,N_18399);
or U25253 (N_25253,N_18032,N_22280);
nand U25254 (N_25254,N_21193,N_21985);
xnor U25255 (N_25255,N_18560,N_20437);
nor U25256 (N_25256,N_23510,N_21834);
and U25257 (N_25257,N_22184,N_23263);
and U25258 (N_25258,N_22916,N_20191);
nor U25259 (N_25259,N_23788,N_21445);
and U25260 (N_25260,N_23754,N_23819);
or U25261 (N_25261,N_23286,N_22654);
nand U25262 (N_25262,N_20785,N_20573);
nor U25263 (N_25263,N_23143,N_23558);
nand U25264 (N_25264,N_20088,N_18434);
xor U25265 (N_25265,N_19710,N_21058);
nand U25266 (N_25266,N_23439,N_22489);
or U25267 (N_25267,N_20500,N_19758);
nor U25268 (N_25268,N_20485,N_22655);
xor U25269 (N_25269,N_18790,N_22333);
and U25270 (N_25270,N_23130,N_22519);
and U25271 (N_25271,N_23885,N_18996);
or U25272 (N_25272,N_21306,N_19636);
and U25273 (N_25273,N_23691,N_19157);
nor U25274 (N_25274,N_21293,N_22472);
xor U25275 (N_25275,N_22585,N_22629);
and U25276 (N_25276,N_19374,N_19053);
xnor U25277 (N_25277,N_23272,N_20113);
nand U25278 (N_25278,N_19515,N_23680);
or U25279 (N_25279,N_19729,N_20635);
or U25280 (N_25280,N_22908,N_18974);
or U25281 (N_25281,N_20311,N_21051);
nor U25282 (N_25282,N_21738,N_22027);
xnor U25283 (N_25283,N_22891,N_21223);
or U25284 (N_25284,N_21415,N_20386);
and U25285 (N_25285,N_18355,N_23380);
nand U25286 (N_25286,N_19062,N_19617);
nand U25287 (N_25287,N_18280,N_20653);
and U25288 (N_25288,N_20186,N_19972);
or U25289 (N_25289,N_23455,N_18160);
xor U25290 (N_25290,N_22965,N_19200);
or U25291 (N_25291,N_20717,N_19994);
or U25292 (N_25292,N_18361,N_20996);
nand U25293 (N_25293,N_23041,N_18469);
nand U25294 (N_25294,N_22626,N_20510);
nand U25295 (N_25295,N_22198,N_19626);
nand U25296 (N_25296,N_19172,N_23600);
nand U25297 (N_25297,N_21248,N_21680);
or U25298 (N_25298,N_22684,N_18651);
nor U25299 (N_25299,N_18167,N_21042);
nand U25300 (N_25300,N_23716,N_23270);
nor U25301 (N_25301,N_23228,N_22825);
nand U25302 (N_25302,N_23088,N_18897);
and U25303 (N_25303,N_22291,N_22070);
nor U25304 (N_25304,N_22945,N_19422);
nand U25305 (N_25305,N_19685,N_21605);
xor U25306 (N_25306,N_22325,N_19343);
nand U25307 (N_25307,N_21128,N_20009);
and U25308 (N_25308,N_20387,N_19185);
nor U25309 (N_25309,N_22428,N_19619);
nor U25310 (N_25310,N_19755,N_23632);
nor U25311 (N_25311,N_20554,N_18086);
nand U25312 (N_25312,N_20190,N_23519);
and U25313 (N_25313,N_22706,N_20721);
or U25314 (N_25314,N_23027,N_22998);
and U25315 (N_25315,N_22361,N_23465);
and U25316 (N_25316,N_18490,N_19739);
nor U25317 (N_25317,N_23031,N_21933);
nor U25318 (N_25318,N_20321,N_22885);
nand U25319 (N_25319,N_21721,N_23295);
nand U25320 (N_25320,N_23337,N_20127);
nor U25321 (N_25321,N_20092,N_22844);
nand U25322 (N_25322,N_19704,N_23054);
or U25323 (N_25323,N_23784,N_21949);
and U25324 (N_25324,N_19578,N_18148);
or U25325 (N_25325,N_20068,N_19554);
nand U25326 (N_25326,N_20122,N_19042);
or U25327 (N_25327,N_23268,N_19394);
nor U25328 (N_25328,N_20198,N_22445);
or U25329 (N_25329,N_20921,N_22422);
or U25330 (N_25330,N_21245,N_22592);
nor U25331 (N_25331,N_19748,N_22467);
and U25332 (N_25332,N_23963,N_18740);
and U25333 (N_25333,N_23553,N_23608);
and U25334 (N_25334,N_19051,N_23222);
nor U25335 (N_25335,N_18607,N_18157);
nor U25336 (N_25336,N_23648,N_22672);
or U25337 (N_25337,N_20322,N_21880);
nand U25338 (N_25338,N_19241,N_21637);
nor U25339 (N_25339,N_22803,N_19589);
or U25340 (N_25340,N_22372,N_22196);
nand U25341 (N_25341,N_22210,N_18676);
xor U25342 (N_25342,N_22444,N_23412);
xor U25343 (N_25343,N_22720,N_18260);
and U25344 (N_25344,N_20603,N_18753);
xor U25345 (N_25345,N_21858,N_23758);
or U25346 (N_25346,N_23580,N_19982);
or U25347 (N_25347,N_23460,N_21777);
nand U25348 (N_25348,N_19299,N_21257);
and U25349 (N_25349,N_23778,N_18344);
nor U25350 (N_25350,N_23978,N_21475);
nor U25351 (N_25351,N_23620,N_18979);
or U25352 (N_25352,N_18886,N_20617);
nor U25353 (N_25353,N_23532,N_22847);
and U25354 (N_25354,N_18290,N_19603);
and U25355 (N_25355,N_18305,N_20836);
nand U25356 (N_25356,N_21007,N_21750);
nor U25357 (N_25357,N_22096,N_21339);
and U25358 (N_25358,N_23131,N_18493);
and U25359 (N_25359,N_20188,N_21328);
or U25360 (N_25360,N_20526,N_21460);
and U25361 (N_25361,N_18438,N_21408);
xor U25362 (N_25362,N_21155,N_19934);
nand U25363 (N_25363,N_21630,N_22051);
nor U25364 (N_25364,N_22558,N_20022);
nor U25365 (N_25365,N_22502,N_18462);
nor U25366 (N_25366,N_23868,N_22514);
or U25367 (N_25367,N_18390,N_20171);
nor U25368 (N_25368,N_18767,N_21001);
or U25369 (N_25369,N_20308,N_23991);
nand U25370 (N_25370,N_19148,N_19750);
nand U25371 (N_25371,N_18503,N_19908);
or U25372 (N_25372,N_20583,N_22150);
and U25373 (N_25373,N_20385,N_23073);
or U25374 (N_25374,N_18327,N_20325);
nor U25375 (N_25375,N_22967,N_22077);
or U25376 (N_25376,N_20411,N_18375);
nand U25377 (N_25377,N_21196,N_18166);
or U25378 (N_25378,N_19292,N_21171);
nand U25379 (N_25379,N_19356,N_20210);
and U25380 (N_25380,N_21540,N_18652);
nand U25381 (N_25381,N_20358,N_23982);
nor U25382 (N_25382,N_19721,N_21747);
or U25383 (N_25383,N_23636,N_21428);
and U25384 (N_25384,N_23044,N_19334);
xor U25385 (N_25385,N_18726,N_20246);
and U25386 (N_25386,N_19521,N_22910);
or U25387 (N_25387,N_22370,N_22762);
nand U25388 (N_25388,N_22899,N_19271);
or U25389 (N_25389,N_23873,N_22123);
or U25390 (N_25390,N_22949,N_18822);
nor U25391 (N_25391,N_19958,N_22968);
xor U25392 (N_25392,N_23771,N_18965);
nor U25393 (N_25393,N_21946,N_20406);
nand U25394 (N_25394,N_22804,N_22008);
nand U25395 (N_25395,N_20598,N_18392);
and U25396 (N_25396,N_18873,N_20391);
nor U25397 (N_25397,N_20725,N_22779);
or U25398 (N_25398,N_20787,N_20702);
or U25399 (N_25399,N_18883,N_21517);
nand U25400 (N_25400,N_19205,N_20438);
nand U25401 (N_25401,N_22279,N_19581);
and U25402 (N_25402,N_20906,N_20517);
and U25403 (N_25403,N_18223,N_20215);
nand U25404 (N_25404,N_22869,N_20450);
nand U25405 (N_25405,N_21696,N_20153);
xnor U25406 (N_25406,N_18501,N_21125);
xnor U25407 (N_25407,N_18391,N_23033);
nor U25408 (N_25408,N_21952,N_23324);
and U25409 (N_25409,N_20503,N_22234);
xor U25410 (N_25410,N_22015,N_23378);
nor U25411 (N_25411,N_21730,N_19215);
or U25412 (N_25412,N_21308,N_22430);
nand U25413 (N_25413,N_21655,N_19135);
nor U25414 (N_25414,N_23058,N_22510);
and U25415 (N_25415,N_23020,N_20025);
or U25416 (N_25416,N_18672,N_21664);
nor U25417 (N_25417,N_18418,N_21961);
or U25418 (N_25418,N_22960,N_22800);
nor U25419 (N_25419,N_21174,N_18288);
nor U25420 (N_25420,N_18880,N_21623);
nand U25421 (N_25421,N_19278,N_18681);
nor U25422 (N_25422,N_22917,N_22207);
nand U25423 (N_25423,N_23291,N_20616);
nor U25424 (N_25424,N_23679,N_18985);
nor U25425 (N_25425,N_20466,N_21819);
xor U25426 (N_25426,N_23004,N_23257);
and U25427 (N_25427,N_18846,N_20402);
nand U25428 (N_25428,N_21959,N_23056);
or U25429 (N_25429,N_19675,N_22047);
or U25430 (N_25430,N_18749,N_18885);
and U25431 (N_25431,N_21148,N_20379);
and U25432 (N_25432,N_23140,N_22225);
or U25433 (N_25433,N_18464,N_21828);
nor U25434 (N_25434,N_23149,N_22637);
xor U25435 (N_25435,N_20594,N_23015);
and U25436 (N_25436,N_19012,N_21609);
nor U25437 (N_25437,N_22237,N_20455);
nand U25438 (N_25438,N_20330,N_23422);
or U25439 (N_25439,N_20460,N_20518);
nor U25440 (N_25440,N_22261,N_21561);
and U25441 (N_25441,N_20038,N_21230);
and U25442 (N_25442,N_18053,N_23096);
and U25443 (N_25443,N_23711,N_18583);
nor U25444 (N_25444,N_20559,N_20610);
or U25445 (N_25445,N_23718,N_21502);
or U25446 (N_25446,N_23987,N_21032);
or U25447 (N_25447,N_22830,N_22722);
or U25448 (N_25448,N_20351,N_20494);
and U25449 (N_25449,N_20273,N_20388);
or U25450 (N_25450,N_20255,N_20777);
or U25451 (N_25451,N_21572,N_23289);
nor U25452 (N_25452,N_20588,N_18068);
and U25453 (N_25453,N_22019,N_22556);
nand U25454 (N_25454,N_18052,N_18529);
nor U25455 (N_25455,N_19242,N_20291);
nand U25456 (N_25456,N_23804,N_19428);
nor U25457 (N_25457,N_23583,N_19533);
xnor U25458 (N_25458,N_18855,N_23520);
nand U25459 (N_25459,N_18124,N_22493);
nor U25460 (N_25460,N_21433,N_19363);
and U25461 (N_25461,N_19706,N_23436);
and U25462 (N_25462,N_19885,N_21524);
and U25463 (N_25463,N_18968,N_21190);
or U25464 (N_25464,N_21278,N_21219);
and U25465 (N_25465,N_19360,N_20953);
nand U25466 (N_25466,N_21814,N_19225);
and U25467 (N_25467,N_20342,N_18232);
or U25468 (N_25468,N_18776,N_23018);
nand U25469 (N_25469,N_18689,N_21292);
and U25470 (N_25470,N_22723,N_22362);
nand U25471 (N_25471,N_20850,N_21775);
or U25472 (N_25472,N_18156,N_18134);
or U25473 (N_25473,N_20070,N_19346);
and U25474 (N_25474,N_19811,N_20633);
or U25475 (N_25475,N_22969,N_19884);
nand U25476 (N_25476,N_19714,N_23912);
nor U25477 (N_25477,N_19503,N_22187);
nor U25478 (N_25478,N_18204,N_18509);
and U25479 (N_25479,N_21619,N_22662);
nor U25480 (N_25480,N_18542,N_20378);
nand U25481 (N_25481,N_19110,N_18825);
nor U25482 (N_25482,N_19539,N_22425);
nand U25483 (N_25483,N_22454,N_20794);
or U25484 (N_25484,N_22751,N_18333);
xnor U25485 (N_25485,N_20852,N_18665);
or U25486 (N_25486,N_22382,N_19132);
or U25487 (N_25487,N_20066,N_19133);
or U25488 (N_25488,N_23546,N_22293);
and U25489 (N_25489,N_19707,N_19183);
nand U25490 (N_25490,N_22487,N_22120);
and U25491 (N_25491,N_20600,N_22328);
xnor U25492 (N_25492,N_21929,N_18862);
xnor U25493 (N_25493,N_23273,N_20731);
or U25494 (N_25494,N_18442,N_23445);
xnor U25495 (N_25495,N_21487,N_23619);
xnor U25496 (N_25496,N_23153,N_20204);
xnor U25497 (N_25497,N_23301,N_23389);
and U25498 (N_25498,N_21327,N_20991);
nand U25499 (N_25499,N_19203,N_23895);
and U25500 (N_25500,N_21532,N_18599);
and U25501 (N_25501,N_19835,N_21398);
xnor U25502 (N_25502,N_18035,N_23013);
nor U25503 (N_25503,N_23190,N_21218);
nor U25504 (N_25504,N_23242,N_21260);
nand U25505 (N_25505,N_19130,N_19444);
nand U25506 (N_25506,N_19566,N_22775);
nor U25507 (N_25507,N_19642,N_20345);
and U25508 (N_25508,N_19768,N_21511);
nand U25509 (N_25509,N_22470,N_22227);
and U25510 (N_25510,N_23362,N_21273);
nor U25511 (N_25511,N_23927,N_22991);
xnor U25512 (N_25512,N_18105,N_22400);
nor U25513 (N_25513,N_18248,N_19930);
nor U25514 (N_25514,N_22704,N_19391);
and U25515 (N_25515,N_23491,N_22712);
xor U25516 (N_25516,N_18537,N_19819);
nand U25517 (N_25517,N_18210,N_21401);
or U25518 (N_25518,N_22839,N_22327);
xnor U25519 (N_25519,N_20182,N_19128);
nand U25520 (N_25520,N_21761,N_21591);
and U25521 (N_25521,N_23407,N_21377);
or U25522 (N_25522,N_21481,N_19049);
and U25523 (N_25523,N_18713,N_18381);
nor U25524 (N_25524,N_19955,N_23835);
xor U25525 (N_25525,N_18450,N_22903);
nor U25526 (N_25526,N_19026,N_22850);
nand U25527 (N_25527,N_20400,N_19584);
or U25528 (N_25528,N_20621,N_20910);
nand U25529 (N_25529,N_19277,N_20150);
and U25530 (N_25530,N_20430,N_18680);
nor U25531 (N_25531,N_21310,N_20015);
nand U25532 (N_25532,N_23083,N_22781);
or U25533 (N_25533,N_20712,N_22795);
or U25534 (N_25534,N_22000,N_18494);
or U25535 (N_25535,N_22250,N_22022);
or U25536 (N_25536,N_19865,N_22544);
nor U25537 (N_25537,N_18181,N_18329);
or U25538 (N_25538,N_21667,N_19487);
nand U25539 (N_25539,N_20898,N_18369);
xnor U25540 (N_25540,N_21321,N_22902);
and U25541 (N_25541,N_22734,N_20279);
and U25542 (N_25542,N_19666,N_19935);
or U25543 (N_25543,N_18800,N_20250);
xnor U25544 (N_25544,N_19243,N_20507);
or U25545 (N_25545,N_22026,N_18851);
xor U25546 (N_25546,N_18083,N_18945);
and U25547 (N_25547,N_19808,N_21074);
or U25548 (N_25548,N_22086,N_19001);
nand U25549 (N_25549,N_19341,N_22314);
nor U25550 (N_25550,N_22632,N_18948);
nor U25551 (N_25551,N_19509,N_18937);
nand U25552 (N_25552,N_22560,N_22392);
or U25553 (N_25553,N_21409,N_20086);
and U25554 (N_25554,N_21817,N_23779);
xor U25555 (N_25555,N_22011,N_22862);
xnor U25556 (N_25556,N_18727,N_23089);
and U25557 (N_25557,N_18235,N_22892);
or U25558 (N_25558,N_19351,N_22025);
nand U25559 (N_25559,N_21826,N_23893);
or U25560 (N_25560,N_18019,N_23303);
and U25561 (N_25561,N_20930,N_20452);
and U25562 (N_25562,N_18762,N_22764);
or U25563 (N_25563,N_19485,N_22935);
xnor U25564 (N_25564,N_20551,N_18093);
nand U25565 (N_25565,N_21861,N_19496);
nand U25566 (N_25566,N_18639,N_20172);
and U25567 (N_25567,N_18804,N_20472);
and U25568 (N_25568,N_18352,N_22905);
and U25569 (N_25569,N_18312,N_19659);
or U25570 (N_25570,N_23166,N_19003);
and U25571 (N_25571,N_23762,N_20864);
or U25572 (N_25572,N_18330,N_23828);
nor U25573 (N_25573,N_19604,N_18380);
nor U25574 (N_25574,N_23757,N_18194);
or U25575 (N_25575,N_21145,N_22331);
nor U25576 (N_25576,N_21968,N_18200);
or U25577 (N_25577,N_22390,N_19275);
or U25578 (N_25578,N_22594,N_22177);
xor U25579 (N_25579,N_22555,N_18499);
nand U25580 (N_25580,N_20532,N_23676);
and U25581 (N_25581,N_19433,N_19549);
and U25582 (N_25582,N_21112,N_23831);
nand U25583 (N_25583,N_23447,N_18824);
or U25584 (N_25584,N_23571,N_18414);
nor U25585 (N_25585,N_21011,N_19947);
and U25586 (N_25586,N_23278,N_22062);
nand U25587 (N_25587,N_20185,N_22213);
xnor U25588 (N_25588,N_23708,N_22845);
xnor U25589 (N_25589,N_19897,N_23392);
and U25590 (N_25590,N_18925,N_23355);
and U25591 (N_25591,N_23206,N_18827);
and U25592 (N_25592,N_23352,N_18488);
and U25593 (N_25593,N_23427,N_18513);
or U25594 (N_25594,N_21955,N_20599);
and U25595 (N_25595,N_19201,N_22175);
xor U25596 (N_25596,N_20200,N_22075);
and U25597 (N_25597,N_21136,N_19421);
and U25598 (N_25598,N_18687,N_19104);
xnor U25599 (N_25599,N_22736,N_21253);
nand U25600 (N_25600,N_19437,N_19456);
and U25601 (N_25601,N_21424,N_18321);
nand U25602 (N_25602,N_22315,N_19565);
or U25603 (N_25603,N_22855,N_18813);
nor U25604 (N_25604,N_20881,N_23547);
nor U25605 (N_25605,N_19732,N_20302);
nand U25606 (N_25606,N_22630,N_19610);
nor U25607 (N_25607,N_20513,N_23097);
and U25608 (N_25608,N_23184,N_20278);
nor U25609 (N_25609,N_21063,N_18255);
nand U25610 (N_25610,N_23613,N_23177);
or U25611 (N_25611,N_21486,N_22671);
nand U25612 (N_25612,N_23781,N_20091);
nor U25613 (N_25613,N_20811,N_20090);
nor U25614 (N_25614,N_19301,N_19637);
and U25615 (N_25615,N_21852,N_22603);
nor U25616 (N_25616,N_21244,N_23432);
nand U25617 (N_25617,N_19386,N_21576);
and U25618 (N_25618,N_23816,N_21070);
or U25619 (N_25619,N_21096,N_18780);
or U25620 (N_25620,N_23923,N_18443);
or U25621 (N_25621,N_23208,N_19508);
nand U25622 (N_25622,N_23314,N_22131);
nand U25623 (N_25623,N_23142,N_21752);
nand U25624 (N_25624,N_19936,N_20071);
and U25625 (N_25625,N_19286,N_18721);
or U25626 (N_25626,N_23495,N_20859);
xnor U25627 (N_25627,N_22356,N_18281);
nand U25628 (N_25628,N_18018,N_19358);
xnor U25629 (N_25629,N_20096,N_23948);
or U25630 (N_25630,N_20410,N_22285);
nand U25631 (N_25631,N_21707,N_23764);
or U25632 (N_25632,N_19145,N_23361);
and U25633 (N_25633,N_20568,N_23504);
and U25634 (N_25634,N_21427,N_22936);
and U25635 (N_25635,N_18642,N_21914);
nor U25636 (N_25636,N_22615,N_20754);
and U25637 (N_25637,N_20668,N_18203);
xor U25638 (N_25638,N_20100,N_22912);
nand U25639 (N_25639,N_21274,N_23860);
nand U25640 (N_25640,N_19806,N_23588);
and U25641 (N_25641,N_19213,N_23883);
nor U25642 (N_25642,N_20723,N_18070);
nor U25643 (N_25643,N_23878,N_22743);
xnor U25644 (N_25644,N_23734,N_18901);
nand U25645 (N_25645,N_19764,N_21393);
or U25646 (N_25646,N_19681,N_18524);
and U25647 (N_25647,N_20844,N_19670);
xnor U25648 (N_25648,N_22765,N_18497);
and U25649 (N_25649,N_23062,N_22494);
or U25650 (N_25650,N_22048,N_20258);
nand U25651 (N_25651,N_20314,N_20672);
or U25652 (N_25652,N_21715,N_20644);
nand U25653 (N_25653,N_20298,N_20818);
nor U25654 (N_25654,N_23561,N_22232);
and U25655 (N_25655,N_22517,N_19534);
or U25656 (N_25656,N_23349,N_20260);
or U25657 (N_25657,N_21871,N_22870);
nor U25658 (N_25658,N_20980,N_23681);
or U25659 (N_25659,N_19093,N_19639);
nand U25660 (N_25660,N_22596,N_22725);
and U25661 (N_25661,N_19027,N_18395);
or U25662 (N_25662,N_21943,N_20937);
nor U25663 (N_25663,N_18857,N_19911);
nor U25664 (N_25664,N_19388,N_18214);
nor U25665 (N_25665,N_20916,N_23330);
xnor U25666 (N_25666,N_19664,N_18815);
nor U25667 (N_25667,N_23105,N_23851);
nor U25668 (N_25668,N_21441,N_22049);
or U25669 (N_25669,N_22255,N_18793);
nor U25670 (N_25670,N_23178,N_23087);
or U25671 (N_25671,N_18960,N_19378);
nand U25672 (N_25672,N_19858,N_18031);
nor U25673 (N_25673,N_23843,N_22305);
nand U25674 (N_25674,N_18870,N_18121);
xnor U25675 (N_25675,N_18039,N_19267);
or U25676 (N_25676,N_20124,N_20254);
nor U25677 (N_25677,N_18449,N_23918);
nor U25678 (N_25678,N_22119,N_19459);
and U25679 (N_25679,N_22641,N_21701);
and U25680 (N_25680,N_22399,N_20420);
or U25681 (N_25681,N_22168,N_18350);
nor U25682 (N_25682,N_23090,N_20964);
xor U25683 (N_25683,N_20023,N_22414);
nand U25684 (N_25684,N_20271,N_18426);
and U25685 (N_25685,N_19655,N_18910);
nand U25686 (N_25686,N_20786,N_19899);
and U25687 (N_25687,N_19711,N_22407);
or U25688 (N_25688,N_18928,N_22821);
and U25689 (N_25689,N_23994,N_21438);
nor U25690 (N_25690,N_18765,N_23787);
xnor U25691 (N_25691,N_18199,N_20840);
nand U25692 (N_25692,N_20301,N_23489);
or U25693 (N_25693,N_20132,N_21984);
nand U25694 (N_25694,N_23946,N_23026);
nand U25695 (N_25695,N_19072,N_23591);
nand U25696 (N_25696,N_21440,N_21978);
nand U25697 (N_25697,N_21399,N_21371);
nor U25698 (N_25698,N_18576,N_20448);
xnor U25699 (N_25699,N_22172,N_19407);
or U25700 (N_25700,N_18037,N_18853);
or U25701 (N_25701,N_19307,N_19094);
nand U25702 (N_25702,N_19348,N_20268);
nand U25703 (N_25703,N_21290,N_18775);
nor U25704 (N_25704,N_20231,N_20499);
nand U25705 (N_25705,N_19108,N_23098);
or U25706 (N_25706,N_23634,N_21823);
nand U25707 (N_25707,N_20492,N_21085);
and U25708 (N_25708,N_18527,N_18661);
and U25709 (N_25709,N_19272,N_20867);
nand U25710 (N_25710,N_18951,N_23298);
and U25711 (N_25711,N_19953,N_22272);
and U25712 (N_25712,N_23840,N_18206);
xnor U25713 (N_25713,N_20512,N_20248);
nand U25714 (N_25714,N_18635,N_20399);
nor U25715 (N_25715,N_19111,N_18921);
or U25716 (N_25716,N_23276,N_19974);
nor U25717 (N_25717,N_23334,N_22265);
nor U25718 (N_25718,N_23813,N_20509);
or U25719 (N_25719,N_18340,N_22735);
or U25720 (N_25720,N_22697,N_21865);
nor U25721 (N_25721,N_18611,N_18304);
xnor U25722 (N_25722,N_19288,N_22259);
and U25723 (N_25723,N_19677,N_20315);
nor U25724 (N_25724,N_19260,N_20667);
xor U25725 (N_25725,N_20942,N_23609);
nand U25726 (N_25726,N_21461,N_18619);
and U25727 (N_25727,N_22909,N_23225);
nor U25728 (N_25728,N_18733,N_21601);
or U25729 (N_25729,N_21551,N_22094);
xnor U25730 (N_25730,N_22017,N_22718);
and U25731 (N_25731,N_19171,N_23194);
or U25732 (N_25732,N_18739,N_23726);
nand U25733 (N_25733,N_19834,N_23379);
nand U25734 (N_25734,N_22462,N_19405);
and U25735 (N_25735,N_19098,N_21388);
xnor U25736 (N_25736,N_23397,N_23859);
and U25737 (N_25737,N_21932,N_23235);
nor U25738 (N_25738,N_18010,N_19715);
and U25739 (N_25739,N_18371,N_21312);
nor U25740 (N_25740,N_21396,N_21536);
nand U25741 (N_25741,N_23593,N_18624);
nor U25742 (N_25742,N_23312,N_19014);
nor U25743 (N_25743,N_18865,N_21175);
nor U25744 (N_25744,N_20976,N_22233);
or U25745 (N_25745,N_21557,N_23134);
xnor U25746 (N_25746,N_20194,N_20896);
nor U25747 (N_25747,N_20203,N_19925);
xor U25748 (N_25748,N_20795,N_18306);
nand U25749 (N_25749,N_21518,N_20478);
xor U25750 (N_25750,N_21990,N_18120);
xnor U25751 (N_25751,N_22934,N_22836);
nor U25752 (N_25752,N_20202,N_22947);
and U25753 (N_25753,N_23322,N_19719);
and U25754 (N_25754,N_20110,N_19742);
nand U25755 (N_25755,N_22640,N_19749);
nor U25756 (N_25756,N_23543,N_23829);
and U25757 (N_25757,N_20947,N_23234);
nand U25758 (N_25758,N_19840,N_20669);
and U25759 (N_25759,N_21728,N_19575);
and U25760 (N_25760,N_22879,N_19663);
nand U25761 (N_25761,N_20580,N_22609);
and U25762 (N_25762,N_22742,N_21935);
nor U25763 (N_25763,N_23165,N_23229);
xor U25764 (N_25764,N_19864,N_21304);
or U25765 (N_25765,N_18803,N_20530);
nor U25766 (N_25766,N_18284,N_21220);
and U25767 (N_25767,N_23339,N_22106);
and U25768 (N_25768,N_21425,N_20157);
and U25769 (N_25769,N_21521,N_22092);
nand U25770 (N_25770,N_19206,N_21233);
nor U25771 (N_25771,N_20637,N_20340);
or U25772 (N_25772,N_23802,N_18012);
nand U25773 (N_25773,N_20252,N_23818);
and U25774 (N_25774,N_18274,N_22760);
nand U25775 (N_25775,N_19199,N_23375);
nand U25776 (N_25776,N_21358,N_22732);
nor U25777 (N_25777,N_23683,N_22055);
and U25778 (N_25778,N_20822,N_19121);
nor U25779 (N_25779,N_18291,N_22449);
xor U25780 (N_25780,N_19289,N_20950);
nor U25781 (N_25781,N_23958,N_21299);
xor U25782 (N_25782,N_23328,N_20374);
nor U25783 (N_25783,N_20891,N_22943);
or U25784 (N_25784,N_23319,N_20770);
or U25785 (N_25785,N_21940,N_19882);
and U25786 (N_25786,N_21212,N_18253);
or U25787 (N_25787,N_23226,N_22490);
or U25788 (N_25788,N_21181,N_18796);
nor U25789 (N_25789,N_22176,N_20948);
or U25790 (N_25790,N_23641,N_22696);
nor U25791 (N_25791,N_20317,N_20945);
nor U25792 (N_25792,N_19967,N_21987);
nor U25793 (N_25793,N_18359,N_23955);
or U25794 (N_25794,N_23549,N_23443);
and U25795 (N_25795,N_19676,N_21277);
nand U25796 (N_25796,N_19247,N_20601);
and U25797 (N_25797,N_21868,N_20561);
nand U25798 (N_25798,N_21716,N_19088);
or U25799 (N_25799,N_23466,N_22703);
nor U25800 (N_25800,N_20565,N_22387);
and U25801 (N_25801,N_20892,N_20524);
nand U25802 (N_25802,N_19209,N_22427);
and U25803 (N_25803,N_20685,N_20303);
and U25804 (N_25804,N_18958,N_21799);
or U25805 (N_25805,N_23664,N_19684);
nor U25806 (N_25806,N_20424,N_19517);
nor U25807 (N_25807,N_22872,N_19924);
and U25808 (N_25808,N_19429,N_22191);
nand U25809 (N_25809,N_21234,N_21179);
nand U25810 (N_25810,N_20884,N_19671);
nor U25811 (N_25811,N_22581,N_21247);
nand U25812 (N_25812,N_20862,N_20596);
nor U25813 (N_25813,N_19216,N_19336);
and U25814 (N_25814,N_18127,N_19970);
nor U25815 (N_25815,N_22160,N_21134);
or U25816 (N_25816,N_20137,N_23611);
nor U25817 (N_25817,N_21342,N_21207);
or U25818 (N_25818,N_21974,N_22944);
and U25819 (N_25819,N_20057,N_19693);
nor U25820 (N_25820,N_18207,N_18060);
nand U25821 (N_25821,N_22873,N_20209);
nor U25822 (N_25822,N_20232,N_21261);
nand U25823 (N_25823,N_23869,N_22816);
nand U25824 (N_25824,N_23906,N_23028);
and U25825 (N_25825,N_19624,N_20367);
nand U25826 (N_25826,N_22823,N_18929);
and U25827 (N_25827,N_21544,N_18709);
and U25828 (N_25828,N_23396,N_23744);
nand U25829 (N_25829,N_23865,N_22946);
or U25830 (N_25830,N_20696,N_22852);
and U25831 (N_25831,N_18694,N_21208);
or U25832 (N_25832,N_22887,N_18118);
and U25833 (N_25833,N_21782,N_23703);
nor U25834 (N_25834,N_20629,N_18342);
xor U25835 (N_25835,N_19629,N_19527);
or U25836 (N_25836,N_19873,N_20363);
or U25837 (N_25837,N_20283,N_22705);
and U25838 (N_25838,N_20960,N_20249);
nor U25839 (N_25839,N_23039,N_22966);
nand U25840 (N_25840,N_19887,N_18294);
or U25841 (N_25841,N_18514,N_19968);
nor U25842 (N_25842,N_19593,N_19413);
nor U25843 (N_25843,N_18328,N_20675);
nand U25844 (N_25844,N_20468,N_19724);
nand U25845 (N_25845,N_21335,N_22014);
and U25846 (N_25846,N_20730,N_19090);
xor U25847 (N_25847,N_18102,N_22929);
nor U25848 (N_25848,N_19722,N_21132);
and U25849 (N_25849,N_23743,N_21522);
and U25850 (N_25850,N_19118,N_23562);
nand U25851 (N_25851,N_19727,N_23402);
and U25852 (N_25852,N_18620,N_21331);
nand U25853 (N_25853,N_18267,N_23949);
and U25854 (N_25854,N_22687,N_20697);
xor U25855 (N_25855,N_23403,N_21917);
or U25856 (N_25856,N_23051,N_20065);
and U25857 (N_25857,N_23038,N_18216);
xnor U25858 (N_25858,N_23320,N_22665);
and U25859 (N_25859,N_21942,N_22838);
nand U25860 (N_25860,N_20483,N_18132);
nor U25861 (N_25861,N_19211,N_22894);
nand U25862 (N_25862,N_20010,N_22579);
and U25863 (N_25863,N_22420,N_23036);
or U25864 (N_25864,N_21770,N_23981);
and U25865 (N_25865,N_22895,N_19571);
nand U25866 (N_25866,N_23741,N_21843);
and U25867 (N_25867,N_18523,N_18912);
and U25868 (N_25868,N_20476,N_18177);
nand U25869 (N_25869,N_18174,N_21298);
or U25870 (N_25870,N_18401,N_22683);
and U25871 (N_25871,N_23252,N_18874);
nand U25872 (N_25872,N_23530,N_22918);
and U25873 (N_25873,N_22496,N_19280);
or U25874 (N_25874,N_19809,N_22713);
nand U25875 (N_25875,N_18129,N_19166);
nor U25876 (N_25876,N_22591,N_18674);
nand U25877 (N_25877,N_18864,N_18145);
or U25878 (N_25878,N_23753,N_19914);
or U25879 (N_25879,N_20547,N_23892);
xor U25880 (N_25880,N_22474,N_19031);
or U25881 (N_25881,N_23682,N_23827);
or U25882 (N_25882,N_21139,N_20623);
nand U25883 (N_25883,N_19520,N_20940);
nor U25884 (N_25884,N_18341,N_18386);
xor U25885 (N_25885,N_20952,N_23176);
nand U25886 (N_25886,N_20282,N_23941);
and U25887 (N_25887,N_20701,N_22572);
or U25888 (N_25888,N_21483,N_21732);
or U25889 (N_25889,N_18218,N_22667);
or U25890 (N_25890,N_21964,N_22169);
nor U25891 (N_25891,N_18887,N_19245);
or U25892 (N_25892,N_18699,N_23508);
nand U25893 (N_25893,N_23267,N_19667);
and U25894 (N_25894,N_20765,N_19100);
or U25895 (N_25895,N_20861,N_23074);
xor U25896 (N_25896,N_21712,N_21374);
nand U25897 (N_25897,N_18396,N_19613);
and U25898 (N_25898,N_22484,N_21141);
xnor U25899 (N_25899,N_20939,N_18303);
or U25900 (N_25900,N_18832,N_23011);
or U25901 (N_25901,N_22750,N_23920);
xor U25902 (N_25902,N_20490,N_22208);
and U25903 (N_25903,N_21123,N_21703);
nor U25904 (N_25904,N_20225,N_23673);
nor U25905 (N_25905,N_20155,N_20067);
or U25906 (N_25906,N_23256,N_22345);
and U25907 (N_25907,N_18009,N_23219);
nor U25908 (N_25908,N_21739,N_22593);
nand U25909 (N_25909,N_21505,N_22195);
xor U25910 (N_25910,N_23902,N_18048);
xor U25911 (N_25911,N_19805,N_20695);
nand U25912 (N_25912,N_19532,N_22297);
and U25913 (N_25913,N_23989,N_20619);
nor U25914 (N_25914,N_23662,N_22863);
nand U25915 (N_25915,N_20889,N_23922);
nor U25916 (N_25916,N_21563,N_22618);
xor U25917 (N_25917,N_18628,N_22792);
nand U25918 (N_25918,N_19735,N_19169);
xor U25919 (N_25919,N_22532,N_22782);
or U25920 (N_25920,N_18249,N_20848);
nor U25921 (N_25921,N_19770,N_19282);
xor U25922 (N_25922,N_20280,N_18831);
nor U25923 (N_25923,N_18320,N_18407);
nand U25924 (N_25924,N_20119,N_21736);
and U25925 (N_25925,N_23506,N_23577);
xor U25926 (N_25926,N_21185,N_22831);
nor U25927 (N_25927,N_22997,N_21705);
and U25928 (N_25928,N_22957,N_19237);
nand U25929 (N_25929,N_18481,N_23642);
xnor U25930 (N_25930,N_20001,N_21625);
nor U25931 (N_25931,N_20810,N_18444);
or U25932 (N_25932,N_23316,N_18125);
xnor U25933 (N_25933,N_20488,N_23570);
nand U25934 (N_25934,N_19129,N_20829);
xor U25935 (N_25935,N_20927,N_18424);
nor U25936 (N_25936,N_21520,N_21090);
nor U25937 (N_25937,N_21037,N_22036);
nand U25938 (N_25938,N_18107,N_20680);
nor U25939 (N_25939,N_23490,N_23969);
or U25940 (N_25940,N_23093,N_18895);
or U25941 (N_25941,N_19167,N_19543);
and U25942 (N_25942,N_20733,N_21317);
or U25943 (N_25943,N_19845,N_19836);
or U25944 (N_25944,N_21472,N_20719);
nor U25945 (N_25945,N_21333,N_23068);
and U25946 (N_25946,N_21787,N_22353);
nand U25947 (N_25947,N_20094,N_21928);
nand U25948 (N_25948,N_18109,N_22564);
and U25949 (N_25949,N_20035,N_19537);
or U25950 (N_25950,N_20045,N_23585);
or U25951 (N_25951,N_22757,N_20089);
or U25952 (N_25952,N_23428,N_19117);
nor U25953 (N_25953,N_23492,N_18168);
nor U25954 (N_25954,N_21620,N_19406);
or U25955 (N_25955,N_21884,N_22659);
nand U25956 (N_25956,N_22481,N_18417);
xor U25957 (N_25957,N_18205,N_21122);
nor U25958 (N_25958,N_20181,N_19650);
and U25959 (N_25959,N_22955,N_19785);
or U25960 (N_25960,N_22539,N_22389);
nor U25961 (N_25961,N_21973,N_20061);
and U25962 (N_25962,N_18878,N_23671);
or U25963 (N_25963,N_19266,N_21764);
and U25964 (N_25964,N_19192,N_20404);
or U25965 (N_25965,N_19138,N_19119);
nor U25966 (N_25966,N_18835,N_21767);
nand U25967 (N_25967,N_21697,N_22087);
or U25968 (N_25968,N_22848,N_18598);
nor U25969 (N_25969,N_22304,N_23581);
and U25970 (N_25970,N_20759,N_21315);
nor U25971 (N_25971,N_22286,N_23476);
nand U25972 (N_25972,N_22926,N_18040);
nand U25973 (N_25973,N_20728,N_21660);
and U25974 (N_25974,N_23663,N_22529);
or U25975 (N_25975,N_18563,N_18113);
nand U25976 (N_25976,N_19381,N_18612);
and U25977 (N_25977,N_20523,N_23808);
xnor U25978 (N_25978,N_23233,N_18600);
or U25979 (N_25979,N_19083,N_19536);
nor U25980 (N_25980,N_23430,N_21876);
and U25981 (N_25981,N_20079,N_22635);
and U25982 (N_25982,N_19186,N_23079);
xnor U25983 (N_25983,N_20817,N_19587);
nand U25984 (N_25984,N_21115,N_19178);
or U25985 (N_25985,N_21963,N_23104);
nor U25986 (N_25986,N_19784,N_19855);
and U25987 (N_25987,N_20929,N_18541);
xnor U25988 (N_25988,N_19397,N_19432);
nand U25989 (N_25989,N_23740,N_21981);
and U25990 (N_25990,N_19325,N_18389);
or U25991 (N_25991,N_22312,N_21029);
and U25992 (N_25992,N_18978,N_21309);
or U25993 (N_25993,N_23610,N_18225);
nand U25994 (N_25994,N_21005,N_19122);
nor U25995 (N_25995,N_18755,N_22921);
and U25996 (N_25996,N_19473,N_22552);
or U25997 (N_25997,N_23668,N_23034);
or U25998 (N_25998,N_18903,N_23964);
or U25999 (N_25999,N_23282,N_20550);
or U26000 (N_26000,N_21533,N_19011);
nor U26001 (N_26001,N_19238,N_21386);
nor U26002 (N_26002,N_22859,N_18135);
xnor U26003 (N_26003,N_19035,N_18451);
and U26004 (N_26004,N_23221,N_18289);
xnor U26005 (N_26005,N_23300,N_21723);
nand U26006 (N_26006,N_20441,N_21116);
or U26007 (N_26007,N_21288,N_23810);
or U26008 (N_26008,N_19728,N_19525);
or U26009 (N_26009,N_22041,N_18922);
and U26010 (N_26010,N_19890,N_21894);
and U26011 (N_26011,N_19614,N_19175);
xnor U26012 (N_26012,N_22358,N_23678);
nor U26013 (N_26013,N_20752,N_23288);
xnor U26014 (N_26014,N_18116,N_19573);
or U26015 (N_26015,N_18977,N_20920);
nand U26016 (N_26016,N_21435,N_22230);
nand U26017 (N_26017,N_19973,N_20706);
nand U26018 (N_26018,N_19868,N_18076);
or U26019 (N_26019,N_21791,N_23646);
or U26020 (N_26020,N_18187,N_20756);
xnor U26021 (N_26021,N_18058,N_21776);
nand U26022 (N_26022,N_21027,N_23705);
nand U26023 (N_26023,N_18099,N_22753);
nand U26024 (N_26024,N_22739,N_23129);
nand U26025 (N_26025,N_22179,N_20661);
and U26026 (N_26026,N_20607,N_21503);
and U26027 (N_26027,N_23066,N_19112);
and U26028 (N_26028,N_22466,N_19579);
or U26029 (N_26029,N_18876,N_19481);
nor U26030 (N_26030,N_22508,N_18567);
nand U26031 (N_26031,N_21235,N_23277);
or U26032 (N_26032,N_22813,N_19919);
and U26033 (N_26033,N_22012,N_23812);
nor U26034 (N_26034,N_19153,N_18067);
nand U26035 (N_26035,N_20592,N_22538);
nor U26036 (N_26036,N_22018,N_20403);
and U26037 (N_26037,N_19580,N_19162);
nand U26038 (N_26038,N_21492,N_21992);
nand U26039 (N_26039,N_21781,N_20443);
or U26040 (N_26040,N_18792,N_19479);
nand U26041 (N_26041,N_23972,N_21394);
nor U26042 (N_26042,N_22550,N_23067);
or U26043 (N_26043,N_19917,N_23884);
nand U26044 (N_26044,N_18540,N_21855);
or U26045 (N_26045,N_20310,N_23872);
and U26046 (N_26046,N_21195,N_23347);
nor U26047 (N_26047,N_23657,N_19458);
or U26048 (N_26048,N_20473,N_22647);
xnor U26049 (N_26049,N_22769,N_23694);
and U26050 (N_26050,N_18419,N_18933);
or U26051 (N_26051,N_20579,N_18528);
nand U26052 (N_26052,N_21340,N_19311);
or U26053 (N_26053,N_18483,N_20170);
or U26054 (N_26054,N_19647,N_19857);
and U26055 (N_26055,N_21547,N_23985);
or U26056 (N_26056,N_20977,N_21762);
and U26057 (N_26057,N_22344,N_19740);
nand U26058 (N_26058,N_22820,N_21663);
xnor U26059 (N_26059,N_23408,N_20771);
nand U26060 (N_26060,N_21539,N_18686);
and U26061 (N_26061,N_18884,N_19403);
nand U26062 (N_26062,N_20775,N_19006);
and U26063 (N_26063,N_19763,N_20030);
nand U26064 (N_26064,N_20799,N_21276);
and U26065 (N_26065,N_18439,N_18098);
nor U26066 (N_26066,N_18816,N_23496);
nand U26067 (N_26067,N_20748,N_23509);
nor U26068 (N_26068,N_21645,N_19871);
or U26069 (N_26069,N_22566,N_19915);
nand U26070 (N_26070,N_18751,N_21923);
or U26071 (N_26071,N_21225,N_19849);
and U26072 (N_26072,N_19725,N_21698);
and U26073 (N_26073,N_18272,N_20141);
and U26074 (N_26074,N_22453,N_20368);
nor U26075 (N_26075,N_19453,N_21743);
nand U26076 (N_26076,N_22091,N_22611);
and U26077 (N_26077,N_22835,N_21452);
nor U26078 (N_26078,N_22081,N_18949);
or U26079 (N_26079,N_19435,N_18175);
nand U26080 (N_26080,N_23952,N_19124);
nor U26081 (N_26081,N_20195,N_19147);
or U26082 (N_26082,N_19426,N_18760);
nand U26083 (N_26083,N_21323,N_20949);
nor U26084 (N_26084,N_22080,N_19985);
and U26085 (N_26085,N_20577,N_21509);
nand U26086 (N_26086,N_23957,N_18808);
nand U26087 (N_26087,N_19222,N_22442);
nor U26088 (N_26088,N_23327,N_20451);
and U26089 (N_26089,N_19661,N_21349);
xnor U26090 (N_26090,N_23653,N_20758);
nand U26091 (N_26091,N_20006,N_21606);
nor U26092 (N_26092,N_20908,N_18810);
and U26093 (N_26093,N_22639,N_23487);
nor U26094 (N_26094,N_18007,N_20453);
nand U26095 (N_26095,N_19139,N_21039);
nand U26096 (N_26096,N_20860,N_19874);
nor U26097 (N_26097,N_20060,N_19252);
nand U26098 (N_26098,N_23231,N_22954);
or U26099 (N_26099,N_18716,N_19259);
nand U26100 (N_26100,N_18092,N_23567);
and U26101 (N_26101,N_21580,N_23933);
nand U26102 (N_26102,N_23420,N_22352);
or U26103 (N_26103,N_20703,N_21893);
xnor U26104 (N_26104,N_19030,N_20741);
or U26105 (N_26105,N_18256,N_22064);
or U26106 (N_26106,N_20755,N_23280);
nand U26107 (N_26107,N_21907,N_23472);
and U26108 (N_26108,N_18597,N_22246);
or U26109 (N_26109,N_19799,N_23916);
nor U26110 (N_26110,N_19324,N_22660);
nor U26111 (N_26111,N_18100,N_19838);
nand U26112 (N_26112,N_23410,N_19290);
or U26113 (N_26113,N_20087,N_22981);
nor U26114 (N_26114,N_21621,N_23511);
and U26115 (N_26115,N_19844,N_20238);
nor U26116 (N_26116,N_22043,N_19368);
nor U26117 (N_26117,N_18065,N_23625);
or U26118 (N_26118,N_20560,N_21788);
nor U26119 (N_26119,N_23942,N_20871);
or U26120 (N_26120,N_21938,N_20918);
and U26121 (N_26121,N_19837,N_23746);
nor U26122 (N_26122,N_19605,N_23590);
xnor U26123 (N_26123,N_22309,N_20348);
nand U26124 (N_26124,N_22569,N_20174);
nand U26125 (N_26125,N_23996,N_18584);
nor U26126 (N_26126,N_22436,N_20464);
nand U26127 (N_26127,N_21569,N_23698);
or U26128 (N_26128,N_21343,N_20781);
nor U26129 (N_26129,N_22201,N_21153);
or U26130 (N_26130,N_19491,N_23805);
nand U26131 (N_26131,N_21977,N_23308);
or U26132 (N_26132,N_18788,N_18084);
or U26133 (N_26133,N_21231,N_20266);
and U26134 (N_26134,N_18953,N_18573);
or U26135 (N_26135,N_21829,N_23118);
and U26136 (N_26136,N_18574,N_20963);
or U26137 (N_26137,N_19709,N_22772);
xnor U26138 (N_26138,N_18844,N_19366);
nor U26139 (N_26139,N_22450,N_22052);
nand U26140 (N_26140,N_18564,N_23800);
or U26141 (N_26141,N_19273,N_18510);
nand U26142 (N_26142,N_22351,N_19651);
nor U26143 (N_26143,N_19150,N_22001);
and U26144 (N_26144,N_18615,N_22330);
or U26145 (N_26145,N_18867,N_18646);
and U26146 (N_26146,N_22473,N_23772);
nand U26147 (N_26147,N_22521,N_21647);
nand U26148 (N_26148,N_23522,N_23007);
nor U26149 (N_26149,N_19815,N_21066);
nand U26150 (N_26150,N_18472,N_22679);
nor U26151 (N_26151,N_21669,N_18242);
nor U26152 (N_26152,N_20099,N_19143);
and U26153 (N_26153,N_18034,N_18277);
or U26154 (N_26154,N_23894,N_21281);
and U26155 (N_26155,N_19361,N_22950);
xor U26156 (N_26156,N_18159,N_22192);
and U26157 (N_26157,N_23493,N_18315);
and U26158 (N_26158,N_18526,N_19000);
xor U26159 (N_26159,N_20218,N_20988);
xnor U26160 (N_26160,N_20354,N_18382);
nor U26161 (N_26161,N_18579,N_21803);
nand U26162 (N_26162,N_18664,N_18847);
nor U26163 (N_26163,N_22007,N_23521);
or U26164 (N_26164,N_20658,N_23449);
or U26165 (N_26165,N_19847,N_20290);
or U26166 (N_26166,N_20780,N_19788);
nand U26167 (N_26167,N_22366,N_21406);
or U26168 (N_26168,N_21410,N_21854);
nand U26169 (N_26169,N_21766,N_23622);
or U26170 (N_26170,N_20237,N_22506);
nand U26171 (N_26171,N_21143,N_21543);
xor U26172 (N_26172,N_18941,N_22802);
nor U26173 (N_26173,N_20595,N_21215);
xnor U26174 (N_26174,N_18190,N_19673);
and U26175 (N_26175,N_22973,N_21046);
and U26176 (N_26176,N_18061,N_19095);
and U26177 (N_26177,N_22045,N_23238);
or U26178 (N_26178,N_22625,N_18261);
and U26179 (N_26179,N_20632,N_20826);
nand U26180 (N_26180,N_20763,N_23274);
nand U26181 (N_26181,N_21469,N_20804);
nor U26182 (N_26182,N_18269,N_22786);
and U26183 (N_26183,N_18758,N_18408);
nor U26184 (N_26184,N_23720,N_22999);
nor U26185 (N_26185,N_21945,N_21785);
nor U26186 (N_26186,N_23839,N_21873);
or U26187 (N_26187,N_20842,N_22423);
nand U26188 (N_26188,N_22837,N_18955);
and U26189 (N_26189,N_19632,N_19705);
and U26190 (N_26190,N_19627,N_19945);
and U26191 (N_26191,N_20827,N_18931);
and U26192 (N_26192,N_20427,N_21994);
and U26193 (N_26193,N_20984,N_21381);
and U26194 (N_26194,N_19631,N_19013);
and U26195 (N_26195,N_20024,N_20076);
nand U26196 (N_26196,N_20711,N_19567);
and U26197 (N_26197,N_18211,N_21013);
or U26198 (N_26198,N_20954,N_19210);
and U26199 (N_26199,N_21018,N_21264);
and U26200 (N_26200,N_23161,N_23995);
xnor U26201 (N_26201,N_18771,N_22103);
xor U26202 (N_26202,N_18547,N_20604);
xor U26203 (N_26203,N_19040,N_18819);
or U26204 (N_26204,N_20985,N_22284);
and U26205 (N_26205,N_22171,N_21326);
and U26206 (N_26206,N_20227,N_21783);
nand U26207 (N_26207,N_20419,N_20957);
or U26208 (N_26208,N_23782,N_20628);
nor U26209 (N_26209,N_22754,N_21602);
or U26210 (N_26210,N_21921,N_23409);
or U26211 (N_26211,N_21612,N_21025);
xor U26212 (N_26212,N_18718,N_21991);
nor U26213 (N_26213,N_18603,N_22818);
nand U26214 (N_26214,N_23021,N_18307);
nand U26215 (N_26215,N_18585,N_18149);
nor U26216 (N_26216,N_21429,N_21719);
nand U26217 (N_26217,N_23801,N_18770);
nand U26218 (N_26218,N_22439,N_19372);
and U26219 (N_26219,N_23910,N_18554);
xor U26220 (N_26220,N_20331,N_20915);
or U26221 (N_26221,N_19400,N_19244);
and U26222 (N_26222,N_22457,N_23921);
and U26223 (N_26223,N_21259,N_20445);
or U26224 (N_26224,N_21380,N_20876);
and U26225 (N_26225,N_23155,N_18973);
nor U26226 (N_26226,N_21373,N_20339);
xor U26227 (N_26227,N_21771,N_21255);
nand U26228 (N_26228,N_19123,N_20169);
and U26229 (N_26229,N_20932,N_22397);
nor U26230 (N_26230,N_23214,N_19701);
xnor U26231 (N_26231,N_23002,N_18711);
xnor U26232 (N_26232,N_21083,N_23456);
xor U26233 (N_26233,N_18346,N_23943);
or U26234 (N_26234,N_21052,N_21897);
or U26235 (N_26235,N_22597,N_20306);
or U26236 (N_26236,N_19544,N_20766);
nand U26237 (N_26237,N_19048,N_20586);
or U26238 (N_26238,N_19608,N_19718);
nor U26239 (N_26239,N_22565,N_20520);
and U26240 (N_26240,N_18446,N_23846);
or U26241 (N_26241,N_22189,N_22771);
nand U26242 (N_26242,N_20381,N_21405);
or U26243 (N_26243,N_22459,N_23559);
nand U26244 (N_26244,N_22384,N_21797);
or U26245 (N_26245,N_21319,N_22976);
nand U26246 (N_26246,N_19979,N_22796);
nand U26247 (N_26247,N_19345,N_18595);
nor U26248 (N_26248,N_18692,N_19022);
nand U26249 (N_26249,N_21699,N_19660);
nor U26250 (N_26250,N_22223,N_22308);
and U26251 (N_26251,N_18431,N_21639);
nor U26252 (N_26252,N_20104,N_18217);
xor U26253 (N_26253,N_20359,N_22748);
nor U26254 (N_26254,N_22904,N_19523);
nor U26255 (N_26255,N_19340,N_19263);
nand U26256 (N_26256,N_19638,N_20396);
or U26257 (N_26257,N_20205,N_20149);
nand U26258 (N_26258,N_19848,N_22512);
or U26259 (N_26259,N_19058,N_19009);
nor U26260 (N_26260,N_23281,N_21008);
and U26261 (N_26261,N_21686,N_19017);
or U26262 (N_26262,N_23645,N_18894);
nand U26263 (N_26263,N_22282,N_19767);
or U26264 (N_26264,N_22907,N_21038);
nand U26265 (N_26265,N_18764,N_20244);
nand U26266 (N_26266,N_19265,N_21903);
xor U26267 (N_26267,N_23464,N_19160);
nor U26268 (N_26268,N_20145,N_20102);
nand U26269 (N_26269,N_22548,N_21451);
nor U26270 (N_26270,N_22940,N_21531);
or U26271 (N_26271,N_22928,N_21711);
or U26272 (N_26272,N_20486,N_21862);
or U26273 (N_26273,N_18807,N_19814);
nor U26274 (N_26274,N_21351,N_18298);
nand U26275 (N_26275,N_23605,N_19050);
nor U26276 (N_26276,N_23081,N_19641);
and U26277 (N_26277,N_22368,N_18397);
and U26278 (N_26278,N_21614,N_23735);
xor U26279 (N_26279,N_23820,N_21779);
nor U26280 (N_26280,N_19445,N_22360);
and U26281 (N_26281,N_20474,N_21584);
nand U26282 (N_26282,N_21666,N_22440);
and U26283 (N_26283,N_21022,N_22549);
nand U26284 (N_26284,N_19738,N_22199);
or U26285 (N_26285,N_20529,N_23151);
nor U26286 (N_26286,N_20082,N_18221);
nor U26287 (N_26287,N_21581,N_23399);
nand U26288 (N_26288,N_18594,N_23821);
nor U26289 (N_26289,N_19450,N_23959);
or U26290 (N_26290,N_19268,N_19158);
nor U26291 (N_26291,N_22562,N_18766);
nor U26292 (N_26292,N_18658,N_19643);
nor U26293 (N_26293,N_21632,N_19956);
and U26294 (N_26294,N_23824,N_20355);
and U26295 (N_26295,N_20270,N_19420);
nor U26296 (N_26296,N_18275,N_23459);
or U26297 (N_26297,N_20764,N_22083);
nand U26298 (N_26298,N_21093,N_21805);
and U26299 (N_26299,N_23874,N_18020);
and U26300 (N_26300,N_18577,N_22101);
nand U26301 (N_26301,N_23727,N_18393);
nand U26302 (N_26302,N_19467,N_19779);
nand U26303 (N_26303,N_21227,N_18485);
or U26304 (N_26304,N_21359,N_20414);
nand U26305 (N_26305,N_23435,N_21484);
xnor U26306 (N_26306,N_22030,N_18892);
nand U26307 (N_26307,N_21197,N_18252);
nor U26308 (N_26308,N_19552,N_23518);
or U26309 (N_26309,N_22778,N_20116);
nor U26310 (N_26310,N_21657,N_18283);
or U26311 (N_26311,N_23452,N_18087);
and U26312 (N_26312,N_19822,N_20938);
and U26313 (N_26313,N_19512,N_18123);
xor U26314 (N_26314,N_20465,N_21421);
or U26315 (N_26315,N_19056,N_18582);
nor U26316 (N_26316,N_19219,N_18729);
and U26317 (N_26317,N_19442,N_18353);
and U26318 (N_26318,N_20390,N_20536);
nand U26319 (N_26319,N_19180,N_20251);
nand U26320 (N_26320,N_19383,N_21590);
and U26321 (N_26321,N_21242,N_21995);
and U26322 (N_26322,N_23144,N_23170);
xnor U26323 (N_26323,N_22707,N_20622);
nand U26324 (N_26324,N_19019,N_21979);
nor U26325 (N_26325,N_22468,N_23264);
and U26326 (N_26326,N_18416,N_18821);
and U26327 (N_26327,N_22107,N_23309);
nor U26328 (N_26328,N_18000,N_23411);
nand U26329 (N_26329,N_19507,N_21859);
xnor U26330 (N_26330,N_19455,N_22958);
nand U26331 (N_26331,N_20934,N_19823);
nor U26332 (N_26332,N_19988,N_23875);
or U26333 (N_26333,N_20828,N_22865);
xor U26334 (N_26334,N_21216,N_20423);
and U26335 (N_26335,N_18088,N_22067);
and U26336 (N_26336,N_18544,N_23326);
nand U26337 (N_26337,N_19436,N_23797);
nor U26338 (N_26338,N_23168,N_20689);
nor U26339 (N_26339,N_19929,N_20247);
and U26340 (N_26340,N_21226,N_22128);
and U26341 (N_26341,N_23292,N_21002);
nand U26342 (N_26342,N_23340,N_23325);
nor U26343 (N_26343,N_22752,N_22157);
and U26344 (N_26344,N_18090,N_20736);
and U26345 (N_26345,N_21993,N_21597);
nand U26346 (N_26346,N_20477,N_19004);
nand U26347 (N_26347,N_21631,N_23236);
nand U26348 (N_26348,N_18016,N_20042);
nand U26349 (N_26349,N_23615,N_19080);
nand U26350 (N_26350,N_22888,N_23441);
or U26351 (N_26351,N_18271,N_19430);
and U26352 (N_26352,N_18975,N_23749);
or U26353 (N_26353,N_20651,N_20329);
nand U26354 (N_26354,N_23924,N_22050);
nor U26355 (N_26355,N_19931,N_21578);
and U26356 (N_26356,N_22561,N_19234);
xnor U26357 (N_26357,N_22963,N_20753);
or U26358 (N_26358,N_23908,N_22485);
nor U26359 (N_26359,N_21129,N_22930);
and U26360 (N_26360,N_22807,N_22173);
and U26361 (N_26361,N_22295,N_21407);
nor U26362 (N_26362,N_21758,N_18787);
nand U26363 (N_26363,N_23377,N_18245);
and U26364 (N_26364,N_22897,N_19737);
and U26365 (N_26365,N_22526,N_19630);
nand U26366 (N_26366,N_21822,N_23858);
nor U26367 (N_26367,N_20746,N_18475);
and U26368 (N_26368,N_22948,N_23507);
and U26369 (N_26369,N_22543,N_20002);
or U26370 (N_26370,N_23059,N_21379);
nand U26371 (N_26371,N_19472,N_23630);
nand U26372 (N_26372,N_22190,N_21835);
or U26373 (N_26373,N_22580,N_23183);
and U26374 (N_26374,N_23029,N_21983);
nor U26375 (N_26375,N_22215,N_20013);
nor U26376 (N_26376,N_18616,N_23896);
nand U26377 (N_26377,N_23498,N_18017);
nand U26378 (N_26378,N_18559,N_20641);
nor U26379 (N_26379,N_20845,N_23111);
and U26380 (N_26380,N_23706,N_23578);
nor U26381 (N_26381,N_21646,N_18626);
and U26382 (N_26382,N_21209,N_23796);
and U26383 (N_26383,N_23154,N_20129);
nor U26384 (N_26384,N_18666,N_23404);
and U26385 (N_26385,N_22700,N_22355);
and U26386 (N_26386,N_18492,N_23126);
nor U26387 (N_26387,N_20106,N_23939);
or U26388 (N_26388,N_18376,N_19734);
or U26389 (N_26389,N_23329,N_22520);
nor U26390 (N_26390,N_18747,N_19695);
xor U26391 (N_26391,N_22127,N_22089);
nand U26392 (N_26392,N_21416,N_23940);
and U26393 (N_26393,N_18103,N_23175);
or U26394 (N_26394,N_23092,N_21086);
and U26395 (N_26395,N_22159,N_21654);
xor U26396 (N_26396,N_21447,N_23601);
or U26397 (N_26397,N_22183,N_20553);
and U26398 (N_26398,N_21599,N_19699);
nand U26399 (N_26399,N_20085,N_23685);
and U26400 (N_26400,N_19294,N_18546);
or U26401 (N_26401,N_23953,N_22951);
or U26402 (N_26402,N_18215,N_23216);
nand U26403 (N_26403,N_19644,N_22871);
nor U26404 (N_26404,N_18323,N_21392);
or U26405 (N_26405,N_20502,N_21763);
and U26406 (N_26406,N_21444,N_21760);
and U26407 (N_26407,N_20421,N_20882);
xor U26408 (N_26408,N_18802,N_19686);
and U26409 (N_26409,N_23650,N_23237);
and U26410 (N_26410,N_22693,N_18310);
nand U26411 (N_26411,N_21658,N_23444);
nor U26412 (N_26412,N_22165,N_18437);
or U26413 (N_26413,N_23302,N_21168);
and U26414 (N_26414,N_20048,N_18378);
xor U26415 (N_26415,N_18063,N_22884);
or U26416 (N_26416,N_20645,N_21450);
nor U26417 (N_26417,N_20125,N_19218);
and U26418 (N_26418,N_22856,N_20784);
or U26419 (N_26419,N_21311,N_22379);
or U26420 (N_26420,N_22726,N_19937);
xnor U26421 (N_26421,N_21420,N_23082);
and U26422 (N_26422,N_21714,N_21283);
nand U26423 (N_26423,N_18182,N_22777);
nand U26424 (N_26424,N_19498,N_23462);
and U26425 (N_26425,N_19829,N_22371);
xnor U26426 (N_26426,N_20101,N_20973);
nor U26427 (N_26427,N_20749,N_22270);
and U26428 (N_26428,N_21878,N_22398);
and U26429 (N_26429,N_20570,N_22511);
or U26430 (N_26430,N_22643,N_22993);
nor U26431 (N_26431,N_22741,N_19141);
and U26432 (N_26432,N_18115,N_20487);
and U26433 (N_26433,N_20426,N_22979);
nand U26434 (N_26434,N_19395,N_19084);
nand U26435 (N_26435,N_20760,N_19932);
or U26436 (N_26436,N_19384,N_22290);
nor U26437 (N_26437,N_20972,N_22645);
or U26438 (N_26438,N_23102,N_23393);
and U26439 (N_26439,N_18240,N_22292);
and U26440 (N_26440,N_18868,N_20815);
nor U26441 (N_26441,N_23296,N_18690);
nor U26442 (N_26442,N_20158,N_20772);
xnor U26443 (N_26443,N_22875,N_19692);
xor U26444 (N_26444,N_19551,N_21443);
or U26445 (N_26445,N_23947,N_23930);
or U26446 (N_26446,N_21040,N_19648);
xnor U26447 (N_26447,N_18717,N_23937);
or U26448 (N_26448,N_19783,N_19853);
and U26449 (N_26449,N_18679,N_23555);
or U26450 (N_26450,N_23451,N_21726);
nand U26451 (N_26451,N_18580,N_20989);
or U26452 (N_26452,N_20164,N_19516);
and U26453 (N_26453,N_18698,N_23535);
nand U26454 (N_26454,N_20112,N_20868);
xor U26455 (N_26455,N_21700,N_21941);
or U26456 (N_26456,N_22394,N_18568);
or U26457 (N_26457,N_22535,N_23714);
nor U26458 (N_26458,N_19355,N_23022);
nor U26459 (N_26459,N_23387,N_23061);
nand U26460 (N_26460,N_23988,N_22651);
nand U26461 (N_26461,N_23065,N_18833);
nor U26462 (N_26462,N_20783,N_22154);
and U26463 (N_26463,N_19231,N_22676);
or U26464 (N_26464,N_23687,N_23713);
and U26465 (N_26465,N_23586,N_23145);
and U26466 (N_26466,N_20392,N_23579);
or U26467 (N_26467,N_19298,N_21370);
or U26468 (N_26468,N_19804,N_20691);
nor U26469 (N_26469,N_21892,N_22102);
or U26470 (N_26470,N_19550,N_19949);
nor U26471 (N_26471,N_22338,N_22621);
nor U26472 (N_26472,N_21149,N_18336);
or U26473 (N_26473,N_21135,N_18202);
and U26474 (N_26474,N_22524,N_22815);
nor U26475 (N_26475,N_23617,N_20005);
or U26476 (N_26476,N_18939,N_23962);
and U26477 (N_26477,N_22497,N_23592);
nor U26478 (N_26478,N_22274,N_23830);
or U26479 (N_26479,N_18029,N_21154);
or U26480 (N_26480,N_18593,N_18398);
or U26481 (N_26481,N_19196,N_23179);
nor U26482 (N_26482,N_21710,N_19540);
and U26483 (N_26483,N_19793,N_23792);
and U26484 (N_26484,N_23006,N_20223);
and U26485 (N_26485,N_19802,N_19257);
xnor U26486 (N_26486,N_21546,N_23348);
and U26487 (N_26487,N_18036,N_22257);
and U26488 (N_26488,N_22006,N_23855);
nor U26489 (N_26489,N_21477,N_22606);
or U26490 (N_26490,N_18781,N_23269);
nor U26491 (N_26491,N_21413,N_18448);
or U26492 (N_26492,N_23305,N_22456);
or U26493 (N_26493,N_23193,N_22893);
or U26494 (N_26494,N_18653,N_19499);
nand U26495 (N_26495,N_20075,N_22340);
nor U26496 (N_26496,N_22211,N_23499);
nor U26497 (N_26497,N_22938,N_22996);
xnor U26498 (N_26498,N_19302,N_22065);
nand U26499 (N_26499,N_18517,N_23928);
and U26500 (N_26500,N_21458,N_20841);
nor U26501 (N_26501,N_21254,N_23360);
and U26502 (N_26502,N_19315,N_21177);
nor U26503 (N_26503,N_23185,N_23956);
nor U26504 (N_26504,N_22809,N_18561);
or U26505 (N_26505,N_21383,N_18262);
nand U26506 (N_26506,N_20496,N_19564);
or U26507 (N_26507,N_19969,N_22321);
xor U26508 (N_26508,N_23245,N_23934);
or U26509 (N_26509,N_20769,N_22622);
and U26510 (N_26510,N_21482,N_19621);
and U26511 (N_26511,N_23001,N_18096);
xnor U26512 (N_26512,N_18539,N_20108);
and U26513 (N_26513,N_20557,N_23047);
nand U26514 (N_26514,N_20757,N_20901);
and U26515 (N_26515,N_19504,N_18569);
nor U26516 (N_26516,N_19682,N_18119);
nor U26517 (N_26517,N_20370,N_22805);
nand U26518 (N_26518,N_23542,N_19731);
nand U26519 (N_26519,N_22269,N_18144);
or U26520 (N_26520,N_19082,N_18072);
nand U26521 (N_26521,N_22010,N_21355);
nand U26522 (N_26522,N_18158,N_20470);
or U26523 (N_26523,N_19876,N_23524);
or U26524 (N_26524,N_22601,N_20044);
nand U26525 (N_26525,N_20979,N_19227);
nand U26526 (N_26526,N_22125,N_22575);
or U26527 (N_26527,N_22441,N_21140);
xnor U26528 (N_26528,N_20235,N_18360);
or U26529 (N_26529,N_18106,N_18938);
and U26530 (N_26530,N_22268,N_22634);
or U26531 (N_26531,N_22364,N_21670);
nand U26532 (N_26532,N_22068,N_20877);
and U26533 (N_26533,N_22465,N_18332);
or U26534 (N_26534,N_22303,N_23040);
and U26535 (N_26535,N_22435,N_22073);
nand U26536 (N_26536,N_19866,N_19480);
nor U26537 (N_26537,N_23854,N_18045);
nand U26538 (N_26538,N_22139,N_18164);
nand U26539 (N_26539,N_23950,N_21036);
and U26540 (N_26540,N_18556,N_22461);
and U26541 (N_26541,N_19689,N_23880);
and U26542 (N_26542,N_18634,N_22424);
and U26543 (N_26543,N_19223,N_19762);
and U26544 (N_26544,N_20307,N_22785);
or U26545 (N_26545,N_22956,N_18587);
and U26546 (N_26546,N_19399,N_23970);
and U26547 (N_26547,N_22689,N_21857);
and U26548 (N_26548,N_19044,N_22116);
or U26549 (N_26549,N_22861,N_18111);
nor U26550 (N_26550,N_20707,N_20285);
or U26551 (N_26551,N_20319,N_23075);
and U26552 (N_26552,N_20907,N_20147);
xnor U26553 (N_26553,N_18959,N_21442);
or U26554 (N_26554,N_21702,N_19657);
xnor U26555 (N_26555,N_20886,N_18062);
or U26556 (N_26556,N_19754,N_21679);
nand U26557 (N_26557,N_18179,N_21927);
nor U26558 (N_26558,N_22235,N_19069);
nand U26559 (N_26559,N_22100,N_18478);
and U26560 (N_26560,N_22584,N_19191);
nor U26561 (N_26561,N_18334,N_19880);
or U26562 (N_26562,N_18456,N_18308);
and U26563 (N_26563,N_20955,N_23833);
and U26564 (N_26564,N_21570,N_21178);
nor U26565 (N_26565,N_20506,N_23725);
nor U26566 (N_26566,N_21678,N_22276);
nor U26567 (N_26567,N_21474,N_21049);
nand U26568 (N_26568,N_19454,N_20865);
nor U26569 (N_26569,N_20458,N_23401);
or U26570 (N_26570,N_21491,N_18772);
and U26571 (N_26571,N_22479,N_19269);
and U26572 (N_26572,N_19038,N_19484);
xnor U26573 (N_26573,N_21041,N_19414);
or U26574 (N_26574,N_19161,N_20475);
and U26575 (N_26575,N_22578,N_23005);
nor U26576 (N_26576,N_21028,N_18172);
xor U26577 (N_26577,N_19745,N_18313);
and U26578 (N_26578,N_23739,N_21694);
and U26579 (N_26579,N_21287,N_20609);
nor U26580 (N_26580,N_23429,N_21905);
and U26581 (N_26581,N_20166,N_22296);
and U26582 (N_26582,N_23862,N_19662);
nor U26583 (N_26583,N_18213,N_19300);
and U26584 (N_26584,N_20997,N_21305);
nand U26585 (N_26585,N_23369,N_20224);
xnor U26586 (N_26586,N_21986,N_22531);
nor U26587 (N_26587,N_20440,N_18259);
and U26588 (N_26588,N_18691,N_22846);
nor U26589 (N_26589,N_18014,N_18685);
and U26590 (N_26590,N_22507,N_18491);
and U26591 (N_26591,N_18025,N_21121);
nand U26592 (N_26592,N_19425,N_23468);
nor U26593 (N_26593,N_21500,N_22590);
and U26594 (N_26594,N_23434,N_22488);
or U26595 (N_26595,N_22686,N_20874);
and U26596 (N_26596,N_20679,N_23127);
nor U26597 (N_26597,N_23786,N_22088);
nor U26598 (N_26598,N_19312,N_21496);
nand U26599 (N_26599,N_22889,N_21815);
nor U26600 (N_26600,N_23250,N_18219);
nand U26601 (N_26601,N_18314,N_19895);
or U26602 (N_26602,N_19941,N_22986);
xor U26603 (N_26603,N_18532,N_23425);
nor U26604 (N_26604,N_23774,N_20905);
nand U26605 (N_26605,N_18643,N_18441);
nor U26606 (N_26606,N_23523,N_22984);
nand U26607 (N_26607,N_20909,N_19902);
nor U26608 (N_26608,N_18543,N_18051);
nor U26609 (N_26609,N_18468,N_19513);
and U26610 (N_26610,N_22381,N_19382);
nor U26611 (N_26611,N_23722,N_23162);
nor U26612 (N_26612,N_19790,N_23891);
nor U26613 (N_26613,N_23016,N_19295);
or U26614 (N_26614,N_19831,N_19329);
nand U26615 (N_26615,N_18195,N_23419);
or U26616 (N_26616,N_21784,N_19424);
nor U26617 (N_26617,N_20993,N_23686);
and U26618 (N_26618,N_23936,N_19369);
nor U26619 (N_26619,N_19061,N_18551);
nand U26620 (N_26620,N_19816,N_18535);
or U26621 (N_26621,N_23200,N_20334);
and U26622 (N_26622,N_20961,N_18311);
or U26623 (N_26623,N_18777,N_18480);
xor U26624 (N_26624,N_22767,N_23789);
xor U26625 (N_26625,N_21124,N_20143);
or U26626 (N_26626,N_22273,N_20987);
or U26627 (N_26627,N_20026,N_20111);
or U26628 (N_26628,N_21356,N_18909);
xnor U26629 (N_26629,N_22138,N_23213);
nor U26630 (N_26630,N_20187,N_20059);
nand U26631 (N_26631,N_23977,N_20750);
nand U26632 (N_26632,N_18988,N_21545);
nand U26633 (N_26633,N_18610,N_18902);
nand U26634 (N_26634,N_18385,N_23438);
or U26635 (N_26635,N_21956,N_19297);
nor U26636 (N_26636,N_18300,N_21653);
and U26637 (N_26637,N_21202,N_18027);
and U26638 (N_26638,N_20259,N_20511);
or U26639 (N_26639,N_20664,N_20591);
nor U26640 (N_26640,N_23992,N_21389);
or U26641 (N_26641,N_19065,N_22990);
xor U26642 (N_26642,N_21422,N_22876);
and U26643 (N_26643,N_23114,N_23032);
or U26644 (N_26644,N_19362,N_23124);
nor U26645 (N_26645,N_19602,N_20457);
xnor U26646 (N_26646,N_21385,N_19046);
nand U26647 (N_26647,N_21187,N_18668);
nor U26648 (N_26648,N_20812,N_19338);
nor U26649 (N_26649,N_20709,N_18511);
or U26650 (N_26650,N_23697,N_22801);
and U26651 (N_26651,N_23876,N_19010);
nand U26652 (N_26652,N_23132,N_22612);
nor U26653 (N_26653,N_21585,N_21138);
nor U26654 (N_26654,N_22299,N_21390);
nand U26655 (N_26655,N_21372,N_18848);
nand U26656 (N_26656,N_23115,N_20666);
xor U26657 (N_26657,N_22181,N_21332);
nor U26658 (N_26658,N_20941,N_22451);
nor U26659 (N_26659,N_23342,N_22266);
nand U26660 (N_26660,N_18811,N_22443);
nor U26661 (N_26661,N_18317,N_20969);
or U26662 (N_26662,N_19313,N_23870);
or U26663 (N_26663,N_20761,N_21661);
and U26664 (N_26664,N_23966,N_20053);
or U26665 (N_26665,N_22649,N_18082);
or U26666 (N_26666,N_21080,N_20418);
nor U26667 (N_26667,N_21951,N_22896);
nor U26668 (N_26668,N_23534,N_18695);
nor U26669 (N_26669,N_22267,N_22919);
or U26670 (N_26670,N_21515,N_22434);
or U26671 (N_26671,N_20241,N_18697);
or U26672 (N_26672,N_23388,N_21384);
nand U26673 (N_26673,N_21031,N_21853);
nor U26674 (N_26674,N_19283,N_20401);
or U26675 (N_26675,N_18161,N_18575);
and U26676 (N_26676,N_21357,N_22688);
or U26677 (N_26677,N_21077,N_19350);
and U26678 (N_26678,N_20534,N_21863);
nor U26679 (N_26679,N_19795,N_23666);
and U26680 (N_26680,N_21098,N_18507);
nand U26681 (N_26681,N_20052,N_18997);
xnor U26682 (N_26682,N_19116,N_20745);
xnor U26683 (N_26683,N_21279,N_22247);
and U26684 (N_26684,N_20778,N_20413);
nor U26685 (N_26685,N_23195,N_23742);
nand U26686 (N_26686,N_18667,N_21282);
or U26687 (N_26687,N_18899,N_21285);
or U26688 (N_26688,N_18021,N_22249);
nand U26689 (N_26689,N_18239,N_22200);
or U26690 (N_26690,N_18882,N_22668);
xnor U26691 (N_26691,N_21684,N_23138);
and U26692 (N_26692,N_19940,N_19546);
or U26693 (N_26693,N_19321,N_18629);
nand U26694 (N_26694,N_22336,N_20288);
nor U26695 (N_26695,N_20431,N_20007);
xnor U26696 (N_26696,N_19385,N_21681);
nor U26697 (N_26697,N_22680,N_19645);
and U26698 (N_26698,N_23372,N_23614);
nand U26699 (N_26699,N_19332,N_21241);
and U26700 (N_26700,N_21270,N_18094);
xor U26701 (N_26701,N_19891,N_22252);
or U26702 (N_26702,N_23217,N_18552);
and U26703 (N_26703,N_22901,N_23086);
or U26704 (N_26704,N_23469,N_22275);
or U26705 (N_26705,N_20175,N_22505);
nand U26706 (N_26706,N_22911,N_22577);
or U26707 (N_26707,N_22193,N_23699);
nand U26708 (N_26708,N_21280,N_23502);
nor U26709 (N_26709,N_23770,N_18006);
or U26710 (N_26710,N_22024,N_21899);
nand U26711 (N_26711,N_19708,N_21033);
and U26712 (N_26712,N_22619,N_22784);
nand U26713 (N_26713,N_20924,N_22695);
and U26714 (N_26714,N_20063,N_23383);
nand U26715 (N_26715,N_18400,N_21840);
or U26716 (N_26716,N_21222,N_22306);
nand U26717 (N_26717,N_19066,N_18826);
nor U26718 (N_26718,N_18055,N_23513);
xnor U26719 (N_26719,N_18845,N_23385);
xor U26720 (N_26720,N_19419,N_21130);
xnor U26721 (N_26721,N_20462,N_19765);
nand U26722 (N_26722,N_19018,N_21972);
nand U26723 (N_26723,N_18823,N_21636);
or U26724 (N_26724,N_23667,N_20095);
and U26725 (N_26725,N_18293,N_23431);
nor U26726 (N_26726,N_22332,N_20597);
nor U26727 (N_26727,N_23975,N_19688);
xor U26728 (N_26728,N_18558,N_19261);
or U26729 (N_26729,N_23356,N_21414);
and U26730 (N_26730,N_22311,N_20738);
xor U26731 (N_26731,N_20429,N_23109);
or U26732 (N_26732,N_20642,N_22464);
and U26733 (N_26733,N_23338,N_22178);
nand U26734 (N_26734,N_19144,N_21953);
nor U26735 (N_26735,N_23528,N_18657);
or U26736 (N_26736,N_23621,N_20011);
xor U26737 (N_26737,N_19861,N_19633);
xor U26738 (N_26738,N_19954,N_23552);
and U26739 (N_26739,N_23693,N_20548);
nand U26740 (N_26740,N_20040,N_18655);
or U26741 (N_26741,N_22143,N_18994);
nand U26742 (N_26742,N_20284,N_22860);
nor U26743 (N_26743,N_23715,N_22797);
nand U26744 (N_26744,N_23202,N_18750);
xnor U26745 (N_26745,N_23471,N_22721);
nor U26746 (N_26746,N_21200,N_21119);
nand U26747 (N_26747,N_23205,N_19212);
or U26748 (N_26748,N_20974,N_22209);
nand U26749 (N_26749,N_19817,N_22711);
and U26750 (N_26750,N_23849,N_23898);
or U26751 (N_26751,N_21297,N_18566);
nand U26752 (N_26752,N_23364,N_20525);
xor U26753 (N_26753,N_20207,N_18731);
nand U26754 (N_26754,N_23670,N_18754);
xor U26755 (N_26755,N_22134,N_20676);
nand U26756 (N_26756,N_18188,N_19152);
or U26757 (N_26757,N_22536,N_22716);
and U26758 (N_26758,N_19401,N_23248);
or U26759 (N_26759,N_20103,N_20257);
nor U26760 (N_26760,N_21238,N_19310);
and U26761 (N_26761,N_22417,N_19842);
nor U26762 (N_26762,N_19772,N_22878);
xor U26763 (N_26763,N_18818,N_20350);
or U26764 (N_26764,N_23598,N_23569);
nand U26765 (N_26765,N_20434,N_22447);
xor U26766 (N_26766,N_18258,N_21217);
or U26767 (N_26767,N_22320,N_23009);
and U26768 (N_26768,N_22602,N_21004);
nand U26769 (N_26769,N_20699,N_19519);
or U26770 (N_26770,N_18425,N_18173);
or U26771 (N_26771,N_21045,N_22204);
nand U26772 (N_26772,N_20556,N_19591);
nor U26773 (N_26773,N_19448,N_18586);
nand U26774 (N_26774,N_18101,N_22756);
nand U26775 (N_26775,N_22129,N_23763);
xnor U26776 (N_26776,N_19905,N_20287);
nor U26777 (N_26777,N_19423,N_23759);
nand U26778 (N_26778,N_21170,N_20163);
nand U26779 (N_26779,N_22053,N_21104);
and U26780 (N_26780,N_21084,N_21203);
nand U26781 (N_26781,N_22604,N_20519);
or U26782 (N_26782,N_21329,N_22302);
and U26783 (N_26783,N_22118,N_20853);
or U26784 (N_26784,N_18180,N_23669);
and U26785 (N_26785,N_22738,N_18872);
or U26786 (N_26786,N_19674,N_23414);
or U26787 (N_26787,N_18201,N_19658);
nand U26788 (N_26788,N_19999,N_21610);
nor U26789 (N_26789,N_20890,N_23113);
nor U26790 (N_26790,N_23331,N_19441);
nor U26791 (N_26791,N_18748,N_23806);
or U26792 (N_26792,N_20713,N_20819);
nor U26793 (N_26793,N_18015,N_21957);
nand U26794 (N_26794,N_23483,N_19826);
nand U26795 (N_26795,N_20975,N_18946);
and U26796 (N_26796,N_22613,N_21635);
and U26797 (N_26797,N_19220,N_21378);
xnor U26798 (N_26798,N_18265,N_18678);
nor U26799 (N_26799,N_22658,N_21936);
or U26800 (N_26800,N_18809,N_23239);
nor U26801 (N_26801,N_22074,N_19446);
nand U26802 (N_26802,N_21519,N_18623);
and U26803 (N_26803,N_20855,N_18592);
and U26804 (N_26804,N_20138,N_18963);
and U26805 (N_26805,N_23315,N_19597);
and U26806 (N_26806,N_18893,N_20803);
nand U26807 (N_26807,N_19854,N_22770);
xnor U26808 (N_26808,N_22347,N_21595);
nor U26809 (N_26809,N_18422,N_20047);
or U26810 (N_26810,N_20267,N_21391);
xnor U26811 (N_26811,N_23440,N_21347);
and U26812 (N_26812,N_18429,N_18406);
nor U26813 (N_26813,N_22239,N_23544);
or U26814 (N_26814,N_18970,N_21996);
or U26815 (N_26815,N_23359,N_22737);
nand U26816 (N_26816,N_21072,N_18732);
and U26817 (N_26817,N_18155,N_19984);
or U26818 (N_26818,N_19778,N_19155);
and U26819 (N_26819,N_20951,N_18420);
xor U26820 (N_26820,N_21682,N_20318);
xnor U26821 (N_26821,N_19354,N_19254);
nand U26822 (N_26822,N_19164,N_19555);
nand U26823 (N_26823,N_20914,N_20281);
nand U26824 (N_26824,N_21252,N_21364);
nor U26825 (N_26825,N_19904,N_23596);
nand U26826 (N_26826,N_21263,N_23769);
or U26827 (N_26827,N_22964,N_22685);
and U26828 (N_26828,N_21603,N_21024);
and U26829 (N_26829,N_23776,N_22300);
and U26830 (N_26830,N_23035,N_19514);
or U26831 (N_26831,N_23052,N_22152);
or U26832 (N_26832,N_23147,N_22262);
xnor U26833 (N_26833,N_22287,N_19531);
nor U26834 (N_26834,N_23844,N_20657);
nor U26835 (N_26835,N_19964,N_23888);
nor U26836 (N_26836,N_21455,N_23063);
nand U26837 (N_26837,N_18625,N_19700);
nand U26838 (N_26838,N_22806,N_20747);
and U26839 (N_26839,N_20639,N_23332);
and U26840 (N_26840,N_18043,N_20585);
nand U26841 (N_26841,N_21495,N_19089);
nand U26842 (N_26842,N_23765,N_21501);
xor U26843 (N_26843,N_19464,N_19997);
or U26844 (N_26844,N_23799,N_23160);
nand U26845 (N_26845,N_21023,N_19556);
and U26846 (N_26846,N_22161,N_23433);
nand U26847 (N_26847,N_22614,N_20269);
or U26848 (N_26848,N_22334,N_20541);
and U26849 (N_26849,N_19021,N_21962);
nand U26850 (N_26850,N_18363,N_20346);
or U26851 (N_26851,N_18707,N_20640);
or U26852 (N_26852,N_18095,N_22471);
nand U26853 (N_26853,N_21047,N_23424);
nor U26854 (N_26854,N_18479,N_23857);
and U26855 (N_26855,N_20627,N_18433);
and U26856 (N_26856,N_20123,N_21448);
and U26857 (N_26857,N_22607,N_23626);
nor U26858 (N_26858,N_23442,N_20636);
nand U26859 (N_26859,N_21811,N_18962);
and U26860 (N_26860,N_20115,N_22789);
and U26861 (N_26861,N_23914,N_22416);
nand U26862 (N_26862,N_19054,N_21796);
xor U26863 (N_26863,N_19331,N_23045);
nand U26864 (N_26864,N_19501,N_20652);
nor U26865 (N_26865,N_22824,N_22599);
nor U26866 (N_26866,N_19024,N_18459);
and U26867 (N_26867,N_22404,N_22421);
nor U26868 (N_26868,N_19276,N_18531);
nand U26869 (N_26869,N_21100,N_22283);
nand U26870 (N_26870,N_22515,N_22715);
nor U26871 (N_26871,N_23576,N_23103);
and U26872 (N_26872,N_18700,N_18906);
or U26873 (N_26873,N_20800,N_20793);
nor U26874 (N_26874,N_22745,N_23163);
and U26875 (N_26875,N_21081,N_21341);
nor U26876 (N_26876,N_21014,N_18046);
nand U26877 (N_26877,N_19483,N_23760);
xor U26878 (N_26878,N_18486,N_22260);
nand U26879 (N_26879,N_18954,N_18089);
nand U26880 (N_26880,N_19005,N_22289);
nand U26881 (N_26881,N_20782,N_20700);
and U26882 (N_26882,N_19114,N_21344);
nor U26883 (N_26883,N_18237,N_22141);
or U26884 (N_26884,N_20459,N_18295);
and U26885 (N_26885,N_22513,N_20362);
or U26886 (N_26886,N_22620,N_23363);
nor U26887 (N_26887,N_21064,N_18590);
xnor U26888 (N_26888,N_18080,N_18455);
or U26889 (N_26889,N_22554,N_21573);
and U26890 (N_26890,N_18519,N_18104);
nor U26891 (N_26891,N_20029,N_20461);
nand U26892 (N_26892,N_20409,N_22214);
nor U26893 (N_26893,N_23112,N_19250);
and U26894 (N_26894,N_20922,N_18287);
or U26895 (N_26895,N_18976,N_20020);
and U26896 (N_26896,N_22498,N_23304);
and U26897 (N_26897,N_22155,N_22708);
nor U26898 (N_26898,N_22386,N_20097);
and U26899 (N_26899,N_20212,N_22881);
nor U26900 (N_26900,N_18534,N_23556);
nand U26901 (N_26901,N_19032,N_23373);
or U26902 (N_26902,N_21015,N_18495);
and U26903 (N_26903,N_21541,N_21611);
and U26904 (N_26904,N_22263,N_22108);
nand U26905 (N_26905,N_21523,N_19452);
nand U26906 (N_26906,N_19041,N_19921);
nor U26907 (N_26907,N_22504,N_18993);
nand U26908 (N_26908,N_22631,N_19204);
nand U26909 (N_26909,N_19992,N_19015);
or U26910 (N_26910,N_18133,N_21832);
nor U26911 (N_26911,N_18550,N_18852);
or U26912 (N_26912,N_21205,N_23246);
nor U26913 (N_26913,N_23488,N_20683);
nor U26914 (N_26914,N_18791,N_18285);
nand U26915 (N_26915,N_21030,N_18863);
and U26916 (N_26916,N_21589,N_20498);
nand U26917 (N_26917,N_22858,N_18649);
and U26918 (N_26918,N_22408,N_22714);
and U26919 (N_26919,N_21902,N_23834);
nand U26920 (N_26920,N_22158,N_22849);
nor U26921 (N_26921,N_20630,N_20693);
or U26922 (N_26922,N_20219,N_19938);
or U26923 (N_26923,N_20762,N_21318);
nand U26924 (N_26924,N_21403,N_23091);
or U26925 (N_26925,N_22378,N_20377);
xor U26926 (N_26926,N_19606,N_22137);
nand U26927 (N_26927,N_19037,N_18073);
and U26928 (N_26928,N_19248,N_23203);
and U26929 (N_26929,N_21751,N_23391);
nand U26930 (N_26930,N_20027,N_22681);
and U26931 (N_26931,N_22115,N_23095);
nand U26932 (N_26932,N_23258,N_22915);
nand U26933 (N_26933,N_18351,N_21915);
xor U26934 (N_26934,N_18515,N_21912);
and U26935 (N_26935,N_20863,N_22509);
and U26936 (N_26936,N_19526,N_20535);
or U26937 (N_26937,N_18005,N_18984);
nor U26938 (N_26938,N_19775,N_21577);
nand U26939 (N_26939,N_22072,N_20968);
nand U26940 (N_26940,N_20105,N_22142);
nor U26941 (N_26941,N_19059,N_23976);
nand U26942 (N_26942,N_23251,N_23832);
or U26943 (N_26943,N_23712,N_18908);
nand U26944 (N_26944,N_23370,N_23199);
nor U26945 (N_26945,N_23215,N_21967);
and U26946 (N_26946,N_20000,N_18349);
xnor U26947 (N_26947,N_20965,N_20838);
nand U26948 (N_26948,N_19173,N_20563);
nor U26949 (N_26949,N_20618,N_23917);
nor U26950 (N_26950,N_22983,N_19188);
or U26951 (N_26951,N_23189,N_19494);
and U26952 (N_26952,N_18662,N_18605);
or U26953 (N_26953,N_21512,N_23497);
xor U26954 (N_26954,N_20272,N_20327);
nor U26955 (N_26955,N_20069,N_22170);
nor U26956 (N_26956,N_23971,N_21906);
or U26957 (N_26957,N_18533,N_18632);
and U26958 (N_26958,N_19528,N_21671);
nand U26959 (N_26959,N_21324,N_21554);
and U26960 (N_26960,N_19229,N_21749);
or U26961 (N_26961,N_18487,N_20504);
xor U26962 (N_26962,N_23999,N_22694);
nor U26963 (N_26963,N_20790,N_19337);
nand U26964 (N_26964,N_21704,N_23761);
and U26965 (N_26965,N_19922,N_20998);
nand U26966 (N_26966,N_21003,N_22542);
xor U26967 (N_26967,N_21537,N_22833);
nand U26968 (N_26968,N_22970,N_21733);
and U26969 (N_26969,N_18193,N_23069);
nand U26970 (N_26970,N_18504,N_22186);
or U26971 (N_26971,N_21105,N_23790);
or U26972 (N_26972,N_18888,N_23244);
nor U26973 (N_26973,N_19558,N_19588);
nand U26974 (N_26974,N_21286,N_18279);
xor U26975 (N_26975,N_18952,N_22677);
nand U26976 (N_26976,N_21176,N_23864);
or U26977 (N_26977,N_22038,N_23254);
and U26978 (N_26978,N_21808,N_19409);
nor U26979 (N_26979,N_22701,N_22412);
and U26980 (N_26980,N_22774,N_18141);
xnor U26981 (N_26981,N_21061,N_18924);
xnor U26982 (N_26982,N_20454,N_22920);
nand U26983 (N_26983,N_18860,N_23573);
and U26984 (N_26984,N_18117,N_21613);
or U26985 (N_26985,N_23863,N_21454);
and U26986 (N_26986,N_22343,N_21494);
nor U26987 (N_26987,N_22822,N_21146);
or U26988 (N_26988,N_18302,N_21624);
nor U26989 (N_26989,N_20323,N_18165);
and U26990 (N_26990,N_22766,N_21348);
and U26991 (N_26991,N_20516,N_21224);
and U26992 (N_26992,N_21729,N_19987);
or U26993 (N_26993,N_20888,N_23538);
or U26994 (N_26994,N_19726,N_23817);
and U26995 (N_26995,N_21642,N_19077);
or U26996 (N_26996,N_18854,N_20361);
xor U26997 (N_26997,N_21284,N_23729);
nand U26998 (N_26998,N_22278,N_19364);
and U26999 (N_26999,N_21806,N_20522);
nand U27000 (N_27000,N_18227,N_18419);
nand U27001 (N_27001,N_23470,N_21736);
nand U27002 (N_27002,N_22886,N_23026);
nor U27003 (N_27003,N_21668,N_23356);
or U27004 (N_27004,N_23144,N_19638);
or U27005 (N_27005,N_23611,N_21942);
nand U27006 (N_27006,N_19445,N_22920);
nand U27007 (N_27007,N_22753,N_19738);
or U27008 (N_27008,N_21783,N_22684);
or U27009 (N_27009,N_20291,N_19742);
nand U27010 (N_27010,N_22771,N_23599);
nand U27011 (N_27011,N_19491,N_21090);
and U27012 (N_27012,N_23781,N_21292);
nand U27013 (N_27013,N_22690,N_23682);
nor U27014 (N_27014,N_19346,N_18505);
nand U27015 (N_27015,N_18188,N_20771);
nand U27016 (N_27016,N_23912,N_22155);
nand U27017 (N_27017,N_18309,N_20053);
nor U27018 (N_27018,N_20920,N_22996);
nand U27019 (N_27019,N_23695,N_21174);
nand U27020 (N_27020,N_22866,N_23048);
and U27021 (N_27021,N_21173,N_19032);
or U27022 (N_27022,N_18286,N_19055);
and U27023 (N_27023,N_22739,N_23882);
nor U27024 (N_27024,N_18544,N_23369);
and U27025 (N_27025,N_19530,N_21999);
and U27026 (N_27026,N_20927,N_22127);
and U27027 (N_27027,N_18809,N_23112);
nor U27028 (N_27028,N_19750,N_23222);
or U27029 (N_27029,N_20737,N_20641);
and U27030 (N_27030,N_19176,N_23468);
or U27031 (N_27031,N_22075,N_21367);
and U27032 (N_27032,N_22493,N_21967);
and U27033 (N_27033,N_21881,N_20131);
and U27034 (N_27034,N_20434,N_20616);
nand U27035 (N_27035,N_21058,N_20431);
or U27036 (N_27036,N_22226,N_21373);
nand U27037 (N_27037,N_18098,N_20318);
or U27038 (N_27038,N_19368,N_18330);
nand U27039 (N_27039,N_23759,N_20415);
nand U27040 (N_27040,N_19430,N_19459);
nor U27041 (N_27041,N_21667,N_20598);
and U27042 (N_27042,N_22875,N_19456);
xnor U27043 (N_27043,N_21349,N_18276);
and U27044 (N_27044,N_19068,N_21141);
nor U27045 (N_27045,N_23506,N_23856);
or U27046 (N_27046,N_21547,N_21315);
nor U27047 (N_27047,N_20989,N_18862);
nor U27048 (N_27048,N_22244,N_18647);
or U27049 (N_27049,N_19327,N_20166);
nand U27050 (N_27050,N_19653,N_22620);
and U27051 (N_27051,N_23273,N_23299);
xor U27052 (N_27052,N_22771,N_21487);
nor U27053 (N_27053,N_21615,N_19073);
nand U27054 (N_27054,N_22184,N_22516);
or U27055 (N_27055,N_18731,N_20603);
or U27056 (N_27056,N_21638,N_21884);
and U27057 (N_27057,N_19685,N_21367);
nand U27058 (N_27058,N_20618,N_18657);
nand U27059 (N_27059,N_23027,N_20888);
nor U27060 (N_27060,N_22224,N_22689);
nor U27061 (N_27061,N_18147,N_18928);
nor U27062 (N_27062,N_19575,N_19785);
or U27063 (N_27063,N_23948,N_23382);
or U27064 (N_27064,N_20751,N_18172);
xnor U27065 (N_27065,N_23301,N_19929);
nor U27066 (N_27066,N_23620,N_23822);
nor U27067 (N_27067,N_23544,N_22394);
nor U27068 (N_27068,N_23046,N_23017);
nand U27069 (N_27069,N_20463,N_19847);
or U27070 (N_27070,N_21237,N_19015);
and U27071 (N_27071,N_20016,N_21626);
xor U27072 (N_27072,N_23791,N_21196);
xor U27073 (N_27073,N_22192,N_22556);
nor U27074 (N_27074,N_18685,N_21579);
xnor U27075 (N_27075,N_21270,N_19629);
or U27076 (N_27076,N_22213,N_23614);
nor U27077 (N_27077,N_21262,N_20589);
and U27078 (N_27078,N_19494,N_19845);
and U27079 (N_27079,N_19583,N_20323);
or U27080 (N_27080,N_18120,N_22335);
nand U27081 (N_27081,N_21817,N_23232);
and U27082 (N_27082,N_20167,N_21193);
nor U27083 (N_27083,N_23282,N_20057);
xor U27084 (N_27084,N_20236,N_20534);
nor U27085 (N_27085,N_23383,N_23118);
nor U27086 (N_27086,N_21744,N_20016);
nand U27087 (N_27087,N_19326,N_18020);
xor U27088 (N_27088,N_23157,N_19168);
nand U27089 (N_27089,N_19156,N_18137);
or U27090 (N_27090,N_19295,N_22757);
and U27091 (N_27091,N_18799,N_20795);
and U27092 (N_27092,N_22642,N_18101);
nand U27093 (N_27093,N_18091,N_18633);
nand U27094 (N_27094,N_19251,N_20797);
or U27095 (N_27095,N_19413,N_23846);
nor U27096 (N_27096,N_20701,N_21496);
nor U27097 (N_27097,N_20065,N_21843);
or U27098 (N_27098,N_21397,N_18440);
or U27099 (N_27099,N_22274,N_22873);
nor U27100 (N_27100,N_21004,N_18033);
nand U27101 (N_27101,N_19570,N_21020);
or U27102 (N_27102,N_19492,N_18318);
nor U27103 (N_27103,N_19179,N_21910);
and U27104 (N_27104,N_18452,N_19963);
nand U27105 (N_27105,N_18554,N_20214);
nor U27106 (N_27106,N_22540,N_19748);
xnor U27107 (N_27107,N_21812,N_20959);
nand U27108 (N_27108,N_19192,N_22838);
and U27109 (N_27109,N_23357,N_23772);
nand U27110 (N_27110,N_22429,N_22957);
nand U27111 (N_27111,N_22345,N_22906);
and U27112 (N_27112,N_19972,N_19626);
nor U27113 (N_27113,N_20439,N_23460);
xor U27114 (N_27114,N_22651,N_18110);
and U27115 (N_27115,N_20379,N_19708);
nand U27116 (N_27116,N_23829,N_19443);
xor U27117 (N_27117,N_23606,N_22996);
and U27118 (N_27118,N_20797,N_18361);
nor U27119 (N_27119,N_18445,N_22422);
nand U27120 (N_27120,N_18606,N_23090);
or U27121 (N_27121,N_21692,N_21605);
nor U27122 (N_27122,N_21037,N_23348);
and U27123 (N_27123,N_19809,N_23733);
nor U27124 (N_27124,N_22901,N_20673);
nor U27125 (N_27125,N_23090,N_21637);
or U27126 (N_27126,N_21937,N_19315);
and U27127 (N_27127,N_22574,N_18644);
nor U27128 (N_27128,N_22977,N_19376);
or U27129 (N_27129,N_20674,N_22383);
and U27130 (N_27130,N_22651,N_21787);
or U27131 (N_27131,N_18358,N_21120);
and U27132 (N_27132,N_18163,N_19191);
or U27133 (N_27133,N_19417,N_19828);
or U27134 (N_27134,N_21447,N_18064);
nor U27135 (N_27135,N_22260,N_21042);
nor U27136 (N_27136,N_22170,N_20879);
and U27137 (N_27137,N_18305,N_18297);
or U27138 (N_27138,N_21785,N_22377);
and U27139 (N_27139,N_20021,N_20363);
nor U27140 (N_27140,N_21599,N_22935);
nor U27141 (N_27141,N_19007,N_23681);
and U27142 (N_27142,N_23328,N_18078);
and U27143 (N_27143,N_22533,N_22634);
xnor U27144 (N_27144,N_23877,N_22231);
and U27145 (N_27145,N_20957,N_20188);
and U27146 (N_27146,N_21864,N_18459);
nand U27147 (N_27147,N_22633,N_18931);
or U27148 (N_27148,N_23811,N_22480);
nor U27149 (N_27149,N_20995,N_23906);
nand U27150 (N_27150,N_19539,N_23625);
nor U27151 (N_27151,N_23762,N_21660);
or U27152 (N_27152,N_22874,N_18326);
xor U27153 (N_27153,N_23016,N_20432);
nor U27154 (N_27154,N_19349,N_19789);
nor U27155 (N_27155,N_18258,N_22369);
nor U27156 (N_27156,N_19901,N_21729);
nor U27157 (N_27157,N_21760,N_18477);
and U27158 (N_27158,N_22010,N_22046);
xnor U27159 (N_27159,N_21543,N_23309);
nand U27160 (N_27160,N_23922,N_18734);
and U27161 (N_27161,N_20586,N_18246);
nand U27162 (N_27162,N_23351,N_23816);
nand U27163 (N_27163,N_22568,N_22293);
nand U27164 (N_27164,N_21666,N_18458);
nand U27165 (N_27165,N_18299,N_21329);
nor U27166 (N_27166,N_18692,N_21407);
and U27167 (N_27167,N_19125,N_18069);
and U27168 (N_27168,N_21559,N_23925);
nand U27169 (N_27169,N_23170,N_19097);
or U27170 (N_27170,N_19924,N_19980);
or U27171 (N_27171,N_18569,N_19580);
nor U27172 (N_27172,N_22777,N_20428);
xor U27173 (N_27173,N_20718,N_22835);
nor U27174 (N_27174,N_20117,N_20189);
xnor U27175 (N_27175,N_20243,N_18500);
nand U27176 (N_27176,N_21579,N_22335);
and U27177 (N_27177,N_18114,N_22222);
nor U27178 (N_27178,N_18990,N_22926);
or U27179 (N_27179,N_18157,N_22795);
and U27180 (N_27180,N_20584,N_19449);
nand U27181 (N_27181,N_21812,N_21948);
xnor U27182 (N_27182,N_23935,N_22368);
xor U27183 (N_27183,N_20491,N_20592);
nor U27184 (N_27184,N_22442,N_22293);
nor U27185 (N_27185,N_20657,N_18981);
xor U27186 (N_27186,N_21828,N_19320);
or U27187 (N_27187,N_20742,N_22787);
or U27188 (N_27188,N_18919,N_22623);
nand U27189 (N_27189,N_19513,N_18319);
nor U27190 (N_27190,N_23374,N_19370);
and U27191 (N_27191,N_20929,N_22026);
nand U27192 (N_27192,N_18701,N_22527);
or U27193 (N_27193,N_21132,N_21743);
or U27194 (N_27194,N_22262,N_20666);
nor U27195 (N_27195,N_19912,N_18034);
xor U27196 (N_27196,N_22344,N_22044);
xnor U27197 (N_27197,N_22436,N_20901);
xnor U27198 (N_27198,N_22610,N_21199);
nor U27199 (N_27199,N_21715,N_19050);
nor U27200 (N_27200,N_22706,N_23749);
xnor U27201 (N_27201,N_18755,N_21547);
nand U27202 (N_27202,N_23468,N_18277);
and U27203 (N_27203,N_20035,N_19454);
nand U27204 (N_27204,N_23291,N_22918);
nand U27205 (N_27205,N_21174,N_18214);
and U27206 (N_27206,N_21218,N_20491);
or U27207 (N_27207,N_23778,N_21988);
nor U27208 (N_27208,N_20953,N_20239);
nand U27209 (N_27209,N_21557,N_19543);
nor U27210 (N_27210,N_19342,N_21738);
and U27211 (N_27211,N_22668,N_18224);
nor U27212 (N_27212,N_21340,N_19277);
or U27213 (N_27213,N_21450,N_20330);
nand U27214 (N_27214,N_19534,N_20170);
or U27215 (N_27215,N_20741,N_18317);
nand U27216 (N_27216,N_20536,N_21849);
nand U27217 (N_27217,N_19153,N_20462);
and U27218 (N_27218,N_18391,N_22586);
nor U27219 (N_27219,N_22739,N_19161);
xor U27220 (N_27220,N_19973,N_19665);
xor U27221 (N_27221,N_23233,N_19117);
and U27222 (N_27222,N_23223,N_23670);
nor U27223 (N_27223,N_20340,N_19461);
and U27224 (N_27224,N_22098,N_22072);
xor U27225 (N_27225,N_18588,N_18822);
nand U27226 (N_27226,N_20350,N_22971);
and U27227 (N_27227,N_18855,N_20233);
or U27228 (N_27228,N_22286,N_23152);
or U27229 (N_27229,N_21965,N_21500);
xnor U27230 (N_27230,N_18093,N_22849);
nand U27231 (N_27231,N_19622,N_23379);
nand U27232 (N_27232,N_18783,N_23625);
and U27233 (N_27233,N_18887,N_22485);
and U27234 (N_27234,N_20507,N_20869);
nand U27235 (N_27235,N_19141,N_18249);
and U27236 (N_27236,N_21326,N_23147);
xor U27237 (N_27237,N_19513,N_19074);
and U27238 (N_27238,N_21115,N_20661);
nor U27239 (N_27239,N_23117,N_20889);
and U27240 (N_27240,N_20287,N_18241);
xor U27241 (N_27241,N_18829,N_21413);
xor U27242 (N_27242,N_20296,N_18702);
and U27243 (N_27243,N_20420,N_22457);
and U27244 (N_27244,N_21585,N_19649);
xor U27245 (N_27245,N_21478,N_22979);
nand U27246 (N_27246,N_19058,N_22473);
xnor U27247 (N_27247,N_21146,N_20236);
nand U27248 (N_27248,N_18896,N_20599);
nor U27249 (N_27249,N_20343,N_21048);
nand U27250 (N_27250,N_18930,N_21247);
nand U27251 (N_27251,N_20053,N_18802);
nand U27252 (N_27252,N_23737,N_21222);
xor U27253 (N_27253,N_22449,N_21537);
nor U27254 (N_27254,N_21951,N_21702);
and U27255 (N_27255,N_20177,N_18079);
nand U27256 (N_27256,N_23205,N_22033);
nand U27257 (N_27257,N_21342,N_21818);
nand U27258 (N_27258,N_19466,N_22365);
xnor U27259 (N_27259,N_23947,N_20580);
or U27260 (N_27260,N_22408,N_23674);
nand U27261 (N_27261,N_21602,N_18424);
nor U27262 (N_27262,N_21612,N_18362);
xnor U27263 (N_27263,N_22019,N_19187);
xor U27264 (N_27264,N_20096,N_21937);
or U27265 (N_27265,N_18231,N_23875);
or U27266 (N_27266,N_23173,N_21098);
and U27267 (N_27267,N_22915,N_18028);
nor U27268 (N_27268,N_18161,N_23261);
nor U27269 (N_27269,N_18966,N_19489);
or U27270 (N_27270,N_23724,N_20818);
xor U27271 (N_27271,N_18459,N_18047);
nand U27272 (N_27272,N_22460,N_23459);
nor U27273 (N_27273,N_23837,N_18840);
nor U27274 (N_27274,N_20967,N_18530);
xnor U27275 (N_27275,N_19748,N_23056);
or U27276 (N_27276,N_22121,N_19940);
or U27277 (N_27277,N_19705,N_19976);
or U27278 (N_27278,N_21154,N_23109);
nand U27279 (N_27279,N_20805,N_21847);
or U27280 (N_27280,N_20840,N_22081);
nand U27281 (N_27281,N_20467,N_20555);
and U27282 (N_27282,N_20849,N_20751);
nor U27283 (N_27283,N_20020,N_23978);
nand U27284 (N_27284,N_22858,N_23164);
nor U27285 (N_27285,N_22766,N_18696);
xor U27286 (N_27286,N_22636,N_23439);
xnor U27287 (N_27287,N_18719,N_21501);
nor U27288 (N_27288,N_18128,N_20238);
xor U27289 (N_27289,N_21690,N_21272);
or U27290 (N_27290,N_20991,N_19107);
and U27291 (N_27291,N_21769,N_19842);
or U27292 (N_27292,N_23807,N_18041);
xor U27293 (N_27293,N_23639,N_22861);
nand U27294 (N_27294,N_23728,N_18889);
or U27295 (N_27295,N_22513,N_18120);
or U27296 (N_27296,N_21238,N_20847);
nor U27297 (N_27297,N_23709,N_21254);
nand U27298 (N_27298,N_19657,N_22358);
nor U27299 (N_27299,N_18722,N_19773);
nand U27300 (N_27300,N_18802,N_18979);
or U27301 (N_27301,N_23454,N_22261);
nand U27302 (N_27302,N_22260,N_22779);
or U27303 (N_27303,N_23618,N_18691);
and U27304 (N_27304,N_21135,N_21748);
or U27305 (N_27305,N_19818,N_21504);
nor U27306 (N_27306,N_19465,N_19292);
xnor U27307 (N_27307,N_21867,N_22657);
nor U27308 (N_27308,N_18765,N_22565);
xnor U27309 (N_27309,N_23361,N_20155);
and U27310 (N_27310,N_21867,N_19347);
nor U27311 (N_27311,N_20426,N_21662);
nand U27312 (N_27312,N_19267,N_22795);
or U27313 (N_27313,N_19090,N_23709);
nand U27314 (N_27314,N_18542,N_23743);
nor U27315 (N_27315,N_18315,N_20537);
xor U27316 (N_27316,N_19795,N_21138);
and U27317 (N_27317,N_23820,N_21901);
nand U27318 (N_27318,N_23264,N_23711);
or U27319 (N_27319,N_20633,N_23636);
and U27320 (N_27320,N_18556,N_18394);
or U27321 (N_27321,N_23797,N_21444);
nor U27322 (N_27322,N_18940,N_22195);
xnor U27323 (N_27323,N_23294,N_19937);
nor U27324 (N_27324,N_22466,N_23195);
or U27325 (N_27325,N_23491,N_18172);
or U27326 (N_27326,N_22644,N_21991);
nor U27327 (N_27327,N_20446,N_19698);
nor U27328 (N_27328,N_19430,N_21851);
or U27329 (N_27329,N_22539,N_19264);
and U27330 (N_27330,N_21491,N_21295);
and U27331 (N_27331,N_18290,N_18429);
nand U27332 (N_27332,N_19579,N_22715);
and U27333 (N_27333,N_20979,N_22845);
xnor U27334 (N_27334,N_21679,N_18580);
nand U27335 (N_27335,N_21484,N_19251);
nand U27336 (N_27336,N_22746,N_22601);
or U27337 (N_27337,N_22648,N_21849);
nor U27338 (N_27338,N_22463,N_22714);
nor U27339 (N_27339,N_22462,N_22344);
nand U27340 (N_27340,N_22379,N_23237);
and U27341 (N_27341,N_23666,N_22217);
nor U27342 (N_27342,N_20095,N_21543);
nor U27343 (N_27343,N_22527,N_21902);
or U27344 (N_27344,N_18761,N_21263);
nand U27345 (N_27345,N_21673,N_20672);
and U27346 (N_27346,N_23038,N_23711);
nor U27347 (N_27347,N_22398,N_22359);
or U27348 (N_27348,N_22837,N_21872);
nand U27349 (N_27349,N_21564,N_21722);
and U27350 (N_27350,N_20802,N_21144);
and U27351 (N_27351,N_19516,N_19110);
nand U27352 (N_27352,N_20997,N_21599);
xor U27353 (N_27353,N_18150,N_22421);
or U27354 (N_27354,N_18719,N_20155);
and U27355 (N_27355,N_22658,N_19614);
and U27356 (N_27356,N_22887,N_22311);
nor U27357 (N_27357,N_19905,N_23034);
nor U27358 (N_27358,N_20305,N_22318);
or U27359 (N_27359,N_23704,N_19207);
nor U27360 (N_27360,N_22167,N_23361);
nand U27361 (N_27361,N_19441,N_23539);
or U27362 (N_27362,N_20072,N_18850);
or U27363 (N_27363,N_19809,N_18282);
nor U27364 (N_27364,N_21461,N_23193);
or U27365 (N_27365,N_19265,N_22647);
or U27366 (N_27366,N_22606,N_21708);
or U27367 (N_27367,N_22210,N_21203);
and U27368 (N_27368,N_21395,N_20325);
nor U27369 (N_27369,N_19518,N_22784);
xnor U27370 (N_27370,N_21986,N_19890);
or U27371 (N_27371,N_19581,N_21700);
and U27372 (N_27372,N_18596,N_23830);
nor U27373 (N_27373,N_19215,N_19272);
xnor U27374 (N_27374,N_22592,N_21261);
nor U27375 (N_27375,N_19286,N_23754);
xor U27376 (N_27376,N_19487,N_19806);
and U27377 (N_27377,N_22307,N_22835);
xor U27378 (N_27378,N_20076,N_18612);
and U27379 (N_27379,N_21804,N_21717);
or U27380 (N_27380,N_23682,N_19358);
xnor U27381 (N_27381,N_22542,N_19414);
nand U27382 (N_27382,N_21740,N_19266);
nand U27383 (N_27383,N_23614,N_22137);
and U27384 (N_27384,N_21012,N_22931);
xor U27385 (N_27385,N_21189,N_18667);
and U27386 (N_27386,N_21916,N_23172);
nand U27387 (N_27387,N_20754,N_23733);
and U27388 (N_27388,N_23187,N_23763);
or U27389 (N_27389,N_19715,N_20567);
or U27390 (N_27390,N_23699,N_22825);
nand U27391 (N_27391,N_23417,N_20945);
nand U27392 (N_27392,N_20987,N_23192);
nand U27393 (N_27393,N_18431,N_22206);
and U27394 (N_27394,N_19960,N_20817);
nor U27395 (N_27395,N_20901,N_20175);
xnor U27396 (N_27396,N_22141,N_21300);
nor U27397 (N_27397,N_18048,N_20452);
nand U27398 (N_27398,N_21274,N_18472);
nand U27399 (N_27399,N_20489,N_19215);
and U27400 (N_27400,N_22534,N_22339);
nor U27401 (N_27401,N_22331,N_18818);
nor U27402 (N_27402,N_18918,N_20405);
and U27403 (N_27403,N_22139,N_20018);
and U27404 (N_27404,N_19669,N_23482);
and U27405 (N_27405,N_18848,N_22906);
and U27406 (N_27406,N_21580,N_22987);
nand U27407 (N_27407,N_21815,N_19569);
or U27408 (N_27408,N_19514,N_19390);
nand U27409 (N_27409,N_21447,N_20821);
nor U27410 (N_27410,N_19830,N_23951);
nand U27411 (N_27411,N_21082,N_20585);
nor U27412 (N_27412,N_19503,N_19402);
or U27413 (N_27413,N_20785,N_22102);
or U27414 (N_27414,N_23991,N_21479);
or U27415 (N_27415,N_19626,N_22205);
nand U27416 (N_27416,N_18131,N_19449);
xor U27417 (N_27417,N_21914,N_20106);
nand U27418 (N_27418,N_22709,N_18651);
nor U27419 (N_27419,N_20177,N_20730);
nor U27420 (N_27420,N_22033,N_22789);
or U27421 (N_27421,N_22896,N_18526);
and U27422 (N_27422,N_21579,N_22150);
nand U27423 (N_27423,N_21957,N_22045);
nor U27424 (N_27424,N_19296,N_22569);
and U27425 (N_27425,N_20054,N_21229);
xor U27426 (N_27426,N_18891,N_20015);
nand U27427 (N_27427,N_21944,N_19764);
and U27428 (N_27428,N_18730,N_21934);
xor U27429 (N_27429,N_20934,N_22731);
nand U27430 (N_27430,N_18597,N_21147);
or U27431 (N_27431,N_18972,N_22811);
nand U27432 (N_27432,N_22551,N_19886);
and U27433 (N_27433,N_19008,N_23165);
xor U27434 (N_27434,N_20289,N_18982);
and U27435 (N_27435,N_21806,N_18321);
or U27436 (N_27436,N_21927,N_22860);
nor U27437 (N_27437,N_22823,N_19086);
and U27438 (N_27438,N_22706,N_23014);
or U27439 (N_27439,N_18478,N_18841);
xnor U27440 (N_27440,N_20710,N_18152);
xnor U27441 (N_27441,N_18618,N_22738);
xor U27442 (N_27442,N_23011,N_21865);
nor U27443 (N_27443,N_18950,N_21855);
or U27444 (N_27444,N_20750,N_21426);
and U27445 (N_27445,N_22150,N_23036);
or U27446 (N_27446,N_21012,N_18204);
xor U27447 (N_27447,N_20544,N_20264);
nor U27448 (N_27448,N_22676,N_18135);
nand U27449 (N_27449,N_20589,N_21478);
nor U27450 (N_27450,N_23685,N_21938);
and U27451 (N_27451,N_23027,N_23099);
and U27452 (N_27452,N_23986,N_21842);
xor U27453 (N_27453,N_22116,N_23326);
and U27454 (N_27454,N_20182,N_23938);
nor U27455 (N_27455,N_18846,N_18101);
nor U27456 (N_27456,N_18220,N_21653);
nand U27457 (N_27457,N_23335,N_21311);
nor U27458 (N_27458,N_19027,N_22215);
and U27459 (N_27459,N_22971,N_23893);
nor U27460 (N_27460,N_20987,N_18624);
nor U27461 (N_27461,N_23902,N_18938);
and U27462 (N_27462,N_23288,N_19444);
nand U27463 (N_27463,N_23208,N_19992);
xnor U27464 (N_27464,N_18395,N_18881);
nor U27465 (N_27465,N_18864,N_20166);
xnor U27466 (N_27466,N_20230,N_18164);
nor U27467 (N_27467,N_23435,N_20890);
nand U27468 (N_27468,N_19222,N_22176);
xnor U27469 (N_27469,N_22062,N_19273);
xnor U27470 (N_27470,N_20716,N_23241);
or U27471 (N_27471,N_19235,N_22856);
xnor U27472 (N_27472,N_19661,N_20579);
nand U27473 (N_27473,N_22225,N_21306);
and U27474 (N_27474,N_21803,N_22183);
nor U27475 (N_27475,N_19365,N_23584);
xor U27476 (N_27476,N_20158,N_21501);
nand U27477 (N_27477,N_22247,N_20774);
nand U27478 (N_27478,N_23460,N_20533);
nor U27479 (N_27479,N_23013,N_20624);
nand U27480 (N_27480,N_19798,N_20646);
and U27481 (N_27481,N_21334,N_22568);
nand U27482 (N_27482,N_19046,N_20291);
nor U27483 (N_27483,N_19851,N_21653);
nand U27484 (N_27484,N_23389,N_21318);
nor U27485 (N_27485,N_21764,N_21533);
and U27486 (N_27486,N_19476,N_22909);
nor U27487 (N_27487,N_20878,N_19343);
nor U27488 (N_27488,N_19551,N_22862);
or U27489 (N_27489,N_20546,N_20721);
nor U27490 (N_27490,N_18080,N_22850);
or U27491 (N_27491,N_22084,N_23333);
nand U27492 (N_27492,N_20226,N_21501);
and U27493 (N_27493,N_20180,N_19126);
nor U27494 (N_27494,N_23342,N_19748);
or U27495 (N_27495,N_19649,N_22238);
and U27496 (N_27496,N_18561,N_21303);
xnor U27497 (N_27497,N_23449,N_20160);
nand U27498 (N_27498,N_20241,N_20390);
nand U27499 (N_27499,N_23445,N_19457);
nand U27500 (N_27500,N_23100,N_21743);
and U27501 (N_27501,N_21334,N_23352);
or U27502 (N_27502,N_23280,N_21250);
or U27503 (N_27503,N_18737,N_20429);
nor U27504 (N_27504,N_23011,N_20079);
nor U27505 (N_27505,N_21069,N_20773);
and U27506 (N_27506,N_18121,N_21159);
nand U27507 (N_27507,N_19138,N_19436);
and U27508 (N_27508,N_20321,N_21797);
nand U27509 (N_27509,N_22596,N_23197);
or U27510 (N_27510,N_21265,N_23615);
xnor U27511 (N_27511,N_21740,N_21817);
nand U27512 (N_27512,N_22849,N_18415);
or U27513 (N_27513,N_18119,N_19207);
nand U27514 (N_27514,N_21544,N_21939);
xnor U27515 (N_27515,N_21526,N_19836);
and U27516 (N_27516,N_23617,N_18584);
and U27517 (N_27517,N_19288,N_23116);
nor U27518 (N_27518,N_19690,N_22793);
xnor U27519 (N_27519,N_22201,N_22490);
or U27520 (N_27520,N_18537,N_21204);
nand U27521 (N_27521,N_23236,N_20829);
nand U27522 (N_27522,N_22297,N_20641);
nand U27523 (N_27523,N_18502,N_20013);
and U27524 (N_27524,N_19805,N_18841);
and U27525 (N_27525,N_21812,N_21867);
nor U27526 (N_27526,N_18574,N_19390);
nor U27527 (N_27527,N_19996,N_21269);
nand U27528 (N_27528,N_20292,N_18651);
nor U27529 (N_27529,N_20522,N_23005);
or U27530 (N_27530,N_18332,N_21531);
nand U27531 (N_27531,N_18429,N_21270);
xnor U27532 (N_27532,N_21738,N_20094);
nor U27533 (N_27533,N_23248,N_20018);
xnor U27534 (N_27534,N_20659,N_23493);
and U27535 (N_27535,N_20210,N_21991);
and U27536 (N_27536,N_19542,N_18830);
nand U27537 (N_27537,N_19313,N_23235);
nand U27538 (N_27538,N_20686,N_22857);
nor U27539 (N_27539,N_23458,N_19088);
nand U27540 (N_27540,N_18286,N_21048);
and U27541 (N_27541,N_21293,N_18407);
or U27542 (N_27542,N_19601,N_20010);
nor U27543 (N_27543,N_19341,N_21552);
nor U27544 (N_27544,N_19479,N_20581);
and U27545 (N_27545,N_19178,N_23222);
and U27546 (N_27546,N_21411,N_19527);
nand U27547 (N_27547,N_21949,N_22812);
nor U27548 (N_27548,N_20735,N_20903);
and U27549 (N_27549,N_19863,N_21053);
and U27550 (N_27550,N_20755,N_20553);
or U27551 (N_27551,N_21450,N_23563);
and U27552 (N_27552,N_23398,N_18334);
and U27553 (N_27553,N_23946,N_23824);
nor U27554 (N_27554,N_21897,N_20042);
or U27555 (N_27555,N_21510,N_18992);
xor U27556 (N_27556,N_18754,N_18549);
or U27557 (N_27557,N_22507,N_21009);
and U27558 (N_27558,N_21880,N_19253);
or U27559 (N_27559,N_20937,N_22463);
or U27560 (N_27560,N_20892,N_20381);
nand U27561 (N_27561,N_20880,N_22174);
or U27562 (N_27562,N_21719,N_18637);
and U27563 (N_27563,N_20667,N_20584);
or U27564 (N_27564,N_22763,N_23107);
or U27565 (N_27565,N_19850,N_19839);
nand U27566 (N_27566,N_21951,N_19669);
or U27567 (N_27567,N_22359,N_18100);
nand U27568 (N_27568,N_18392,N_22442);
nand U27569 (N_27569,N_22964,N_19881);
or U27570 (N_27570,N_22454,N_23844);
nand U27571 (N_27571,N_20952,N_20670);
nor U27572 (N_27572,N_23284,N_19923);
or U27573 (N_27573,N_23112,N_22530);
and U27574 (N_27574,N_18683,N_19855);
nor U27575 (N_27575,N_23784,N_22152);
nand U27576 (N_27576,N_22547,N_22271);
or U27577 (N_27577,N_21388,N_21560);
nor U27578 (N_27578,N_18578,N_21927);
nand U27579 (N_27579,N_21281,N_18699);
nand U27580 (N_27580,N_18028,N_20848);
xnor U27581 (N_27581,N_21836,N_18698);
or U27582 (N_27582,N_20242,N_21443);
nor U27583 (N_27583,N_23915,N_20776);
and U27584 (N_27584,N_19796,N_18405);
or U27585 (N_27585,N_19457,N_22355);
nor U27586 (N_27586,N_21311,N_21573);
nor U27587 (N_27587,N_21133,N_22787);
nand U27588 (N_27588,N_21578,N_19991);
and U27589 (N_27589,N_22864,N_19379);
and U27590 (N_27590,N_22599,N_19617);
or U27591 (N_27591,N_18118,N_23854);
nor U27592 (N_27592,N_19386,N_19760);
or U27593 (N_27593,N_21432,N_19627);
xnor U27594 (N_27594,N_21624,N_20665);
nor U27595 (N_27595,N_22199,N_23478);
nor U27596 (N_27596,N_19408,N_19288);
or U27597 (N_27597,N_21803,N_21924);
nor U27598 (N_27598,N_22306,N_22403);
xnor U27599 (N_27599,N_22873,N_22769);
nor U27600 (N_27600,N_19371,N_19664);
nor U27601 (N_27601,N_22685,N_22090);
xnor U27602 (N_27602,N_20554,N_21341);
or U27603 (N_27603,N_20027,N_18912);
and U27604 (N_27604,N_21908,N_18006);
and U27605 (N_27605,N_21529,N_23970);
or U27606 (N_27606,N_20567,N_18842);
and U27607 (N_27607,N_21416,N_20526);
xor U27608 (N_27608,N_19573,N_22298);
nand U27609 (N_27609,N_18049,N_19079);
nor U27610 (N_27610,N_23848,N_22802);
nor U27611 (N_27611,N_23997,N_21652);
xnor U27612 (N_27612,N_19999,N_20296);
xnor U27613 (N_27613,N_18352,N_23171);
nor U27614 (N_27614,N_23869,N_23525);
and U27615 (N_27615,N_23980,N_21406);
nand U27616 (N_27616,N_18324,N_18221);
or U27617 (N_27617,N_18879,N_19629);
nor U27618 (N_27618,N_23392,N_22146);
nand U27619 (N_27619,N_19876,N_19653);
nor U27620 (N_27620,N_23814,N_21896);
and U27621 (N_27621,N_20295,N_19905);
or U27622 (N_27622,N_20148,N_23767);
xor U27623 (N_27623,N_22147,N_23220);
and U27624 (N_27624,N_23474,N_23062);
nand U27625 (N_27625,N_18784,N_18421);
and U27626 (N_27626,N_21935,N_20714);
nand U27627 (N_27627,N_18011,N_19050);
and U27628 (N_27628,N_20238,N_22027);
and U27629 (N_27629,N_20305,N_22541);
and U27630 (N_27630,N_19931,N_20309);
xnor U27631 (N_27631,N_23686,N_23123);
nand U27632 (N_27632,N_22197,N_23127);
nand U27633 (N_27633,N_23289,N_20810);
nand U27634 (N_27634,N_22279,N_20775);
nand U27635 (N_27635,N_18265,N_21328);
nor U27636 (N_27636,N_23252,N_19290);
nor U27637 (N_27637,N_23841,N_18002);
and U27638 (N_27638,N_23072,N_22586);
and U27639 (N_27639,N_23382,N_20613);
and U27640 (N_27640,N_20944,N_18985);
or U27641 (N_27641,N_21534,N_18522);
nor U27642 (N_27642,N_20247,N_19652);
nor U27643 (N_27643,N_19776,N_23922);
or U27644 (N_27644,N_20780,N_18283);
and U27645 (N_27645,N_18373,N_21105);
and U27646 (N_27646,N_18851,N_19132);
nand U27647 (N_27647,N_22677,N_21744);
or U27648 (N_27648,N_20499,N_18942);
nand U27649 (N_27649,N_20844,N_18319);
xnor U27650 (N_27650,N_21931,N_20280);
or U27651 (N_27651,N_19605,N_18655);
or U27652 (N_27652,N_23266,N_23798);
and U27653 (N_27653,N_21390,N_18585);
or U27654 (N_27654,N_19836,N_21338);
nor U27655 (N_27655,N_22443,N_23615);
or U27656 (N_27656,N_21950,N_18695);
and U27657 (N_27657,N_22454,N_20884);
and U27658 (N_27658,N_19248,N_21444);
nor U27659 (N_27659,N_20375,N_23998);
xor U27660 (N_27660,N_23633,N_22620);
nand U27661 (N_27661,N_22556,N_18865);
xnor U27662 (N_27662,N_19403,N_20685);
nand U27663 (N_27663,N_23620,N_21327);
nand U27664 (N_27664,N_21111,N_21982);
nand U27665 (N_27665,N_18740,N_22741);
nor U27666 (N_27666,N_21751,N_20557);
nand U27667 (N_27667,N_21243,N_18646);
nand U27668 (N_27668,N_18027,N_22358);
nor U27669 (N_27669,N_23140,N_19094);
xnor U27670 (N_27670,N_23312,N_23201);
nor U27671 (N_27671,N_18054,N_18019);
or U27672 (N_27672,N_19907,N_23924);
or U27673 (N_27673,N_20583,N_22047);
nor U27674 (N_27674,N_22146,N_21633);
nand U27675 (N_27675,N_22173,N_21221);
xnor U27676 (N_27676,N_22225,N_20324);
and U27677 (N_27677,N_21778,N_21712);
xnor U27678 (N_27678,N_18775,N_23355);
xor U27679 (N_27679,N_18493,N_19169);
nor U27680 (N_27680,N_18410,N_21461);
nor U27681 (N_27681,N_18256,N_22258);
or U27682 (N_27682,N_18217,N_18959);
or U27683 (N_27683,N_21711,N_19232);
or U27684 (N_27684,N_20294,N_18279);
nand U27685 (N_27685,N_22623,N_20428);
nor U27686 (N_27686,N_22356,N_22191);
nor U27687 (N_27687,N_18296,N_20463);
nor U27688 (N_27688,N_18819,N_23822);
or U27689 (N_27689,N_21382,N_21344);
nand U27690 (N_27690,N_23530,N_20919);
nor U27691 (N_27691,N_18012,N_19134);
or U27692 (N_27692,N_23313,N_19656);
and U27693 (N_27693,N_21260,N_21355);
or U27694 (N_27694,N_23459,N_18032);
and U27695 (N_27695,N_18658,N_21156);
nand U27696 (N_27696,N_18528,N_22395);
and U27697 (N_27697,N_23035,N_22744);
or U27698 (N_27698,N_20025,N_20624);
nor U27699 (N_27699,N_19522,N_23021);
nor U27700 (N_27700,N_18893,N_18765);
nor U27701 (N_27701,N_19658,N_21871);
nor U27702 (N_27702,N_21077,N_21425);
nor U27703 (N_27703,N_20537,N_21155);
nand U27704 (N_27704,N_21140,N_21791);
and U27705 (N_27705,N_23021,N_20414);
and U27706 (N_27706,N_19999,N_18753);
nor U27707 (N_27707,N_20484,N_23474);
and U27708 (N_27708,N_19270,N_20675);
nor U27709 (N_27709,N_20466,N_20970);
nor U27710 (N_27710,N_20644,N_21890);
nor U27711 (N_27711,N_20079,N_22714);
nor U27712 (N_27712,N_23533,N_21734);
nor U27713 (N_27713,N_21889,N_21177);
and U27714 (N_27714,N_20922,N_23782);
xnor U27715 (N_27715,N_21483,N_22885);
or U27716 (N_27716,N_21807,N_21625);
nor U27717 (N_27717,N_21621,N_18957);
or U27718 (N_27718,N_18576,N_19684);
nor U27719 (N_27719,N_20706,N_20366);
nand U27720 (N_27720,N_23846,N_21414);
and U27721 (N_27721,N_23754,N_21836);
and U27722 (N_27722,N_23933,N_22442);
nand U27723 (N_27723,N_18800,N_20741);
nand U27724 (N_27724,N_18764,N_18773);
nand U27725 (N_27725,N_23195,N_21414);
or U27726 (N_27726,N_22915,N_18151);
xor U27727 (N_27727,N_20250,N_19838);
and U27728 (N_27728,N_21346,N_18120);
nor U27729 (N_27729,N_21186,N_22095);
nor U27730 (N_27730,N_18247,N_20810);
or U27731 (N_27731,N_20734,N_21124);
nand U27732 (N_27732,N_21974,N_20904);
and U27733 (N_27733,N_23647,N_20789);
and U27734 (N_27734,N_20343,N_22609);
or U27735 (N_27735,N_20235,N_20660);
and U27736 (N_27736,N_20503,N_21420);
nor U27737 (N_27737,N_22058,N_18267);
nor U27738 (N_27738,N_19470,N_23730);
nor U27739 (N_27739,N_21674,N_23594);
xnor U27740 (N_27740,N_18519,N_18234);
xnor U27741 (N_27741,N_18738,N_23751);
nor U27742 (N_27742,N_23853,N_22496);
or U27743 (N_27743,N_18998,N_18044);
and U27744 (N_27744,N_21823,N_21615);
nor U27745 (N_27745,N_23498,N_19298);
or U27746 (N_27746,N_22486,N_20768);
nand U27747 (N_27747,N_21635,N_21097);
nand U27748 (N_27748,N_23196,N_19320);
or U27749 (N_27749,N_19933,N_20986);
and U27750 (N_27750,N_20462,N_18644);
or U27751 (N_27751,N_21926,N_21719);
nor U27752 (N_27752,N_22840,N_23128);
nand U27753 (N_27753,N_22651,N_22023);
xor U27754 (N_27754,N_23412,N_23222);
xnor U27755 (N_27755,N_23263,N_19112);
and U27756 (N_27756,N_22489,N_22721);
nand U27757 (N_27757,N_20088,N_21570);
xor U27758 (N_27758,N_18248,N_22518);
or U27759 (N_27759,N_18625,N_18707);
xnor U27760 (N_27760,N_20886,N_21966);
nand U27761 (N_27761,N_18136,N_21463);
nor U27762 (N_27762,N_20682,N_19809);
xor U27763 (N_27763,N_22389,N_19300);
nor U27764 (N_27764,N_18120,N_22025);
or U27765 (N_27765,N_21622,N_19384);
nor U27766 (N_27766,N_19805,N_18849);
or U27767 (N_27767,N_21321,N_19913);
nor U27768 (N_27768,N_22165,N_20162);
or U27769 (N_27769,N_22862,N_18215);
nor U27770 (N_27770,N_18166,N_18556);
and U27771 (N_27771,N_23253,N_23407);
nor U27772 (N_27772,N_18186,N_20295);
or U27773 (N_27773,N_18054,N_20111);
or U27774 (N_27774,N_22205,N_19981);
nor U27775 (N_27775,N_19198,N_18915);
nand U27776 (N_27776,N_22974,N_22086);
or U27777 (N_27777,N_22695,N_20766);
nand U27778 (N_27778,N_20475,N_22634);
and U27779 (N_27779,N_23865,N_19007);
or U27780 (N_27780,N_20791,N_19983);
and U27781 (N_27781,N_20563,N_20634);
and U27782 (N_27782,N_19478,N_23043);
nand U27783 (N_27783,N_19053,N_22577);
and U27784 (N_27784,N_22445,N_19361);
nor U27785 (N_27785,N_23142,N_21936);
nand U27786 (N_27786,N_18760,N_22642);
nand U27787 (N_27787,N_19739,N_23231);
nor U27788 (N_27788,N_21115,N_21531);
and U27789 (N_27789,N_18525,N_22296);
or U27790 (N_27790,N_23806,N_23183);
nand U27791 (N_27791,N_18900,N_21849);
nand U27792 (N_27792,N_21773,N_19323);
and U27793 (N_27793,N_20268,N_21709);
or U27794 (N_27794,N_20928,N_18594);
and U27795 (N_27795,N_23870,N_20751);
or U27796 (N_27796,N_20884,N_20995);
and U27797 (N_27797,N_23753,N_20160);
or U27798 (N_27798,N_20174,N_23360);
nor U27799 (N_27799,N_21093,N_19938);
xnor U27800 (N_27800,N_23346,N_18792);
and U27801 (N_27801,N_22336,N_20871);
or U27802 (N_27802,N_22708,N_23932);
and U27803 (N_27803,N_18246,N_22227);
and U27804 (N_27804,N_22315,N_21606);
nor U27805 (N_27805,N_20502,N_18678);
nor U27806 (N_27806,N_22615,N_18450);
nand U27807 (N_27807,N_23102,N_20600);
or U27808 (N_27808,N_19278,N_20982);
nand U27809 (N_27809,N_21241,N_20960);
and U27810 (N_27810,N_20306,N_21975);
or U27811 (N_27811,N_19439,N_18341);
or U27812 (N_27812,N_21032,N_18715);
and U27813 (N_27813,N_19925,N_21797);
or U27814 (N_27814,N_23489,N_22893);
nor U27815 (N_27815,N_18430,N_23358);
nand U27816 (N_27816,N_19181,N_23462);
or U27817 (N_27817,N_19579,N_22734);
xor U27818 (N_27818,N_20571,N_19917);
nand U27819 (N_27819,N_20868,N_23827);
nor U27820 (N_27820,N_19627,N_22075);
nand U27821 (N_27821,N_22399,N_19305);
or U27822 (N_27822,N_23595,N_21344);
xor U27823 (N_27823,N_19038,N_22569);
nor U27824 (N_27824,N_21930,N_18417);
and U27825 (N_27825,N_20987,N_21466);
or U27826 (N_27826,N_19666,N_22483);
nor U27827 (N_27827,N_18368,N_23754);
and U27828 (N_27828,N_18757,N_18815);
and U27829 (N_27829,N_20331,N_20340);
nand U27830 (N_27830,N_19742,N_23612);
or U27831 (N_27831,N_21555,N_19676);
or U27832 (N_27832,N_19210,N_22303);
nand U27833 (N_27833,N_18903,N_23310);
nand U27834 (N_27834,N_21494,N_22501);
or U27835 (N_27835,N_20566,N_23365);
xnor U27836 (N_27836,N_23648,N_22400);
or U27837 (N_27837,N_20079,N_21905);
and U27838 (N_27838,N_19011,N_23191);
nand U27839 (N_27839,N_18615,N_18944);
nand U27840 (N_27840,N_18927,N_21848);
nand U27841 (N_27841,N_21880,N_20989);
xor U27842 (N_27842,N_23028,N_23479);
nor U27843 (N_27843,N_22051,N_20890);
nand U27844 (N_27844,N_18013,N_23195);
nor U27845 (N_27845,N_19792,N_23641);
nor U27846 (N_27846,N_21442,N_18187);
nand U27847 (N_27847,N_18075,N_23062);
nor U27848 (N_27848,N_22787,N_18930);
xor U27849 (N_27849,N_18870,N_21441);
nand U27850 (N_27850,N_20366,N_23199);
or U27851 (N_27851,N_20158,N_22087);
nor U27852 (N_27852,N_18989,N_22456);
and U27853 (N_27853,N_18696,N_20240);
nor U27854 (N_27854,N_18155,N_23804);
and U27855 (N_27855,N_19036,N_19770);
and U27856 (N_27856,N_19877,N_22785);
or U27857 (N_27857,N_21057,N_22728);
nand U27858 (N_27858,N_23647,N_21694);
and U27859 (N_27859,N_23067,N_18845);
or U27860 (N_27860,N_23524,N_18708);
nand U27861 (N_27861,N_19429,N_23368);
nand U27862 (N_27862,N_21915,N_18296);
nor U27863 (N_27863,N_22062,N_21574);
nor U27864 (N_27864,N_18711,N_23854);
or U27865 (N_27865,N_22444,N_21495);
nand U27866 (N_27866,N_21554,N_20247);
nand U27867 (N_27867,N_22325,N_23038);
or U27868 (N_27868,N_20722,N_19956);
nand U27869 (N_27869,N_19440,N_23158);
or U27870 (N_27870,N_21029,N_18366);
and U27871 (N_27871,N_23833,N_22694);
or U27872 (N_27872,N_20424,N_20023);
or U27873 (N_27873,N_20350,N_18382);
and U27874 (N_27874,N_20964,N_23663);
and U27875 (N_27875,N_18474,N_23460);
or U27876 (N_27876,N_19830,N_20892);
and U27877 (N_27877,N_18395,N_21985);
and U27878 (N_27878,N_20592,N_20295);
or U27879 (N_27879,N_22107,N_22677);
or U27880 (N_27880,N_21921,N_20739);
xor U27881 (N_27881,N_19597,N_22753);
and U27882 (N_27882,N_20806,N_21435);
xnor U27883 (N_27883,N_20993,N_23713);
xor U27884 (N_27884,N_21262,N_21740);
xor U27885 (N_27885,N_18680,N_18628);
nand U27886 (N_27886,N_19115,N_19871);
nand U27887 (N_27887,N_20424,N_20722);
xor U27888 (N_27888,N_22900,N_21385);
nand U27889 (N_27889,N_18321,N_21501);
or U27890 (N_27890,N_21125,N_21885);
or U27891 (N_27891,N_23996,N_22882);
or U27892 (N_27892,N_19922,N_21878);
or U27893 (N_27893,N_19076,N_21217);
nor U27894 (N_27894,N_21215,N_23760);
nand U27895 (N_27895,N_19424,N_23763);
nor U27896 (N_27896,N_20166,N_21787);
xor U27897 (N_27897,N_23827,N_20061);
nand U27898 (N_27898,N_23312,N_20221);
nor U27899 (N_27899,N_18446,N_21466);
and U27900 (N_27900,N_20165,N_21158);
or U27901 (N_27901,N_19892,N_22019);
nor U27902 (N_27902,N_23798,N_22747);
nand U27903 (N_27903,N_23786,N_22266);
or U27904 (N_27904,N_23272,N_21431);
nor U27905 (N_27905,N_19575,N_22458);
nand U27906 (N_27906,N_20352,N_18477);
nor U27907 (N_27907,N_22269,N_19930);
and U27908 (N_27908,N_18553,N_23334);
nand U27909 (N_27909,N_18848,N_22140);
and U27910 (N_27910,N_19526,N_22968);
xnor U27911 (N_27911,N_18369,N_20418);
nand U27912 (N_27912,N_18010,N_20318);
nor U27913 (N_27913,N_20170,N_21876);
or U27914 (N_27914,N_20164,N_20665);
or U27915 (N_27915,N_21212,N_19874);
nor U27916 (N_27916,N_21083,N_20721);
and U27917 (N_27917,N_20770,N_18244);
nand U27918 (N_27918,N_22075,N_22514);
nand U27919 (N_27919,N_19732,N_23539);
nor U27920 (N_27920,N_22853,N_23342);
nor U27921 (N_27921,N_21997,N_18040);
or U27922 (N_27922,N_20428,N_22595);
xnor U27923 (N_27923,N_23765,N_22907);
xor U27924 (N_27924,N_20919,N_19418);
or U27925 (N_27925,N_19576,N_21376);
and U27926 (N_27926,N_22385,N_20641);
and U27927 (N_27927,N_21750,N_21338);
or U27928 (N_27928,N_22091,N_22160);
or U27929 (N_27929,N_21958,N_20762);
nor U27930 (N_27930,N_19949,N_19911);
and U27931 (N_27931,N_20414,N_22389);
and U27932 (N_27932,N_22682,N_23584);
and U27933 (N_27933,N_20885,N_20293);
nor U27934 (N_27934,N_21398,N_22026);
xor U27935 (N_27935,N_23295,N_21853);
or U27936 (N_27936,N_22778,N_20190);
or U27937 (N_27937,N_19906,N_23817);
nor U27938 (N_27938,N_20883,N_19083);
xor U27939 (N_27939,N_19927,N_20599);
xor U27940 (N_27940,N_18396,N_23608);
nor U27941 (N_27941,N_23267,N_21691);
nand U27942 (N_27942,N_19735,N_23598);
and U27943 (N_27943,N_20066,N_20467);
nor U27944 (N_27944,N_20775,N_18599);
and U27945 (N_27945,N_18724,N_18111);
or U27946 (N_27946,N_21493,N_23439);
or U27947 (N_27947,N_23696,N_23678);
and U27948 (N_27948,N_18267,N_19036);
nor U27949 (N_27949,N_18718,N_22821);
nand U27950 (N_27950,N_22525,N_23811);
nand U27951 (N_27951,N_22918,N_21167);
nand U27952 (N_27952,N_19015,N_23980);
nand U27953 (N_27953,N_22701,N_20556);
or U27954 (N_27954,N_20002,N_19129);
or U27955 (N_27955,N_19678,N_20685);
and U27956 (N_27956,N_19476,N_23563);
nand U27957 (N_27957,N_19987,N_20907);
and U27958 (N_27958,N_20663,N_20551);
nor U27959 (N_27959,N_23657,N_18290);
nor U27960 (N_27960,N_20835,N_21969);
nand U27961 (N_27961,N_19569,N_23004);
nor U27962 (N_27962,N_21692,N_23100);
nand U27963 (N_27963,N_22465,N_19464);
nor U27964 (N_27964,N_23605,N_22088);
and U27965 (N_27965,N_23142,N_19248);
or U27966 (N_27966,N_20153,N_19215);
or U27967 (N_27967,N_21555,N_22348);
nand U27968 (N_27968,N_22112,N_21069);
or U27969 (N_27969,N_21661,N_19239);
nand U27970 (N_27970,N_20162,N_23664);
or U27971 (N_27971,N_23921,N_22901);
nand U27972 (N_27972,N_20797,N_23282);
xor U27973 (N_27973,N_22089,N_18817);
and U27974 (N_27974,N_19956,N_21178);
and U27975 (N_27975,N_20868,N_22706);
xnor U27976 (N_27976,N_21480,N_18086);
nand U27977 (N_27977,N_20582,N_18346);
nand U27978 (N_27978,N_18055,N_20627);
nor U27979 (N_27979,N_22847,N_19561);
or U27980 (N_27980,N_19057,N_18770);
and U27981 (N_27981,N_19623,N_18391);
or U27982 (N_27982,N_22921,N_18303);
or U27983 (N_27983,N_18425,N_19587);
nor U27984 (N_27984,N_20743,N_18159);
or U27985 (N_27985,N_19571,N_19580);
xor U27986 (N_27986,N_23148,N_18488);
nor U27987 (N_27987,N_18260,N_18854);
and U27988 (N_27988,N_19397,N_19880);
nor U27989 (N_27989,N_23428,N_23465);
nor U27990 (N_27990,N_20906,N_22386);
or U27991 (N_27991,N_22985,N_23249);
or U27992 (N_27992,N_21304,N_21993);
or U27993 (N_27993,N_18067,N_23783);
nand U27994 (N_27994,N_23180,N_21496);
nand U27995 (N_27995,N_21851,N_20785);
nor U27996 (N_27996,N_21830,N_18997);
or U27997 (N_27997,N_18244,N_22246);
xor U27998 (N_27998,N_20683,N_21019);
nor U27999 (N_27999,N_21821,N_23605);
nand U28000 (N_28000,N_21476,N_23065);
nor U28001 (N_28001,N_18934,N_20120);
nand U28002 (N_28002,N_20800,N_20775);
nor U28003 (N_28003,N_19648,N_20981);
and U28004 (N_28004,N_22475,N_23619);
nand U28005 (N_28005,N_21007,N_18287);
or U28006 (N_28006,N_20020,N_22332);
nor U28007 (N_28007,N_21264,N_22931);
or U28008 (N_28008,N_18863,N_23526);
or U28009 (N_28009,N_21419,N_19505);
nand U28010 (N_28010,N_21262,N_23921);
nor U28011 (N_28011,N_18787,N_18909);
nand U28012 (N_28012,N_22446,N_21063);
or U28013 (N_28013,N_21712,N_22388);
and U28014 (N_28014,N_20460,N_23309);
or U28015 (N_28015,N_19663,N_21914);
xnor U28016 (N_28016,N_20222,N_21086);
nand U28017 (N_28017,N_18080,N_22776);
or U28018 (N_28018,N_18011,N_21763);
nor U28019 (N_28019,N_20531,N_19299);
nand U28020 (N_28020,N_19596,N_18558);
nor U28021 (N_28021,N_22999,N_21118);
and U28022 (N_28022,N_18496,N_18486);
or U28023 (N_28023,N_20059,N_20836);
or U28024 (N_28024,N_21846,N_20681);
or U28025 (N_28025,N_21093,N_19999);
nor U28026 (N_28026,N_23890,N_19160);
nand U28027 (N_28027,N_21117,N_20006);
nor U28028 (N_28028,N_19923,N_23449);
or U28029 (N_28029,N_19912,N_20447);
and U28030 (N_28030,N_18589,N_21519);
nor U28031 (N_28031,N_19949,N_21129);
nor U28032 (N_28032,N_20841,N_22945);
and U28033 (N_28033,N_21194,N_22573);
nand U28034 (N_28034,N_22772,N_18140);
and U28035 (N_28035,N_21277,N_20388);
nor U28036 (N_28036,N_18923,N_22689);
and U28037 (N_28037,N_18085,N_18081);
or U28038 (N_28038,N_20324,N_23398);
nor U28039 (N_28039,N_19218,N_20192);
and U28040 (N_28040,N_22393,N_21572);
nor U28041 (N_28041,N_18084,N_23205);
and U28042 (N_28042,N_21275,N_18753);
and U28043 (N_28043,N_20812,N_23549);
nand U28044 (N_28044,N_22699,N_20983);
or U28045 (N_28045,N_20420,N_18580);
nor U28046 (N_28046,N_20665,N_23095);
and U28047 (N_28047,N_19337,N_20734);
nand U28048 (N_28048,N_21996,N_19792);
nor U28049 (N_28049,N_23881,N_21934);
nand U28050 (N_28050,N_19244,N_22497);
or U28051 (N_28051,N_21238,N_20928);
xor U28052 (N_28052,N_21136,N_20508);
or U28053 (N_28053,N_18743,N_18302);
nor U28054 (N_28054,N_22293,N_19338);
and U28055 (N_28055,N_22031,N_20783);
nand U28056 (N_28056,N_20394,N_23456);
nor U28057 (N_28057,N_19208,N_21214);
or U28058 (N_28058,N_19823,N_19153);
nor U28059 (N_28059,N_22285,N_21336);
xnor U28060 (N_28060,N_23989,N_19468);
xnor U28061 (N_28061,N_20089,N_22201);
and U28062 (N_28062,N_22355,N_23442);
nand U28063 (N_28063,N_22178,N_22153);
xnor U28064 (N_28064,N_21211,N_18048);
nand U28065 (N_28065,N_19008,N_22200);
or U28066 (N_28066,N_20607,N_22014);
nand U28067 (N_28067,N_20846,N_23722);
or U28068 (N_28068,N_19617,N_20119);
nor U28069 (N_28069,N_20215,N_23779);
xnor U28070 (N_28070,N_19916,N_19698);
and U28071 (N_28071,N_19854,N_23658);
nand U28072 (N_28072,N_22504,N_22616);
nor U28073 (N_28073,N_18438,N_18196);
nand U28074 (N_28074,N_22228,N_22222);
nand U28075 (N_28075,N_21046,N_20936);
and U28076 (N_28076,N_18537,N_18840);
xor U28077 (N_28077,N_20436,N_21363);
xnor U28078 (N_28078,N_22717,N_21049);
or U28079 (N_28079,N_19951,N_19963);
nor U28080 (N_28080,N_23919,N_19796);
xnor U28081 (N_28081,N_19634,N_18885);
and U28082 (N_28082,N_18821,N_20210);
nand U28083 (N_28083,N_23582,N_23029);
and U28084 (N_28084,N_23826,N_20287);
or U28085 (N_28085,N_19930,N_21471);
xnor U28086 (N_28086,N_21361,N_18787);
and U28087 (N_28087,N_21207,N_19006);
xnor U28088 (N_28088,N_18251,N_21801);
nor U28089 (N_28089,N_19152,N_18748);
nand U28090 (N_28090,N_19207,N_22204);
and U28091 (N_28091,N_19230,N_23724);
or U28092 (N_28092,N_21392,N_20006);
and U28093 (N_28093,N_20072,N_22882);
and U28094 (N_28094,N_22178,N_21993);
nor U28095 (N_28095,N_23656,N_19065);
nand U28096 (N_28096,N_19412,N_20832);
nand U28097 (N_28097,N_20079,N_22120);
nand U28098 (N_28098,N_22352,N_20371);
and U28099 (N_28099,N_22754,N_19159);
and U28100 (N_28100,N_20528,N_19130);
nand U28101 (N_28101,N_19154,N_20905);
nor U28102 (N_28102,N_21193,N_19867);
nor U28103 (N_28103,N_18608,N_18086);
nor U28104 (N_28104,N_20792,N_23002);
nor U28105 (N_28105,N_22227,N_18474);
nor U28106 (N_28106,N_19223,N_21657);
nor U28107 (N_28107,N_23299,N_21764);
xor U28108 (N_28108,N_20865,N_21428);
xor U28109 (N_28109,N_19127,N_19834);
nand U28110 (N_28110,N_20408,N_22374);
and U28111 (N_28111,N_20047,N_18617);
nand U28112 (N_28112,N_19653,N_23529);
and U28113 (N_28113,N_18734,N_20055);
nand U28114 (N_28114,N_18132,N_23408);
xor U28115 (N_28115,N_20619,N_19356);
nand U28116 (N_28116,N_22012,N_22431);
or U28117 (N_28117,N_20414,N_18216);
and U28118 (N_28118,N_21149,N_20464);
and U28119 (N_28119,N_21196,N_20255);
nand U28120 (N_28120,N_22508,N_22229);
and U28121 (N_28121,N_18907,N_19301);
and U28122 (N_28122,N_21105,N_19900);
xor U28123 (N_28123,N_23212,N_22695);
nand U28124 (N_28124,N_21243,N_22331);
nor U28125 (N_28125,N_23240,N_22138);
nand U28126 (N_28126,N_22988,N_21930);
or U28127 (N_28127,N_18324,N_23662);
or U28128 (N_28128,N_21895,N_18450);
xnor U28129 (N_28129,N_18138,N_20790);
or U28130 (N_28130,N_23928,N_20304);
and U28131 (N_28131,N_19865,N_21927);
or U28132 (N_28132,N_23301,N_22195);
nand U28133 (N_28133,N_20581,N_18919);
nor U28134 (N_28134,N_23230,N_23886);
xor U28135 (N_28135,N_22898,N_22680);
nand U28136 (N_28136,N_18775,N_20874);
or U28137 (N_28137,N_21967,N_19886);
or U28138 (N_28138,N_23273,N_22907);
nor U28139 (N_28139,N_23788,N_20728);
and U28140 (N_28140,N_23407,N_19259);
nor U28141 (N_28141,N_19538,N_23995);
xnor U28142 (N_28142,N_21212,N_18444);
nor U28143 (N_28143,N_20229,N_19896);
nor U28144 (N_28144,N_22380,N_22702);
or U28145 (N_28145,N_20121,N_23555);
and U28146 (N_28146,N_18219,N_19952);
and U28147 (N_28147,N_22164,N_20090);
and U28148 (N_28148,N_18148,N_20566);
nor U28149 (N_28149,N_18494,N_18904);
or U28150 (N_28150,N_19458,N_21127);
and U28151 (N_28151,N_20760,N_19922);
nand U28152 (N_28152,N_18839,N_22301);
or U28153 (N_28153,N_22321,N_23284);
nor U28154 (N_28154,N_22952,N_20643);
or U28155 (N_28155,N_19877,N_23665);
nor U28156 (N_28156,N_18185,N_18566);
xor U28157 (N_28157,N_20108,N_19961);
and U28158 (N_28158,N_19722,N_21812);
or U28159 (N_28159,N_21211,N_22699);
and U28160 (N_28160,N_18944,N_22944);
nand U28161 (N_28161,N_19542,N_20030);
or U28162 (N_28162,N_22018,N_21808);
nor U28163 (N_28163,N_20010,N_19792);
or U28164 (N_28164,N_18365,N_22232);
and U28165 (N_28165,N_23026,N_22960);
or U28166 (N_28166,N_19277,N_22717);
or U28167 (N_28167,N_21574,N_21239);
nor U28168 (N_28168,N_22138,N_23311);
or U28169 (N_28169,N_22972,N_22195);
nand U28170 (N_28170,N_20403,N_19361);
or U28171 (N_28171,N_18643,N_21053);
nand U28172 (N_28172,N_19223,N_18897);
xnor U28173 (N_28173,N_22380,N_19777);
nand U28174 (N_28174,N_19418,N_18298);
nand U28175 (N_28175,N_18565,N_19672);
nor U28176 (N_28176,N_19241,N_20129);
or U28177 (N_28177,N_22636,N_22648);
or U28178 (N_28178,N_20147,N_18771);
nand U28179 (N_28179,N_19130,N_21524);
xnor U28180 (N_28180,N_19345,N_18331);
nor U28181 (N_28181,N_18856,N_23803);
nand U28182 (N_28182,N_18594,N_23175);
and U28183 (N_28183,N_18744,N_19517);
nor U28184 (N_28184,N_19827,N_19125);
and U28185 (N_28185,N_21025,N_18971);
nor U28186 (N_28186,N_18402,N_20171);
or U28187 (N_28187,N_18515,N_20894);
nand U28188 (N_28188,N_21755,N_19162);
and U28189 (N_28189,N_22801,N_21176);
xor U28190 (N_28190,N_21266,N_20294);
nor U28191 (N_28191,N_20694,N_22110);
and U28192 (N_28192,N_23245,N_22077);
or U28193 (N_28193,N_20524,N_22480);
nand U28194 (N_28194,N_20740,N_22884);
nand U28195 (N_28195,N_23752,N_22867);
nand U28196 (N_28196,N_18958,N_19006);
nor U28197 (N_28197,N_22528,N_22050);
nor U28198 (N_28198,N_23871,N_19316);
nand U28199 (N_28199,N_20407,N_20896);
nand U28200 (N_28200,N_19785,N_23497);
xnor U28201 (N_28201,N_22621,N_22242);
nor U28202 (N_28202,N_19131,N_19915);
and U28203 (N_28203,N_21400,N_23515);
and U28204 (N_28204,N_18430,N_23419);
or U28205 (N_28205,N_19133,N_22566);
or U28206 (N_28206,N_21443,N_23955);
nor U28207 (N_28207,N_19521,N_18708);
nor U28208 (N_28208,N_20076,N_21737);
nor U28209 (N_28209,N_20887,N_19517);
nor U28210 (N_28210,N_22283,N_22077);
nor U28211 (N_28211,N_18175,N_21076);
nand U28212 (N_28212,N_23388,N_21124);
nand U28213 (N_28213,N_19925,N_22289);
and U28214 (N_28214,N_18875,N_20703);
nand U28215 (N_28215,N_21802,N_20142);
or U28216 (N_28216,N_21091,N_20213);
nand U28217 (N_28217,N_19196,N_23868);
nor U28218 (N_28218,N_23093,N_22624);
xnor U28219 (N_28219,N_20188,N_20641);
and U28220 (N_28220,N_23907,N_18190);
or U28221 (N_28221,N_22846,N_19791);
or U28222 (N_28222,N_19261,N_20419);
or U28223 (N_28223,N_23801,N_21010);
xor U28224 (N_28224,N_19592,N_23764);
nand U28225 (N_28225,N_22229,N_19036);
nor U28226 (N_28226,N_19248,N_20149);
nor U28227 (N_28227,N_20469,N_22475);
or U28228 (N_28228,N_23724,N_23052);
nor U28229 (N_28229,N_22302,N_18436);
nand U28230 (N_28230,N_18364,N_20042);
nor U28231 (N_28231,N_19525,N_20498);
and U28232 (N_28232,N_22112,N_21854);
nor U28233 (N_28233,N_20955,N_22065);
or U28234 (N_28234,N_22141,N_19088);
nand U28235 (N_28235,N_20418,N_23251);
and U28236 (N_28236,N_21888,N_23153);
or U28237 (N_28237,N_23497,N_21016);
and U28238 (N_28238,N_21643,N_20833);
or U28239 (N_28239,N_20282,N_23684);
nand U28240 (N_28240,N_20976,N_21093);
nor U28241 (N_28241,N_19895,N_22044);
or U28242 (N_28242,N_21547,N_23517);
nor U28243 (N_28243,N_23451,N_22797);
or U28244 (N_28244,N_22513,N_20452);
or U28245 (N_28245,N_22954,N_22530);
nor U28246 (N_28246,N_22520,N_21678);
and U28247 (N_28247,N_20914,N_23301);
and U28248 (N_28248,N_23744,N_20878);
nor U28249 (N_28249,N_23377,N_20495);
xor U28250 (N_28250,N_18294,N_23671);
and U28251 (N_28251,N_18789,N_21799);
and U28252 (N_28252,N_18183,N_23060);
nor U28253 (N_28253,N_22646,N_20174);
xnor U28254 (N_28254,N_18806,N_18635);
nor U28255 (N_28255,N_23126,N_19487);
nor U28256 (N_28256,N_22514,N_19360);
nand U28257 (N_28257,N_23838,N_19191);
and U28258 (N_28258,N_22457,N_18359);
and U28259 (N_28259,N_18103,N_19605);
or U28260 (N_28260,N_23137,N_23217);
or U28261 (N_28261,N_23045,N_19480);
or U28262 (N_28262,N_20422,N_23833);
nand U28263 (N_28263,N_18101,N_21183);
xnor U28264 (N_28264,N_23428,N_22198);
or U28265 (N_28265,N_20703,N_20539);
or U28266 (N_28266,N_19085,N_18665);
nand U28267 (N_28267,N_22659,N_23990);
xor U28268 (N_28268,N_19840,N_21916);
and U28269 (N_28269,N_23294,N_20540);
or U28270 (N_28270,N_19488,N_18691);
nor U28271 (N_28271,N_21441,N_19812);
or U28272 (N_28272,N_23485,N_22720);
or U28273 (N_28273,N_18730,N_18434);
or U28274 (N_28274,N_21188,N_23186);
and U28275 (N_28275,N_20174,N_20018);
nor U28276 (N_28276,N_21533,N_23361);
nand U28277 (N_28277,N_23021,N_18545);
nand U28278 (N_28278,N_22674,N_20977);
nor U28279 (N_28279,N_18881,N_23957);
nand U28280 (N_28280,N_20543,N_21497);
and U28281 (N_28281,N_21344,N_18479);
nor U28282 (N_28282,N_21764,N_18034);
or U28283 (N_28283,N_20502,N_19404);
and U28284 (N_28284,N_19678,N_19462);
nor U28285 (N_28285,N_19639,N_19720);
and U28286 (N_28286,N_23967,N_19038);
and U28287 (N_28287,N_21384,N_18181);
nor U28288 (N_28288,N_21564,N_20387);
nor U28289 (N_28289,N_23417,N_22407);
nand U28290 (N_28290,N_22321,N_19712);
nand U28291 (N_28291,N_22110,N_19715);
nor U28292 (N_28292,N_20599,N_18961);
nand U28293 (N_28293,N_19602,N_20517);
xnor U28294 (N_28294,N_20053,N_20355);
nand U28295 (N_28295,N_22586,N_22259);
and U28296 (N_28296,N_19577,N_22915);
xnor U28297 (N_28297,N_18436,N_18451);
and U28298 (N_28298,N_18381,N_23616);
and U28299 (N_28299,N_23221,N_23080);
and U28300 (N_28300,N_23824,N_22049);
and U28301 (N_28301,N_23526,N_21719);
xnor U28302 (N_28302,N_18969,N_20060);
or U28303 (N_28303,N_22097,N_20822);
nand U28304 (N_28304,N_18409,N_23281);
or U28305 (N_28305,N_23720,N_19926);
nand U28306 (N_28306,N_22446,N_20842);
nor U28307 (N_28307,N_22782,N_22254);
and U28308 (N_28308,N_21092,N_22505);
or U28309 (N_28309,N_23187,N_20233);
nor U28310 (N_28310,N_18180,N_21925);
nor U28311 (N_28311,N_22707,N_20209);
nand U28312 (N_28312,N_19268,N_21407);
nand U28313 (N_28313,N_18577,N_23465);
and U28314 (N_28314,N_18946,N_23555);
nor U28315 (N_28315,N_20983,N_21583);
nand U28316 (N_28316,N_19056,N_21101);
or U28317 (N_28317,N_23657,N_18973);
or U28318 (N_28318,N_23784,N_22066);
or U28319 (N_28319,N_21376,N_22079);
or U28320 (N_28320,N_22406,N_19800);
nand U28321 (N_28321,N_18461,N_19597);
and U28322 (N_28322,N_21883,N_21627);
nor U28323 (N_28323,N_22840,N_19581);
and U28324 (N_28324,N_18074,N_18587);
or U28325 (N_28325,N_19522,N_23266);
nand U28326 (N_28326,N_22915,N_22225);
or U28327 (N_28327,N_20790,N_18871);
or U28328 (N_28328,N_22926,N_21703);
nand U28329 (N_28329,N_20784,N_20014);
and U28330 (N_28330,N_21244,N_21628);
xor U28331 (N_28331,N_21820,N_21644);
or U28332 (N_28332,N_22772,N_18895);
nand U28333 (N_28333,N_23576,N_22121);
nor U28334 (N_28334,N_18218,N_18151);
or U28335 (N_28335,N_22951,N_20012);
and U28336 (N_28336,N_23978,N_19280);
nand U28337 (N_28337,N_22734,N_20050);
nor U28338 (N_28338,N_22473,N_22025);
or U28339 (N_28339,N_22263,N_20414);
nor U28340 (N_28340,N_20122,N_23269);
or U28341 (N_28341,N_20055,N_19309);
and U28342 (N_28342,N_19964,N_23645);
or U28343 (N_28343,N_20638,N_21665);
and U28344 (N_28344,N_20370,N_22182);
and U28345 (N_28345,N_23179,N_18980);
or U28346 (N_28346,N_18246,N_21405);
or U28347 (N_28347,N_18910,N_22422);
nor U28348 (N_28348,N_19943,N_20211);
nor U28349 (N_28349,N_22558,N_19067);
nor U28350 (N_28350,N_19887,N_21938);
and U28351 (N_28351,N_21251,N_22900);
xor U28352 (N_28352,N_23564,N_20815);
nand U28353 (N_28353,N_19198,N_18643);
nand U28354 (N_28354,N_19199,N_18412);
nand U28355 (N_28355,N_21817,N_20822);
nor U28356 (N_28356,N_18528,N_19342);
and U28357 (N_28357,N_18932,N_20004);
nand U28358 (N_28358,N_19540,N_19012);
and U28359 (N_28359,N_23585,N_19527);
and U28360 (N_28360,N_21986,N_20264);
or U28361 (N_28361,N_23027,N_19565);
or U28362 (N_28362,N_21159,N_22777);
or U28363 (N_28363,N_19825,N_21068);
and U28364 (N_28364,N_21278,N_20031);
or U28365 (N_28365,N_20842,N_22888);
nand U28366 (N_28366,N_22170,N_22555);
and U28367 (N_28367,N_20623,N_18255);
or U28368 (N_28368,N_22171,N_18872);
and U28369 (N_28369,N_22384,N_21807);
and U28370 (N_28370,N_21176,N_19534);
nor U28371 (N_28371,N_21747,N_21738);
nand U28372 (N_28372,N_19851,N_20955);
xor U28373 (N_28373,N_22625,N_22304);
nor U28374 (N_28374,N_20354,N_20764);
xnor U28375 (N_28375,N_18327,N_19209);
xor U28376 (N_28376,N_18148,N_18707);
nor U28377 (N_28377,N_23460,N_22154);
nor U28378 (N_28378,N_21139,N_22705);
xnor U28379 (N_28379,N_21423,N_21967);
or U28380 (N_28380,N_20203,N_18348);
nor U28381 (N_28381,N_19828,N_23540);
nor U28382 (N_28382,N_20540,N_23382);
or U28383 (N_28383,N_21204,N_22287);
xnor U28384 (N_28384,N_23151,N_21589);
and U28385 (N_28385,N_20766,N_20539);
nand U28386 (N_28386,N_21236,N_22523);
nor U28387 (N_28387,N_20153,N_19139);
nor U28388 (N_28388,N_20755,N_21103);
nor U28389 (N_28389,N_23270,N_21633);
xnor U28390 (N_28390,N_18032,N_23195);
nor U28391 (N_28391,N_21729,N_22504);
nand U28392 (N_28392,N_20750,N_18823);
nand U28393 (N_28393,N_23652,N_22361);
nor U28394 (N_28394,N_21217,N_18301);
or U28395 (N_28395,N_21211,N_20506);
or U28396 (N_28396,N_22946,N_21799);
and U28397 (N_28397,N_18075,N_21017);
or U28398 (N_28398,N_19230,N_18107);
and U28399 (N_28399,N_22806,N_20964);
nor U28400 (N_28400,N_21587,N_18593);
nand U28401 (N_28401,N_21680,N_21619);
and U28402 (N_28402,N_21841,N_18400);
nor U28403 (N_28403,N_23696,N_20258);
nor U28404 (N_28404,N_23112,N_23083);
and U28405 (N_28405,N_20571,N_20666);
and U28406 (N_28406,N_20414,N_20087);
nor U28407 (N_28407,N_19006,N_18837);
and U28408 (N_28408,N_18320,N_20879);
nand U28409 (N_28409,N_23123,N_18057);
nand U28410 (N_28410,N_21873,N_20602);
nand U28411 (N_28411,N_22495,N_23407);
xor U28412 (N_28412,N_21490,N_20609);
xnor U28413 (N_28413,N_21469,N_18656);
nor U28414 (N_28414,N_19738,N_21943);
nor U28415 (N_28415,N_22951,N_20623);
or U28416 (N_28416,N_22113,N_23387);
or U28417 (N_28417,N_20246,N_23600);
nand U28418 (N_28418,N_23032,N_19524);
and U28419 (N_28419,N_20532,N_23550);
xnor U28420 (N_28420,N_20408,N_18353);
nand U28421 (N_28421,N_23530,N_18182);
nor U28422 (N_28422,N_23829,N_22981);
and U28423 (N_28423,N_20276,N_19428);
or U28424 (N_28424,N_23410,N_23460);
and U28425 (N_28425,N_20139,N_21023);
nor U28426 (N_28426,N_19418,N_23863);
nand U28427 (N_28427,N_23121,N_21861);
and U28428 (N_28428,N_18897,N_23131);
nand U28429 (N_28429,N_21865,N_18278);
or U28430 (N_28430,N_22884,N_20132);
nand U28431 (N_28431,N_22922,N_20802);
and U28432 (N_28432,N_22865,N_19904);
xor U28433 (N_28433,N_22535,N_18546);
and U28434 (N_28434,N_19210,N_23591);
and U28435 (N_28435,N_20523,N_21255);
nand U28436 (N_28436,N_23518,N_23305);
xor U28437 (N_28437,N_19204,N_20655);
and U28438 (N_28438,N_18545,N_23452);
xor U28439 (N_28439,N_19813,N_19589);
or U28440 (N_28440,N_22512,N_21229);
or U28441 (N_28441,N_23906,N_23346);
nand U28442 (N_28442,N_22499,N_22517);
or U28443 (N_28443,N_22005,N_22615);
or U28444 (N_28444,N_22559,N_20314);
and U28445 (N_28445,N_18766,N_21706);
nor U28446 (N_28446,N_19173,N_23994);
nand U28447 (N_28447,N_20772,N_18601);
nor U28448 (N_28448,N_22437,N_20619);
nand U28449 (N_28449,N_21984,N_23761);
nand U28450 (N_28450,N_22379,N_23610);
or U28451 (N_28451,N_23385,N_19807);
nor U28452 (N_28452,N_21044,N_23324);
and U28453 (N_28453,N_18855,N_22108);
nor U28454 (N_28454,N_19624,N_20906);
and U28455 (N_28455,N_20230,N_18514);
or U28456 (N_28456,N_22532,N_18680);
and U28457 (N_28457,N_22053,N_21173);
nand U28458 (N_28458,N_20723,N_19740);
xor U28459 (N_28459,N_19475,N_23942);
nand U28460 (N_28460,N_19004,N_19729);
or U28461 (N_28461,N_18991,N_22628);
xnor U28462 (N_28462,N_20347,N_20353);
nand U28463 (N_28463,N_23275,N_21950);
nand U28464 (N_28464,N_22676,N_23688);
nor U28465 (N_28465,N_23468,N_19419);
nand U28466 (N_28466,N_23184,N_21024);
nor U28467 (N_28467,N_21308,N_23868);
or U28468 (N_28468,N_23806,N_23432);
or U28469 (N_28469,N_18718,N_19388);
nor U28470 (N_28470,N_20736,N_23007);
nand U28471 (N_28471,N_18844,N_19940);
or U28472 (N_28472,N_23517,N_22945);
or U28473 (N_28473,N_19934,N_19153);
nor U28474 (N_28474,N_23754,N_21512);
or U28475 (N_28475,N_18832,N_23086);
xnor U28476 (N_28476,N_20095,N_22802);
and U28477 (N_28477,N_18765,N_23971);
xnor U28478 (N_28478,N_18360,N_18067);
or U28479 (N_28479,N_22269,N_18286);
nand U28480 (N_28480,N_20575,N_19323);
and U28481 (N_28481,N_22089,N_18573);
xnor U28482 (N_28482,N_23667,N_20181);
or U28483 (N_28483,N_19316,N_20166);
nor U28484 (N_28484,N_19326,N_20149);
and U28485 (N_28485,N_23968,N_22473);
nor U28486 (N_28486,N_21375,N_21181);
and U28487 (N_28487,N_18649,N_23548);
nand U28488 (N_28488,N_21494,N_19544);
nand U28489 (N_28489,N_20153,N_22970);
nor U28490 (N_28490,N_19253,N_23330);
and U28491 (N_28491,N_22385,N_19022);
xor U28492 (N_28492,N_19449,N_22593);
nor U28493 (N_28493,N_20978,N_22840);
nor U28494 (N_28494,N_19152,N_23581);
nand U28495 (N_28495,N_21849,N_23089);
xnor U28496 (N_28496,N_22519,N_20535);
nor U28497 (N_28497,N_20941,N_22226);
xnor U28498 (N_28498,N_18975,N_19286);
nor U28499 (N_28499,N_22610,N_19040);
and U28500 (N_28500,N_21281,N_20865);
nor U28501 (N_28501,N_19232,N_20256);
and U28502 (N_28502,N_23346,N_19585);
xor U28503 (N_28503,N_19248,N_23294);
nor U28504 (N_28504,N_19742,N_22351);
or U28505 (N_28505,N_22227,N_23135);
or U28506 (N_28506,N_22474,N_21834);
nand U28507 (N_28507,N_22481,N_20954);
and U28508 (N_28508,N_22680,N_19211);
and U28509 (N_28509,N_21707,N_20478);
xor U28510 (N_28510,N_20084,N_21756);
nor U28511 (N_28511,N_18640,N_20361);
nand U28512 (N_28512,N_20057,N_21021);
nor U28513 (N_28513,N_23953,N_18548);
nor U28514 (N_28514,N_19226,N_21695);
or U28515 (N_28515,N_18995,N_22614);
nor U28516 (N_28516,N_19231,N_22933);
and U28517 (N_28517,N_22785,N_19005);
nand U28518 (N_28518,N_18210,N_19077);
nand U28519 (N_28519,N_19314,N_19274);
nor U28520 (N_28520,N_20305,N_20372);
or U28521 (N_28521,N_22173,N_23048);
nand U28522 (N_28522,N_18719,N_22417);
and U28523 (N_28523,N_21025,N_18491);
or U28524 (N_28524,N_22921,N_21209);
nand U28525 (N_28525,N_19364,N_22619);
nor U28526 (N_28526,N_18571,N_21494);
or U28527 (N_28527,N_18370,N_23874);
nand U28528 (N_28528,N_20898,N_23122);
nor U28529 (N_28529,N_18245,N_20731);
and U28530 (N_28530,N_20691,N_23798);
or U28531 (N_28531,N_21536,N_18348);
nor U28532 (N_28532,N_20364,N_20860);
nand U28533 (N_28533,N_19084,N_21437);
nor U28534 (N_28534,N_23212,N_22729);
xor U28535 (N_28535,N_23412,N_22878);
nand U28536 (N_28536,N_23997,N_23431);
or U28537 (N_28537,N_21300,N_20300);
or U28538 (N_28538,N_19242,N_19751);
or U28539 (N_28539,N_22219,N_19555);
nand U28540 (N_28540,N_23128,N_22545);
nor U28541 (N_28541,N_19721,N_19844);
and U28542 (N_28542,N_19375,N_20242);
or U28543 (N_28543,N_20997,N_21349);
nand U28544 (N_28544,N_19428,N_20629);
nand U28545 (N_28545,N_18683,N_23853);
or U28546 (N_28546,N_18828,N_22397);
nor U28547 (N_28547,N_23347,N_19223);
nor U28548 (N_28548,N_21106,N_20706);
nand U28549 (N_28549,N_18810,N_18402);
nor U28550 (N_28550,N_20905,N_23072);
or U28551 (N_28551,N_22371,N_20700);
or U28552 (N_28552,N_18642,N_19856);
nor U28553 (N_28553,N_19197,N_18306);
nor U28554 (N_28554,N_18368,N_23381);
and U28555 (N_28555,N_18294,N_23882);
or U28556 (N_28556,N_23926,N_20875);
nor U28557 (N_28557,N_20268,N_23824);
and U28558 (N_28558,N_20233,N_18292);
or U28559 (N_28559,N_18414,N_22064);
nor U28560 (N_28560,N_22314,N_18148);
or U28561 (N_28561,N_18316,N_18380);
and U28562 (N_28562,N_22916,N_18150);
nor U28563 (N_28563,N_21613,N_18056);
nand U28564 (N_28564,N_19977,N_20637);
nand U28565 (N_28565,N_18032,N_23752);
or U28566 (N_28566,N_19678,N_21058);
nor U28567 (N_28567,N_23825,N_20573);
and U28568 (N_28568,N_20964,N_19329);
or U28569 (N_28569,N_23625,N_21214);
and U28570 (N_28570,N_18081,N_19426);
nand U28571 (N_28571,N_23022,N_23147);
nand U28572 (N_28572,N_23847,N_19976);
or U28573 (N_28573,N_21202,N_18856);
nand U28574 (N_28574,N_19794,N_19861);
nor U28575 (N_28575,N_20089,N_20610);
nand U28576 (N_28576,N_20395,N_18513);
or U28577 (N_28577,N_21791,N_22814);
and U28578 (N_28578,N_19510,N_21215);
nor U28579 (N_28579,N_22219,N_19993);
or U28580 (N_28580,N_21146,N_20217);
nor U28581 (N_28581,N_18438,N_20449);
and U28582 (N_28582,N_19148,N_22436);
nand U28583 (N_28583,N_19649,N_20198);
nor U28584 (N_28584,N_22972,N_20843);
nor U28585 (N_28585,N_19106,N_23561);
nor U28586 (N_28586,N_19527,N_23675);
or U28587 (N_28587,N_22063,N_23631);
or U28588 (N_28588,N_19397,N_21707);
and U28589 (N_28589,N_19572,N_23886);
xnor U28590 (N_28590,N_18192,N_23764);
nand U28591 (N_28591,N_19299,N_18238);
nor U28592 (N_28592,N_21334,N_20469);
nor U28593 (N_28593,N_22786,N_18188);
nand U28594 (N_28594,N_21399,N_20183);
nand U28595 (N_28595,N_22324,N_19794);
nor U28596 (N_28596,N_20171,N_22867);
xor U28597 (N_28597,N_23549,N_21660);
xnor U28598 (N_28598,N_23935,N_21078);
nor U28599 (N_28599,N_19151,N_20944);
xnor U28600 (N_28600,N_21995,N_21174);
nor U28601 (N_28601,N_18586,N_22175);
nor U28602 (N_28602,N_19216,N_18855);
nand U28603 (N_28603,N_19447,N_18602);
nor U28604 (N_28604,N_22931,N_20704);
nand U28605 (N_28605,N_20656,N_22896);
nand U28606 (N_28606,N_21435,N_19839);
nor U28607 (N_28607,N_18396,N_22795);
and U28608 (N_28608,N_21257,N_23087);
or U28609 (N_28609,N_18288,N_21970);
nor U28610 (N_28610,N_22880,N_21909);
nor U28611 (N_28611,N_20534,N_21225);
nor U28612 (N_28612,N_19259,N_18771);
nor U28613 (N_28613,N_20642,N_18364);
or U28614 (N_28614,N_18632,N_22892);
nand U28615 (N_28615,N_20135,N_20614);
nand U28616 (N_28616,N_20000,N_18581);
and U28617 (N_28617,N_23940,N_18016);
or U28618 (N_28618,N_20672,N_23666);
and U28619 (N_28619,N_18398,N_18001);
nor U28620 (N_28620,N_18502,N_22048);
and U28621 (N_28621,N_19961,N_22534);
nand U28622 (N_28622,N_21316,N_21956);
and U28623 (N_28623,N_18733,N_22622);
and U28624 (N_28624,N_23443,N_21664);
xnor U28625 (N_28625,N_23310,N_23487);
nand U28626 (N_28626,N_23960,N_18533);
and U28627 (N_28627,N_21027,N_18189);
nor U28628 (N_28628,N_20212,N_22119);
nand U28629 (N_28629,N_19799,N_22218);
nor U28630 (N_28630,N_18705,N_21365);
nand U28631 (N_28631,N_19827,N_22029);
nand U28632 (N_28632,N_23832,N_19801);
nor U28633 (N_28633,N_23867,N_18876);
nand U28634 (N_28634,N_20168,N_19833);
or U28635 (N_28635,N_19499,N_23647);
nor U28636 (N_28636,N_19505,N_23345);
nor U28637 (N_28637,N_21091,N_23071);
and U28638 (N_28638,N_20201,N_23286);
or U28639 (N_28639,N_20347,N_22078);
xnor U28640 (N_28640,N_20587,N_20361);
nand U28641 (N_28641,N_20594,N_21534);
xor U28642 (N_28642,N_21586,N_23513);
and U28643 (N_28643,N_18181,N_20144);
nor U28644 (N_28644,N_20170,N_19484);
nand U28645 (N_28645,N_21275,N_19827);
or U28646 (N_28646,N_23691,N_19551);
nand U28647 (N_28647,N_19464,N_21608);
or U28648 (N_28648,N_21977,N_23699);
or U28649 (N_28649,N_20288,N_20504);
nor U28650 (N_28650,N_23581,N_18366);
xor U28651 (N_28651,N_21210,N_22782);
nor U28652 (N_28652,N_20821,N_22309);
nor U28653 (N_28653,N_22032,N_19743);
nor U28654 (N_28654,N_20986,N_18915);
xor U28655 (N_28655,N_21684,N_20543);
nand U28656 (N_28656,N_19713,N_20881);
and U28657 (N_28657,N_22492,N_23647);
nor U28658 (N_28658,N_22769,N_23579);
and U28659 (N_28659,N_22038,N_21232);
and U28660 (N_28660,N_20145,N_19946);
nand U28661 (N_28661,N_19242,N_20612);
xnor U28662 (N_28662,N_22231,N_22545);
and U28663 (N_28663,N_19574,N_18358);
or U28664 (N_28664,N_22591,N_19789);
nor U28665 (N_28665,N_21741,N_19446);
nand U28666 (N_28666,N_22807,N_23240);
xor U28667 (N_28667,N_21118,N_22821);
nand U28668 (N_28668,N_21702,N_19702);
and U28669 (N_28669,N_20099,N_20167);
nor U28670 (N_28670,N_19573,N_20125);
nor U28671 (N_28671,N_23991,N_22695);
nor U28672 (N_28672,N_19640,N_22966);
or U28673 (N_28673,N_22705,N_22564);
nand U28674 (N_28674,N_22450,N_19320);
nand U28675 (N_28675,N_20009,N_19323);
and U28676 (N_28676,N_19332,N_20782);
or U28677 (N_28677,N_20570,N_19333);
and U28678 (N_28678,N_20589,N_23882);
nor U28679 (N_28679,N_18816,N_20266);
or U28680 (N_28680,N_21903,N_23395);
and U28681 (N_28681,N_22166,N_19280);
nor U28682 (N_28682,N_18103,N_22030);
nand U28683 (N_28683,N_23511,N_18985);
or U28684 (N_28684,N_21102,N_19307);
and U28685 (N_28685,N_18664,N_22198);
and U28686 (N_28686,N_19828,N_18259);
and U28687 (N_28687,N_22348,N_21097);
nor U28688 (N_28688,N_19996,N_22263);
nor U28689 (N_28689,N_18765,N_23642);
or U28690 (N_28690,N_18696,N_19083);
or U28691 (N_28691,N_21496,N_21981);
xor U28692 (N_28692,N_22733,N_23321);
and U28693 (N_28693,N_22494,N_21649);
nor U28694 (N_28694,N_20023,N_19340);
or U28695 (N_28695,N_23535,N_21422);
or U28696 (N_28696,N_23180,N_18134);
nor U28697 (N_28697,N_19425,N_22737);
nand U28698 (N_28698,N_23082,N_18605);
and U28699 (N_28699,N_18797,N_20191);
nor U28700 (N_28700,N_19734,N_23564);
nand U28701 (N_28701,N_20163,N_20012);
or U28702 (N_28702,N_19036,N_20015);
nand U28703 (N_28703,N_19889,N_18839);
nand U28704 (N_28704,N_18233,N_19309);
and U28705 (N_28705,N_18112,N_19572);
nand U28706 (N_28706,N_20771,N_21942);
nand U28707 (N_28707,N_18564,N_22328);
and U28708 (N_28708,N_20654,N_20083);
and U28709 (N_28709,N_20972,N_21387);
xnor U28710 (N_28710,N_19400,N_23816);
xnor U28711 (N_28711,N_18931,N_21898);
nand U28712 (N_28712,N_19099,N_21929);
xnor U28713 (N_28713,N_19278,N_18246);
and U28714 (N_28714,N_18258,N_23402);
xor U28715 (N_28715,N_20038,N_18829);
and U28716 (N_28716,N_18599,N_23798);
nand U28717 (N_28717,N_22435,N_23197);
or U28718 (N_28718,N_18061,N_20693);
nand U28719 (N_28719,N_19211,N_20883);
or U28720 (N_28720,N_23028,N_22844);
and U28721 (N_28721,N_23920,N_19385);
nand U28722 (N_28722,N_19180,N_21623);
or U28723 (N_28723,N_21948,N_19561);
nor U28724 (N_28724,N_20518,N_20578);
nand U28725 (N_28725,N_20443,N_21502);
or U28726 (N_28726,N_19755,N_21741);
or U28727 (N_28727,N_18109,N_22881);
and U28728 (N_28728,N_18971,N_22221);
xor U28729 (N_28729,N_19225,N_19697);
or U28730 (N_28730,N_21606,N_23517);
nor U28731 (N_28731,N_21519,N_23919);
or U28732 (N_28732,N_20264,N_22830);
and U28733 (N_28733,N_21366,N_23586);
or U28734 (N_28734,N_19231,N_23942);
nor U28735 (N_28735,N_18004,N_22804);
and U28736 (N_28736,N_23715,N_18540);
nand U28737 (N_28737,N_22625,N_20215);
nor U28738 (N_28738,N_23805,N_20037);
or U28739 (N_28739,N_22135,N_20743);
or U28740 (N_28740,N_20204,N_22467);
or U28741 (N_28741,N_23059,N_21764);
and U28742 (N_28742,N_20416,N_22418);
nor U28743 (N_28743,N_21780,N_18032);
xor U28744 (N_28744,N_19865,N_19292);
and U28745 (N_28745,N_21048,N_20712);
nand U28746 (N_28746,N_19471,N_23787);
nor U28747 (N_28747,N_21560,N_19574);
and U28748 (N_28748,N_18645,N_23144);
and U28749 (N_28749,N_23016,N_20802);
nand U28750 (N_28750,N_18789,N_20504);
nand U28751 (N_28751,N_23270,N_22405);
nor U28752 (N_28752,N_22218,N_21846);
nor U28753 (N_28753,N_18717,N_22368);
or U28754 (N_28754,N_23347,N_22403);
nor U28755 (N_28755,N_18927,N_18651);
or U28756 (N_28756,N_18912,N_22944);
and U28757 (N_28757,N_22572,N_22329);
nand U28758 (N_28758,N_18208,N_19337);
nand U28759 (N_28759,N_21835,N_21365);
or U28760 (N_28760,N_19585,N_20799);
and U28761 (N_28761,N_19215,N_21089);
nand U28762 (N_28762,N_21252,N_20252);
nand U28763 (N_28763,N_18091,N_22535);
nor U28764 (N_28764,N_21135,N_23999);
or U28765 (N_28765,N_19497,N_20450);
nand U28766 (N_28766,N_19218,N_19465);
and U28767 (N_28767,N_21512,N_18600);
and U28768 (N_28768,N_23095,N_22857);
nand U28769 (N_28769,N_22674,N_21936);
and U28770 (N_28770,N_21949,N_23298);
or U28771 (N_28771,N_23525,N_23435);
nor U28772 (N_28772,N_18510,N_22645);
nor U28773 (N_28773,N_23877,N_22981);
nor U28774 (N_28774,N_23910,N_19110);
nand U28775 (N_28775,N_23450,N_19948);
xnor U28776 (N_28776,N_19356,N_19368);
or U28777 (N_28777,N_18199,N_21351);
nand U28778 (N_28778,N_20763,N_21558);
or U28779 (N_28779,N_18281,N_19996);
or U28780 (N_28780,N_21084,N_22223);
and U28781 (N_28781,N_20328,N_22339);
and U28782 (N_28782,N_23242,N_22918);
xnor U28783 (N_28783,N_23057,N_22270);
xnor U28784 (N_28784,N_19616,N_22878);
or U28785 (N_28785,N_21919,N_18892);
nor U28786 (N_28786,N_21254,N_23882);
nand U28787 (N_28787,N_19765,N_20052);
and U28788 (N_28788,N_19873,N_21447);
nor U28789 (N_28789,N_19545,N_22562);
nand U28790 (N_28790,N_22917,N_18355);
and U28791 (N_28791,N_19929,N_18805);
or U28792 (N_28792,N_22447,N_18065);
nand U28793 (N_28793,N_18421,N_20549);
and U28794 (N_28794,N_18833,N_20069);
and U28795 (N_28795,N_22552,N_19988);
or U28796 (N_28796,N_18306,N_19125);
and U28797 (N_28797,N_20713,N_21565);
or U28798 (N_28798,N_21341,N_18877);
nand U28799 (N_28799,N_19005,N_18279);
or U28800 (N_28800,N_22493,N_22153);
and U28801 (N_28801,N_21032,N_22140);
nor U28802 (N_28802,N_18322,N_20977);
or U28803 (N_28803,N_20446,N_19540);
nand U28804 (N_28804,N_18942,N_20639);
nand U28805 (N_28805,N_22038,N_18054);
and U28806 (N_28806,N_21543,N_20199);
or U28807 (N_28807,N_21632,N_21766);
nor U28808 (N_28808,N_20843,N_18330);
nand U28809 (N_28809,N_23546,N_21141);
or U28810 (N_28810,N_20746,N_18926);
and U28811 (N_28811,N_22154,N_20270);
or U28812 (N_28812,N_23055,N_19837);
nand U28813 (N_28813,N_21319,N_18039);
nand U28814 (N_28814,N_21274,N_23468);
nand U28815 (N_28815,N_19435,N_19565);
nor U28816 (N_28816,N_21071,N_19881);
nor U28817 (N_28817,N_20447,N_19188);
and U28818 (N_28818,N_20858,N_23813);
nand U28819 (N_28819,N_18573,N_21987);
xnor U28820 (N_28820,N_19139,N_22866);
nand U28821 (N_28821,N_21958,N_23837);
nor U28822 (N_28822,N_19556,N_19713);
nor U28823 (N_28823,N_23110,N_23334);
nand U28824 (N_28824,N_21316,N_20204);
and U28825 (N_28825,N_19028,N_21350);
xnor U28826 (N_28826,N_22873,N_23473);
or U28827 (N_28827,N_21552,N_23569);
nand U28828 (N_28828,N_20577,N_19967);
nand U28829 (N_28829,N_19436,N_21945);
nor U28830 (N_28830,N_22226,N_23245);
or U28831 (N_28831,N_19332,N_20203);
nor U28832 (N_28832,N_23030,N_21815);
nor U28833 (N_28833,N_19703,N_19076);
and U28834 (N_28834,N_18639,N_19738);
nand U28835 (N_28835,N_18998,N_23934);
and U28836 (N_28836,N_22824,N_18851);
xnor U28837 (N_28837,N_21226,N_23542);
or U28838 (N_28838,N_19386,N_20315);
and U28839 (N_28839,N_23510,N_23134);
nand U28840 (N_28840,N_18863,N_23096);
or U28841 (N_28841,N_18877,N_22512);
or U28842 (N_28842,N_21130,N_23033);
nand U28843 (N_28843,N_18069,N_19103);
nor U28844 (N_28844,N_22827,N_19429);
nand U28845 (N_28845,N_22879,N_18195);
xnor U28846 (N_28846,N_21064,N_19493);
or U28847 (N_28847,N_23397,N_21150);
nand U28848 (N_28848,N_18161,N_18015);
nor U28849 (N_28849,N_23108,N_21189);
nor U28850 (N_28850,N_21266,N_23396);
xor U28851 (N_28851,N_23507,N_18456);
and U28852 (N_28852,N_21621,N_19865);
nand U28853 (N_28853,N_22269,N_18543);
xnor U28854 (N_28854,N_18574,N_19668);
and U28855 (N_28855,N_23134,N_21353);
nor U28856 (N_28856,N_19823,N_18678);
or U28857 (N_28857,N_18340,N_20204);
and U28858 (N_28858,N_18633,N_18192);
nand U28859 (N_28859,N_21888,N_20008);
or U28860 (N_28860,N_18048,N_19668);
and U28861 (N_28861,N_22387,N_23007);
and U28862 (N_28862,N_19334,N_21429);
nor U28863 (N_28863,N_21087,N_18690);
or U28864 (N_28864,N_21969,N_18248);
nand U28865 (N_28865,N_22007,N_21967);
nor U28866 (N_28866,N_23280,N_22984);
or U28867 (N_28867,N_22020,N_18025);
or U28868 (N_28868,N_19793,N_23825);
nand U28869 (N_28869,N_23094,N_22629);
nor U28870 (N_28870,N_19150,N_23833);
nand U28871 (N_28871,N_21261,N_21879);
and U28872 (N_28872,N_23766,N_19475);
and U28873 (N_28873,N_22078,N_22403);
or U28874 (N_28874,N_21785,N_21039);
or U28875 (N_28875,N_19802,N_20842);
and U28876 (N_28876,N_19044,N_23973);
nor U28877 (N_28877,N_19339,N_21137);
and U28878 (N_28878,N_18750,N_21472);
nor U28879 (N_28879,N_23734,N_18446);
and U28880 (N_28880,N_18330,N_19461);
nor U28881 (N_28881,N_20502,N_20116);
nor U28882 (N_28882,N_20225,N_18014);
nand U28883 (N_28883,N_23425,N_22499);
or U28884 (N_28884,N_19102,N_20934);
nor U28885 (N_28885,N_22906,N_19295);
and U28886 (N_28886,N_23364,N_19950);
nor U28887 (N_28887,N_18497,N_20838);
nand U28888 (N_28888,N_20581,N_22224);
nand U28889 (N_28889,N_19464,N_22895);
and U28890 (N_28890,N_23696,N_21515);
nor U28891 (N_28891,N_20934,N_18759);
and U28892 (N_28892,N_22217,N_20526);
and U28893 (N_28893,N_23393,N_22913);
nor U28894 (N_28894,N_22207,N_22746);
or U28895 (N_28895,N_19757,N_20104);
nand U28896 (N_28896,N_22047,N_18651);
nand U28897 (N_28897,N_19881,N_19953);
nor U28898 (N_28898,N_22489,N_23105);
nor U28899 (N_28899,N_22616,N_19645);
nor U28900 (N_28900,N_19742,N_18150);
nor U28901 (N_28901,N_21682,N_23371);
nor U28902 (N_28902,N_21879,N_19405);
nor U28903 (N_28903,N_22420,N_20714);
nand U28904 (N_28904,N_18849,N_23782);
xnor U28905 (N_28905,N_19985,N_20218);
nor U28906 (N_28906,N_23429,N_19352);
nand U28907 (N_28907,N_23113,N_23447);
nor U28908 (N_28908,N_23600,N_20407);
nand U28909 (N_28909,N_18238,N_21928);
or U28910 (N_28910,N_21603,N_19381);
or U28911 (N_28911,N_20547,N_21804);
and U28912 (N_28912,N_19152,N_18607);
or U28913 (N_28913,N_23079,N_19171);
and U28914 (N_28914,N_19343,N_21392);
or U28915 (N_28915,N_20985,N_21118);
or U28916 (N_28916,N_23059,N_22977);
and U28917 (N_28917,N_22900,N_23804);
nor U28918 (N_28918,N_21187,N_20452);
or U28919 (N_28919,N_23544,N_23653);
nor U28920 (N_28920,N_23873,N_19482);
nor U28921 (N_28921,N_20411,N_23341);
or U28922 (N_28922,N_18821,N_22370);
nor U28923 (N_28923,N_20890,N_19560);
and U28924 (N_28924,N_18921,N_19284);
xor U28925 (N_28925,N_19121,N_18678);
or U28926 (N_28926,N_20694,N_20466);
nor U28927 (N_28927,N_19747,N_20345);
nor U28928 (N_28928,N_21814,N_22778);
nand U28929 (N_28929,N_19414,N_19581);
or U28930 (N_28930,N_19339,N_18683);
nor U28931 (N_28931,N_18766,N_20527);
xor U28932 (N_28932,N_18173,N_20649);
or U28933 (N_28933,N_20484,N_18234);
nand U28934 (N_28934,N_18234,N_19976);
and U28935 (N_28935,N_22199,N_22011);
and U28936 (N_28936,N_18048,N_22054);
nand U28937 (N_28937,N_22417,N_18897);
nor U28938 (N_28938,N_23239,N_22182);
and U28939 (N_28939,N_21204,N_22181);
and U28940 (N_28940,N_21613,N_22485);
and U28941 (N_28941,N_20421,N_18030);
nand U28942 (N_28942,N_18128,N_19339);
nor U28943 (N_28943,N_18639,N_19399);
nand U28944 (N_28944,N_23942,N_23452);
nor U28945 (N_28945,N_21536,N_19049);
nor U28946 (N_28946,N_20034,N_22316);
nand U28947 (N_28947,N_21401,N_20854);
nor U28948 (N_28948,N_19532,N_22116);
or U28949 (N_28949,N_23002,N_21889);
and U28950 (N_28950,N_23904,N_23359);
nor U28951 (N_28951,N_21273,N_19145);
nor U28952 (N_28952,N_20570,N_18886);
nor U28953 (N_28953,N_19763,N_22866);
and U28954 (N_28954,N_23269,N_18804);
nand U28955 (N_28955,N_22254,N_20234);
and U28956 (N_28956,N_19991,N_23310);
nor U28957 (N_28957,N_23829,N_22451);
and U28958 (N_28958,N_21066,N_18475);
or U28959 (N_28959,N_18652,N_21887);
nor U28960 (N_28960,N_18334,N_19151);
nand U28961 (N_28961,N_20497,N_23578);
nor U28962 (N_28962,N_18870,N_18149);
nand U28963 (N_28963,N_18179,N_19068);
and U28964 (N_28964,N_23468,N_22379);
xnor U28965 (N_28965,N_19366,N_19225);
nand U28966 (N_28966,N_21232,N_20158);
and U28967 (N_28967,N_23932,N_21642);
nor U28968 (N_28968,N_18064,N_18726);
nand U28969 (N_28969,N_18193,N_23690);
nor U28970 (N_28970,N_21358,N_19004);
or U28971 (N_28971,N_20802,N_20959);
nand U28972 (N_28972,N_21144,N_19284);
and U28973 (N_28973,N_18948,N_20029);
xor U28974 (N_28974,N_21244,N_19600);
and U28975 (N_28975,N_21297,N_20779);
nand U28976 (N_28976,N_19392,N_20118);
and U28977 (N_28977,N_23962,N_22492);
xnor U28978 (N_28978,N_18173,N_19137);
nor U28979 (N_28979,N_19264,N_21928);
nor U28980 (N_28980,N_22815,N_21976);
nand U28981 (N_28981,N_20543,N_20345);
nand U28982 (N_28982,N_18073,N_21278);
and U28983 (N_28983,N_20314,N_20154);
or U28984 (N_28984,N_20923,N_18445);
or U28985 (N_28985,N_23393,N_19040);
nand U28986 (N_28986,N_23180,N_23606);
nand U28987 (N_28987,N_19755,N_18759);
nand U28988 (N_28988,N_20693,N_19910);
and U28989 (N_28989,N_19355,N_21772);
nor U28990 (N_28990,N_22962,N_21024);
nand U28991 (N_28991,N_21334,N_18595);
nor U28992 (N_28992,N_21166,N_22339);
nand U28993 (N_28993,N_20145,N_18306);
nor U28994 (N_28994,N_18255,N_23796);
nand U28995 (N_28995,N_21068,N_19839);
nor U28996 (N_28996,N_20789,N_19246);
and U28997 (N_28997,N_21755,N_18433);
or U28998 (N_28998,N_20132,N_22404);
xnor U28999 (N_28999,N_20102,N_18276);
nor U29000 (N_29000,N_18449,N_18050);
nand U29001 (N_29001,N_20209,N_23685);
nor U29002 (N_29002,N_21162,N_19323);
nor U29003 (N_29003,N_18385,N_22728);
nor U29004 (N_29004,N_22969,N_20712);
nor U29005 (N_29005,N_19397,N_23061);
xor U29006 (N_29006,N_22830,N_20584);
or U29007 (N_29007,N_23690,N_20734);
nor U29008 (N_29008,N_20463,N_21369);
nor U29009 (N_29009,N_19171,N_22959);
and U29010 (N_29010,N_23058,N_19435);
nand U29011 (N_29011,N_22306,N_18299);
or U29012 (N_29012,N_21754,N_22555);
nor U29013 (N_29013,N_19372,N_22029);
or U29014 (N_29014,N_21965,N_18652);
and U29015 (N_29015,N_23395,N_20015);
nor U29016 (N_29016,N_23410,N_23164);
or U29017 (N_29017,N_22560,N_22486);
and U29018 (N_29018,N_19925,N_18199);
or U29019 (N_29019,N_20160,N_20630);
or U29020 (N_29020,N_22343,N_18185);
nand U29021 (N_29021,N_18982,N_23344);
or U29022 (N_29022,N_19863,N_18216);
nand U29023 (N_29023,N_19166,N_21592);
and U29024 (N_29024,N_23701,N_22421);
and U29025 (N_29025,N_20364,N_18777);
and U29026 (N_29026,N_18478,N_23193);
nor U29027 (N_29027,N_21530,N_18891);
xor U29028 (N_29028,N_23595,N_22164);
nor U29029 (N_29029,N_22238,N_19984);
and U29030 (N_29030,N_23784,N_19082);
nor U29031 (N_29031,N_21943,N_22227);
or U29032 (N_29032,N_20960,N_20163);
or U29033 (N_29033,N_23274,N_18131);
or U29034 (N_29034,N_18706,N_18936);
nor U29035 (N_29035,N_21879,N_22031);
and U29036 (N_29036,N_23407,N_21376);
or U29037 (N_29037,N_22273,N_23651);
xor U29038 (N_29038,N_19172,N_19431);
nand U29039 (N_29039,N_23470,N_19325);
or U29040 (N_29040,N_22959,N_21961);
nor U29041 (N_29041,N_23373,N_20348);
nor U29042 (N_29042,N_18929,N_22350);
and U29043 (N_29043,N_21852,N_18457);
and U29044 (N_29044,N_23982,N_21724);
xor U29045 (N_29045,N_18113,N_18320);
nand U29046 (N_29046,N_20080,N_21304);
or U29047 (N_29047,N_18488,N_20140);
nor U29048 (N_29048,N_20465,N_21458);
nor U29049 (N_29049,N_21972,N_19947);
or U29050 (N_29050,N_20219,N_18574);
nor U29051 (N_29051,N_20236,N_20023);
xor U29052 (N_29052,N_22532,N_18129);
nand U29053 (N_29053,N_18328,N_23456);
nand U29054 (N_29054,N_20309,N_20937);
and U29055 (N_29055,N_20170,N_23744);
nor U29056 (N_29056,N_20332,N_21987);
and U29057 (N_29057,N_23116,N_20142);
xor U29058 (N_29058,N_22053,N_22998);
or U29059 (N_29059,N_21332,N_20830);
nand U29060 (N_29060,N_22670,N_22081);
nand U29061 (N_29061,N_21874,N_19028);
nor U29062 (N_29062,N_21470,N_22601);
nor U29063 (N_29063,N_19174,N_20014);
nor U29064 (N_29064,N_23368,N_21834);
or U29065 (N_29065,N_22135,N_21332);
nor U29066 (N_29066,N_23412,N_20622);
and U29067 (N_29067,N_18598,N_23370);
xor U29068 (N_29068,N_22958,N_21221);
nand U29069 (N_29069,N_18940,N_20124);
nand U29070 (N_29070,N_23801,N_21208);
and U29071 (N_29071,N_20003,N_22756);
or U29072 (N_29072,N_23773,N_20221);
nor U29073 (N_29073,N_20176,N_19804);
or U29074 (N_29074,N_18359,N_22271);
nand U29075 (N_29075,N_19951,N_20710);
xor U29076 (N_29076,N_22546,N_20659);
and U29077 (N_29077,N_20579,N_19078);
nor U29078 (N_29078,N_19645,N_20619);
nand U29079 (N_29079,N_20624,N_21051);
nor U29080 (N_29080,N_21701,N_18537);
nor U29081 (N_29081,N_19021,N_22631);
and U29082 (N_29082,N_21157,N_22629);
or U29083 (N_29083,N_19596,N_22497);
nor U29084 (N_29084,N_20893,N_21839);
nand U29085 (N_29085,N_22744,N_22312);
nand U29086 (N_29086,N_21121,N_23724);
nor U29087 (N_29087,N_18704,N_22249);
nand U29088 (N_29088,N_19867,N_20172);
or U29089 (N_29089,N_18915,N_22871);
and U29090 (N_29090,N_21724,N_21343);
nor U29091 (N_29091,N_22690,N_19397);
or U29092 (N_29092,N_20092,N_20604);
or U29093 (N_29093,N_22235,N_20919);
or U29094 (N_29094,N_19876,N_23078);
nor U29095 (N_29095,N_18032,N_21336);
and U29096 (N_29096,N_21943,N_18893);
or U29097 (N_29097,N_23669,N_21928);
nand U29098 (N_29098,N_19495,N_23987);
xnor U29099 (N_29099,N_19299,N_21816);
nand U29100 (N_29100,N_22751,N_23449);
or U29101 (N_29101,N_19476,N_21556);
or U29102 (N_29102,N_22434,N_23536);
and U29103 (N_29103,N_23403,N_19370);
and U29104 (N_29104,N_18059,N_22160);
or U29105 (N_29105,N_22277,N_23004);
xor U29106 (N_29106,N_20450,N_20053);
or U29107 (N_29107,N_22050,N_21317);
nor U29108 (N_29108,N_20793,N_21171);
nand U29109 (N_29109,N_18026,N_21931);
nand U29110 (N_29110,N_18873,N_18777);
or U29111 (N_29111,N_19034,N_18706);
xnor U29112 (N_29112,N_23005,N_19884);
and U29113 (N_29113,N_23692,N_22641);
or U29114 (N_29114,N_22485,N_23978);
or U29115 (N_29115,N_22386,N_19060);
nand U29116 (N_29116,N_19787,N_21906);
nor U29117 (N_29117,N_18783,N_20615);
nor U29118 (N_29118,N_20619,N_19278);
or U29119 (N_29119,N_19629,N_23659);
or U29120 (N_29120,N_23682,N_20963);
nand U29121 (N_29121,N_20428,N_20033);
nor U29122 (N_29122,N_18456,N_22910);
and U29123 (N_29123,N_18769,N_19188);
nand U29124 (N_29124,N_19903,N_21048);
and U29125 (N_29125,N_19577,N_23857);
nor U29126 (N_29126,N_19266,N_22544);
or U29127 (N_29127,N_18741,N_22315);
nand U29128 (N_29128,N_19335,N_22317);
nand U29129 (N_29129,N_20298,N_18927);
or U29130 (N_29130,N_21084,N_19892);
nand U29131 (N_29131,N_20876,N_19279);
and U29132 (N_29132,N_22705,N_20509);
or U29133 (N_29133,N_21333,N_20504);
nand U29134 (N_29134,N_19240,N_19005);
nor U29135 (N_29135,N_20476,N_21972);
or U29136 (N_29136,N_23123,N_20381);
nor U29137 (N_29137,N_18622,N_21312);
or U29138 (N_29138,N_20036,N_20061);
nand U29139 (N_29139,N_21214,N_22938);
nand U29140 (N_29140,N_23553,N_19883);
or U29141 (N_29141,N_19982,N_20537);
nor U29142 (N_29142,N_22607,N_19621);
xnor U29143 (N_29143,N_21393,N_23492);
and U29144 (N_29144,N_23452,N_18913);
nand U29145 (N_29145,N_20545,N_18455);
nor U29146 (N_29146,N_20914,N_19294);
and U29147 (N_29147,N_22124,N_22469);
nor U29148 (N_29148,N_23612,N_21413);
and U29149 (N_29149,N_19322,N_22884);
and U29150 (N_29150,N_19487,N_22423);
nor U29151 (N_29151,N_22973,N_21715);
nand U29152 (N_29152,N_18431,N_18250);
or U29153 (N_29153,N_23736,N_18399);
and U29154 (N_29154,N_18890,N_20185);
and U29155 (N_29155,N_23440,N_23876);
nand U29156 (N_29156,N_18234,N_23066);
or U29157 (N_29157,N_21393,N_20074);
and U29158 (N_29158,N_20056,N_20277);
nor U29159 (N_29159,N_23717,N_19063);
and U29160 (N_29160,N_18091,N_19318);
and U29161 (N_29161,N_20403,N_19989);
nor U29162 (N_29162,N_21329,N_19441);
nand U29163 (N_29163,N_22017,N_19178);
nor U29164 (N_29164,N_19029,N_18600);
or U29165 (N_29165,N_19141,N_18477);
and U29166 (N_29166,N_23919,N_18488);
nand U29167 (N_29167,N_23135,N_19867);
nand U29168 (N_29168,N_20786,N_22969);
and U29169 (N_29169,N_20185,N_23390);
xnor U29170 (N_29170,N_20614,N_23141);
nor U29171 (N_29171,N_18755,N_21487);
nor U29172 (N_29172,N_18909,N_19003);
nor U29173 (N_29173,N_23018,N_19918);
nand U29174 (N_29174,N_21859,N_19503);
nor U29175 (N_29175,N_23507,N_19251);
nand U29176 (N_29176,N_22191,N_20748);
xor U29177 (N_29177,N_23202,N_22582);
xor U29178 (N_29178,N_18172,N_20583);
nor U29179 (N_29179,N_20426,N_19425);
or U29180 (N_29180,N_19635,N_21741);
and U29181 (N_29181,N_18079,N_18615);
or U29182 (N_29182,N_19120,N_18713);
nand U29183 (N_29183,N_22039,N_20611);
nor U29184 (N_29184,N_19707,N_19161);
xor U29185 (N_29185,N_20126,N_21750);
xor U29186 (N_29186,N_21653,N_22148);
and U29187 (N_29187,N_18006,N_19537);
nor U29188 (N_29188,N_22782,N_20500);
and U29189 (N_29189,N_21353,N_18457);
nand U29190 (N_29190,N_18119,N_23925);
and U29191 (N_29191,N_23922,N_20866);
nand U29192 (N_29192,N_19830,N_18701);
and U29193 (N_29193,N_18565,N_19532);
nand U29194 (N_29194,N_21430,N_19309);
or U29195 (N_29195,N_21224,N_19422);
or U29196 (N_29196,N_18282,N_23455);
xor U29197 (N_29197,N_18204,N_18169);
xor U29198 (N_29198,N_18516,N_21509);
or U29199 (N_29199,N_20990,N_18101);
and U29200 (N_29200,N_22952,N_22065);
and U29201 (N_29201,N_19295,N_23588);
and U29202 (N_29202,N_23246,N_19284);
and U29203 (N_29203,N_19426,N_22297);
or U29204 (N_29204,N_20814,N_22092);
or U29205 (N_29205,N_22884,N_18097);
and U29206 (N_29206,N_21752,N_18459);
nand U29207 (N_29207,N_21088,N_23891);
and U29208 (N_29208,N_18533,N_22748);
and U29209 (N_29209,N_21542,N_20114);
and U29210 (N_29210,N_21168,N_19690);
and U29211 (N_29211,N_19611,N_22173);
nor U29212 (N_29212,N_19112,N_22035);
and U29213 (N_29213,N_23402,N_22802);
nor U29214 (N_29214,N_23480,N_19285);
and U29215 (N_29215,N_20627,N_18482);
and U29216 (N_29216,N_19386,N_21888);
xor U29217 (N_29217,N_18049,N_18833);
nand U29218 (N_29218,N_20954,N_20793);
nor U29219 (N_29219,N_19244,N_18423);
and U29220 (N_29220,N_22461,N_18489);
nor U29221 (N_29221,N_19298,N_23035);
nand U29222 (N_29222,N_22765,N_23056);
and U29223 (N_29223,N_23251,N_18508);
nor U29224 (N_29224,N_19491,N_18111);
or U29225 (N_29225,N_20995,N_19839);
nor U29226 (N_29226,N_21576,N_20055);
nand U29227 (N_29227,N_23560,N_22470);
or U29228 (N_29228,N_23195,N_21595);
nor U29229 (N_29229,N_18755,N_22183);
and U29230 (N_29230,N_20011,N_23330);
or U29231 (N_29231,N_21442,N_19451);
and U29232 (N_29232,N_23557,N_19005);
nand U29233 (N_29233,N_20762,N_19945);
nor U29234 (N_29234,N_22437,N_18465);
nor U29235 (N_29235,N_21582,N_19452);
or U29236 (N_29236,N_20372,N_23710);
xor U29237 (N_29237,N_18657,N_18053);
and U29238 (N_29238,N_22710,N_22803);
and U29239 (N_29239,N_18090,N_22882);
xor U29240 (N_29240,N_23176,N_18546);
or U29241 (N_29241,N_22013,N_22759);
and U29242 (N_29242,N_18588,N_21949);
nor U29243 (N_29243,N_22811,N_21418);
nor U29244 (N_29244,N_23329,N_22259);
and U29245 (N_29245,N_19117,N_20963);
and U29246 (N_29246,N_22525,N_23116);
nor U29247 (N_29247,N_22791,N_23297);
nand U29248 (N_29248,N_21399,N_19949);
and U29249 (N_29249,N_19415,N_20334);
and U29250 (N_29250,N_20039,N_18433);
xor U29251 (N_29251,N_21999,N_21708);
or U29252 (N_29252,N_22443,N_19120);
or U29253 (N_29253,N_18688,N_23967);
or U29254 (N_29254,N_18594,N_22052);
nor U29255 (N_29255,N_18283,N_19978);
and U29256 (N_29256,N_21367,N_20690);
nand U29257 (N_29257,N_19534,N_20994);
nand U29258 (N_29258,N_20072,N_21675);
nor U29259 (N_29259,N_21330,N_21079);
nor U29260 (N_29260,N_19473,N_18980);
nor U29261 (N_29261,N_22891,N_21317);
nand U29262 (N_29262,N_23148,N_23062);
or U29263 (N_29263,N_20473,N_18119);
nor U29264 (N_29264,N_20092,N_21665);
xnor U29265 (N_29265,N_21720,N_22892);
and U29266 (N_29266,N_20479,N_18881);
and U29267 (N_29267,N_22844,N_18544);
or U29268 (N_29268,N_18677,N_21007);
or U29269 (N_29269,N_19116,N_22171);
or U29270 (N_29270,N_18912,N_23598);
or U29271 (N_29271,N_21995,N_22955);
nor U29272 (N_29272,N_23410,N_18024);
and U29273 (N_29273,N_22561,N_21669);
and U29274 (N_29274,N_21648,N_21411);
nand U29275 (N_29275,N_18207,N_22683);
nor U29276 (N_29276,N_20934,N_20866);
or U29277 (N_29277,N_22348,N_19122);
xor U29278 (N_29278,N_19098,N_21835);
nand U29279 (N_29279,N_22721,N_20487);
xor U29280 (N_29280,N_21982,N_20629);
xnor U29281 (N_29281,N_20465,N_18295);
or U29282 (N_29282,N_22150,N_23226);
nand U29283 (N_29283,N_22534,N_22081);
or U29284 (N_29284,N_18108,N_20541);
and U29285 (N_29285,N_18085,N_22801);
and U29286 (N_29286,N_21200,N_21786);
and U29287 (N_29287,N_21238,N_19968);
nor U29288 (N_29288,N_21847,N_21269);
and U29289 (N_29289,N_23785,N_21610);
or U29290 (N_29290,N_23709,N_19663);
or U29291 (N_29291,N_21584,N_21408);
xor U29292 (N_29292,N_19540,N_18146);
xor U29293 (N_29293,N_18181,N_23998);
or U29294 (N_29294,N_21406,N_22593);
nor U29295 (N_29295,N_19296,N_22054);
or U29296 (N_29296,N_19113,N_20236);
or U29297 (N_29297,N_22097,N_19493);
or U29298 (N_29298,N_23959,N_19797);
nor U29299 (N_29299,N_22127,N_20484);
or U29300 (N_29300,N_21081,N_19769);
nor U29301 (N_29301,N_21336,N_23179);
or U29302 (N_29302,N_21289,N_23640);
and U29303 (N_29303,N_22623,N_21703);
nand U29304 (N_29304,N_18819,N_19329);
and U29305 (N_29305,N_18913,N_18050);
nor U29306 (N_29306,N_19857,N_19374);
and U29307 (N_29307,N_21880,N_21435);
or U29308 (N_29308,N_22673,N_19167);
and U29309 (N_29309,N_20996,N_23142);
or U29310 (N_29310,N_22925,N_23740);
xnor U29311 (N_29311,N_19477,N_19228);
nand U29312 (N_29312,N_19437,N_22653);
xor U29313 (N_29313,N_23591,N_22821);
xor U29314 (N_29314,N_19799,N_18221);
nor U29315 (N_29315,N_19031,N_21528);
nand U29316 (N_29316,N_22545,N_18199);
nand U29317 (N_29317,N_19074,N_23007);
or U29318 (N_29318,N_21935,N_18206);
and U29319 (N_29319,N_21973,N_19595);
and U29320 (N_29320,N_18089,N_20476);
nor U29321 (N_29321,N_22039,N_22451);
nand U29322 (N_29322,N_18005,N_21439);
or U29323 (N_29323,N_21885,N_23571);
nand U29324 (N_29324,N_20067,N_20154);
nor U29325 (N_29325,N_18400,N_23529);
nand U29326 (N_29326,N_22182,N_21674);
or U29327 (N_29327,N_22492,N_22220);
nor U29328 (N_29328,N_20819,N_21491);
or U29329 (N_29329,N_20176,N_22825);
nand U29330 (N_29330,N_20869,N_18950);
xnor U29331 (N_29331,N_21806,N_22729);
xnor U29332 (N_29332,N_19553,N_20702);
or U29333 (N_29333,N_23830,N_20355);
nor U29334 (N_29334,N_22585,N_21424);
nand U29335 (N_29335,N_18807,N_18987);
or U29336 (N_29336,N_20147,N_22948);
xor U29337 (N_29337,N_21631,N_19428);
xnor U29338 (N_29338,N_23298,N_19376);
or U29339 (N_29339,N_23375,N_23680);
nor U29340 (N_29340,N_19696,N_23768);
and U29341 (N_29341,N_18476,N_22947);
nand U29342 (N_29342,N_20005,N_19936);
nand U29343 (N_29343,N_18899,N_22593);
xnor U29344 (N_29344,N_20684,N_23683);
nor U29345 (N_29345,N_20562,N_20015);
or U29346 (N_29346,N_19963,N_19939);
or U29347 (N_29347,N_20183,N_22883);
nand U29348 (N_29348,N_21993,N_19120);
and U29349 (N_29349,N_18695,N_18341);
or U29350 (N_29350,N_21322,N_19757);
and U29351 (N_29351,N_19773,N_23994);
or U29352 (N_29352,N_19094,N_19122);
and U29353 (N_29353,N_21153,N_22755);
and U29354 (N_29354,N_23683,N_18692);
or U29355 (N_29355,N_20635,N_20101);
nor U29356 (N_29356,N_18862,N_19642);
nor U29357 (N_29357,N_20989,N_20820);
and U29358 (N_29358,N_18558,N_20587);
nand U29359 (N_29359,N_20573,N_23646);
or U29360 (N_29360,N_19796,N_18008);
nand U29361 (N_29361,N_23451,N_18100);
or U29362 (N_29362,N_23338,N_20884);
nand U29363 (N_29363,N_22801,N_21265);
nor U29364 (N_29364,N_22174,N_23098);
nor U29365 (N_29365,N_20665,N_23880);
or U29366 (N_29366,N_18706,N_18834);
or U29367 (N_29367,N_18697,N_18801);
or U29368 (N_29368,N_21521,N_22492);
xor U29369 (N_29369,N_21411,N_23248);
or U29370 (N_29370,N_22183,N_19705);
nor U29371 (N_29371,N_23100,N_18126);
nand U29372 (N_29372,N_23227,N_19648);
nor U29373 (N_29373,N_22444,N_19721);
xnor U29374 (N_29374,N_19167,N_22376);
and U29375 (N_29375,N_21261,N_21890);
nand U29376 (N_29376,N_20571,N_20409);
or U29377 (N_29377,N_21316,N_22721);
nand U29378 (N_29378,N_22911,N_20333);
nand U29379 (N_29379,N_21365,N_22696);
and U29380 (N_29380,N_22359,N_21873);
and U29381 (N_29381,N_18577,N_23538);
and U29382 (N_29382,N_18019,N_22285);
or U29383 (N_29383,N_22090,N_21866);
and U29384 (N_29384,N_21001,N_20778);
nand U29385 (N_29385,N_19984,N_21459);
and U29386 (N_29386,N_21048,N_22431);
or U29387 (N_29387,N_21553,N_18157);
and U29388 (N_29388,N_23647,N_21494);
and U29389 (N_29389,N_20706,N_23578);
nand U29390 (N_29390,N_21438,N_23618);
nor U29391 (N_29391,N_20546,N_23982);
or U29392 (N_29392,N_18983,N_18363);
xnor U29393 (N_29393,N_22877,N_19784);
and U29394 (N_29394,N_23635,N_23244);
nand U29395 (N_29395,N_22308,N_19258);
or U29396 (N_29396,N_20352,N_20296);
nand U29397 (N_29397,N_18301,N_22714);
and U29398 (N_29398,N_22769,N_18393);
nor U29399 (N_29399,N_22262,N_19154);
nor U29400 (N_29400,N_18375,N_18104);
nand U29401 (N_29401,N_20422,N_20608);
or U29402 (N_29402,N_21606,N_22407);
nand U29403 (N_29403,N_19804,N_23223);
or U29404 (N_29404,N_19097,N_23323);
or U29405 (N_29405,N_23760,N_21497);
and U29406 (N_29406,N_18770,N_22990);
or U29407 (N_29407,N_18322,N_19382);
xnor U29408 (N_29408,N_23085,N_20771);
or U29409 (N_29409,N_22985,N_22757);
nand U29410 (N_29410,N_19848,N_22844);
nor U29411 (N_29411,N_21505,N_23588);
nor U29412 (N_29412,N_21921,N_20693);
nand U29413 (N_29413,N_23447,N_23943);
and U29414 (N_29414,N_20873,N_19619);
nor U29415 (N_29415,N_19836,N_21216);
nand U29416 (N_29416,N_19826,N_23811);
and U29417 (N_29417,N_22820,N_18224);
xnor U29418 (N_29418,N_19375,N_21850);
xor U29419 (N_29419,N_18085,N_18916);
nand U29420 (N_29420,N_20122,N_22968);
or U29421 (N_29421,N_23937,N_21479);
and U29422 (N_29422,N_20737,N_19235);
and U29423 (N_29423,N_18109,N_18368);
or U29424 (N_29424,N_18124,N_22960);
xnor U29425 (N_29425,N_20307,N_21233);
and U29426 (N_29426,N_19296,N_20470);
and U29427 (N_29427,N_23336,N_22252);
and U29428 (N_29428,N_21398,N_22220);
xor U29429 (N_29429,N_18447,N_21251);
and U29430 (N_29430,N_22974,N_19338);
or U29431 (N_29431,N_18479,N_23718);
or U29432 (N_29432,N_20318,N_19739);
nor U29433 (N_29433,N_20387,N_23614);
nand U29434 (N_29434,N_22867,N_23416);
or U29435 (N_29435,N_19051,N_23233);
nor U29436 (N_29436,N_21328,N_21838);
nor U29437 (N_29437,N_21121,N_22709);
nand U29438 (N_29438,N_21614,N_18040);
nor U29439 (N_29439,N_19274,N_20990);
nand U29440 (N_29440,N_18656,N_23064);
and U29441 (N_29441,N_18762,N_21184);
and U29442 (N_29442,N_21127,N_22749);
xnor U29443 (N_29443,N_20999,N_20646);
nand U29444 (N_29444,N_23032,N_19254);
nor U29445 (N_29445,N_22098,N_22897);
or U29446 (N_29446,N_22299,N_23329);
nor U29447 (N_29447,N_20860,N_22307);
xnor U29448 (N_29448,N_18576,N_20771);
and U29449 (N_29449,N_18868,N_20841);
and U29450 (N_29450,N_22809,N_19399);
nor U29451 (N_29451,N_19925,N_19962);
or U29452 (N_29452,N_20972,N_20989);
xor U29453 (N_29453,N_22057,N_21384);
or U29454 (N_29454,N_21215,N_23069);
and U29455 (N_29455,N_20146,N_19287);
nor U29456 (N_29456,N_21674,N_21787);
or U29457 (N_29457,N_19814,N_22578);
nor U29458 (N_29458,N_21680,N_21901);
xnor U29459 (N_29459,N_21313,N_22740);
nor U29460 (N_29460,N_19784,N_23175);
and U29461 (N_29461,N_23800,N_19066);
or U29462 (N_29462,N_21292,N_22991);
or U29463 (N_29463,N_23065,N_22303);
nand U29464 (N_29464,N_19545,N_20807);
nand U29465 (N_29465,N_22980,N_19734);
nor U29466 (N_29466,N_22127,N_22395);
or U29467 (N_29467,N_19890,N_18149);
xor U29468 (N_29468,N_21154,N_20464);
and U29469 (N_29469,N_19406,N_20742);
nand U29470 (N_29470,N_18998,N_22778);
or U29471 (N_29471,N_21017,N_20655);
nor U29472 (N_29472,N_18210,N_20972);
and U29473 (N_29473,N_20423,N_21913);
or U29474 (N_29474,N_20753,N_20485);
nor U29475 (N_29475,N_19744,N_20337);
nand U29476 (N_29476,N_18869,N_19300);
nor U29477 (N_29477,N_22024,N_22032);
or U29478 (N_29478,N_23011,N_22354);
and U29479 (N_29479,N_23425,N_19848);
nand U29480 (N_29480,N_18760,N_19374);
nand U29481 (N_29481,N_19512,N_21799);
or U29482 (N_29482,N_21003,N_22380);
nand U29483 (N_29483,N_19361,N_19022);
nor U29484 (N_29484,N_22998,N_23673);
and U29485 (N_29485,N_19677,N_20993);
nor U29486 (N_29486,N_19477,N_20687);
or U29487 (N_29487,N_21698,N_20727);
xor U29488 (N_29488,N_20215,N_21291);
and U29489 (N_29489,N_20870,N_21740);
nand U29490 (N_29490,N_23044,N_21663);
nand U29491 (N_29491,N_19994,N_18853);
and U29492 (N_29492,N_23558,N_19798);
and U29493 (N_29493,N_22879,N_19172);
xnor U29494 (N_29494,N_19296,N_18408);
nand U29495 (N_29495,N_22226,N_22395);
nor U29496 (N_29496,N_21986,N_20337);
nor U29497 (N_29497,N_23976,N_23173);
nor U29498 (N_29498,N_18142,N_21292);
nand U29499 (N_29499,N_22911,N_22985);
or U29500 (N_29500,N_20241,N_22063);
and U29501 (N_29501,N_23462,N_21525);
nand U29502 (N_29502,N_23929,N_21731);
nand U29503 (N_29503,N_21460,N_22345);
and U29504 (N_29504,N_18449,N_19483);
nand U29505 (N_29505,N_20243,N_20667);
or U29506 (N_29506,N_23045,N_20103);
or U29507 (N_29507,N_21141,N_20662);
nor U29508 (N_29508,N_23923,N_22209);
and U29509 (N_29509,N_19228,N_19834);
xnor U29510 (N_29510,N_18739,N_23906);
xnor U29511 (N_29511,N_22480,N_22211);
and U29512 (N_29512,N_21488,N_18588);
and U29513 (N_29513,N_18674,N_23993);
nor U29514 (N_29514,N_19998,N_21723);
nand U29515 (N_29515,N_18688,N_21411);
nand U29516 (N_29516,N_19094,N_19993);
nor U29517 (N_29517,N_23473,N_21543);
nor U29518 (N_29518,N_23463,N_22196);
nand U29519 (N_29519,N_20810,N_22567);
nor U29520 (N_29520,N_18744,N_20571);
and U29521 (N_29521,N_19078,N_18800);
and U29522 (N_29522,N_19211,N_21878);
nor U29523 (N_29523,N_18880,N_21706);
nand U29524 (N_29524,N_22734,N_18533);
and U29525 (N_29525,N_22608,N_21189);
xnor U29526 (N_29526,N_20066,N_21033);
xnor U29527 (N_29527,N_22844,N_23656);
or U29528 (N_29528,N_19293,N_20472);
and U29529 (N_29529,N_20732,N_23870);
or U29530 (N_29530,N_21576,N_18965);
nor U29531 (N_29531,N_19733,N_21532);
nor U29532 (N_29532,N_23190,N_23026);
and U29533 (N_29533,N_18269,N_20247);
and U29534 (N_29534,N_19664,N_18055);
nor U29535 (N_29535,N_18326,N_23540);
or U29536 (N_29536,N_23532,N_21811);
or U29537 (N_29537,N_23376,N_18120);
xor U29538 (N_29538,N_19986,N_23337);
xnor U29539 (N_29539,N_18581,N_19926);
and U29540 (N_29540,N_21569,N_20562);
nand U29541 (N_29541,N_22961,N_22669);
and U29542 (N_29542,N_22359,N_21243);
and U29543 (N_29543,N_23154,N_19050);
xnor U29544 (N_29544,N_20578,N_19911);
and U29545 (N_29545,N_21587,N_18058);
xor U29546 (N_29546,N_18440,N_23330);
or U29547 (N_29547,N_20333,N_22097);
nor U29548 (N_29548,N_22068,N_19893);
nor U29549 (N_29549,N_18160,N_19250);
xor U29550 (N_29550,N_23225,N_20369);
nor U29551 (N_29551,N_19866,N_18818);
nor U29552 (N_29552,N_18430,N_22354);
xor U29553 (N_29553,N_20045,N_22222);
nand U29554 (N_29554,N_23304,N_20825);
and U29555 (N_29555,N_18394,N_19768);
nor U29556 (N_29556,N_18451,N_18825);
nand U29557 (N_29557,N_18592,N_19805);
xnor U29558 (N_29558,N_23234,N_20522);
and U29559 (N_29559,N_20757,N_18840);
nor U29560 (N_29560,N_20388,N_21099);
xnor U29561 (N_29561,N_23363,N_23728);
or U29562 (N_29562,N_18081,N_19743);
or U29563 (N_29563,N_21992,N_18852);
nand U29564 (N_29564,N_19119,N_23799);
xnor U29565 (N_29565,N_23500,N_22201);
nor U29566 (N_29566,N_23814,N_22412);
or U29567 (N_29567,N_22905,N_19715);
xnor U29568 (N_29568,N_23604,N_22302);
and U29569 (N_29569,N_23037,N_23476);
xnor U29570 (N_29570,N_22159,N_22225);
or U29571 (N_29571,N_20534,N_23457);
xnor U29572 (N_29572,N_18619,N_19151);
or U29573 (N_29573,N_18029,N_23248);
nor U29574 (N_29574,N_20896,N_22614);
or U29575 (N_29575,N_19024,N_19407);
nor U29576 (N_29576,N_18866,N_19198);
and U29577 (N_29577,N_22392,N_18955);
nand U29578 (N_29578,N_21892,N_22712);
and U29579 (N_29579,N_21450,N_19630);
nand U29580 (N_29580,N_18433,N_18293);
or U29581 (N_29581,N_22934,N_20685);
nor U29582 (N_29582,N_21750,N_20945);
and U29583 (N_29583,N_18001,N_19008);
nor U29584 (N_29584,N_18754,N_18004);
nand U29585 (N_29585,N_21449,N_19627);
and U29586 (N_29586,N_18150,N_22426);
and U29587 (N_29587,N_19625,N_23445);
and U29588 (N_29588,N_22346,N_21969);
xor U29589 (N_29589,N_21615,N_19051);
nor U29590 (N_29590,N_20117,N_22272);
xor U29591 (N_29591,N_18804,N_20795);
xnor U29592 (N_29592,N_22335,N_21315);
nor U29593 (N_29593,N_22690,N_18527);
xor U29594 (N_29594,N_22232,N_22727);
nand U29595 (N_29595,N_21623,N_21332);
or U29596 (N_29596,N_18524,N_23353);
nor U29597 (N_29597,N_18180,N_20633);
and U29598 (N_29598,N_20433,N_21074);
nand U29599 (N_29599,N_20603,N_18332);
xor U29600 (N_29600,N_20539,N_18365);
xnor U29601 (N_29601,N_20369,N_18171);
or U29602 (N_29602,N_22941,N_21732);
nor U29603 (N_29603,N_23373,N_23360);
nand U29604 (N_29604,N_19966,N_20633);
nor U29605 (N_29605,N_22755,N_21978);
and U29606 (N_29606,N_22053,N_19443);
and U29607 (N_29607,N_22066,N_21783);
nor U29608 (N_29608,N_21225,N_20033);
nand U29609 (N_29609,N_18646,N_23213);
nand U29610 (N_29610,N_18860,N_19281);
and U29611 (N_29611,N_18005,N_19797);
or U29612 (N_29612,N_18693,N_20242);
or U29613 (N_29613,N_21337,N_21467);
nand U29614 (N_29614,N_20266,N_22433);
xnor U29615 (N_29615,N_18760,N_18648);
xnor U29616 (N_29616,N_22427,N_20750);
nor U29617 (N_29617,N_21343,N_22757);
nand U29618 (N_29618,N_18327,N_23142);
xnor U29619 (N_29619,N_22911,N_20869);
nand U29620 (N_29620,N_20462,N_23072);
nand U29621 (N_29621,N_21789,N_18192);
nor U29622 (N_29622,N_22568,N_21921);
and U29623 (N_29623,N_18401,N_21275);
and U29624 (N_29624,N_23566,N_23925);
or U29625 (N_29625,N_20626,N_20532);
or U29626 (N_29626,N_21777,N_23681);
or U29627 (N_29627,N_21474,N_22895);
nand U29628 (N_29628,N_21277,N_18969);
xor U29629 (N_29629,N_18434,N_20383);
or U29630 (N_29630,N_20135,N_23586);
xor U29631 (N_29631,N_23695,N_23852);
and U29632 (N_29632,N_19040,N_18319);
xor U29633 (N_29633,N_18513,N_21828);
nand U29634 (N_29634,N_23094,N_19681);
nor U29635 (N_29635,N_19684,N_21016);
or U29636 (N_29636,N_18077,N_18036);
and U29637 (N_29637,N_19062,N_22371);
or U29638 (N_29638,N_18259,N_22553);
and U29639 (N_29639,N_21229,N_21301);
xor U29640 (N_29640,N_21884,N_20899);
xor U29641 (N_29641,N_21695,N_18854);
and U29642 (N_29642,N_21067,N_20093);
and U29643 (N_29643,N_21053,N_21402);
xor U29644 (N_29644,N_18606,N_20107);
and U29645 (N_29645,N_23728,N_19916);
and U29646 (N_29646,N_22968,N_20952);
and U29647 (N_29647,N_19698,N_18789);
or U29648 (N_29648,N_19758,N_21729);
nor U29649 (N_29649,N_21716,N_22277);
xnor U29650 (N_29650,N_19126,N_18772);
xor U29651 (N_29651,N_20171,N_22589);
and U29652 (N_29652,N_20984,N_22026);
and U29653 (N_29653,N_22324,N_23525);
nor U29654 (N_29654,N_20615,N_23616);
nor U29655 (N_29655,N_21448,N_21261);
nand U29656 (N_29656,N_19278,N_22277);
and U29657 (N_29657,N_23858,N_22215);
and U29658 (N_29658,N_19704,N_20473);
and U29659 (N_29659,N_22273,N_20595);
nand U29660 (N_29660,N_19372,N_20249);
xnor U29661 (N_29661,N_19187,N_19510);
or U29662 (N_29662,N_23815,N_21609);
and U29663 (N_29663,N_22800,N_19309);
or U29664 (N_29664,N_21565,N_19409);
and U29665 (N_29665,N_19627,N_20021);
nand U29666 (N_29666,N_18577,N_18757);
nand U29667 (N_29667,N_22571,N_18931);
nand U29668 (N_29668,N_18836,N_22665);
or U29669 (N_29669,N_22090,N_18687);
or U29670 (N_29670,N_18554,N_20065);
and U29671 (N_29671,N_18140,N_21452);
and U29672 (N_29672,N_20775,N_21508);
or U29673 (N_29673,N_22176,N_19599);
and U29674 (N_29674,N_22419,N_18349);
nor U29675 (N_29675,N_21929,N_23012);
xnor U29676 (N_29676,N_20129,N_20142);
and U29677 (N_29677,N_20185,N_18967);
and U29678 (N_29678,N_19705,N_18249);
or U29679 (N_29679,N_18682,N_18675);
xor U29680 (N_29680,N_23948,N_19754);
or U29681 (N_29681,N_23116,N_19678);
or U29682 (N_29682,N_19629,N_18381);
nor U29683 (N_29683,N_23063,N_22129);
nor U29684 (N_29684,N_23355,N_20295);
and U29685 (N_29685,N_19995,N_21322);
and U29686 (N_29686,N_18636,N_20402);
nor U29687 (N_29687,N_20861,N_22394);
and U29688 (N_29688,N_23325,N_22876);
nor U29689 (N_29689,N_20373,N_21199);
and U29690 (N_29690,N_21616,N_20098);
and U29691 (N_29691,N_18096,N_19565);
or U29692 (N_29692,N_21238,N_20464);
or U29693 (N_29693,N_20798,N_20593);
or U29694 (N_29694,N_20695,N_18072);
or U29695 (N_29695,N_20764,N_20557);
or U29696 (N_29696,N_18911,N_18289);
and U29697 (N_29697,N_19120,N_19544);
nand U29698 (N_29698,N_19679,N_19770);
and U29699 (N_29699,N_19777,N_22016);
nor U29700 (N_29700,N_21736,N_19879);
nand U29701 (N_29701,N_18644,N_22910);
nand U29702 (N_29702,N_19387,N_19971);
xnor U29703 (N_29703,N_22171,N_21445);
or U29704 (N_29704,N_19719,N_23436);
nand U29705 (N_29705,N_18637,N_22953);
and U29706 (N_29706,N_18530,N_21730);
nor U29707 (N_29707,N_22796,N_19432);
nor U29708 (N_29708,N_20232,N_23176);
nand U29709 (N_29709,N_21631,N_19199);
or U29710 (N_29710,N_21740,N_22638);
nor U29711 (N_29711,N_19622,N_22046);
nand U29712 (N_29712,N_20096,N_22088);
or U29713 (N_29713,N_20933,N_18507);
nor U29714 (N_29714,N_22005,N_23930);
nand U29715 (N_29715,N_23191,N_20327);
or U29716 (N_29716,N_19726,N_21377);
and U29717 (N_29717,N_20378,N_22639);
nor U29718 (N_29718,N_23227,N_22688);
nand U29719 (N_29719,N_18590,N_19317);
and U29720 (N_29720,N_23165,N_23188);
or U29721 (N_29721,N_18288,N_20986);
nand U29722 (N_29722,N_23243,N_19329);
and U29723 (N_29723,N_21454,N_22169);
nor U29724 (N_29724,N_20073,N_19969);
nand U29725 (N_29725,N_22296,N_21114);
nand U29726 (N_29726,N_22729,N_19734);
and U29727 (N_29727,N_22315,N_22537);
or U29728 (N_29728,N_21885,N_19398);
nand U29729 (N_29729,N_23124,N_19910);
nor U29730 (N_29730,N_23604,N_20515);
nor U29731 (N_29731,N_22619,N_19457);
nor U29732 (N_29732,N_22563,N_21822);
nand U29733 (N_29733,N_20285,N_23291);
nor U29734 (N_29734,N_23001,N_19406);
and U29735 (N_29735,N_21603,N_22673);
nand U29736 (N_29736,N_22424,N_20352);
nor U29737 (N_29737,N_21079,N_22658);
and U29738 (N_29738,N_22237,N_19242);
or U29739 (N_29739,N_20164,N_22125);
or U29740 (N_29740,N_22116,N_19538);
nor U29741 (N_29741,N_21271,N_22864);
nand U29742 (N_29742,N_20630,N_23503);
and U29743 (N_29743,N_20634,N_20481);
and U29744 (N_29744,N_18738,N_20810);
nand U29745 (N_29745,N_23833,N_23308);
nor U29746 (N_29746,N_21502,N_22675);
or U29747 (N_29747,N_19324,N_21676);
or U29748 (N_29748,N_18112,N_23641);
nor U29749 (N_29749,N_19291,N_19628);
nor U29750 (N_29750,N_18502,N_22737);
or U29751 (N_29751,N_23539,N_19658);
xnor U29752 (N_29752,N_20840,N_21446);
or U29753 (N_29753,N_22365,N_20825);
nand U29754 (N_29754,N_19358,N_20522);
xnor U29755 (N_29755,N_23137,N_22834);
or U29756 (N_29756,N_20665,N_22349);
and U29757 (N_29757,N_19475,N_23463);
or U29758 (N_29758,N_23019,N_20210);
nand U29759 (N_29759,N_21476,N_23776);
nand U29760 (N_29760,N_21401,N_18346);
and U29761 (N_29761,N_19732,N_22663);
or U29762 (N_29762,N_23869,N_22431);
or U29763 (N_29763,N_23146,N_22225);
xnor U29764 (N_29764,N_21158,N_20120);
and U29765 (N_29765,N_22124,N_19600);
nor U29766 (N_29766,N_19540,N_22622);
nand U29767 (N_29767,N_21617,N_23388);
or U29768 (N_29768,N_20947,N_19119);
nor U29769 (N_29769,N_21678,N_20383);
or U29770 (N_29770,N_23156,N_19048);
nor U29771 (N_29771,N_23305,N_23714);
nor U29772 (N_29772,N_23354,N_22874);
nor U29773 (N_29773,N_22992,N_18053);
and U29774 (N_29774,N_23867,N_21669);
nand U29775 (N_29775,N_18767,N_20022);
and U29776 (N_29776,N_21375,N_21855);
nor U29777 (N_29777,N_23301,N_21407);
and U29778 (N_29778,N_19550,N_20045);
nand U29779 (N_29779,N_22344,N_21346);
and U29780 (N_29780,N_22310,N_22986);
xnor U29781 (N_29781,N_20156,N_20752);
or U29782 (N_29782,N_18454,N_23021);
nand U29783 (N_29783,N_20994,N_23105);
and U29784 (N_29784,N_23788,N_22520);
nor U29785 (N_29785,N_20369,N_21157);
or U29786 (N_29786,N_21399,N_22183);
xor U29787 (N_29787,N_23219,N_19708);
or U29788 (N_29788,N_20413,N_22146);
nor U29789 (N_29789,N_23946,N_22084);
nand U29790 (N_29790,N_22950,N_19774);
nand U29791 (N_29791,N_23740,N_20301);
nand U29792 (N_29792,N_23520,N_18686);
or U29793 (N_29793,N_20915,N_22030);
and U29794 (N_29794,N_19018,N_21321);
and U29795 (N_29795,N_19605,N_19372);
xor U29796 (N_29796,N_20905,N_21139);
and U29797 (N_29797,N_18521,N_18512);
nor U29798 (N_29798,N_21071,N_19731);
and U29799 (N_29799,N_20514,N_22761);
and U29800 (N_29800,N_21922,N_18913);
nand U29801 (N_29801,N_20814,N_19698);
or U29802 (N_29802,N_21847,N_21951);
nor U29803 (N_29803,N_18279,N_20679);
or U29804 (N_29804,N_23226,N_21209);
or U29805 (N_29805,N_19345,N_22239);
and U29806 (N_29806,N_18451,N_22413);
nand U29807 (N_29807,N_21215,N_19996);
and U29808 (N_29808,N_23931,N_21811);
and U29809 (N_29809,N_18982,N_23331);
nor U29810 (N_29810,N_18753,N_23173);
nor U29811 (N_29811,N_22967,N_19005);
or U29812 (N_29812,N_18537,N_22717);
nor U29813 (N_29813,N_21021,N_21361);
nor U29814 (N_29814,N_23026,N_21572);
xor U29815 (N_29815,N_23417,N_23104);
nor U29816 (N_29816,N_21531,N_20754);
or U29817 (N_29817,N_23293,N_18150);
nand U29818 (N_29818,N_22225,N_19346);
nand U29819 (N_29819,N_22429,N_22650);
nand U29820 (N_29820,N_18812,N_23258);
or U29821 (N_29821,N_23431,N_20980);
nor U29822 (N_29822,N_19055,N_18896);
or U29823 (N_29823,N_18087,N_18043);
and U29824 (N_29824,N_19633,N_22591);
nand U29825 (N_29825,N_22906,N_22557);
nand U29826 (N_29826,N_18917,N_19452);
nand U29827 (N_29827,N_23572,N_20525);
nor U29828 (N_29828,N_23043,N_21841);
or U29829 (N_29829,N_18135,N_18565);
nand U29830 (N_29830,N_20371,N_20607);
or U29831 (N_29831,N_23917,N_20904);
xnor U29832 (N_29832,N_19040,N_22684);
nand U29833 (N_29833,N_21197,N_20162);
nand U29834 (N_29834,N_21890,N_20048);
and U29835 (N_29835,N_20486,N_23152);
or U29836 (N_29836,N_23500,N_21071);
nor U29837 (N_29837,N_22895,N_22417);
and U29838 (N_29838,N_20682,N_18797);
or U29839 (N_29839,N_23908,N_19106);
nand U29840 (N_29840,N_21661,N_21906);
and U29841 (N_29841,N_18821,N_23894);
and U29842 (N_29842,N_23414,N_19296);
or U29843 (N_29843,N_22889,N_21235);
xor U29844 (N_29844,N_23751,N_23130);
nor U29845 (N_29845,N_21990,N_20107);
nand U29846 (N_29846,N_22005,N_23292);
nand U29847 (N_29847,N_20914,N_23452);
xor U29848 (N_29848,N_20164,N_23301);
and U29849 (N_29849,N_23807,N_21832);
and U29850 (N_29850,N_20028,N_22915);
and U29851 (N_29851,N_22891,N_23592);
or U29852 (N_29852,N_22278,N_19384);
and U29853 (N_29853,N_21109,N_18141);
xnor U29854 (N_29854,N_20777,N_19068);
and U29855 (N_29855,N_18771,N_19393);
nor U29856 (N_29856,N_22558,N_21238);
or U29857 (N_29857,N_18540,N_21508);
or U29858 (N_29858,N_19527,N_23127);
nand U29859 (N_29859,N_23636,N_19630);
nand U29860 (N_29860,N_20802,N_20202);
or U29861 (N_29861,N_21570,N_18609);
or U29862 (N_29862,N_20645,N_21443);
nor U29863 (N_29863,N_20414,N_21646);
or U29864 (N_29864,N_19947,N_22619);
nand U29865 (N_29865,N_22316,N_21614);
and U29866 (N_29866,N_22677,N_21095);
nand U29867 (N_29867,N_23688,N_21926);
nor U29868 (N_29868,N_20985,N_21240);
or U29869 (N_29869,N_21950,N_23636);
nor U29870 (N_29870,N_19624,N_23948);
nand U29871 (N_29871,N_19537,N_21373);
nand U29872 (N_29872,N_20910,N_20301);
nand U29873 (N_29873,N_21947,N_23837);
nand U29874 (N_29874,N_18504,N_23973);
xnor U29875 (N_29875,N_21121,N_20532);
nand U29876 (N_29876,N_23175,N_23850);
xnor U29877 (N_29877,N_22849,N_18528);
and U29878 (N_29878,N_22804,N_21749);
xnor U29879 (N_29879,N_22823,N_22759);
nand U29880 (N_29880,N_21592,N_23263);
nand U29881 (N_29881,N_22940,N_19839);
or U29882 (N_29882,N_20124,N_19525);
nor U29883 (N_29883,N_18022,N_20875);
nand U29884 (N_29884,N_21390,N_18554);
or U29885 (N_29885,N_20303,N_23997);
nand U29886 (N_29886,N_22693,N_22424);
nand U29887 (N_29887,N_22064,N_18732);
nand U29888 (N_29888,N_20611,N_21294);
nor U29889 (N_29889,N_22514,N_19580);
xnor U29890 (N_29890,N_18020,N_19721);
and U29891 (N_29891,N_19968,N_22014);
nor U29892 (N_29892,N_22907,N_22637);
or U29893 (N_29893,N_20815,N_23348);
or U29894 (N_29894,N_18293,N_23374);
nor U29895 (N_29895,N_23993,N_23272);
xor U29896 (N_29896,N_23228,N_21962);
or U29897 (N_29897,N_19733,N_20316);
nor U29898 (N_29898,N_22370,N_23342);
nor U29899 (N_29899,N_19479,N_22078);
and U29900 (N_29900,N_22833,N_19682);
and U29901 (N_29901,N_19135,N_20755);
and U29902 (N_29902,N_22032,N_20011);
nor U29903 (N_29903,N_19592,N_20747);
nor U29904 (N_29904,N_18804,N_20169);
nor U29905 (N_29905,N_18405,N_21616);
or U29906 (N_29906,N_21090,N_22612);
nor U29907 (N_29907,N_18031,N_23737);
or U29908 (N_29908,N_18107,N_21404);
or U29909 (N_29909,N_21772,N_18195);
and U29910 (N_29910,N_18026,N_21597);
nand U29911 (N_29911,N_22764,N_20966);
xnor U29912 (N_29912,N_18538,N_22727);
and U29913 (N_29913,N_18298,N_18359);
nand U29914 (N_29914,N_21795,N_21505);
or U29915 (N_29915,N_21572,N_19283);
and U29916 (N_29916,N_22167,N_19933);
or U29917 (N_29917,N_18336,N_21008);
or U29918 (N_29918,N_22749,N_23631);
nand U29919 (N_29919,N_22749,N_19877);
and U29920 (N_29920,N_20035,N_18518);
xnor U29921 (N_29921,N_22333,N_19036);
or U29922 (N_29922,N_23221,N_19441);
or U29923 (N_29923,N_19408,N_23461);
nor U29924 (N_29924,N_22298,N_21356);
and U29925 (N_29925,N_23024,N_19974);
xnor U29926 (N_29926,N_20849,N_21970);
nand U29927 (N_29927,N_22566,N_22140);
or U29928 (N_29928,N_21435,N_18381);
nor U29929 (N_29929,N_22040,N_18099);
and U29930 (N_29930,N_22715,N_23872);
or U29931 (N_29931,N_23730,N_23721);
nor U29932 (N_29932,N_18868,N_19998);
nor U29933 (N_29933,N_22891,N_20708);
xnor U29934 (N_29934,N_20036,N_23868);
and U29935 (N_29935,N_21252,N_21546);
and U29936 (N_29936,N_19329,N_22158);
and U29937 (N_29937,N_21289,N_21467);
nor U29938 (N_29938,N_18389,N_20196);
nand U29939 (N_29939,N_18064,N_22927);
or U29940 (N_29940,N_23329,N_20387);
and U29941 (N_29941,N_18559,N_20622);
and U29942 (N_29942,N_22733,N_21619);
and U29943 (N_29943,N_23821,N_18695);
nor U29944 (N_29944,N_19424,N_23502);
xor U29945 (N_29945,N_19958,N_19472);
nor U29946 (N_29946,N_18802,N_22084);
nand U29947 (N_29947,N_21985,N_21946);
nor U29948 (N_29948,N_19476,N_20964);
nor U29949 (N_29949,N_21420,N_20564);
nand U29950 (N_29950,N_18615,N_22969);
and U29951 (N_29951,N_22356,N_20681);
nand U29952 (N_29952,N_19824,N_20696);
and U29953 (N_29953,N_22881,N_18649);
xor U29954 (N_29954,N_23787,N_18878);
nand U29955 (N_29955,N_19251,N_20540);
nand U29956 (N_29956,N_21972,N_23809);
and U29957 (N_29957,N_20457,N_19079);
and U29958 (N_29958,N_19760,N_23195);
nor U29959 (N_29959,N_22146,N_23360);
and U29960 (N_29960,N_22469,N_18448);
nand U29961 (N_29961,N_21524,N_19398);
or U29962 (N_29962,N_21335,N_23537);
or U29963 (N_29963,N_18972,N_20288);
nor U29964 (N_29964,N_18842,N_20428);
or U29965 (N_29965,N_18888,N_22378);
nand U29966 (N_29966,N_20724,N_18564);
nand U29967 (N_29967,N_18441,N_19478);
or U29968 (N_29968,N_20842,N_20984);
and U29969 (N_29969,N_23703,N_21588);
and U29970 (N_29970,N_19098,N_19349);
nand U29971 (N_29971,N_18421,N_23804);
xor U29972 (N_29972,N_21869,N_21961);
nand U29973 (N_29973,N_20239,N_18379);
nor U29974 (N_29974,N_23408,N_22676);
nand U29975 (N_29975,N_21562,N_21897);
nand U29976 (N_29976,N_20658,N_23254);
or U29977 (N_29977,N_21114,N_22169);
xnor U29978 (N_29978,N_18635,N_18277);
or U29979 (N_29979,N_21196,N_21284);
and U29980 (N_29980,N_22757,N_21906);
nand U29981 (N_29981,N_23177,N_21083);
nor U29982 (N_29982,N_18379,N_23466);
or U29983 (N_29983,N_21139,N_23285);
nand U29984 (N_29984,N_22431,N_21616);
nor U29985 (N_29985,N_19282,N_21092);
or U29986 (N_29986,N_19278,N_19325);
nand U29987 (N_29987,N_18993,N_19743);
nor U29988 (N_29988,N_23083,N_22091);
nor U29989 (N_29989,N_21595,N_20979);
nand U29990 (N_29990,N_21344,N_18688);
nand U29991 (N_29991,N_21835,N_18269);
nand U29992 (N_29992,N_19240,N_19346);
or U29993 (N_29993,N_22103,N_20915);
and U29994 (N_29994,N_22851,N_21822);
nor U29995 (N_29995,N_22350,N_20038);
and U29996 (N_29996,N_23862,N_23645);
nor U29997 (N_29997,N_18113,N_20638);
or U29998 (N_29998,N_23030,N_19992);
and U29999 (N_29999,N_23086,N_22096);
nand UO_0 (O_0,N_29013,N_27001);
nand UO_1 (O_1,N_25639,N_24825);
or UO_2 (O_2,N_26511,N_24590);
and UO_3 (O_3,N_25679,N_25224);
or UO_4 (O_4,N_29772,N_27777);
and UO_5 (O_5,N_29914,N_28812);
or UO_6 (O_6,N_29808,N_24781);
and UO_7 (O_7,N_26420,N_24346);
and UO_8 (O_8,N_27527,N_26415);
or UO_9 (O_9,N_28709,N_25862);
and UO_10 (O_10,N_26468,N_24973);
or UO_11 (O_11,N_27277,N_28669);
or UO_12 (O_12,N_24833,N_29874);
nand UO_13 (O_13,N_27886,N_25201);
and UO_14 (O_14,N_24921,N_28501);
nor UO_15 (O_15,N_24910,N_27599);
or UO_16 (O_16,N_26845,N_27171);
and UO_17 (O_17,N_25252,N_27487);
and UO_18 (O_18,N_26327,N_28701);
xnor UO_19 (O_19,N_27500,N_28279);
or UO_20 (O_20,N_24625,N_24519);
or UO_21 (O_21,N_28602,N_24255);
nand UO_22 (O_22,N_27858,N_28537);
xor UO_23 (O_23,N_24858,N_25002);
and UO_24 (O_24,N_27451,N_28853);
nand UO_25 (O_25,N_29235,N_28273);
or UO_26 (O_26,N_28771,N_28754);
or UO_27 (O_27,N_27908,N_29942);
xnor UO_28 (O_28,N_25307,N_25243);
or UO_29 (O_29,N_28059,N_27581);
nand UO_30 (O_30,N_26212,N_24767);
or UO_31 (O_31,N_28046,N_27540);
xor UO_32 (O_32,N_27133,N_29453);
xnor UO_33 (O_33,N_26432,N_24139);
and UO_34 (O_34,N_29331,N_29594);
and UO_35 (O_35,N_29075,N_27262);
and UO_36 (O_36,N_29306,N_24669);
nor UO_37 (O_37,N_24812,N_28755);
nand UO_38 (O_38,N_28057,N_29302);
nor UO_39 (O_39,N_24146,N_27427);
nor UO_40 (O_40,N_25532,N_28841);
nor UO_41 (O_41,N_26742,N_25955);
nand UO_42 (O_42,N_27663,N_26142);
nand UO_43 (O_43,N_25550,N_25754);
and UO_44 (O_44,N_29139,N_27424);
or UO_45 (O_45,N_25757,N_29563);
or UO_46 (O_46,N_26119,N_28278);
nand UO_47 (O_47,N_26770,N_25063);
and UO_48 (O_48,N_26840,N_29744);
and UO_49 (O_49,N_27218,N_26897);
nand UO_50 (O_50,N_26346,N_27559);
and UO_51 (O_51,N_27420,N_26718);
and UO_52 (O_52,N_26589,N_26905);
nand UO_53 (O_53,N_24309,N_28799);
and UO_54 (O_54,N_28840,N_24397);
and UO_55 (O_55,N_25001,N_28287);
nand UO_56 (O_56,N_27790,N_24140);
nor UO_57 (O_57,N_24680,N_29766);
xnor UO_58 (O_58,N_26019,N_26505);
nand UO_59 (O_59,N_24892,N_29136);
nand UO_60 (O_60,N_27762,N_28026);
nand UO_61 (O_61,N_26532,N_29433);
xor UO_62 (O_62,N_27006,N_28526);
and UO_63 (O_63,N_24211,N_25655);
nor UO_64 (O_64,N_28401,N_27433);
and UO_65 (O_65,N_26210,N_24646);
nand UO_66 (O_66,N_25662,N_24729);
and UO_67 (O_67,N_29183,N_29245);
or UO_68 (O_68,N_29647,N_28130);
and UO_69 (O_69,N_27187,N_29201);
nand UO_70 (O_70,N_27727,N_28941);
nand UO_71 (O_71,N_26353,N_29026);
nand UO_72 (O_72,N_26097,N_27655);
and UO_73 (O_73,N_24580,N_29709);
or UO_74 (O_74,N_28355,N_24064);
or UO_75 (O_75,N_28651,N_29972);
and UO_76 (O_76,N_24434,N_29068);
xor UO_77 (O_77,N_26245,N_29912);
or UO_78 (O_78,N_28164,N_26088);
and UO_79 (O_79,N_25940,N_28765);
or UO_80 (O_80,N_29494,N_29123);
or UO_81 (O_81,N_29582,N_24049);
nor UO_82 (O_82,N_28158,N_27403);
or UO_83 (O_83,N_26025,N_24305);
nor UO_84 (O_84,N_29314,N_27924);
and UO_85 (O_85,N_25588,N_29735);
nand UO_86 (O_86,N_26132,N_26282);
xnor UO_87 (O_87,N_28378,N_27382);
or UO_88 (O_88,N_24558,N_25022);
or UO_89 (O_89,N_24742,N_28752);
xor UO_90 (O_90,N_26670,N_24644);
or UO_91 (O_91,N_28636,N_24935);
xnor UO_92 (O_92,N_28134,N_26572);
nand UO_93 (O_93,N_25815,N_27932);
nor UO_94 (O_94,N_25875,N_25137);
nand UO_95 (O_95,N_24520,N_27351);
xor UO_96 (O_96,N_24642,N_29198);
and UO_97 (O_97,N_27968,N_29910);
nand UO_98 (O_98,N_24426,N_29960);
nor UO_99 (O_99,N_25156,N_25515);
nand UO_100 (O_100,N_29944,N_29679);
and UO_101 (O_101,N_27164,N_24059);
nor UO_102 (O_102,N_28574,N_29119);
nor UO_103 (O_103,N_29603,N_27131);
and UO_104 (O_104,N_28813,N_24659);
or UO_105 (O_105,N_24727,N_25263);
and UO_106 (O_106,N_26872,N_27117);
nand UO_107 (O_107,N_26696,N_29357);
xnor UO_108 (O_108,N_29185,N_25092);
and UO_109 (O_109,N_26404,N_24159);
or UO_110 (O_110,N_27712,N_27666);
nand UO_111 (O_111,N_28339,N_27766);
nand UO_112 (O_112,N_24572,N_25574);
nor UO_113 (O_113,N_25157,N_27544);
xnor UO_114 (O_114,N_24191,N_28247);
xor UO_115 (O_115,N_29963,N_25052);
nor UO_116 (O_116,N_26022,N_25717);
xnor UO_117 (O_117,N_27819,N_29590);
nor UO_118 (O_118,N_24431,N_27018);
nor UO_119 (O_119,N_24410,N_27112);
and UO_120 (O_120,N_27895,N_25682);
or UO_121 (O_121,N_29202,N_26043);
nor UO_122 (O_122,N_28457,N_25031);
xor UO_123 (O_123,N_25169,N_29572);
or UO_124 (O_124,N_28286,N_25238);
nand UO_125 (O_125,N_26943,N_24268);
nand UO_126 (O_126,N_25820,N_28465);
nand UO_127 (O_127,N_27731,N_27838);
and UO_128 (O_128,N_26174,N_27029);
nand UO_129 (O_129,N_26576,N_29975);
and UO_130 (O_130,N_26751,N_28790);
and UO_131 (O_131,N_27616,N_27338);
xnor UO_132 (O_132,N_28095,N_28964);
nor UO_133 (O_133,N_26020,N_26487);
and UO_134 (O_134,N_26545,N_28316);
nand UO_135 (O_135,N_24279,N_27030);
nand UO_136 (O_136,N_27372,N_28647);
nor UO_137 (O_137,N_26323,N_27507);
or UO_138 (O_138,N_28533,N_27169);
nor UO_139 (O_139,N_24396,N_27812);
nor UO_140 (O_140,N_26180,N_26612);
and UO_141 (O_141,N_29806,N_29482);
nor UO_142 (O_142,N_24818,N_24190);
xnor UO_143 (O_143,N_29380,N_26497);
and UO_144 (O_144,N_28528,N_24319);
nand UO_145 (O_145,N_29547,N_27588);
or UO_146 (O_146,N_24399,N_25922);
nand UO_147 (O_147,N_25636,N_27975);
nand UO_148 (O_148,N_27859,N_29058);
and UO_149 (O_149,N_27319,N_25237);
xor UO_150 (O_150,N_25721,N_28221);
or UO_151 (O_151,N_25453,N_27184);
nand UO_152 (O_152,N_29096,N_27677);
and UO_153 (O_153,N_29923,N_27659);
nand UO_154 (O_154,N_24354,N_27770);
or UO_155 (O_155,N_27329,N_27406);
and UO_156 (O_156,N_24372,N_28565);
xnor UO_157 (O_157,N_29631,N_25667);
nor UO_158 (O_158,N_27412,N_26010);
or UO_159 (O_159,N_26396,N_28944);
nor UO_160 (O_160,N_27384,N_26087);
and UO_161 (O_161,N_27037,N_29079);
or UO_162 (O_162,N_28716,N_28139);
nor UO_163 (O_163,N_27389,N_25360);
nor UO_164 (O_164,N_25934,N_25434);
nand UO_165 (O_165,N_25267,N_26229);
xnor UO_166 (O_166,N_24492,N_29325);
nor UO_167 (O_167,N_28326,N_27726);
xor UO_168 (O_168,N_27826,N_26554);
nor UO_169 (O_169,N_24045,N_29409);
xor UO_170 (O_170,N_28567,N_27468);
xor UO_171 (O_171,N_24071,N_29574);
nor UO_172 (O_172,N_29776,N_28855);
nor UO_173 (O_173,N_26832,N_27314);
and UO_174 (O_174,N_29063,N_24238);
nand UO_175 (O_175,N_26739,N_24752);
and UO_176 (O_176,N_29087,N_25025);
or UO_177 (O_177,N_28627,N_26333);
nor UO_178 (O_178,N_25884,N_28118);
nand UO_179 (O_179,N_26698,N_25072);
and UO_180 (O_180,N_25101,N_28839);
or UO_181 (O_181,N_24808,N_27914);
nor UO_182 (O_182,N_26459,N_28746);
nand UO_183 (O_183,N_24289,N_29654);
nor UO_184 (O_184,N_28053,N_26369);
nor UO_185 (O_185,N_27536,N_29286);
and UO_186 (O_186,N_29176,N_24691);
nor UO_187 (O_187,N_24712,N_28304);
nor UO_188 (O_188,N_24814,N_25368);
nor UO_189 (O_189,N_24933,N_29134);
nand UO_190 (O_190,N_26844,N_25767);
nor UO_191 (O_191,N_26846,N_24143);
nor UO_192 (O_192,N_25308,N_25122);
or UO_193 (O_193,N_29977,N_25946);
nor UO_194 (O_194,N_25440,N_27820);
nor UO_195 (O_195,N_26760,N_28676);
nand UO_196 (O_196,N_24504,N_27964);
and UO_197 (O_197,N_26783,N_29738);
nand UO_198 (O_198,N_25818,N_25189);
nor UO_199 (O_199,N_25781,N_25328);
or UO_200 (O_200,N_28129,N_29714);
and UO_201 (O_201,N_25615,N_29678);
nand UO_202 (O_202,N_25829,N_29591);
and UO_203 (O_203,N_28217,N_24332);
nor UO_204 (O_204,N_24724,N_28687);
nand UO_205 (O_205,N_25321,N_25469);
nor UO_206 (O_206,N_26109,N_29150);
or UO_207 (O_207,N_27062,N_29195);
nor UO_208 (O_208,N_28170,N_29327);
nor UO_209 (O_209,N_24710,N_29883);
nor UO_210 (O_210,N_25883,N_27380);
nand UO_211 (O_211,N_29388,N_29816);
or UO_212 (O_212,N_26835,N_24873);
or UO_213 (O_213,N_28033,N_28886);
nor UO_214 (O_214,N_27988,N_25731);
xnor UO_215 (O_215,N_26188,N_24573);
nor UO_216 (O_216,N_28876,N_24650);
nand UO_217 (O_217,N_26304,N_28064);
nor UO_218 (O_218,N_24150,N_27746);
nand UO_219 (O_219,N_29697,N_27682);
nor UO_220 (O_220,N_24389,N_26913);
or UO_221 (O_221,N_25713,N_27881);
nor UO_222 (O_222,N_26699,N_25298);
nor UO_223 (O_223,N_26914,N_24082);
nand UO_224 (O_224,N_29040,N_26221);
nand UO_225 (O_225,N_25316,N_29871);
xnor UO_226 (O_226,N_28420,N_25960);
and UO_227 (O_227,N_25046,N_24334);
nor UO_228 (O_228,N_27723,N_26761);
nor UO_229 (O_229,N_26598,N_24366);
nor UO_230 (O_230,N_29727,N_27186);
nor UO_231 (O_231,N_29199,N_29203);
and UO_232 (O_232,N_29757,N_29720);
and UO_233 (O_233,N_29916,N_29059);
nand UO_234 (O_234,N_26697,N_24732);
nand UO_235 (O_235,N_29159,N_27444);
xnor UO_236 (O_236,N_25044,N_28127);
nor UO_237 (O_237,N_28807,N_29224);
xor UO_238 (O_238,N_27250,N_29476);
or UO_239 (O_239,N_24273,N_25477);
or UO_240 (O_240,N_24666,N_28311);
nor UO_241 (O_241,N_24595,N_26350);
xor UO_242 (O_242,N_29643,N_28830);
or UO_243 (O_243,N_29712,N_29567);
or UO_244 (O_244,N_26652,N_27807);
nor UO_245 (O_245,N_28140,N_25527);
nand UO_246 (O_246,N_25746,N_26377);
nor UO_247 (O_247,N_25782,N_26854);
or UO_248 (O_248,N_24900,N_27260);
and UO_249 (O_249,N_24382,N_24882);
or UO_250 (O_250,N_26682,N_26820);
or UO_251 (O_251,N_25812,N_27896);
nor UO_252 (O_252,N_24805,N_27060);
nand UO_253 (O_253,N_26156,N_24958);
or UO_254 (O_254,N_24367,N_27969);
nor UO_255 (O_255,N_27477,N_24654);
nand UO_256 (O_256,N_26957,N_24117);
nor UO_257 (O_257,N_29905,N_27823);
nand UO_258 (O_258,N_26692,N_28456);
xnor UO_259 (O_259,N_24269,N_26979);
or UO_260 (O_260,N_29921,N_29682);
nand UO_261 (O_261,N_29652,N_28739);
or UO_262 (O_262,N_27765,N_25806);
nor UO_263 (O_263,N_28797,N_25483);
nor UO_264 (O_264,N_27634,N_24097);
nor UO_265 (O_265,N_28280,N_25420);
and UO_266 (O_266,N_25276,N_25445);
or UO_267 (O_267,N_29230,N_29930);
or UO_268 (O_268,N_28474,N_26743);
nor UO_269 (O_269,N_28389,N_25647);
and UO_270 (O_270,N_26825,N_28541);
or UO_271 (O_271,N_25701,N_29463);
or UO_272 (O_272,N_28085,N_28706);
nand UO_273 (O_273,N_26877,N_24449);
nand UO_274 (O_274,N_28804,N_24645);
nand UO_275 (O_275,N_24507,N_29791);
nor UO_276 (O_276,N_26364,N_29098);
or UO_277 (O_277,N_26249,N_25787);
nor UO_278 (O_278,N_25219,N_24701);
nor UO_279 (O_279,N_29022,N_26707);
nand UO_280 (O_280,N_24292,N_24864);
and UO_281 (O_281,N_27108,N_28857);
and UO_282 (O_282,N_25347,N_26449);
nor UO_283 (O_283,N_24824,N_29070);
or UO_284 (O_284,N_27442,N_28897);
and UO_285 (O_285,N_26805,N_28283);
nand UO_286 (O_286,N_26531,N_24920);
nor UO_287 (O_287,N_25974,N_27280);
or UO_288 (O_288,N_26779,N_25043);
nand UO_289 (O_289,N_24158,N_25207);
xnor UO_290 (O_290,N_27463,N_24879);
xor UO_291 (O_291,N_26154,N_27148);
xnor UO_292 (O_292,N_24459,N_25999);
nor UO_293 (O_293,N_25329,N_24829);
nor UO_294 (O_294,N_25489,N_26410);
nand UO_295 (O_295,N_28614,N_25744);
and UO_296 (O_296,N_29583,N_25530);
and UO_297 (O_297,N_29369,N_28492);
and UO_298 (O_298,N_28508,N_28022);
xnor UO_299 (O_299,N_26069,N_25397);
and UO_300 (O_300,N_27097,N_26978);
nor UO_301 (O_301,N_24875,N_28992);
nand UO_302 (O_302,N_29989,N_29089);
nor UO_303 (O_303,N_27564,N_26711);
or UO_304 (O_304,N_25213,N_26349);
nor UO_305 (O_305,N_25649,N_29177);
nand UO_306 (O_306,N_25241,N_25595);
or UO_307 (O_307,N_28579,N_28773);
xnor UO_308 (O_308,N_29876,N_27408);
or UO_309 (O_309,N_25658,N_27920);
or UO_310 (O_310,N_27633,N_26574);
or UO_311 (O_311,N_29609,N_25674);
nand UO_312 (O_312,N_27501,N_26930);
xor UO_313 (O_313,N_25299,N_25763);
nor UO_314 (O_314,N_27627,N_24083);
nand UO_315 (O_315,N_27439,N_26688);
and UO_316 (O_316,N_28106,N_28119);
nand UO_317 (O_317,N_27251,N_28011);
xor UO_318 (O_318,N_29406,N_27789);
nand UO_319 (O_319,N_26970,N_25415);
or UO_320 (O_320,N_29033,N_26057);
nor UO_321 (O_321,N_25194,N_29354);
and UO_322 (O_322,N_27296,N_27566);
nand UO_323 (O_323,N_26360,N_24462);
nor UO_324 (O_324,N_24339,N_28634);
and UO_325 (O_325,N_25210,N_28766);
nand UO_326 (O_326,N_29984,N_26858);
nand UO_327 (O_327,N_28487,N_28268);
and UO_328 (O_328,N_24104,N_29328);
nor UO_329 (O_329,N_24197,N_28562);
nor UO_330 (O_330,N_28785,N_28535);
or UO_331 (O_331,N_25332,N_24192);
nand UO_332 (O_332,N_29676,N_28360);
nor UO_333 (O_333,N_24498,N_27548);
nand UO_334 (O_334,N_24607,N_26017);
xnor UO_335 (O_335,N_24897,N_27786);
nor UO_336 (O_336,N_27986,N_25013);
and UO_337 (O_337,N_24416,N_24976);
nor UO_338 (O_338,N_27554,N_24374);
and UO_339 (O_339,N_28730,N_28426);
or UO_340 (O_340,N_26726,N_29153);
nor UO_341 (O_341,N_25604,N_28100);
and UO_342 (O_342,N_27174,N_25970);
or UO_343 (O_343,N_25150,N_27871);
xnor UO_344 (O_344,N_29379,N_24253);
nand UO_345 (O_345,N_28391,N_28014);
nand UO_346 (O_346,N_24061,N_24582);
nor UO_347 (O_347,N_25467,N_26170);
nand UO_348 (O_348,N_29280,N_25225);
nor UO_349 (O_349,N_29438,N_28851);
nor UO_350 (O_350,N_27537,N_26317);
and UO_351 (O_351,N_28540,N_29037);
nor UO_352 (O_352,N_27707,N_28469);
nor UO_353 (O_353,N_28157,N_25221);
nand UO_354 (O_354,N_24009,N_28743);
nor UO_355 (O_355,N_28073,N_27031);
nor UO_356 (O_356,N_25800,N_28354);
nor UO_357 (O_357,N_25593,N_27341);
or UO_358 (O_358,N_28909,N_28193);
nand UO_359 (O_359,N_25986,N_25838);
nor UO_360 (O_360,N_28173,N_26653);
and UO_361 (O_361,N_27580,N_25660);
nand UO_362 (O_362,N_27141,N_25535);
nand UO_363 (O_363,N_24201,N_25140);
and UO_364 (O_364,N_28745,N_29827);
xor UO_365 (O_365,N_28550,N_25534);
or UO_366 (O_366,N_28156,N_27851);
or UO_367 (O_367,N_29193,N_29394);
and UO_368 (O_368,N_25968,N_26622);
nand UO_369 (O_369,N_24226,N_26237);
nand UO_370 (O_370,N_29352,N_29677);
nor UO_371 (O_371,N_26810,N_29821);
or UO_372 (O_372,N_29725,N_29624);
nor UO_373 (O_373,N_26134,N_29285);
nand UO_374 (O_374,N_24135,N_25635);
or UO_375 (O_375,N_27294,N_29300);
nand UO_376 (O_376,N_29137,N_25661);
and UO_377 (O_377,N_28973,N_26026);
nor UO_378 (O_378,N_27664,N_24916);
and UO_379 (O_379,N_24853,N_25198);
xnor UO_380 (O_380,N_28318,N_28793);
xor UO_381 (O_381,N_26773,N_25878);
nand UO_382 (O_382,N_26721,N_24898);
xnor UO_383 (O_383,N_29383,N_24930);
or UO_384 (O_384,N_25982,N_26150);
and UO_385 (O_385,N_28344,N_28962);
xnor UO_386 (O_386,N_27390,N_25886);
nor UO_387 (O_387,N_28595,N_27149);
and UO_388 (O_388,N_28563,N_27780);
and UO_389 (O_389,N_26626,N_27891);
nor UO_390 (O_390,N_28605,N_26982);
or UO_391 (O_391,N_25645,N_29700);
xor UO_392 (O_392,N_27704,N_28098);
nand UO_393 (O_393,N_25461,N_27953);
nand UO_394 (O_394,N_26926,N_24280);
nand UO_395 (O_395,N_29043,N_26708);
or UO_396 (O_396,N_27009,N_28831);
nor UO_397 (O_397,N_28988,N_26515);
and UO_398 (O_398,N_28892,N_25694);
or UO_399 (O_399,N_26312,N_28586);
nand UO_400 (O_400,N_27379,N_29011);
nand UO_401 (O_401,N_29027,N_29083);
nand UO_402 (O_402,N_28801,N_28300);
nand UO_403 (O_403,N_25866,N_27374);
nor UO_404 (O_404,N_28176,N_25921);
xor UO_405 (O_405,N_29743,N_29852);
nor UO_406 (O_406,N_28809,N_26593);
xor UO_407 (O_407,N_29495,N_24236);
and UO_408 (O_408,N_26544,N_26704);
nor UO_409 (O_409,N_24361,N_28303);
and UO_410 (O_410,N_29164,N_25432);
nand UO_411 (O_411,N_26195,N_27392);
and UO_412 (O_412,N_26512,N_25473);
or UO_413 (O_413,N_27154,N_24544);
or UO_414 (O_414,N_26709,N_26031);
or UO_415 (O_415,N_26809,N_26220);
and UO_416 (O_416,N_28336,N_25429);
nand UO_417 (O_417,N_28088,N_28659);
or UO_418 (O_418,N_29264,N_29315);
and UO_419 (O_419,N_25629,N_26300);
nor UO_420 (O_420,N_28949,N_26651);
nor UO_421 (O_421,N_25652,N_25745);
and UO_422 (O_422,N_28265,N_29407);
or UO_423 (O_423,N_29432,N_29915);
or UO_424 (O_424,N_28001,N_24997);
and UO_425 (O_425,N_25124,N_25363);
xor UO_426 (O_426,N_28666,N_25314);
or UO_427 (O_427,N_29243,N_29389);
nor UO_428 (O_428,N_24835,N_25414);
and UO_429 (O_429,N_27773,N_27049);
and UO_430 (O_430,N_27352,N_27792);
nor UO_431 (O_431,N_29351,N_25438);
xnor UO_432 (O_432,N_24627,N_29387);
nand UO_433 (O_433,N_28428,N_25718);
or UO_434 (O_434,N_29122,N_26103);
nand UO_435 (O_435,N_29219,N_26331);
nor UO_436 (O_436,N_25312,N_25323);
nor UO_437 (O_437,N_26358,N_29667);
nand UO_438 (O_438,N_26680,N_27330);
and UO_439 (O_439,N_27877,N_29061);
or UO_440 (O_440,N_24819,N_27764);
nor UO_441 (O_441,N_29489,N_25603);
nor UO_442 (O_442,N_27729,N_26289);
nand UO_443 (O_443,N_24568,N_24454);
xnor UO_444 (O_444,N_25853,N_26931);
nor UO_445 (O_445,N_25129,N_24993);
and UO_446 (O_446,N_29343,N_27038);
or UO_447 (O_447,N_24421,N_28580);
nor UO_448 (O_448,N_28227,N_28321);
nor UO_449 (O_449,N_26836,N_28864);
and UO_450 (O_450,N_29437,N_27535);
nor UO_451 (O_451,N_29073,N_27606);
or UO_452 (O_452,N_28399,N_25382);
xor UO_453 (O_453,N_28471,N_26984);
nand UO_454 (O_454,N_24092,N_25177);
nand UO_455 (O_455,N_27391,N_27013);
or UO_456 (O_456,N_24424,N_24130);
or UO_457 (O_457,N_25170,N_24655);
nand UO_458 (O_458,N_25117,N_25648);
or UO_459 (O_459,N_29543,N_26351);
nand UO_460 (O_460,N_25497,N_29749);
and UO_461 (O_461,N_24725,N_24484);
and UO_462 (O_462,N_29885,N_24658);
or UO_463 (O_463,N_24551,N_24653);
nor UO_464 (O_464,N_26411,N_26956);
nor UO_465 (O_465,N_25991,N_29307);
and UO_466 (O_466,N_27388,N_26202);
xor UO_467 (O_467,N_25120,N_27309);
nand UO_468 (O_468,N_26679,N_28315);
nor UO_469 (O_469,N_26441,N_25867);
and UO_470 (O_470,N_26038,N_26480);
xor UO_471 (O_471,N_24762,N_24624);
nand UO_472 (O_472,N_24222,N_26791);
or UO_473 (O_473,N_27996,N_26977);
nor UO_474 (O_474,N_27378,N_28932);
nor UO_475 (O_475,N_24861,N_29418);
and UO_476 (O_476,N_25217,N_27364);
nor UO_477 (O_477,N_28365,N_28942);
nor UO_478 (O_478,N_28664,N_27876);
and UO_479 (O_479,N_24053,N_27387);
nor UO_480 (O_480,N_24588,N_29005);
xor UO_481 (O_481,N_27565,N_26246);
nand UO_482 (O_482,N_27063,N_27353);
nand UO_483 (O_483,N_26427,N_26919);
nand UO_484 (O_484,N_28695,N_24657);
or UO_485 (O_485,N_25895,N_29653);
or UO_486 (O_486,N_25011,N_26822);
or UO_487 (O_487,N_24148,N_28343);
or UO_488 (O_488,N_26419,N_27583);
and UO_489 (O_489,N_28685,N_26133);
nand UO_490 (O_490,N_26605,N_24867);
and UO_491 (O_491,N_25919,N_28199);
nand UO_492 (O_492,N_29416,N_28010);
nand UO_493 (O_493,N_27929,N_28258);
and UO_494 (O_494,N_28075,N_28919);
or UO_495 (O_495,N_29329,N_26000);
nand UO_496 (O_496,N_25003,N_27959);
nor UO_497 (O_497,N_27743,N_29324);
or UO_498 (O_498,N_27867,N_27073);
nand UO_499 (O_499,N_25455,N_26291);
nand UO_500 (O_500,N_29943,N_29439);
and UO_501 (O_501,N_25580,N_26391);
nand UO_502 (O_502,N_26586,N_26885);
and UO_503 (O_503,N_29657,N_29385);
and UO_504 (O_504,N_27231,N_27751);
or UO_505 (O_505,N_26749,N_29705);
or UO_506 (O_506,N_26703,N_24084);
or UO_507 (O_507,N_26091,N_28778);
nand UO_508 (O_508,N_26489,N_28214);
or UO_509 (O_509,N_26305,N_24224);
nor UO_510 (O_510,N_28920,N_28103);
xnor UO_511 (O_511,N_25692,N_24055);
nand UO_512 (O_512,N_24038,N_26029);
or UO_513 (O_513,N_26744,N_28259);
and UO_514 (O_514,N_26011,N_29525);
nand UO_515 (O_515,N_29449,N_27472);
and UO_516 (O_516,N_28017,N_29490);
nor UO_517 (O_517,N_29269,N_28111);
nand UO_518 (O_518,N_26082,N_27774);
or UO_519 (O_519,N_25204,N_26362);
or UO_520 (O_520,N_24675,N_28047);
and UO_521 (O_521,N_24744,N_24977);
and UO_522 (O_522,N_24290,N_27703);
nand UO_523 (O_523,N_29655,N_24816);
or UO_524 (O_524,N_25442,N_24510);
or UO_525 (O_525,N_25424,N_27511);
or UO_526 (O_526,N_29411,N_26466);
or UO_527 (O_527,N_26955,N_28043);
nand UO_528 (O_528,N_29771,N_28871);
nor UO_529 (O_529,N_25542,N_28031);
and UO_530 (O_530,N_27356,N_26882);
or UO_531 (O_531,N_27796,N_29443);
and UO_532 (O_532,N_28226,N_26254);
xor UO_533 (O_533,N_29585,N_26128);
and UO_534 (O_534,N_27216,N_25617);
and UO_535 (O_535,N_25049,N_26987);
or UO_536 (O_536,N_29633,N_27393);
nand UO_537 (O_537,N_28246,N_26260);
nand UO_538 (O_538,N_25048,N_24433);
xnor UO_539 (O_539,N_26599,N_27370);
nor UO_540 (O_540,N_27441,N_24872);
nand UO_541 (O_541,N_26204,N_29220);
xnor UO_542 (O_542,N_27575,N_28800);
and UO_543 (O_543,N_26663,N_24956);
nand UO_544 (O_544,N_29455,N_26442);
nand UO_545 (O_545,N_25752,N_29731);
and UO_546 (O_546,N_24960,N_29604);
nor UO_547 (O_547,N_26372,N_27515);
nand UO_548 (O_548,N_25041,N_27652);
nor UO_549 (O_549,N_28067,N_26160);
nor UO_550 (O_550,N_28489,N_28891);
or UO_551 (O_551,N_27948,N_25536);
and UO_552 (O_552,N_24250,N_27022);
nor UO_553 (O_553,N_27613,N_29499);
and UO_554 (O_554,N_24750,N_27455);
nor UO_555 (O_555,N_28546,N_27176);
xor UO_556 (O_556,N_29971,N_28077);
nand UO_557 (O_557,N_28097,N_25641);
or UO_558 (O_558,N_24136,N_27573);
nand UO_559 (O_559,N_29419,N_28682);
or UO_560 (O_560,N_29571,N_28645);
and UO_561 (O_561,N_26898,N_26394);
xor UO_562 (O_562,N_26627,N_28373);
xor UO_563 (O_563,N_26070,N_26929);
or UO_564 (O_564,N_25589,N_28930);
nor UO_565 (O_565,N_27101,N_27568);
and UO_566 (O_566,N_25006,N_28000);
nor UO_567 (O_567,N_25927,N_25923);
and UO_568 (O_568,N_27005,N_29475);
nand UO_569 (O_569,N_27668,N_26365);
xor UO_570 (O_570,N_25582,N_24964);
nand UO_571 (O_571,N_25769,N_25562);
xor UO_572 (O_572,N_25341,N_27274);
nand UO_573 (O_573,N_29382,N_28603);
xnor UO_574 (O_574,N_26499,N_26823);
nand UO_575 (O_575,N_29641,N_28063);
or UO_576 (O_576,N_26073,N_26271);
and UO_577 (O_577,N_26556,N_25309);
nor UO_578 (O_578,N_28460,N_25901);
nor UO_579 (O_579,N_28635,N_24690);
nor UO_580 (O_580,N_24219,N_24941);
and UO_581 (O_581,N_26694,N_28449);
nand UO_582 (O_582,N_29998,N_28548);
or UO_583 (O_583,N_24043,N_25261);
or UO_584 (O_584,N_24783,N_27075);
and UO_585 (O_585,N_26200,N_24472);
nand UO_586 (O_586,N_26722,N_25512);
nand UO_587 (O_587,N_26794,N_24134);
nor UO_588 (O_588,N_24039,N_28314);
nor UO_589 (O_589,N_27227,N_24852);
nor UO_590 (O_590,N_27011,N_25310);
xnor UO_591 (O_591,N_25186,N_28213);
and UO_592 (O_592,N_27856,N_24508);
nor UO_593 (O_593,N_24664,N_24615);
nor UO_594 (O_594,N_27685,N_27576);
nor UO_595 (O_595,N_28609,N_28424);
or UO_596 (O_596,N_25084,N_24463);
and UO_597 (O_597,N_24184,N_26710);
nor UO_598 (O_598,N_28970,N_27878);
and UO_599 (O_599,N_28953,N_29052);
nor UO_600 (O_600,N_28727,N_24788);
nand UO_601 (O_601,N_28590,N_25995);
and UO_602 (O_602,N_29421,N_29355);
nand UO_603 (O_603,N_26398,N_27680);
or UO_604 (O_604,N_28885,N_29162);
nand UO_605 (O_605,N_25872,N_26027);
or UO_606 (O_606,N_24214,N_29982);
or UO_607 (O_607,N_24208,N_25222);
or UO_608 (O_608,N_24357,N_24515);
and UO_609 (O_609,N_28008,N_27153);
nor UO_610 (O_610,N_27273,N_25422);
or UO_611 (O_611,N_26616,N_29229);
nand UO_612 (O_612,N_29194,N_25395);
or UO_613 (O_613,N_28496,N_29822);
nor UO_614 (O_614,N_27990,N_24843);
or UO_615 (O_615,N_29309,N_27542);
nand UO_616 (O_616,N_28589,N_27497);
nand UO_617 (O_617,N_28241,N_27522);
xor UO_618 (O_618,N_27696,N_26129);
nor UO_619 (O_619,N_25680,N_24711);
xnor UO_620 (O_620,N_26386,N_27822);
and UO_621 (O_621,N_28699,N_24436);
and UO_622 (O_622,N_25496,N_27912);
and UO_623 (O_623,N_26460,N_27071);
or UO_624 (O_624,N_28122,N_27242);
xor UO_625 (O_625,N_25778,N_27688);
and UO_626 (O_626,N_24232,N_24423);
nor UO_627 (O_627,N_28395,N_29055);
nor UO_628 (O_628,N_28473,N_25561);
nand UO_629 (O_629,N_25909,N_26437);
nand UO_630 (O_630,N_29875,N_25055);
nand UO_631 (O_631,N_29537,N_27055);
and UO_632 (O_632,N_25608,N_27963);
or UO_633 (O_633,N_29665,N_24322);
or UO_634 (O_634,N_26329,N_27617);
or UO_635 (O_635,N_28498,N_24784);
and UO_636 (O_636,N_28978,N_29492);
or UO_637 (O_637,N_27521,N_27447);
or UO_638 (O_638,N_24975,N_26382);
nor UO_639 (O_639,N_26390,N_29623);
and UO_640 (O_640,N_28741,N_28209);
or UO_641 (O_641,N_24102,N_27753);
and UO_642 (O_642,N_26524,N_26008);
or UO_643 (O_643,N_29114,N_24142);
or UO_644 (O_644,N_24183,N_27452);
and UO_645 (O_645,N_29261,N_25196);
nand UO_646 (O_646,N_28842,N_28517);
nor UO_647 (O_647,N_29393,N_29007);
xor UO_648 (O_648,N_28952,N_27551);
xor UO_649 (O_649,N_24501,N_24164);
nand UO_650 (O_650,N_25231,N_24610);
nand UO_651 (O_651,N_28195,N_27139);
and UO_652 (O_652,N_24386,N_29216);
or UO_653 (O_653,N_25859,N_26002);
xnor UO_654 (O_654,N_26101,N_26403);
or UO_655 (O_655,N_27673,N_26745);
nand UO_656 (O_656,N_25935,N_28215);
or UO_657 (O_657,N_28668,N_25108);
and UO_658 (O_658,N_24700,N_27638);
xnor UO_659 (O_659,N_29844,N_27244);
nand UO_660 (O_660,N_24385,N_28285);
or UO_661 (O_661,N_25594,N_26625);
and UO_662 (O_662,N_28673,N_28686);
or UO_663 (O_663,N_27069,N_26600);
and UO_664 (O_664,N_29505,N_27737);
nor UO_665 (O_665,N_28019,N_25162);
and UO_666 (O_666,N_29105,N_27830);
xnor UO_667 (O_667,N_24972,N_27032);
nor UO_668 (O_668,N_26908,N_25926);
nor UO_669 (O_669,N_25600,N_29884);
nand UO_670 (O_670,N_25475,N_25969);
and UO_671 (O_671,N_27776,N_28431);
nor UO_672 (O_672,N_26159,N_27550);
or UO_673 (O_673,N_29242,N_25056);
xnor UO_674 (O_674,N_29305,N_26378);
nand UO_675 (O_675,N_24632,N_27449);
nand UO_676 (O_676,N_24801,N_24467);
and UO_677 (O_677,N_26292,N_25495);
or UO_678 (O_678,N_27437,N_25032);
or UO_679 (O_679,N_24482,N_26666);
or UO_680 (O_680,N_25180,N_24506);
nand UO_681 (O_681,N_29180,N_29946);
or UO_682 (O_682,N_29395,N_26110);
xor UO_683 (O_683,N_26638,N_28331);
or UO_684 (O_684,N_29637,N_25500);
nand UO_685 (O_685,N_26941,N_29658);
nor UO_686 (O_686,N_28147,N_27313);
nor UO_687 (O_687,N_26602,N_25839);
and UO_688 (O_688,N_24040,N_26958);
or UO_689 (O_689,N_25111,N_28131);
xnor UO_690 (O_690,N_26932,N_29866);
and UO_691 (O_691,N_27930,N_24381);
nand UO_692 (O_692,N_24234,N_27355);
nand UO_693 (O_693,N_28203,N_25856);
nand UO_694 (O_694,N_29131,N_26063);
nand UO_695 (O_695,N_24929,N_26226);
nor UO_696 (O_696,N_29932,N_25961);
and UO_697 (O_697,N_27464,N_25253);
nand UO_698 (O_698,N_25696,N_29190);
nand UO_699 (O_699,N_28994,N_28916);
nand UO_700 (O_700,N_24591,N_25924);
nand UO_701 (O_701,N_26754,N_28534);
nand UO_702 (O_702,N_25824,N_26399);
or UO_703 (O_703,N_26284,N_25739);
xor UO_704 (O_704,N_25064,N_29270);
and UO_705 (O_705,N_29964,N_24612);
nor UO_706 (O_706,N_25411,N_24665);
xor UO_707 (O_707,N_25587,N_26737);
nand UO_708 (O_708,N_29817,N_28881);
and UO_709 (O_709,N_29497,N_26071);
or UO_710 (O_710,N_25791,N_29577);
nor UO_711 (O_711,N_25080,N_24987);
or UO_712 (O_712,N_24739,N_29870);
and UO_713 (O_713,N_26239,N_28704);
nor UO_714 (O_714,N_26776,N_29333);
or UO_715 (O_715,N_27919,N_28822);
and UO_716 (O_716,N_25110,N_24263);
or UO_717 (O_717,N_24266,N_28229);
nor UO_718 (O_718,N_28108,N_24777);
nand UO_719 (O_719,N_27459,N_29109);
xnor UO_720 (O_720,N_28515,N_27697);
or UO_721 (O_721,N_29974,N_27359);
or UO_722 (O_722,N_28132,N_26199);
and UO_723 (O_723,N_25555,N_26185);
and UO_724 (O_724,N_25348,N_28613);
or UO_725 (O_725,N_29528,N_29645);
nand UO_726 (O_726,N_27539,N_24857);
and UO_727 (O_727,N_27208,N_27593);
nor UO_728 (O_728,N_28204,N_26623);
nor UO_729 (O_729,N_24796,N_29689);
and UO_730 (O_730,N_26406,N_28530);
or UO_731 (O_731,N_26764,N_27719);
nand UO_732 (O_732,N_27713,N_25671);
or UO_733 (O_733,N_24817,N_27587);
xor UO_734 (O_734,N_26991,N_29549);
nor UO_735 (O_735,N_28620,N_28197);
and UO_736 (O_736,N_29496,N_25357);
xor UO_737 (O_737,N_25632,N_25279);
or UO_738 (O_738,N_29940,N_26514);
and UO_739 (O_739,N_24791,N_24393);
nand UO_740 (O_740,N_25021,N_29363);
nor UO_741 (O_741,N_25794,N_25342);
and UO_742 (O_742,N_25292,N_29621);
and UO_743 (O_743,N_24155,N_29361);
nor UO_744 (O_744,N_27855,N_28041);
and UO_745 (O_745,N_26853,N_26194);
nand UO_746 (O_746,N_26968,N_29882);
or UO_747 (O_747,N_24233,N_27875);
nand UO_748 (O_748,N_28770,N_28907);
or UO_749 (O_749,N_29523,N_25454);
and UO_750 (O_750,N_26286,N_24713);
xor UO_751 (O_751,N_27426,N_25646);
nand UO_752 (O_752,N_28531,N_25408);
nor UO_753 (O_753,N_25474,N_24850);
and UO_754 (O_754,N_25245,N_24025);
nand UO_755 (O_755,N_27651,N_26322);
or UO_756 (O_756,N_29857,N_25450);
nor UO_757 (O_757,N_26207,N_27937);
and UO_758 (O_758,N_28302,N_26345);
or UO_759 (O_759,N_24167,N_24016);
or UO_760 (O_760,N_24596,N_26062);
or UO_761 (O_761,N_25173,N_24948);
nand UO_762 (O_762,N_29550,N_24517);
or UO_763 (O_763,N_25079,N_26831);
or UO_764 (O_764,N_26829,N_29034);
xnor UO_765 (O_765,N_24493,N_28357);
and UO_766 (O_766,N_29509,N_24387);
nor UO_767 (O_767,N_26232,N_25612);
nor UO_768 (O_768,N_28396,N_24400);
nor UO_769 (O_769,N_27047,N_28025);
nand UO_770 (O_770,N_29558,N_26189);
nand UO_771 (O_771,N_24583,N_26771);
xnor UO_772 (O_772,N_25985,N_29233);
nor UO_773 (O_773,N_26591,N_29398);
and UO_774 (O_774,N_26992,N_29125);
xor UO_775 (O_775,N_27706,N_29763);
and UO_776 (O_776,N_24904,N_26961);
and UO_777 (O_777,N_27124,N_27648);
nor UO_778 (O_778,N_27275,N_27046);
and UO_779 (O_779,N_25010,N_29581);
and UO_780 (O_780,N_28086,N_26099);
and UO_781 (O_781,N_26550,N_28376);
and UO_782 (O_782,N_26479,N_24422);
or UO_783 (O_783,N_27785,N_27065);
and UO_784 (O_784,N_25751,N_25585);
nand UO_785 (O_785,N_26893,N_28600);
or UO_786 (O_786,N_25626,N_27971);
nor UO_787 (O_787,N_27357,N_27629);
and UO_788 (O_788,N_28610,N_25039);
or UO_789 (O_789,N_25758,N_25688);
nand UO_790 (O_790,N_29587,N_27350);
and UO_791 (O_791,N_28044,N_27724);
xor UO_792 (O_792,N_25876,N_25821);
nor UO_793 (O_793,N_26527,N_26861);
or UO_794 (O_794,N_26277,N_27215);
nand UO_795 (O_795,N_27970,N_24660);
nand UO_796 (O_796,N_24513,N_26876);
and UO_797 (O_797,N_24536,N_25159);
or UO_798 (O_798,N_25508,N_24753);
nor UO_799 (O_799,N_24021,N_27041);
and UO_800 (O_800,N_26100,N_27004);
and UO_801 (O_801,N_24859,N_24126);
or UO_802 (O_802,N_29592,N_27135);
xor UO_803 (O_803,N_28838,N_25206);
xor UO_804 (O_804,N_27467,N_24110);
xnor UO_805 (O_805,N_25214,N_27594);
nand UO_806 (O_806,N_28939,N_29559);
xnor UO_807 (O_807,N_28611,N_28738);
and UO_808 (O_808,N_29301,N_27305);
nor UO_809 (O_809,N_26066,N_26243);
nor UO_810 (O_810,N_27730,N_28633);
and UO_811 (O_811,N_25121,N_25619);
nand UO_812 (O_812,N_25716,N_24967);
and UO_813 (O_813,N_28558,N_28958);
and UO_814 (O_814,N_27405,N_28640);
and UO_815 (O_815,N_27528,N_26417);
or UO_816 (O_816,N_27484,N_26308);
and UO_817 (O_817,N_26044,N_25278);
or UO_818 (O_818,N_28547,N_28505);
and UO_819 (O_819,N_26090,N_25601);
and UO_820 (O_820,N_27657,N_25584);
or UO_821 (O_821,N_25401,N_28244);
xor UO_822 (O_822,N_24285,N_29783);
nor UO_823 (O_823,N_26052,N_26018);
nor UO_824 (O_824,N_25766,N_29381);
nand UO_825 (O_825,N_27586,N_28231);
nand UO_826 (O_826,N_24689,N_26227);
xor UO_827 (O_827,N_24810,N_28027);
xor UO_828 (O_828,N_26481,N_28107);
nand UO_829 (O_829,N_25962,N_26015);
nor UO_830 (O_830,N_28753,N_24161);
and UO_831 (O_831,N_26795,N_25714);
and UO_832 (O_832,N_25402,N_25466);
nand UO_833 (O_833,N_24754,N_26454);
nand UO_834 (O_834,N_29601,N_26098);
or UO_835 (O_835,N_28889,N_25786);
nor UO_836 (O_836,N_26533,N_29212);
or UO_837 (O_837,N_24876,N_25834);
and UO_838 (O_838,N_27067,N_29028);
or UO_839 (O_839,N_28594,N_26130);
nand UO_840 (O_840,N_26671,N_25271);
and UO_841 (O_841,N_29196,N_27127);
or UO_842 (O_842,N_28325,N_28358);
xor UO_843 (O_843,N_29717,N_26793);
or UO_844 (O_844,N_24220,N_24878);
xor UO_845 (O_845,N_26388,N_25577);
and UO_846 (O_846,N_26817,N_28912);
and UO_847 (O_847,N_29668,N_24747);
nand UO_848 (O_848,N_26607,N_26092);
nand UO_849 (O_849,N_28710,N_28999);
or UO_850 (O_850,N_28657,N_25825);
nor UO_851 (O_851,N_26565,N_25732);
nand UO_852 (O_852,N_26705,N_24636);
nor UO_853 (O_853,N_28245,N_28732);
nand UO_854 (O_854,N_29427,N_25830);
nor UO_855 (O_855,N_26471,N_26706);
nor UO_856 (O_856,N_26948,N_26314);
xnor UO_857 (O_857,N_25708,N_28483);
nand UO_858 (O_858,N_28989,N_29117);
and UO_859 (O_859,N_24702,N_25605);
or UO_860 (O_860,N_27957,N_28225);
nand UO_861 (O_861,N_29576,N_29755);
and UO_862 (O_862,N_28545,N_28402);
and UO_863 (O_863,N_27577,N_29597);
nand UO_864 (O_864,N_29949,N_28403);
nand UO_865 (O_865,N_27371,N_25836);
nor UO_866 (O_866,N_28649,N_28429);
nand UO_867 (O_867,N_27715,N_27864);
nand UO_868 (O_868,N_29696,N_25695);
nand UO_869 (O_869,N_26393,N_25572);
xnor UO_870 (O_870,N_24453,N_29990);
nand UO_871 (O_871,N_27526,N_27267);
nand UO_872 (O_872,N_28684,N_25967);
or UO_873 (O_873,N_24670,N_24093);
xnor UO_874 (O_874,N_26431,N_24601);
nor UO_875 (O_875,N_28607,N_27222);
and UO_876 (O_876,N_27034,N_27440);
nand UO_877 (O_877,N_27889,N_29672);
and UO_878 (O_878,N_26690,N_27115);
nand UO_879 (O_879,N_27748,N_28322);
xor UO_880 (O_880,N_25272,N_27520);
or UO_881 (O_881,N_27255,N_27331);
nor UO_882 (O_882,N_27519,N_26857);
or UO_883 (O_883,N_27100,N_28142);
or UO_884 (O_884,N_29962,N_29674);
and UO_885 (O_885,N_27888,N_26994);
and UO_886 (O_886,N_26522,N_27532);
nand UO_887 (O_887,N_25760,N_28539);
or UO_888 (O_888,N_25462,N_25089);
nand UO_889 (O_889,N_26476,N_25540);
nand UO_890 (O_890,N_29573,N_27234);
nand UO_891 (O_891,N_29234,N_24345);
nor UO_892 (O_892,N_25560,N_26562);
or UO_893 (O_893,N_26409,N_29046);
nand UO_894 (O_894,N_28954,N_25914);
nor UO_895 (O_895,N_24077,N_29064);
nor UO_896 (O_896,N_29924,N_29215);
nor UO_897 (O_897,N_28705,N_28367);
nand UO_898 (O_898,N_29568,N_26946);
nor UO_899 (O_899,N_26518,N_26149);
or UO_900 (O_900,N_29802,N_25097);
xor UO_901 (O_901,N_29174,N_27805);
xor UO_902 (O_902,N_28291,N_24223);
nand UO_903 (O_903,N_25247,N_25346);
or UO_904 (O_904,N_24838,N_24107);
nor UO_905 (O_905,N_26413,N_25852);
and UO_906 (O_906,N_24602,N_26716);
nand UO_907 (O_907,N_28927,N_24311);
and UO_908 (O_908,N_25663,N_27831);
and UO_909 (O_909,N_25571,N_28902);
or UO_910 (O_910,N_28144,N_28593);
nor UO_911 (O_911,N_24030,N_28650);
and UO_912 (O_912,N_29656,N_26736);
and UO_913 (O_913,N_28836,N_27578);
and UO_914 (O_914,N_29110,N_25803);
and UO_915 (O_915,N_29431,N_25391);
xnor UO_916 (O_916,N_27846,N_26884);
or UO_917 (O_917,N_29630,N_27561);
nor UO_918 (O_918,N_26604,N_26936);
or UO_919 (O_919,N_24687,N_27534);
nor UO_920 (O_920,N_26996,N_27143);
and UO_921 (O_921,N_27717,N_27843);
nor UO_922 (O_922,N_29602,N_28582);
nand UO_923 (O_923,N_26190,N_27934);
nor UO_924 (O_924,N_27460,N_26054);
xnor UO_925 (O_925,N_27798,N_28835);
nor UO_926 (O_926,N_24668,N_25932);
and UO_927 (O_927,N_25707,N_24738);
nand UO_928 (O_928,N_25335,N_27070);
nand UO_929 (O_929,N_24763,N_28604);
and UO_930 (O_930,N_25693,N_29961);
xor UO_931 (O_931,N_29578,N_28368);
nand UO_932 (O_932,N_25738,N_24052);
nand UO_933 (O_933,N_25993,N_24518);
and UO_934 (O_934,N_24696,N_28307);
or UO_935 (O_935,N_29106,N_29742);
or UO_936 (O_936,N_26819,N_28993);
or UO_937 (O_937,N_29464,N_26967);
nor UO_938 (O_938,N_27897,N_28638);
nand UO_939 (O_939,N_29865,N_27755);
and UO_940 (O_940,N_27556,N_28656);
nor UO_941 (O_941,N_24577,N_26023);
nand UO_942 (O_942,N_27192,N_24915);
or UO_943 (O_943,N_27738,N_25524);
nand UO_944 (O_944,N_26715,N_28591);
and UO_945 (O_945,N_29927,N_26414);
nor UO_946 (O_946,N_27960,N_28917);
or UO_947 (O_947,N_24649,N_24047);
nor UO_948 (O_948,N_24537,N_27456);
nor UO_949 (O_949,N_26421,N_28787);
or UO_950 (O_950,N_26049,N_28023);
xor UO_951 (O_951,N_27525,N_29435);
or UO_952 (O_952,N_26267,N_28201);
nor UO_953 (O_953,N_24792,N_24066);
and UO_954 (O_954,N_26513,N_28569);
and UO_955 (O_955,N_24114,N_26974);
and UO_956 (O_956,N_29391,N_29897);
nand UO_957 (O_957,N_24634,N_26186);
nor UO_958 (O_958,N_25069,N_24121);
nand UO_959 (O_959,N_28015,N_28045);
or UO_960 (O_960,N_26447,N_25460);
nor UO_961 (O_961,N_29706,N_29787);
xnor UO_962 (O_962,N_25350,N_25774);
and UO_963 (O_963,N_24974,N_25565);
or UO_964 (O_964,N_27945,N_28516);
nand UO_965 (O_965,N_24476,N_26975);
xnor UO_966 (O_966,N_27835,N_29425);
nand UO_967 (O_967,N_27495,N_26534);
nand UO_968 (O_968,N_28653,N_27861);
and UO_969 (O_969,N_28955,N_29562);
or UO_970 (O_970,N_24619,N_26580);
nor UO_971 (O_971,N_28472,N_25076);
nor UO_972 (O_972,N_27027,N_26564);
xnor UO_973 (O_973,N_27619,N_29794);
nor UO_974 (O_974,N_24428,N_26108);
nor UO_975 (O_975,N_29342,N_29730);
nand UO_976 (O_976,N_27362,N_25487);
nor UO_977 (O_977,N_28342,N_27346);
and UO_978 (O_978,N_24120,N_28925);
and UO_979 (O_979,N_28340,N_26862);
xor UO_980 (O_980,N_28538,N_27611);
and UO_981 (O_981,N_29462,N_24342);
nor UO_982 (O_982,N_24432,N_25863);
or UO_983 (O_983,N_29057,N_24212);
and UO_984 (O_984,N_24001,N_29085);
nand UO_985 (O_985,N_29020,N_27078);
xnor UO_986 (O_986,N_29214,N_28722);
xnor UO_987 (O_987,N_27567,N_28691);
and UO_988 (O_988,N_27496,N_27621);
and UO_989 (O_989,N_24514,N_26916);
nand UO_990 (O_990,N_25447,N_27647);
nand UO_991 (O_991,N_24586,N_26842);
and UO_992 (O_992,N_24041,N_25631);
nand UO_993 (O_993,N_26664,N_25322);
or UO_994 (O_994,N_28646,N_27824);
nor UO_995 (O_995,N_29716,N_24243);
nand UO_996 (O_996,N_29545,N_28102);
nor UO_997 (O_997,N_27003,N_24002);
nand UO_998 (O_998,N_25012,N_26727);
or UO_999 (O_999,N_28443,N_29797);
nand UO_1000 (O_1000,N_28821,N_28254);
nor UO_1001 (O_1001,N_27284,N_26570);
nand UO_1002 (O_1002,N_27498,N_28566);
or UO_1003 (O_1003,N_29246,N_29364);
nor UO_1004 (O_1004,N_25877,N_27524);
and UO_1005 (O_1005,N_25388,N_25390);
nor UO_1006 (O_1006,N_24228,N_26917);
and UO_1007 (O_1007,N_29133,N_27373);
and UO_1008 (O_1008,N_24251,N_25366);
nor UO_1009 (O_1009,N_26944,N_29375);
nand UO_1010 (O_1010,N_26856,N_27081);
and UO_1011 (O_1011,N_25374,N_25179);
and UO_1012 (O_1012,N_27162,N_29769);
nand UO_1013 (O_1013,N_24109,N_27686);
or UO_1014 (O_1014,N_26548,N_27941);
nor UO_1015 (O_1015,N_29127,N_28154);
or UO_1016 (O_1016,N_29831,N_26689);
nor UO_1017 (O_1017,N_24026,N_27584);
nor UO_1018 (O_1018,N_24087,N_24419);
nand UO_1019 (O_1019,N_25065,N_28873);
or UO_1020 (O_1020,N_29588,N_25212);
nor UO_1021 (O_1021,N_29466,N_27221);
nor UO_1022 (O_1022,N_27226,N_27993);
nand UO_1023 (O_1023,N_28629,N_24313);
xor UO_1024 (O_1024,N_29241,N_24769);
nand UO_1025 (O_1025,N_28803,N_24703);
and UO_1026 (O_1026,N_25297,N_24072);
xnor UO_1027 (O_1027,N_26813,N_25433);
nor UO_1028 (O_1028,N_25345,N_28514);
or UO_1029 (O_1029,N_27050,N_29336);
nor UO_1030 (O_1030,N_27560,N_28080);
xor UO_1031 (O_1031,N_25624,N_26559);
nor UO_1032 (O_1032,N_27290,N_24471);
or UO_1033 (O_1033,N_28815,N_28398);
nand UO_1034 (O_1034,N_26297,N_29842);
nor UO_1035 (O_1035,N_27130,N_24237);
and UO_1036 (O_1036,N_26766,N_24605);
nand UO_1037 (O_1037,N_27806,N_27490);
nand UO_1038 (O_1038,N_27312,N_28984);
and UO_1039 (O_1039,N_26553,N_29788);
nand UO_1040 (O_1040,N_28969,N_26552);
nand UO_1041 (O_1041,N_29534,N_27076);
and UO_1042 (O_1042,N_29140,N_29958);
and UO_1043 (O_1043,N_26105,N_28677);
xor UO_1044 (O_1044,N_25592,N_28040);
and UO_1045 (O_1045,N_28500,N_29138);
nand UO_1046 (O_1046,N_28612,N_27269);
xor UO_1047 (O_1047,N_24202,N_28692);
and UO_1048 (O_1048,N_24995,N_27401);
and UO_1049 (O_1049,N_24395,N_25656);
and UO_1050 (O_1050,N_28772,N_24417);
nor UO_1051 (O_1051,N_26950,N_28276);
nand UO_1052 (O_1052,N_26347,N_28592);
nand UO_1053 (O_1053,N_24171,N_29957);
nor UO_1054 (O_1054,N_27261,N_27898);
and UO_1055 (O_1055,N_28135,N_27502);
nor UO_1056 (O_1056,N_25193,N_28105);
or UO_1057 (O_1057,N_25313,N_26136);
or UO_1058 (O_1058,N_24418,N_29488);
nor UO_1059 (O_1059,N_26804,N_24949);
or UO_1060 (O_1060,N_24560,N_27483);
and UO_1061 (O_1061,N_25146,N_25367);
nand UO_1062 (O_1062,N_24466,N_29426);
xor UO_1063 (O_1063,N_25994,N_24896);
or UO_1064 (O_1064,N_28811,N_25490);
nand UO_1065 (O_1065,N_26258,N_27961);
xor UO_1066 (O_1066,N_27955,N_26486);
and UO_1067 (O_1067,N_26535,N_24500);
and UO_1068 (O_1068,N_26077,N_29287);
or UO_1069 (O_1069,N_29413,N_27622);
or UO_1070 (O_1070,N_24926,N_24324);
nand UO_1071 (O_1071,N_25526,N_24343);
nand UO_1072 (O_1072,N_25944,N_28066);
nand UO_1073 (O_1073,N_26678,N_25972);
xor UO_1074 (O_1074,N_29707,N_24398);
or UO_1075 (O_1075,N_27381,N_26458);
nor UO_1076 (O_1076,N_27066,N_29244);
or UO_1077 (O_1077,N_25672,N_27870);
xnor UO_1078 (O_1078,N_29918,N_26597);
or UO_1079 (O_1079,N_27129,N_24782);
and UO_1080 (O_1080,N_28728,N_24841);
nand UO_1081 (O_1081,N_24341,N_27714);
and UO_1082 (O_1082,N_25485,N_28324);
nand UO_1083 (O_1083,N_24272,N_25887);
nand UO_1084 (O_1084,N_27007,N_27292);
nor UO_1085 (O_1085,N_24491,N_24965);
or UO_1086 (O_1086,N_24249,N_26219);
nor UO_1087 (O_1087,N_24478,N_25936);
nor UO_1088 (O_1088,N_27771,N_26288);
nand UO_1089 (O_1089,N_29688,N_26750);
or UO_1090 (O_1090,N_25568,N_29937);
nor UO_1091 (O_1091,N_24057,N_25199);
or UO_1092 (O_1092,N_26763,N_28740);
or UO_1093 (O_1093,N_28731,N_24007);
nand UO_1094 (O_1094,N_28606,N_28751);
xor UO_1095 (O_1095,N_29130,N_25439);
xor UO_1096 (O_1096,N_26102,N_27589);
and UO_1097 (O_1097,N_24592,N_29823);
or UO_1098 (O_1098,N_29856,N_26269);
nor UO_1099 (O_1099,N_24187,N_28419);
or UO_1100 (O_1100,N_26541,N_25128);
or UO_1101 (O_1101,N_28392,N_28940);
nand UO_1102 (O_1102,N_28532,N_25765);
nand UO_1103 (O_1103,N_29761,N_26355);
or UO_1104 (O_1104,N_25285,N_27094);
and UO_1105 (O_1105,N_26865,N_28452);
and UO_1106 (O_1106,N_24800,N_27395);
nand UO_1107 (O_1107,N_27918,N_27344);
or UO_1108 (O_1108,N_24452,N_28165);
and UO_1109 (O_1109,N_27612,N_24244);
or UO_1110 (O_1110,N_28720,N_25274);
and UO_1111 (O_1111,N_28346,N_24248);
and UO_1112 (O_1112,N_24316,N_29877);
nor UO_1113 (O_1113,N_25591,N_29526);
or UO_1114 (O_1114,N_26816,N_24094);
and UO_1115 (O_1115,N_24663,N_25333);
nor UO_1116 (O_1116,N_25358,N_28585);
or UO_1117 (O_1117,N_28824,N_26303);
or UO_1118 (O_1118,N_25220,N_28931);
nand UO_1119 (O_1119,N_24122,N_29044);
nand UO_1120 (O_1120,N_26601,N_28407);
nor UO_1121 (O_1121,N_25814,N_27109);
and UO_1122 (O_1122,N_27833,N_26452);
nor UO_1123 (O_1123,N_24978,N_27596);
and UO_1124 (O_1124,N_26299,N_24137);
and UO_1125 (O_1125,N_28327,N_26575);
or UO_1126 (O_1126,N_29149,N_24524);
nor UO_1127 (O_1127,N_24957,N_24674);
or UO_1128 (O_1128,N_28624,N_29191);
nor UO_1129 (O_1129,N_25393,N_29530);
nand UO_1130 (O_1130,N_27705,N_29423);
and UO_1131 (O_1131,N_27107,N_24199);
xor UO_1132 (O_1132,N_27662,N_28090);
or UO_1133 (O_1133,N_25334,N_25288);
nor UO_1134 (O_1134,N_24027,N_25771);
or UO_1135 (O_1135,N_29451,N_25024);
nand UO_1136 (O_1136,N_27476,N_29554);
and UO_1137 (O_1137,N_29948,N_25865);
nand UO_1138 (O_1138,N_26942,N_24773);
and UO_1139 (O_1139,N_27797,N_29290);
nand UO_1140 (O_1140,N_27874,N_27750);
nand UO_1141 (O_1141,N_26517,N_27473);
xor UO_1142 (O_1142,N_25743,N_24811);
nor UO_1143 (O_1143,N_24401,N_26988);
or UO_1144 (O_1144,N_27400,N_26218);
or UO_1145 (O_1145,N_28002,N_25009);
and UO_1146 (O_1146,N_25563,N_29723);
nor UO_1147 (O_1147,N_25230,N_29186);
and UO_1148 (O_1148,N_24465,N_29900);
and UO_1149 (O_1149,N_29151,N_29084);
nor UO_1150 (O_1150,N_28587,N_25755);
or UO_1151 (O_1151,N_25376,N_28412);
nor UO_1152 (O_1152,N_28178,N_27817);
nand UO_1153 (O_1153,N_24277,N_25318);
nor UO_1154 (O_1154,N_27803,N_24940);
and UO_1155 (O_1155,N_26061,N_27194);
or UO_1156 (O_1156,N_27933,N_25687);
nor UO_1157 (O_1157,N_29440,N_27414);
xnor UO_1158 (O_1158,N_26660,N_25037);
and UO_1159 (O_1159,N_24917,N_24326);
xnor UO_1160 (O_1160,N_25051,N_26191);
xnor UO_1161 (O_1161,N_28110,N_24606);
and UO_1162 (O_1162,N_27513,N_24218);
nor UO_1163 (O_1163,N_28742,N_27821);
nand UO_1164 (O_1164,N_28557,N_27402);
nor UO_1165 (O_1165,N_27615,N_27302);
or UO_1166 (O_1166,N_29935,N_29129);
nor UO_1167 (O_1167,N_26933,N_27479);
or UO_1168 (O_1168,N_24694,N_26283);
xnor UO_1169 (O_1169,N_24221,N_26560);
and UO_1170 (O_1170,N_27946,N_27728);
and UO_1171 (O_1171,N_24446,N_26892);
or UO_1172 (O_1172,N_26266,N_27436);
or UO_1173 (O_1173,N_29751,N_29993);
or UO_1174 (O_1174,N_26045,N_24789);
nand UO_1175 (O_1175,N_29907,N_27811);
nand UO_1176 (O_1176,N_26138,N_26483);
nand UO_1177 (O_1177,N_25392,N_28120);
xnor UO_1178 (O_1178,N_27358,N_24806);
nor UO_1179 (O_1179,N_28869,N_26435);
nand UO_1180 (O_1180,N_26649,N_24023);
nor UO_1181 (O_1181,N_24106,N_27976);
or UO_1182 (O_1182,N_26683,N_26561);
and UO_1183 (O_1183,N_24894,N_26096);
nand UO_1184 (O_1184,N_24716,N_29546);
or UO_1185 (O_1185,N_28083,N_25657);
nor UO_1186 (O_1186,N_25354,N_26168);
xor UO_1187 (O_1187,N_27711,N_29182);
and UO_1188 (O_1188,N_29555,N_24733);
nor UO_1189 (O_1189,N_26500,N_28523);
nor UO_1190 (O_1190,N_24748,N_24240);
or UO_1191 (O_1191,N_27252,N_28832);
and UO_1192 (O_1192,N_26573,N_24242);
nand UO_1193 (O_1193,N_25045,N_28663);
nand UO_1194 (O_1194,N_29206,N_24598);
or UO_1195 (O_1195,N_25950,N_27448);
or UO_1196 (O_1196,N_27386,N_29612);
and UO_1197 (O_1197,N_29811,N_28951);
xor UO_1198 (O_1198,N_26255,N_24616);
nand UO_1199 (O_1199,N_24761,N_28578);
or UO_1200 (O_1200,N_28138,N_29452);
nand UO_1201 (O_1201,N_28476,N_24566);
nand UO_1202 (O_1202,N_26296,N_29729);
and UO_1203 (O_1203,N_27839,N_27377);
xnor UO_1204 (O_1204,N_24304,N_27676);
nor UO_1205 (O_1205,N_24405,N_25183);
or UO_1206 (O_1206,N_28826,N_27745);
nor UO_1207 (O_1207,N_29458,N_24552);
xor UO_1208 (O_1208,N_25522,N_29737);
and UO_1209 (O_1209,N_27678,N_26247);
nor UO_1210 (O_1210,N_26634,N_25819);
or UO_1211 (O_1211,N_24745,N_26046);
nand UO_1212 (O_1212,N_25523,N_29872);
and UO_1213 (O_1213,N_27694,N_25870);
and UO_1214 (O_1214,N_27904,N_26964);
and UO_1215 (O_1215,N_27173,N_29995);
nand UO_1216 (O_1216,N_27229,N_25075);
nand UO_1217 (O_1217,N_29584,N_28126);
or UO_1218 (O_1218,N_27335,N_29893);
and UO_1219 (O_1219,N_24206,N_25899);
or UO_1220 (O_1220,N_26179,N_27533);
and UO_1221 (O_1221,N_29062,N_27253);
nor UO_1222 (O_1222,N_24877,N_26887);
nor UO_1223 (O_1223,N_28104,N_29107);
nand UO_1224 (O_1224,N_26903,N_28099);
and UO_1225 (O_1225,N_25144,N_28658);
nor UO_1226 (O_1226,N_27428,N_28257);
nand UO_1227 (O_1227,N_25706,N_25200);
or UO_1228 (O_1228,N_29892,N_27752);
or UO_1229 (O_1229,N_29818,N_24661);
or UO_1230 (O_1230,N_26492,N_28512);
xnor UO_1231 (O_1231,N_29648,N_26024);
nand UO_1232 (O_1232,N_24581,N_24794);
and UO_1233 (O_1233,N_29168,N_24278);
nand UO_1234 (O_1234,N_24042,N_29289);
nand UO_1235 (O_1235,N_25705,N_24390);
or UO_1236 (O_1236,N_27546,N_25874);
and UO_1237 (O_1237,N_27051,N_26746);
nor UO_1238 (O_1238,N_24575,N_25616);
and UO_1239 (O_1239,N_25416,N_26321);
and UO_1240 (O_1240,N_29113,N_28861);
nand UO_1241 (O_1241,N_28671,N_26089);
and UO_1242 (O_1242,N_28445,N_24578);
xor UO_1243 (O_1243,N_28652,N_28185);
and UO_1244 (O_1244,N_25054,N_25176);
and UO_1245 (O_1245,N_29401,N_24258);
nand UO_1246 (O_1246,N_25407,N_25215);
xor UO_1247 (O_1247,N_26290,N_26843);
and UO_1248 (O_1248,N_29898,N_29311);
or UO_1249 (O_1249,N_25033,N_25971);
nor UO_1250 (O_1250,N_28458,N_24584);
or UO_1251 (O_1251,N_26392,N_24988);
and UO_1252 (O_1252,N_26818,N_29366);
nand UO_1253 (O_1253,N_24011,N_25338);
nor UO_1254 (O_1254,N_29936,N_29675);
and UO_1255 (O_1255,N_25902,N_29158);
nor UO_1256 (O_1256,N_29467,N_24152);
nor UO_1257 (O_1257,N_29666,N_29849);
xor UO_1258 (O_1258,N_24695,N_25690);
xnor UO_1259 (O_1259,N_29260,N_24509);
and UO_1260 (O_1260,N_29634,N_28181);
nand UO_1261 (O_1261,N_27126,N_27572);
nor UO_1262 (O_1262,N_27980,N_24543);
nand UO_1263 (O_1263,N_26401,N_29340);
nor UO_1264 (O_1264,N_29807,N_26332);
nor UO_1265 (O_1265,N_24336,N_28981);
nor UO_1266 (O_1266,N_24626,N_24427);
and UO_1267 (O_1267,N_29448,N_24826);
and UO_1268 (O_1268,N_24299,N_28654);
nand UO_1269 (O_1269,N_24096,N_24490);
or UO_1270 (O_1270,N_26482,N_26960);
nor UO_1271 (O_1271,N_25937,N_24837);
nor UO_1272 (O_1272,N_27396,N_29181);
or UO_1273 (O_1273,N_29500,N_25336);
and UO_1274 (O_1274,N_28136,N_26939);
nor UO_1275 (O_1275,N_26839,N_29446);
and UO_1276 (O_1276,N_29613,N_25471);
or UO_1277 (O_1277,N_27170,N_27104);
xnor UO_1278 (O_1278,N_27695,N_24112);
and UO_1279 (O_1279,N_26808,N_26337);
xor UO_1280 (O_1280,N_29520,N_27906);
nand UO_1281 (O_1281,N_28847,N_28519);
nand UO_1282 (O_1282,N_26782,N_28430);
or UO_1283 (O_1283,N_29535,N_25851);
nor UO_1284 (O_1284,N_26728,N_28141);
or UO_1285 (O_1285,N_28016,N_24648);
or UO_1286 (O_1286,N_26423,N_26259);
nand UO_1287 (O_1287,N_24443,N_24091);
or UO_1288 (O_1288,N_28529,N_24075);
xnor UO_1289 (O_1289,N_25300,N_27445);
or UO_1290 (O_1290,N_29710,N_29460);
nand UO_1291 (O_1291,N_29638,N_28967);
nand UO_1292 (O_1292,N_28418,N_28877);
nand UO_1293 (O_1293,N_27285,N_26446);
nand UO_1294 (O_1294,N_25811,N_25090);
nand UO_1295 (O_1295,N_24899,N_29773);
nor UO_1296 (O_1296,N_24360,N_26445);
and UO_1297 (O_1297,N_26016,N_25651);
or UO_1298 (O_1298,N_25484,N_27214);
nand UO_1299 (O_1299,N_27431,N_24557);
and UO_1300 (O_1300,N_24555,N_24755);
or UO_1301 (O_1301,N_29824,N_24528);
nand UO_1302 (O_1302,N_27421,N_24613);
nor UO_1303 (O_1303,N_28466,N_25029);
or UO_1304 (O_1304,N_27210,N_26055);
nor UO_1305 (O_1305,N_25216,N_25158);
or UO_1306 (O_1306,N_28049,N_25492);
nor UO_1307 (O_1307,N_24085,N_26429);
xor UO_1308 (O_1308,N_28896,N_24018);
nor UO_1309 (O_1309,N_26222,N_29468);
or UO_1310 (O_1310,N_25892,N_27188);
or UO_1311 (O_1311,N_26519,N_28175);
xnor UO_1312 (O_1312,N_25062,N_26792);
or UO_1313 (O_1313,N_27547,N_25242);
and UO_1314 (O_1314,N_27410,N_27983);
nor UO_1315 (O_1315,N_27429,N_26920);
and UO_1316 (O_1316,N_24550,N_24261);
nand UO_1317 (O_1317,N_28924,N_24526);
and UO_1318 (O_1318,N_28513,N_26899);
or UO_1319 (O_1319,N_25913,N_27416);
nor UO_1320 (O_1320,N_26632,N_26863);
nor UO_1321 (O_1321,N_27493,N_28230);
nand UO_1322 (O_1322,N_24618,N_26784);
and UO_1323 (O_1323,N_24488,N_25034);
nor UO_1324 (O_1324,N_25344,N_26693);
or UO_1325 (O_1325,N_25827,N_24731);
nor UO_1326 (O_1326,N_27689,N_24271);
nor UO_1327 (O_1327,N_25700,N_26389);
nand UO_1328 (O_1328,N_26912,N_24477);
and UO_1329 (O_1329,N_28182,N_24029);
nand UO_1330 (O_1330,N_24377,N_25239);
and UO_1331 (O_1331,N_25807,N_25109);
nor UO_1332 (O_1332,N_27570,N_29702);
and UO_1333 (O_1333,N_27317,N_24681);
nor UO_1334 (O_1334,N_24505,N_26336);
and UO_1335 (O_1335,N_26523,N_27880);
or UO_1336 (O_1336,N_29258,N_29257);
nor UO_1337 (O_1337,N_24288,N_25280);
nand UO_1338 (O_1338,N_28935,N_28433);
nor UO_1339 (O_1339,N_28277,N_29367);
nand UO_1340 (O_1340,N_29952,N_25817);
xor UO_1341 (O_1341,N_29548,N_29890);
xnor UO_1342 (O_1342,N_29746,N_27667);
nand UO_1343 (O_1343,N_28467,N_27122);
nand UO_1344 (O_1344,N_25879,N_28884);
and UO_1345 (O_1345,N_27140,N_24260);
or UO_1346 (O_1346,N_27160,N_24499);
nor UO_1347 (O_1347,N_25900,N_25964);
nand UO_1348 (O_1348,N_24028,N_25127);
nor UO_1349 (O_1349,N_29208,N_28721);
nor UO_1350 (O_1350,N_25956,N_29207);
or UO_1351 (O_1351,N_27660,N_28400);
nor UO_1352 (O_1352,N_27213,N_26083);
nor UO_1353 (O_1353,N_24235,N_27791);
nor UO_1354 (O_1354,N_29862,N_29225);
or UO_1355 (O_1355,N_26896,N_28698);
and UO_1356 (O_1356,N_27035,N_28079);
nand UO_1357 (O_1357,N_26280,N_25511);
and UO_1358 (O_1358,N_29323,N_24065);
or UO_1359 (O_1359,N_24356,N_29478);
nand UO_1360 (O_1360,N_27637,N_25893);
or UO_1361 (O_1361,N_25864,N_24969);
nor UO_1362 (O_1362,N_27942,N_29031);
nand UO_1363 (O_1363,N_24746,N_27913);
or UO_1364 (O_1364,N_24576,N_27943);
and UO_1365 (O_1365,N_24868,N_28509);
and UO_1366 (O_1366,N_26583,N_27902);
nor UO_1367 (O_1367,N_24787,N_25529);
nor UO_1368 (O_1368,N_25142,N_27432);
nor UO_1369 (O_1369,N_25134,N_26475);
nand UO_1370 (O_1370,N_25638,N_25949);
nor UO_1371 (O_1371,N_25810,N_26724);
or UO_1372 (O_1372,N_28643,N_29326);
or UO_1373 (O_1373,N_25599,N_28494);
or UO_1374 (O_1374,N_26231,N_28125);
and UO_1375 (O_1375,N_24531,N_28425);
nor UO_1376 (O_1376,N_24032,N_28794);
nor UO_1377 (O_1377,N_29544,N_24726);
and UO_1378 (O_1378,N_27310,N_29891);
nor UO_1379 (O_1379,N_28880,N_26691);
nor UO_1380 (O_1380,N_28555,N_26645);
nand UO_1381 (O_1381,N_24275,N_27481);
xnor UO_1382 (O_1382,N_28037,N_25254);
xnor UO_1383 (O_1383,N_27591,N_29321);
xor UO_1384 (O_1384,N_25640,N_24925);
nor UO_1385 (O_1385,N_26470,N_27965);
and UO_1386 (O_1386,N_26644,N_26662);
or UO_1387 (O_1387,N_28071,N_24352);
and UO_1388 (O_1388,N_29170,N_26748);
nand UO_1389 (O_1389,N_24563,N_26609);
nand UO_1390 (O_1390,N_26344,N_28637);
nand UO_1391 (O_1391,N_26176,N_27759);
nor UO_1392 (O_1392,N_27692,N_25479);
nor UO_1393 (O_1393,N_26335,N_28038);
xnor UO_1394 (O_1394,N_25653,N_24775);
nand UO_1395 (O_1395,N_26086,N_29812);
nand UO_1396 (O_1396,N_24404,N_29909);
nand UO_1397 (O_1397,N_24456,N_26238);
nand UO_1398 (O_1398,N_24060,N_24323);
nor UO_1399 (O_1399,N_27021,N_24939);
nor UO_1400 (O_1400,N_24743,N_24533);
nor UO_1401 (O_1401,N_28190,N_27538);
and UO_1402 (O_1402,N_25833,N_28556);
xor UO_1403 (O_1403,N_29481,N_24790);
nand UO_1404 (O_1404,N_29332,N_29564);
or UO_1405 (O_1405,N_28439,N_29863);
nor UO_1406 (O_1406,N_26436,N_27772);
and UO_1407 (O_1407,N_29619,N_25038);
and UO_1408 (O_1408,N_29832,N_25973);
nand UO_1409 (O_1409,N_27119,N_28507);
nand UO_1410 (O_1410,N_25236,N_25244);
nor UO_1411 (O_1411,N_29200,N_27739);
nor UO_1412 (O_1412,N_25930,N_26440);
and UO_1413 (O_1413,N_25081,N_28329);
and UO_1414 (O_1414,N_27905,N_27607);
or UO_1415 (O_1415,N_28520,N_25197);
nor UO_1416 (O_1416,N_27799,N_25502);
and UO_1417 (O_1417,N_27300,N_28054);
nor UO_1418 (O_1418,N_28678,N_29828);
and UO_1419 (O_1419,N_24908,N_28461);
or UO_1420 (O_1420,N_25195,N_29670);
xor UO_1421 (O_1421,N_29012,N_27057);
and UO_1422 (O_1422,N_25983,N_29429);
or UO_1423 (O_1423,N_27868,N_29570);
xor UO_1424 (O_1424,N_26650,N_27211);
or UO_1425 (O_1425,N_24539,N_29038);
or UO_1426 (O_1426,N_25351,N_29886);
nand UO_1427 (O_1427,N_24617,N_27925);
or UO_1428 (O_1428,N_24370,N_24966);
nor UO_1429 (O_1429,N_26131,N_28661);
xor UO_1430 (O_1430,N_24996,N_24153);
nor UO_1431 (O_1431,N_27863,N_24932);
nand UO_1432 (O_1432,N_25724,N_26140);
or UO_1433 (O_1433,N_24749,N_24901);
and UO_1434 (O_1434,N_29349,N_29093);
or UO_1435 (O_1435,N_26040,N_26042);
nand UO_1436 (O_1436,N_25737,N_27768);
or UO_1437 (O_1437,N_29298,N_24284);
xnor UO_1438 (O_1438,N_24413,N_26095);
nor UO_1439 (O_1439,N_28261,N_29734);
and UO_1440 (O_1440,N_29690,N_28299);
nand UO_1441 (O_1441,N_28601,N_29695);
nor UO_1442 (O_1442,N_24314,N_26669);
nand UO_1443 (O_1443,N_26569,N_26012);
or UO_1444 (O_1444,N_25664,N_27800);
nor UO_1445 (O_1445,N_29006,N_29896);
nor UO_1446 (O_1446,N_28829,N_25284);
xnor UO_1447 (O_1447,N_26201,N_29210);
nor UO_1448 (O_1448,N_24353,N_29268);
nand UO_1449 (O_1449,N_26208,N_29978);
and UO_1450 (O_1450,N_26610,N_24705);
nor UO_1451 (O_1451,N_29204,N_24779);
or UO_1452 (O_1452,N_26367,N_29386);
xor UO_1453 (O_1453,N_25070,N_25355);
or UO_1454 (O_1454,N_28518,N_26568);
and UO_1455 (O_1455,N_26585,N_24734);
nand UO_1456 (O_1456,N_27926,N_27967);
nor UO_1457 (O_1457,N_26734,N_26381);
or UO_1458 (O_1458,N_24145,N_28422);
and UO_1459 (O_1459,N_26039,N_29580);
and UO_1460 (O_1460,N_24267,N_26253);
xnor UO_1461 (O_1461,N_27563,N_27235);
nand UO_1462 (O_1462,N_25035,N_28784);
or UO_1463 (O_1463,N_28042,N_26426);
nor UO_1464 (O_1464,N_25953,N_25896);
nand UO_1465 (O_1465,N_25578,N_26370);
nor UO_1466 (O_1466,N_27569,N_28296);
xor UO_1467 (O_1467,N_26641,N_24154);
and UO_1468 (O_1468,N_24081,N_27910);
or UO_1469 (O_1469,N_24162,N_26959);
or UO_1470 (O_1470,N_28972,N_24205);
nor UO_1471 (O_1471,N_27123,N_29662);
nor UO_1472 (O_1472,N_25016,N_26262);
or UO_1473 (O_1473,N_29798,N_29188);
nand UO_1474 (O_1474,N_28957,N_25844);
or UO_1475 (O_1475,N_29250,N_29785);
nor UO_1476 (O_1476,N_25226,N_26951);
nand UO_1477 (O_1477,N_25775,N_29649);
or UO_1478 (O_1478,N_25759,N_28087);
or UO_1479 (O_1479,N_26578,N_26273);
nand UO_1480 (O_1480,N_28697,N_26786);
and UO_1481 (O_1481,N_26973,N_27778);
nor UO_1482 (O_1482,N_26068,N_28341);
nand UO_1483 (O_1483,N_28975,N_24495);
nand UO_1484 (O_1484,N_26059,N_29142);
xnor UO_1485 (O_1485,N_28390,N_28352);
or UO_1486 (O_1486,N_27590,N_27494);
or UO_1487 (O_1487,N_25740,N_24830);
and UO_1488 (O_1488,N_26430,N_28928);
and UO_1489 (O_1489,N_26463,N_28405);
nand UO_1490 (O_1490,N_29002,N_28112);
nand UO_1491 (O_1491,N_28124,N_28511);
nand UO_1492 (O_1492,N_29904,N_25290);
nand UO_1493 (O_1493,N_24848,N_24820);
and UO_1494 (O_1494,N_25918,N_24662);
xor UO_1495 (O_1495,N_28484,N_24686);
nor UO_1496 (O_1496,N_24329,N_28274);
or UO_1497 (O_1497,N_29310,N_29541);
nor UO_1498 (O_1498,N_27080,N_28366);
or UO_1499 (O_1499,N_28890,N_27665);
nor UO_1500 (O_1500,N_27340,N_24795);
or UO_1501 (O_1501,N_29889,N_27092);
xor UO_1502 (O_1502,N_25083,N_29925);
nand UO_1503 (O_1503,N_25510,N_28155);
nor UO_1504 (O_1504,N_29777,N_28377);
and UO_1505 (O_1505,N_29899,N_29377);
nor UO_1506 (O_1506,N_28089,N_26874);
or UO_1507 (O_1507,N_25232,N_26617);
nand UO_1508 (O_1508,N_26424,N_26324);
nor UO_1509 (O_1509,N_26759,N_24562);
nor UO_1510 (O_1510,N_29965,N_25683);
xnor UO_1511 (O_1511,N_26654,N_29154);
nor UO_1512 (O_1512,N_29753,N_25268);
nand UO_1513 (O_1513,N_28883,N_25925);
nand UO_1514 (O_1514,N_24384,N_27610);
nand UO_1515 (O_1515,N_26477,N_26268);
nand UO_1516 (O_1516,N_28717,N_27237);
and UO_1517 (O_1517,N_24213,N_25734);
or UO_1518 (O_1518,N_29502,N_28560);
and UO_1519 (O_1519,N_29341,N_27857);
or UO_1520 (O_1520,N_27672,N_26985);
nand UO_1521 (O_1521,N_26251,N_25659);
nor UO_1522 (O_1522,N_26047,N_25106);
nor UO_1523 (O_1523,N_24822,N_27802);
nor UO_1524 (O_1524,N_26157,N_29192);
or UO_1525 (O_1525,N_26735,N_24469);
and UO_1526 (O_1526,N_27332,N_27118);
nand UO_1527 (O_1527,N_27978,N_24480);
nor UO_1528 (O_1528,N_28295,N_26741);
nand UO_1529 (O_1529,N_24447,N_24757);
nand UO_1530 (O_1530,N_25251,N_27360);
xor UO_1531 (O_1531,N_29894,N_27079);
nor UO_1532 (O_1532,N_27734,N_26772);
xor UO_1533 (O_1533,N_24737,N_26536);
and UO_1534 (O_1534,N_28464,N_24310);
nor UO_1535 (O_1535,N_29259,N_27349);
and UO_1536 (O_1536,N_28029,N_28823);
nand UO_1537 (O_1537,N_27058,N_24274);
or UO_1538 (O_1538,N_24283,N_24141);
nand UO_1539 (O_1539,N_24494,N_29887);
nand UO_1540 (O_1540,N_29589,N_28570);
and UO_1541 (O_1541,N_26455,N_25980);
and UO_1542 (O_1542,N_28233,N_25203);
and UO_1543 (O_1543,N_24893,N_29596);
xor UO_1544 (O_1544,N_25613,N_25860);
nand UO_1545 (O_1545,N_24151,N_25843);
nand UO_1546 (O_1546,N_29605,N_25104);
and UO_1547 (O_1547,N_26787,N_25008);
xor UO_1548 (O_1548,N_28253,N_24937);
or UO_1549 (O_1549,N_28091,N_25208);
nand UO_1550 (O_1550,N_28848,N_24246);
nand UO_1551 (O_1551,N_25123,N_24365);
nand UO_1552 (O_1552,N_25644,N_28893);
nand UO_1553 (O_1553,N_28825,N_27669);
and UO_1554 (O_1554,N_28270,N_24196);
nor UO_1555 (O_1555,N_27632,N_24672);
nand UO_1556 (O_1556,N_24545,N_25282);
nand UO_1557 (O_1557,N_26647,N_26701);
or UO_1558 (O_1558,N_27219,N_25929);
nand UO_1559 (O_1559,N_28294,N_24599);
nand UO_1560 (O_1560,N_25381,N_29080);
nor UO_1561 (O_1561,N_27008,N_25979);
nor UO_1562 (O_1562,N_24540,N_26525);
or UO_1563 (O_1563,N_25491,N_29507);
nor UO_1564 (O_1564,N_27128,N_24845);
nor UO_1565 (O_1565,N_27749,N_24936);
or UO_1566 (O_1566,N_29078,N_28255);
nor UO_1567 (O_1567,N_26161,N_24736);
xnor UO_1568 (O_1568,N_24772,N_27549);
nand UO_1569 (O_1569,N_29527,N_24127);
and UO_1570 (O_1570,N_26104,N_29281);
or UO_1571 (O_1571,N_24439,N_29847);
or UO_1572 (O_1572,N_28113,N_29522);
or UO_1573 (O_1573,N_28145,N_26551);
nand UO_1574 (O_1574,N_24312,N_26900);
nand UO_1575 (O_1575,N_28061,N_25315);
nand UO_1576 (O_1576,N_24647,N_29968);
nand UO_1577 (O_1577,N_27947,N_27635);
nand UO_1578 (O_1578,N_24185,N_29686);
or UO_1579 (O_1579,N_24635,N_25609);
and UO_1580 (O_1580,N_29021,N_24344);
or UO_1581 (O_1581,N_25171,N_25435);
and UO_1582 (O_1582,N_29945,N_29108);
nor UO_1583 (O_1583,N_28694,N_29838);
xor UO_1584 (O_1584,N_27316,N_29931);
nor UO_1585 (O_1585,N_25119,N_28703);
nor UO_1586 (O_1586,N_25398,N_24403);
nand UO_1587 (O_1587,N_29420,N_26257);
nor UO_1588 (O_1588,N_28966,N_25098);
nor UO_1589 (O_1589,N_24683,N_24780);
nor UO_1590 (O_1590,N_26673,N_25464);
nor UO_1591 (O_1591,N_25463,N_27202);
nand UO_1592 (O_1592,N_27220,N_25246);
nand UO_1593 (O_1593,N_26279,N_25845);
nand UO_1594 (O_1594,N_28048,N_25795);
nor UO_1595 (O_1595,N_24362,N_28282);
xor UO_1596 (O_1596,N_27175,N_28568);
nor UO_1597 (O_1597,N_28672,N_25164);
nand UO_1598 (O_1598,N_25015,N_26037);
nand UO_1599 (O_1599,N_28081,N_25798);
or UO_1600 (O_1600,N_26789,N_27670);
or UO_1601 (O_1601,N_29615,N_24090);
nor UO_1602 (O_1602,N_24388,N_24193);
nand UO_1603 (O_1603,N_26752,N_28914);
and UO_1604 (O_1604,N_26824,N_25412);
and UO_1605 (O_1605,N_24629,N_27201);
nand UO_1606 (O_1606,N_28631,N_26584);
nor UO_1607 (O_1607,N_27512,N_26849);
and UO_1608 (O_1608,N_24944,N_24024);
nor UO_1609 (O_1609,N_25132,N_25678);
and UO_1610 (O_1610,N_25269,N_25686);
or UO_1611 (O_1611,N_27394,N_24884);
nand UO_1612 (O_1612,N_27758,N_29239);
or UO_1613 (O_1613,N_24149,N_29599);
nor UO_1614 (O_1614,N_29238,N_25770);
or UO_1615 (O_1615,N_28806,N_26339);
nand UO_1616 (O_1616,N_24450,N_26261);
nor UO_1617 (O_1617,N_24771,N_26294);
nand UO_1618 (O_1618,N_28148,N_25155);
nor UO_1619 (O_1619,N_28266,N_24174);
and UO_1620 (O_1620,N_24682,N_25059);
xnor UO_1621 (O_1621,N_27120,N_25855);
nor UO_1622 (O_1622,N_29091,N_24270);
xor UO_1623 (O_1623,N_28843,N_25389);
and UO_1624 (O_1624,N_28769,N_29092);
or UO_1625 (O_1625,N_28945,N_24676);
or UO_1626 (O_1626,N_27168,N_25073);
nand UO_1627 (O_1627,N_26256,N_25139);
nor UO_1628 (O_1628,N_28051,N_26060);
or UO_1629 (O_1629,N_28151,N_27852);
xnor UO_1630 (O_1630,N_28290,N_29996);
nor UO_1631 (O_1631,N_28409,N_27740);
nor UO_1632 (O_1632,N_24070,N_29477);
nand UO_1633 (O_1633,N_25868,N_24123);
or UO_1634 (O_1634,N_24521,N_26530);
or UO_1635 (O_1635,N_25832,N_26886);
or UO_1636 (O_1636,N_26837,N_27200);
or UO_1637 (O_1637,N_27788,N_28323);
nand UO_1638 (O_1638,N_25096,N_27417);
and UO_1639 (O_1639,N_27241,N_24986);
nand UO_1640 (O_1640,N_29708,N_28735);
and UO_1641 (O_1641,N_29635,N_27952);
nor UO_1642 (O_1642,N_24842,N_26949);
nand UO_1643 (O_1643,N_26798,N_27911);
nand UO_1644 (O_1644,N_25725,N_27653);
or UO_1645 (O_1645,N_28985,N_24115);
and UO_1646 (O_1646,N_25637,N_27649);
nor UO_1647 (O_1647,N_26281,N_27997);
nand UO_1648 (O_1648,N_28350,N_27137);
and UO_1649 (O_1649,N_29969,N_25669);
nand UO_1650 (O_1650,N_27105,N_24865);
nand UO_1651 (O_1651,N_26416,N_24909);
and UO_1652 (O_1652,N_28180,N_25480);
nand UO_1653 (O_1653,N_28767,N_26363);
nand UO_1654 (O_1654,N_28724,N_24373);
or UO_1655 (O_1655,N_24302,N_27763);
or UO_1656 (O_1656,N_29650,N_27056);
and UO_1657 (O_1657,N_27020,N_29392);
nor UO_1658 (O_1658,N_27474,N_26080);
or UO_1659 (O_1659,N_24963,N_28482);
and UO_1660 (O_1660,N_27232,N_24849);
and UO_1661 (O_1661,N_26004,N_27530);
or UO_1662 (O_1662,N_25957,N_28188);
nand UO_1663 (O_1663,N_28055,N_26675);
nand UO_1664 (O_1664,N_25620,N_27339);
xnor UO_1665 (O_1665,N_24994,N_24295);
nor UO_1666 (O_1666,N_24679,N_26453);
nor UO_1667 (O_1667,N_28117,N_25726);
xnor UO_1668 (O_1668,N_25697,N_26166);
nor UO_1669 (O_1669,N_24802,N_25319);
nand UO_1670 (O_1670,N_28499,N_26547);
nor UO_1671 (O_1671,N_27600,N_24486);
nand UO_1672 (O_1672,N_26113,N_24815);
and UO_1673 (O_1673,N_27039,N_24347);
and UO_1674 (O_1674,N_25148,N_24105);
and UO_1675 (O_1675,N_29209,N_25305);
nand UO_1676 (O_1676,N_28337,N_29338);
or UO_1677 (O_1677,N_26747,N_25790);
and UO_1678 (O_1678,N_26407,N_28434);
nand UO_1679 (O_1679,N_24058,N_29424);
nor UO_1680 (O_1680,N_28068,N_25703);
and UO_1681 (O_1681,N_25185,N_24069);
or UO_1682 (O_1682,N_24215,N_24086);
nand UO_1683 (O_1683,N_26330,N_27475);
or UO_1684 (O_1684,N_27315,N_28693);
nor UO_1685 (O_1685,N_28288,N_29651);
nand UO_1686 (O_1686,N_26592,N_29826);
and UO_1687 (O_1687,N_26348,N_24051);
xor UO_1688 (O_1688,N_26433,N_26516);
and UO_1689 (O_1689,N_27064,N_26981);
or UO_1690 (O_1690,N_26540,N_25793);
nor UO_1691 (O_1691,N_29684,N_29441);
nor UO_1692 (O_1692,N_29404,N_29456);
and UO_1693 (O_1693,N_24375,N_28702);
or UO_1694 (O_1694,N_26828,N_25047);
or UO_1695 (O_1695,N_24692,N_28356);
nand UO_1696 (O_1696,N_26383,N_24855);
xnor UO_1697 (O_1697,N_25784,N_25729);
or UO_1698 (O_1698,N_28416,N_25014);
and UO_1699 (O_1699,N_27199,N_28242);
nor UO_1700 (O_1700,N_24173,N_29799);
xnor UO_1701 (O_1701,N_29317,N_26603);
and UO_1702 (O_1702,N_24229,N_28581);
and UO_1703 (O_1703,N_24886,N_27036);
and UO_1704 (O_1704,N_29322,N_27674);
and UO_1705 (O_1705,N_28712,N_24889);
nor UO_1706 (O_1706,N_28882,N_29479);
or UO_1707 (O_1707,N_28447,N_29506);
nand UO_1708 (O_1708,N_26855,N_24905);
and UO_1709 (O_1709,N_29732,N_26509);
and UO_1710 (O_1710,N_29353,N_26549);
xnor UO_1711 (O_1711,N_24473,N_29346);
nand UO_1712 (O_1712,N_28486,N_27981);
and UO_1713 (O_1713,N_24496,N_25854);
and UO_1714 (O_1714,N_25799,N_27026);
nand UO_1715 (O_1715,N_26827,N_27605);
and UO_1716 (O_1716,N_28524,N_28333);
nand UO_1717 (O_1717,N_24005,N_29701);
or UO_1718 (O_1718,N_29853,N_29422);
nor UO_1719 (O_1719,N_24809,N_24614);
or UO_1720 (O_1720,N_25250,N_27183);
xor UO_1721 (O_1721,N_25518,N_28320);
nand UO_1722 (O_1722,N_27083,N_28887);
or UO_1723 (O_1723,N_25175,N_24391);
nor UO_1724 (O_1724,N_24715,N_27989);
nand UO_1725 (O_1725,N_29607,N_29009);
and UO_1726 (O_1726,N_27506,N_25990);
or UO_1727 (O_1727,N_26034,N_26490);
or UO_1728 (O_1728,N_27645,N_25353);
nand UO_1729 (O_1729,N_24080,N_25406);
or UO_1730 (O_1730,N_25715,N_29157);
nor UO_1731 (O_1731,N_28628,N_28018);
or UO_1732 (O_1732,N_27190,N_25331);
nor UO_1733 (O_1733,N_28867,N_28859);
nor UO_1734 (O_1734,N_24803,N_26732);
nand UO_1735 (O_1735,N_29959,N_26796);
or UO_1736 (O_1736,N_24723,N_28901);
and UO_1737 (O_1737,N_29316,N_28013);
nand UO_1738 (O_1738,N_29348,N_28865);
or UO_1739 (O_1739,N_26801,N_28619);
xnor UO_1740 (O_1740,N_24813,N_25618);
or UO_1741 (O_1741,N_24227,N_24320);
nor UO_1742 (O_1742,N_26577,N_25709);
and UO_1743 (O_1743,N_24631,N_29169);
and UO_1744 (O_1744,N_29680,N_25273);
nand UO_1745 (O_1745,N_29999,N_26889);
and UO_1746 (O_1746,N_26065,N_27940);
nand UO_1747 (O_1747,N_24188,N_29878);
xnor UO_1748 (O_1748,N_24350,N_29767);
nor UO_1749 (O_1749,N_27193,N_28252);
nor UO_1750 (O_1750,N_28559,N_24034);
and UO_1751 (O_1751,N_29814,N_28202);
nor UO_1752 (O_1752,N_27258,N_24807);
nor UO_1753 (O_1753,N_28065,N_29227);
and UO_1754 (O_1754,N_25294,N_28271);
nor UO_1755 (O_1755,N_26579,N_25405);
or UO_1756 (O_1756,N_25552,N_24298);
nor UO_1757 (O_1757,N_29784,N_29846);
nor UO_1758 (O_1758,N_26028,N_29039);
or UO_1759 (O_1759,N_24245,N_25517);
nand UO_1760 (O_1760,N_27985,N_27873);
or UO_1761 (O_1761,N_28232,N_25911);
or UO_1762 (O_1762,N_26225,N_26484);
and UO_1763 (O_1763,N_26343,N_29175);
and UO_1764 (O_1764,N_26223,N_27142);
xnor UO_1765 (O_1765,N_26814,N_28777);
or UO_1766 (O_1766,N_26927,N_28459);
nor UO_1767 (O_1767,N_29627,N_27203);
and UO_1768 (O_1768,N_28306,N_25352);
and UO_1769 (O_1769,N_27189,N_26380);
nor UO_1770 (O_1770,N_25498,N_26563);
nand UO_1771 (O_1771,N_26295,N_28372);
xnor UO_1772 (O_1772,N_29810,N_27700);
and UO_1773 (O_1773,N_29736,N_25167);
or UO_1774 (O_1774,N_29487,N_25952);
or UO_1775 (O_1775,N_28481,N_28860);
nor UO_1776 (O_1776,N_25801,N_25229);
and UO_1777 (O_1777,N_28723,N_24325);
or UO_1778 (O_1778,N_25472,N_24445);
or UO_1779 (O_1779,N_26450,N_28036);
nor UO_1780 (O_1780,N_24667,N_28910);
nand UO_1781 (O_1781,N_27698,N_26145);
or UO_1782 (O_1782,N_28084,N_27482);
or UO_1783 (O_1783,N_25187,N_26093);
and UO_1784 (O_1784,N_25948,N_26272);
or UO_1785 (O_1785,N_25304,N_27721);
xnor UO_1786 (O_1786,N_25521,N_25228);
or UO_1787 (O_1787,N_27639,N_25004);
or UO_1788 (O_1788,N_29803,N_24256);
nand UO_1789 (O_1789,N_26621,N_27756);
xor UO_1790 (O_1790,N_25525,N_27679);
nor UO_1791 (O_1791,N_26757,N_29251);
or UO_1792 (O_1792,N_28072,N_27722);
and UO_1793 (O_1793,N_26135,N_28301);
and UO_1794 (O_1794,N_26233,N_28028);
and UO_1795 (O_1795,N_24633,N_25741);
or UO_1796 (O_1796,N_28963,N_25802);
xor UO_1797 (O_1797,N_24656,N_29845);
or UO_1798 (O_1798,N_24293,N_25147);
and UO_1799 (O_1799,N_29056,N_29226);
and UO_1800 (O_1800,N_26875,N_28264);
nand UO_1801 (O_1801,N_27369,N_27010);
or UO_1802 (O_1802,N_25575,N_27291);
xnor UO_1803 (O_1803,N_25804,N_24006);
nor UO_1804 (O_1804,N_24180,N_28454);
nor UO_1805 (O_1805,N_26209,N_27281);
and UO_1806 (O_1806,N_25436,N_24331);
or UO_1807 (O_1807,N_27247,N_29032);
or UO_1808 (O_1808,N_27054,N_25378);
or UO_1809 (O_1809,N_26755,N_29277);
and UO_1810 (O_1810,N_26762,N_28415);
or UO_1811 (O_1811,N_24888,N_26173);
and UO_1812 (O_1812,N_24869,N_29739);
or UO_1813 (O_1813,N_25082,N_29805);
nor UO_1814 (O_1814,N_27869,N_24394);
or UO_1815 (O_1815,N_26368,N_24014);
and UO_1816 (O_1816,N_26557,N_28237);
or UO_1817 (O_1817,N_27841,N_26740);
nand UO_1818 (O_1818,N_27415,N_29428);
nand UO_1819 (O_1819,N_26167,N_24998);
nand UO_1820 (O_1820,N_29146,N_28186);
or UO_1821 (O_1821,N_29249,N_26164);
or UO_1822 (O_1822,N_29774,N_27409);
xnor UO_1823 (O_1823,N_29760,N_24020);
nand UO_1824 (O_1824,N_29661,N_27825);
nor UO_1825 (O_1825,N_29754,N_26538);
and UO_1826 (O_1826,N_26485,N_29010);
or UO_1827 (O_1827,N_29370,N_24862);
or UO_1828 (O_1828,N_27462,N_29465);
and UO_1829 (O_1829,N_25670,N_27334);
or UO_1830 (O_1830,N_26211,N_26883);
and UO_1831 (O_1831,N_28667,N_26815);
nand UO_1832 (O_1832,N_25449,N_25933);
nand UO_1833 (O_1833,N_26637,N_27991);
and UO_1834 (O_1834,N_26546,N_29373);
or UO_1835 (O_1835,N_26375,N_25785);
or UO_1836 (O_1836,N_28281,N_25576);
or UO_1837 (O_1837,N_28211,N_25419);
or UO_1838 (O_1838,N_27025,N_29850);
or UO_1839 (O_1839,N_25339,N_24951);
nand UO_1840 (O_1840,N_29095,N_25370);
nor UO_1841 (O_1841,N_29879,N_25506);
nor UO_1842 (O_1842,N_24265,N_28775);
nor UO_1843 (O_1843,N_26117,N_27928);
nor UO_1844 (O_1844,N_29719,N_27814);
or UO_1845 (O_1845,N_24230,N_27423);
nor UO_1846 (O_1846,N_27769,N_24116);
nand UO_1847 (O_1847,N_29330,N_27994);
or UO_1848 (O_1848,N_29160,N_28060);
and UO_1849 (O_1849,N_24179,N_25050);
nand UO_1850 (O_1850,N_27623,N_28284);
xnor UO_1851 (O_1851,N_28410,N_26451);
nand UO_1852 (O_1852,N_28411,N_24678);
nor UO_1853 (O_1853,N_27618,N_27882);
and UO_1854 (O_1854,N_24276,N_24943);
xnor UO_1855 (O_1855,N_29617,N_27972);
and UO_1856 (O_1856,N_27053,N_29081);
or UO_1857 (O_1857,N_28933,N_29782);
xor UO_1858 (O_1858,N_29205,N_25581);
nand UO_1859 (O_1859,N_25340,N_27691);
or UO_1860 (O_1860,N_29740,N_25546);
xor UO_1861 (O_1861,N_27998,N_26587);
nand UO_1862 (O_1862,N_24111,N_24912);
or UO_1863 (O_1863,N_28379,N_24786);
nor UO_1864 (O_1864,N_26935,N_26175);
and UO_1865 (O_1865,N_24437,N_28980);
xnor UO_1866 (O_1866,N_24535,N_28816);
nor UO_1867 (O_1867,N_26064,N_25566);
nor UO_1868 (O_1868,N_26838,N_25000);
nor UO_1869 (O_1869,N_24799,N_24408);
xnor UO_1870 (O_1870,N_25885,N_28251);
nor UO_1871 (O_1871,N_24125,N_26193);
and UO_1872 (O_1872,N_25113,N_25543);
nand UO_1873 (O_1873,N_27113,N_24999);
or UO_1874 (O_1874,N_28196,N_24306);
nand UO_1875 (O_1875,N_28846,N_28622);
or UO_1876 (O_1876,N_27236,N_28383);
and UO_1877 (O_1877,N_26169,N_25349);
or UO_1878 (O_1878,N_24489,N_28708);
and UO_1879 (O_1879,N_25514,N_26834);
nor UO_1880 (O_1880,N_25611,N_25634);
nand UO_1881 (O_1881,N_25377,N_25665);
and UO_1882 (O_1882,N_27106,N_27320);
xnor UO_1883 (O_1883,N_27111,N_29378);
xor UO_1884 (O_1884,N_25606,N_25303);
nor UO_1885 (O_1885,N_27757,N_25421);
nor UO_1886 (O_1886,N_25907,N_28442);
nand UO_1887 (O_1887,N_28542,N_24992);
or UO_1888 (O_1888,N_27681,N_24409);
or UO_1889 (O_1889,N_27470,N_27602);
nor UO_1890 (O_1890,N_24451,N_28923);
and UO_1891 (O_1891,N_27899,N_29474);
or UO_1892 (O_1892,N_27592,N_29538);
nor UO_1893 (O_1893,N_29986,N_29956);
or UO_1894 (O_1894,N_24851,N_24475);
nand UO_1895 (O_1895,N_26387,N_29271);
and UO_1896 (O_1896,N_28384,N_25265);
and UO_1897 (O_1897,N_28854,N_25992);
or UO_1898 (O_1898,N_27979,N_26075);
and UO_1899 (O_1899,N_27625,N_25257);
and UO_1900 (O_1900,N_29575,N_27640);
and UO_1901 (O_1901,N_29622,N_28544);
nand UO_1902 (O_1902,N_29284,N_24198);
nand UO_1903 (O_1903,N_29953,N_29121);
nor UO_1904 (O_1904,N_29836,N_29800);
nand UO_1905 (O_1905,N_28670,N_27508);
nand UO_1906 (O_1906,N_27935,N_24371);
nand UO_1907 (O_1907,N_27684,N_26529);
nor UO_1908 (O_1908,N_26643,N_24637);
xor UO_1909 (O_1909,N_29313,N_29486);
nor UO_1910 (O_1910,N_24913,N_29713);
nor UO_1911 (O_1911,N_29397,N_29618);
nand UO_1912 (O_1912,N_26830,N_28584);
xor UO_1913 (O_1913,N_24770,N_25622);
xor UO_1914 (O_1914,N_29840,N_26338);
nor UO_1915 (O_1915,N_25209,N_25165);
and UO_1916 (O_1916,N_28875,N_26873);
or UO_1917 (O_1917,N_29632,N_29152);
nor UO_1918 (O_1918,N_29663,N_24751);
xnor UO_1919 (O_1919,N_24593,N_24330);
and UO_1920 (O_1920,N_28922,N_28381);
or UO_1921 (O_1921,N_27266,N_27061);
or UO_1922 (O_1922,N_25978,N_27327);
or UO_1923 (O_1923,N_26035,N_26685);
and UO_1924 (O_1924,N_26111,N_29408);
nand UO_1925 (O_1925,N_27909,N_29339);
xor UO_1926 (O_1926,N_26639,N_25789);
and UO_1927 (O_1927,N_29231,N_26738);
and UO_1928 (O_1928,N_24641,N_27944);
nand UO_1929 (O_1929,N_29628,N_25747);
and UO_1930 (O_1930,N_29405,N_29839);
nor UO_1931 (O_1931,N_28349,N_24182);
nor UO_1932 (O_1932,N_25888,N_27230);
nor UO_1933 (O_1933,N_26940,N_28267);
nand UO_1934 (O_1934,N_25602,N_27295);
xnor UO_1935 (O_1935,N_28837,N_27720);
nor UO_1936 (O_1936,N_29459,N_28200);
and UO_1937 (O_1937,N_27145,N_29778);
nor UO_1938 (O_1938,N_26373,N_29337);
or UO_1939 (O_1939,N_24147,N_28335);
nand UO_1940 (O_1940,N_29992,N_24379);
nand UO_1941 (O_1941,N_24652,N_29362);
or UO_1942 (O_1942,N_28572,N_26733);
xnor UO_1943 (O_1943,N_28490,N_24297);
or UO_1944 (O_1944,N_29094,N_25997);
nand UO_1945 (O_1945,N_26126,N_25275);
nand UO_1946 (O_1946,N_26965,N_29724);
nor UO_1947 (O_1947,N_26780,N_29556);
nand UO_1948 (O_1948,N_27068,N_26613);
or UO_1949 (O_1949,N_25730,N_27308);
nand UO_1950 (O_1950,N_29025,N_24170);
and UO_1951 (O_1951,N_28493,N_25519);
and UO_1952 (O_1952,N_29759,N_24881);
nand UO_1953 (O_1953,N_26642,N_24048);
nor UO_1954 (O_1954,N_28926,N_27716);
and UO_1955 (O_1955,N_27240,N_25143);
xnor UO_1956 (O_1956,N_25426,N_25027);
nor UO_1957 (O_1957,N_29664,N_25871);
and UO_1958 (O_1958,N_24124,N_28289);
xnor UO_1959 (O_1959,N_26214,N_28440);
and UO_1960 (O_1960,N_28414,N_27747);
and UO_1961 (O_1961,N_25093,N_28764);
nand UO_1962 (O_1962,N_29758,N_28364);
nor UO_1963 (O_1963,N_24991,N_24088);
or UO_1964 (O_1964,N_25975,N_24529);
nor UO_1965 (O_1965,N_26462,N_24166);
nand UO_1966 (O_1966,N_24195,N_25413);
or UO_1967 (O_1967,N_28979,N_28681);
xor UO_1968 (O_1968,N_27503,N_25327);
and UO_1969 (O_1969,N_26922,N_25431);
and UO_1970 (O_1970,N_28437,N_29997);
or UO_1971 (O_1971,N_25136,N_29673);
or UO_1972 (O_1972,N_25586,N_24554);
or UO_1973 (O_1973,N_26986,N_25116);
nand UO_1974 (O_1974,N_25188,N_25583);
nor UO_1975 (O_1975,N_27636,N_26488);
nor UO_1976 (O_1976,N_24903,N_24793);
and UO_1977 (O_1977,N_29023,N_26510);
nor UO_1978 (O_1978,N_24721,N_24561);
and UO_1979 (O_1979,N_28679,N_27810);
or UO_1980 (O_1980,N_26116,N_25078);
and UO_1981 (O_1981,N_25722,N_24522);
and UO_1982 (O_1982,N_26162,N_28427);
xnor UO_1983 (O_1983,N_25403,N_26325);
nor UO_1984 (O_1984,N_26947,N_29065);
nand UO_1985 (O_1985,N_28791,N_26241);
xor UO_1986 (O_1986,N_25809,N_26503);
xnor UO_1987 (O_1987,N_24010,N_29966);
xnor UO_1988 (O_1988,N_27562,N_26206);
and UO_1989 (O_1989,N_27853,N_25727);
or UO_1990 (O_1990,N_24673,N_29928);
or UO_1991 (O_1991,N_26802,N_27152);
or UO_1992 (O_1992,N_29008,N_24719);
or UO_1993 (O_1993,N_28218,N_26352);
nor UO_1994 (O_1994,N_26228,N_27782);
or UO_1995 (O_1995,N_24100,N_24067);
nand UO_1996 (O_1996,N_24931,N_29167);
nand UO_1997 (O_1997,N_29855,N_27809);
and UO_1998 (O_1998,N_24351,N_28527);
and UO_1999 (O_1999,N_28238,N_25625);
and UO_2000 (O_2000,N_27254,N_29320);
and UO_2001 (O_2001,N_26833,N_24286);
nor UO_2002 (O_2002,N_28436,N_29920);
and UO_2003 (O_2003,N_24542,N_24036);
or UO_2004 (O_2004,N_29344,N_28675);
nor UO_2005 (O_2005,N_26318,N_29692);
nand UO_2006 (O_2006,N_26953,N_27430);
and UO_2007 (O_2007,N_24328,N_26611);
and UO_2008 (O_2008,N_27040,N_29184);
nor UO_2009 (O_2009,N_27523,N_26250);
nor UO_2010 (O_2010,N_29851,N_24128);
xor UO_2011 (O_2011,N_28899,N_26252);
nand UO_2012 (O_2012,N_27816,N_27541);
nor UO_2013 (O_2013,N_28774,N_27966);
and UO_2014 (O_2014,N_28929,N_27553);
xor UO_2015 (O_2015,N_24044,N_27191);
nand UO_2016 (O_2016,N_27102,N_28408);
nand UO_2017 (O_2017,N_27849,N_28915);
or UO_2018 (O_2018,N_25516,N_28748);
nor UO_2019 (O_2019,N_26112,N_29072);
nor UO_2020 (O_2020,N_26767,N_29228);
nor UO_2021 (O_2021,N_28781,N_26316);
nand UO_2022 (O_2022,N_29371,N_24209);
nor UO_2023 (O_2023,N_29173,N_28317);
or UO_2024 (O_2024,N_26457,N_24008);
nor UO_2025 (O_2025,N_25190,N_24457);
xnor UO_2026 (O_2026,N_29524,N_29929);
nand UO_2027 (O_2027,N_28455,N_26152);
nor UO_2028 (O_2028,N_28248,N_26841);
and UO_2029 (O_2029,N_25556,N_26434);
or UO_2030 (O_2030,N_28564,N_24470);
or UO_2031 (O_2031,N_28719,N_25998);
nand UO_2032 (O_2032,N_26474,N_26465);
and UO_2033 (O_2033,N_26005,N_25912);
nor UO_2034 (O_2034,N_28353,N_25889);
nor UO_2035 (O_2035,N_29088,N_28189);
nand UO_2036 (O_2036,N_27348,N_24355);
nand UO_2037 (O_2037,N_25579,N_26963);
xnor UO_2038 (O_2038,N_27900,N_28210);
nand UO_2039 (O_2039,N_27399,N_26878);
nor UO_2040 (O_2040,N_24282,N_27407);
nand UO_2041 (O_2041,N_27276,N_24883);
nand UO_2042 (O_2042,N_25086,N_29825);
xor UO_2043 (O_2043,N_28451,N_29274);
nand UO_2044 (O_2044,N_27693,N_26172);
and UO_2045 (O_2045,N_26891,N_24181);
xnor UO_2046 (O_2046,N_28432,N_24923);
nand UO_2047 (O_2047,N_26498,N_29086);
and UO_2048 (O_2048,N_27787,N_25399);
nand UO_2049 (O_2049,N_24440,N_27023);
nor UO_2050 (O_2050,N_29813,N_24003);
or UO_2051 (O_2051,N_25539,N_27093);
nand UO_2052 (O_2052,N_28937,N_26684);
nand UO_2053 (O_2053,N_25842,N_26983);
nand UO_2054 (O_2054,N_27086,N_26655);
or UO_2055 (O_2055,N_25846,N_29036);
and UO_2056 (O_2056,N_24296,N_24947);
and UO_2057 (O_2057,N_26041,N_24693);
and UO_2058 (O_2058,N_25905,N_28143);
nand UO_2059 (O_2059,N_24132,N_26850);
nor UO_2060 (O_2060,N_28298,N_27283);
nand UO_2061 (O_2061,N_26558,N_27628);
or UO_2062 (O_2062,N_27984,N_25184);
nor UO_2063 (O_2063,N_29318,N_24708);
or UO_2064 (O_2064,N_26171,N_24481);
or UO_2065 (O_2065,N_29041,N_28762);
xor UO_2066 (O_2066,N_24204,N_27950);
nor UO_2067 (O_2067,N_29415,N_25060);
nor UO_2068 (O_2068,N_28351,N_29786);
and UO_2069 (O_2069,N_27518,N_28477);
nor UO_2070 (O_2070,N_25448,N_27917);
or UO_2071 (O_2071,N_26590,N_26581);
or UO_2072 (O_2072,N_26906,N_29519);
nand UO_2073 (O_2073,N_27425,N_26443);
nor UO_2074 (O_2074,N_29434,N_28012);
xor UO_2075 (O_2075,N_29560,N_24704);
nand UO_2076 (O_2076,N_26051,N_29820);
and UO_2077 (O_2077,N_27894,N_26106);
and UO_2078 (O_2078,N_25141,N_24464);
nand UO_2079 (O_2079,N_24839,N_24890);
nand UO_2080 (O_2080,N_25255,N_27804);
and UO_2081 (O_2081,N_29835,N_28030);
and UO_2082 (O_2082,N_27884,N_26357);
nor UO_2083 (O_2083,N_26676,N_28934);
and UO_2084 (O_2084,N_27398,N_29741);
or UO_2085 (O_2085,N_27922,N_26980);
and UO_2086 (O_2086,N_24368,N_28024);
nand UO_2087 (O_2087,N_29660,N_28506);
and UO_2088 (O_2088,N_25768,N_28577);
or UO_2089 (O_2089,N_29833,N_26315);
xor UO_2090 (O_2090,N_29770,N_24990);
nor UO_2091 (O_2091,N_25301,N_25095);
nor UO_2092 (O_2092,N_26631,N_29273);
nand UO_2093 (O_2093,N_26234,N_24327);
or UO_2094 (O_2094,N_28990,N_29115);
nand UO_2095 (O_2095,N_26139,N_25780);
and UO_2096 (O_2096,N_27206,N_24571);
nand UO_2097 (O_2097,N_27272,N_26307);
nand UO_2098 (O_2098,N_28236,N_28239);
nand UO_2099 (O_2099,N_24291,N_29141);
nand UO_2100 (O_2100,N_29135,N_29417);
nand UO_2101 (O_2101,N_27249,N_24938);
nor UO_2102 (O_2102,N_24448,N_24564);
nor UO_2103 (O_2103,N_28369,N_29747);
and UO_2104 (O_2104,N_29511,N_24022);
nor UO_2105 (O_2105,N_25476,N_28293);
and UO_2106 (O_2106,N_27180,N_25085);
nand UO_2107 (O_2107,N_24348,N_29934);
or UO_2108 (O_2108,N_26756,N_28553);
nor UO_2109 (O_2109,N_26276,N_24168);
and UO_2110 (O_2110,N_26851,N_25650);
xor UO_2111 (O_2111,N_25873,N_28003);
nand UO_2112 (O_2112,N_25931,N_25295);
or UO_2113 (O_2113,N_25174,N_28485);
or UO_2114 (O_2114,N_29536,N_28438);
nand UO_2115 (O_2115,N_25881,N_27157);
nand UO_2116 (O_2116,N_26995,N_25248);
nand UO_2117 (O_2117,N_27259,N_28234);
nor UO_2118 (O_2118,N_27099,N_26714);
and UO_2119 (O_2119,N_26264,N_24706);
nor UO_2120 (O_2120,N_25951,N_26205);
and UO_2121 (O_2121,N_28852,N_28212);
nor UO_2122 (O_2122,N_24804,N_24425);
or UO_2123 (O_2123,N_25850,N_29111);
xor UO_2124 (O_2124,N_29299,N_24144);
and UO_2125 (O_2125,N_29625,N_24474);
nand UO_2126 (O_2126,N_29954,N_27091);
xnor UO_2127 (O_2127,N_24740,N_27354);
and UO_2128 (O_2128,N_26934,N_26009);
nand UO_2129 (O_2129,N_26215,N_29049);
and UO_2130 (O_2130,N_27012,N_24685);
or UO_2131 (O_2131,N_29358,N_25976);
or UO_2132 (O_2132,N_26528,N_28058);
xnor UO_2133 (O_2133,N_29762,N_27238);
nand UO_2134 (O_2134,N_24337,N_26567);
or UO_2135 (O_2135,N_26456,N_24982);
nor UO_2136 (O_2136,N_24438,N_25533);
and UO_2137 (O_2137,N_24455,N_24303);
or UO_2138 (O_2138,N_26659,N_29294);
nand UO_2139 (O_2139,N_25826,N_24157);
or UO_2140 (O_2140,N_29640,N_29926);
nand UO_2141 (O_2141,N_27072,N_26379);
and UO_2142 (O_2142,N_28133,N_25691);
xor UO_2143 (O_2143,N_26192,N_26672);
xor UO_2144 (O_2144,N_29801,N_26868);
or UO_2145 (O_2145,N_24079,N_28707);
nand UO_2146 (O_2146,N_24017,N_25642);
nand UO_2147 (O_2147,N_24068,N_27761);
nand UO_2148 (O_2148,N_26870,N_28662);
and UO_2149 (O_2149,N_29218,N_24985);
nand UO_2150 (O_2150,N_28789,N_26725);
and UO_2151 (O_2151,N_26438,N_28359);
or UO_2152 (O_2152,N_26467,N_26313);
nand UO_2153 (O_2153,N_24101,N_28006);
xnor UO_2154 (O_2154,N_24113,N_27443);
or UO_2155 (O_2155,N_26966,N_24981);
nor UO_2156 (O_2156,N_29569,N_27927);
or UO_2157 (O_2157,N_25020,N_26526);
nor UO_2158 (O_2158,N_28479,N_29704);
and UO_2159 (O_2159,N_29457,N_29595);
xor UO_2160 (O_2160,N_25456,N_28959);
nand UO_2161 (O_2161,N_24547,N_25287);
nor UO_2162 (O_2162,N_26240,N_27121);
nand UO_2163 (O_2163,N_29491,N_25942);
nand UO_2164 (O_2164,N_27783,N_24383);
nand UO_2165 (O_2165,N_27019,N_25628);
and UO_2166 (O_2166,N_26624,N_27397);
or UO_2167 (O_2167,N_28082,N_26648);
nand UO_2168 (O_2168,N_29854,N_29165);
nand UO_2169 (O_2169,N_29843,N_25130);
xnor UO_2170 (O_2170,N_28450,N_28056);
xor UO_2171 (O_2171,N_27735,N_28642);
or UO_2172 (O_2172,N_26923,N_24608);
xor UO_2173 (O_2173,N_24828,N_24497);
and UO_2174 (O_2174,N_26439,N_26418);
or UO_2175 (O_2175,N_28502,N_29715);
and UO_2176 (O_2176,N_25943,N_24095);
xnor UO_2177 (O_2177,N_24970,N_25554);
or UO_2178 (O_2178,N_28137,N_27701);
or UO_2179 (O_2179,N_26989,N_26155);
and UO_2180 (O_2180,N_26894,N_28711);
and UO_2181 (O_2181,N_25938,N_26319);
and UO_2182 (O_2182,N_25373,N_25756);
nor UO_2183 (O_2183,N_28849,N_24169);
nor UO_2184 (O_2184,N_28665,N_26248);
nor UO_2185 (O_2185,N_27654,N_25486);
or UO_2186 (O_2186,N_29498,N_29947);
nand UO_2187 (O_2187,N_24364,N_25126);
nand UO_2188 (O_2188,N_24961,N_25131);
and UO_2189 (O_2189,N_27461,N_28393);
or UO_2190 (O_2190,N_28328,N_25343);
and UO_2191 (O_2191,N_25481,N_26478);
nand UO_2192 (O_2192,N_29985,N_28397);
and UO_2193 (O_2193,N_29295,N_25947);
nand UO_2194 (O_2194,N_28596,N_29809);
nor UO_2195 (O_2195,N_27336,N_28744);
or UO_2196 (O_2196,N_25361,N_26428);
nor UO_2197 (O_2197,N_25153,N_28062);
nand UO_2198 (O_2198,N_25384,N_29112);
or UO_2199 (O_2199,N_29118,N_25711);
nand UO_2200 (O_2200,N_25621,N_29869);
nor UO_2201 (O_2201,N_24050,N_27643);
xnor UO_2202 (O_2202,N_28191,N_28780);
and UO_2203 (O_2203,N_29267,N_25831);
nor UO_2204 (O_2204,N_26366,N_26990);
nand UO_2205 (O_2205,N_29473,N_27263);
or UO_2206 (O_2206,N_25205,N_25005);
or UO_2207 (O_2207,N_26278,N_26790);
nand UO_2208 (O_2208,N_29513,N_25551);
nand UO_2209 (O_2209,N_26712,N_27207);
nand UO_2210 (O_2210,N_24262,N_26275);
and UO_2211 (O_2211,N_24953,N_26993);
nor UO_2212 (O_2212,N_27159,N_27829);
nor UO_2213 (O_2213,N_25163,N_29396);
and UO_2214 (O_2214,N_26921,N_26700);
and UO_2215 (O_2215,N_28388,N_27709);
and UO_2216 (O_2216,N_28868,N_24407);
nor UO_2217 (O_2217,N_25291,N_26614);
and UO_2218 (O_2218,N_28655,N_25091);
nand UO_2219 (O_2219,N_26869,N_25504);
xnor UO_2220 (O_2220,N_24623,N_27158);
and UO_2221 (O_2221,N_26640,N_27767);
or UO_2222 (O_2222,N_25840,N_26217);
xnor UO_2223 (O_2223,N_28101,N_25689);
or UO_2224 (O_2224,N_24885,N_28976);
nand UO_2225 (O_2225,N_27801,N_24776);
nor UO_2226 (O_2226,N_25920,N_26807);
or UO_2227 (O_2227,N_28641,N_26014);
or UO_2228 (O_2228,N_28345,N_29939);
nand UO_2229 (O_2229,N_25857,N_27779);
nor UO_2230 (O_2230,N_27601,N_27434);
nor UO_2231 (O_2231,N_28169,N_25673);
nand UO_2232 (O_2232,N_25783,N_28798);
nand UO_2233 (O_2233,N_28750,N_26376);
xor UO_2234 (O_2234,N_27603,N_27245);
nor UO_2235 (O_2235,N_28862,N_27760);
and UO_2236 (O_2236,N_27217,N_27177);
nand UO_2237 (O_2237,N_24458,N_24380);
and UO_2238 (O_2238,N_25019,N_27181);
nor UO_2239 (O_2239,N_24919,N_24569);
and UO_2240 (O_2240,N_25598,N_24924);
or UO_2241 (O_2241,N_26520,N_27923);
nand UO_2242 (O_2242,N_29360,N_26555);
and UO_2243 (O_2243,N_25451,N_28608);
and UO_2244 (O_2244,N_24918,N_29646);
and UO_2245 (O_2245,N_28413,N_27322);
and UO_2246 (O_2246,N_25509,N_26124);
nand UO_2247 (O_2247,N_29756,N_27784);
and UO_2248 (O_2248,N_29444,N_27224);
nand UO_2249 (O_2249,N_29919,N_29600);
nand UO_2250 (O_2250,N_26702,N_28713);
nand UO_2251 (O_2251,N_25890,N_27995);
or UO_2252 (O_2252,N_27286,N_28032);
and UO_2253 (O_2253,N_26633,N_28522);
nand UO_2254 (O_2254,N_25668,N_29752);
nand UO_2255 (O_2255,N_25779,N_27471);
or UO_2256 (O_2256,N_28116,N_28224);
nand UO_2257 (O_2257,N_27278,N_28406);
and UO_2258 (O_2258,N_25218,N_26340);
nand UO_2259 (O_2259,N_29859,N_27555);
or UO_2260 (O_2260,N_28874,N_25917);
and UO_2261 (O_2261,N_28782,N_26397);
nand UO_2262 (O_2262,N_24435,N_24378);
or UO_2263 (O_2263,N_28921,N_25302);
or UO_2264 (O_2264,N_28361,N_28906);
and UO_2265 (O_2265,N_28908,N_25676);
and UO_2266 (O_2266,N_29829,N_24765);
xor UO_2267 (O_2267,N_27225,N_24559);
xnor UO_2268 (O_2268,N_28161,N_28904);
xnor UO_2269 (O_2269,N_24863,N_29504);
nor UO_2270 (O_2270,N_26342,N_28475);
nand UO_2271 (O_2271,N_26812,N_26354);
nand UO_2272 (O_2272,N_29552,N_27687);
and UO_2273 (O_2273,N_26067,N_26635);
nor UO_2274 (O_2274,N_27510,N_28726);
nor UO_2275 (O_2275,N_24012,N_28235);
nor UO_2276 (O_2276,N_28150,N_27813);
and UO_2277 (O_2277,N_27342,N_26596);
xnor UO_2278 (O_2278,N_29514,N_27307);
xnor UO_2279 (O_2279,N_25067,N_24376);
or UO_2280 (O_2280,N_25040,N_24630);
or UO_2281 (O_2281,N_25262,N_29531);
and UO_2282 (O_2282,N_25549,N_27848);
and UO_2283 (O_2283,N_26050,N_28313);
nor UO_2284 (O_2284,N_29848,N_29365);
nand UO_2285 (O_2285,N_26907,N_25428);
and UO_2286 (O_2286,N_27363,N_25537);
and UO_2287 (O_2287,N_28039,N_27741);
nor UO_2288 (O_2288,N_25427,N_29532);
nand UO_2289 (O_2289,N_29471,N_29102);
xnor UO_2290 (O_2290,N_27815,N_28828);
or UO_2291 (O_2291,N_24989,N_24415);
or UO_2292 (O_2292,N_24709,N_24429);
xor UO_2293 (O_2293,N_27505,N_25847);
or UO_2294 (O_2294,N_29016,N_25493);
and UO_2295 (O_2295,N_27865,N_24176);
nand UO_2296 (O_2296,N_29262,N_26758);
nand UO_2297 (O_2297,N_25387,N_24952);
or UO_2298 (O_2298,N_24640,N_29566);
or UO_2299 (O_2299,N_29503,N_26765);
or UO_2300 (O_2300,N_25234,N_27656);
nor UO_2301 (O_2301,N_25058,N_26146);
nand UO_2302 (O_2302,N_26507,N_29090);
nand UO_2303 (O_2303,N_26768,N_29620);
nand UO_2304 (O_2304,N_24847,N_27293);
and UO_2305 (O_2305,N_26615,N_29145);
nand UO_2306 (O_2306,N_28243,N_28571);
nand UO_2307 (O_2307,N_25094,N_24718);
and UO_2308 (O_2308,N_28747,N_24078);
and UO_2309 (O_2309,N_28480,N_28491);
or UO_2310 (O_2310,N_24914,N_29906);
nand UO_2311 (O_2311,N_28096,N_24165);
or UO_2312 (O_2312,N_24035,N_25569);
nor UO_2313 (O_2313,N_27059,N_24392);
or UO_2314 (O_2314,N_24530,N_24609);
nand UO_2315 (O_2315,N_26236,N_27368);
xor UO_2316 (O_2316,N_25538,N_28269);
nor UO_2317 (O_2317,N_29237,N_27499);
nor UO_2318 (O_2318,N_26720,N_27987);
nand UO_2319 (O_2319,N_25430,N_27185);
xor UO_2320 (O_2320,N_28206,N_29450);
or UO_2321 (O_2321,N_28760,N_29868);
and UO_2322 (O_2322,N_27347,N_29148);
or UO_2323 (O_2323,N_29069,N_26320);
and UO_2324 (O_2324,N_27147,N_29430);
nor UO_2325 (O_2325,N_29410,N_27458);
or UO_2326 (O_2326,N_27854,N_25753);
and UO_2327 (O_2327,N_26151,N_26032);
nor UO_2328 (O_2328,N_28961,N_28370);
or UO_2329 (O_2329,N_24177,N_27418);
nor UO_2330 (O_2330,N_25418,N_26013);
xnor UO_2331 (O_2331,N_24089,N_29750);
nor UO_2332 (O_2332,N_28737,N_27205);
or UO_2333 (O_2333,N_27289,N_26847);
nand UO_2334 (O_2334,N_27949,N_25266);
and UO_2335 (O_2335,N_28898,N_24369);
or UO_2336 (O_2336,N_26502,N_29132);
nand UO_2337 (O_2337,N_24968,N_26799);
or UO_2338 (O_2338,N_25441,N_25596);
nor UO_2339 (O_2339,N_24720,N_29745);
nor UO_2340 (O_2340,N_29014,N_24340);
nand UO_2341 (O_2341,N_29681,N_25666);
nand UO_2342 (O_2342,N_27837,N_28680);
nand UO_2343 (O_2343,N_25772,N_28374);
and UO_2344 (O_2344,N_28905,N_24671);
or UO_2345 (O_2345,N_26695,N_25858);
nand UO_2346 (O_2346,N_29128,N_26464);
nand UO_2347 (O_2347,N_27641,N_25837);
xnor UO_2348 (O_2348,N_27271,N_28795);
nor UO_2349 (O_2349,N_26998,N_26881);
and UO_2350 (O_2350,N_25841,N_27492);
or UO_2351 (O_2351,N_27196,N_28504);
xor UO_2352 (O_2352,N_28615,N_24511);
nor UO_2353 (O_2353,N_26084,N_28648);
nand UO_2354 (O_2354,N_24874,N_26888);
nor UO_2355 (O_2355,N_25125,N_29987);
and UO_2356 (O_2356,N_27435,N_24611);
and UO_2357 (O_2357,N_26141,N_26400);
nor UO_2358 (O_2358,N_25915,N_25372);
and UO_2359 (O_2359,N_28503,N_27209);
nand UO_2360 (O_2360,N_24301,N_25452);
xnor UO_2361 (O_2361,N_27306,N_27710);
or UO_2362 (O_2362,N_24074,N_26496);
nand UO_2363 (O_2363,N_25152,N_25965);
xor UO_2364 (O_2364,N_29639,N_27956);
nand UO_2365 (O_2365,N_26594,N_28172);
and UO_2366 (O_2366,N_28844,N_29003);
nand UO_2367 (O_2367,N_29659,N_29722);
nand UO_2368 (O_2368,N_29071,N_27936);
nor UO_2369 (O_2369,N_25181,N_25074);
or UO_2370 (O_2370,N_26165,N_24119);
or UO_2371 (O_2371,N_27298,N_24962);
nor UO_2372 (O_2372,N_27973,N_29017);
and UO_2373 (O_2373,N_28808,N_29335);
and UO_2374 (O_2374,N_25541,N_24523);
and UO_2375 (O_2375,N_29296,N_24108);
and UO_2376 (O_2376,N_26508,N_28094);
xor UO_2377 (O_2377,N_24160,N_24823);
and UO_2378 (O_2378,N_27630,N_27939);
nor UO_2379 (O_2379,N_24950,N_24651);
xor UO_2380 (O_2380,N_24774,N_25762);
or UO_2381 (O_2381,N_25805,N_24483);
and UO_2382 (O_2382,N_29796,N_25371);
and UO_2383 (O_2383,N_27893,N_28588);
xor UO_2384 (O_2384,N_27834,N_29074);
or UO_2385 (O_2385,N_25066,N_28198);
xor UO_2386 (O_2386,N_28168,N_27504);
nor UO_2387 (O_2387,N_25264,N_25654);
xor UO_2388 (O_2388,N_25720,N_27671);
or UO_2389 (O_2389,N_29312,N_29189);
nor UO_2390 (O_2390,N_29913,N_25764);
or UO_2391 (O_2391,N_24131,N_29356);
or UO_2392 (O_2392,N_29901,N_27514);
and UO_2393 (O_2393,N_25233,N_24887);
nor UO_2394 (O_2394,N_29000,N_24699);
nor UO_2395 (O_2395,N_24722,N_29606);
or UO_2396 (O_2396,N_29076,N_28900);
and UO_2397 (O_2397,N_25630,N_29636);
or UO_2398 (O_2398,N_24133,N_25258);
xor UO_2399 (O_2399,N_28160,N_27702);
nor UO_2400 (O_2400,N_28309,N_24844);
nor UO_2401 (O_2401,N_25698,N_28583);
nor UO_2402 (O_2402,N_25710,N_28250);
xor UO_2403 (O_2403,N_26114,N_25610);
or UO_2404 (O_2404,N_24479,N_27892);
xor UO_2405 (O_2405,N_25643,N_28736);
nor UO_2406 (O_2406,N_27155,N_25380);
nor UO_2407 (O_2407,N_24579,N_24546);
or UO_2408 (O_2408,N_27571,N_28417);
and UO_2409 (O_2409,N_24414,N_27324);
nor UO_2410 (O_2410,N_29561,N_26148);
or UO_2411 (O_2411,N_27304,N_29938);
or UO_2412 (O_2412,N_27264,N_27239);
nor UO_2413 (O_2413,N_27543,N_29979);
nand UO_2414 (O_2414,N_26719,N_29881);
or UO_2415 (O_2415,N_24954,N_29436);
and UO_2416 (O_2416,N_27096,N_29980);
xor UO_2417 (O_2417,N_29748,N_26674);
and UO_2418 (O_2418,N_26081,N_27163);
and UO_2419 (O_2419,N_24063,N_29155);
nor UO_2420 (O_2420,N_26115,N_28788);
and UO_2421 (O_2421,N_28947,N_24871);
or UO_2422 (O_2422,N_28733,N_25761);
nand UO_2423 (O_2423,N_24203,N_25966);
nor UO_2424 (O_2424,N_27866,N_27650);
nand UO_2425 (O_2425,N_25223,N_26461);
or UO_2426 (O_2426,N_24860,N_26901);
and UO_2427 (O_2427,N_26717,N_29179);
and UO_2428 (O_2428,N_24420,N_25520);
and UO_2429 (O_2429,N_27000,N_26469);
and UO_2430 (O_2430,N_27725,N_29521);
nor UO_2431 (O_2431,N_28759,N_28435);
or UO_2432 (O_2432,N_27326,N_25507);
nor UO_2433 (O_2433,N_29248,N_29066);
nand UO_2434 (O_2434,N_26213,N_25880);
nor UO_2435 (O_2435,N_24363,N_25166);
and UO_2436 (O_2436,N_27489,N_28617);
and UO_2437 (O_2437,N_27301,N_26774);
or UO_2438 (O_2438,N_29211,N_27683);
nand UO_2439 (O_2439,N_26224,N_25259);
or UO_2440 (O_2440,N_28918,N_24567);
nand UO_2441 (O_2441,N_27052,N_29347);
xor UO_2442 (O_2442,N_25071,N_28468);
xor UO_2443 (O_2443,N_29213,N_27921);
nand UO_2444 (O_2444,N_29903,N_27585);
and UO_2445 (O_2445,N_27089,N_26775);
nand UO_2446 (O_2446,N_29669,N_25458);
and UO_2447 (O_2447,N_27557,N_24553);
nand UO_2448 (O_2448,N_29501,N_26879);
or UO_2449 (O_2449,N_28228,N_25988);
or UO_2450 (O_2450,N_26048,N_27982);
or UO_2451 (O_2451,N_26127,N_24294);
xor UO_2452 (O_2452,N_28879,N_28827);
nor UO_2453 (O_2453,N_25227,N_29240);
nand UO_2454 (O_2454,N_24013,N_29610);
or UO_2455 (O_2455,N_25364,N_26003);
and UO_2456 (O_2456,N_29101,N_29764);
or UO_2457 (O_2457,N_24764,N_28153);
and UO_2458 (O_2458,N_24891,N_27454);
and UO_2459 (O_2459,N_26677,N_24444);
and UO_2460 (O_2460,N_28863,N_24549);
and UO_2461 (O_2461,N_24834,N_29171);
or UO_2462 (O_2462,N_28249,N_29308);
nor UO_2463 (O_2463,N_29001,N_28938);
or UO_2464 (O_2464,N_25712,N_25916);
nand UO_2465 (O_2465,N_27438,N_27265);
and UO_2466 (O_2466,N_27246,N_29508);
xor UO_2467 (O_2467,N_26661,N_27375);
or UO_2468 (O_2468,N_28986,N_27478);
xor UO_2469 (O_2469,N_26636,N_27243);
or UO_2470 (O_2470,N_26630,N_24532);
or UO_2471 (O_2471,N_28872,N_28700);
nor UO_2472 (O_2472,N_27223,N_27178);
nor UO_2473 (O_2473,N_28194,N_29768);
nor UO_2474 (O_2474,N_29050,N_29976);
and UO_2475 (O_2475,N_29557,N_29616);
nand UO_2476 (O_2476,N_27268,N_25409);
nand UO_2477 (O_2477,N_26293,N_29733);
and UO_2478 (O_2478,N_27279,N_24955);
nand UO_2479 (O_2479,N_28977,N_24411);
and UO_2480 (O_2480,N_26803,N_29598);
and UO_2481 (O_2481,N_27311,N_26769);
and UO_2482 (O_2482,N_25100,N_27323);
xor UO_2483 (O_2483,N_29163,N_25211);
nor UO_2484 (O_2484,N_24308,N_24046);
nand UO_2485 (O_2485,N_28035,N_29699);
and UO_2486 (O_2486,N_28362,N_28894);
or UO_2487 (O_2487,N_27179,N_24178);
xnor UO_2488 (O_2488,N_24073,N_25105);
nor UO_2489 (O_2489,N_24207,N_29161);
nor UO_2490 (O_2490,N_29830,N_24922);
nand UO_2491 (O_2491,N_24287,N_25423);
nand UO_2492 (O_2492,N_28888,N_26542);
and UO_2493 (O_2493,N_26606,N_27742);
nor UO_2494 (O_2494,N_28146,N_26686);
nor UO_2495 (O_2495,N_26120,N_29703);
xnor UO_2496 (O_2496,N_29512,N_29247);
nor UO_2497 (O_2497,N_27598,N_24846);
or UO_2498 (O_2498,N_29608,N_28552);
xor UO_2499 (O_2499,N_24502,N_29485);
and UO_2500 (O_2500,N_28216,N_28858);
xnor UO_2501 (O_2501,N_25906,N_25178);
nor UO_2502 (O_2502,N_24210,N_29236);
xor UO_2503 (O_2503,N_27775,N_24254);
or UO_2504 (O_2504,N_28319,N_24247);
nand UO_2505 (O_2505,N_25240,N_24983);
nand UO_2506 (O_2506,N_28688,N_24037);
nor UO_2507 (O_2507,N_28223,N_28404);
and UO_2508 (O_2508,N_25077,N_28347);
and UO_2509 (O_2509,N_27885,N_28192);
nor UO_2510 (O_2510,N_24485,N_25482);
and UO_2511 (O_2511,N_27974,N_24031);
nor UO_2512 (O_2512,N_24516,N_24118);
xnor UO_2513 (O_2513,N_28152,N_28495);
nor UO_2514 (O_2514,N_29217,N_28179);
nand UO_2515 (O_2515,N_27517,N_24015);
and UO_2516 (O_2516,N_28573,N_28007);
and UO_2517 (O_2517,N_25749,N_25941);
nor UO_2518 (O_2518,N_26797,N_29272);
and UO_2519 (O_2519,N_24461,N_29222);
nand UO_2520 (O_2520,N_26216,N_27574);
nand UO_2521 (O_2521,N_24538,N_28996);
or UO_2522 (O_2522,N_29048,N_25777);
nand UO_2523 (O_2523,N_28312,N_25385);
nand UO_2524 (O_2524,N_24231,N_25277);
or UO_2525 (O_2525,N_27818,N_24895);
or UO_2526 (O_2526,N_27413,N_28690);
or UO_2527 (O_2527,N_25776,N_24512);
nor UO_2528 (O_2528,N_29685,N_28385);
or UO_2529 (O_2529,N_29539,N_28714);
nand UO_2530 (O_2530,N_27793,N_25365);
nor UO_2531 (O_2531,N_26235,N_27270);
xnor UO_2532 (O_2532,N_24402,N_24441);
nor UO_2533 (O_2533,N_28470,N_28960);
nor UO_2534 (O_2534,N_27457,N_27114);
nor UO_2535 (O_2535,N_26608,N_26537);
nor UO_2536 (O_2536,N_27992,N_27794);
or UO_2537 (O_2537,N_29790,N_25026);
nor UO_2538 (O_2538,N_24760,N_27024);
nor UO_2539 (O_2539,N_24335,N_24979);
or UO_2540 (O_2540,N_26723,N_27642);
and UO_2541 (O_2541,N_27620,N_25099);
xor UO_2542 (O_2542,N_24798,N_24821);
nand UO_2543 (O_2543,N_28818,N_28375);
nand UO_2544 (O_2544,N_27836,N_25145);
or UO_2545 (O_2545,N_28371,N_25573);
xnor UO_2546 (O_2546,N_24194,N_29611);
and UO_2547 (O_2547,N_29275,N_24735);
xor UO_2548 (O_2548,N_28786,N_25750);
nor UO_2549 (O_2549,N_26184,N_29626);
nor UO_2550 (O_2550,N_24907,N_29493);
or UO_2551 (O_2551,N_25437,N_27367);
and UO_2552 (O_2552,N_26618,N_26777);
nor UO_2553 (O_2553,N_25107,N_27134);
nor UO_2554 (O_2554,N_26306,N_25897);
and UO_2555 (O_2555,N_25813,N_29614);
nor UO_2556 (O_2556,N_26311,N_29126);
xnor UO_2557 (O_2557,N_24840,N_28616);
and UO_2558 (O_2558,N_25293,N_25894);
and UO_2559 (O_2559,N_26309,N_24412);
and UO_2560 (O_2560,N_29399,N_27042);
or UO_2561 (O_2561,N_25337,N_24534);
nor UO_2562 (O_2562,N_28776,N_27182);
nand UO_2563 (O_2563,N_24759,N_29988);
nor UO_2564 (O_2564,N_28444,N_25112);
xnor UO_2565 (O_2565,N_29950,N_24836);
or UO_2566 (O_2566,N_29120,N_29350);
or UO_2567 (O_2567,N_24621,N_25362);
or UO_2568 (O_2568,N_24778,N_26495);
xor UO_2569 (O_2569,N_26860,N_27087);
nand UO_2570 (O_2570,N_27516,N_26033);
nor UO_2571 (O_2571,N_26918,N_24677);
nor UO_2572 (O_2572,N_27958,N_26848);
or UO_2573 (O_2573,N_27916,N_25470);
or UO_2574 (O_2574,N_26448,N_27343);
and UO_2575 (O_2575,N_28159,N_26118);
nor UO_2576 (O_2576,N_25773,N_27907);
nor UO_2577 (O_2577,N_28903,N_29442);
and UO_2578 (O_2578,N_28598,N_27552);
xor UO_2579 (O_2579,N_29908,N_29147);
nor UO_2580 (O_2580,N_25260,N_27204);
and UO_2581 (O_2581,N_26326,N_25386);
nor UO_2582 (O_2582,N_27732,N_24756);
nor UO_2583 (O_2583,N_27028,N_24698);
nand UO_2584 (O_2584,N_25114,N_24728);
nor UO_2585 (O_2585,N_25882,N_29967);
xor UO_2586 (O_2586,N_25928,N_29390);
or UO_2587 (O_2587,N_24707,N_28948);
and UO_2588 (O_2588,N_26871,N_27257);
nand UO_2589 (O_2589,N_27014,N_29765);
xnor UO_2590 (O_2590,N_26494,N_25311);
or UO_2591 (O_2591,N_29461,N_29728);
and UO_2592 (O_2592,N_24714,N_29077);
and UO_2593 (O_2593,N_24056,N_28093);
nand UO_2594 (O_2594,N_25400,N_27156);
or UO_2595 (O_2595,N_25459,N_24717);
nand UO_2596 (O_2596,N_25151,N_25958);
and UO_2597 (O_2597,N_28998,N_27465);
nor UO_2598 (O_2598,N_28166,N_29293);
or UO_2599 (O_2599,N_27146,N_27074);
nor UO_2600 (O_2600,N_29933,N_28802);
nand UO_2601 (O_2601,N_24797,N_24945);
nand UO_2602 (O_2602,N_27781,N_24315);
nor UO_2603 (O_2603,N_26107,N_25135);
nor UO_2604 (O_2604,N_29542,N_25987);
xnor UO_2605 (O_2605,N_25557,N_25945);
nand UO_2606 (O_2606,N_29518,N_26778);
nand UO_2607 (O_2607,N_26668,N_28630);
nor UO_2608 (O_2608,N_29045,N_25468);
or UO_2609 (O_2609,N_27872,N_24163);
or UO_2610 (O_2610,N_26713,N_28208);
nand UO_2611 (O_2611,N_27509,N_25796);
nand UO_2612 (O_2612,N_29124,N_25478);
nand UO_2613 (O_2613,N_29873,N_26263);
nand UO_2614 (O_2614,N_27614,N_27132);
and UO_2615 (O_2615,N_26198,N_24300);
xor UO_2616 (O_2616,N_29263,N_28768);
nand UO_2617 (O_2617,N_27842,N_26588);
and UO_2618 (O_2618,N_25685,N_28911);
and UO_2619 (O_2619,N_28334,N_24984);
nand UO_2620 (O_2620,N_24902,N_25030);
xnor UO_2621 (O_2621,N_26328,N_28551);
nor UO_2622 (O_2622,N_26628,N_24600);
nor UO_2623 (O_2623,N_27404,N_26867);
nand UO_2624 (O_2624,N_25699,N_26687);
nand UO_2625 (O_2625,N_28639,N_25898);
or UO_2626 (O_2626,N_28074,N_27840);
or UO_2627 (O_2627,N_29837,N_27754);
nand UO_2628 (O_2628,N_27125,N_26539);
and UO_2629 (O_2629,N_26928,N_26788);
or UO_2630 (O_2630,N_28380,N_27198);
or UO_2631 (O_2631,N_28792,N_24033);
and UO_2632 (O_2632,N_26753,N_25558);
or UO_2633 (O_2633,N_28625,N_29683);
and UO_2634 (O_2634,N_25028,N_29172);
and UO_2635 (O_2635,N_28597,N_24620);
and UO_2636 (O_2636,N_26408,N_27480);
nand UO_2637 (O_2637,N_25330,N_27228);
xnor UO_2638 (O_2638,N_24570,N_27545);
and UO_2639 (O_2639,N_25168,N_24172);
nand UO_2640 (O_2640,N_26058,N_29288);
nand UO_2641 (O_2641,N_29911,N_29359);
and UO_2642 (O_2642,N_26909,N_29054);
and UO_2643 (O_2643,N_26904,N_24138);
nand UO_2644 (O_2644,N_25324,N_29414);
nand UO_2645 (O_2645,N_25736,N_26997);
or UO_2646 (O_2646,N_29711,N_25559);
and UO_2647 (O_2647,N_28478,N_25963);
nand UO_2648 (O_2648,N_28718,N_27646);
nand UO_2649 (O_2649,N_29035,N_28219);
and UO_2650 (O_2650,N_26053,N_25270);
xor UO_2651 (O_2651,N_26030,N_24785);
nand UO_2652 (O_2652,N_29902,N_26341);
nand UO_2653 (O_2653,N_29412,N_29586);
xnor UO_2654 (O_2654,N_25249,N_29533);
xnor UO_2655 (O_2655,N_26158,N_24866);
or UO_2656 (O_2656,N_26301,N_27446);
nand UO_2657 (O_2657,N_28021,N_25742);
or UO_2658 (O_2658,N_29941,N_29266);
and UO_2659 (O_2659,N_29265,N_28543);
and UO_2660 (O_2660,N_28332,N_26730);
and UO_2661 (O_2661,N_26359,N_26999);
nand UO_2662 (O_2662,N_29232,N_26969);
nand UO_2663 (O_2663,N_25306,N_24688);
and UO_2664 (O_2664,N_25501,N_26196);
or UO_2665 (O_2665,N_24004,N_27256);
or UO_2666 (O_2666,N_27328,N_27951);
nand UO_2667 (O_2667,N_24487,N_29384);
nor UO_2668 (O_2668,N_24307,N_25154);
nor UO_2669 (O_2669,N_27690,N_27150);
nor UO_2670 (O_2670,N_29718,N_28510);
nor UO_2671 (O_2671,N_27529,N_28020);
and UO_2672 (O_2672,N_29515,N_26125);
and UO_2673 (O_2673,N_27808,N_28997);
or UO_2674 (O_2674,N_26954,N_27082);
nand UO_2675 (O_2675,N_27318,N_26962);
nand UO_2676 (O_2676,N_27085,N_28856);
and UO_2677 (O_2677,N_27608,N_29841);
or UO_2678 (O_2678,N_25317,N_29221);
and UO_2679 (O_2679,N_27303,N_24589);
nor UO_2680 (O_2680,N_28009,N_26472);
nand UO_2681 (O_2681,N_29283,N_24349);
or UO_2682 (O_2682,N_27485,N_27090);
and UO_2683 (O_2683,N_25954,N_26078);
and UO_2684 (O_2684,N_27166,N_24156);
and UO_2685 (O_2685,N_25977,N_27901);
and UO_2686 (O_2686,N_27558,N_24768);
nand UO_2687 (O_2687,N_25256,N_28348);
and UO_2688 (O_2688,N_26302,N_25984);
xnor UO_2689 (O_2689,N_25908,N_24980);
nand UO_2690 (O_2690,N_25822,N_25513);
xor UO_2691 (O_2691,N_26781,N_24827);
or UO_2692 (O_2692,N_27288,N_25359);
nor UO_2693 (O_2693,N_24831,N_27736);
nor UO_2694 (O_2694,N_26800,N_26298);
and UO_2695 (O_2695,N_25607,N_29100);
xnor UO_2696 (O_2696,N_29970,N_28895);
or UO_2697 (O_2697,N_26395,N_27718);
and UO_2698 (O_2698,N_25835,N_29781);
or UO_2699 (O_2699,N_24019,N_25627);
and UO_2700 (O_2700,N_27077,N_27098);
xor UO_2701 (O_2701,N_24597,N_26895);
and UO_2702 (O_2702,N_26729,N_26287);
and UO_2703 (O_2703,N_27744,N_26006);
and UO_2704 (O_2704,N_24832,N_29345);
and UO_2705 (O_2705,N_26076,N_26182);
or UO_2706 (O_2706,N_29721,N_24927);
xor UO_2707 (O_2707,N_29864,N_29178);
nand UO_2708 (O_2708,N_29565,N_24697);
or UO_2709 (O_2709,N_27845,N_24928);
nand UO_2710 (O_2710,N_27531,N_24189);
nor UO_2711 (O_2711,N_29082,N_29955);
nand UO_2712 (O_2712,N_27212,N_26187);
and UO_2713 (O_2713,N_26385,N_29819);
nand UO_2714 (O_2714,N_27850,N_27658);
nand UO_2715 (O_2715,N_29368,N_29644);
or UO_2716 (O_2716,N_29279,N_25828);
nand UO_2717 (O_2717,N_24643,N_26826);
xnor UO_2718 (O_2718,N_24639,N_27879);
nor UO_2719 (O_2719,N_28561,N_24934);
nor UO_2720 (O_2720,N_24321,N_27365);
nor UO_2721 (O_2721,N_25007,N_24946);
and UO_2722 (O_2722,N_27708,N_28991);
nand UO_2723 (O_2723,N_25017,N_25553);
and UO_2724 (O_2724,N_28174,N_26911);
or UO_2725 (O_2725,N_26491,N_27172);
nor UO_2726 (O_2726,N_29103,N_28453);
or UO_2727 (O_2727,N_27579,N_24971);
or UO_2728 (O_2728,N_24241,N_29029);
nor UO_2729 (O_2729,N_26952,N_24766);
nor UO_2730 (O_2730,N_24622,N_25939);
and UO_2731 (O_2731,N_26521,N_25202);
or UO_2732 (O_2732,N_26681,N_28497);
and UO_2733 (O_2733,N_29860,N_29895);
and UO_2734 (O_2734,N_24217,N_29374);
nor UO_2735 (O_2735,N_24333,N_25053);
or UO_2736 (O_2736,N_28205,N_29254);
nand UO_2737 (O_2737,N_27915,N_28382);
nand UO_2738 (O_2738,N_28338,N_26334);
nor UO_2739 (O_2739,N_29470,N_26230);
xnor UO_2740 (O_2740,N_25182,N_27299);
and UO_2741 (O_2741,N_29099,N_25728);
and UO_2742 (O_2742,N_28305,N_28783);
and UO_2743 (O_2743,N_26566,N_25283);
nand UO_2744 (O_2744,N_25719,N_29403);
nand UO_2745 (O_2745,N_27419,N_24741);
nor UO_2746 (O_2746,N_25488,N_25018);
and UO_2747 (O_2747,N_26244,N_28262);
or UO_2748 (O_2748,N_29447,N_27167);
and UO_2749 (O_2749,N_25023,N_26074);
and UO_2750 (O_2750,N_26595,N_25623);
and UO_2751 (O_2751,N_24854,N_28599);
nand UO_2752 (O_2752,N_29400,N_26056);
nand UO_2753 (O_2753,N_27016,N_28394);
xor UO_2754 (O_2754,N_26177,N_27954);
or UO_2755 (O_2755,N_25425,N_25849);
or UO_2756 (O_2756,N_29671,N_29510);
or UO_2757 (O_2757,N_26203,N_28076);
nor UO_2758 (O_2758,N_29804,N_25702);
nand UO_2759 (O_2759,N_25545,N_24911);
and UO_2760 (O_2760,N_27962,N_26972);
or UO_2761 (O_2761,N_28575,N_29983);
or UO_2762 (O_2762,N_26021,N_28050);
or UO_2763 (O_2763,N_27138,N_28363);
nand UO_2764 (O_2764,N_27116,N_26852);
and UO_2765 (O_2765,N_27469,N_24574);
or UO_2766 (O_2766,N_25369,N_24959);
nor UO_2767 (O_2767,N_28387,N_29469);
or UO_2768 (O_2768,N_29480,N_28725);
nand UO_2769 (O_2769,N_27999,N_27048);
or UO_2770 (O_2770,N_27626,N_25286);
nand UO_2771 (O_2771,N_25320,N_24942);
or UO_2772 (O_2772,N_24062,N_29858);
and UO_2773 (O_2773,N_26658,N_27466);
or UO_2774 (O_2774,N_28995,N_25547);
and UO_2775 (O_2775,N_25989,N_28834);
nand UO_2776 (O_2776,N_29291,N_29104);
nand UO_2777 (O_2777,N_29775,N_25564);
and UO_2778 (O_2778,N_26122,N_29694);
or UO_2779 (O_2779,N_26493,N_28292);
and UO_2780 (O_2780,N_27044,N_27366);
and UO_2781 (O_2781,N_26821,N_27103);
or UO_2782 (O_2782,N_25959,N_28950);
or UO_2783 (O_2783,N_25681,N_28913);
and UO_2784 (O_2784,N_26085,N_25792);
nor UO_2785 (O_2785,N_24200,N_28220);
and UO_2786 (O_2786,N_27282,N_28936);
and UO_2787 (O_2787,N_28761,N_29779);
and UO_2788 (O_2788,N_29792,N_29795);
or UO_2789 (O_2789,N_24604,N_27287);
and UO_2790 (O_2790,N_25797,N_25848);
xor UO_2791 (O_2791,N_28423,N_29516);
or UO_2792 (O_2792,N_27385,N_26665);
nand UO_2793 (O_2793,N_28796,N_24556);
nand UO_2794 (O_2794,N_24430,N_27733);
nor UO_2795 (O_2795,N_26859,N_27795);
or UO_2796 (O_2796,N_24730,N_25281);
nor UO_2797 (O_2797,N_27631,N_28441);
or UO_2798 (O_2798,N_26143,N_25675);
nand UO_2799 (O_2799,N_26137,N_28833);
and UO_2800 (O_2800,N_28965,N_28069);
nor UO_2801 (O_2801,N_25499,N_28330);
or UO_2802 (O_2802,N_24186,N_26971);
nor UO_2803 (O_2803,N_26937,N_29861);
nand UO_2804 (O_2804,N_24548,N_28729);
or UO_2805 (O_2805,N_26153,N_28946);
xnor UO_2806 (O_2806,N_27033,N_28660);
nand UO_2807 (O_2807,N_27337,N_28968);
nand UO_2808 (O_2808,N_29454,N_25684);
and UO_2809 (O_2809,N_24565,N_29116);
or UO_2810 (O_2810,N_24880,N_27491);
or UO_2811 (O_2811,N_26374,N_29304);
or UO_2812 (O_2812,N_28536,N_29629);
xor UO_2813 (O_2813,N_24585,N_29483);
nand UO_2814 (O_2814,N_24442,N_26361);
or UO_2815 (O_2815,N_26270,N_27197);
and UO_2816 (O_2816,N_27938,N_25192);
and UO_2817 (O_2817,N_25443,N_28943);
xnor UO_2818 (O_2818,N_24468,N_27977);
xnor UO_2819 (O_2819,N_28297,N_26094);
nor UO_2820 (O_2820,N_25356,N_29551);
and UO_2821 (O_2821,N_26197,N_24541);
nand UO_2822 (O_2822,N_25503,N_28240);
and UO_2823 (O_2823,N_29372,N_28779);
or UO_2824 (O_2824,N_29292,N_28446);
xnor UO_2825 (O_2825,N_28109,N_28078);
or UO_2826 (O_2826,N_24129,N_29019);
nand UO_2827 (O_2827,N_26405,N_28263);
and UO_2828 (O_2828,N_28521,N_28674);
nor UO_2829 (O_2829,N_29024,N_27450);
nor UO_2830 (O_2830,N_29726,N_29018);
and UO_2831 (O_2831,N_29256,N_28983);
or UO_2832 (O_2832,N_25869,N_29143);
nor UO_2833 (O_2833,N_24318,N_25910);
or UO_2834 (O_2834,N_27860,N_26402);
and UO_2835 (O_2835,N_25494,N_27699);
and UO_2836 (O_2836,N_24460,N_29144);
or UO_2837 (O_2837,N_24603,N_28974);
nand UO_2838 (O_2838,N_27903,N_27144);
or UO_2839 (O_2839,N_28971,N_27604);
and UO_2840 (O_2840,N_28621,N_24527);
nand UO_2841 (O_2841,N_25138,N_24259);
or UO_2842 (O_2842,N_24503,N_26785);
and UO_2843 (O_2843,N_27345,N_26422);
xnor UO_2844 (O_2844,N_29276,N_28052);
or UO_2845 (O_2845,N_26582,N_27422);
nand UO_2846 (O_2846,N_25042,N_29981);
nor UO_2847 (O_2847,N_28817,N_26242);
nand UO_2848 (O_2848,N_25149,N_24338);
nand UO_2849 (O_2849,N_28162,N_25904);
or UO_2850 (O_2850,N_28183,N_29060);
nor UO_2851 (O_2851,N_25505,N_28167);
nor UO_2852 (O_2852,N_28696,N_29030);
nand UO_2853 (O_2853,N_29223,N_28956);
nor UO_2854 (O_2854,N_25087,N_24103);
or UO_2855 (O_2855,N_24000,N_27095);
or UO_2856 (O_2856,N_29815,N_29445);
or UO_2857 (O_2857,N_27136,N_28763);
nand UO_2858 (O_2858,N_29593,N_28734);
or UO_2859 (O_2859,N_25088,N_28819);
nand UO_2860 (O_2860,N_24870,N_24594);
or UO_2861 (O_2861,N_25375,N_26880);
and UO_2862 (O_2862,N_29917,N_27002);
nor UO_2863 (O_2863,N_24281,N_25118);
nor UO_2864 (O_2864,N_26285,N_25036);
nor UO_2865 (O_2865,N_25396,N_28177);
xnor UO_2866 (O_2866,N_24359,N_25808);
or UO_2867 (O_2867,N_29051,N_28004);
xor UO_2868 (O_2868,N_28272,N_26178);
nor UO_2869 (O_2869,N_25465,N_28070);
nand UO_2870 (O_2870,N_28184,N_24406);
nor UO_2871 (O_2871,N_28870,N_26619);
nand UO_2872 (O_2872,N_28207,N_26072);
nand UO_2873 (O_2873,N_25326,N_29529);
nand UO_2874 (O_2874,N_28757,N_29642);
nand UO_2875 (O_2875,N_27110,N_29793);
or UO_2876 (O_2876,N_24257,N_29197);
xnor UO_2877 (O_2877,N_28626,N_26181);
nand UO_2878 (O_2878,N_28260,N_27161);
and UO_2879 (O_2879,N_28756,N_29693);
and UO_2880 (O_2880,N_25379,N_27847);
and UO_2881 (O_2881,N_27486,N_25735);
and UO_2882 (O_2882,N_25903,N_26501);
and UO_2883 (O_2883,N_27624,N_27582);
and UO_2884 (O_2884,N_24358,N_29053);
or UO_2885 (O_2885,N_27333,N_29282);
or UO_2886 (O_2886,N_29156,N_27597);
nand UO_2887 (O_2887,N_26310,N_28758);
xnor UO_2888 (O_2888,N_29303,N_25981);
or UO_2889 (O_2889,N_26890,N_26473);
or UO_2890 (O_2890,N_29888,N_24239);
or UO_2891 (O_2891,N_26147,N_25677);
nand UO_2892 (O_2892,N_29187,N_24099);
nand UO_2893 (O_2893,N_27151,N_28128);
xor UO_2894 (O_2894,N_25528,N_29834);
or UO_2895 (O_2895,N_27015,N_29687);
or UO_2896 (O_2896,N_25444,N_28623);
xor UO_2897 (O_2897,N_28034,N_27844);
and UO_2898 (O_2898,N_28386,N_29278);
xnor UO_2899 (O_2899,N_26265,N_26079);
and UO_2900 (O_2900,N_28005,N_29867);
nand UO_2901 (O_2901,N_27931,N_26121);
nor UO_2902 (O_2902,N_26731,N_27248);
nor UO_2903 (O_2903,N_26811,N_25891);
and UO_2904 (O_2904,N_28115,N_26007);
nand UO_2905 (O_2905,N_29166,N_27862);
xor UO_2906 (O_2906,N_28554,N_28421);
or UO_2907 (O_2907,N_25061,N_29319);
and UO_2908 (O_2908,N_25704,N_28149);
nand UO_2909 (O_2909,N_29297,N_24225);
nor UO_2910 (O_2910,N_26412,N_28310);
and UO_2911 (O_2911,N_24628,N_27609);
nand UO_2912 (O_2912,N_27233,N_27828);
and UO_2913 (O_2913,N_28689,N_27887);
nor UO_2914 (O_2914,N_25996,N_29922);
nand UO_2915 (O_2915,N_28805,N_26656);
nand UO_2916 (O_2916,N_28187,N_28644);
or UO_2917 (O_2917,N_28549,N_25544);
or UO_2918 (O_2918,N_26036,N_26925);
nor UO_2919 (O_2919,N_27832,N_28814);
nor UO_2920 (O_2920,N_27045,N_26504);
xor UO_2921 (O_2921,N_26123,N_29517);
nand UO_2922 (O_2922,N_26425,N_26001);
nor UO_2923 (O_2923,N_27661,N_25590);
and UO_2924 (O_2924,N_29880,N_26910);
or UO_2925 (O_2925,N_25191,N_25597);
xnor UO_2926 (O_2926,N_27383,N_26915);
nand UO_2927 (O_2927,N_26506,N_29780);
or UO_2928 (O_2928,N_28092,N_25531);
and UO_2929 (O_2929,N_26646,N_29047);
or UO_2930 (O_2930,N_26144,N_26371);
or UO_2931 (O_2931,N_26444,N_25567);
xor UO_2932 (O_2932,N_26976,N_25161);
or UO_2933 (O_2933,N_27488,N_24758);
nand UO_2934 (O_2934,N_26543,N_25296);
nand UO_2935 (O_2935,N_28683,N_27043);
nor UO_2936 (O_2936,N_25103,N_25160);
xnor UO_2937 (O_2937,N_28463,N_26629);
and UO_2938 (O_2938,N_28448,N_28715);
nand UO_2939 (O_2939,N_26620,N_27675);
nand UO_2940 (O_2940,N_29951,N_29472);
xnor UO_2941 (O_2941,N_29067,N_24587);
nor UO_2942 (O_2942,N_29015,N_24525);
and UO_2943 (O_2943,N_28987,N_25823);
or UO_2944 (O_2944,N_25417,N_26902);
and UO_2945 (O_2945,N_24252,N_25325);
nand UO_2946 (O_2946,N_25404,N_28850);
nand UO_2947 (O_2947,N_28576,N_27453);
and UO_2948 (O_2948,N_28121,N_25068);
or UO_2949 (O_2949,N_29097,N_28123);
nor UO_2950 (O_2950,N_25723,N_27017);
and UO_2951 (O_2951,N_27165,N_25289);
nor UO_2952 (O_2952,N_25816,N_26667);
and UO_2953 (O_2953,N_28820,N_25733);
xnor UO_2954 (O_2954,N_24264,N_29042);
nor UO_2955 (O_2955,N_26945,N_28525);
nand UO_2956 (O_2956,N_26356,N_24906);
nand UO_2957 (O_2957,N_26866,N_26924);
and UO_2958 (O_2958,N_29376,N_28749);
nand UO_2959 (O_2959,N_27644,N_29484);
nor UO_2960 (O_2960,N_25446,N_25057);
xor UO_2961 (O_2961,N_25548,N_25410);
and UO_2962 (O_2962,N_24317,N_28163);
nand UO_2963 (O_2963,N_29691,N_25633);
nand UO_2964 (O_2964,N_26657,N_28632);
nor UO_2965 (O_2965,N_26864,N_26384);
or UO_2966 (O_2966,N_29994,N_29540);
and UO_2967 (O_2967,N_27890,N_28222);
or UO_2968 (O_2968,N_29252,N_24054);
and UO_2969 (O_2969,N_29255,N_28275);
nor UO_2970 (O_2970,N_27088,N_27195);
and UO_2971 (O_2971,N_29579,N_29253);
or UO_2972 (O_2972,N_25861,N_28618);
nor UO_2973 (O_2973,N_27883,N_25172);
and UO_2974 (O_2974,N_24856,N_26163);
nand UO_2975 (O_2975,N_25102,N_28114);
nand UO_2976 (O_2976,N_29973,N_24216);
or UO_2977 (O_2977,N_28171,N_26806);
nand UO_2978 (O_2978,N_25235,N_24098);
nor UO_2979 (O_2979,N_25748,N_26938);
nor UO_2980 (O_2980,N_28982,N_28462);
and UO_2981 (O_2981,N_27297,N_25133);
and UO_2982 (O_2982,N_25383,N_25570);
nand UO_2983 (O_2983,N_29334,N_25788);
nor UO_2984 (O_2984,N_29402,N_29553);
nor UO_2985 (O_2985,N_27321,N_26274);
and UO_2986 (O_2986,N_28878,N_28810);
and UO_2987 (O_2987,N_24684,N_28256);
or UO_2988 (O_2988,N_25115,N_27084);
xor UO_2989 (O_2989,N_28845,N_27325);
nand UO_2990 (O_2990,N_27361,N_24175);
and UO_2991 (O_2991,N_27595,N_25457);
nand UO_2992 (O_2992,N_27411,N_28308);
xnor UO_2993 (O_2993,N_29698,N_29004);
nor UO_2994 (O_2994,N_27376,N_28866);
or UO_2995 (O_2995,N_25394,N_24638);
and UO_2996 (O_2996,N_29789,N_27827);
and UO_2997 (O_2997,N_24076,N_28488);
and UO_2998 (O_2998,N_26571,N_26183);
and UO_2999 (O_2999,N_29991,N_25614);
nand UO_3000 (O_3000,N_26150,N_25332);
nor UO_3001 (O_3001,N_25009,N_26375);
nor UO_3002 (O_3002,N_28810,N_27353);
and UO_3003 (O_3003,N_26127,N_27949);
or UO_3004 (O_3004,N_27444,N_24516);
or UO_3005 (O_3005,N_24050,N_27933);
xnor UO_3006 (O_3006,N_25552,N_27789);
nand UO_3007 (O_3007,N_27809,N_28459);
and UO_3008 (O_3008,N_24656,N_29908);
nand UO_3009 (O_3009,N_27814,N_29535);
nor UO_3010 (O_3010,N_29760,N_24796);
nand UO_3011 (O_3011,N_29969,N_28251);
nor UO_3012 (O_3012,N_24410,N_24325);
xnor UO_3013 (O_3013,N_24038,N_29736);
and UO_3014 (O_3014,N_25106,N_24170);
xor UO_3015 (O_3015,N_29257,N_24542);
nand UO_3016 (O_3016,N_24747,N_27499);
nand UO_3017 (O_3017,N_28204,N_26598);
nand UO_3018 (O_3018,N_24430,N_28587);
and UO_3019 (O_3019,N_28066,N_27469);
xor UO_3020 (O_3020,N_28962,N_28490);
nand UO_3021 (O_3021,N_27217,N_24443);
or UO_3022 (O_3022,N_27776,N_28295);
nand UO_3023 (O_3023,N_25176,N_25645);
and UO_3024 (O_3024,N_24751,N_27412);
or UO_3025 (O_3025,N_25235,N_27825);
nand UO_3026 (O_3026,N_28344,N_27801);
nor UO_3027 (O_3027,N_24270,N_24384);
nand UO_3028 (O_3028,N_29956,N_24271);
nand UO_3029 (O_3029,N_29355,N_24057);
or UO_3030 (O_3030,N_28865,N_25018);
nand UO_3031 (O_3031,N_26447,N_29031);
xor UO_3032 (O_3032,N_24407,N_27692);
or UO_3033 (O_3033,N_29190,N_29180);
nor UO_3034 (O_3034,N_25367,N_25896);
or UO_3035 (O_3035,N_26314,N_26881);
and UO_3036 (O_3036,N_26543,N_28229);
or UO_3037 (O_3037,N_27190,N_26152);
nand UO_3038 (O_3038,N_26162,N_27654);
or UO_3039 (O_3039,N_24821,N_25708);
or UO_3040 (O_3040,N_25064,N_25008);
or UO_3041 (O_3041,N_26480,N_29098);
nand UO_3042 (O_3042,N_24943,N_24157);
nor UO_3043 (O_3043,N_29870,N_29030);
and UO_3044 (O_3044,N_24636,N_27714);
and UO_3045 (O_3045,N_24428,N_28796);
nand UO_3046 (O_3046,N_26373,N_27287);
or UO_3047 (O_3047,N_27924,N_25147);
and UO_3048 (O_3048,N_28399,N_24996);
or UO_3049 (O_3049,N_26108,N_27216);
or UO_3050 (O_3050,N_24012,N_28866);
or UO_3051 (O_3051,N_28142,N_29958);
or UO_3052 (O_3052,N_24023,N_27600);
or UO_3053 (O_3053,N_28090,N_25054);
xnor UO_3054 (O_3054,N_24079,N_28690);
and UO_3055 (O_3055,N_26733,N_28594);
xor UO_3056 (O_3056,N_24862,N_29838);
nand UO_3057 (O_3057,N_29794,N_28176);
nand UO_3058 (O_3058,N_26741,N_29409);
nor UO_3059 (O_3059,N_28189,N_24531);
xnor UO_3060 (O_3060,N_29992,N_28708);
or UO_3061 (O_3061,N_24669,N_28189);
nand UO_3062 (O_3062,N_26010,N_24079);
nand UO_3063 (O_3063,N_27732,N_28009);
nor UO_3064 (O_3064,N_24179,N_27096);
and UO_3065 (O_3065,N_26326,N_26463);
nand UO_3066 (O_3066,N_25333,N_28936);
nand UO_3067 (O_3067,N_29126,N_27454);
and UO_3068 (O_3068,N_27942,N_25911);
nand UO_3069 (O_3069,N_26316,N_24561);
xor UO_3070 (O_3070,N_28231,N_26390);
xnor UO_3071 (O_3071,N_25223,N_24475);
or UO_3072 (O_3072,N_27459,N_26128);
nor UO_3073 (O_3073,N_26486,N_24213);
or UO_3074 (O_3074,N_27041,N_25133);
or UO_3075 (O_3075,N_25446,N_28923);
or UO_3076 (O_3076,N_24910,N_25156);
nor UO_3077 (O_3077,N_27180,N_24980);
or UO_3078 (O_3078,N_29074,N_27102);
nor UO_3079 (O_3079,N_29915,N_29361);
or UO_3080 (O_3080,N_27665,N_26483);
and UO_3081 (O_3081,N_27159,N_26210);
and UO_3082 (O_3082,N_28119,N_29381);
nand UO_3083 (O_3083,N_26146,N_25588);
and UO_3084 (O_3084,N_27425,N_26258);
nand UO_3085 (O_3085,N_25476,N_26214);
nor UO_3086 (O_3086,N_29771,N_25296);
and UO_3087 (O_3087,N_25426,N_25373);
nor UO_3088 (O_3088,N_24804,N_29881);
or UO_3089 (O_3089,N_24421,N_27218);
nand UO_3090 (O_3090,N_27686,N_26456);
nand UO_3091 (O_3091,N_24870,N_25622);
nand UO_3092 (O_3092,N_28523,N_29846);
or UO_3093 (O_3093,N_24176,N_28579);
nand UO_3094 (O_3094,N_29672,N_24990);
or UO_3095 (O_3095,N_24707,N_29011);
nor UO_3096 (O_3096,N_29742,N_28913);
xor UO_3097 (O_3097,N_28943,N_29708);
xnor UO_3098 (O_3098,N_29621,N_26585);
or UO_3099 (O_3099,N_26290,N_27341);
and UO_3100 (O_3100,N_24205,N_27435);
and UO_3101 (O_3101,N_27659,N_29614);
xor UO_3102 (O_3102,N_27619,N_25181);
nand UO_3103 (O_3103,N_26930,N_29131);
xor UO_3104 (O_3104,N_29734,N_29729);
and UO_3105 (O_3105,N_27319,N_27936);
or UO_3106 (O_3106,N_24651,N_28842);
nand UO_3107 (O_3107,N_29779,N_28836);
nor UO_3108 (O_3108,N_27986,N_24627);
nor UO_3109 (O_3109,N_28276,N_24121);
nand UO_3110 (O_3110,N_27647,N_28443);
or UO_3111 (O_3111,N_29850,N_27029);
nand UO_3112 (O_3112,N_28569,N_26857);
and UO_3113 (O_3113,N_24433,N_28706);
nand UO_3114 (O_3114,N_25772,N_27226);
and UO_3115 (O_3115,N_25002,N_28562);
nand UO_3116 (O_3116,N_27282,N_26773);
nand UO_3117 (O_3117,N_26619,N_28379);
and UO_3118 (O_3118,N_25056,N_25412);
nand UO_3119 (O_3119,N_25341,N_27993);
and UO_3120 (O_3120,N_27783,N_28226);
and UO_3121 (O_3121,N_25713,N_26744);
and UO_3122 (O_3122,N_25635,N_24162);
and UO_3123 (O_3123,N_26749,N_25493);
or UO_3124 (O_3124,N_24288,N_27384);
nand UO_3125 (O_3125,N_26708,N_26209);
or UO_3126 (O_3126,N_25224,N_27220);
nor UO_3127 (O_3127,N_27245,N_27416);
or UO_3128 (O_3128,N_29363,N_26671);
or UO_3129 (O_3129,N_24297,N_28985);
and UO_3130 (O_3130,N_27453,N_25889);
or UO_3131 (O_3131,N_29034,N_26626);
or UO_3132 (O_3132,N_26554,N_25206);
and UO_3133 (O_3133,N_29212,N_25040);
and UO_3134 (O_3134,N_29347,N_27726);
nor UO_3135 (O_3135,N_27632,N_28620);
nor UO_3136 (O_3136,N_29646,N_29963);
nand UO_3137 (O_3137,N_27930,N_26999);
and UO_3138 (O_3138,N_29083,N_27011);
nor UO_3139 (O_3139,N_27736,N_29076);
or UO_3140 (O_3140,N_26385,N_24129);
nor UO_3141 (O_3141,N_25504,N_24887);
or UO_3142 (O_3142,N_28757,N_29624);
or UO_3143 (O_3143,N_28857,N_24317);
xor UO_3144 (O_3144,N_28518,N_27725);
and UO_3145 (O_3145,N_27824,N_28744);
nand UO_3146 (O_3146,N_28101,N_26890);
xor UO_3147 (O_3147,N_24542,N_26594);
nor UO_3148 (O_3148,N_26328,N_26026);
or UO_3149 (O_3149,N_26259,N_24907);
nand UO_3150 (O_3150,N_29516,N_25344);
nand UO_3151 (O_3151,N_27958,N_24120);
nand UO_3152 (O_3152,N_24680,N_26752);
xor UO_3153 (O_3153,N_24917,N_26545);
nor UO_3154 (O_3154,N_26826,N_29006);
nand UO_3155 (O_3155,N_28526,N_26147);
and UO_3156 (O_3156,N_28053,N_29818);
or UO_3157 (O_3157,N_28854,N_28784);
nor UO_3158 (O_3158,N_28258,N_25881);
nand UO_3159 (O_3159,N_29623,N_28111);
or UO_3160 (O_3160,N_26316,N_24135);
or UO_3161 (O_3161,N_27888,N_25892);
nand UO_3162 (O_3162,N_24636,N_24387);
or UO_3163 (O_3163,N_26918,N_24993);
nand UO_3164 (O_3164,N_28075,N_29914);
and UO_3165 (O_3165,N_28532,N_24008);
nor UO_3166 (O_3166,N_28576,N_28928);
or UO_3167 (O_3167,N_26448,N_29354);
nand UO_3168 (O_3168,N_28626,N_29325);
nand UO_3169 (O_3169,N_25711,N_29106);
or UO_3170 (O_3170,N_24524,N_29764);
nor UO_3171 (O_3171,N_24582,N_28390);
or UO_3172 (O_3172,N_29816,N_29562);
nand UO_3173 (O_3173,N_29664,N_25103);
and UO_3174 (O_3174,N_27701,N_24572);
nor UO_3175 (O_3175,N_28088,N_25880);
xnor UO_3176 (O_3176,N_25767,N_28274);
nor UO_3177 (O_3177,N_25643,N_28316);
nand UO_3178 (O_3178,N_26839,N_29007);
nand UO_3179 (O_3179,N_27602,N_24276);
nand UO_3180 (O_3180,N_24886,N_28958);
or UO_3181 (O_3181,N_28623,N_26858);
and UO_3182 (O_3182,N_27994,N_28796);
or UO_3183 (O_3183,N_28060,N_27736);
and UO_3184 (O_3184,N_29538,N_24282);
or UO_3185 (O_3185,N_29584,N_25206);
nand UO_3186 (O_3186,N_25078,N_25142);
nor UO_3187 (O_3187,N_27076,N_25733);
nor UO_3188 (O_3188,N_29353,N_29069);
and UO_3189 (O_3189,N_26949,N_29439);
and UO_3190 (O_3190,N_25202,N_28789);
or UO_3191 (O_3191,N_26352,N_24835);
nor UO_3192 (O_3192,N_25515,N_27961);
and UO_3193 (O_3193,N_24048,N_25137);
or UO_3194 (O_3194,N_24670,N_24725);
and UO_3195 (O_3195,N_26454,N_24966);
nand UO_3196 (O_3196,N_28761,N_27176);
and UO_3197 (O_3197,N_25612,N_25825);
or UO_3198 (O_3198,N_29658,N_28833);
or UO_3199 (O_3199,N_27605,N_25736);
xnor UO_3200 (O_3200,N_29587,N_25591);
and UO_3201 (O_3201,N_24946,N_27119);
xor UO_3202 (O_3202,N_25362,N_24030);
or UO_3203 (O_3203,N_28836,N_24988);
xnor UO_3204 (O_3204,N_29512,N_26785);
nor UO_3205 (O_3205,N_28716,N_27829);
nand UO_3206 (O_3206,N_29211,N_28741);
nand UO_3207 (O_3207,N_28510,N_25593);
xor UO_3208 (O_3208,N_28603,N_28515);
and UO_3209 (O_3209,N_29384,N_28633);
xor UO_3210 (O_3210,N_26182,N_25539);
nor UO_3211 (O_3211,N_29224,N_26740);
nand UO_3212 (O_3212,N_29264,N_27465);
and UO_3213 (O_3213,N_25278,N_28186);
nor UO_3214 (O_3214,N_24465,N_24694);
nor UO_3215 (O_3215,N_26174,N_29404);
nor UO_3216 (O_3216,N_26869,N_28727);
or UO_3217 (O_3217,N_28717,N_28876);
nor UO_3218 (O_3218,N_26736,N_29778);
or UO_3219 (O_3219,N_29316,N_28097);
and UO_3220 (O_3220,N_28985,N_27398);
or UO_3221 (O_3221,N_26790,N_29894);
nand UO_3222 (O_3222,N_25994,N_28690);
nor UO_3223 (O_3223,N_26494,N_24758);
or UO_3224 (O_3224,N_24950,N_29253);
and UO_3225 (O_3225,N_26029,N_28185);
and UO_3226 (O_3226,N_24739,N_25942);
nor UO_3227 (O_3227,N_28326,N_29890);
or UO_3228 (O_3228,N_28109,N_26647);
nor UO_3229 (O_3229,N_24982,N_29299);
nand UO_3230 (O_3230,N_29954,N_25141);
or UO_3231 (O_3231,N_24726,N_27431);
nor UO_3232 (O_3232,N_26191,N_29053);
nand UO_3233 (O_3233,N_24349,N_29838);
and UO_3234 (O_3234,N_24316,N_27991);
nor UO_3235 (O_3235,N_28815,N_26136);
or UO_3236 (O_3236,N_29782,N_25918);
nand UO_3237 (O_3237,N_24061,N_26905);
and UO_3238 (O_3238,N_29261,N_24887);
xor UO_3239 (O_3239,N_28512,N_28470);
and UO_3240 (O_3240,N_27902,N_25549);
nor UO_3241 (O_3241,N_26498,N_29386);
or UO_3242 (O_3242,N_27530,N_24604);
xor UO_3243 (O_3243,N_25614,N_29016);
or UO_3244 (O_3244,N_26797,N_24993);
nor UO_3245 (O_3245,N_27823,N_26797);
nand UO_3246 (O_3246,N_26440,N_24124);
and UO_3247 (O_3247,N_26213,N_27921);
xnor UO_3248 (O_3248,N_24759,N_29730);
and UO_3249 (O_3249,N_28089,N_24642);
or UO_3250 (O_3250,N_29710,N_24735);
or UO_3251 (O_3251,N_29481,N_25712);
or UO_3252 (O_3252,N_26152,N_28071);
nor UO_3253 (O_3253,N_25713,N_26420);
and UO_3254 (O_3254,N_27314,N_24711);
nor UO_3255 (O_3255,N_28111,N_28274);
or UO_3256 (O_3256,N_24077,N_25239);
nor UO_3257 (O_3257,N_29306,N_29821);
nand UO_3258 (O_3258,N_25047,N_29387);
or UO_3259 (O_3259,N_26884,N_25518);
nor UO_3260 (O_3260,N_28614,N_27476);
and UO_3261 (O_3261,N_24413,N_25959);
and UO_3262 (O_3262,N_27897,N_27017);
nand UO_3263 (O_3263,N_27137,N_26204);
and UO_3264 (O_3264,N_26091,N_29393);
nand UO_3265 (O_3265,N_26840,N_28416);
or UO_3266 (O_3266,N_28068,N_26938);
xor UO_3267 (O_3267,N_25729,N_26838);
and UO_3268 (O_3268,N_29291,N_24001);
and UO_3269 (O_3269,N_26331,N_27867);
or UO_3270 (O_3270,N_25099,N_29877);
xnor UO_3271 (O_3271,N_29802,N_26764);
or UO_3272 (O_3272,N_28004,N_25467);
and UO_3273 (O_3273,N_27274,N_27583);
xor UO_3274 (O_3274,N_25574,N_29163);
nand UO_3275 (O_3275,N_27872,N_26142);
and UO_3276 (O_3276,N_28192,N_29256);
nor UO_3277 (O_3277,N_26911,N_26993);
or UO_3278 (O_3278,N_26858,N_27448);
and UO_3279 (O_3279,N_25723,N_29803);
nor UO_3280 (O_3280,N_29060,N_25731);
or UO_3281 (O_3281,N_28912,N_24256);
nand UO_3282 (O_3282,N_26924,N_25317);
nor UO_3283 (O_3283,N_27531,N_26909);
xor UO_3284 (O_3284,N_24413,N_29076);
or UO_3285 (O_3285,N_27033,N_29525);
or UO_3286 (O_3286,N_26413,N_27544);
nor UO_3287 (O_3287,N_26565,N_29539);
and UO_3288 (O_3288,N_26453,N_29051);
nor UO_3289 (O_3289,N_28894,N_25188);
nand UO_3290 (O_3290,N_28850,N_27665);
nand UO_3291 (O_3291,N_25959,N_25775);
and UO_3292 (O_3292,N_28285,N_27884);
xor UO_3293 (O_3293,N_28147,N_24455);
and UO_3294 (O_3294,N_28964,N_28136);
or UO_3295 (O_3295,N_26741,N_26038);
nand UO_3296 (O_3296,N_28129,N_24949);
nand UO_3297 (O_3297,N_25636,N_27269);
nor UO_3298 (O_3298,N_27803,N_24923);
nand UO_3299 (O_3299,N_24211,N_25399);
nor UO_3300 (O_3300,N_28233,N_29472);
and UO_3301 (O_3301,N_28337,N_24906);
and UO_3302 (O_3302,N_24672,N_27173);
or UO_3303 (O_3303,N_24473,N_29723);
and UO_3304 (O_3304,N_26986,N_28423);
xor UO_3305 (O_3305,N_26224,N_27998);
and UO_3306 (O_3306,N_28434,N_26257);
nor UO_3307 (O_3307,N_28744,N_29357);
nor UO_3308 (O_3308,N_24770,N_29008);
nor UO_3309 (O_3309,N_26618,N_27376);
nand UO_3310 (O_3310,N_29338,N_27283);
and UO_3311 (O_3311,N_24883,N_26604);
nand UO_3312 (O_3312,N_26232,N_24052);
nand UO_3313 (O_3313,N_24261,N_26026);
or UO_3314 (O_3314,N_29538,N_27537);
nor UO_3315 (O_3315,N_27748,N_27642);
nand UO_3316 (O_3316,N_27818,N_25875);
and UO_3317 (O_3317,N_26913,N_26025);
and UO_3318 (O_3318,N_27316,N_26813);
nand UO_3319 (O_3319,N_24845,N_27800);
or UO_3320 (O_3320,N_25203,N_25803);
nor UO_3321 (O_3321,N_25454,N_27281);
nand UO_3322 (O_3322,N_25551,N_28097);
nand UO_3323 (O_3323,N_28204,N_27432);
nor UO_3324 (O_3324,N_29206,N_26732);
nand UO_3325 (O_3325,N_26573,N_24207);
nor UO_3326 (O_3326,N_24476,N_26154);
nor UO_3327 (O_3327,N_29801,N_26415);
nor UO_3328 (O_3328,N_27967,N_25201);
nor UO_3329 (O_3329,N_28701,N_28247);
or UO_3330 (O_3330,N_28788,N_29099);
xor UO_3331 (O_3331,N_25281,N_27300);
or UO_3332 (O_3332,N_25400,N_26648);
and UO_3333 (O_3333,N_25605,N_24800);
or UO_3334 (O_3334,N_26583,N_25633);
nor UO_3335 (O_3335,N_26440,N_26589);
nand UO_3336 (O_3336,N_26007,N_24351);
or UO_3337 (O_3337,N_24410,N_28241);
nand UO_3338 (O_3338,N_27700,N_24843);
xor UO_3339 (O_3339,N_27052,N_25131);
nor UO_3340 (O_3340,N_28693,N_28489);
or UO_3341 (O_3341,N_24693,N_25190);
nor UO_3342 (O_3342,N_28527,N_24732);
nand UO_3343 (O_3343,N_25267,N_25960);
nor UO_3344 (O_3344,N_28843,N_26409);
and UO_3345 (O_3345,N_27221,N_26013);
or UO_3346 (O_3346,N_25156,N_26371);
nor UO_3347 (O_3347,N_27039,N_28358);
xor UO_3348 (O_3348,N_26295,N_28307);
nor UO_3349 (O_3349,N_26493,N_26573);
or UO_3350 (O_3350,N_25447,N_24576);
or UO_3351 (O_3351,N_29090,N_27715);
nor UO_3352 (O_3352,N_27612,N_25807);
and UO_3353 (O_3353,N_29446,N_29889);
nand UO_3354 (O_3354,N_24487,N_29646);
xor UO_3355 (O_3355,N_29707,N_24490);
and UO_3356 (O_3356,N_24639,N_28826);
and UO_3357 (O_3357,N_28692,N_27975);
and UO_3358 (O_3358,N_27045,N_24754);
nor UO_3359 (O_3359,N_25914,N_28805);
and UO_3360 (O_3360,N_26240,N_29715);
xor UO_3361 (O_3361,N_26728,N_27908);
nand UO_3362 (O_3362,N_29390,N_26983);
nand UO_3363 (O_3363,N_26111,N_27792);
and UO_3364 (O_3364,N_27579,N_24754);
nor UO_3365 (O_3365,N_25713,N_28128);
xnor UO_3366 (O_3366,N_29572,N_25616);
and UO_3367 (O_3367,N_26609,N_29470);
nand UO_3368 (O_3368,N_24049,N_29173);
or UO_3369 (O_3369,N_24979,N_29755);
nand UO_3370 (O_3370,N_28500,N_25034);
nor UO_3371 (O_3371,N_26872,N_24755);
nand UO_3372 (O_3372,N_24010,N_25842);
nor UO_3373 (O_3373,N_26581,N_26730);
nor UO_3374 (O_3374,N_29326,N_24449);
and UO_3375 (O_3375,N_24097,N_29748);
and UO_3376 (O_3376,N_26552,N_26067);
and UO_3377 (O_3377,N_26948,N_24235);
or UO_3378 (O_3378,N_29365,N_24552);
nor UO_3379 (O_3379,N_27723,N_26333);
and UO_3380 (O_3380,N_28923,N_26586);
nor UO_3381 (O_3381,N_25129,N_28418);
xor UO_3382 (O_3382,N_24468,N_28329);
nand UO_3383 (O_3383,N_28620,N_25764);
nand UO_3384 (O_3384,N_28450,N_24906);
or UO_3385 (O_3385,N_27828,N_27009);
xor UO_3386 (O_3386,N_27760,N_25651);
or UO_3387 (O_3387,N_29068,N_27202);
nor UO_3388 (O_3388,N_25910,N_27575);
or UO_3389 (O_3389,N_27399,N_25171);
and UO_3390 (O_3390,N_28816,N_27934);
or UO_3391 (O_3391,N_27534,N_24483);
xor UO_3392 (O_3392,N_25445,N_28250);
nand UO_3393 (O_3393,N_27532,N_29485);
and UO_3394 (O_3394,N_25314,N_27662);
and UO_3395 (O_3395,N_24229,N_29815);
or UO_3396 (O_3396,N_29065,N_29350);
and UO_3397 (O_3397,N_24523,N_29793);
nand UO_3398 (O_3398,N_29962,N_25175);
nor UO_3399 (O_3399,N_28483,N_28473);
or UO_3400 (O_3400,N_25529,N_27350);
nor UO_3401 (O_3401,N_25187,N_26493);
and UO_3402 (O_3402,N_28285,N_27300);
nand UO_3403 (O_3403,N_28658,N_25573);
and UO_3404 (O_3404,N_29149,N_27043);
or UO_3405 (O_3405,N_25488,N_25626);
nand UO_3406 (O_3406,N_28155,N_28060);
or UO_3407 (O_3407,N_24223,N_29167);
nand UO_3408 (O_3408,N_24146,N_26961);
nand UO_3409 (O_3409,N_28045,N_29670);
and UO_3410 (O_3410,N_29786,N_24554);
and UO_3411 (O_3411,N_26713,N_25856);
nand UO_3412 (O_3412,N_25860,N_25949);
xor UO_3413 (O_3413,N_26131,N_25506);
nand UO_3414 (O_3414,N_29485,N_26510);
nor UO_3415 (O_3415,N_28768,N_29220);
or UO_3416 (O_3416,N_29427,N_28331);
and UO_3417 (O_3417,N_28840,N_26261);
nor UO_3418 (O_3418,N_27560,N_29175);
nor UO_3419 (O_3419,N_26382,N_27154);
nor UO_3420 (O_3420,N_29239,N_26911);
nand UO_3421 (O_3421,N_29322,N_28996);
nand UO_3422 (O_3422,N_25305,N_26242);
or UO_3423 (O_3423,N_26263,N_28039);
and UO_3424 (O_3424,N_24432,N_28680);
or UO_3425 (O_3425,N_27797,N_25177);
or UO_3426 (O_3426,N_28337,N_24524);
or UO_3427 (O_3427,N_24149,N_24885);
and UO_3428 (O_3428,N_28062,N_27151);
and UO_3429 (O_3429,N_27015,N_27733);
and UO_3430 (O_3430,N_29890,N_28912);
and UO_3431 (O_3431,N_26535,N_28494);
and UO_3432 (O_3432,N_26246,N_29213);
nor UO_3433 (O_3433,N_25099,N_29627);
nor UO_3434 (O_3434,N_27242,N_28293);
and UO_3435 (O_3435,N_28916,N_27902);
nor UO_3436 (O_3436,N_29829,N_29782);
nor UO_3437 (O_3437,N_26159,N_29364);
nand UO_3438 (O_3438,N_27912,N_29450);
nand UO_3439 (O_3439,N_29423,N_25589);
and UO_3440 (O_3440,N_25783,N_26810);
and UO_3441 (O_3441,N_29047,N_27305);
and UO_3442 (O_3442,N_29982,N_29418);
and UO_3443 (O_3443,N_26335,N_25450);
nand UO_3444 (O_3444,N_25223,N_29602);
nand UO_3445 (O_3445,N_24177,N_28437);
nand UO_3446 (O_3446,N_28985,N_25570);
nor UO_3447 (O_3447,N_26103,N_24329);
xor UO_3448 (O_3448,N_29526,N_28113);
nor UO_3449 (O_3449,N_28073,N_28015);
and UO_3450 (O_3450,N_28750,N_26927);
and UO_3451 (O_3451,N_29266,N_24007);
or UO_3452 (O_3452,N_28624,N_29192);
or UO_3453 (O_3453,N_26986,N_24288);
nor UO_3454 (O_3454,N_27035,N_29356);
or UO_3455 (O_3455,N_26840,N_26690);
nand UO_3456 (O_3456,N_24905,N_24330);
or UO_3457 (O_3457,N_25223,N_28615);
nor UO_3458 (O_3458,N_29784,N_26794);
nand UO_3459 (O_3459,N_26570,N_26606);
nor UO_3460 (O_3460,N_24263,N_24687);
and UO_3461 (O_3461,N_28419,N_24789);
nor UO_3462 (O_3462,N_28918,N_28334);
and UO_3463 (O_3463,N_28270,N_24160);
nor UO_3464 (O_3464,N_24191,N_24458);
and UO_3465 (O_3465,N_25044,N_27447);
nor UO_3466 (O_3466,N_25605,N_28909);
or UO_3467 (O_3467,N_29977,N_24990);
nand UO_3468 (O_3468,N_29781,N_29713);
and UO_3469 (O_3469,N_27347,N_25872);
nor UO_3470 (O_3470,N_27342,N_25280);
nor UO_3471 (O_3471,N_29047,N_25874);
or UO_3472 (O_3472,N_28453,N_26537);
nand UO_3473 (O_3473,N_26529,N_26373);
nor UO_3474 (O_3474,N_27921,N_26555);
nor UO_3475 (O_3475,N_24316,N_24188);
nand UO_3476 (O_3476,N_26344,N_25080);
or UO_3477 (O_3477,N_26232,N_27242);
nand UO_3478 (O_3478,N_24214,N_26584);
xor UO_3479 (O_3479,N_26261,N_28973);
and UO_3480 (O_3480,N_29036,N_24685);
or UO_3481 (O_3481,N_24592,N_24067);
nor UO_3482 (O_3482,N_29450,N_29845);
nand UO_3483 (O_3483,N_25007,N_28338);
nand UO_3484 (O_3484,N_26774,N_24244);
and UO_3485 (O_3485,N_29022,N_25732);
and UO_3486 (O_3486,N_28892,N_29914);
nor UO_3487 (O_3487,N_28069,N_28805);
nand UO_3488 (O_3488,N_26989,N_28318);
nand UO_3489 (O_3489,N_24816,N_26757);
nand UO_3490 (O_3490,N_27704,N_24893);
or UO_3491 (O_3491,N_25665,N_29672);
and UO_3492 (O_3492,N_26253,N_28102);
nor UO_3493 (O_3493,N_28747,N_29520);
xor UO_3494 (O_3494,N_26624,N_27377);
nor UO_3495 (O_3495,N_26650,N_27324);
or UO_3496 (O_3496,N_27014,N_27907);
nor UO_3497 (O_3497,N_24286,N_24136);
nand UO_3498 (O_3498,N_29721,N_25628);
nor UO_3499 (O_3499,N_27746,N_24594);
endmodule