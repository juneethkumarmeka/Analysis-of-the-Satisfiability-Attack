module basic_750_5000_1000_50_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_372,In_587);
nand U1 (N_1,In_41,In_168);
or U2 (N_2,In_490,In_63);
xor U3 (N_3,In_698,In_197);
nor U4 (N_4,In_86,In_282);
nand U5 (N_5,In_248,In_87);
and U6 (N_6,In_458,In_457);
nand U7 (N_7,In_465,In_169);
and U8 (N_8,In_747,In_231);
and U9 (N_9,In_68,In_193);
nand U10 (N_10,In_230,In_551);
nor U11 (N_11,In_390,In_331);
nor U12 (N_12,In_410,In_638);
nor U13 (N_13,In_147,In_164);
nor U14 (N_14,In_515,In_318);
nor U15 (N_15,In_275,In_603);
and U16 (N_16,In_313,In_46);
xor U17 (N_17,In_292,In_732);
or U18 (N_18,In_257,In_262);
or U19 (N_19,In_142,In_353);
nand U20 (N_20,In_583,In_427);
and U21 (N_21,In_133,In_308);
and U22 (N_22,In_88,In_101);
nand U23 (N_23,In_12,In_527);
nand U24 (N_24,In_42,In_387);
xnor U25 (N_25,In_389,In_417);
nor U26 (N_26,In_192,In_366);
nand U27 (N_27,In_272,In_98);
nand U28 (N_28,In_478,In_489);
nor U29 (N_29,In_109,In_117);
nand U30 (N_30,In_559,In_243);
xor U31 (N_31,In_582,In_635);
nor U32 (N_32,In_64,In_425);
nor U33 (N_33,In_496,In_207);
nand U34 (N_34,In_202,In_150);
or U35 (N_35,In_391,In_524);
and U36 (N_36,In_49,In_153);
or U37 (N_37,In_615,In_20);
or U38 (N_38,In_556,In_344);
nor U39 (N_39,In_673,In_362);
or U40 (N_40,In_36,In_421);
nand U41 (N_41,In_249,In_370);
nand U42 (N_42,In_376,In_60);
xor U43 (N_43,In_704,In_10);
nand U44 (N_44,In_212,In_729);
or U45 (N_45,In_735,In_518);
or U46 (N_46,In_359,In_349);
nor U47 (N_47,In_360,In_239);
or U48 (N_48,In_595,In_283);
nor U49 (N_49,In_552,In_733);
nand U50 (N_50,In_691,In_663);
nor U51 (N_51,In_497,In_251);
nor U52 (N_52,In_462,In_121);
or U53 (N_53,In_204,In_571);
or U54 (N_54,In_45,In_166);
or U55 (N_55,In_707,In_232);
nand U56 (N_56,In_53,In_529);
and U57 (N_57,In_383,In_554);
or U58 (N_58,In_711,In_434);
or U59 (N_59,In_633,In_709);
xor U60 (N_60,In_67,In_560);
and U61 (N_61,In_599,In_306);
nor U62 (N_62,In_361,In_543);
and U63 (N_63,In_508,In_749);
and U64 (N_64,In_244,In_575);
nor U65 (N_65,In_75,In_72);
nor U66 (N_66,In_548,In_172);
or U67 (N_67,In_473,In_509);
nand U68 (N_68,In_126,In_165);
and U69 (N_69,In_734,In_499);
and U70 (N_70,In_507,In_184);
or U71 (N_71,In_480,In_640);
nor U72 (N_72,In_6,In_468);
and U73 (N_73,In_479,In_430);
nor U74 (N_74,In_661,In_189);
or U75 (N_75,In_301,In_606);
or U76 (N_76,In_748,In_65);
nand U77 (N_77,In_510,In_82);
xnor U78 (N_78,In_284,In_122);
and U79 (N_79,In_1,In_89);
nand U80 (N_80,In_608,In_297);
and U81 (N_81,In_73,In_211);
and U82 (N_82,In_415,In_450);
or U83 (N_83,In_352,In_135);
and U84 (N_84,In_550,In_423);
and U85 (N_85,In_697,In_573);
and U86 (N_86,In_668,In_354);
nor U87 (N_87,In_336,In_69);
or U88 (N_88,In_738,In_730);
nand U89 (N_89,In_238,In_157);
or U90 (N_90,In_144,In_25);
nor U91 (N_91,In_541,In_534);
and U92 (N_92,In_482,In_335);
and U93 (N_93,In_500,In_14);
and U94 (N_94,In_128,In_31);
nor U95 (N_95,In_676,In_535);
nor U96 (N_96,In_130,In_652);
nand U97 (N_97,In_356,In_302);
and U98 (N_98,In_409,In_127);
or U99 (N_99,In_487,In_286);
nor U100 (N_100,In_634,In_23);
nor U101 (N_101,N_39,In_287);
nand U102 (N_102,In_293,N_53);
and U103 (N_103,N_90,N_54);
and U104 (N_104,N_42,N_64);
or U105 (N_105,In_276,In_371);
nand U106 (N_106,In_213,In_520);
nor U107 (N_107,N_83,In_437);
and U108 (N_108,In_728,In_546);
nand U109 (N_109,N_85,N_61);
nand U110 (N_110,In_96,N_88);
nand U111 (N_111,In_493,In_446);
or U112 (N_112,In_722,In_432);
nor U113 (N_113,In_50,In_667);
and U114 (N_114,In_62,In_317);
or U115 (N_115,In_187,In_623);
nand U116 (N_116,In_481,In_324);
nand U117 (N_117,In_201,In_616);
xnor U118 (N_118,In_678,In_210);
and U119 (N_119,In_38,In_483);
nand U120 (N_120,In_537,N_43);
nand U121 (N_121,In_99,In_669);
xnor U122 (N_122,In_312,In_588);
nor U123 (N_123,N_82,N_8);
and U124 (N_124,In_449,In_630);
and U125 (N_125,In_355,In_93);
nand U126 (N_126,N_28,N_73);
nand U127 (N_127,In_268,In_622);
nand U128 (N_128,In_382,In_627);
xnor U129 (N_129,In_555,In_112);
and U130 (N_130,In_533,In_338);
nor U131 (N_131,In_158,N_71);
or U132 (N_132,In_380,In_628);
nor U133 (N_133,In_436,In_717);
and U134 (N_134,In_593,In_680);
and U135 (N_135,In_137,In_584);
nand U136 (N_136,In_447,N_65);
nand U137 (N_137,In_596,In_162);
and U138 (N_138,N_6,In_525);
nor U139 (N_139,In_377,In_245);
and U140 (N_140,In_107,In_206);
nor U141 (N_141,In_196,In_672);
nor U142 (N_142,In_102,N_30);
and U143 (N_143,In_506,In_28);
and U144 (N_144,In_636,In_580);
and U145 (N_145,In_208,N_27);
or U146 (N_146,In_674,In_670);
nor U147 (N_147,N_16,In_439);
and U148 (N_148,In_666,In_547);
and U149 (N_149,In_739,In_81);
nand U150 (N_150,In_474,In_33);
nor U151 (N_151,In_186,In_532);
or U152 (N_152,N_50,In_624);
and U153 (N_153,In_11,In_565);
or U154 (N_154,In_339,In_92);
and U155 (N_155,In_263,In_330);
and U156 (N_156,In_725,In_205);
nand U157 (N_157,In_323,In_74);
nand U158 (N_158,N_10,In_646);
or U159 (N_159,In_71,N_26);
nor U160 (N_160,In_332,N_47);
nor U161 (N_161,In_326,N_29);
or U162 (N_162,In_113,In_270);
and U163 (N_163,In_316,In_718);
nor U164 (N_164,In_281,In_348);
or U165 (N_165,In_104,In_378);
or U166 (N_166,In_413,In_77);
or U167 (N_167,In_218,In_236);
nor U168 (N_168,N_20,In_440);
nor U169 (N_169,In_684,In_598);
and U170 (N_170,In_305,In_374);
or U171 (N_171,In_737,In_601);
nor U172 (N_172,In_645,In_219);
nand U173 (N_173,In_328,N_79);
or U174 (N_174,In_295,In_265);
and U175 (N_175,In_18,N_77);
nand U176 (N_176,In_341,N_56);
and U177 (N_177,N_14,In_574);
nand U178 (N_178,In_176,N_7);
and U179 (N_179,In_76,N_94);
and U180 (N_180,In_629,In_394);
nor U181 (N_181,In_225,In_146);
nor U182 (N_182,In_47,In_54);
nand U183 (N_183,In_91,In_505);
nand U184 (N_184,In_40,In_492);
or U185 (N_185,In_736,In_369);
nor U186 (N_186,In_160,In_229);
and U187 (N_187,In_3,N_44);
or U188 (N_188,In_405,In_719);
nand U189 (N_189,In_381,In_716);
nand U190 (N_190,In_141,In_407);
nand U191 (N_191,In_456,In_151);
nand U192 (N_192,In_644,N_40);
nand U193 (N_193,In_343,In_228);
xnor U194 (N_194,In_538,In_291);
nor U195 (N_195,In_161,In_241);
nand U196 (N_196,In_264,In_626);
nand U197 (N_197,In_589,In_617);
xnor U198 (N_198,In_149,In_513);
and U199 (N_199,N_92,In_119);
and U200 (N_200,In_428,In_375);
and U201 (N_201,N_166,In_303);
nor U202 (N_202,N_74,In_233);
nand U203 (N_203,In_654,In_105);
nor U204 (N_204,In_677,In_411);
and U205 (N_205,In_124,N_180);
nand U206 (N_206,In_521,N_190);
nor U207 (N_207,N_60,In_118);
nand U208 (N_208,In_591,N_150);
nand U209 (N_209,In_22,In_424);
nand U210 (N_210,In_278,N_55);
or U211 (N_211,In_30,In_731);
nand U212 (N_212,In_299,In_442);
and U213 (N_213,In_319,In_581);
nand U214 (N_214,N_66,In_116);
nor U215 (N_215,In_191,N_96);
nor U216 (N_216,N_57,In_234);
and U217 (N_217,N_140,In_727);
or U218 (N_218,In_246,In_198);
nor U219 (N_219,In_200,N_106);
or U220 (N_220,In_743,In_441);
or U221 (N_221,In_544,In_134);
nand U222 (N_222,N_187,In_215);
nor U223 (N_223,N_161,In_259);
and U224 (N_224,In_167,N_136);
and U225 (N_225,N_170,In_396);
nor U226 (N_226,In_594,N_67);
xor U227 (N_227,In_123,In_611);
and U228 (N_228,In_511,In_679);
or U229 (N_229,In_563,N_138);
nor U230 (N_230,In_138,N_36);
nor U231 (N_231,In_177,N_182);
or U232 (N_232,In_37,N_4);
nand U233 (N_233,In_252,N_80);
nor U234 (N_234,In_604,N_68);
or U235 (N_235,N_23,In_643);
or U236 (N_236,N_5,N_38);
and U237 (N_237,In_452,In_83);
and U238 (N_238,In_346,In_240);
nand U239 (N_239,In_700,In_55);
nand U240 (N_240,In_685,N_45);
xor U241 (N_241,In_609,N_1);
and U242 (N_242,N_179,In_435);
nand U243 (N_243,In_539,In_656);
and U244 (N_244,In_84,In_683);
xor U245 (N_245,In_398,N_99);
nand U246 (N_246,In_715,In_742);
nand U247 (N_247,In_620,In_406);
or U248 (N_248,N_124,In_576);
and U249 (N_249,In_364,N_111);
nand U250 (N_250,In_572,In_562);
nor U251 (N_251,In_618,In_746);
and U252 (N_252,In_693,In_702);
and U253 (N_253,N_87,In_558);
nand U254 (N_254,In_400,N_192);
nand U255 (N_255,N_160,In_567);
and U256 (N_256,In_528,N_112);
and U257 (N_257,N_35,In_269);
and U258 (N_258,N_153,N_165);
nor U259 (N_259,In_460,In_311);
or U260 (N_260,N_152,N_157);
and U261 (N_261,In_592,N_18);
nor U262 (N_262,N_146,In_597);
and U263 (N_263,In_498,In_57);
nor U264 (N_264,N_169,N_75);
or U265 (N_265,In_255,In_561);
and U266 (N_266,In_0,In_58);
nand U267 (N_267,In_132,In_108);
xnor U268 (N_268,N_13,In_358);
nor U269 (N_269,In_300,In_687);
nand U270 (N_270,N_91,In_488);
and U271 (N_271,N_9,N_143);
nand U272 (N_272,In_433,N_175);
nand U273 (N_273,In_185,In_512);
nand U274 (N_274,In_621,In_170);
nand U275 (N_275,N_119,In_298);
or U276 (N_276,In_531,In_723);
nor U277 (N_277,In_214,In_494);
or U278 (N_278,In_59,In_614);
and U279 (N_279,N_125,In_106);
or U280 (N_280,In_545,In_256);
and U281 (N_281,N_193,N_188);
or U282 (N_282,N_162,In_414);
nor U283 (N_283,In_392,In_412);
nor U284 (N_284,In_342,In_540);
or U285 (N_285,In_664,In_688);
or U286 (N_286,N_21,N_113);
or U287 (N_287,In_431,N_116);
and U288 (N_288,N_155,N_158);
and U289 (N_289,In_173,In_470);
nand U290 (N_290,N_103,In_464);
nor U291 (N_291,N_22,In_156);
nor U292 (N_292,N_11,N_59);
xor U293 (N_293,In_475,In_451);
nand U294 (N_294,In_29,N_148);
nor U295 (N_295,N_164,N_122);
or U296 (N_296,N_151,In_152);
or U297 (N_297,In_397,In_665);
and U298 (N_298,In_115,In_315);
or U299 (N_299,In_27,N_135);
nand U300 (N_300,N_232,N_105);
and U301 (N_301,N_81,In_386);
or U302 (N_302,In_662,In_337);
nand U303 (N_303,In_517,N_227);
and U304 (N_304,N_263,N_97);
nor U305 (N_305,In_222,N_274);
nand U306 (N_306,In_70,N_267);
xor U307 (N_307,N_256,In_741);
nand U308 (N_308,In_129,In_4);
and U309 (N_309,In_658,N_273);
xnor U310 (N_310,In_103,N_194);
or U311 (N_311,In_659,In_461);
and U312 (N_312,N_284,In_174);
nand U313 (N_313,N_149,In_347);
nor U314 (N_314,In_448,In_477);
or U315 (N_315,In_395,N_108);
nor U316 (N_316,In_250,N_132);
or U317 (N_317,N_63,In_689);
or U318 (N_318,In_110,In_469);
nand U319 (N_319,N_218,In_61);
and U320 (N_320,N_202,N_104);
or U321 (N_321,N_24,N_250);
nor U322 (N_322,N_261,N_255);
or U323 (N_323,In_9,In_463);
nor U324 (N_324,N_117,N_209);
or U325 (N_325,N_196,In_221);
nand U326 (N_326,In_296,N_120);
or U327 (N_327,In_17,N_72);
nand U328 (N_328,N_212,N_230);
and U329 (N_329,In_714,In_639);
or U330 (N_330,In_280,In_13);
nor U331 (N_331,In_519,N_34);
nor U332 (N_332,N_183,N_228);
nor U333 (N_333,N_290,In_329);
and U334 (N_334,In_159,In_351);
and U335 (N_335,In_388,N_134);
or U336 (N_336,N_251,In_675);
nor U337 (N_337,N_174,In_80);
and U338 (N_338,In_651,In_368);
or U339 (N_339,In_642,In_586);
or U340 (N_340,N_292,N_197);
and U341 (N_341,In_379,N_115);
and U342 (N_342,In_579,N_185);
or U343 (N_343,In_217,In_273);
or U344 (N_344,N_118,In_694);
nand U345 (N_345,N_260,In_699);
and U346 (N_346,N_127,In_471);
or U347 (N_347,In_569,N_206);
or U348 (N_348,In_226,N_195);
and U349 (N_349,N_239,N_213);
and U350 (N_350,N_171,N_177);
or U351 (N_351,N_217,N_109);
and U352 (N_352,In_455,In_564);
and U353 (N_353,N_244,N_142);
and U354 (N_354,In_467,N_139);
or U355 (N_355,In_472,N_31);
or U356 (N_356,In_454,In_223);
or U357 (N_357,In_365,In_237);
and U358 (N_358,In_43,In_503);
nand U359 (N_359,N_76,In_304);
or U360 (N_360,In_209,In_536);
nor U361 (N_361,N_298,In_612);
or U362 (N_362,In_66,N_121);
and U363 (N_363,N_236,In_285);
xnor U364 (N_364,In_476,In_648);
xnor U365 (N_365,In_274,In_502);
nand U366 (N_366,In_632,In_114);
or U367 (N_367,In_570,In_602);
nand U368 (N_368,N_225,In_51);
nand U369 (N_369,In_24,In_310);
nand U370 (N_370,N_51,In_557);
nand U371 (N_371,N_12,In_485);
or U372 (N_372,In_466,N_101);
nor U373 (N_373,In_290,N_129);
nor U374 (N_374,In_100,N_272);
nor U375 (N_375,In_314,In_35);
or U376 (N_376,In_325,In_671);
and U377 (N_377,In_294,N_128);
nor U378 (N_378,N_287,In_553);
nor U379 (N_379,In_95,In_203);
and U380 (N_380,In_429,N_264);
nor U381 (N_381,In_271,In_655);
and U382 (N_382,In_566,N_198);
and U383 (N_383,N_168,In_178);
or U384 (N_384,In_542,In_418);
nand U385 (N_385,In_26,In_199);
nand U386 (N_386,In_44,In_708);
or U387 (N_387,In_637,In_404);
and U388 (N_388,N_216,N_289);
and U389 (N_389,In_163,N_280);
and U390 (N_390,In_7,In_695);
nor U391 (N_391,In_607,In_393);
or U392 (N_392,N_268,N_237);
and U393 (N_393,In_705,In_327);
or U394 (N_394,N_89,In_48);
nand U395 (N_395,In_254,N_141);
and U396 (N_396,In_610,In_131);
and U397 (N_397,In_307,In_97);
and U398 (N_398,In_309,In_261);
or U399 (N_399,In_227,In_641);
xnor U400 (N_400,N_397,N_352);
nor U401 (N_401,In_363,N_130);
nand U402 (N_402,In_181,In_690);
and U403 (N_403,In_385,N_234);
and U404 (N_404,In_657,N_242);
or U405 (N_405,N_176,N_70);
nand U406 (N_406,N_224,In_422);
nor U407 (N_407,N_381,N_341);
nand U408 (N_408,N_254,In_484);
nor U409 (N_409,N_326,In_486);
and U410 (N_410,N_310,In_578);
or U411 (N_411,N_383,In_111);
or U412 (N_412,In_745,In_577);
nor U413 (N_413,In_5,N_208);
and U414 (N_414,N_346,In_523);
nand U415 (N_415,N_304,In_180);
nand U416 (N_416,N_144,N_210);
nor U417 (N_417,N_282,In_52);
nor U418 (N_418,In_568,In_85);
xnor U419 (N_419,In_322,N_221);
and U420 (N_420,N_375,N_324);
and U421 (N_421,N_219,N_283);
or U422 (N_422,N_399,N_46);
or U423 (N_423,In_120,N_243);
nor U424 (N_424,N_371,In_516);
and U425 (N_425,N_207,In_625);
nand U426 (N_426,N_396,In_258);
or U427 (N_427,In_367,N_3);
and U428 (N_428,N_154,N_306);
nand U429 (N_429,In_288,In_143);
or U430 (N_430,N_235,In_79);
xor U431 (N_431,N_300,In_78);
nor U432 (N_432,In_216,N_388);
nor U433 (N_433,N_328,N_211);
and U434 (N_434,N_281,N_58);
nor U435 (N_435,N_350,N_333);
and U436 (N_436,In_267,In_660);
or U437 (N_437,N_329,In_224);
or U438 (N_438,In_459,In_320);
nand U439 (N_439,N_33,In_504);
nor U440 (N_440,In_253,In_720);
nor U441 (N_441,In_220,In_139);
or U442 (N_442,In_631,In_713);
nor U443 (N_443,N_191,N_214);
and U444 (N_444,N_342,N_370);
or U445 (N_445,In_653,N_189);
or U446 (N_446,In_426,N_258);
and U447 (N_447,N_181,In_491);
and U448 (N_448,In_247,N_215);
nor U449 (N_449,N_245,N_316);
and U450 (N_450,N_238,In_345);
or U451 (N_451,In_235,N_295);
and U452 (N_452,N_265,N_137);
and U453 (N_453,N_159,In_420);
and U454 (N_454,N_285,N_49);
nor U455 (N_455,N_395,N_384);
or U456 (N_456,In_402,N_252);
nor U457 (N_457,N_368,N_311);
or U458 (N_458,N_291,N_379);
and U459 (N_459,N_355,N_363);
nand U460 (N_460,N_378,N_296);
and U461 (N_461,N_327,In_19);
or U462 (N_462,In_613,In_647);
nor U463 (N_463,N_394,N_147);
and U464 (N_464,N_41,N_344);
and U465 (N_465,N_376,In_34);
nor U466 (N_466,In_21,In_495);
and U467 (N_467,N_110,In_681);
nand U468 (N_468,N_331,In_445);
nor U469 (N_469,In_32,In_530);
nand U470 (N_470,In_94,In_148);
nor U471 (N_471,N_361,N_84);
and U472 (N_472,N_365,In_408);
nand U473 (N_473,N_332,In_585);
and U474 (N_474,N_248,In_453);
nor U475 (N_475,N_294,In_260);
or U476 (N_476,N_380,In_321);
nand U477 (N_477,N_357,In_600);
or U478 (N_478,N_241,In_444);
or U479 (N_479,N_107,N_323);
nand U480 (N_480,In_549,In_190);
and U481 (N_481,N_318,In_194);
or U482 (N_482,In_16,In_403);
nor U483 (N_483,In_522,N_330);
xor U484 (N_484,N_48,In_340);
nor U485 (N_485,In_712,In_56);
nor U486 (N_486,N_37,In_136);
and U487 (N_487,In_514,N_391);
nor U488 (N_488,N_226,N_362);
and U489 (N_489,N_247,In_179);
or U490 (N_490,N_203,In_39);
or U491 (N_491,N_367,In_438);
or U492 (N_492,N_301,N_69);
nor U493 (N_493,N_322,N_100);
and U494 (N_494,N_385,N_313);
xnor U495 (N_495,N_133,In_703);
nor U496 (N_496,N_348,In_279);
or U497 (N_497,N_276,In_333);
nor U498 (N_498,In_15,N_269);
or U499 (N_499,N_257,N_319);
nand U500 (N_500,N_495,N_484);
nor U501 (N_501,N_404,N_201);
nor U502 (N_502,N_356,N_456);
nand U503 (N_503,N_443,N_2);
nand U504 (N_504,N_123,N_489);
or U505 (N_505,In_90,N_413);
or U506 (N_506,In_2,N_433);
or U507 (N_507,N_460,N_492);
or U508 (N_508,N_421,N_434);
or U509 (N_509,N_266,N_497);
and U510 (N_510,In_419,N_366);
and U511 (N_511,In_696,N_249);
nor U512 (N_512,N_354,N_390);
and U513 (N_513,N_482,N_436);
or U514 (N_514,N_455,N_451);
or U515 (N_515,N_25,N_167);
nand U516 (N_516,N_372,N_307);
or U517 (N_517,N_425,N_427);
nor U518 (N_518,In_183,N_373);
nor U519 (N_519,N_479,N_473);
nor U520 (N_520,In_692,N_317);
or U521 (N_521,N_345,N_297);
or U522 (N_522,N_418,In_686);
and U523 (N_523,In_195,N_52);
nand U524 (N_524,In_682,In_726);
nand U525 (N_525,N_481,In_125);
xor U526 (N_526,N_173,N_448);
or U527 (N_527,N_314,N_93);
or U528 (N_528,N_449,N_308);
nor U529 (N_529,N_465,N_398);
or U530 (N_530,In_373,N_335);
and U531 (N_531,N_312,In_145);
xnor U532 (N_532,N_431,N_321);
nand U533 (N_533,In_443,N_486);
or U534 (N_534,N_114,In_619);
or U535 (N_535,N_491,N_240);
and U536 (N_536,N_411,N_454);
and U537 (N_537,N_469,In_242);
or U538 (N_538,N_415,N_416);
nand U539 (N_539,In_350,N_461);
xor U540 (N_540,N_420,N_369);
and U541 (N_541,N_259,N_472);
and U542 (N_542,N_102,In_710);
xor U543 (N_543,N_468,N_403);
and U544 (N_544,N_477,N_17);
and U545 (N_545,N_470,N_442);
xor U546 (N_546,In_289,N_374);
nor U547 (N_547,N_325,N_359);
nand U548 (N_548,N_457,N_409);
and U549 (N_549,In_744,N_377);
nor U550 (N_550,N_498,N_62);
and U551 (N_551,N_334,N_494);
nand U552 (N_552,In_605,N_464);
nand U553 (N_553,N_315,N_32);
nand U554 (N_554,N_445,N_126);
nor U555 (N_555,N_336,N_302);
nand U556 (N_556,N_410,In_175);
xnor U557 (N_557,N_419,N_408);
and U558 (N_558,In_182,N_286);
or U559 (N_559,In_650,N_422);
nor U560 (N_560,N_347,In_526);
nor U561 (N_561,N_358,N_309);
nor U562 (N_562,N_204,N_490);
nor U563 (N_563,N_429,N_222);
or U564 (N_564,In_8,N_441);
nand U565 (N_565,N_220,N_320);
and U566 (N_566,N_386,N_86);
or U567 (N_567,N_496,N_424);
or U568 (N_568,N_279,N_438);
and U569 (N_569,N_156,In_701);
and U570 (N_570,N_459,N_205);
nor U571 (N_571,N_471,N_343);
xor U572 (N_572,N_485,N_349);
or U573 (N_573,In_188,N_262);
and U574 (N_574,N_351,In_334);
nand U575 (N_575,N_406,N_423);
and U576 (N_576,N_303,N_253);
nand U577 (N_577,In_649,In_171);
or U578 (N_578,N_402,In_384);
nand U579 (N_579,In_724,N_483);
nand U580 (N_580,N_338,N_499);
nor U581 (N_581,In_721,N_475);
and U582 (N_582,N_467,N_393);
or U583 (N_583,N_145,N_78);
nand U584 (N_584,In_706,N_426);
nand U585 (N_585,N_476,N_488);
nor U586 (N_586,N_439,N_432);
nand U587 (N_587,N_462,N_487);
nor U588 (N_588,N_382,N_288);
nor U589 (N_589,In_590,N_271);
or U590 (N_590,N_246,N_353);
or U591 (N_591,In_401,N_199);
nor U592 (N_592,In_154,N_437);
and U593 (N_593,N_453,N_447);
or U594 (N_594,N_184,N_435);
or U595 (N_595,N_131,N_200);
or U596 (N_596,N_392,In_277);
or U597 (N_597,N_163,In_357);
or U598 (N_598,In_266,N_186);
xor U599 (N_599,N_405,N_270);
or U600 (N_600,N_444,N_533);
or U601 (N_601,N_562,N_571);
nand U602 (N_602,N_579,In_740);
or U603 (N_603,N_510,N_480);
and U604 (N_604,N_599,N_507);
nor U605 (N_605,N_535,N_231);
and U606 (N_606,N_466,N_505);
xor U607 (N_607,N_517,N_587);
or U608 (N_608,N_519,N_594);
nand U609 (N_609,N_576,N_589);
or U610 (N_610,N_563,N_474);
and U611 (N_611,N_440,N_229);
nor U612 (N_612,N_387,N_545);
or U613 (N_613,N_592,N_588);
and U614 (N_614,N_565,N_400);
or U615 (N_615,N_578,N_339);
and U616 (N_616,N_478,N_572);
or U617 (N_617,N_506,N_417);
nand U618 (N_618,N_514,N_178);
and U619 (N_619,N_598,N_596);
nor U620 (N_620,N_458,N_539);
and U621 (N_621,N_98,N_573);
nor U622 (N_622,N_452,N_570);
or U623 (N_623,N_305,N_566);
nand U624 (N_624,N_554,N_340);
nand U625 (N_625,In_399,N_575);
and U626 (N_626,N_556,N_593);
nor U627 (N_627,In_501,N_538);
and U628 (N_628,N_299,N_559);
or U629 (N_629,N_450,N_597);
nand U630 (N_630,N_568,N_548);
nand U631 (N_631,N_513,N_508);
and U632 (N_632,N_511,N_407);
xnor U633 (N_633,N_529,N_537);
and U634 (N_634,N_504,N_564);
or U635 (N_635,N_549,N_560);
nor U636 (N_636,N_590,N_15);
nor U637 (N_637,N_503,N_515);
and U638 (N_638,N_223,N_512);
nor U639 (N_639,N_581,N_463);
nand U640 (N_640,N_502,N_557);
or U641 (N_641,N_547,N_277);
or U642 (N_642,N_567,N_561);
or U643 (N_643,N_520,N_528);
or U644 (N_644,N_574,N_428);
or U645 (N_645,N_360,N_516);
nand U646 (N_646,N_532,N_555);
and U647 (N_647,N_584,N_364);
nand U648 (N_648,N_293,N_522);
and U649 (N_649,N_412,In_155);
or U650 (N_650,N_558,N_172);
or U651 (N_651,N_544,N_540);
or U652 (N_652,In_416,N_583);
nor U653 (N_653,N_531,N_518);
nand U654 (N_654,N_275,N_534);
and U655 (N_655,N_553,N_526);
nand U656 (N_656,N_530,N_580);
nor U657 (N_657,N_541,N_525);
and U658 (N_658,N_523,N_582);
and U659 (N_659,N_278,N_509);
or U660 (N_660,N_595,N_521);
nand U661 (N_661,N_546,N_536);
and U662 (N_662,N_552,N_501);
and U663 (N_663,N_569,N_414);
nand U664 (N_664,N_551,N_493);
nand U665 (N_665,N_446,N_527);
nand U666 (N_666,N_430,N_550);
nand U667 (N_667,N_233,N_401);
or U668 (N_668,N_337,N_585);
or U669 (N_669,N_542,N_524);
and U670 (N_670,N_19,N_543);
and U671 (N_671,N_591,N_95);
or U672 (N_672,In_140,N_577);
nand U673 (N_673,N_500,N_0);
nor U674 (N_674,N_586,N_389);
and U675 (N_675,N_563,N_580);
xor U676 (N_676,N_542,N_523);
nand U677 (N_677,N_493,N_450);
nand U678 (N_678,N_172,N_530);
nand U679 (N_679,N_231,N_517);
nor U680 (N_680,N_564,N_532);
and U681 (N_681,N_360,N_541);
nand U682 (N_682,N_511,N_588);
and U683 (N_683,N_229,N_430);
and U684 (N_684,N_531,N_574);
or U685 (N_685,N_544,N_560);
nor U686 (N_686,N_561,N_571);
or U687 (N_687,N_233,N_520);
nand U688 (N_688,N_531,N_458);
nand U689 (N_689,N_535,N_518);
or U690 (N_690,N_278,N_596);
or U691 (N_691,N_360,N_517);
nor U692 (N_692,N_587,N_567);
and U693 (N_693,N_521,N_293);
nor U694 (N_694,N_553,N_528);
or U695 (N_695,N_569,N_474);
and U696 (N_696,N_545,N_507);
nor U697 (N_697,N_539,N_552);
and U698 (N_698,N_584,N_586);
or U699 (N_699,N_520,N_527);
or U700 (N_700,N_638,N_639);
nand U701 (N_701,N_689,N_674);
nand U702 (N_702,N_643,N_655);
nand U703 (N_703,N_677,N_679);
or U704 (N_704,N_640,N_605);
or U705 (N_705,N_635,N_630);
or U706 (N_706,N_632,N_671);
nor U707 (N_707,N_682,N_610);
nand U708 (N_708,N_628,N_603);
and U709 (N_709,N_623,N_668);
nand U710 (N_710,N_654,N_684);
and U711 (N_711,N_685,N_606);
and U712 (N_712,N_670,N_613);
or U713 (N_713,N_645,N_680);
nand U714 (N_714,N_612,N_622);
and U715 (N_715,N_694,N_667);
or U716 (N_716,N_699,N_600);
nand U717 (N_717,N_618,N_690);
nand U718 (N_718,N_659,N_678);
or U719 (N_719,N_616,N_681);
and U720 (N_720,N_601,N_625);
or U721 (N_721,N_697,N_649);
nor U722 (N_722,N_661,N_698);
or U723 (N_723,N_693,N_626);
or U724 (N_724,N_609,N_656);
and U725 (N_725,N_683,N_675);
or U726 (N_726,N_687,N_664);
nor U727 (N_727,N_663,N_627);
and U728 (N_728,N_669,N_629);
and U729 (N_729,N_686,N_644);
and U730 (N_730,N_617,N_647);
and U731 (N_731,N_620,N_633);
nor U732 (N_732,N_657,N_653);
nor U733 (N_733,N_666,N_652);
and U734 (N_734,N_695,N_676);
nand U735 (N_735,N_641,N_611);
nand U736 (N_736,N_621,N_692);
nor U737 (N_737,N_608,N_624);
nand U738 (N_738,N_646,N_665);
nor U739 (N_739,N_688,N_602);
and U740 (N_740,N_607,N_614);
nand U741 (N_741,N_651,N_637);
nand U742 (N_742,N_691,N_658);
nand U743 (N_743,N_636,N_619);
or U744 (N_744,N_615,N_696);
nor U745 (N_745,N_673,N_672);
xor U746 (N_746,N_642,N_662);
or U747 (N_747,N_634,N_650);
nand U748 (N_748,N_604,N_660);
nor U749 (N_749,N_648,N_631);
xor U750 (N_750,N_669,N_691);
and U751 (N_751,N_628,N_625);
and U752 (N_752,N_696,N_650);
or U753 (N_753,N_620,N_692);
or U754 (N_754,N_630,N_626);
nand U755 (N_755,N_666,N_615);
and U756 (N_756,N_602,N_665);
or U757 (N_757,N_605,N_636);
or U758 (N_758,N_678,N_677);
and U759 (N_759,N_654,N_668);
nor U760 (N_760,N_651,N_676);
or U761 (N_761,N_680,N_627);
and U762 (N_762,N_649,N_693);
nor U763 (N_763,N_681,N_662);
or U764 (N_764,N_629,N_654);
xor U765 (N_765,N_650,N_635);
nand U766 (N_766,N_667,N_657);
nor U767 (N_767,N_692,N_631);
and U768 (N_768,N_619,N_677);
nand U769 (N_769,N_653,N_609);
nor U770 (N_770,N_628,N_665);
nand U771 (N_771,N_633,N_655);
or U772 (N_772,N_691,N_682);
nand U773 (N_773,N_678,N_613);
nor U774 (N_774,N_679,N_681);
nand U775 (N_775,N_622,N_634);
nand U776 (N_776,N_639,N_674);
or U777 (N_777,N_633,N_696);
and U778 (N_778,N_604,N_681);
or U779 (N_779,N_608,N_676);
nor U780 (N_780,N_692,N_681);
or U781 (N_781,N_681,N_695);
or U782 (N_782,N_652,N_609);
nor U783 (N_783,N_608,N_671);
or U784 (N_784,N_694,N_684);
and U785 (N_785,N_628,N_614);
xor U786 (N_786,N_675,N_657);
and U787 (N_787,N_679,N_641);
nand U788 (N_788,N_660,N_653);
nand U789 (N_789,N_675,N_603);
or U790 (N_790,N_661,N_656);
nand U791 (N_791,N_631,N_632);
nor U792 (N_792,N_635,N_691);
or U793 (N_793,N_613,N_614);
or U794 (N_794,N_606,N_674);
and U795 (N_795,N_641,N_671);
nand U796 (N_796,N_616,N_628);
nor U797 (N_797,N_619,N_667);
nor U798 (N_798,N_643,N_666);
nand U799 (N_799,N_639,N_630);
and U800 (N_800,N_778,N_780);
nor U801 (N_801,N_706,N_797);
nor U802 (N_802,N_701,N_725);
nor U803 (N_803,N_720,N_791);
or U804 (N_804,N_790,N_746);
nand U805 (N_805,N_742,N_789);
nand U806 (N_806,N_728,N_748);
nand U807 (N_807,N_755,N_765);
or U808 (N_808,N_783,N_710);
and U809 (N_809,N_731,N_771);
nand U810 (N_810,N_732,N_786);
and U811 (N_811,N_757,N_722);
nor U812 (N_812,N_747,N_704);
and U813 (N_813,N_711,N_781);
nor U814 (N_814,N_730,N_772);
or U815 (N_815,N_712,N_719);
nand U816 (N_816,N_792,N_705);
or U817 (N_817,N_773,N_759);
and U818 (N_818,N_727,N_702);
nand U819 (N_819,N_767,N_793);
nand U820 (N_820,N_751,N_799);
and U821 (N_821,N_738,N_735);
nor U822 (N_822,N_745,N_777);
nand U823 (N_823,N_794,N_788);
or U824 (N_824,N_784,N_779);
or U825 (N_825,N_769,N_774);
or U826 (N_826,N_764,N_775);
nand U827 (N_827,N_734,N_796);
nor U828 (N_828,N_721,N_770);
and U829 (N_829,N_750,N_707);
nand U830 (N_830,N_787,N_729);
and U831 (N_831,N_726,N_744);
nand U832 (N_832,N_737,N_753);
or U833 (N_833,N_782,N_762);
nand U834 (N_834,N_766,N_749);
and U835 (N_835,N_714,N_760);
nor U836 (N_836,N_700,N_763);
and U837 (N_837,N_733,N_752);
or U838 (N_838,N_716,N_724);
nor U839 (N_839,N_776,N_758);
or U840 (N_840,N_715,N_708);
nor U841 (N_841,N_785,N_736);
and U842 (N_842,N_795,N_740);
and U843 (N_843,N_754,N_739);
xor U844 (N_844,N_756,N_768);
nand U845 (N_845,N_717,N_709);
or U846 (N_846,N_723,N_741);
nand U847 (N_847,N_761,N_713);
and U848 (N_848,N_703,N_743);
or U849 (N_849,N_718,N_798);
nor U850 (N_850,N_792,N_794);
nor U851 (N_851,N_737,N_762);
or U852 (N_852,N_713,N_722);
nor U853 (N_853,N_727,N_755);
or U854 (N_854,N_779,N_729);
nor U855 (N_855,N_718,N_788);
and U856 (N_856,N_757,N_747);
and U857 (N_857,N_740,N_756);
nand U858 (N_858,N_706,N_747);
nor U859 (N_859,N_785,N_749);
nor U860 (N_860,N_722,N_786);
nor U861 (N_861,N_745,N_722);
xor U862 (N_862,N_755,N_772);
and U863 (N_863,N_763,N_706);
and U864 (N_864,N_724,N_745);
or U865 (N_865,N_746,N_715);
or U866 (N_866,N_778,N_785);
and U867 (N_867,N_710,N_797);
and U868 (N_868,N_744,N_742);
nor U869 (N_869,N_790,N_717);
or U870 (N_870,N_707,N_731);
nor U871 (N_871,N_734,N_798);
or U872 (N_872,N_729,N_762);
nand U873 (N_873,N_726,N_747);
and U874 (N_874,N_782,N_774);
nand U875 (N_875,N_792,N_740);
and U876 (N_876,N_705,N_797);
and U877 (N_877,N_751,N_725);
nand U878 (N_878,N_750,N_745);
or U879 (N_879,N_757,N_751);
and U880 (N_880,N_739,N_769);
or U881 (N_881,N_752,N_757);
and U882 (N_882,N_752,N_779);
and U883 (N_883,N_794,N_742);
and U884 (N_884,N_752,N_754);
or U885 (N_885,N_709,N_786);
nand U886 (N_886,N_705,N_760);
or U887 (N_887,N_716,N_766);
nor U888 (N_888,N_739,N_761);
and U889 (N_889,N_742,N_773);
nand U890 (N_890,N_743,N_793);
nor U891 (N_891,N_784,N_738);
or U892 (N_892,N_718,N_764);
and U893 (N_893,N_790,N_723);
or U894 (N_894,N_713,N_740);
and U895 (N_895,N_752,N_724);
and U896 (N_896,N_776,N_726);
nand U897 (N_897,N_750,N_731);
or U898 (N_898,N_700,N_766);
or U899 (N_899,N_709,N_756);
nand U900 (N_900,N_892,N_840);
nand U901 (N_901,N_895,N_877);
and U902 (N_902,N_819,N_807);
and U903 (N_903,N_845,N_881);
and U904 (N_904,N_891,N_854);
or U905 (N_905,N_883,N_841);
nor U906 (N_906,N_843,N_823);
or U907 (N_907,N_830,N_880);
nand U908 (N_908,N_878,N_848);
nor U909 (N_909,N_821,N_802);
nand U910 (N_910,N_827,N_865);
and U911 (N_911,N_837,N_875);
or U912 (N_912,N_871,N_805);
nand U913 (N_913,N_868,N_894);
nor U914 (N_914,N_859,N_818);
or U915 (N_915,N_814,N_851);
or U916 (N_916,N_857,N_835);
or U917 (N_917,N_867,N_898);
nand U918 (N_918,N_817,N_862);
or U919 (N_919,N_864,N_809);
and U920 (N_920,N_801,N_844);
nand U921 (N_921,N_842,N_800);
nor U922 (N_922,N_828,N_869);
or U923 (N_923,N_824,N_873);
nor U924 (N_924,N_803,N_889);
or U925 (N_925,N_806,N_861);
nor U926 (N_926,N_850,N_872);
or U927 (N_927,N_884,N_808);
and U928 (N_928,N_888,N_887);
or U929 (N_929,N_822,N_893);
nand U930 (N_930,N_846,N_874);
or U931 (N_931,N_813,N_882);
nand U932 (N_932,N_826,N_886);
or U933 (N_933,N_834,N_863);
or U934 (N_934,N_812,N_829);
nor U935 (N_935,N_815,N_896);
nor U936 (N_936,N_879,N_885);
nand U937 (N_937,N_866,N_833);
nand U938 (N_938,N_860,N_839);
nor U939 (N_939,N_820,N_897);
or U940 (N_940,N_852,N_853);
nand U941 (N_941,N_838,N_810);
or U942 (N_942,N_890,N_804);
nor U943 (N_943,N_858,N_849);
nor U944 (N_944,N_832,N_870);
nor U945 (N_945,N_825,N_876);
and U946 (N_946,N_816,N_847);
nand U947 (N_947,N_811,N_831);
nor U948 (N_948,N_836,N_856);
and U949 (N_949,N_855,N_899);
or U950 (N_950,N_819,N_811);
or U951 (N_951,N_895,N_822);
or U952 (N_952,N_811,N_868);
or U953 (N_953,N_879,N_878);
nor U954 (N_954,N_893,N_888);
or U955 (N_955,N_844,N_881);
nor U956 (N_956,N_806,N_814);
and U957 (N_957,N_861,N_839);
or U958 (N_958,N_859,N_887);
and U959 (N_959,N_836,N_859);
or U960 (N_960,N_890,N_818);
or U961 (N_961,N_862,N_863);
nor U962 (N_962,N_889,N_824);
nand U963 (N_963,N_825,N_885);
nor U964 (N_964,N_844,N_856);
and U965 (N_965,N_853,N_891);
and U966 (N_966,N_874,N_894);
and U967 (N_967,N_885,N_808);
nand U968 (N_968,N_841,N_869);
and U969 (N_969,N_827,N_866);
and U970 (N_970,N_858,N_828);
or U971 (N_971,N_833,N_811);
nor U972 (N_972,N_853,N_825);
or U973 (N_973,N_805,N_809);
or U974 (N_974,N_850,N_857);
and U975 (N_975,N_878,N_802);
and U976 (N_976,N_875,N_832);
nand U977 (N_977,N_800,N_817);
nor U978 (N_978,N_868,N_826);
nand U979 (N_979,N_881,N_874);
or U980 (N_980,N_826,N_816);
nand U981 (N_981,N_820,N_880);
or U982 (N_982,N_858,N_899);
and U983 (N_983,N_872,N_832);
nand U984 (N_984,N_863,N_867);
and U985 (N_985,N_837,N_866);
and U986 (N_986,N_854,N_819);
nand U987 (N_987,N_883,N_836);
or U988 (N_988,N_834,N_892);
xnor U989 (N_989,N_894,N_828);
or U990 (N_990,N_841,N_800);
or U991 (N_991,N_853,N_863);
or U992 (N_992,N_802,N_842);
and U993 (N_993,N_871,N_876);
nor U994 (N_994,N_835,N_846);
nor U995 (N_995,N_862,N_864);
nand U996 (N_996,N_802,N_875);
and U997 (N_997,N_811,N_890);
nor U998 (N_998,N_884,N_881);
nor U999 (N_999,N_800,N_863);
nor U1000 (N_1000,N_969,N_935);
or U1001 (N_1001,N_987,N_955);
or U1002 (N_1002,N_981,N_925);
or U1003 (N_1003,N_929,N_906);
and U1004 (N_1004,N_932,N_985);
nor U1005 (N_1005,N_909,N_976);
nor U1006 (N_1006,N_951,N_933);
and U1007 (N_1007,N_954,N_992);
nand U1008 (N_1008,N_936,N_924);
and U1009 (N_1009,N_953,N_904);
and U1010 (N_1010,N_916,N_996);
nand U1011 (N_1011,N_957,N_959);
or U1012 (N_1012,N_999,N_977);
or U1013 (N_1013,N_973,N_901);
and U1014 (N_1014,N_905,N_980);
or U1015 (N_1015,N_967,N_910);
and U1016 (N_1016,N_920,N_934);
or U1017 (N_1017,N_979,N_918);
or U1018 (N_1018,N_900,N_983);
nand U1019 (N_1019,N_968,N_937);
nor U1020 (N_1020,N_972,N_902);
and U1021 (N_1021,N_989,N_990);
nand U1022 (N_1022,N_911,N_956);
and U1023 (N_1023,N_944,N_962);
or U1024 (N_1024,N_913,N_988);
xor U1025 (N_1025,N_993,N_961);
xnor U1026 (N_1026,N_966,N_942);
nand U1027 (N_1027,N_915,N_919);
nor U1028 (N_1028,N_970,N_971);
nor U1029 (N_1029,N_998,N_914);
or U1030 (N_1030,N_926,N_921);
or U1031 (N_1031,N_931,N_994);
or U1032 (N_1032,N_917,N_948);
and U1033 (N_1033,N_938,N_952);
and U1034 (N_1034,N_941,N_986);
nand U1035 (N_1035,N_995,N_958);
or U1036 (N_1036,N_949,N_982);
nand U1037 (N_1037,N_991,N_903);
or U1038 (N_1038,N_965,N_912);
or U1039 (N_1039,N_943,N_927);
nor U1040 (N_1040,N_947,N_930);
nor U1041 (N_1041,N_974,N_946);
nor U1042 (N_1042,N_908,N_964);
nor U1043 (N_1043,N_997,N_923);
nand U1044 (N_1044,N_939,N_928);
nor U1045 (N_1045,N_940,N_907);
and U1046 (N_1046,N_960,N_922);
nor U1047 (N_1047,N_978,N_963);
nand U1048 (N_1048,N_975,N_945);
or U1049 (N_1049,N_984,N_950);
nand U1050 (N_1050,N_941,N_939);
or U1051 (N_1051,N_902,N_983);
nand U1052 (N_1052,N_976,N_985);
xor U1053 (N_1053,N_912,N_955);
nor U1054 (N_1054,N_917,N_985);
nand U1055 (N_1055,N_901,N_907);
nand U1056 (N_1056,N_976,N_953);
and U1057 (N_1057,N_923,N_966);
and U1058 (N_1058,N_954,N_955);
and U1059 (N_1059,N_938,N_931);
and U1060 (N_1060,N_996,N_930);
nor U1061 (N_1061,N_944,N_915);
nor U1062 (N_1062,N_900,N_992);
xor U1063 (N_1063,N_992,N_951);
and U1064 (N_1064,N_932,N_961);
nor U1065 (N_1065,N_926,N_983);
nor U1066 (N_1066,N_976,N_906);
or U1067 (N_1067,N_986,N_909);
nand U1068 (N_1068,N_933,N_937);
nand U1069 (N_1069,N_950,N_952);
or U1070 (N_1070,N_984,N_956);
and U1071 (N_1071,N_932,N_951);
or U1072 (N_1072,N_960,N_954);
nor U1073 (N_1073,N_959,N_903);
nor U1074 (N_1074,N_992,N_934);
or U1075 (N_1075,N_906,N_975);
or U1076 (N_1076,N_996,N_962);
nand U1077 (N_1077,N_910,N_983);
nor U1078 (N_1078,N_966,N_958);
nor U1079 (N_1079,N_979,N_941);
nand U1080 (N_1080,N_981,N_928);
nor U1081 (N_1081,N_925,N_997);
nor U1082 (N_1082,N_904,N_926);
nand U1083 (N_1083,N_932,N_939);
or U1084 (N_1084,N_940,N_993);
nand U1085 (N_1085,N_939,N_921);
and U1086 (N_1086,N_937,N_930);
nor U1087 (N_1087,N_931,N_947);
and U1088 (N_1088,N_949,N_905);
or U1089 (N_1089,N_927,N_969);
nand U1090 (N_1090,N_963,N_925);
nand U1091 (N_1091,N_923,N_963);
and U1092 (N_1092,N_992,N_945);
nor U1093 (N_1093,N_949,N_918);
and U1094 (N_1094,N_943,N_956);
nand U1095 (N_1095,N_999,N_983);
or U1096 (N_1096,N_900,N_979);
nand U1097 (N_1097,N_992,N_903);
nor U1098 (N_1098,N_945,N_977);
nor U1099 (N_1099,N_991,N_964);
nor U1100 (N_1100,N_1086,N_1018);
and U1101 (N_1101,N_1071,N_1041);
or U1102 (N_1102,N_1051,N_1052);
nor U1103 (N_1103,N_1077,N_1056);
nor U1104 (N_1104,N_1045,N_1053);
nor U1105 (N_1105,N_1088,N_1002);
and U1106 (N_1106,N_1063,N_1027);
nand U1107 (N_1107,N_1044,N_1000);
and U1108 (N_1108,N_1016,N_1080);
and U1109 (N_1109,N_1098,N_1050);
or U1110 (N_1110,N_1039,N_1046);
and U1111 (N_1111,N_1065,N_1078);
and U1112 (N_1112,N_1087,N_1031);
nor U1113 (N_1113,N_1008,N_1007);
nand U1114 (N_1114,N_1014,N_1021);
nor U1115 (N_1115,N_1054,N_1067);
nand U1116 (N_1116,N_1010,N_1048);
nand U1117 (N_1117,N_1062,N_1025);
or U1118 (N_1118,N_1064,N_1058);
and U1119 (N_1119,N_1072,N_1042);
or U1120 (N_1120,N_1057,N_1012);
or U1121 (N_1121,N_1020,N_1081);
and U1122 (N_1122,N_1040,N_1099);
nand U1123 (N_1123,N_1076,N_1089);
nand U1124 (N_1124,N_1022,N_1090);
nor U1125 (N_1125,N_1017,N_1096);
or U1126 (N_1126,N_1084,N_1037);
and U1127 (N_1127,N_1055,N_1033);
or U1128 (N_1128,N_1030,N_1034);
nor U1129 (N_1129,N_1068,N_1036);
and U1130 (N_1130,N_1061,N_1085);
or U1131 (N_1131,N_1083,N_1097);
nor U1132 (N_1132,N_1035,N_1092);
and U1133 (N_1133,N_1079,N_1006);
or U1134 (N_1134,N_1093,N_1013);
nor U1135 (N_1135,N_1059,N_1009);
or U1136 (N_1136,N_1026,N_1032);
nor U1137 (N_1137,N_1011,N_1019);
or U1138 (N_1138,N_1075,N_1003);
and U1139 (N_1139,N_1015,N_1047);
and U1140 (N_1140,N_1069,N_1091);
and U1141 (N_1141,N_1038,N_1023);
nand U1142 (N_1142,N_1073,N_1070);
nor U1143 (N_1143,N_1060,N_1043);
nor U1144 (N_1144,N_1074,N_1049);
nand U1145 (N_1145,N_1029,N_1001);
and U1146 (N_1146,N_1066,N_1028);
and U1147 (N_1147,N_1024,N_1095);
or U1148 (N_1148,N_1094,N_1004);
or U1149 (N_1149,N_1082,N_1005);
nor U1150 (N_1150,N_1028,N_1085);
nor U1151 (N_1151,N_1003,N_1027);
nand U1152 (N_1152,N_1046,N_1035);
or U1153 (N_1153,N_1002,N_1070);
nand U1154 (N_1154,N_1045,N_1036);
and U1155 (N_1155,N_1002,N_1044);
xor U1156 (N_1156,N_1026,N_1030);
nand U1157 (N_1157,N_1017,N_1073);
or U1158 (N_1158,N_1031,N_1028);
or U1159 (N_1159,N_1090,N_1081);
nand U1160 (N_1160,N_1083,N_1056);
xnor U1161 (N_1161,N_1080,N_1073);
and U1162 (N_1162,N_1003,N_1061);
or U1163 (N_1163,N_1073,N_1003);
and U1164 (N_1164,N_1088,N_1012);
or U1165 (N_1165,N_1015,N_1086);
or U1166 (N_1166,N_1032,N_1094);
xnor U1167 (N_1167,N_1046,N_1088);
and U1168 (N_1168,N_1002,N_1096);
or U1169 (N_1169,N_1037,N_1020);
nand U1170 (N_1170,N_1005,N_1027);
or U1171 (N_1171,N_1004,N_1006);
nand U1172 (N_1172,N_1074,N_1040);
nor U1173 (N_1173,N_1053,N_1036);
nand U1174 (N_1174,N_1042,N_1064);
or U1175 (N_1175,N_1093,N_1001);
and U1176 (N_1176,N_1012,N_1008);
nor U1177 (N_1177,N_1046,N_1017);
nand U1178 (N_1178,N_1005,N_1095);
and U1179 (N_1179,N_1085,N_1044);
nand U1180 (N_1180,N_1042,N_1039);
and U1181 (N_1181,N_1013,N_1043);
nand U1182 (N_1182,N_1099,N_1089);
or U1183 (N_1183,N_1025,N_1055);
nand U1184 (N_1184,N_1089,N_1034);
nand U1185 (N_1185,N_1049,N_1010);
nand U1186 (N_1186,N_1007,N_1001);
nand U1187 (N_1187,N_1046,N_1036);
and U1188 (N_1188,N_1093,N_1007);
and U1189 (N_1189,N_1038,N_1053);
nor U1190 (N_1190,N_1045,N_1085);
and U1191 (N_1191,N_1032,N_1065);
nor U1192 (N_1192,N_1008,N_1086);
or U1193 (N_1193,N_1056,N_1005);
and U1194 (N_1194,N_1030,N_1051);
nand U1195 (N_1195,N_1062,N_1023);
and U1196 (N_1196,N_1065,N_1051);
nor U1197 (N_1197,N_1088,N_1085);
or U1198 (N_1198,N_1003,N_1054);
and U1199 (N_1199,N_1073,N_1093);
nor U1200 (N_1200,N_1101,N_1108);
and U1201 (N_1201,N_1164,N_1111);
or U1202 (N_1202,N_1104,N_1151);
and U1203 (N_1203,N_1149,N_1117);
and U1204 (N_1204,N_1114,N_1129);
or U1205 (N_1205,N_1115,N_1178);
and U1206 (N_1206,N_1126,N_1145);
nor U1207 (N_1207,N_1142,N_1130);
or U1208 (N_1208,N_1136,N_1156);
or U1209 (N_1209,N_1106,N_1181);
nor U1210 (N_1210,N_1155,N_1127);
or U1211 (N_1211,N_1121,N_1122);
nand U1212 (N_1212,N_1123,N_1184);
nor U1213 (N_1213,N_1144,N_1153);
nand U1214 (N_1214,N_1187,N_1163);
or U1215 (N_1215,N_1165,N_1138);
and U1216 (N_1216,N_1162,N_1119);
or U1217 (N_1217,N_1134,N_1190);
or U1218 (N_1218,N_1161,N_1135);
nand U1219 (N_1219,N_1159,N_1133);
nor U1220 (N_1220,N_1172,N_1176);
and U1221 (N_1221,N_1179,N_1139);
nor U1222 (N_1222,N_1197,N_1124);
nor U1223 (N_1223,N_1158,N_1180);
nor U1224 (N_1224,N_1198,N_1183);
nand U1225 (N_1225,N_1177,N_1107);
nand U1226 (N_1226,N_1175,N_1173);
nor U1227 (N_1227,N_1195,N_1116);
or U1228 (N_1228,N_1168,N_1199);
and U1229 (N_1229,N_1169,N_1102);
or U1230 (N_1230,N_1112,N_1157);
and U1231 (N_1231,N_1171,N_1191);
nor U1232 (N_1232,N_1167,N_1160);
nor U1233 (N_1233,N_1182,N_1125);
or U1234 (N_1234,N_1146,N_1189);
and U1235 (N_1235,N_1152,N_1137);
and U1236 (N_1236,N_1174,N_1140);
nor U1237 (N_1237,N_1110,N_1196);
and U1238 (N_1238,N_1188,N_1185);
nand U1239 (N_1239,N_1103,N_1143);
and U1240 (N_1240,N_1186,N_1193);
nand U1241 (N_1241,N_1113,N_1132);
nor U1242 (N_1242,N_1120,N_1194);
xor U1243 (N_1243,N_1166,N_1118);
nor U1244 (N_1244,N_1105,N_1131);
nand U1245 (N_1245,N_1148,N_1150);
nor U1246 (N_1246,N_1128,N_1192);
nor U1247 (N_1247,N_1170,N_1141);
nand U1248 (N_1248,N_1109,N_1100);
nand U1249 (N_1249,N_1154,N_1147);
or U1250 (N_1250,N_1124,N_1127);
nor U1251 (N_1251,N_1142,N_1101);
nand U1252 (N_1252,N_1125,N_1127);
or U1253 (N_1253,N_1130,N_1178);
or U1254 (N_1254,N_1128,N_1116);
xnor U1255 (N_1255,N_1105,N_1149);
or U1256 (N_1256,N_1190,N_1185);
or U1257 (N_1257,N_1185,N_1156);
nand U1258 (N_1258,N_1171,N_1199);
nand U1259 (N_1259,N_1151,N_1178);
or U1260 (N_1260,N_1174,N_1179);
nor U1261 (N_1261,N_1143,N_1181);
nor U1262 (N_1262,N_1172,N_1188);
nand U1263 (N_1263,N_1137,N_1101);
and U1264 (N_1264,N_1185,N_1119);
xnor U1265 (N_1265,N_1185,N_1145);
or U1266 (N_1266,N_1157,N_1143);
nand U1267 (N_1267,N_1187,N_1127);
nor U1268 (N_1268,N_1111,N_1178);
and U1269 (N_1269,N_1178,N_1169);
and U1270 (N_1270,N_1161,N_1153);
nor U1271 (N_1271,N_1104,N_1191);
or U1272 (N_1272,N_1121,N_1103);
and U1273 (N_1273,N_1196,N_1145);
nor U1274 (N_1274,N_1149,N_1168);
and U1275 (N_1275,N_1185,N_1144);
and U1276 (N_1276,N_1159,N_1142);
nand U1277 (N_1277,N_1160,N_1173);
nand U1278 (N_1278,N_1150,N_1156);
xnor U1279 (N_1279,N_1165,N_1195);
and U1280 (N_1280,N_1169,N_1172);
and U1281 (N_1281,N_1173,N_1108);
nand U1282 (N_1282,N_1110,N_1107);
or U1283 (N_1283,N_1151,N_1109);
and U1284 (N_1284,N_1194,N_1154);
or U1285 (N_1285,N_1169,N_1166);
nor U1286 (N_1286,N_1173,N_1168);
and U1287 (N_1287,N_1199,N_1105);
nand U1288 (N_1288,N_1157,N_1146);
and U1289 (N_1289,N_1186,N_1131);
nor U1290 (N_1290,N_1135,N_1148);
and U1291 (N_1291,N_1186,N_1142);
nor U1292 (N_1292,N_1199,N_1101);
or U1293 (N_1293,N_1151,N_1169);
nor U1294 (N_1294,N_1177,N_1164);
and U1295 (N_1295,N_1115,N_1170);
nor U1296 (N_1296,N_1185,N_1152);
nor U1297 (N_1297,N_1193,N_1149);
nor U1298 (N_1298,N_1186,N_1139);
nor U1299 (N_1299,N_1191,N_1173);
and U1300 (N_1300,N_1243,N_1212);
nand U1301 (N_1301,N_1277,N_1256);
nor U1302 (N_1302,N_1272,N_1262);
and U1303 (N_1303,N_1286,N_1244);
nor U1304 (N_1304,N_1213,N_1295);
and U1305 (N_1305,N_1293,N_1268);
nor U1306 (N_1306,N_1290,N_1205);
and U1307 (N_1307,N_1267,N_1201);
nor U1308 (N_1308,N_1279,N_1207);
or U1309 (N_1309,N_1206,N_1236);
or U1310 (N_1310,N_1219,N_1264);
xnor U1311 (N_1311,N_1276,N_1216);
xor U1312 (N_1312,N_1202,N_1273);
or U1313 (N_1313,N_1227,N_1237);
and U1314 (N_1314,N_1239,N_1281);
and U1315 (N_1315,N_1284,N_1250);
nor U1316 (N_1316,N_1231,N_1263);
nor U1317 (N_1317,N_1274,N_1208);
nor U1318 (N_1318,N_1278,N_1288);
and U1319 (N_1319,N_1291,N_1230);
or U1320 (N_1320,N_1215,N_1298);
nor U1321 (N_1321,N_1228,N_1257);
and U1322 (N_1322,N_1234,N_1283);
nand U1323 (N_1323,N_1204,N_1233);
and U1324 (N_1324,N_1265,N_1221);
xor U1325 (N_1325,N_1218,N_1299);
or U1326 (N_1326,N_1259,N_1220);
nand U1327 (N_1327,N_1240,N_1269);
or U1328 (N_1328,N_1280,N_1248);
nand U1329 (N_1329,N_1229,N_1200);
nand U1330 (N_1330,N_1238,N_1266);
nor U1331 (N_1331,N_1289,N_1211);
nor U1332 (N_1332,N_1292,N_1247);
and U1333 (N_1333,N_1214,N_1242);
and U1334 (N_1334,N_1210,N_1203);
and U1335 (N_1335,N_1285,N_1246);
and U1336 (N_1336,N_1225,N_1217);
or U1337 (N_1337,N_1271,N_1249);
or U1338 (N_1338,N_1245,N_1252);
and U1339 (N_1339,N_1209,N_1297);
and U1340 (N_1340,N_1235,N_1282);
and U1341 (N_1341,N_1223,N_1275);
nand U1342 (N_1342,N_1294,N_1224);
nand U1343 (N_1343,N_1270,N_1241);
or U1344 (N_1344,N_1222,N_1255);
and U1345 (N_1345,N_1258,N_1296);
or U1346 (N_1346,N_1260,N_1251);
or U1347 (N_1347,N_1232,N_1254);
nand U1348 (N_1348,N_1226,N_1261);
and U1349 (N_1349,N_1253,N_1287);
nand U1350 (N_1350,N_1204,N_1282);
or U1351 (N_1351,N_1217,N_1220);
nand U1352 (N_1352,N_1276,N_1288);
nor U1353 (N_1353,N_1227,N_1275);
and U1354 (N_1354,N_1202,N_1296);
or U1355 (N_1355,N_1235,N_1266);
or U1356 (N_1356,N_1211,N_1255);
nor U1357 (N_1357,N_1276,N_1231);
and U1358 (N_1358,N_1288,N_1292);
nand U1359 (N_1359,N_1276,N_1274);
or U1360 (N_1360,N_1236,N_1218);
nand U1361 (N_1361,N_1277,N_1239);
nand U1362 (N_1362,N_1222,N_1257);
and U1363 (N_1363,N_1298,N_1294);
and U1364 (N_1364,N_1264,N_1228);
or U1365 (N_1365,N_1299,N_1219);
and U1366 (N_1366,N_1297,N_1240);
or U1367 (N_1367,N_1235,N_1232);
nor U1368 (N_1368,N_1273,N_1236);
or U1369 (N_1369,N_1260,N_1206);
nand U1370 (N_1370,N_1218,N_1234);
xnor U1371 (N_1371,N_1242,N_1288);
and U1372 (N_1372,N_1206,N_1232);
nand U1373 (N_1373,N_1276,N_1277);
nor U1374 (N_1374,N_1297,N_1290);
xnor U1375 (N_1375,N_1265,N_1227);
nor U1376 (N_1376,N_1284,N_1225);
and U1377 (N_1377,N_1250,N_1230);
and U1378 (N_1378,N_1204,N_1205);
nand U1379 (N_1379,N_1266,N_1289);
or U1380 (N_1380,N_1252,N_1249);
nand U1381 (N_1381,N_1209,N_1288);
or U1382 (N_1382,N_1290,N_1226);
or U1383 (N_1383,N_1228,N_1223);
nor U1384 (N_1384,N_1221,N_1239);
nand U1385 (N_1385,N_1270,N_1257);
nor U1386 (N_1386,N_1275,N_1212);
nand U1387 (N_1387,N_1225,N_1259);
or U1388 (N_1388,N_1241,N_1254);
nand U1389 (N_1389,N_1206,N_1233);
and U1390 (N_1390,N_1213,N_1239);
and U1391 (N_1391,N_1289,N_1226);
and U1392 (N_1392,N_1205,N_1257);
and U1393 (N_1393,N_1286,N_1243);
nand U1394 (N_1394,N_1200,N_1236);
or U1395 (N_1395,N_1254,N_1296);
or U1396 (N_1396,N_1281,N_1217);
and U1397 (N_1397,N_1284,N_1206);
or U1398 (N_1398,N_1207,N_1212);
or U1399 (N_1399,N_1222,N_1218);
nand U1400 (N_1400,N_1394,N_1334);
or U1401 (N_1401,N_1356,N_1316);
nor U1402 (N_1402,N_1302,N_1392);
or U1403 (N_1403,N_1364,N_1352);
nor U1404 (N_1404,N_1330,N_1381);
and U1405 (N_1405,N_1388,N_1305);
xor U1406 (N_1406,N_1340,N_1345);
nand U1407 (N_1407,N_1375,N_1374);
and U1408 (N_1408,N_1353,N_1396);
nor U1409 (N_1409,N_1377,N_1313);
or U1410 (N_1410,N_1386,N_1303);
and U1411 (N_1411,N_1346,N_1398);
nand U1412 (N_1412,N_1342,N_1304);
or U1413 (N_1413,N_1309,N_1344);
xnor U1414 (N_1414,N_1339,N_1329);
nor U1415 (N_1415,N_1367,N_1378);
or U1416 (N_1416,N_1328,N_1358);
and U1417 (N_1417,N_1327,N_1371);
nor U1418 (N_1418,N_1369,N_1397);
and U1419 (N_1419,N_1372,N_1361);
nor U1420 (N_1420,N_1376,N_1382);
and U1421 (N_1421,N_1357,N_1387);
nor U1422 (N_1422,N_1399,N_1336);
or U1423 (N_1423,N_1337,N_1324);
or U1424 (N_1424,N_1354,N_1335);
and U1425 (N_1425,N_1366,N_1384);
nor U1426 (N_1426,N_1391,N_1379);
and U1427 (N_1427,N_1317,N_1355);
or U1428 (N_1428,N_1306,N_1314);
or U1429 (N_1429,N_1322,N_1311);
or U1430 (N_1430,N_1390,N_1307);
nand U1431 (N_1431,N_1321,N_1362);
nand U1432 (N_1432,N_1301,N_1373);
nand U1433 (N_1433,N_1347,N_1319);
and U1434 (N_1434,N_1318,N_1332);
nor U1435 (N_1435,N_1343,N_1333);
nand U1436 (N_1436,N_1351,N_1389);
nand U1437 (N_1437,N_1363,N_1383);
and U1438 (N_1438,N_1325,N_1308);
nand U1439 (N_1439,N_1300,N_1341);
and U1440 (N_1440,N_1380,N_1323);
nor U1441 (N_1441,N_1348,N_1365);
nor U1442 (N_1442,N_1331,N_1370);
nand U1443 (N_1443,N_1350,N_1320);
nor U1444 (N_1444,N_1338,N_1368);
and U1445 (N_1445,N_1395,N_1349);
nor U1446 (N_1446,N_1315,N_1393);
or U1447 (N_1447,N_1385,N_1360);
nor U1448 (N_1448,N_1359,N_1326);
and U1449 (N_1449,N_1312,N_1310);
nand U1450 (N_1450,N_1375,N_1367);
nor U1451 (N_1451,N_1371,N_1325);
or U1452 (N_1452,N_1393,N_1375);
and U1453 (N_1453,N_1321,N_1359);
and U1454 (N_1454,N_1391,N_1313);
xor U1455 (N_1455,N_1322,N_1371);
nand U1456 (N_1456,N_1311,N_1376);
nor U1457 (N_1457,N_1355,N_1378);
and U1458 (N_1458,N_1385,N_1309);
nand U1459 (N_1459,N_1306,N_1394);
and U1460 (N_1460,N_1310,N_1352);
nand U1461 (N_1461,N_1360,N_1398);
nand U1462 (N_1462,N_1383,N_1329);
nor U1463 (N_1463,N_1311,N_1333);
nor U1464 (N_1464,N_1350,N_1347);
nand U1465 (N_1465,N_1321,N_1378);
nand U1466 (N_1466,N_1308,N_1377);
nor U1467 (N_1467,N_1301,N_1309);
nor U1468 (N_1468,N_1303,N_1310);
and U1469 (N_1469,N_1350,N_1366);
nor U1470 (N_1470,N_1389,N_1358);
and U1471 (N_1471,N_1399,N_1389);
and U1472 (N_1472,N_1389,N_1319);
or U1473 (N_1473,N_1373,N_1337);
or U1474 (N_1474,N_1394,N_1337);
and U1475 (N_1475,N_1318,N_1387);
nand U1476 (N_1476,N_1357,N_1352);
nor U1477 (N_1477,N_1313,N_1390);
nand U1478 (N_1478,N_1324,N_1305);
nor U1479 (N_1479,N_1387,N_1378);
nor U1480 (N_1480,N_1325,N_1346);
and U1481 (N_1481,N_1329,N_1372);
nor U1482 (N_1482,N_1326,N_1394);
and U1483 (N_1483,N_1322,N_1397);
or U1484 (N_1484,N_1370,N_1373);
nor U1485 (N_1485,N_1352,N_1321);
nand U1486 (N_1486,N_1359,N_1302);
nor U1487 (N_1487,N_1331,N_1318);
nand U1488 (N_1488,N_1329,N_1314);
and U1489 (N_1489,N_1343,N_1366);
nor U1490 (N_1490,N_1375,N_1356);
and U1491 (N_1491,N_1382,N_1352);
or U1492 (N_1492,N_1325,N_1335);
nand U1493 (N_1493,N_1319,N_1395);
nor U1494 (N_1494,N_1308,N_1347);
nor U1495 (N_1495,N_1388,N_1329);
nand U1496 (N_1496,N_1320,N_1376);
and U1497 (N_1497,N_1368,N_1397);
nand U1498 (N_1498,N_1360,N_1312);
or U1499 (N_1499,N_1366,N_1381);
or U1500 (N_1500,N_1477,N_1445);
nand U1501 (N_1501,N_1415,N_1466);
nand U1502 (N_1502,N_1493,N_1414);
and U1503 (N_1503,N_1448,N_1494);
nor U1504 (N_1504,N_1438,N_1463);
or U1505 (N_1505,N_1490,N_1418);
or U1506 (N_1506,N_1421,N_1482);
or U1507 (N_1507,N_1433,N_1412);
xnor U1508 (N_1508,N_1444,N_1458);
and U1509 (N_1509,N_1439,N_1400);
and U1510 (N_1510,N_1429,N_1434);
nand U1511 (N_1511,N_1405,N_1496);
and U1512 (N_1512,N_1422,N_1441);
and U1513 (N_1513,N_1471,N_1436);
or U1514 (N_1514,N_1487,N_1459);
and U1515 (N_1515,N_1498,N_1440);
nand U1516 (N_1516,N_1451,N_1413);
and U1517 (N_1517,N_1492,N_1416);
nand U1518 (N_1518,N_1480,N_1454);
nor U1519 (N_1519,N_1473,N_1428);
nor U1520 (N_1520,N_1425,N_1423);
and U1521 (N_1521,N_1467,N_1462);
and U1522 (N_1522,N_1474,N_1435);
or U1523 (N_1523,N_1402,N_1455);
nor U1524 (N_1524,N_1443,N_1408);
nand U1525 (N_1525,N_1486,N_1452);
nand U1526 (N_1526,N_1460,N_1407);
nand U1527 (N_1527,N_1457,N_1420);
nand U1528 (N_1528,N_1417,N_1485);
or U1529 (N_1529,N_1419,N_1489);
nand U1530 (N_1530,N_1450,N_1499);
and U1531 (N_1531,N_1424,N_1446);
nand U1532 (N_1532,N_1464,N_1437);
nand U1533 (N_1533,N_1449,N_1409);
nand U1534 (N_1534,N_1461,N_1497);
nor U1535 (N_1535,N_1456,N_1431);
and U1536 (N_1536,N_1427,N_1442);
nand U1537 (N_1537,N_1488,N_1470);
nand U1538 (N_1538,N_1469,N_1411);
and U1539 (N_1539,N_1472,N_1430);
or U1540 (N_1540,N_1426,N_1410);
and U1541 (N_1541,N_1495,N_1406);
nor U1542 (N_1542,N_1481,N_1447);
or U1543 (N_1543,N_1483,N_1453);
nor U1544 (N_1544,N_1479,N_1404);
nor U1545 (N_1545,N_1475,N_1484);
or U1546 (N_1546,N_1468,N_1401);
or U1547 (N_1547,N_1478,N_1403);
xor U1548 (N_1548,N_1465,N_1491);
and U1549 (N_1549,N_1432,N_1476);
nor U1550 (N_1550,N_1462,N_1465);
nor U1551 (N_1551,N_1452,N_1461);
nor U1552 (N_1552,N_1404,N_1466);
and U1553 (N_1553,N_1437,N_1405);
or U1554 (N_1554,N_1492,N_1455);
or U1555 (N_1555,N_1470,N_1466);
or U1556 (N_1556,N_1439,N_1409);
nand U1557 (N_1557,N_1430,N_1456);
and U1558 (N_1558,N_1479,N_1423);
or U1559 (N_1559,N_1446,N_1449);
xor U1560 (N_1560,N_1455,N_1431);
nor U1561 (N_1561,N_1494,N_1466);
nand U1562 (N_1562,N_1427,N_1469);
or U1563 (N_1563,N_1408,N_1462);
and U1564 (N_1564,N_1428,N_1414);
nand U1565 (N_1565,N_1443,N_1413);
and U1566 (N_1566,N_1484,N_1443);
nor U1567 (N_1567,N_1403,N_1422);
nand U1568 (N_1568,N_1419,N_1440);
nor U1569 (N_1569,N_1476,N_1428);
and U1570 (N_1570,N_1455,N_1437);
or U1571 (N_1571,N_1474,N_1406);
or U1572 (N_1572,N_1457,N_1476);
or U1573 (N_1573,N_1458,N_1431);
nor U1574 (N_1574,N_1475,N_1449);
or U1575 (N_1575,N_1446,N_1494);
and U1576 (N_1576,N_1406,N_1421);
and U1577 (N_1577,N_1462,N_1497);
nand U1578 (N_1578,N_1489,N_1454);
nor U1579 (N_1579,N_1422,N_1404);
or U1580 (N_1580,N_1440,N_1487);
nor U1581 (N_1581,N_1402,N_1460);
nand U1582 (N_1582,N_1447,N_1422);
or U1583 (N_1583,N_1493,N_1451);
or U1584 (N_1584,N_1492,N_1428);
and U1585 (N_1585,N_1450,N_1448);
or U1586 (N_1586,N_1434,N_1457);
nor U1587 (N_1587,N_1428,N_1432);
xor U1588 (N_1588,N_1480,N_1490);
nand U1589 (N_1589,N_1413,N_1432);
nor U1590 (N_1590,N_1450,N_1461);
or U1591 (N_1591,N_1470,N_1439);
nor U1592 (N_1592,N_1454,N_1446);
or U1593 (N_1593,N_1451,N_1439);
nand U1594 (N_1594,N_1483,N_1458);
and U1595 (N_1595,N_1450,N_1409);
nand U1596 (N_1596,N_1443,N_1462);
nand U1597 (N_1597,N_1486,N_1442);
nand U1598 (N_1598,N_1412,N_1470);
and U1599 (N_1599,N_1434,N_1488);
nor U1600 (N_1600,N_1592,N_1537);
and U1601 (N_1601,N_1527,N_1528);
or U1602 (N_1602,N_1591,N_1510);
nor U1603 (N_1603,N_1547,N_1512);
nand U1604 (N_1604,N_1541,N_1586);
and U1605 (N_1605,N_1575,N_1535);
nand U1606 (N_1606,N_1577,N_1599);
nor U1607 (N_1607,N_1584,N_1587);
nand U1608 (N_1608,N_1589,N_1544);
or U1609 (N_1609,N_1580,N_1560);
and U1610 (N_1610,N_1519,N_1506);
nand U1611 (N_1611,N_1596,N_1517);
nor U1612 (N_1612,N_1593,N_1546);
nor U1613 (N_1613,N_1511,N_1568);
nand U1614 (N_1614,N_1501,N_1516);
and U1615 (N_1615,N_1563,N_1574);
xor U1616 (N_1616,N_1529,N_1551);
nor U1617 (N_1617,N_1559,N_1538);
nor U1618 (N_1618,N_1571,N_1554);
and U1619 (N_1619,N_1515,N_1508);
and U1620 (N_1620,N_1582,N_1509);
nor U1621 (N_1621,N_1556,N_1564);
or U1622 (N_1622,N_1533,N_1558);
or U1623 (N_1623,N_1518,N_1543);
or U1624 (N_1624,N_1525,N_1505);
or U1625 (N_1625,N_1531,N_1520);
nor U1626 (N_1626,N_1576,N_1548);
or U1627 (N_1627,N_1570,N_1545);
nor U1628 (N_1628,N_1539,N_1550);
and U1629 (N_1629,N_1590,N_1567);
nand U1630 (N_1630,N_1566,N_1552);
nor U1631 (N_1631,N_1536,N_1503);
nor U1632 (N_1632,N_1598,N_1504);
nand U1633 (N_1633,N_1581,N_1557);
or U1634 (N_1634,N_1513,N_1555);
nor U1635 (N_1635,N_1578,N_1524);
nand U1636 (N_1636,N_1595,N_1585);
nand U1637 (N_1637,N_1540,N_1561);
and U1638 (N_1638,N_1521,N_1562);
or U1639 (N_1639,N_1502,N_1583);
nand U1640 (N_1640,N_1500,N_1526);
or U1641 (N_1641,N_1565,N_1569);
and U1642 (N_1642,N_1514,N_1542);
nor U1643 (N_1643,N_1573,N_1522);
xnor U1644 (N_1644,N_1572,N_1532);
xnor U1645 (N_1645,N_1530,N_1507);
and U1646 (N_1646,N_1534,N_1588);
and U1647 (N_1647,N_1579,N_1553);
nor U1648 (N_1648,N_1597,N_1594);
nand U1649 (N_1649,N_1549,N_1523);
or U1650 (N_1650,N_1582,N_1593);
nand U1651 (N_1651,N_1588,N_1531);
and U1652 (N_1652,N_1517,N_1502);
and U1653 (N_1653,N_1555,N_1523);
and U1654 (N_1654,N_1571,N_1529);
and U1655 (N_1655,N_1504,N_1529);
nand U1656 (N_1656,N_1523,N_1593);
nor U1657 (N_1657,N_1576,N_1532);
and U1658 (N_1658,N_1599,N_1516);
nor U1659 (N_1659,N_1583,N_1550);
or U1660 (N_1660,N_1557,N_1531);
and U1661 (N_1661,N_1559,N_1543);
and U1662 (N_1662,N_1537,N_1514);
nand U1663 (N_1663,N_1584,N_1525);
nand U1664 (N_1664,N_1558,N_1591);
and U1665 (N_1665,N_1523,N_1553);
or U1666 (N_1666,N_1565,N_1509);
xor U1667 (N_1667,N_1548,N_1583);
nand U1668 (N_1668,N_1501,N_1574);
xnor U1669 (N_1669,N_1560,N_1562);
and U1670 (N_1670,N_1548,N_1553);
or U1671 (N_1671,N_1541,N_1571);
nand U1672 (N_1672,N_1529,N_1575);
and U1673 (N_1673,N_1529,N_1599);
nor U1674 (N_1674,N_1552,N_1577);
nor U1675 (N_1675,N_1560,N_1506);
nor U1676 (N_1676,N_1509,N_1528);
and U1677 (N_1677,N_1563,N_1576);
nor U1678 (N_1678,N_1585,N_1569);
and U1679 (N_1679,N_1552,N_1578);
and U1680 (N_1680,N_1504,N_1531);
and U1681 (N_1681,N_1540,N_1554);
and U1682 (N_1682,N_1548,N_1599);
and U1683 (N_1683,N_1581,N_1596);
nor U1684 (N_1684,N_1562,N_1597);
nand U1685 (N_1685,N_1591,N_1549);
or U1686 (N_1686,N_1525,N_1510);
and U1687 (N_1687,N_1589,N_1563);
nand U1688 (N_1688,N_1589,N_1516);
nor U1689 (N_1689,N_1595,N_1579);
nor U1690 (N_1690,N_1578,N_1527);
nor U1691 (N_1691,N_1562,N_1538);
and U1692 (N_1692,N_1590,N_1570);
or U1693 (N_1693,N_1539,N_1536);
or U1694 (N_1694,N_1592,N_1594);
nand U1695 (N_1695,N_1584,N_1512);
nor U1696 (N_1696,N_1506,N_1554);
nand U1697 (N_1697,N_1563,N_1520);
nor U1698 (N_1698,N_1588,N_1579);
nand U1699 (N_1699,N_1578,N_1553);
and U1700 (N_1700,N_1683,N_1615);
or U1701 (N_1701,N_1643,N_1630);
nor U1702 (N_1702,N_1682,N_1612);
nor U1703 (N_1703,N_1696,N_1658);
nor U1704 (N_1704,N_1623,N_1653);
and U1705 (N_1705,N_1621,N_1674);
or U1706 (N_1706,N_1636,N_1688);
nand U1707 (N_1707,N_1619,N_1691);
or U1708 (N_1708,N_1634,N_1660);
nand U1709 (N_1709,N_1605,N_1600);
or U1710 (N_1710,N_1699,N_1606);
nand U1711 (N_1711,N_1628,N_1626);
and U1712 (N_1712,N_1690,N_1687);
and U1713 (N_1713,N_1659,N_1620);
and U1714 (N_1714,N_1645,N_1616);
nand U1715 (N_1715,N_1602,N_1613);
and U1716 (N_1716,N_1625,N_1631);
and U1717 (N_1717,N_1654,N_1675);
and U1718 (N_1718,N_1676,N_1681);
and U1719 (N_1719,N_1665,N_1641);
nor U1720 (N_1720,N_1697,N_1684);
and U1721 (N_1721,N_1646,N_1642);
and U1722 (N_1722,N_1607,N_1648);
and U1723 (N_1723,N_1652,N_1655);
nor U1724 (N_1724,N_1637,N_1695);
or U1725 (N_1725,N_1694,N_1664);
nand U1726 (N_1726,N_1671,N_1698);
or U1727 (N_1727,N_1651,N_1666);
nor U1728 (N_1728,N_1647,N_1629);
nor U1729 (N_1729,N_1692,N_1689);
or U1730 (N_1730,N_1618,N_1686);
or U1731 (N_1731,N_1601,N_1668);
nand U1732 (N_1732,N_1650,N_1608);
and U1733 (N_1733,N_1640,N_1662);
or U1734 (N_1734,N_1624,N_1611);
nand U1735 (N_1735,N_1669,N_1617);
nand U1736 (N_1736,N_1663,N_1649);
nor U1737 (N_1737,N_1685,N_1673);
nand U1738 (N_1738,N_1678,N_1677);
nor U1739 (N_1739,N_1670,N_1638);
nand U1740 (N_1740,N_1610,N_1604);
or U1741 (N_1741,N_1657,N_1609);
or U1742 (N_1742,N_1644,N_1656);
or U1743 (N_1743,N_1661,N_1680);
nor U1744 (N_1744,N_1639,N_1635);
nand U1745 (N_1745,N_1627,N_1693);
or U1746 (N_1746,N_1633,N_1667);
or U1747 (N_1747,N_1603,N_1632);
or U1748 (N_1748,N_1614,N_1679);
or U1749 (N_1749,N_1622,N_1672);
nor U1750 (N_1750,N_1606,N_1678);
nor U1751 (N_1751,N_1605,N_1606);
and U1752 (N_1752,N_1651,N_1695);
nand U1753 (N_1753,N_1673,N_1650);
nor U1754 (N_1754,N_1647,N_1675);
nor U1755 (N_1755,N_1619,N_1666);
nand U1756 (N_1756,N_1647,N_1636);
or U1757 (N_1757,N_1605,N_1656);
nor U1758 (N_1758,N_1618,N_1699);
or U1759 (N_1759,N_1655,N_1651);
and U1760 (N_1760,N_1640,N_1647);
nand U1761 (N_1761,N_1617,N_1674);
nor U1762 (N_1762,N_1603,N_1694);
nor U1763 (N_1763,N_1661,N_1602);
or U1764 (N_1764,N_1668,N_1617);
or U1765 (N_1765,N_1671,N_1695);
and U1766 (N_1766,N_1655,N_1673);
nand U1767 (N_1767,N_1662,N_1698);
nor U1768 (N_1768,N_1644,N_1684);
xnor U1769 (N_1769,N_1675,N_1678);
nor U1770 (N_1770,N_1642,N_1677);
nand U1771 (N_1771,N_1626,N_1635);
or U1772 (N_1772,N_1624,N_1617);
nand U1773 (N_1773,N_1699,N_1695);
nand U1774 (N_1774,N_1647,N_1643);
nand U1775 (N_1775,N_1695,N_1638);
and U1776 (N_1776,N_1605,N_1696);
nand U1777 (N_1777,N_1687,N_1665);
nor U1778 (N_1778,N_1644,N_1661);
xnor U1779 (N_1779,N_1619,N_1603);
and U1780 (N_1780,N_1698,N_1634);
and U1781 (N_1781,N_1651,N_1616);
nand U1782 (N_1782,N_1694,N_1660);
or U1783 (N_1783,N_1653,N_1697);
nor U1784 (N_1784,N_1692,N_1650);
and U1785 (N_1785,N_1676,N_1631);
or U1786 (N_1786,N_1611,N_1691);
and U1787 (N_1787,N_1630,N_1659);
nor U1788 (N_1788,N_1698,N_1692);
or U1789 (N_1789,N_1666,N_1691);
xnor U1790 (N_1790,N_1628,N_1685);
nor U1791 (N_1791,N_1666,N_1634);
or U1792 (N_1792,N_1668,N_1655);
and U1793 (N_1793,N_1685,N_1607);
nand U1794 (N_1794,N_1698,N_1601);
and U1795 (N_1795,N_1611,N_1625);
nor U1796 (N_1796,N_1617,N_1675);
nand U1797 (N_1797,N_1623,N_1680);
nand U1798 (N_1798,N_1651,N_1632);
nand U1799 (N_1799,N_1608,N_1602);
and U1800 (N_1800,N_1720,N_1767);
or U1801 (N_1801,N_1773,N_1779);
or U1802 (N_1802,N_1701,N_1703);
nor U1803 (N_1803,N_1757,N_1786);
or U1804 (N_1804,N_1775,N_1710);
and U1805 (N_1805,N_1755,N_1741);
nand U1806 (N_1806,N_1748,N_1729);
or U1807 (N_1807,N_1764,N_1787);
and U1808 (N_1808,N_1736,N_1771);
nand U1809 (N_1809,N_1705,N_1790);
or U1810 (N_1810,N_1716,N_1739);
nand U1811 (N_1811,N_1785,N_1776);
or U1812 (N_1812,N_1706,N_1782);
and U1813 (N_1813,N_1784,N_1735);
or U1814 (N_1814,N_1788,N_1722);
nor U1815 (N_1815,N_1744,N_1732);
nor U1816 (N_1816,N_1737,N_1734);
and U1817 (N_1817,N_1752,N_1763);
and U1818 (N_1818,N_1747,N_1733);
or U1819 (N_1819,N_1774,N_1731);
nand U1820 (N_1820,N_1768,N_1772);
xor U1821 (N_1821,N_1702,N_1726);
nor U1822 (N_1822,N_1797,N_1709);
nand U1823 (N_1823,N_1758,N_1789);
and U1824 (N_1824,N_1714,N_1794);
nand U1825 (N_1825,N_1791,N_1730);
nand U1826 (N_1826,N_1700,N_1761);
and U1827 (N_1827,N_1708,N_1718);
or U1828 (N_1828,N_1712,N_1745);
nand U1829 (N_1829,N_1725,N_1760);
nor U1830 (N_1830,N_1721,N_1738);
and U1831 (N_1831,N_1769,N_1749);
or U1832 (N_1832,N_1799,N_1753);
nand U1833 (N_1833,N_1783,N_1740);
nand U1834 (N_1834,N_1750,N_1746);
and U1835 (N_1835,N_1762,N_1728);
or U1836 (N_1836,N_1770,N_1704);
or U1837 (N_1837,N_1798,N_1711);
or U1838 (N_1838,N_1795,N_1759);
or U1839 (N_1839,N_1715,N_1754);
nor U1840 (N_1840,N_1756,N_1777);
nand U1841 (N_1841,N_1766,N_1719);
or U1842 (N_1842,N_1743,N_1723);
nand U1843 (N_1843,N_1751,N_1727);
or U1844 (N_1844,N_1792,N_1781);
and U1845 (N_1845,N_1724,N_1793);
and U1846 (N_1846,N_1713,N_1765);
and U1847 (N_1847,N_1778,N_1707);
or U1848 (N_1848,N_1717,N_1796);
and U1849 (N_1849,N_1742,N_1780);
or U1850 (N_1850,N_1789,N_1798);
or U1851 (N_1851,N_1744,N_1723);
or U1852 (N_1852,N_1769,N_1794);
nor U1853 (N_1853,N_1799,N_1787);
xnor U1854 (N_1854,N_1745,N_1738);
or U1855 (N_1855,N_1713,N_1718);
nand U1856 (N_1856,N_1749,N_1799);
or U1857 (N_1857,N_1793,N_1761);
or U1858 (N_1858,N_1752,N_1736);
nor U1859 (N_1859,N_1797,N_1767);
and U1860 (N_1860,N_1712,N_1759);
and U1861 (N_1861,N_1704,N_1784);
nor U1862 (N_1862,N_1722,N_1736);
or U1863 (N_1863,N_1781,N_1797);
nor U1864 (N_1864,N_1781,N_1724);
and U1865 (N_1865,N_1772,N_1748);
nand U1866 (N_1866,N_1790,N_1731);
or U1867 (N_1867,N_1728,N_1715);
and U1868 (N_1868,N_1789,N_1756);
or U1869 (N_1869,N_1727,N_1768);
nand U1870 (N_1870,N_1778,N_1738);
nand U1871 (N_1871,N_1714,N_1730);
nor U1872 (N_1872,N_1742,N_1770);
xor U1873 (N_1873,N_1719,N_1758);
or U1874 (N_1874,N_1770,N_1739);
or U1875 (N_1875,N_1790,N_1709);
nor U1876 (N_1876,N_1715,N_1766);
and U1877 (N_1877,N_1713,N_1775);
or U1878 (N_1878,N_1771,N_1733);
and U1879 (N_1879,N_1775,N_1701);
or U1880 (N_1880,N_1771,N_1727);
and U1881 (N_1881,N_1767,N_1757);
and U1882 (N_1882,N_1785,N_1737);
and U1883 (N_1883,N_1768,N_1788);
or U1884 (N_1884,N_1705,N_1799);
or U1885 (N_1885,N_1752,N_1704);
nor U1886 (N_1886,N_1751,N_1731);
nor U1887 (N_1887,N_1798,N_1780);
nor U1888 (N_1888,N_1773,N_1796);
nand U1889 (N_1889,N_1743,N_1799);
nand U1890 (N_1890,N_1723,N_1772);
and U1891 (N_1891,N_1773,N_1735);
nor U1892 (N_1892,N_1737,N_1763);
xor U1893 (N_1893,N_1779,N_1768);
and U1894 (N_1894,N_1764,N_1735);
nand U1895 (N_1895,N_1721,N_1724);
or U1896 (N_1896,N_1784,N_1766);
nand U1897 (N_1897,N_1762,N_1790);
nand U1898 (N_1898,N_1763,N_1740);
and U1899 (N_1899,N_1784,N_1741);
xor U1900 (N_1900,N_1819,N_1842);
and U1901 (N_1901,N_1876,N_1893);
or U1902 (N_1902,N_1869,N_1851);
and U1903 (N_1903,N_1839,N_1896);
and U1904 (N_1904,N_1879,N_1880);
nor U1905 (N_1905,N_1837,N_1800);
or U1906 (N_1906,N_1832,N_1888);
and U1907 (N_1907,N_1867,N_1886);
nor U1908 (N_1908,N_1897,N_1887);
and U1909 (N_1909,N_1890,N_1866);
nand U1910 (N_1910,N_1822,N_1877);
or U1911 (N_1911,N_1874,N_1854);
nor U1912 (N_1912,N_1848,N_1827);
and U1913 (N_1913,N_1857,N_1838);
nand U1914 (N_1914,N_1809,N_1878);
nor U1915 (N_1915,N_1823,N_1808);
nor U1916 (N_1916,N_1813,N_1847);
nand U1917 (N_1917,N_1850,N_1840);
nor U1918 (N_1918,N_1891,N_1883);
xnor U1919 (N_1919,N_1895,N_1859);
nor U1920 (N_1920,N_1814,N_1844);
nand U1921 (N_1921,N_1870,N_1889);
and U1922 (N_1922,N_1861,N_1820);
or U1923 (N_1923,N_1871,N_1864);
and U1924 (N_1924,N_1810,N_1855);
or U1925 (N_1925,N_1860,N_1853);
nand U1926 (N_1926,N_1815,N_1824);
nand U1927 (N_1927,N_1845,N_1807);
or U1928 (N_1928,N_1821,N_1868);
nor U1929 (N_1929,N_1801,N_1884);
nor U1930 (N_1930,N_1831,N_1862);
and U1931 (N_1931,N_1852,N_1863);
or U1932 (N_1932,N_1881,N_1829);
xnor U1933 (N_1933,N_1825,N_1894);
and U1934 (N_1934,N_1856,N_1872);
or U1935 (N_1935,N_1841,N_1806);
nor U1936 (N_1936,N_1873,N_1882);
or U1937 (N_1937,N_1803,N_1843);
and U1938 (N_1938,N_1833,N_1817);
or U1939 (N_1939,N_1836,N_1805);
nor U1940 (N_1940,N_1899,N_1818);
nor U1941 (N_1941,N_1885,N_1816);
or U1942 (N_1942,N_1858,N_1865);
and U1943 (N_1943,N_1828,N_1875);
and U1944 (N_1944,N_1812,N_1835);
or U1945 (N_1945,N_1898,N_1849);
and U1946 (N_1946,N_1826,N_1804);
and U1947 (N_1947,N_1846,N_1834);
or U1948 (N_1948,N_1830,N_1811);
nand U1949 (N_1949,N_1802,N_1892);
nand U1950 (N_1950,N_1886,N_1846);
or U1951 (N_1951,N_1810,N_1880);
or U1952 (N_1952,N_1829,N_1879);
or U1953 (N_1953,N_1894,N_1817);
nor U1954 (N_1954,N_1805,N_1887);
nor U1955 (N_1955,N_1853,N_1851);
and U1956 (N_1956,N_1811,N_1874);
nand U1957 (N_1957,N_1838,N_1842);
nor U1958 (N_1958,N_1881,N_1800);
or U1959 (N_1959,N_1808,N_1801);
nand U1960 (N_1960,N_1851,N_1858);
and U1961 (N_1961,N_1896,N_1809);
or U1962 (N_1962,N_1813,N_1870);
nor U1963 (N_1963,N_1857,N_1890);
xor U1964 (N_1964,N_1888,N_1872);
or U1965 (N_1965,N_1879,N_1878);
nor U1966 (N_1966,N_1806,N_1808);
nor U1967 (N_1967,N_1882,N_1835);
nor U1968 (N_1968,N_1843,N_1895);
or U1969 (N_1969,N_1817,N_1849);
or U1970 (N_1970,N_1839,N_1841);
or U1971 (N_1971,N_1891,N_1818);
or U1972 (N_1972,N_1836,N_1884);
and U1973 (N_1973,N_1822,N_1899);
and U1974 (N_1974,N_1860,N_1870);
or U1975 (N_1975,N_1801,N_1810);
or U1976 (N_1976,N_1880,N_1889);
nor U1977 (N_1977,N_1823,N_1853);
and U1978 (N_1978,N_1865,N_1875);
and U1979 (N_1979,N_1821,N_1843);
or U1980 (N_1980,N_1891,N_1857);
and U1981 (N_1981,N_1823,N_1813);
or U1982 (N_1982,N_1841,N_1896);
or U1983 (N_1983,N_1850,N_1812);
and U1984 (N_1984,N_1842,N_1878);
nand U1985 (N_1985,N_1870,N_1835);
nor U1986 (N_1986,N_1880,N_1804);
and U1987 (N_1987,N_1801,N_1874);
or U1988 (N_1988,N_1891,N_1831);
nand U1989 (N_1989,N_1894,N_1800);
nand U1990 (N_1990,N_1855,N_1894);
nor U1991 (N_1991,N_1872,N_1854);
and U1992 (N_1992,N_1825,N_1827);
or U1993 (N_1993,N_1897,N_1868);
and U1994 (N_1994,N_1892,N_1815);
and U1995 (N_1995,N_1848,N_1818);
or U1996 (N_1996,N_1847,N_1872);
nor U1997 (N_1997,N_1839,N_1853);
nor U1998 (N_1998,N_1842,N_1880);
nor U1999 (N_1999,N_1829,N_1883);
and U2000 (N_2000,N_1928,N_1900);
and U2001 (N_2001,N_1911,N_1996);
or U2002 (N_2002,N_1945,N_1978);
and U2003 (N_2003,N_1913,N_1985);
or U2004 (N_2004,N_1990,N_1971);
and U2005 (N_2005,N_1956,N_1926);
nand U2006 (N_2006,N_1950,N_1989);
and U2007 (N_2007,N_1942,N_1962);
and U2008 (N_2008,N_1954,N_1917);
nor U2009 (N_2009,N_1955,N_1959);
nor U2010 (N_2010,N_1952,N_1919);
nor U2011 (N_2011,N_1933,N_1904);
nand U2012 (N_2012,N_1970,N_1997);
nor U2013 (N_2013,N_1908,N_1958);
and U2014 (N_2014,N_1992,N_1976);
xnor U2015 (N_2015,N_1982,N_1924);
nor U2016 (N_2016,N_1964,N_1920);
and U2017 (N_2017,N_1972,N_1902);
nor U2018 (N_2018,N_1969,N_1995);
nand U2019 (N_2019,N_1903,N_1977);
and U2020 (N_2020,N_1941,N_1947);
or U2021 (N_2021,N_1927,N_1966);
nand U2022 (N_2022,N_1931,N_1993);
and U2023 (N_2023,N_1979,N_1988);
or U2024 (N_2024,N_1914,N_1937);
or U2025 (N_2025,N_1986,N_1980);
nand U2026 (N_2026,N_1943,N_1906);
or U2027 (N_2027,N_1929,N_1932);
and U2028 (N_2028,N_1973,N_1949);
and U2029 (N_2029,N_1963,N_1946);
nand U2030 (N_2030,N_1922,N_1925);
nor U2031 (N_2031,N_1916,N_1944);
nor U2032 (N_2032,N_1953,N_1951);
and U2033 (N_2033,N_1901,N_1923);
xor U2034 (N_2034,N_1934,N_1915);
or U2035 (N_2035,N_1968,N_1961);
or U2036 (N_2036,N_1960,N_1936);
nor U2037 (N_2037,N_1921,N_1905);
nor U2038 (N_2038,N_1975,N_1912);
and U2039 (N_2039,N_1974,N_1984);
nor U2040 (N_2040,N_1935,N_1918);
or U2041 (N_2041,N_1991,N_1998);
and U2042 (N_2042,N_1940,N_1965);
and U2043 (N_2043,N_1957,N_1983);
and U2044 (N_2044,N_1938,N_1930);
or U2045 (N_2045,N_1910,N_1907);
and U2046 (N_2046,N_1999,N_1987);
and U2047 (N_2047,N_1981,N_1948);
or U2048 (N_2048,N_1939,N_1909);
nor U2049 (N_2049,N_1967,N_1994);
nand U2050 (N_2050,N_1994,N_1933);
or U2051 (N_2051,N_1979,N_1989);
nand U2052 (N_2052,N_1958,N_1928);
and U2053 (N_2053,N_1985,N_1954);
nand U2054 (N_2054,N_1981,N_1986);
and U2055 (N_2055,N_1909,N_1968);
and U2056 (N_2056,N_1954,N_1946);
or U2057 (N_2057,N_1980,N_1944);
or U2058 (N_2058,N_1912,N_1916);
or U2059 (N_2059,N_1984,N_1995);
or U2060 (N_2060,N_1999,N_1906);
nor U2061 (N_2061,N_1969,N_1928);
nand U2062 (N_2062,N_1911,N_1932);
or U2063 (N_2063,N_1939,N_1958);
nand U2064 (N_2064,N_1964,N_1931);
nand U2065 (N_2065,N_1980,N_1993);
nor U2066 (N_2066,N_1914,N_1917);
nor U2067 (N_2067,N_1920,N_1986);
nand U2068 (N_2068,N_1961,N_1978);
and U2069 (N_2069,N_1909,N_1947);
nand U2070 (N_2070,N_1982,N_1900);
nand U2071 (N_2071,N_1953,N_1926);
nand U2072 (N_2072,N_1901,N_1987);
and U2073 (N_2073,N_1974,N_1981);
or U2074 (N_2074,N_1976,N_1954);
or U2075 (N_2075,N_1941,N_1938);
nor U2076 (N_2076,N_1954,N_1918);
nor U2077 (N_2077,N_1905,N_1954);
nand U2078 (N_2078,N_1987,N_1956);
nor U2079 (N_2079,N_1953,N_1944);
nand U2080 (N_2080,N_1986,N_1944);
or U2081 (N_2081,N_1983,N_1956);
nand U2082 (N_2082,N_1996,N_1934);
xnor U2083 (N_2083,N_1909,N_1903);
nor U2084 (N_2084,N_1964,N_1956);
nand U2085 (N_2085,N_1951,N_1957);
nor U2086 (N_2086,N_1928,N_1996);
or U2087 (N_2087,N_1910,N_1982);
nor U2088 (N_2088,N_1955,N_1905);
or U2089 (N_2089,N_1934,N_1952);
nand U2090 (N_2090,N_1990,N_1981);
and U2091 (N_2091,N_1920,N_1902);
nor U2092 (N_2092,N_1951,N_1995);
and U2093 (N_2093,N_1914,N_1980);
nand U2094 (N_2094,N_1919,N_1941);
nor U2095 (N_2095,N_1974,N_1978);
and U2096 (N_2096,N_1992,N_1967);
and U2097 (N_2097,N_1971,N_1992);
xor U2098 (N_2098,N_1924,N_1933);
or U2099 (N_2099,N_1932,N_1931);
or U2100 (N_2100,N_2061,N_2028);
or U2101 (N_2101,N_2076,N_2096);
or U2102 (N_2102,N_2060,N_2014);
and U2103 (N_2103,N_2021,N_2052);
nor U2104 (N_2104,N_2062,N_2099);
or U2105 (N_2105,N_2011,N_2094);
and U2106 (N_2106,N_2022,N_2008);
or U2107 (N_2107,N_2066,N_2064);
or U2108 (N_2108,N_2049,N_2092);
and U2109 (N_2109,N_2025,N_2009);
or U2110 (N_2110,N_2074,N_2081);
and U2111 (N_2111,N_2029,N_2097);
xor U2112 (N_2112,N_2006,N_2077);
nand U2113 (N_2113,N_2016,N_2095);
and U2114 (N_2114,N_2053,N_2044);
or U2115 (N_2115,N_2072,N_2089);
or U2116 (N_2116,N_2069,N_2055);
or U2117 (N_2117,N_2015,N_2056);
xor U2118 (N_2118,N_2043,N_2087);
nand U2119 (N_2119,N_2051,N_2079);
and U2120 (N_2120,N_2039,N_2032);
or U2121 (N_2121,N_2057,N_2042);
or U2122 (N_2122,N_2068,N_2027);
xnor U2123 (N_2123,N_2054,N_2088);
nand U2124 (N_2124,N_2019,N_2048);
nor U2125 (N_2125,N_2059,N_2020);
nor U2126 (N_2126,N_2084,N_2073);
nand U2127 (N_2127,N_2046,N_2047);
nand U2128 (N_2128,N_2031,N_2010);
or U2129 (N_2129,N_2004,N_2041);
nand U2130 (N_2130,N_2065,N_2078);
and U2131 (N_2131,N_2036,N_2075);
nor U2132 (N_2132,N_2086,N_2082);
nand U2133 (N_2133,N_2090,N_2063);
nand U2134 (N_2134,N_2080,N_2093);
nand U2135 (N_2135,N_2005,N_2000);
xnor U2136 (N_2136,N_2071,N_2007);
or U2137 (N_2137,N_2034,N_2030);
nor U2138 (N_2138,N_2026,N_2003);
and U2139 (N_2139,N_2033,N_2024);
and U2140 (N_2140,N_2001,N_2040);
and U2141 (N_2141,N_2045,N_2067);
or U2142 (N_2142,N_2002,N_2013);
or U2143 (N_2143,N_2085,N_2091);
or U2144 (N_2144,N_2037,N_2012);
or U2145 (N_2145,N_2017,N_2038);
nor U2146 (N_2146,N_2018,N_2058);
and U2147 (N_2147,N_2083,N_2070);
and U2148 (N_2148,N_2023,N_2050);
nor U2149 (N_2149,N_2035,N_2098);
or U2150 (N_2150,N_2097,N_2086);
and U2151 (N_2151,N_2074,N_2076);
nand U2152 (N_2152,N_2003,N_2043);
and U2153 (N_2153,N_2024,N_2070);
or U2154 (N_2154,N_2072,N_2006);
and U2155 (N_2155,N_2029,N_2082);
nor U2156 (N_2156,N_2080,N_2028);
nor U2157 (N_2157,N_2062,N_2025);
nand U2158 (N_2158,N_2098,N_2057);
or U2159 (N_2159,N_2099,N_2090);
nand U2160 (N_2160,N_2083,N_2066);
and U2161 (N_2161,N_2082,N_2012);
nand U2162 (N_2162,N_2095,N_2043);
nor U2163 (N_2163,N_2093,N_2064);
and U2164 (N_2164,N_2010,N_2059);
and U2165 (N_2165,N_2024,N_2013);
nor U2166 (N_2166,N_2045,N_2047);
and U2167 (N_2167,N_2074,N_2015);
nor U2168 (N_2168,N_2004,N_2095);
nor U2169 (N_2169,N_2038,N_2027);
nand U2170 (N_2170,N_2095,N_2076);
nand U2171 (N_2171,N_2054,N_2070);
and U2172 (N_2172,N_2044,N_2096);
nor U2173 (N_2173,N_2086,N_2030);
and U2174 (N_2174,N_2081,N_2089);
nor U2175 (N_2175,N_2018,N_2044);
and U2176 (N_2176,N_2058,N_2052);
or U2177 (N_2177,N_2047,N_2004);
or U2178 (N_2178,N_2075,N_2016);
or U2179 (N_2179,N_2049,N_2085);
nor U2180 (N_2180,N_2061,N_2074);
nand U2181 (N_2181,N_2028,N_2032);
and U2182 (N_2182,N_2010,N_2004);
nand U2183 (N_2183,N_2015,N_2065);
or U2184 (N_2184,N_2033,N_2028);
and U2185 (N_2185,N_2028,N_2078);
and U2186 (N_2186,N_2033,N_2027);
and U2187 (N_2187,N_2086,N_2015);
and U2188 (N_2188,N_2081,N_2067);
nand U2189 (N_2189,N_2091,N_2019);
nand U2190 (N_2190,N_2080,N_2010);
nor U2191 (N_2191,N_2024,N_2023);
nand U2192 (N_2192,N_2044,N_2027);
and U2193 (N_2193,N_2096,N_2084);
nor U2194 (N_2194,N_2004,N_2070);
and U2195 (N_2195,N_2089,N_2088);
and U2196 (N_2196,N_2097,N_2096);
nor U2197 (N_2197,N_2084,N_2037);
or U2198 (N_2198,N_2068,N_2061);
and U2199 (N_2199,N_2036,N_2003);
and U2200 (N_2200,N_2140,N_2142);
and U2201 (N_2201,N_2176,N_2190);
nand U2202 (N_2202,N_2164,N_2192);
nand U2203 (N_2203,N_2122,N_2110);
nand U2204 (N_2204,N_2172,N_2106);
nor U2205 (N_2205,N_2146,N_2163);
nand U2206 (N_2206,N_2195,N_2141);
nor U2207 (N_2207,N_2139,N_2159);
or U2208 (N_2208,N_2152,N_2132);
and U2209 (N_2209,N_2133,N_2111);
and U2210 (N_2210,N_2119,N_2130);
nor U2211 (N_2211,N_2124,N_2136);
nand U2212 (N_2212,N_2162,N_2128);
or U2213 (N_2213,N_2125,N_2134);
nand U2214 (N_2214,N_2104,N_2103);
and U2215 (N_2215,N_2184,N_2149);
nor U2216 (N_2216,N_2171,N_2182);
nor U2217 (N_2217,N_2198,N_2179);
nand U2218 (N_2218,N_2188,N_2154);
nand U2219 (N_2219,N_2145,N_2153);
nor U2220 (N_2220,N_2177,N_2151);
nor U2221 (N_2221,N_2118,N_2155);
nand U2222 (N_2222,N_2158,N_2197);
or U2223 (N_2223,N_2187,N_2169);
and U2224 (N_2224,N_2117,N_2112);
nor U2225 (N_2225,N_2160,N_2113);
and U2226 (N_2226,N_2108,N_2109);
nor U2227 (N_2227,N_2199,N_2191);
xnor U2228 (N_2228,N_2193,N_2114);
or U2229 (N_2229,N_2185,N_2143);
or U2230 (N_2230,N_2183,N_2175);
and U2231 (N_2231,N_2156,N_2148);
and U2232 (N_2232,N_2157,N_2166);
or U2233 (N_2233,N_2131,N_2144);
or U2234 (N_2234,N_2174,N_2127);
nor U2235 (N_2235,N_2181,N_2121);
and U2236 (N_2236,N_2138,N_2107);
and U2237 (N_2237,N_2100,N_2168);
and U2238 (N_2238,N_2147,N_2194);
or U2239 (N_2239,N_2120,N_2161);
and U2240 (N_2240,N_2170,N_2126);
nand U2241 (N_2241,N_2180,N_2167);
nand U2242 (N_2242,N_2137,N_2105);
and U2243 (N_2243,N_2189,N_2165);
nand U2244 (N_2244,N_2178,N_2101);
nand U2245 (N_2245,N_2135,N_2123);
or U2246 (N_2246,N_2115,N_2186);
nand U2247 (N_2247,N_2102,N_2129);
nor U2248 (N_2248,N_2196,N_2150);
and U2249 (N_2249,N_2173,N_2116);
and U2250 (N_2250,N_2120,N_2133);
and U2251 (N_2251,N_2197,N_2131);
nor U2252 (N_2252,N_2137,N_2175);
nand U2253 (N_2253,N_2195,N_2116);
and U2254 (N_2254,N_2171,N_2162);
or U2255 (N_2255,N_2142,N_2125);
or U2256 (N_2256,N_2194,N_2154);
nand U2257 (N_2257,N_2111,N_2199);
or U2258 (N_2258,N_2159,N_2114);
or U2259 (N_2259,N_2182,N_2104);
nor U2260 (N_2260,N_2152,N_2136);
or U2261 (N_2261,N_2160,N_2166);
nor U2262 (N_2262,N_2106,N_2188);
nor U2263 (N_2263,N_2143,N_2190);
and U2264 (N_2264,N_2147,N_2107);
or U2265 (N_2265,N_2146,N_2112);
nor U2266 (N_2266,N_2123,N_2197);
nand U2267 (N_2267,N_2169,N_2179);
and U2268 (N_2268,N_2130,N_2169);
nand U2269 (N_2269,N_2187,N_2101);
nand U2270 (N_2270,N_2136,N_2170);
and U2271 (N_2271,N_2187,N_2183);
and U2272 (N_2272,N_2196,N_2103);
or U2273 (N_2273,N_2176,N_2188);
or U2274 (N_2274,N_2136,N_2133);
and U2275 (N_2275,N_2174,N_2185);
or U2276 (N_2276,N_2152,N_2178);
or U2277 (N_2277,N_2138,N_2183);
and U2278 (N_2278,N_2188,N_2151);
and U2279 (N_2279,N_2170,N_2125);
or U2280 (N_2280,N_2129,N_2122);
nor U2281 (N_2281,N_2101,N_2117);
or U2282 (N_2282,N_2115,N_2180);
nand U2283 (N_2283,N_2123,N_2166);
or U2284 (N_2284,N_2105,N_2168);
nand U2285 (N_2285,N_2109,N_2167);
and U2286 (N_2286,N_2155,N_2122);
and U2287 (N_2287,N_2139,N_2186);
or U2288 (N_2288,N_2147,N_2168);
and U2289 (N_2289,N_2182,N_2112);
nor U2290 (N_2290,N_2104,N_2156);
nor U2291 (N_2291,N_2144,N_2185);
nand U2292 (N_2292,N_2103,N_2163);
nor U2293 (N_2293,N_2177,N_2159);
and U2294 (N_2294,N_2127,N_2153);
and U2295 (N_2295,N_2139,N_2185);
nor U2296 (N_2296,N_2127,N_2115);
nor U2297 (N_2297,N_2113,N_2174);
nor U2298 (N_2298,N_2111,N_2184);
xor U2299 (N_2299,N_2112,N_2116);
or U2300 (N_2300,N_2214,N_2220);
nor U2301 (N_2301,N_2218,N_2271);
nand U2302 (N_2302,N_2290,N_2266);
nand U2303 (N_2303,N_2236,N_2222);
or U2304 (N_2304,N_2263,N_2204);
and U2305 (N_2305,N_2212,N_2225);
xnor U2306 (N_2306,N_2232,N_2258);
nor U2307 (N_2307,N_2260,N_2238);
and U2308 (N_2308,N_2257,N_2297);
xnor U2309 (N_2309,N_2209,N_2241);
nor U2310 (N_2310,N_2216,N_2235);
nor U2311 (N_2311,N_2207,N_2256);
and U2312 (N_2312,N_2203,N_2205);
or U2313 (N_2313,N_2245,N_2278);
nand U2314 (N_2314,N_2239,N_2282);
nor U2315 (N_2315,N_2215,N_2228);
or U2316 (N_2316,N_2277,N_2206);
nand U2317 (N_2317,N_2233,N_2243);
and U2318 (N_2318,N_2286,N_2227);
and U2319 (N_2319,N_2237,N_2299);
nand U2320 (N_2320,N_2211,N_2247);
and U2321 (N_2321,N_2281,N_2223);
or U2322 (N_2322,N_2250,N_2242);
nand U2323 (N_2323,N_2251,N_2272);
or U2324 (N_2324,N_2283,N_2259);
and U2325 (N_2325,N_2249,N_2219);
nand U2326 (N_2326,N_2224,N_2202);
or U2327 (N_2327,N_2221,N_2248);
nand U2328 (N_2328,N_2270,N_2289);
nor U2329 (N_2329,N_2213,N_2296);
nor U2330 (N_2330,N_2264,N_2210);
or U2331 (N_2331,N_2269,N_2244);
and U2332 (N_2332,N_2293,N_2273);
nor U2333 (N_2333,N_2246,N_2274);
and U2334 (N_2334,N_2265,N_2261);
nor U2335 (N_2335,N_2268,N_2255);
nand U2336 (N_2336,N_2291,N_2240);
and U2337 (N_2337,N_2231,N_2253);
or U2338 (N_2338,N_2279,N_2280);
nor U2339 (N_2339,N_2234,N_2294);
nor U2340 (N_2340,N_2275,N_2208);
nand U2341 (N_2341,N_2252,N_2226);
nand U2342 (N_2342,N_2292,N_2229);
nor U2343 (N_2343,N_2230,N_2254);
nand U2344 (N_2344,N_2295,N_2285);
nor U2345 (N_2345,N_2267,N_2298);
nor U2346 (N_2346,N_2276,N_2217);
nand U2347 (N_2347,N_2201,N_2288);
nand U2348 (N_2348,N_2200,N_2262);
nand U2349 (N_2349,N_2284,N_2287);
and U2350 (N_2350,N_2223,N_2294);
nand U2351 (N_2351,N_2251,N_2233);
and U2352 (N_2352,N_2219,N_2230);
nor U2353 (N_2353,N_2286,N_2237);
nor U2354 (N_2354,N_2216,N_2243);
or U2355 (N_2355,N_2218,N_2252);
or U2356 (N_2356,N_2263,N_2217);
nor U2357 (N_2357,N_2282,N_2211);
nor U2358 (N_2358,N_2272,N_2224);
or U2359 (N_2359,N_2270,N_2242);
nand U2360 (N_2360,N_2272,N_2298);
and U2361 (N_2361,N_2234,N_2285);
nor U2362 (N_2362,N_2242,N_2241);
nand U2363 (N_2363,N_2276,N_2237);
nor U2364 (N_2364,N_2252,N_2211);
or U2365 (N_2365,N_2213,N_2254);
or U2366 (N_2366,N_2261,N_2241);
or U2367 (N_2367,N_2297,N_2234);
xor U2368 (N_2368,N_2292,N_2283);
and U2369 (N_2369,N_2246,N_2290);
nand U2370 (N_2370,N_2257,N_2225);
nor U2371 (N_2371,N_2291,N_2277);
or U2372 (N_2372,N_2216,N_2232);
nand U2373 (N_2373,N_2207,N_2248);
or U2374 (N_2374,N_2254,N_2229);
nand U2375 (N_2375,N_2228,N_2251);
or U2376 (N_2376,N_2238,N_2259);
or U2377 (N_2377,N_2290,N_2216);
or U2378 (N_2378,N_2237,N_2243);
or U2379 (N_2379,N_2253,N_2260);
or U2380 (N_2380,N_2226,N_2251);
nand U2381 (N_2381,N_2233,N_2288);
and U2382 (N_2382,N_2230,N_2276);
and U2383 (N_2383,N_2270,N_2286);
nand U2384 (N_2384,N_2256,N_2205);
nand U2385 (N_2385,N_2294,N_2201);
nor U2386 (N_2386,N_2241,N_2244);
and U2387 (N_2387,N_2257,N_2216);
nand U2388 (N_2388,N_2297,N_2265);
nor U2389 (N_2389,N_2267,N_2241);
nor U2390 (N_2390,N_2214,N_2256);
and U2391 (N_2391,N_2215,N_2237);
or U2392 (N_2392,N_2252,N_2295);
nor U2393 (N_2393,N_2253,N_2274);
and U2394 (N_2394,N_2208,N_2228);
or U2395 (N_2395,N_2239,N_2229);
or U2396 (N_2396,N_2228,N_2217);
xnor U2397 (N_2397,N_2244,N_2242);
nor U2398 (N_2398,N_2266,N_2291);
and U2399 (N_2399,N_2203,N_2272);
and U2400 (N_2400,N_2388,N_2354);
or U2401 (N_2401,N_2371,N_2303);
nand U2402 (N_2402,N_2360,N_2396);
and U2403 (N_2403,N_2369,N_2373);
and U2404 (N_2404,N_2320,N_2340);
nor U2405 (N_2405,N_2319,N_2337);
or U2406 (N_2406,N_2317,N_2346);
and U2407 (N_2407,N_2358,N_2321);
and U2408 (N_2408,N_2310,N_2306);
or U2409 (N_2409,N_2386,N_2339);
nand U2410 (N_2410,N_2392,N_2382);
nand U2411 (N_2411,N_2355,N_2381);
nand U2412 (N_2412,N_2377,N_2387);
and U2413 (N_2413,N_2335,N_2353);
xnor U2414 (N_2414,N_2397,N_2375);
and U2415 (N_2415,N_2325,N_2326);
or U2416 (N_2416,N_2372,N_2364);
or U2417 (N_2417,N_2332,N_2395);
and U2418 (N_2418,N_2367,N_2370);
nand U2419 (N_2419,N_2398,N_2301);
nand U2420 (N_2420,N_2349,N_2351);
nor U2421 (N_2421,N_2342,N_2368);
nor U2422 (N_2422,N_2341,N_2393);
and U2423 (N_2423,N_2313,N_2347);
and U2424 (N_2424,N_2390,N_2348);
nand U2425 (N_2425,N_2331,N_2330);
nor U2426 (N_2426,N_2352,N_2374);
nor U2427 (N_2427,N_2328,N_2394);
xnor U2428 (N_2428,N_2350,N_2338);
nor U2429 (N_2429,N_2344,N_2309);
or U2430 (N_2430,N_2389,N_2302);
or U2431 (N_2431,N_2356,N_2305);
and U2432 (N_2432,N_2308,N_2300);
nand U2433 (N_2433,N_2345,N_2333);
nand U2434 (N_2434,N_2312,N_2316);
and U2435 (N_2435,N_2311,N_2324);
and U2436 (N_2436,N_2362,N_2399);
nor U2437 (N_2437,N_2379,N_2322);
and U2438 (N_2438,N_2361,N_2376);
or U2439 (N_2439,N_2307,N_2314);
nand U2440 (N_2440,N_2329,N_2318);
and U2441 (N_2441,N_2365,N_2366);
nor U2442 (N_2442,N_2304,N_2327);
and U2443 (N_2443,N_2315,N_2384);
and U2444 (N_2444,N_2336,N_2359);
nand U2445 (N_2445,N_2385,N_2391);
and U2446 (N_2446,N_2343,N_2323);
and U2447 (N_2447,N_2383,N_2363);
or U2448 (N_2448,N_2380,N_2334);
and U2449 (N_2449,N_2378,N_2357);
nor U2450 (N_2450,N_2368,N_2304);
nand U2451 (N_2451,N_2347,N_2395);
or U2452 (N_2452,N_2391,N_2319);
and U2453 (N_2453,N_2385,N_2367);
nand U2454 (N_2454,N_2384,N_2334);
and U2455 (N_2455,N_2363,N_2324);
and U2456 (N_2456,N_2353,N_2333);
nor U2457 (N_2457,N_2353,N_2309);
or U2458 (N_2458,N_2350,N_2363);
nor U2459 (N_2459,N_2331,N_2319);
nor U2460 (N_2460,N_2317,N_2398);
nor U2461 (N_2461,N_2333,N_2313);
and U2462 (N_2462,N_2388,N_2347);
or U2463 (N_2463,N_2378,N_2331);
nor U2464 (N_2464,N_2338,N_2310);
nor U2465 (N_2465,N_2321,N_2325);
nand U2466 (N_2466,N_2302,N_2387);
and U2467 (N_2467,N_2309,N_2325);
or U2468 (N_2468,N_2355,N_2370);
nand U2469 (N_2469,N_2309,N_2331);
nor U2470 (N_2470,N_2378,N_2339);
or U2471 (N_2471,N_2349,N_2383);
nor U2472 (N_2472,N_2374,N_2317);
nor U2473 (N_2473,N_2324,N_2359);
nand U2474 (N_2474,N_2334,N_2394);
nand U2475 (N_2475,N_2390,N_2327);
and U2476 (N_2476,N_2308,N_2321);
or U2477 (N_2477,N_2378,N_2377);
nand U2478 (N_2478,N_2374,N_2353);
and U2479 (N_2479,N_2322,N_2380);
and U2480 (N_2480,N_2314,N_2320);
xnor U2481 (N_2481,N_2396,N_2384);
or U2482 (N_2482,N_2391,N_2317);
nand U2483 (N_2483,N_2325,N_2311);
and U2484 (N_2484,N_2380,N_2376);
nand U2485 (N_2485,N_2333,N_2388);
nor U2486 (N_2486,N_2317,N_2383);
nor U2487 (N_2487,N_2328,N_2318);
nor U2488 (N_2488,N_2390,N_2329);
xnor U2489 (N_2489,N_2391,N_2383);
nand U2490 (N_2490,N_2316,N_2322);
or U2491 (N_2491,N_2375,N_2346);
nand U2492 (N_2492,N_2306,N_2374);
or U2493 (N_2493,N_2313,N_2394);
nor U2494 (N_2494,N_2361,N_2329);
or U2495 (N_2495,N_2308,N_2314);
nand U2496 (N_2496,N_2376,N_2362);
nor U2497 (N_2497,N_2353,N_2396);
xnor U2498 (N_2498,N_2328,N_2346);
and U2499 (N_2499,N_2315,N_2387);
nor U2500 (N_2500,N_2469,N_2438);
nor U2501 (N_2501,N_2409,N_2444);
nor U2502 (N_2502,N_2453,N_2433);
and U2503 (N_2503,N_2454,N_2484);
nand U2504 (N_2504,N_2481,N_2498);
or U2505 (N_2505,N_2414,N_2422);
and U2506 (N_2506,N_2429,N_2448);
and U2507 (N_2507,N_2485,N_2405);
nand U2508 (N_2508,N_2434,N_2497);
or U2509 (N_2509,N_2499,N_2447);
nor U2510 (N_2510,N_2431,N_2491);
or U2511 (N_2511,N_2449,N_2442);
nor U2512 (N_2512,N_2432,N_2459);
and U2513 (N_2513,N_2426,N_2441);
xor U2514 (N_2514,N_2492,N_2402);
nand U2515 (N_2515,N_2452,N_2451);
nand U2516 (N_2516,N_2430,N_2486);
nor U2517 (N_2517,N_2472,N_2471);
or U2518 (N_2518,N_2439,N_2416);
or U2519 (N_2519,N_2421,N_2417);
and U2520 (N_2520,N_2482,N_2455);
and U2521 (N_2521,N_2456,N_2468);
or U2522 (N_2522,N_2477,N_2413);
and U2523 (N_2523,N_2445,N_2403);
or U2524 (N_2524,N_2490,N_2496);
nand U2525 (N_2525,N_2435,N_2464);
or U2526 (N_2526,N_2458,N_2450);
or U2527 (N_2527,N_2408,N_2461);
nor U2528 (N_2528,N_2424,N_2475);
nor U2529 (N_2529,N_2495,N_2443);
nor U2530 (N_2530,N_2420,N_2411);
and U2531 (N_2531,N_2400,N_2476);
nor U2532 (N_2532,N_2479,N_2412);
nor U2533 (N_2533,N_2446,N_2406);
and U2534 (N_2534,N_2460,N_2437);
xor U2535 (N_2535,N_2404,N_2494);
nor U2536 (N_2536,N_2467,N_2407);
or U2537 (N_2537,N_2487,N_2428);
or U2538 (N_2538,N_2462,N_2489);
nand U2539 (N_2539,N_2427,N_2480);
nand U2540 (N_2540,N_2488,N_2493);
or U2541 (N_2541,N_2457,N_2466);
nor U2542 (N_2542,N_2425,N_2474);
or U2543 (N_2543,N_2483,N_2478);
nor U2544 (N_2544,N_2470,N_2423);
nor U2545 (N_2545,N_2440,N_2419);
nand U2546 (N_2546,N_2465,N_2473);
and U2547 (N_2547,N_2401,N_2463);
xnor U2548 (N_2548,N_2436,N_2410);
and U2549 (N_2549,N_2418,N_2415);
or U2550 (N_2550,N_2494,N_2498);
nor U2551 (N_2551,N_2492,N_2456);
nor U2552 (N_2552,N_2403,N_2428);
nor U2553 (N_2553,N_2460,N_2494);
or U2554 (N_2554,N_2405,N_2426);
and U2555 (N_2555,N_2410,N_2434);
and U2556 (N_2556,N_2454,N_2457);
nand U2557 (N_2557,N_2420,N_2413);
nor U2558 (N_2558,N_2448,N_2493);
or U2559 (N_2559,N_2444,N_2416);
or U2560 (N_2560,N_2438,N_2403);
nand U2561 (N_2561,N_2450,N_2414);
nand U2562 (N_2562,N_2499,N_2414);
nand U2563 (N_2563,N_2482,N_2495);
nand U2564 (N_2564,N_2447,N_2485);
and U2565 (N_2565,N_2435,N_2437);
and U2566 (N_2566,N_2468,N_2409);
nor U2567 (N_2567,N_2466,N_2412);
and U2568 (N_2568,N_2410,N_2470);
and U2569 (N_2569,N_2460,N_2401);
nand U2570 (N_2570,N_2428,N_2455);
and U2571 (N_2571,N_2481,N_2499);
nor U2572 (N_2572,N_2424,N_2450);
or U2573 (N_2573,N_2400,N_2412);
nand U2574 (N_2574,N_2468,N_2429);
and U2575 (N_2575,N_2456,N_2460);
xor U2576 (N_2576,N_2480,N_2408);
nor U2577 (N_2577,N_2480,N_2474);
nand U2578 (N_2578,N_2441,N_2416);
and U2579 (N_2579,N_2458,N_2456);
nor U2580 (N_2580,N_2412,N_2423);
nand U2581 (N_2581,N_2477,N_2450);
and U2582 (N_2582,N_2444,N_2432);
nor U2583 (N_2583,N_2487,N_2460);
nor U2584 (N_2584,N_2458,N_2448);
or U2585 (N_2585,N_2450,N_2418);
nand U2586 (N_2586,N_2440,N_2446);
or U2587 (N_2587,N_2455,N_2415);
nor U2588 (N_2588,N_2482,N_2408);
nand U2589 (N_2589,N_2418,N_2452);
nand U2590 (N_2590,N_2481,N_2431);
and U2591 (N_2591,N_2411,N_2452);
and U2592 (N_2592,N_2428,N_2459);
and U2593 (N_2593,N_2436,N_2406);
and U2594 (N_2594,N_2484,N_2402);
nor U2595 (N_2595,N_2431,N_2498);
and U2596 (N_2596,N_2426,N_2438);
or U2597 (N_2597,N_2426,N_2446);
or U2598 (N_2598,N_2421,N_2430);
or U2599 (N_2599,N_2447,N_2493);
and U2600 (N_2600,N_2519,N_2599);
or U2601 (N_2601,N_2579,N_2520);
nand U2602 (N_2602,N_2565,N_2502);
nor U2603 (N_2603,N_2593,N_2518);
nor U2604 (N_2604,N_2546,N_2561);
or U2605 (N_2605,N_2528,N_2549);
and U2606 (N_2606,N_2512,N_2532);
nand U2607 (N_2607,N_2504,N_2550);
and U2608 (N_2608,N_2539,N_2511);
and U2609 (N_2609,N_2573,N_2576);
nand U2610 (N_2610,N_2580,N_2521);
or U2611 (N_2611,N_2513,N_2592);
and U2612 (N_2612,N_2586,N_2584);
nor U2613 (N_2613,N_2536,N_2548);
or U2614 (N_2614,N_2563,N_2529);
nor U2615 (N_2615,N_2556,N_2575);
nor U2616 (N_2616,N_2501,N_2538);
nand U2617 (N_2617,N_2570,N_2597);
nand U2618 (N_2618,N_2517,N_2596);
and U2619 (N_2619,N_2571,N_2567);
or U2620 (N_2620,N_2560,N_2583);
and U2621 (N_2621,N_2587,N_2594);
nor U2622 (N_2622,N_2506,N_2535);
and U2623 (N_2623,N_2537,N_2582);
or U2624 (N_2624,N_2558,N_2507);
or U2625 (N_2625,N_2574,N_2541);
nand U2626 (N_2626,N_2559,N_2569);
nand U2627 (N_2627,N_2505,N_2545);
and U2628 (N_2628,N_2523,N_2522);
and U2629 (N_2629,N_2503,N_2557);
or U2630 (N_2630,N_2595,N_2526);
nor U2631 (N_2631,N_2540,N_2572);
and U2632 (N_2632,N_2534,N_2530);
xor U2633 (N_2633,N_2598,N_2544);
and U2634 (N_2634,N_2525,N_2552);
and U2635 (N_2635,N_2554,N_2510);
or U2636 (N_2636,N_2591,N_2524);
nor U2637 (N_2637,N_2516,N_2547);
nand U2638 (N_2638,N_2585,N_2578);
and U2639 (N_2639,N_2581,N_2542);
nor U2640 (N_2640,N_2533,N_2588);
nor U2641 (N_2641,N_2562,N_2553);
nand U2642 (N_2642,N_2589,N_2551);
or U2643 (N_2643,N_2566,N_2514);
nand U2644 (N_2644,N_2527,N_2577);
or U2645 (N_2645,N_2531,N_2500);
and U2646 (N_2646,N_2590,N_2508);
and U2647 (N_2647,N_2543,N_2515);
or U2648 (N_2648,N_2509,N_2568);
and U2649 (N_2649,N_2564,N_2555);
nor U2650 (N_2650,N_2563,N_2555);
or U2651 (N_2651,N_2564,N_2517);
or U2652 (N_2652,N_2527,N_2522);
and U2653 (N_2653,N_2580,N_2594);
or U2654 (N_2654,N_2502,N_2587);
nand U2655 (N_2655,N_2518,N_2599);
nand U2656 (N_2656,N_2530,N_2522);
and U2657 (N_2657,N_2594,N_2534);
nor U2658 (N_2658,N_2563,N_2589);
nor U2659 (N_2659,N_2504,N_2554);
or U2660 (N_2660,N_2555,N_2584);
nand U2661 (N_2661,N_2565,N_2551);
nor U2662 (N_2662,N_2585,N_2546);
or U2663 (N_2663,N_2594,N_2535);
nand U2664 (N_2664,N_2579,N_2537);
or U2665 (N_2665,N_2551,N_2585);
and U2666 (N_2666,N_2555,N_2590);
or U2667 (N_2667,N_2544,N_2539);
or U2668 (N_2668,N_2520,N_2594);
nand U2669 (N_2669,N_2525,N_2570);
and U2670 (N_2670,N_2582,N_2587);
or U2671 (N_2671,N_2575,N_2504);
nand U2672 (N_2672,N_2539,N_2512);
or U2673 (N_2673,N_2562,N_2571);
and U2674 (N_2674,N_2552,N_2554);
nor U2675 (N_2675,N_2599,N_2586);
nand U2676 (N_2676,N_2526,N_2590);
or U2677 (N_2677,N_2544,N_2541);
xor U2678 (N_2678,N_2545,N_2585);
nand U2679 (N_2679,N_2588,N_2564);
and U2680 (N_2680,N_2532,N_2522);
and U2681 (N_2681,N_2526,N_2574);
or U2682 (N_2682,N_2597,N_2555);
nor U2683 (N_2683,N_2514,N_2598);
or U2684 (N_2684,N_2535,N_2549);
nand U2685 (N_2685,N_2557,N_2539);
or U2686 (N_2686,N_2592,N_2551);
nor U2687 (N_2687,N_2599,N_2544);
or U2688 (N_2688,N_2589,N_2521);
or U2689 (N_2689,N_2542,N_2538);
and U2690 (N_2690,N_2551,N_2580);
nor U2691 (N_2691,N_2552,N_2526);
nand U2692 (N_2692,N_2585,N_2588);
nand U2693 (N_2693,N_2530,N_2514);
and U2694 (N_2694,N_2564,N_2553);
or U2695 (N_2695,N_2570,N_2521);
and U2696 (N_2696,N_2540,N_2535);
nand U2697 (N_2697,N_2511,N_2503);
and U2698 (N_2698,N_2585,N_2568);
nand U2699 (N_2699,N_2576,N_2523);
xnor U2700 (N_2700,N_2656,N_2676);
nand U2701 (N_2701,N_2648,N_2672);
nor U2702 (N_2702,N_2628,N_2658);
nor U2703 (N_2703,N_2616,N_2650);
nand U2704 (N_2704,N_2694,N_2626);
xor U2705 (N_2705,N_2669,N_2643);
and U2706 (N_2706,N_2634,N_2629);
and U2707 (N_2707,N_2652,N_2620);
nand U2708 (N_2708,N_2660,N_2612);
nor U2709 (N_2709,N_2603,N_2644);
or U2710 (N_2710,N_2680,N_2633);
or U2711 (N_2711,N_2691,N_2601);
or U2712 (N_2712,N_2665,N_2657);
xor U2713 (N_2713,N_2674,N_2614);
or U2714 (N_2714,N_2642,N_2638);
and U2715 (N_2715,N_2627,N_2666);
and U2716 (N_2716,N_2677,N_2622);
nand U2717 (N_2717,N_2687,N_2605);
or U2718 (N_2718,N_2610,N_2697);
nor U2719 (N_2719,N_2623,N_2604);
and U2720 (N_2720,N_2613,N_2690);
or U2721 (N_2721,N_2662,N_2679);
nand U2722 (N_2722,N_2684,N_2671);
and U2723 (N_2723,N_2651,N_2664);
or U2724 (N_2724,N_2632,N_2695);
or U2725 (N_2725,N_2678,N_2608);
nand U2726 (N_2726,N_2646,N_2683);
and U2727 (N_2727,N_2685,N_2673);
or U2728 (N_2728,N_2645,N_2630);
nand U2729 (N_2729,N_2602,N_2631);
xor U2730 (N_2730,N_2667,N_2698);
or U2731 (N_2731,N_2649,N_2692);
or U2732 (N_2732,N_2621,N_2606);
or U2733 (N_2733,N_2615,N_2619);
nor U2734 (N_2734,N_2670,N_2661);
nor U2735 (N_2735,N_2659,N_2607);
or U2736 (N_2736,N_2636,N_2688);
nor U2737 (N_2737,N_2617,N_2693);
nand U2738 (N_2738,N_2609,N_2663);
and U2739 (N_2739,N_2689,N_2635);
nand U2740 (N_2740,N_2639,N_2640);
nor U2741 (N_2741,N_2653,N_2625);
and U2742 (N_2742,N_2600,N_2675);
or U2743 (N_2743,N_2655,N_2647);
xnor U2744 (N_2744,N_2681,N_2611);
or U2745 (N_2745,N_2637,N_2624);
or U2746 (N_2746,N_2668,N_2654);
nor U2747 (N_2747,N_2618,N_2699);
nor U2748 (N_2748,N_2682,N_2641);
nand U2749 (N_2749,N_2686,N_2696);
or U2750 (N_2750,N_2654,N_2685);
nand U2751 (N_2751,N_2689,N_2653);
and U2752 (N_2752,N_2634,N_2627);
nor U2753 (N_2753,N_2632,N_2656);
nand U2754 (N_2754,N_2641,N_2626);
or U2755 (N_2755,N_2650,N_2628);
or U2756 (N_2756,N_2608,N_2612);
or U2757 (N_2757,N_2639,N_2675);
nor U2758 (N_2758,N_2680,N_2681);
and U2759 (N_2759,N_2635,N_2618);
or U2760 (N_2760,N_2607,N_2699);
or U2761 (N_2761,N_2614,N_2628);
nor U2762 (N_2762,N_2618,N_2676);
nor U2763 (N_2763,N_2633,N_2640);
and U2764 (N_2764,N_2667,N_2649);
and U2765 (N_2765,N_2638,N_2686);
nor U2766 (N_2766,N_2685,N_2639);
and U2767 (N_2767,N_2631,N_2611);
or U2768 (N_2768,N_2678,N_2696);
and U2769 (N_2769,N_2655,N_2615);
or U2770 (N_2770,N_2693,N_2600);
or U2771 (N_2771,N_2633,N_2636);
and U2772 (N_2772,N_2642,N_2680);
and U2773 (N_2773,N_2620,N_2699);
nor U2774 (N_2774,N_2669,N_2651);
and U2775 (N_2775,N_2614,N_2690);
nand U2776 (N_2776,N_2640,N_2628);
and U2777 (N_2777,N_2677,N_2656);
and U2778 (N_2778,N_2636,N_2662);
and U2779 (N_2779,N_2614,N_2667);
or U2780 (N_2780,N_2634,N_2674);
and U2781 (N_2781,N_2675,N_2667);
nor U2782 (N_2782,N_2642,N_2648);
or U2783 (N_2783,N_2622,N_2694);
and U2784 (N_2784,N_2638,N_2633);
and U2785 (N_2785,N_2653,N_2621);
and U2786 (N_2786,N_2650,N_2604);
and U2787 (N_2787,N_2685,N_2633);
and U2788 (N_2788,N_2685,N_2619);
and U2789 (N_2789,N_2652,N_2645);
or U2790 (N_2790,N_2645,N_2663);
xnor U2791 (N_2791,N_2669,N_2623);
or U2792 (N_2792,N_2692,N_2603);
or U2793 (N_2793,N_2692,N_2698);
nor U2794 (N_2794,N_2635,N_2625);
nand U2795 (N_2795,N_2670,N_2607);
or U2796 (N_2796,N_2648,N_2624);
or U2797 (N_2797,N_2661,N_2697);
nand U2798 (N_2798,N_2652,N_2695);
nor U2799 (N_2799,N_2635,N_2602);
and U2800 (N_2800,N_2770,N_2779);
nor U2801 (N_2801,N_2731,N_2746);
and U2802 (N_2802,N_2751,N_2726);
or U2803 (N_2803,N_2713,N_2782);
and U2804 (N_2804,N_2734,N_2787);
or U2805 (N_2805,N_2703,N_2774);
and U2806 (N_2806,N_2760,N_2759);
and U2807 (N_2807,N_2743,N_2771);
nand U2808 (N_2808,N_2710,N_2748);
nor U2809 (N_2809,N_2785,N_2772);
and U2810 (N_2810,N_2775,N_2733);
or U2811 (N_2811,N_2777,N_2725);
or U2812 (N_2812,N_2739,N_2730);
nand U2813 (N_2813,N_2780,N_2783);
and U2814 (N_2814,N_2702,N_2718);
or U2815 (N_2815,N_2767,N_2752);
nand U2816 (N_2816,N_2724,N_2778);
or U2817 (N_2817,N_2719,N_2728);
and U2818 (N_2818,N_2792,N_2722);
and U2819 (N_2819,N_2764,N_2788);
or U2820 (N_2820,N_2784,N_2756);
nor U2821 (N_2821,N_2727,N_2737);
and U2822 (N_2822,N_2796,N_2773);
and U2823 (N_2823,N_2706,N_2745);
and U2824 (N_2824,N_2712,N_2729);
nand U2825 (N_2825,N_2735,N_2750);
xnor U2826 (N_2826,N_2701,N_2758);
nor U2827 (N_2827,N_2740,N_2742);
and U2828 (N_2828,N_2769,N_2762);
nor U2829 (N_2829,N_2716,N_2736);
xnor U2830 (N_2830,N_2754,N_2793);
nor U2831 (N_2831,N_2708,N_2747);
xor U2832 (N_2832,N_2781,N_2757);
and U2833 (N_2833,N_2753,N_2797);
and U2834 (N_2834,N_2700,N_2749);
nor U2835 (N_2835,N_2709,N_2776);
and U2836 (N_2836,N_2714,N_2798);
and U2837 (N_2837,N_2738,N_2715);
nand U2838 (N_2838,N_2723,N_2721);
xnor U2839 (N_2839,N_2755,N_2744);
nor U2840 (N_2840,N_2766,N_2794);
and U2841 (N_2841,N_2707,N_2720);
nand U2842 (N_2842,N_2705,N_2732);
nor U2843 (N_2843,N_2741,N_2717);
nor U2844 (N_2844,N_2790,N_2786);
and U2845 (N_2845,N_2768,N_2795);
nor U2846 (N_2846,N_2765,N_2711);
and U2847 (N_2847,N_2791,N_2763);
and U2848 (N_2848,N_2789,N_2704);
and U2849 (N_2849,N_2799,N_2761);
and U2850 (N_2850,N_2701,N_2742);
and U2851 (N_2851,N_2740,N_2769);
and U2852 (N_2852,N_2708,N_2784);
or U2853 (N_2853,N_2757,N_2787);
and U2854 (N_2854,N_2705,N_2763);
nand U2855 (N_2855,N_2761,N_2778);
and U2856 (N_2856,N_2740,N_2705);
nand U2857 (N_2857,N_2709,N_2734);
xnor U2858 (N_2858,N_2751,N_2712);
nand U2859 (N_2859,N_2706,N_2722);
nor U2860 (N_2860,N_2796,N_2725);
nor U2861 (N_2861,N_2701,N_2712);
nor U2862 (N_2862,N_2716,N_2738);
xnor U2863 (N_2863,N_2712,N_2775);
nor U2864 (N_2864,N_2771,N_2726);
xnor U2865 (N_2865,N_2791,N_2784);
and U2866 (N_2866,N_2792,N_2714);
or U2867 (N_2867,N_2794,N_2799);
nor U2868 (N_2868,N_2744,N_2782);
and U2869 (N_2869,N_2792,N_2777);
or U2870 (N_2870,N_2767,N_2726);
and U2871 (N_2871,N_2750,N_2708);
or U2872 (N_2872,N_2761,N_2796);
or U2873 (N_2873,N_2771,N_2763);
or U2874 (N_2874,N_2735,N_2729);
or U2875 (N_2875,N_2771,N_2792);
and U2876 (N_2876,N_2754,N_2779);
and U2877 (N_2877,N_2781,N_2775);
nand U2878 (N_2878,N_2742,N_2717);
xor U2879 (N_2879,N_2788,N_2706);
or U2880 (N_2880,N_2755,N_2793);
and U2881 (N_2881,N_2796,N_2753);
and U2882 (N_2882,N_2762,N_2740);
and U2883 (N_2883,N_2733,N_2797);
nor U2884 (N_2884,N_2771,N_2772);
or U2885 (N_2885,N_2799,N_2714);
or U2886 (N_2886,N_2776,N_2741);
and U2887 (N_2887,N_2759,N_2719);
and U2888 (N_2888,N_2750,N_2776);
or U2889 (N_2889,N_2720,N_2775);
and U2890 (N_2890,N_2792,N_2737);
and U2891 (N_2891,N_2736,N_2772);
xor U2892 (N_2892,N_2743,N_2755);
and U2893 (N_2893,N_2732,N_2771);
or U2894 (N_2894,N_2725,N_2732);
nand U2895 (N_2895,N_2718,N_2794);
nor U2896 (N_2896,N_2776,N_2793);
nor U2897 (N_2897,N_2719,N_2783);
and U2898 (N_2898,N_2784,N_2753);
and U2899 (N_2899,N_2735,N_2761);
or U2900 (N_2900,N_2839,N_2853);
nor U2901 (N_2901,N_2809,N_2808);
nand U2902 (N_2902,N_2817,N_2866);
nor U2903 (N_2903,N_2802,N_2896);
nor U2904 (N_2904,N_2859,N_2814);
nor U2905 (N_2905,N_2882,N_2849);
nand U2906 (N_2906,N_2836,N_2891);
nor U2907 (N_2907,N_2824,N_2845);
or U2908 (N_2908,N_2880,N_2816);
nor U2909 (N_2909,N_2804,N_2870);
nor U2910 (N_2910,N_2848,N_2864);
nand U2911 (N_2911,N_2846,N_2831);
nand U2912 (N_2912,N_2835,N_2803);
or U2913 (N_2913,N_2861,N_2884);
nand U2914 (N_2914,N_2872,N_2813);
nor U2915 (N_2915,N_2879,N_2843);
nand U2916 (N_2916,N_2838,N_2842);
and U2917 (N_2917,N_2885,N_2888);
and U2918 (N_2918,N_2818,N_2810);
or U2919 (N_2919,N_2867,N_2869);
or U2920 (N_2920,N_2822,N_2847);
nor U2921 (N_2921,N_2854,N_2889);
nand U2922 (N_2922,N_2815,N_2890);
nand U2923 (N_2923,N_2819,N_2881);
nor U2924 (N_2924,N_2830,N_2823);
nand U2925 (N_2925,N_2865,N_2828);
nand U2926 (N_2926,N_2820,N_2851);
xnor U2927 (N_2927,N_2898,N_2878);
nor U2928 (N_2928,N_2873,N_2844);
or U2929 (N_2929,N_2886,N_2801);
and U2930 (N_2930,N_2857,N_2893);
nor U2931 (N_2931,N_2821,N_2834);
and U2932 (N_2932,N_2840,N_2811);
nand U2933 (N_2933,N_2895,N_2825);
nand U2934 (N_2934,N_2856,N_2860);
nor U2935 (N_2935,N_2805,N_2899);
nor U2936 (N_2936,N_2841,N_2827);
or U2937 (N_2937,N_2800,N_2807);
nor U2938 (N_2938,N_2876,N_2858);
nand U2939 (N_2939,N_2852,N_2877);
or U2940 (N_2940,N_2833,N_2826);
xor U2941 (N_2941,N_2894,N_2862);
and U2942 (N_2942,N_2874,N_2868);
nand U2943 (N_2943,N_2832,N_2875);
and U2944 (N_2944,N_2829,N_2837);
or U2945 (N_2945,N_2883,N_2892);
nor U2946 (N_2946,N_2806,N_2850);
nand U2947 (N_2947,N_2897,N_2887);
nand U2948 (N_2948,N_2855,N_2871);
and U2949 (N_2949,N_2863,N_2812);
and U2950 (N_2950,N_2883,N_2804);
or U2951 (N_2951,N_2843,N_2871);
nand U2952 (N_2952,N_2820,N_2810);
and U2953 (N_2953,N_2848,N_2899);
nand U2954 (N_2954,N_2804,N_2871);
nand U2955 (N_2955,N_2817,N_2872);
nand U2956 (N_2956,N_2853,N_2832);
and U2957 (N_2957,N_2890,N_2848);
nor U2958 (N_2958,N_2829,N_2864);
xnor U2959 (N_2959,N_2861,N_2831);
or U2960 (N_2960,N_2882,N_2879);
nand U2961 (N_2961,N_2842,N_2809);
nand U2962 (N_2962,N_2815,N_2834);
and U2963 (N_2963,N_2802,N_2885);
and U2964 (N_2964,N_2881,N_2806);
and U2965 (N_2965,N_2872,N_2810);
nand U2966 (N_2966,N_2800,N_2836);
nor U2967 (N_2967,N_2857,N_2844);
or U2968 (N_2968,N_2861,N_2830);
and U2969 (N_2969,N_2887,N_2826);
nand U2970 (N_2970,N_2805,N_2870);
or U2971 (N_2971,N_2829,N_2807);
nand U2972 (N_2972,N_2800,N_2824);
or U2973 (N_2973,N_2813,N_2824);
nand U2974 (N_2974,N_2811,N_2832);
and U2975 (N_2975,N_2820,N_2845);
nor U2976 (N_2976,N_2837,N_2801);
nand U2977 (N_2977,N_2880,N_2874);
nor U2978 (N_2978,N_2856,N_2889);
and U2979 (N_2979,N_2824,N_2872);
and U2980 (N_2980,N_2860,N_2845);
nor U2981 (N_2981,N_2801,N_2810);
or U2982 (N_2982,N_2866,N_2841);
or U2983 (N_2983,N_2825,N_2882);
nor U2984 (N_2984,N_2833,N_2863);
nand U2985 (N_2985,N_2862,N_2842);
nor U2986 (N_2986,N_2829,N_2813);
and U2987 (N_2987,N_2811,N_2845);
or U2988 (N_2988,N_2817,N_2844);
nor U2989 (N_2989,N_2800,N_2853);
or U2990 (N_2990,N_2806,N_2871);
nand U2991 (N_2991,N_2827,N_2829);
or U2992 (N_2992,N_2865,N_2866);
and U2993 (N_2993,N_2874,N_2839);
and U2994 (N_2994,N_2871,N_2863);
and U2995 (N_2995,N_2815,N_2875);
nor U2996 (N_2996,N_2829,N_2845);
and U2997 (N_2997,N_2868,N_2851);
and U2998 (N_2998,N_2808,N_2836);
nor U2999 (N_2999,N_2845,N_2881);
nor U3000 (N_3000,N_2927,N_2901);
or U3001 (N_3001,N_2923,N_2904);
nand U3002 (N_3002,N_2993,N_2972);
nand U3003 (N_3003,N_2952,N_2996);
nor U3004 (N_3004,N_2917,N_2987);
or U3005 (N_3005,N_2982,N_2935);
nor U3006 (N_3006,N_2941,N_2948);
or U3007 (N_3007,N_2929,N_2943);
nand U3008 (N_3008,N_2937,N_2980);
and U3009 (N_3009,N_2950,N_2953);
nand U3010 (N_3010,N_2958,N_2969);
nand U3011 (N_3011,N_2954,N_2946);
or U3012 (N_3012,N_2947,N_2979);
or U3013 (N_3013,N_2903,N_2949);
nor U3014 (N_3014,N_2914,N_2936);
and U3015 (N_3015,N_2930,N_2959);
or U3016 (N_3016,N_2918,N_2964);
and U3017 (N_3017,N_2989,N_2926);
or U3018 (N_3018,N_2921,N_2990);
and U3019 (N_3019,N_2939,N_2933);
or U3020 (N_3020,N_2934,N_2966);
nand U3021 (N_3021,N_2957,N_2945);
nor U3022 (N_3022,N_2922,N_2913);
and U3023 (N_3023,N_2944,N_2960);
nand U3024 (N_3024,N_2955,N_2916);
nor U3025 (N_3025,N_2974,N_2909);
nor U3026 (N_3026,N_2942,N_2977);
and U3027 (N_3027,N_2907,N_2919);
and U3028 (N_3028,N_2992,N_2984);
and U3029 (N_3029,N_2962,N_2976);
and U3030 (N_3030,N_2900,N_2998);
xnor U3031 (N_3031,N_2970,N_2975);
nor U3032 (N_3032,N_2985,N_2905);
and U3033 (N_3033,N_2915,N_2994);
nor U3034 (N_3034,N_2995,N_2908);
and U3035 (N_3035,N_2986,N_2911);
nand U3036 (N_3036,N_2910,N_2931);
nand U3037 (N_3037,N_2940,N_2906);
nand U3038 (N_3038,N_2912,N_2956);
or U3039 (N_3039,N_2932,N_2968);
nor U3040 (N_3040,N_2991,N_2973);
and U3041 (N_3041,N_2920,N_2988);
nor U3042 (N_3042,N_2978,N_2925);
and U3043 (N_3043,N_2999,N_2902);
and U3044 (N_3044,N_2983,N_2951);
nor U3045 (N_3045,N_2981,N_2924);
nor U3046 (N_3046,N_2997,N_2971);
nor U3047 (N_3047,N_2938,N_2961);
nor U3048 (N_3048,N_2965,N_2928);
nor U3049 (N_3049,N_2963,N_2967);
or U3050 (N_3050,N_2961,N_2963);
and U3051 (N_3051,N_2966,N_2919);
nand U3052 (N_3052,N_2946,N_2927);
and U3053 (N_3053,N_2980,N_2958);
nor U3054 (N_3054,N_2979,N_2965);
nor U3055 (N_3055,N_2902,N_2974);
or U3056 (N_3056,N_2992,N_2994);
nand U3057 (N_3057,N_2920,N_2952);
nand U3058 (N_3058,N_2957,N_2950);
or U3059 (N_3059,N_2956,N_2966);
or U3060 (N_3060,N_2957,N_2909);
or U3061 (N_3061,N_2979,N_2985);
and U3062 (N_3062,N_2961,N_2995);
and U3063 (N_3063,N_2966,N_2998);
nand U3064 (N_3064,N_2980,N_2944);
nor U3065 (N_3065,N_2986,N_2966);
nand U3066 (N_3066,N_2999,N_2951);
and U3067 (N_3067,N_2977,N_2918);
nand U3068 (N_3068,N_2964,N_2976);
nor U3069 (N_3069,N_2981,N_2986);
nand U3070 (N_3070,N_2969,N_2997);
and U3071 (N_3071,N_2937,N_2993);
nor U3072 (N_3072,N_2945,N_2962);
or U3073 (N_3073,N_2934,N_2918);
nor U3074 (N_3074,N_2901,N_2980);
nand U3075 (N_3075,N_2968,N_2977);
or U3076 (N_3076,N_2963,N_2947);
and U3077 (N_3077,N_2901,N_2984);
nand U3078 (N_3078,N_2914,N_2916);
nand U3079 (N_3079,N_2968,N_2922);
nand U3080 (N_3080,N_2949,N_2969);
nand U3081 (N_3081,N_2982,N_2946);
nand U3082 (N_3082,N_2996,N_2975);
and U3083 (N_3083,N_2954,N_2902);
nor U3084 (N_3084,N_2985,N_2934);
nor U3085 (N_3085,N_2954,N_2973);
nor U3086 (N_3086,N_2998,N_2994);
or U3087 (N_3087,N_2935,N_2991);
and U3088 (N_3088,N_2986,N_2922);
nand U3089 (N_3089,N_2991,N_2931);
or U3090 (N_3090,N_2997,N_2941);
nand U3091 (N_3091,N_2937,N_2949);
nand U3092 (N_3092,N_2931,N_2944);
and U3093 (N_3093,N_2996,N_2955);
and U3094 (N_3094,N_2998,N_2905);
nor U3095 (N_3095,N_2996,N_2986);
or U3096 (N_3096,N_2984,N_2994);
nor U3097 (N_3097,N_2935,N_2912);
xor U3098 (N_3098,N_2928,N_2996);
and U3099 (N_3099,N_2961,N_2958);
and U3100 (N_3100,N_3013,N_3003);
nor U3101 (N_3101,N_3048,N_3002);
nor U3102 (N_3102,N_3053,N_3089);
or U3103 (N_3103,N_3059,N_3010);
nand U3104 (N_3104,N_3087,N_3097);
or U3105 (N_3105,N_3072,N_3090);
and U3106 (N_3106,N_3026,N_3061);
nand U3107 (N_3107,N_3025,N_3065);
and U3108 (N_3108,N_3024,N_3008);
and U3109 (N_3109,N_3028,N_3030);
or U3110 (N_3110,N_3088,N_3098);
or U3111 (N_3111,N_3068,N_3005);
nor U3112 (N_3112,N_3034,N_3091);
or U3113 (N_3113,N_3044,N_3071);
and U3114 (N_3114,N_3076,N_3085);
or U3115 (N_3115,N_3094,N_3075);
nor U3116 (N_3116,N_3058,N_3062);
nand U3117 (N_3117,N_3055,N_3095);
nor U3118 (N_3118,N_3016,N_3079);
nor U3119 (N_3119,N_3036,N_3096);
nand U3120 (N_3120,N_3007,N_3080);
nand U3121 (N_3121,N_3049,N_3021);
nor U3122 (N_3122,N_3033,N_3018);
and U3123 (N_3123,N_3015,N_3099);
or U3124 (N_3124,N_3066,N_3035);
or U3125 (N_3125,N_3063,N_3052);
nand U3126 (N_3126,N_3029,N_3084);
nor U3127 (N_3127,N_3064,N_3041);
and U3128 (N_3128,N_3039,N_3086);
nor U3129 (N_3129,N_3037,N_3093);
and U3130 (N_3130,N_3078,N_3040);
or U3131 (N_3131,N_3043,N_3092);
nand U3132 (N_3132,N_3023,N_3032);
and U3133 (N_3133,N_3014,N_3054);
or U3134 (N_3134,N_3017,N_3022);
and U3135 (N_3135,N_3050,N_3046);
or U3136 (N_3136,N_3047,N_3011);
and U3137 (N_3137,N_3057,N_3082);
nand U3138 (N_3138,N_3000,N_3019);
and U3139 (N_3139,N_3009,N_3051);
and U3140 (N_3140,N_3006,N_3081);
nor U3141 (N_3141,N_3001,N_3031);
or U3142 (N_3142,N_3074,N_3060);
and U3143 (N_3143,N_3004,N_3056);
nand U3144 (N_3144,N_3020,N_3038);
and U3145 (N_3145,N_3027,N_3067);
or U3146 (N_3146,N_3077,N_3083);
nand U3147 (N_3147,N_3073,N_3012);
nand U3148 (N_3148,N_3045,N_3070);
or U3149 (N_3149,N_3069,N_3042);
xnor U3150 (N_3150,N_3032,N_3083);
nand U3151 (N_3151,N_3094,N_3002);
nor U3152 (N_3152,N_3095,N_3043);
or U3153 (N_3153,N_3057,N_3064);
nor U3154 (N_3154,N_3005,N_3022);
and U3155 (N_3155,N_3062,N_3020);
nand U3156 (N_3156,N_3085,N_3034);
or U3157 (N_3157,N_3008,N_3047);
nor U3158 (N_3158,N_3092,N_3019);
nor U3159 (N_3159,N_3099,N_3023);
nand U3160 (N_3160,N_3080,N_3071);
nand U3161 (N_3161,N_3067,N_3082);
or U3162 (N_3162,N_3059,N_3092);
nor U3163 (N_3163,N_3067,N_3080);
xor U3164 (N_3164,N_3015,N_3044);
or U3165 (N_3165,N_3008,N_3023);
or U3166 (N_3166,N_3093,N_3068);
nand U3167 (N_3167,N_3012,N_3023);
and U3168 (N_3168,N_3001,N_3028);
nand U3169 (N_3169,N_3040,N_3042);
or U3170 (N_3170,N_3089,N_3000);
and U3171 (N_3171,N_3067,N_3028);
or U3172 (N_3172,N_3099,N_3065);
nor U3173 (N_3173,N_3084,N_3044);
xor U3174 (N_3174,N_3099,N_3004);
or U3175 (N_3175,N_3033,N_3020);
xor U3176 (N_3176,N_3074,N_3065);
nor U3177 (N_3177,N_3081,N_3048);
nor U3178 (N_3178,N_3073,N_3077);
nand U3179 (N_3179,N_3020,N_3037);
nand U3180 (N_3180,N_3070,N_3023);
or U3181 (N_3181,N_3015,N_3032);
nand U3182 (N_3182,N_3037,N_3014);
nand U3183 (N_3183,N_3086,N_3016);
and U3184 (N_3184,N_3067,N_3012);
nor U3185 (N_3185,N_3074,N_3069);
nand U3186 (N_3186,N_3008,N_3027);
nand U3187 (N_3187,N_3098,N_3064);
nand U3188 (N_3188,N_3041,N_3075);
nor U3189 (N_3189,N_3058,N_3045);
and U3190 (N_3190,N_3071,N_3003);
or U3191 (N_3191,N_3037,N_3016);
xor U3192 (N_3192,N_3039,N_3006);
and U3193 (N_3193,N_3002,N_3008);
and U3194 (N_3194,N_3006,N_3040);
or U3195 (N_3195,N_3021,N_3095);
and U3196 (N_3196,N_3041,N_3037);
or U3197 (N_3197,N_3000,N_3009);
nand U3198 (N_3198,N_3032,N_3056);
and U3199 (N_3199,N_3081,N_3012);
and U3200 (N_3200,N_3143,N_3108);
nand U3201 (N_3201,N_3150,N_3188);
nor U3202 (N_3202,N_3138,N_3177);
or U3203 (N_3203,N_3128,N_3130);
nand U3204 (N_3204,N_3148,N_3184);
or U3205 (N_3205,N_3124,N_3175);
and U3206 (N_3206,N_3107,N_3163);
or U3207 (N_3207,N_3176,N_3145);
nand U3208 (N_3208,N_3197,N_3117);
nor U3209 (N_3209,N_3137,N_3144);
or U3210 (N_3210,N_3136,N_3127);
and U3211 (N_3211,N_3139,N_3141);
and U3212 (N_3212,N_3102,N_3140);
nor U3213 (N_3213,N_3114,N_3160);
nand U3214 (N_3214,N_3164,N_3103);
nor U3215 (N_3215,N_3166,N_3178);
and U3216 (N_3216,N_3121,N_3129);
nor U3217 (N_3217,N_3158,N_3119);
xor U3218 (N_3218,N_3134,N_3192);
nor U3219 (N_3219,N_3161,N_3171);
nor U3220 (N_3220,N_3151,N_3187);
or U3221 (N_3221,N_3104,N_3106);
nand U3222 (N_3222,N_3155,N_3168);
and U3223 (N_3223,N_3181,N_3154);
xor U3224 (N_3224,N_3198,N_3186);
and U3225 (N_3225,N_3147,N_3170);
nand U3226 (N_3226,N_3116,N_3169);
nor U3227 (N_3227,N_3112,N_3189);
nor U3228 (N_3228,N_3142,N_3133);
and U3229 (N_3229,N_3105,N_3159);
or U3230 (N_3230,N_3149,N_3174);
nand U3231 (N_3231,N_3180,N_3111);
and U3232 (N_3232,N_3100,N_3199);
nand U3233 (N_3233,N_3183,N_3185);
or U3234 (N_3234,N_3182,N_3162);
and U3235 (N_3235,N_3156,N_3190);
or U3236 (N_3236,N_3123,N_3157);
or U3237 (N_3237,N_3135,N_3165);
or U3238 (N_3238,N_3131,N_3173);
nor U3239 (N_3239,N_3167,N_3110);
nor U3240 (N_3240,N_3109,N_3126);
nand U3241 (N_3241,N_3196,N_3118);
and U3242 (N_3242,N_3101,N_3146);
nor U3243 (N_3243,N_3195,N_3132);
or U3244 (N_3244,N_3113,N_3191);
nand U3245 (N_3245,N_3153,N_3115);
nor U3246 (N_3246,N_3172,N_3179);
or U3247 (N_3247,N_3122,N_3193);
nand U3248 (N_3248,N_3120,N_3125);
nand U3249 (N_3249,N_3152,N_3194);
or U3250 (N_3250,N_3193,N_3118);
nor U3251 (N_3251,N_3181,N_3170);
or U3252 (N_3252,N_3131,N_3122);
nor U3253 (N_3253,N_3151,N_3102);
nand U3254 (N_3254,N_3175,N_3128);
nand U3255 (N_3255,N_3198,N_3113);
or U3256 (N_3256,N_3158,N_3157);
nand U3257 (N_3257,N_3111,N_3166);
nor U3258 (N_3258,N_3187,N_3197);
nand U3259 (N_3259,N_3149,N_3108);
and U3260 (N_3260,N_3109,N_3134);
or U3261 (N_3261,N_3145,N_3198);
nand U3262 (N_3262,N_3134,N_3196);
nor U3263 (N_3263,N_3137,N_3160);
nor U3264 (N_3264,N_3117,N_3114);
or U3265 (N_3265,N_3130,N_3162);
nand U3266 (N_3266,N_3173,N_3164);
nor U3267 (N_3267,N_3135,N_3172);
nor U3268 (N_3268,N_3195,N_3180);
nor U3269 (N_3269,N_3162,N_3169);
or U3270 (N_3270,N_3123,N_3109);
or U3271 (N_3271,N_3185,N_3108);
or U3272 (N_3272,N_3131,N_3160);
and U3273 (N_3273,N_3126,N_3189);
and U3274 (N_3274,N_3175,N_3166);
or U3275 (N_3275,N_3166,N_3115);
or U3276 (N_3276,N_3185,N_3131);
nor U3277 (N_3277,N_3115,N_3138);
or U3278 (N_3278,N_3158,N_3189);
and U3279 (N_3279,N_3184,N_3174);
nor U3280 (N_3280,N_3169,N_3125);
and U3281 (N_3281,N_3198,N_3168);
nor U3282 (N_3282,N_3145,N_3117);
or U3283 (N_3283,N_3159,N_3111);
nand U3284 (N_3284,N_3193,N_3197);
nand U3285 (N_3285,N_3179,N_3136);
or U3286 (N_3286,N_3182,N_3177);
nor U3287 (N_3287,N_3183,N_3166);
and U3288 (N_3288,N_3117,N_3184);
or U3289 (N_3289,N_3127,N_3178);
xor U3290 (N_3290,N_3159,N_3173);
nor U3291 (N_3291,N_3169,N_3124);
and U3292 (N_3292,N_3187,N_3116);
nand U3293 (N_3293,N_3111,N_3171);
xor U3294 (N_3294,N_3198,N_3103);
and U3295 (N_3295,N_3198,N_3107);
or U3296 (N_3296,N_3145,N_3128);
or U3297 (N_3297,N_3113,N_3199);
nor U3298 (N_3298,N_3129,N_3180);
nand U3299 (N_3299,N_3125,N_3135);
nor U3300 (N_3300,N_3225,N_3206);
nand U3301 (N_3301,N_3228,N_3258);
or U3302 (N_3302,N_3254,N_3253);
nor U3303 (N_3303,N_3249,N_3292);
or U3304 (N_3304,N_3239,N_3278);
and U3305 (N_3305,N_3209,N_3299);
and U3306 (N_3306,N_3281,N_3240);
and U3307 (N_3307,N_3263,N_3286);
and U3308 (N_3308,N_3247,N_3270);
nand U3309 (N_3309,N_3262,N_3208);
and U3310 (N_3310,N_3274,N_3212);
and U3311 (N_3311,N_3227,N_3229);
nor U3312 (N_3312,N_3238,N_3213);
nor U3313 (N_3313,N_3244,N_3207);
and U3314 (N_3314,N_3211,N_3214);
or U3315 (N_3315,N_3216,N_3260);
nor U3316 (N_3316,N_3268,N_3275);
or U3317 (N_3317,N_3266,N_3203);
nor U3318 (N_3318,N_3201,N_3220);
and U3319 (N_3319,N_3288,N_3200);
and U3320 (N_3320,N_3255,N_3218);
or U3321 (N_3321,N_3232,N_3222);
nand U3322 (N_3322,N_3280,N_3265);
nand U3323 (N_3323,N_3269,N_3248);
and U3324 (N_3324,N_3271,N_3272);
nor U3325 (N_3325,N_3293,N_3287);
nand U3326 (N_3326,N_3285,N_3221);
nand U3327 (N_3327,N_3283,N_3250);
and U3328 (N_3328,N_3282,N_3224);
or U3329 (N_3329,N_3252,N_3291);
xor U3330 (N_3330,N_3277,N_3245);
nor U3331 (N_3331,N_3242,N_3294);
nand U3332 (N_3332,N_3296,N_3290);
nor U3333 (N_3333,N_3241,N_3289);
nand U3334 (N_3334,N_3273,N_3267);
nor U3335 (N_3335,N_3257,N_3215);
nor U3336 (N_3336,N_3233,N_3231);
or U3337 (N_3337,N_3217,N_3276);
or U3338 (N_3338,N_3205,N_3295);
nor U3339 (N_3339,N_3210,N_3279);
nor U3340 (N_3340,N_3219,N_3246);
and U3341 (N_3341,N_3237,N_3264);
nor U3342 (N_3342,N_3256,N_3284);
nand U3343 (N_3343,N_3243,N_3234);
nand U3344 (N_3344,N_3226,N_3204);
or U3345 (N_3345,N_3202,N_3236);
or U3346 (N_3346,N_3259,N_3298);
and U3347 (N_3347,N_3251,N_3223);
nand U3348 (N_3348,N_3235,N_3297);
and U3349 (N_3349,N_3261,N_3230);
nor U3350 (N_3350,N_3282,N_3262);
and U3351 (N_3351,N_3235,N_3242);
nor U3352 (N_3352,N_3275,N_3259);
nand U3353 (N_3353,N_3259,N_3268);
nand U3354 (N_3354,N_3227,N_3266);
or U3355 (N_3355,N_3296,N_3288);
nor U3356 (N_3356,N_3206,N_3294);
or U3357 (N_3357,N_3205,N_3246);
nand U3358 (N_3358,N_3211,N_3296);
nand U3359 (N_3359,N_3277,N_3269);
or U3360 (N_3360,N_3265,N_3270);
nor U3361 (N_3361,N_3250,N_3245);
nor U3362 (N_3362,N_3282,N_3221);
nor U3363 (N_3363,N_3226,N_3297);
nor U3364 (N_3364,N_3246,N_3291);
or U3365 (N_3365,N_3281,N_3244);
or U3366 (N_3366,N_3276,N_3252);
nand U3367 (N_3367,N_3211,N_3290);
nand U3368 (N_3368,N_3217,N_3234);
and U3369 (N_3369,N_3239,N_3277);
and U3370 (N_3370,N_3295,N_3297);
and U3371 (N_3371,N_3254,N_3299);
or U3372 (N_3372,N_3217,N_3202);
nand U3373 (N_3373,N_3277,N_3247);
nor U3374 (N_3374,N_3281,N_3291);
nor U3375 (N_3375,N_3297,N_3233);
nor U3376 (N_3376,N_3257,N_3223);
nand U3377 (N_3377,N_3257,N_3222);
nor U3378 (N_3378,N_3288,N_3268);
nor U3379 (N_3379,N_3270,N_3207);
nor U3380 (N_3380,N_3287,N_3226);
and U3381 (N_3381,N_3289,N_3233);
nor U3382 (N_3382,N_3201,N_3275);
xnor U3383 (N_3383,N_3217,N_3203);
or U3384 (N_3384,N_3250,N_3268);
or U3385 (N_3385,N_3272,N_3206);
nor U3386 (N_3386,N_3229,N_3290);
nand U3387 (N_3387,N_3255,N_3252);
and U3388 (N_3388,N_3296,N_3221);
nor U3389 (N_3389,N_3270,N_3250);
or U3390 (N_3390,N_3210,N_3257);
nand U3391 (N_3391,N_3210,N_3225);
or U3392 (N_3392,N_3223,N_3205);
nor U3393 (N_3393,N_3206,N_3221);
or U3394 (N_3394,N_3248,N_3212);
nor U3395 (N_3395,N_3290,N_3200);
nand U3396 (N_3396,N_3229,N_3270);
xnor U3397 (N_3397,N_3254,N_3281);
and U3398 (N_3398,N_3245,N_3201);
or U3399 (N_3399,N_3246,N_3296);
or U3400 (N_3400,N_3387,N_3320);
nor U3401 (N_3401,N_3304,N_3355);
or U3402 (N_3402,N_3371,N_3341);
and U3403 (N_3403,N_3345,N_3386);
nor U3404 (N_3404,N_3366,N_3312);
and U3405 (N_3405,N_3358,N_3305);
or U3406 (N_3406,N_3310,N_3379);
or U3407 (N_3407,N_3364,N_3350);
or U3408 (N_3408,N_3382,N_3331);
nor U3409 (N_3409,N_3370,N_3389);
or U3410 (N_3410,N_3325,N_3314);
and U3411 (N_3411,N_3353,N_3330);
and U3412 (N_3412,N_3322,N_3388);
or U3413 (N_3413,N_3321,N_3380);
nor U3414 (N_3414,N_3339,N_3391);
and U3415 (N_3415,N_3334,N_3396);
and U3416 (N_3416,N_3363,N_3324);
or U3417 (N_3417,N_3375,N_3395);
nand U3418 (N_3418,N_3369,N_3394);
nand U3419 (N_3419,N_3327,N_3354);
or U3420 (N_3420,N_3313,N_3337);
and U3421 (N_3421,N_3378,N_3311);
nand U3422 (N_3422,N_3392,N_3309);
or U3423 (N_3423,N_3372,N_3376);
nand U3424 (N_3424,N_3343,N_3374);
xor U3425 (N_3425,N_3317,N_3347);
nand U3426 (N_3426,N_3373,N_3368);
or U3427 (N_3427,N_3359,N_3316);
and U3428 (N_3428,N_3361,N_3381);
or U3429 (N_3429,N_3319,N_3344);
and U3430 (N_3430,N_3326,N_3315);
or U3431 (N_3431,N_3360,N_3333);
nand U3432 (N_3432,N_3340,N_3335);
or U3433 (N_3433,N_3346,N_3328);
or U3434 (N_3434,N_3377,N_3351);
or U3435 (N_3435,N_3362,N_3342);
and U3436 (N_3436,N_3329,N_3332);
nand U3437 (N_3437,N_3398,N_3307);
nand U3438 (N_3438,N_3399,N_3301);
nand U3439 (N_3439,N_3318,N_3300);
or U3440 (N_3440,N_3336,N_3349);
or U3441 (N_3441,N_3306,N_3367);
nor U3442 (N_3442,N_3302,N_3390);
nor U3443 (N_3443,N_3348,N_3385);
nand U3444 (N_3444,N_3308,N_3384);
and U3445 (N_3445,N_3352,N_3323);
nand U3446 (N_3446,N_3357,N_3365);
nand U3447 (N_3447,N_3356,N_3397);
or U3448 (N_3448,N_3383,N_3338);
nor U3449 (N_3449,N_3303,N_3393);
nand U3450 (N_3450,N_3302,N_3307);
nor U3451 (N_3451,N_3377,N_3364);
nor U3452 (N_3452,N_3360,N_3326);
nor U3453 (N_3453,N_3336,N_3382);
and U3454 (N_3454,N_3393,N_3380);
or U3455 (N_3455,N_3318,N_3314);
nor U3456 (N_3456,N_3324,N_3367);
nand U3457 (N_3457,N_3326,N_3323);
nor U3458 (N_3458,N_3317,N_3319);
or U3459 (N_3459,N_3332,N_3315);
nand U3460 (N_3460,N_3379,N_3346);
or U3461 (N_3461,N_3303,N_3353);
and U3462 (N_3462,N_3316,N_3312);
and U3463 (N_3463,N_3340,N_3323);
nand U3464 (N_3464,N_3361,N_3344);
or U3465 (N_3465,N_3389,N_3317);
and U3466 (N_3466,N_3314,N_3340);
xnor U3467 (N_3467,N_3377,N_3321);
nor U3468 (N_3468,N_3311,N_3344);
and U3469 (N_3469,N_3309,N_3305);
or U3470 (N_3470,N_3357,N_3319);
or U3471 (N_3471,N_3327,N_3340);
or U3472 (N_3472,N_3344,N_3314);
nor U3473 (N_3473,N_3352,N_3373);
and U3474 (N_3474,N_3324,N_3373);
nor U3475 (N_3475,N_3360,N_3355);
or U3476 (N_3476,N_3397,N_3310);
nand U3477 (N_3477,N_3366,N_3342);
and U3478 (N_3478,N_3342,N_3381);
nand U3479 (N_3479,N_3332,N_3316);
and U3480 (N_3480,N_3395,N_3354);
nand U3481 (N_3481,N_3346,N_3353);
or U3482 (N_3482,N_3328,N_3365);
nor U3483 (N_3483,N_3338,N_3315);
nand U3484 (N_3484,N_3396,N_3391);
nand U3485 (N_3485,N_3359,N_3342);
nor U3486 (N_3486,N_3358,N_3307);
nand U3487 (N_3487,N_3326,N_3335);
nor U3488 (N_3488,N_3396,N_3307);
nor U3489 (N_3489,N_3351,N_3335);
nor U3490 (N_3490,N_3339,N_3303);
or U3491 (N_3491,N_3393,N_3364);
and U3492 (N_3492,N_3371,N_3325);
nand U3493 (N_3493,N_3372,N_3379);
or U3494 (N_3494,N_3386,N_3340);
nor U3495 (N_3495,N_3311,N_3353);
nor U3496 (N_3496,N_3301,N_3306);
nor U3497 (N_3497,N_3354,N_3387);
and U3498 (N_3498,N_3335,N_3385);
and U3499 (N_3499,N_3385,N_3301);
and U3500 (N_3500,N_3462,N_3400);
and U3501 (N_3501,N_3401,N_3495);
or U3502 (N_3502,N_3426,N_3487);
nor U3503 (N_3503,N_3453,N_3467);
or U3504 (N_3504,N_3406,N_3455);
nor U3505 (N_3505,N_3494,N_3496);
nand U3506 (N_3506,N_3418,N_3459);
nand U3507 (N_3507,N_3456,N_3424);
nand U3508 (N_3508,N_3436,N_3482);
or U3509 (N_3509,N_3438,N_3470);
or U3510 (N_3510,N_3485,N_3457);
nand U3511 (N_3511,N_3435,N_3488);
and U3512 (N_3512,N_3480,N_3466);
nor U3513 (N_3513,N_3425,N_3441);
and U3514 (N_3514,N_3458,N_3404);
nand U3515 (N_3515,N_3465,N_3443);
and U3516 (N_3516,N_3410,N_3440);
and U3517 (N_3517,N_3427,N_3432);
and U3518 (N_3518,N_3414,N_3422);
or U3519 (N_3519,N_3492,N_3445);
and U3520 (N_3520,N_3444,N_3433);
nor U3521 (N_3521,N_3449,N_3413);
or U3522 (N_3522,N_3423,N_3472);
nor U3523 (N_3523,N_3489,N_3497);
and U3524 (N_3524,N_3491,N_3408);
and U3525 (N_3525,N_3447,N_3471);
or U3526 (N_3526,N_3461,N_3419);
nor U3527 (N_3527,N_3499,N_3484);
and U3528 (N_3528,N_3469,N_3464);
and U3529 (N_3529,N_3452,N_3474);
nand U3530 (N_3530,N_3448,N_3402);
and U3531 (N_3531,N_3442,N_3428);
or U3532 (N_3532,N_3416,N_3475);
nand U3533 (N_3533,N_3477,N_3407);
nand U3534 (N_3534,N_3454,N_3498);
nand U3535 (N_3535,N_3409,N_3483);
or U3536 (N_3536,N_3468,N_3434);
or U3537 (N_3537,N_3493,N_3415);
and U3538 (N_3538,N_3463,N_3411);
and U3539 (N_3539,N_3460,N_3437);
or U3540 (N_3540,N_3490,N_3478);
and U3541 (N_3541,N_3420,N_3412);
nor U3542 (N_3542,N_3421,N_3446);
xnor U3543 (N_3543,N_3450,N_3439);
and U3544 (N_3544,N_3476,N_3429);
and U3545 (N_3545,N_3431,N_3481);
nand U3546 (N_3546,N_3403,N_3486);
or U3547 (N_3547,N_3473,N_3479);
or U3548 (N_3548,N_3405,N_3451);
or U3549 (N_3549,N_3417,N_3430);
nand U3550 (N_3550,N_3404,N_3444);
or U3551 (N_3551,N_3491,N_3493);
or U3552 (N_3552,N_3473,N_3461);
nor U3553 (N_3553,N_3431,N_3459);
and U3554 (N_3554,N_3492,N_3469);
and U3555 (N_3555,N_3434,N_3401);
nand U3556 (N_3556,N_3412,N_3441);
and U3557 (N_3557,N_3456,N_3482);
nor U3558 (N_3558,N_3472,N_3402);
or U3559 (N_3559,N_3420,N_3460);
or U3560 (N_3560,N_3471,N_3465);
and U3561 (N_3561,N_3478,N_3417);
or U3562 (N_3562,N_3499,N_3431);
and U3563 (N_3563,N_3475,N_3412);
nand U3564 (N_3564,N_3494,N_3416);
nor U3565 (N_3565,N_3498,N_3411);
nand U3566 (N_3566,N_3479,N_3491);
or U3567 (N_3567,N_3490,N_3484);
or U3568 (N_3568,N_3430,N_3456);
nor U3569 (N_3569,N_3481,N_3485);
nor U3570 (N_3570,N_3482,N_3400);
nor U3571 (N_3571,N_3482,N_3439);
and U3572 (N_3572,N_3403,N_3426);
nand U3573 (N_3573,N_3433,N_3472);
or U3574 (N_3574,N_3421,N_3418);
or U3575 (N_3575,N_3494,N_3400);
and U3576 (N_3576,N_3432,N_3405);
nor U3577 (N_3577,N_3460,N_3468);
nor U3578 (N_3578,N_3482,N_3466);
nor U3579 (N_3579,N_3421,N_3409);
nand U3580 (N_3580,N_3480,N_3438);
or U3581 (N_3581,N_3477,N_3408);
nor U3582 (N_3582,N_3459,N_3463);
nand U3583 (N_3583,N_3409,N_3478);
nor U3584 (N_3584,N_3411,N_3427);
nor U3585 (N_3585,N_3478,N_3444);
xnor U3586 (N_3586,N_3411,N_3404);
and U3587 (N_3587,N_3430,N_3438);
or U3588 (N_3588,N_3447,N_3402);
nor U3589 (N_3589,N_3426,N_3435);
and U3590 (N_3590,N_3412,N_3410);
nor U3591 (N_3591,N_3458,N_3475);
or U3592 (N_3592,N_3409,N_3497);
and U3593 (N_3593,N_3466,N_3492);
nor U3594 (N_3594,N_3494,N_3485);
and U3595 (N_3595,N_3444,N_3401);
nor U3596 (N_3596,N_3494,N_3454);
or U3597 (N_3597,N_3423,N_3494);
nor U3598 (N_3598,N_3445,N_3493);
xnor U3599 (N_3599,N_3475,N_3443);
or U3600 (N_3600,N_3522,N_3502);
nor U3601 (N_3601,N_3527,N_3551);
and U3602 (N_3602,N_3529,N_3544);
or U3603 (N_3603,N_3539,N_3516);
nand U3604 (N_3604,N_3543,N_3537);
or U3605 (N_3605,N_3535,N_3530);
nor U3606 (N_3606,N_3513,N_3542);
nor U3607 (N_3607,N_3588,N_3521);
nor U3608 (N_3608,N_3534,N_3509);
or U3609 (N_3609,N_3511,N_3520);
nor U3610 (N_3610,N_3510,N_3562);
and U3611 (N_3611,N_3582,N_3546);
nor U3612 (N_3612,N_3564,N_3512);
and U3613 (N_3613,N_3598,N_3575);
nand U3614 (N_3614,N_3532,N_3599);
nand U3615 (N_3615,N_3525,N_3540);
and U3616 (N_3616,N_3559,N_3504);
nor U3617 (N_3617,N_3515,N_3572);
and U3618 (N_3618,N_3508,N_3549);
xor U3619 (N_3619,N_3507,N_3585);
and U3620 (N_3620,N_3550,N_3500);
and U3621 (N_3621,N_3568,N_3579);
or U3622 (N_3622,N_3523,N_3556);
nand U3623 (N_3623,N_3574,N_3524);
and U3624 (N_3624,N_3591,N_3565);
nand U3625 (N_3625,N_3570,N_3514);
or U3626 (N_3626,N_3597,N_3578);
nand U3627 (N_3627,N_3531,N_3569);
or U3628 (N_3628,N_3553,N_3519);
or U3629 (N_3629,N_3506,N_3548);
and U3630 (N_3630,N_3595,N_3561);
or U3631 (N_3631,N_3566,N_3518);
nand U3632 (N_3632,N_3577,N_3528);
nor U3633 (N_3633,N_3580,N_3563);
or U3634 (N_3634,N_3576,N_3596);
nand U3635 (N_3635,N_3541,N_3587);
nand U3636 (N_3636,N_3586,N_3552);
or U3637 (N_3637,N_3560,N_3584);
or U3638 (N_3638,N_3538,N_3573);
or U3639 (N_3639,N_3547,N_3545);
or U3640 (N_3640,N_3536,N_3505);
and U3641 (N_3641,N_3526,N_3503);
nor U3642 (N_3642,N_3501,N_3594);
nand U3643 (N_3643,N_3581,N_3558);
nand U3644 (N_3644,N_3557,N_3555);
or U3645 (N_3645,N_3571,N_3593);
nor U3646 (N_3646,N_3592,N_3554);
or U3647 (N_3647,N_3590,N_3583);
nor U3648 (N_3648,N_3533,N_3567);
nor U3649 (N_3649,N_3517,N_3589);
or U3650 (N_3650,N_3550,N_3580);
nor U3651 (N_3651,N_3591,N_3511);
nand U3652 (N_3652,N_3529,N_3587);
and U3653 (N_3653,N_3555,N_3501);
nor U3654 (N_3654,N_3564,N_3516);
or U3655 (N_3655,N_3585,N_3532);
or U3656 (N_3656,N_3577,N_3515);
nand U3657 (N_3657,N_3521,N_3589);
nand U3658 (N_3658,N_3500,N_3511);
nand U3659 (N_3659,N_3511,N_3543);
nand U3660 (N_3660,N_3586,N_3525);
nand U3661 (N_3661,N_3572,N_3584);
xor U3662 (N_3662,N_3514,N_3504);
and U3663 (N_3663,N_3554,N_3577);
and U3664 (N_3664,N_3590,N_3540);
nand U3665 (N_3665,N_3505,N_3509);
or U3666 (N_3666,N_3558,N_3564);
xor U3667 (N_3667,N_3507,N_3529);
nand U3668 (N_3668,N_3528,N_3573);
and U3669 (N_3669,N_3593,N_3556);
or U3670 (N_3670,N_3526,N_3518);
or U3671 (N_3671,N_3538,N_3510);
nand U3672 (N_3672,N_3580,N_3549);
or U3673 (N_3673,N_3543,N_3598);
or U3674 (N_3674,N_3589,N_3558);
and U3675 (N_3675,N_3561,N_3588);
xnor U3676 (N_3676,N_3555,N_3534);
nor U3677 (N_3677,N_3561,N_3591);
nand U3678 (N_3678,N_3508,N_3598);
nor U3679 (N_3679,N_3533,N_3547);
nor U3680 (N_3680,N_3550,N_3564);
nor U3681 (N_3681,N_3555,N_3571);
and U3682 (N_3682,N_3573,N_3554);
nor U3683 (N_3683,N_3543,N_3589);
nand U3684 (N_3684,N_3572,N_3529);
and U3685 (N_3685,N_3563,N_3594);
nand U3686 (N_3686,N_3555,N_3524);
nor U3687 (N_3687,N_3562,N_3542);
nor U3688 (N_3688,N_3597,N_3550);
nor U3689 (N_3689,N_3594,N_3556);
and U3690 (N_3690,N_3583,N_3539);
and U3691 (N_3691,N_3581,N_3568);
xnor U3692 (N_3692,N_3550,N_3504);
and U3693 (N_3693,N_3555,N_3539);
and U3694 (N_3694,N_3594,N_3592);
or U3695 (N_3695,N_3542,N_3563);
nor U3696 (N_3696,N_3593,N_3572);
or U3697 (N_3697,N_3565,N_3535);
or U3698 (N_3698,N_3517,N_3572);
and U3699 (N_3699,N_3552,N_3550);
nor U3700 (N_3700,N_3649,N_3688);
nand U3701 (N_3701,N_3611,N_3686);
nor U3702 (N_3702,N_3621,N_3624);
or U3703 (N_3703,N_3664,N_3694);
nor U3704 (N_3704,N_3650,N_3627);
nand U3705 (N_3705,N_3677,N_3632);
or U3706 (N_3706,N_3681,N_3631);
or U3707 (N_3707,N_3600,N_3647);
nor U3708 (N_3708,N_3616,N_3655);
nand U3709 (N_3709,N_3634,N_3608);
or U3710 (N_3710,N_3668,N_3653);
nand U3711 (N_3711,N_3648,N_3629);
or U3712 (N_3712,N_3657,N_3699);
nand U3713 (N_3713,N_3614,N_3618);
nor U3714 (N_3714,N_3656,N_3619);
or U3715 (N_3715,N_3654,N_3607);
nor U3716 (N_3716,N_3671,N_3644);
or U3717 (N_3717,N_3630,N_3620);
or U3718 (N_3718,N_3626,N_3689);
or U3719 (N_3719,N_3662,N_3663);
nand U3720 (N_3720,N_3685,N_3610);
nand U3721 (N_3721,N_3674,N_3625);
nand U3722 (N_3722,N_3683,N_3605);
nand U3723 (N_3723,N_3636,N_3609);
or U3724 (N_3724,N_3682,N_3646);
and U3725 (N_3725,N_3680,N_3697);
nor U3726 (N_3726,N_3604,N_3666);
nand U3727 (N_3727,N_3676,N_3638);
nand U3728 (N_3728,N_3679,N_3642);
nand U3729 (N_3729,N_3633,N_3659);
and U3730 (N_3730,N_3622,N_3643);
nor U3731 (N_3731,N_3603,N_3667);
or U3732 (N_3732,N_3640,N_3635);
and U3733 (N_3733,N_3661,N_3612);
nand U3734 (N_3734,N_3693,N_3698);
nand U3735 (N_3735,N_3628,N_3606);
nor U3736 (N_3736,N_3670,N_3623);
nor U3737 (N_3737,N_3641,N_3669);
nor U3738 (N_3738,N_3684,N_3637);
nand U3739 (N_3739,N_3692,N_3675);
nand U3740 (N_3740,N_3645,N_3652);
nand U3741 (N_3741,N_3678,N_3617);
nand U3742 (N_3742,N_3673,N_3601);
xor U3743 (N_3743,N_3651,N_3665);
nand U3744 (N_3744,N_3615,N_3639);
nand U3745 (N_3745,N_3696,N_3691);
and U3746 (N_3746,N_3690,N_3613);
or U3747 (N_3747,N_3687,N_3672);
xnor U3748 (N_3748,N_3695,N_3602);
or U3749 (N_3749,N_3658,N_3660);
nor U3750 (N_3750,N_3660,N_3688);
nor U3751 (N_3751,N_3636,N_3629);
nand U3752 (N_3752,N_3640,N_3681);
nor U3753 (N_3753,N_3659,N_3634);
or U3754 (N_3754,N_3626,N_3647);
nor U3755 (N_3755,N_3665,N_3691);
and U3756 (N_3756,N_3692,N_3618);
or U3757 (N_3757,N_3667,N_3623);
nor U3758 (N_3758,N_3639,N_3646);
nand U3759 (N_3759,N_3607,N_3611);
or U3760 (N_3760,N_3658,N_3616);
nand U3761 (N_3761,N_3635,N_3621);
nor U3762 (N_3762,N_3638,N_3682);
nor U3763 (N_3763,N_3642,N_3673);
nand U3764 (N_3764,N_3690,N_3682);
nor U3765 (N_3765,N_3636,N_3664);
and U3766 (N_3766,N_3640,N_3628);
and U3767 (N_3767,N_3607,N_3676);
and U3768 (N_3768,N_3644,N_3660);
or U3769 (N_3769,N_3667,N_3650);
or U3770 (N_3770,N_3606,N_3645);
nand U3771 (N_3771,N_3687,N_3660);
nor U3772 (N_3772,N_3675,N_3621);
or U3773 (N_3773,N_3614,N_3666);
nor U3774 (N_3774,N_3689,N_3642);
nand U3775 (N_3775,N_3617,N_3603);
nand U3776 (N_3776,N_3635,N_3617);
nor U3777 (N_3777,N_3667,N_3656);
xor U3778 (N_3778,N_3615,N_3631);
nor U3779 (N_3779,N_3601,N_3638);
or U3780 (N_3780,N_3621,N_3609);
nor U3781 (N_3781,N_3619,N_3686);
nor U3782 (N_3782,N_3697,N_3628);
xnor U3783 (N_3783,N_3657,N_3672);
nor U3784 (N_3784,N_3638,N_3661);
and U3785 (N_3785,N_3675,N_3648);
nand U3786 (N_3786,N_3678,N_3614);
and U3787 (N_3787,N_3690,N_3610);
nand U3788 (N_3788,N_3665,N_3695);
nand U3789 (N_3789,N_3698,N_3616);
and U3790 (N_3790,N_3612,N_3692);
nor U3791 (N_3791,N_3680,N_3695);
and U3792 (N_3792,N_3692,N_3670);
or U3793 (N_3793,N_3647,N_3653);
nor U3794 (N_3794,N_3685,N_3605);
nor U3795 (N_3795,N_3697,N_3635);
or U3796 (N_3796,N_3673,N_3643);
nor U3797 (N_3797,N_3625,N_3633);
and U3798 (N_3798,N_3632,N_3611);
nand U3799 (N_3799,N_3695,N_3687);
nor U3800 (N_3800,N_3777,N_3708);
or U3801 (N_3801,N_3796,N_3779);
nand U3802 (N_3802,N_3714,N_3743);
and U3803 (N_3803,N_3719,N_3718);
nor U3804 (N_3804,N_3786,N_3781);
nand U3805 (N_3805,N_3725,N_3703);
or U3806 (N_3806,N_3755,N_3776);
nor U3807 (N_3807,N_3732,N_3712);
nor U3808 (N_3808,N_3783,N_3764);
xnor U3809 (N_3809,N_3701,N_3726);
and U3810 (N_3810,N_3727,N_3731);
nand U3811 (N_3811,N_3713,N_3790);
and U3812 (N_3812,N_3736,N_3757);
nand U3813 (N_3813,N_3756,N_3758);
nor U3814 (N_3814,N_3761,N_3792);
nor U3815 (N_3815,N_3789,N_3702);
or U3816 (N_3816,N_3770,N_3782);
or U3817 (N_3817,N_3794,N_3728);
nor U3818 (N_3818,N_3722,N_3745);
and U3819 (N_3819,N_3720,N_3753);
nand U3820 (N_3820,N_3739,N_3797);
or U3821 (N_3821,N_3798,N_3734);
or U3822 (N_3822,N_3738,N_3766);
nand U3823 (N_3823,N_3706,N_3747);
nand U3824 (N_3824,N_3780,N_3784);
nor U3825 (N_3825,N_3754,N_3768);
or U3826 (N_3826,N_3704,N_3787);
or U3827 (N_3827,N_3716,N_3778);
nand U3828 (N_3828,N_3715,N_3700);
and U3829 (N_3829,N_3709,N_3733);
and U3830 (N_3830,N_3775,N_3744);
nor U3831 (N_3831,N_3760,N_3741);
and U3832 (N_3832,N_3710,N_3749);
xnor U3833 (N_3833,N_3750,N_3767);
nor U3834 (N_3834,N_3724,N_3785);
and U3835 (N_3835,N_3763,N_3795);
nand U3836 (N_3836,N_3751,N_3746);
nor U3837 (N_3837,N_3774,N_3721);
and U3838 (N_3838,N_3788,N_3772);
and U3839 (N_3839,N_3707,N_3771);
nor U3840 (N_3840,N_3742,N_3729);
and U3841 (N_3841,N_3765,N_3793);
nor U3842 (N_3842,N_3735,N_3752);
nor U3843 (N_3843,N_3717,N_3723);
and U3844 (N_3844,N_3705,N_3748);
nor U3845 (N_3845,N_3740,N_3799);
nand U3846 (N_3846,N_3773,N_3762);
nand U3847 (N_3847,N_3711,N_3730);
and U3848 (N_3848,N_3737,N_3791);
xnor U3849 (N_3849,N_3769,N_3759);
and U3850 (N_3850,N_3747,N_3796);
nand U3851 (N_3851,N_3798,N_3703);
and U3852 (N_3852,N_3719,N_3768);
nor U3853 (N_3853,N_3762,N_3746);
nor U3854 (N_3854,N_3774,N_3731);
or U3855 (N_3855,N_3718,N_3775);
and U3856 (N_3856,N_3775,N_3726);
and U3857 (N_3857,N_3717,N_3714);
nand U3858 (N_3858,N_3703,N_3759);
nor U3859 (N_3859,N_3710,N_3712);
nand U3860 (N_3860,N_3797,N_3785);
nor U3861 (N_3861,N_3746,N_3720);
nand U3862 (N_3862,N_3729,N_3716);
nor U3863 (N_3863,N_3738,N_3716);
or U3864 (N_3864,N_3725,N_3719);
or U3865 (N_3865,N_3765,N_3713);
nor U3866 (N_3866,N_3741,N_3702);
and U3867 (N_3867,N_3756,N_3731);
nor U3868 (N_3868,N_3753,N_3793);
nor U3869 (N_3869,N_3779,N_3701);
nor U3870 (N_3870,N_3798,N_3740);
and U3871 (N_3871,N_3718,N_3751);
or U3872 (N_3872,N_3717,N_3796);
nand U3873 (N_3873,N_3768,N_3758);
nand U3874 (N_3874,N_3759,N_3734);
nor U3875 (N_3875,N_3772,N_3751);
and U3876 (N_3876,N_3713,N_3700);
or U3877 (N_3877,N_3782,N_3745);
nor U3878 (N_3878,N_3758,N_3710);
nand U3879 (N_3879,N_3747,N_3700);
nand U3880 (N_3880,N_3762,N_3747);
or U3881 (N_3881,N_3738,N_3715);
nand U3882 (N_3882,N_3725,N_3780);
or U3883 (N_3883,N_3742,N_3796);
or U3884 (N_3884,N_3727,N_3779);
and U3885 (N_3885,N_3750,N_3759);
and U3886 (N_3886,N_3702,N_3761);
nand U3887 (N_3887,N_3786,N_3727);
or U3888 (N_3888,N_3792,N_3770);
nor U3889 (N_3889,N_3757,N_3786);
nor U3890 (N_3890,N_3713,N_3792);
nor U3891 (N_3891,N_3703,N_3785);
nand U3892 (N_3892,N_3701,N_3796);
nor U3893 (N_3893,N_3718,N_3756);
nand U3894 (N_3894,N_3737,N_3758);
nor U3895 (N_3895,N_3703,N_3714);
nand U3896 (N_3896,N_3737,N_3792);
and U3897 (N_3897,N_3785,N_3773);
nand U3898 (N_3898,N_3791,N_3725);
or U3899 (N_3899,N_3738,N_3763);
and U3900 (N_3900,N_3843,N_3888);
or U3901 (N_3901,N_3846,N_3803);
nand U3902 (N_3902,N_3856,N_3870);
nand U3903 (N_3903,N_3897,N_3894);
or U3904 (N_3904,N_3898,N_3836);
nor U3905 (N_3905,N_3805,N_3848);
and U3906 (N_3906,N_3840,N_3862);
and U3907 (N_3907,N_3877,N_3899);
and U3908 (N_3908,N_3818,N_3872);
or U3909 (N_3909,N_3832,N_3845);
or U3910 (N_3910,N_3821,N_3892);
or U3911 (N_3911,N_3875,N_3831);
nand U3912 (N_3912,N_3824,N_3827);
nor U3913 (N_3913,N_3809,N_3811);
and U3914 (N_3914,N_3857,N_3859);
nor U3915 (N_3915,N_3825,N_3810);
and U3916 (N_3916,N_3860,N_3826);
and U3917 (N_3917,N_3851,N_3867);
nand U3918 (N_3918,N_3889,N_3853);
nand U3919 (N_3919,N_3801,N_3822);
or U3920 (N_3920,N_3883,N_3880);
or U3921 (N_3921,N_3855,N_3838);
and U3922 (N_3922,N_3861,N_3885);
or U3923 (N_3923,N_3871,N_3893);
nor U3924 (N_3924,N_3814,N_3887);
or U3925 (N_3925,N_3830,N_3879);
or U3926 (N_3926,N_3828,N_3852);
nand U3927 (N_3927,N_3817,N_3800);
and U3928 (N_3928,N_3854,N_3841);
nand U3929 (N_3929,N_3882,N_3886);
and U3930 (N_3930,N_3802,N_3858);
or U3931 (N_3931,N_3823,N_3808);
or U3932 (N_3932,N_3847,N_3865);
nand U3933 (N_3933,N_3806,N_3874);
and U3934 (N_3934,N_3833,N_3884);
nand U3935 (N_3935,N_3895,N_3812);
nor U3936 (N_3936,N_3813,N_3829);
nor U3937 (N_3937,N_3876,N_3839);
or U3938 (N_3938,N_3834,N_3820);
or U3939 (N_3939,N_3842,N_3873);
and U3940 (N_3940,N_3837,N_3844);
and U3941 (N_3941,N_3890,N_3816);
nor U3942 (N_3942,N_3881,N_3896);
and U3943 (N_3943,N_3835,N_3850);
or U3944 (N_3944,N_3807,N_3863);
nand U3945 (N_3945,N_3819,N_3815);
nand U3946 (N_3946,N_3891,N_3869);
and U3947 (N_3947,N_3804,N_3864);
and U3948 (N_3948,N_3868,N_3878);
and U3949 (N_3949,N_3849,N_3866);
or U3950 (N_3950,N_3865,N_3802);
or U3951 (N_3951,N_3827,N_3883);
nand U3952 (N_3952,N_3861,N_3849);
nor U3953 (N_3953,N_3834,N_3873);
nor U3954 (N_3954,N_3838,N_3889);
nor U3955 (N_3955,N_3872,N_3841);
and U3956 (N_3956,N_3852,N_3804);
and U3957 (N_3957,N_3887,N_3891);
or U3958 (N_3958,N_3811,N_3857);
or U3959 (N_3959,N_3848,N_3890);
nand U3960 (N_3960,N_3882,N_3878);
or U3961 (N_3961,N_3881,N_3851);
or U3962 (N_3962,N_3833,N_3837);
nand U3963 (N_3963,N_3878,N_3814);
nor U3964 (N_3964,N_3897,N_3814);
nor U3965 (N_3965,N_3806,N_3869);
nor U3966 (N_3966,N_3884,N_3882);
and U3967 (N_3967,N_3899,N_3893);
and U3968 (N_3968,N_3830,N_3837);
and U3969 (N_3969,N_3837,N_3850);
nor U3970 (N_3970,N_3807,N_3853);
and U3971 (N_3971,N_3870,N_3875);
nand U3972 (N_3972,N_3833,N_3835);
nand U3973 (N_3973,N_3826,N_3827);
nor U3974 (N_3974,N_3887,N_3892);
nor U3975 (N_3975,N_3863,N_3826);
and U3976 (N_3976,N_3877,N_3863);
or U3977 (N_3977,N_3853,N_3876);
or U3978 (N_3978,N_3807,N_3882);
nand U3979 (N_3979,N_3843,N_3851);
and U3980 (N_3980,N_3841,N_3857);
or U3981 (N_3981,N_3885,N_3806);
or U3982 (N_3982,N_3891,N_3896);
nor U3983 (N_3983,N_3822,N_3898);
nor U3984 (N_3984,N_3867,N_3872);
nor U3985 (N_3985,N_3896,N_3860);
nor U3986 (N_3986,N_3825,N_3846);
or U3987 (N_3987,N_3839,N_3898);
nand U3988 (N_3988,N_3877,N_3888);
or U3989 (N_3989,N_3826,N_3856);
and U3990 (N_3990,N_3802,N_3809);
or U3991 (N_3991,N_3807,N_3892);
nand U3992 (N_3992,N_3884,N_3810);
nand U3993 (N_3993,N_3813,N_3827);
or U3994 (N_3994,N_3869,N_3811);
nor U3995 (N_3995,N_3850,N_3878);
nor U3996 (N_3996,N_3863,N_3893);
nand U3997 (N_3997,N_3816,N_3811);
nor U3998 (N_3998,N_3821,N_3849);
nor U3999 (N_3999,N_3886,N_3810);
or U4000 (N_4000,N_3940,N_3924);
and U4001 (N_4001,N_3947,N_3960);
or U4002 (N_4002,N_3957,N_3949);
nand U4003 (N_4003,N_3967,N_3988);
and U4004 (N_4004,N_3900,N_3979);
nor U4005 (N_4005,N_3998,N_3970);
and U4006 (N_4006,N_3905,N_3980);
and U4007 (N_4007,N_3938,N_3995);
nor U4008 (N_4008,N_3955,N_3937);
nand U4009 (N_4009,N_3943,N_3952);
nor U4010 (N_4010,N_3935,N_3939);
nor U4011 (N_4011,N_3904,N_3977);
nand U4012 (N_4012,N_3933,N_3963);
nand U4013 (N_4013,N_3912,N_3965);
or U4014 (N_4014,N_3915,N_3999);
nor U4015 (N_4015,N_3956,N_3907);
nor U4016 (N_4016,N_3920,N_3908);
nor U4017 (N_4017,N_3927,N_3916);
xor U4018 (N_4018,N_3981,N_3931);
xor U4019 (N_4019,N_3930,N_3992);
or U4020 (N_4020,N_3928,N_3986);
and U4021 (N_4021,N_3975,N_3922);
nand U4022 (N_4022,N_3913,N_3954);
and U4023 (N_4023,N_3994,N_3991);
or U4024 (N_4024,N_3990,N_3923);
nor U4025 (N_4025,N_3950,N_3984);
and U4026 (N_4026,N_3921,N_3932);
and U4027 (N_4027,N_3958,N_3969);
nand U4028 (N_4028,N_3919,N_3972);
or U4029 (N_4029,N_3968,N_3944);
xnor U4030 (N_4030,N_3945,N_3906);
nor U4031 (N_4031,N_3903,N_3971);
xor U4032 (N_4032,N_3982,N_3964);
and U4033 (N_4033,N_3918,N_3936);
or U4034 (N_4034,N_3902,N_3911);
and U4035 (N_4035,N_3978,N_3951);
nand U4036 (N_4036,N_3925,N_3909);
and U4037 (N_4037,N_3948,N_3996);
nand U4038 (N_4038,N_3985,N_3910);
and U4039 (N_4039,N_3973,N_3993);
nand U4040 (N_4040,N_3974,N_3987);
or U4041 (N_4041,N_3926,N_3953);
and U4042 (N_4042,N_3942,N_3959);
xnor U4043 (N_4043,N_3962,N_3929);
nand U4044 (N_4044,N_3989,N_3914);
nor U4045 (N_4045,N_3934,N_3976);
or U4046 (N_4046,N_3917,N_3946);
nor U4047 (N_4047,N_3997,N_3966);
and U4048 (N_4048,N_3901,N_3983);
and U4049 (N_4049,N_3941,N_3961);
nand U4050 (N_4050,N_3944,N_3900);
or U4051 (N_4051,N_3982,N_3903);
nand U4052 (N_4052,N_3927,N_3914);
or U4053 (N_4053,N_3988,N_3923);
xnor U4054 (N_4054,N_3901,N_3963);
nand U4055 (N_4055,N_3936,N_3955);
and U4056 (N_4056,N_3992,N_3973);
nor U4057 (N_4057,N_3920,N_3930);
nand U4058 (N_4058,N_3924,N_3999);
nand U4059 (N_4059,N_3932,N_3998);
xor U4060 (N_4060,N_3930,N_3952);
nand U4061 (N_4061,N_3920,N_3951);
and U4062 (N_4062,N_3995,N_3924);
nor U4063 (N_4063,N_3916,N_3931);
and U4064 (N_4064,N_3974,N_3970);
or U4065 (N_4065,N_3980,N_3902);
or U4066 (N_4066,N_3976,N_3906);
and U4067 (N_4067,N_3942,N_3988);
or U4068 (N_4068,N_3929,N_3936);
or U4069 (N_4069,N_3973,N_3978);
nor U4070 (N_4070,N_3912,N_3944);
nand U4071 (N_4071,N_3958,N_3973);
or U4072 (N_4072,N_3953,N_3973);
or U4073 (N_4073,N_3955,N_3967);
or U4074 (N_4074,N_3962,N_3970);
nand U4075 (N_4075,N_3922,N_3962);
or U4076 (N_4076,N_3922,N_3963);
xnor U4077 (N_4077,N_3958,N_3960);
nor U4078 (N_4078,N_3904,N_3932);
nor U4079 (N_4079,N_3913,N_3970);
nand U4080 (N_4080,N_3918,N_3960);
or U4081 (N_4081,N_3962,N_3984);
xor U4082 (N_4082,N_3906,N_3978);
and U4083 (N_4083,N_3926,N_3990);
or U4084 (N_4084,N_3922,N_3995);
or U4085 (N_4085,N_3974,N_3998);
and U4086 (N_4086,N_3907,N_3972);
or U4087 (N_4087,N_3938,N_3956);
and U4088 (N_4088,N_3932,N_3961);
and U4089 (N_4089,N_3974,N_3902);
nor U4090 (N_4090,N_3933,N_3992);
nand U4091 (N_4091,N_3940,N_3958);
or U4092 (N_4092,N_3970,N_3983);
nor U4093 (N_4093,N_3905,N_3923);
nand U4094 (N_4094,N_3935,N_3931);
and U4095 (N_4095,N_3948,N_3968);
nand U4096 (N_4096,N_3952,N_3971);
nand U4097 (N_4097,N_3993,N_3943);
or U4098 (N_4098,N_3993,N_3952);
and U4099 (N_4099,N_3940,N_3907);
nand U4100 (N_4100,N_4087,N_4064);
or U4101 (N_4101,N_4054,N_4060);
and U4102 (N_4102,N_4091,N_4076);
and U4103 (N_4103,N_4021,N_4056);
nand U4104 (N_4104,N_4048,N_4012);
nand U4105 (N_4105,N_4031,N_4079);
and U4106 (N_4106,N_4094,N_4029);
nand U4107 (N_4107,N_4083,N_4022);
nand U4108 (N_4108,N_4096,N_4003);
nand U4109 (N_4109,N_4045,N_4080);
nand U4110 (N_4110,N_4024,N_4061);
nand U4111 (N_4111,N_4069,N_4092);
nand U4112 (N_4112,N_4075,N_4038);
nand U4113 (N_4113,N_4010,N_4074);
or U4114 (N_4114,N_4051,N_4077);
nand U4115 (N_4115,N_4039,N_4082);
nand U4116 (N_4116,N_4006,N_4009);
and U4117 (N_4117,N_4063,N_4071);
xor U4118 (N_4118,N_4018,N_4088);
or U4119 (N_4119,N_4053,N_4043);
nand U4120 (N_4120,N_4042,N_4023);
nor U4121 (N_4121,N_4044,N_4057);
nor U4122 (N_4122,N_4017,N_4027);
nand U4123 (N_4123,N_4005,N_4028);
and U4124 (N_4124,N_4065,N_4025);
and U4125 (N_4125,N_4049,N_4046);
or U4126 (N_4126,N_4007,N_4059);
and U4127 (N_4127,N_4072,N_4020);
and U4128 (N_4128,N_4099,N_4078);
and U4129 (N_4129,N_4073,N_4095);
nor U4130 (N_4130,N_4026,N_4052);
or U4131 (N_4131,N_4058,N_4086);
nand U4132 (N_4132,N_4013,N_4019);
nor U4133 (N_4133,N_4090,N_4008);
nand U4134 (N_4134,N_4011,N_4089);
or U4135 (N_4135,N_4085,N_4037);
or U4136 (N_4136,N_4098,N_4016);
and U4137 (N_4137,N_4035,N_4066);
nor U4138 (N_4138,N_4014,N_4067);
nand U4139 (N_4139,N_4030,N_4097);
or U4140 (N_4140,N_4015,N_4001);
or U4141 (N_4141,N_4068,N_4000);
nand U4142 (N_4142,N_4050,N_4047);
nand U4143 (N_4143,N_4081,N_4034);
and U4144 (N_4144,N_4004,N_4041);
or U4145 (N_4145,N_4002,N_4070);
nand U4146 (N_4146,N_4062,N_4084);
nand U4147 (N_4147,N_4040,N_4036);
or U4148 (N_4148,N_4032,N_4093);
nand U4149 (N_4149,N_4033,N_4055);
or U4150 (N_4150,N_4043,N_4049);
nand U4151 (N_4151,N_4036,N_4092);
and U4152 (N_4152,N_4087,N_4093);
nand U4153 (N_4153,N_4056,N_4001);
and U4154 (N_4154,N_4011,N_4008);
nand U4155 (N_4155,N_4044,N_4043);
nand U4156 (N_4156,N_4061,N_4060);
nand U4157 (N_4157,N_4059,N_4027);
nand U4158 (N_4158,N_4021,N_4075);
or U4159 (N_4159,N_4093,N_4027);
or U4160 (N_4160,N_4047,N_4024);
or U4161 (N_4161,N_4082,N_4074);
and U4162 (N_4162,N_4007,N_4075);
nand U4163 (N_4163,N_4023,N_4086);
or U4164 (N_4164,N_4029,N_4079);
nor U4165 (N_4165,N_4090,N_4024);
nor U4166 (N_4166,N_4074,N_4048);
nand U4167 (N_4167,N_4013,N_4078);
nor U4168 (N_4168,N_4032,N_4017);
nor U4169 (N_4169,N_4088,N_4012);
or U4170 (N_4170,N_4023,N_4055);
or U4171 (N_4171,N_4086,N_4048);
and U4172 (N_4172,N_4010,N_4020);
nor U4173 (N_4173,N_4026,N_4083);
nand U4174 (N_4174,N_4046,N_4084);
or U4175 (N_4175,N_4083,N_4077);
nor U4176 (N_4176,N_4048,N_4070);
nor U4177 (N_4177,N_4059,N_4077);
nor U4178 (N_4178,N_4085,N_4007);
nand U4179 (N_4179,N_4035,N_4098);
xor U4180 (N_4180,N_4045,N_4037);
and U4181 (N_4181,N_4040,N_4084);
and U4182 (N_4182,N_4054,N_4036);
and U4183 (N_4183,N_4031,N_4043);
xnor U4184 (N_4184,N_4056,N_4003);
nand U4185 (N_4185,N_4099,N_4067);
nor U4186 (N_4186,N_4065,N_4099);
or U4187 (N_4187,N_4020,N_4027);
and U4188 (N_4188,N_4004,N_4074);
nor U4189 (N_4189,N_4036,N_4027);
nor U4190 (N_4190,N_4083,N_4008);
nand U4191 (N_4191,N_4063,N_4053);
and U4192 (N_4192,N_4059,N_4011);
or U4193 (N_4193,N_4019,N_4051);
nand U4194 (N_4194,N_4076,N_4079);
and U4195 (N_4195,N_4043,N_4011);
and U4196 (N_4196,N_4016,N_4013);
or U4197 (N_4197,N_4045,N_4016);
or U4198 (N_4198,N_4071,N_4003);
and U4199 (N_4199,N_4063,N_4078);
nor U4200 (N_4200,N_4186,N_4164);
and U4201 (N_4201,N_4194,N_4197);
or U4202 (N_4202,N_4154,N_4160);
nor U4203 (N_4203,N_4180,N_4159);
or U4204 (N_4204,N_4175,N_4177);
or U4205 (N_4205,N_4131,N_4130);
and U4206 (N_4206,N_4150,N_4184);
nand U4207 (N_4207,N_4185,N_4101);
and U4208 (N_4208,N_4127,N_4148);
nor U4209 (N_4209,N_4134,N_4119);
and U4210 (N_4210,N_4142,N_4157);
nand U4211 (N_4211,N_4189,N_4178);
nor U4212 (N_4212,N_4141,N_4163);
nor U4213 (N_4213,N_4155,N_4158);
and U4214 (N_4214,N_4162,N_4107);
xnor U4215 (N_4215,N_4199,N_4170);
and U4216 (N_4216,N_4121,N_4128);
nor U4217 (N_4217,N_4195,N_4171);
or U4218 (N_4218,N_4151,N_4123);
nand U4219 (N_4219,N_4135,N_4129);
nand U4220 (N_4220,N_4117,N_4105);
nor U4221 (N_4221,N_4112,N_4114);
nor U4222 (N_4222,N_4169,N_4147);
and U4223 (N_4223,N_4136,N_4110);
or U4224 (N_4224,N_4143,N_4152);
or U4225 (N_4225,N_4104,N_4118);
nand U4226 (N_4226,N_4133,N_4198);
nor U4227 (N_4227,N_4179,N_4176);
nand U4228 (N_4228,N_4144,N_4183);
nor U4229 (N_4229,N_4174,N_4196);
and U4230 (N_4230,N_4122,N_4165);
nor U4231 (N_4231,N_4115,N_4102);
nand U4232 (N_4232,N_4193,N_4173);
or U4233 (N_4233,N_4103,N_4153);
nand U4234 (N_4234,N_4100,N_4113);
nand U4235 (N_4235,N_4181,N_4172);
or U4236 (N_4236,N_4188,N_4139);
nor U4237 (N_4237,N_4108,N_4167);
or U4238 (N_4238,N_4125,N_4161);
or U4239 (N_4239,N_4182,N_4190);
nor U4240 (N_4240,N_4138,N_4192);
or U4241 (N_4241,N_4106,N_4149);
and U4242 (N_4242,N_4132,N_4168);
nand U4243 (N_4243,N_4111,N_4109);
nand U4244 (N_4244,N_4191,N_4137);
nand U4245 (N_4245,N_4116,N_4166);
nand U4246 (N_4246,N_4146,N_4140);
nor U4247 (N_4247,N_4124,N_4187);
and U4248 (N_4248,N_4120,N_4126);
and U4249 (N_4249,N_4156,N_4145);
nor U4250 (N_4250,N_4121,N_4155);
nor U4251 (N_4251,N_4145,N_4147);
or U4252 (N_4252,N_4133,N_4129);
nor U4253 (N_4253,N_4140,N_4199);
nor U4254 (N_4254,N_4152,N_4175);
or U4255 (N_4255,N_4199,N_4196);
and U4256 (N_4256,N_4181,N_4110);
or U4257 (N_4257,N_4132,N_4120);
nand U4258 (N_4258,N_4160,N_4119);
or U4259 (N_4259,N_4135,N_4177);
or U4260 (N_4260,N_4125,N_4151);
nand U4261 (N_4261,N_4119,N_4155);
and U4262 (N_4262,N_4103,N_4176);
nor U4263 (N_4263,N_4108,N_4143);
nand U4264 (N_4264,N_4140,N_4125);
or U4265 (N_4265,N_4125,N_4198);
nor U4266 (N_4266,N_4182,N_4157);
or U4267 (N_4267,N_4154,N_4118);
nor U4268 (N_4268,N_4114,N_4180);
or U4269 (N_4269,N_4143,N_4165);
nor U4270 (N_4270,N_4186,N_4166);
nand U4271 (N_4271,N_4182,N_4193);
nand U4272 (N_4272,N_4171,N_4118);
and U4273 (N_4273,N_4196,N_4150);
and U4274 (N_4274,N_4104,N_4140);
or U4275 (N_4275,N_4119,N_4157);
xor U4276 (N_4276,N_4147,N_4162);
or U4277 (N_4277,N_4115,N_4171);
nand U4278 (N_4278,N_4142,N_4183);
and U4279 (N_4279,N_4103,N_4186);
and U4280 (N_4280,N_4160,N_4150);
nor U4281 (N_4281,N_4122,N_4153);
nand U4282 (N_4282,N_4189,N_4155);
or U4283 (N_4283,N_4191,N_4173);
nor U4284 (N_4284,N_4108,N_4141);
nor U4285 (N_4285,N_4115,N_4195);
nand U4286 (N_4286,N_4103,N_4141);
nand U4287 (N_4287,N_4196,N_4149);
or U4288 (N_4288,N_4175,N_4187);
or U4289 (N_4289,N_4193,N_4162);
xor U4290 (N_4290,N_4181,N_4142);
or U4291 (N_4291,N_4121,N_4171);
nor U4292 (N_4292,N_4132,N_4194);
nand U4293 (N_4293,N_4146,N_4139);
nand U4294 (N_4294,N_4162,N_4135);
nor U4295 (N_4295,N_4156,N_4113);
nand U4296 (N_4296,N_4155,N_4135);
and U4297 (N_4297,N_4130,N_4141);
nor U4298 (N_4298,N_4101,N_4163);
and U4299 (N_4299,N_4109,N_4100);
nor U4300 (N_4300,N_4216,N_4265);
or U4301 (N_4301,N_4273,N_4224);
nand U4302 (N_4302,N_4221,N_4238);
nand U4303 (N_4303,N_4222,N_4268);
nand U4304 (N_4304,N_4240,N_4245);
and U4305 (N_4305,N_4218,N_4211);
and U4306 (N_4306,N_4247,N_4251);
and U4307 (N_4307,N_4242,N_4208);
and U4308 (N_4308,N_4264,N_4283);
or U4309 (N_4309,N_4250,N_4241);
and U4310 (N_4310,N_4263,N_4269);
or U4311 (N_4311,N_4215,N_4243);
nor U4312 (N_4312,N_4223,N_4259);
nor U4313 (N_4313,N_4228,N_4295);
and U4314 (N_4314,N_4257,N_4276);
and U4315 (N_4315,N_4260,N_4262);
and U4316 (N_4316,N_4284,N_4212);
or U4317 (N_4317,N_4226,N_4261);
nor U4318 (N_4318,N_4214,N_4217);
and U4319 (N_4319,N_4274,N_4237);
or U4320 (N_4320,N_4294,N_4275);
nor U4321 (N_4321,N_4246,N_4239);
xor U4322 (N_4322,N_4236,N_4231);
or U4323 (N_4323,N_4256,N_4286);
nand U4324 (N_4324,N_4219,N_4285);
nor U4325 (N_4325,N_4298,N_4277);
or U4326 (N_4326,N_4203,N_4287);
or U4327 (N_4327,N_4249,N_4230);
nand U4328 (N_4328,N_4204,N_4200);
nand U4329 (N_4329,N_4232,N_4291);
and U4330 (N_4330,N_4205,N_4278);
and U4331 (N_4331,N_4254,N_4299);
and U4332 (N_4332,N_4292,N_4225);
or U4333 (N_4333,N_4227,N_4206);
nor U4334 (N_4334,N_4244,N_4288);
nand U4335 (N_4335,N_4220,N_4235);
nor U4336 (N_4336,N_4280,N_4281);
nand U4337 (N_4337,N_4296,N_4229);
and U4338 (N_4338,N_4248,N_4279);
or U4339 (N_4339,N_4267,N_4253);
nor U4340 (N_4340,N_4255,N_4207);
and U4341 (N_4341,N_4272,N_4266);
and U4342 (N_4342,N_4210,N_4271);
nand U4343 (N_4343,N_4282,N_4201);
nor U4344 (N_4344,N_4252,N_4202);
or U4345 (N_4345,N_4270,N_4234);
nor U4346 (N_4346,N_4209,N_4293);
and U4347 (N_4347,N_4258,N_4233);
nor U4348 (N_4348,N_4289,N_4297);
or U4349 (N_4349,N_4290,N_4213);
or U4350 (N_4350,N_4251,N_4227);
and U4351 (N_4351,N_4276,N_4232);
or U4352 (N_4352,N_4285,N_4223);
nand U4353 (N_4353,N_4211,N_4283);
or U4354 (N_4354,N_4290,N_4211);
nor U4355 (N_4355,N_4240,N_4200);
and U4356 (N_4356,N_4298,N_4217);
or U4357 (N_4357,N_4295,N_4252);
or U4358 (N_4358,N_4256,N_4267);
nor U4359 (N_4359,N_4288,N_4238);
or U4360 (N_4360,N_4288,N_4237);
or U4361 (N_4361,N_4298,N_4276);
nand U4362 (N_4362,N_4201,N_4215);
nand U4363 (N_4363,N_4264,N_4208);
or U4364 (N_4364,N_4263,N_4202);
and U4365 (N_4365,N_4281,N_4217);
and U4366 (N_4366,N_4275,N_4211);
nor U4367 (N_4367,N_4271,N_4242);
nand U4368 (N_4368,N_4205,N_4287);
xnor U4369 (N_4369,N_4263,N_4226);
nand U4370 (N_4370,N_4291,N_4225);
nor U4371 (N_4371,N_4283,N_4282);
nor U4372 (N_4372,N_4262,N_4280);
nor U4373 (N_4373,N_4222,N_4227);
and U4374 (N_4374,N_4246,N_4271);
nor U4375 (N_4375,N_4291,N_4202);
xor U4376 (N_4376,N_4248,N_4221);
nor U4377 (N_4377,N_4272,N_4214);
and U4378 (N_4378,N_4283,N_4213);
nand U4379 (N_4379,N_4282,N_4263);
and U4380 (N_4380,N_4236,N_4225);
and U4381 (N_4381,N_4285,N_4265);
and U4382 (N_4382,N_4285,N_4215);
or U4383 (N_4383,N_4260,N_4295);
nand U4384 (N_4384,N_4286,N_4278);
and U4385 (N_4385,N_4266,N_4228);
nor U4386 (N_4386,N_4206,N_4204);
nor U4387 (N_4387,N_4249,N_4248);
and U4388 (N_4388,N_4214,N_4245);
nand U4389 (N_4389,N_4254,N_4200);
or U4390 (N_4390,N_4291,N_4230);
nand U4391 (N_4391,N_4238,N_4299);
nor U4392 (N_4392,N_4208,N_4275);
nor U4393 (N_4393,N_4214,N_4257);
or U4394 (N_4394,N_4243,N_4242);
and U4395 (N_4395,N_4207,N_4246);
nand U4396 (N_4396,N_4200,N_4217);
nand U4397 (N_4397,N_4201,N_4225);
xnor U4398 (N_4398,N_4220,N_4276);
nor U4399 (N_4399,N_4225,N_4244);
nand U4400 (N_4400,N_4376,N_4374);
nor U4401 (N_4401,N_4360,N_4397);
and U4402 (N_4402,N_4383,N_4363);
and U4403 (N_4403,N_4355,N_4317);
xnor U4404 (N_4404,N_4356,N_4375);
or U4405 (N_4405,N_4344,N_4329);
xnor U4406 (N_4406,N_4315,N_4309);
or U4407 (N_4407,N_4366,N_4357);
nor U4408 (N_4408,N_4354,N_4379);
nand U4409 (N_4409,N_4378,N_4393);
nor U4410 (N_4410,N_4332,N_4380);
nor U4411 (N_4411,N_4311,N_4390);
and U4412 (N_4412,N_4326,N_4386);
and U4413 (N_4413,N_4391,N_4305);
or U4414 (N_4414,N_4396,N_4334);
and U4415 (N_4415,N_4385,N_4389);
nor U4416 (N_4416,N_4324,N_4325);
nand U4417 (N_4417,N_4306,N_4312);
nor U4418 (N_4418,N_4384,N_4337);
nor U4419 (N_4419,N_4399,N_4319);
and U4420 (N_4420,N_4343,N_4394);
or U4421 (N_4421,N_4345,N_4364);
nand U4422 (N_4422,N_4370,N_4327);
nand U4423 (N_4423,N_4308,N_4322);
nand U4424 (N_4424,N_4395,N_4362);
or U4425 (N_4425,N_4352,N_4333);
and U4426 (N_4426,N_4307,N_4369);
nor U4427 (N_4427,N_4328,N_4361);
and U4428 (N_4428,N_4341,N_4381);
or U4429 (N_4429,N_4316,N_4365);
and U4430 (N_4430,N_4377,N_4351);
or U4431 (N_4431,N_4372,N_4321);
or U4432 (N_4432,N_4388,N_4339);
or U4433 (N_4433,N_4350,N_4392);
nor U4434 (N_4434,N_4349,N_4346);
nor U4435 (N_4435,N_4368,N_4373);
nand U4436 (N_4436,N_4314,N_4382);
and U4437 (N_4437,N_4398,N_4301);
nor U4438 (N_4438,N_4313,N_4320);
nand U4439 (N_4439,N_4353,N_4367);
and U4440 (N_4440,N_4335,N_4331);
nand U4441 (N_4441,N_4338,N_4303);
and U4442 (N_4442,N_4330,N_4340);
or U4443 (N_4443,N_4318,N_4347);
or U4444 (N_4444,N_4302,N_4358);
and U4445 (N_4445,N_4371,N_4304);
or U4446 (N_4446,N_4359,N_4300);
or U4447 (N_4447,N_4323,N_4310);
or U4448 (N_4448,N_4342,N_4387);
and U4449 (N_4449,N_4348,N_4336);
nor U4450 (N_4450,N_4337,N_4354);
nand U4451 (N_4451,N_4333,N_4377);
nand U4452 (N_4452,N_4344,N_4390);
nand U4453 (N_4453,N_4324,N_4306);
and U4454 (N_4454,N_4380,N_4336);
nand U4455 (N_4455,N_4354,N_4307);
and U4456 (N_4456,N_4360,N_4370);
or U4457 (N_4457,N_4353,N_4384);
or U4458 (N_4458,N_4319,N_4359);
nor U4459 (N_4459,N_4334,N_4346);
and U4460 (N_4460,N_4308,N_4342);
nand U4461 (N_4461,N_4322,N_4346);
or U4462 (N_4462,N_4346,N_4388);
nand U4463 (N_4463,N_4371,N_4381);
nor U4464 (N_4464,N_4382,N_4342);
or U4465 (N_4465,N_4329,N_4346);
nor U4466 (N_4466,N_4364,N_4300);
nor U4467 (N_4467,N_4346,N_4351);
and U4468 (N_4468,N_4347,N_4387);
or U4469 (N_4469,N_4361,N_4310);
nand U4470 (N_4470,N_4307,N_4323);
or U4471 (N_4471,N_4337,N_4359);
nor U4472 (N_4472,N_4363,N_4396);
nand U4473 (N_4473,N_4300,N_4395);
and U4474 (N_4474,N_4381,N_4339);
nor U4475 (N_4475,N_4340,N_4383);
and U4476 (N_4476,N_4392,N_4383);
nand U4477 (N_4477,N_4386,N_4383);
or U4478 (N_4478,N_4309,N_4357);
nand U4479 (N_4479,N_4320,N_4396);
or U4480 (N_4480,N_4303,N_4341);
or U4481 (N_4481,N_4338,N_4378);
nor U4482 (N_4482,N_4334,N_4358);
nor U4483 (N_4483,N_4316,N_4381);
or U4484 (N_4484,N_4375,N_4318);
nor U4485 (N_4485,N_4353,N_4382);
or U4486 (N_4486,N_4323,N_4319);
or U4487 (N_4487,N_4351,N_4375);
or U4488 (N_4488,N_4362,N_4322);
nor U4489 (N_4489,N_4378,N_4313);
or U4490 (N_4490,N_4370,N_4317);
nand U4491 (N_4491,N_4327,N_4335);
nand U4492 (N_4492,N_4325,N_4387);
and U4493 (N_4493,N_4353,N_4398);
or U4494 (N_4494,N_4306,N_4310);
and U4495 (N_4495,N_4344,N_4346);
or U4496 (N_4496,N_4342,N_4306);
and U4497 (N_4497,N_4312,N_4352);
nor U4498 (N_4498,N_4372,N_4381);
or U4499 (N_4499,N_4380,N_4350);
or U4500 (N_4500,N_4442,N_4451);
nand U4501 (N_4501,N_4405,N_4450);
and U4502 (N_4502,N_4454,N_4424);
nor U4503 (N_4503,N_4462,N_4470);
nand U4504 (N_4504,N_4474,N_4495);
nor U4505 (N_4505,N_4438,N_4425);
or U4506 (N_4506,N_4466,N_4414);
nor U4507 (N_4507,N_4464,N_4422);
nor U4508 (N_4508,N_4481,N_4435);
nand U4509 (N_4509,N_4410,N_4465);
nor U4510 (N_4510,N_4413,N_4460);
and U4511 (N_4511,N_4416,N_4403);
nor U4512 (N_4512,N_4487,N_4491);
nand U4513 (N_4513,N_4488,N_4404);
nand U4514 (N_4514,N_4431,N_4494);
nand U4515 (N_4515,N_4428,N_4401);
nand U4516 (N_4516,N_4444,N_4443);
xor U4517 (N_4517,N_4402,N_4400);
nand U4518 (N_4518,N_4420,N_4483);
nand U4519 (N_4519,N_4423,N_4406);
nand U4520 (N_4520,N_4455,N_4469);
nand U4521 (N_4521,N_4445,N_4452);
or U4522 (N_4522,N_4434,N_4473);
or U4523 (N_4523,N_4479,N_4418);
and U4524 (N_4524,N_4419,N_4477);
or U4525 (N_4525,N_4426,N_4478);
xor U4526 (N_4526,N_4446,N_4489);
nand U4527 (N_4527,N_4412,N_4484);
nand U4528 (N_4528,N_4453,N_4440);
and U4529 (N_4529,N_4417,N_4436);
nand U4530 (N_4530,N_4471,N_4496);
nand U4531 (N_4531,N_4441,N_4421);
and U4532 (N_4532,N_4497,N_4456);
nor U4533 (N_4533,N_4476,N_4463);
nor U4534 (N_4534,N_4490,N_4448);
nor U4535 (N_4535,N_4447,N_4415);
and U4536 (N_4536,N_4411,N_4475);
nor U4537 (N_4537,N_4429,N_4409);
or U4538 (N_4538,N_4459,N_4407);
or U4539 (N_4539,N_4432,N_4439);
or U4540 (N_4540,N_4449,N_4467);
and U4541 (N_4541,N_4492,N_4480);
nor U4542 (N_4542,N_4430,N_4408);
and U4543 (N_4543,N_4433,N_4427);
and U4544 (N_4544,N_4472,N_4486);
xor U4545 (N_4545,N_4485,N_4499);
and U4546 (N_4546,N_4493,N_4458);
nand U4547 (N_4547,N_4461,N_4468);
nand U4548 (N_4548,N_4457,N_4498);
and U4549 (N_4549,N_4482,N_4437);
or U4550 (N_4550,N_4424,N_4486);
nand U4551 (N_4551,N_4454,N_4446);
nand U4552 (N_4552,N_4496,N_4498);
and U4553 (N_4553,N_4461,N_4457);
nor U4554 (N_4554,N_4429,N_4472);
or U4555 (N_4555,N_4410,N_4456);
nand U4556 (N_4556,N_4480,N_4490);
or U4557 (N_4557,N_4469,N_4403);
and U4558 (N_4558,N_4475,N_4489);
or U4559 (N_4559,N_4438,N_4472);
nor U4560 (N_4560,N_4415,N_4464);
nand U4561 (N_4561,N_4489,N_4481);
nand U4562 (N_4562,N_4460,N_4431);
nand U4563 (N_4563,N_4474,N_4413);
or U4564 (N_4564,N_4490,N_4474);
and U4565 (N_4565,N_4461,N_4421);
and U4566 (N_4566,N_4475,N_4471);
or U4567 (N_4567,N_4422,N_4436);
and U4568 (N_4568,N_4484,N_4440);
or U4569 (N_4569,N_4427,N_4453);
or U4570 (N_4570,N_4487,N_4421);
or U4571 (N_4571,N_4486,N_4454);
nand U4572 (N_4572,N_4415,N_4450);
or U4573 (N_4573,N_4490,N_4456);
nor U4574 (N_4574,N_4494,N_4457);
nor U4575 (N_4575,N_4444,N_4474);
nand U4576 (N_4576,N_4489,N_4436);
and U4577 (N_4577,N_4437,N_4429);
nand U4578 (N_4578,N_4453,N_4400);
and U4579 (N_4579,N_4463,N_4442);
or U4580 (N_4580,N_4481,N_4403);
nor U4581 (N_4581,N_4480,N_4461);
nor U4582 (N_4582,N_4495,N_4406);
nor U4583 (N_4583,N_4475,N_4413);
nand U4584 (N_4584,N_4426,N_4442);
nand U4585 (N_4585,N_4434,N_4461);
nand U4586 (N_4586,N_4444,N_4462);
or U4587 (N_4587,N_4452,N_4423);
nor U4588 (N_4588,N_4485,N_4422);
nand U4589 (N_4589,N_4492,N_4448);
and U4590 (N_4590,N_4413,N_4436);
nor U4591 (N_4591,N_4440,N_4495);
nand U4592 (N_4592,N_4472,N_4404);
xor U4593 (N_4593,N_4468,N_4493);
nor U4594 (N_4594,N_4472,N_4463);
or U4595 (N_4595,N_4478,N_4436);
nand U4596 (N_4596,N_4493,N_4481);
nand U4597 (N_4597,N_4475,N_4404);
nor U4598 (N_4598,N_4470,N_4466);
or U4599 (N_4599,N_4412,N_4487);
nand U4600 (N_4600,N_4524,N_4589);
nand U4601 (N_4601,N_4562,N_4532);
nand U4602 (N_4602,N_4515,N_4507);
or U4603 (N_4603,N_4558,N_4556);
or U4604 (N_4604,N_4519,N_4549);
or U4605 (N_4605,N_4512,N_4580);
and U4606 (N_4606,N_4547,N_4590);
or U4607 (N_4607,N_4568,N_4505);
nand U4608 (N_4608,N_4594,N_4537);
or U4609 (N_4609,N_4551,N_4536);
xor U4610 (N_4610,N_4591,N_4557);
and U4611 (N_4611,N_4566,N_4542);
and U4612 (N_4612,N_4576,N_4555);
or U4613 (N_4613,N_4593,N_4563);
or U4614 (N_4614,N_4523,N_4578);
or U4615 (N_4615,N_4584,N_4560);
or U4616 (N_4616,N_4569,N_4572);
or U4617 (N_4617,N_4599,N_4503);
nand U4618 (N_4618,N_4574,N_4544);
or U4619 (N_4619,N_4526,N_4518);
xor U4620 (N_4620,N_4514,N_4564);
nand U4621 (N_4621,N_4545,N_4535);
and U4622 (N_4622,N_4529,N_4582);
and U4623 (N_4623,N_4501,N_4531);
nand U4624 (N_4624,N_4504,N_4595);
nor U4625 (N_4625,N_4525,N_4527);
or U4626 (N_4626,N_4534,N_4575);
and U4627 (N_4627,N_4573,N_4543);
or U4628 (N_4628,N_4509,N_4520);
and U4629 (N_4629,N_4521,N_4567);
or U4630 (N_4630,N_4502,N_4596);
nor U4631 (N_4631,N_4539,N_4587);
and U4632 (N_4632,N_4553,N_4554);
nand U4633 (N_4633,N_4516,N_4538);
and U4634 (N_4634,N_4581,N_4579);
nand U4635 (N_4635,N_4541,N_4585);
and U4636 (N_4636,N_4565,N_4597);
nor U4637 (N_4637,N_4508,N_4570);
nor U4638 (N_4638,N_4552,N_4533);
xor U4639 (N_4639,N_4559,N_4546);
or U4640 (N_4640,N_4522,N_4528);
nand U4641 (N_4641,N_4530,N_4588);
and U4642 (N_4642,N_4500,N_4571);
or U4643 (N_4643,N_4510,N_4548);
nor U4644 (N_4644,N_4517,N_4598);
nand U4645 (N_4645,N_4506,N_4586);
and U4646 (N_4646,N_4511,N_4592);
or U4647 (N_4647,N_4513,N_4561);
xnor U4648 (N_4648,N_4577,N_4540);
and U4649 (N_4649,N_4583,N_4550);
or U4650 (N_4650,N_4592,N_4543);
or U4651 (N_4651,N_4560,N_4511);
nor U4652 (N_4652,N_4563,N_4540);
nor U4653 (N_4653,N_4555,N_4553);
or U4654 (N_4654,N_4581,N_4589);
nor U4655 (N_4655,N_4571,N_4555);
nand U4656 (N_4656,N_4561,N_4502);
or U4657 (N_4657,N_4595,N_4555);
and U4658 (N_4658,N_4550,N_4506);
nand U4659 (N_4659,N_4583,N_4507);
nand U4660 (N_4660,N_4590,N_4521);
nor U4661 (N_4661,N_4527,N_4518);
or U4662 (N_4662,N_4588,N_4558);
or U4663 (N_4663,N_4592,N_4548);
nor U4664 (N_4664,N_4544,N_4558);
and U4665 (N_4665,N_4572,N_4520);
nand U4666 (N_4666,N_4535,N_4536);
nand U4667 (N_4667,N_4544,N_4571);
or U4668 (N_4668,N_4520,N_4513);
and U4669 (N_4669,N_4596,N_4583);
and U4670 (N_4670,N_4533,N_4530);
and U4671 (N_4671,N_4599,N_4585);
nand U4672 (N_4672,N_4539,N_4534);
nand U4673 (N_4673,N_4596,N_4514);
and U4674 (N_4674,N_4539,N_4545);
and U4675 (N_4675,N_4522,N_4512);
and U4676 (N_4676,N_4518,N_4541);
nor U4677 (N_4677,N_4599,N_4527);
or U4678 (N_4678,N_4579,N_4592);
and U4679 (N_4679,N_4504,N_4544);
and U4680 (N_4680,N_4555,N_4585);
nor U4681 (N_4681,N_4505,N_4518);
nand U4682 (N_4682,N_4568,N_4538);
nand U4683 (N_4683,N_4541,N_4544);
nand U4684 (N_4684,N_4538,N_4531);
or U4685 (N_4685,N_4560,N_4549);
and U4686 (N_4686,N_4599,N_4520);
nand U4687 (N_4687,N_4534,N_4556);
xnor U4688 (N_4688,N_4575,N_4511);
nand U4689 (N_4689,N_4588,N_4529);
or U4690 (N_4690,N_4567,N_4555);
nor U4691 (N_4691,N_4561,N_4553);
nand U4692 (N_4692,N_4571,N_4581);
and U4693 (N_4693,N_4572,N_4535);
and U4694 (N_4694,N_4517,N_4534);
nor U4695 (N_4695,N_4561,N_4573);
or U4696 (N_4696,N_4562,N_4551);
nand U4697 (N_4697,N_4554,N_4515);
and U4698 (N_4698,N_4540,N_4538);
nor U4699 (N_4699,N_4527,N_4576);
or U4700 (N_4700,N_4671,N_4634);
or U4701 (N_4701,N_4614,N_4662);
nor U4702 (N_4702,N_4696,N_4680);
nor U4703 (N_4703,N_4678,N_4620);
nand U4704 (N_4704,N_4665,N_4639);
and U4705 (N_4705,N_4691,N_4655);
or U4706 (N_4706,N_4643,N_4669);
or U4707 (N_4707,N_4674,N_4605);
nand U4708 (N_4708,N_4627,N_4670);
and U4709 (N_4709,N_4686,N_4623);
nand U4710 (N_4710,N_4641,N_4603);
nand U4711 (N_4711,N_4606,N_4621);
and U4712 (N_4712,N_4663,N_4683);
or U4713 (N_4713,N_4648,N_4612);
and U4714 (N_4714,N_4616,N_4650);
nor U4715 (N_4715,N_4653,N_4672);
or U4716 (N_4716,N_4673,N_4654);
nand U4717 (N_4717,N_4637,N_4636);
and U4718 (N_4718,N_4695,N_4681);
or U4719 (N_4719,N_4689,N_4611);
and U4720 (N_4720,N_4658,N_4600);
nand U4721 (N_4721,N_4630,N_4690);
nor U4722 (N_4722,N_4632,N_4601);
and U4723 (N_4723,N_4624,N_4613);
nor U4724 (N_4724,N_4617,N_4646);
or U4725 (N_4725,N_4607,N_4638);
nand U4726 (N_4726,N_4692,N_4608);
nand U4727 (N_4727,N_4642,N_4640);
or U4728 (N_4728,N_4676,N_4619);
and U4729 (N_4729,N_4664,N_4697);
nor U4730 (N_4730,N_4647,N_4698);
nor U4731 (N_4731,N_4657,N_4661);
nand U4732 (N_4732,N_4625,N_4666);
nor U4733 (N_4733,N_4687,N_4685);
nand U4734 (N_4734,N_4629,N_4610);
or U4735 (N_4735,N_4652,N_4649);
and U4736 (N_4736,N_4659,N_4677);
or U4737 (N_4737,N_4682,N_4618);
and U4738 (N_4738,N_4628,N_4615);
and U4739 (N_4739,N_4604,N_4602);
nand U4740 (N_4740,N_4645,N_4679);
and U4741 (N_4741,N_4675,N_4626);
and U4742 (N_4742,N_4693,N_4694);
and U4743 (N_4743,N_4699,N_4651);
or U4744 (N_4744,N_4631,N_4684);
or U4745 (N_4745,N_4622,N_4633);
or U4746 (N_4746,N_4668,N_4656);
or U4747 (N_4747,N_4635,N_4644);
nand U4748 (N_4748,N_4660,N_4688);
or U4749 (N_4749,N_4609,N_4667);
nand U4750 (N_4750,N_4667,N_4652);
and U4751 (N_4751,N_4697,N_4627);
or U4752 (N_4752,N_4650,N_4685);
nand U4753 (N_4753,N_4614,N_4653);
or U4754 (N_4754,N_4652,N_4621);
nand U4755 (N_4755,N_4689,N_4685);
and U4756 (N_4756,N_4660,N_4618);
or U4757 (N_4757,N_4620,N_4640);
nand U4758 (N_4758,N_4657,N_4629);
nand U4759 (N_4759,N_4614,N_4668);
nand U4760 (N_4760,N_4602,N_4672);
nor U4761 (N_4761,N_4685,N_4642);
or U4762 (N_4762,N_4695,N_4692);
nand U4763 (N_4763,N_4625,N_4676);
and U4764 (N_4764,N_4602,N_4654);
or U4765 (N_4765,N_4666,N_4635);
or U4766 (N_4766,N_4619,N_4631);
nand U4767 (N_4767,N_4699,N_4686);
or U4768 (N_4768,N_4628,N_4683);
nand U4769 (N_4769,N_4642,N_4603);
nor U4770 (N_4770,N_4605,N_4631);
and U4771 (N_4771,N_4633,N_4636);
or U4772 (N_4772,N_4696,N_4654);
or U4773 (N_4773,N_4666,N_4653);
nand U4774 (N_4774,N_4610,N_4684);
and U4775 (N_4775,N_4631,N_4681);
nand U4776 (N_4776,N_4642,N_4609);
or U4777 (N_4777,N_4605,N_4635);
nand U4778 (N_4778,N_4657,N_4620);
nand U4779 (N_4779,N_4645,N_4665);
nand U4780 (N_4780,N_4691,N_4674);
nand U4781 (N_4781,N_4673,N_4619);
nand U4782 (N_4782,N_4600,N_4633);
nand U4783 (N_4783,N_4662,N_4692);
or U4784 (N_4784,N_4628,N_4691);
nand U4785 (N_4785,N_4622,N_4626);
or U4786 (N_4786,N_4691,N_4620);
and U4787 (N_4787,N_4693,N_4662);
nand U4788 (N_4788,N_4603,N_4638);
xor U4789 (N_4789,N_4674,N_4650);
or U4790 (N_4790,N_4654,N_4643);
nand U4791 (N_4791,N_4638,N_4624);
or U4792 (N_4792,N_4697,N_4654);
nor U4793 (N_4793,N_4611,N_4624);
or U4794 (N_4794,N_4651,N_4642);
and U4795 (N_4795,N_4659,N_4643);
nand U4796 (N_4796,N_4664,N_4648);
nor U4797 (N_4797,N_4638,N_4684);
and U4798 (N_4798,N_4680,N_4655);
nand U4799 (N_4799,N_4633,N_4608);
nand U4800 (N_4800,N_4746,N_4705);
or U4801 (N_4801,N_4772,N_4775);
nor U4802 (N_4802,N_4755,N_4756);
or U4803 (N_4803,N_4716,N_4745);
or U4804 (N_4804,N_4764,N_4760);
or U4805 (N_4805,N_4701,N_4717);
and U4806 (N_4806,N_4720,N_4734);
nor U4807 (N_4807,N_4744,N_4795);
or U4808 (N_4808,N_4740,N_4796);
nand U4809 (N_4809,N_4713,N_4769);
or U4810 (N_4810,N_4776,N_4719);
or U4811 (N_4811,N_4786,N_4704);
and U4812 (N_4812,N_4735,N_4798);
nor U4813 (N_4813,N_4784,N_4788);
and U4814 (N_4814,N_4765,N_4709);
and U4815 (N_4815,N_4763,N_4791);
nand U4816 (N_4816,N_4748,N_4758);
nand U4817 (N_4817,N_4707,N_4773);
nor U4818 (N_4818,N_4790,N_4759);
nor U4819 (N_4819,N_4723,N_4751);
or U4820 (N_4820,N_4762,N_4792);
nand U4821 (N_4821,N_4778,N_4767);
nor U4822 (N_4822,N_4726,N_4774);
or U4823 (N_4823,N_4712,N_4711);
or U4824 (N_4824,N_4797,N_4727);
nand U4825 (N_4825,N_4715,N_4789);
xnor U4826 (N_4826,N_4749,N_4737);
nor U4827 (N_4827,N_4700,N_4742);
nor U4828 (N_4828,N_4722,N_4732);
nand U4829 (N_4829,N_4768,N_4757);
and U4830 (N_4830,N_4702,N_4783);
nor U4831 (N_4831,N_4766,N_4771);
nand U4832 (N_4832,N_4787,N_4718);
or U4833 (N_4833,N_4733,N_4714);
and U4834 (N_4834,N_4761,N_4736);
and U4835 (N_4835,N_4779,N_4782);
or U4836 (N_4836,N_4780,N_4793);
xor U4837 (N_4837,N_4724,N_4741);
and U4838 (N_4838,N_4799,N_4731);
or U4839 (N_4839,N_4777,N_4781);
and U4840 (N_4840,N_4750,N_4752);
and U4841 (N_4841,N_4729,N_4703);
nand U4842 (N_4842,N_4725,N_4708);
nand U4843 (N_4843,N_4730,N_4721);
and U4844 (N_4844,N_4794,N_4710);
and U4845 (N_4845,N_4738,N_4728);
and U4846 (N_4846,N_4754,N_4785);
and U4847 (N_4847,N_4747,N_4739);
or U4848 (N_4848,N_4706,N_4770);
nor U4849 (N_4849,N_4743,N_4753);
nand U4850 (N_4850,N_4766,N_4731);
nor U4851 (N_4851,N_4756,N_4712);
and U4852 (N_4852,N_4779,N_4799);
nand U4853 (N_4853,N_4759,N_4708);
nor U4854 (N_4854,N_4773,N_4741);
and U4855 (N_4855,N_4759,N_4761);
and U4856 (N_4856,N_4736,N_4775);
or U4857 (N_4857,N_4765,N_4740);
nand U4858 (N_4858,N_4772,N_4720);
nor U4859 (N_4859,N_4701,N_4723);
and U4860 (N_4860,N_4736,N_4706);
or U4861 (N_4861,N_4728,N_4779);
nand U4862 (N_4862,N_4745,N_4730);
nor U4863 (N_4863,N_4787,N_4772);
and U4864 (N_4864,N_4756,N_4758);
xnor U4865 (N_4865,N_4782,N_4788);
nor U4866 (N_4866,N_4706,N_4725);
nand U4867 (N_4867,N_4764,N_4762);
nand U4868 (N_4868,N_4778,N_4717);
nand U4869 (N_4869,N_4767,N_4719);
nand U4870 (N_4870,N_4778,N_4705);
or U4871 (N_4871,N_4704,N_4719);
nand U4872 (N_4872,N_4716,N_4781);
and U4873 (N_4873,N_4745,N_4796);
and U4874 (N_4874,N_4745,N_4732);
nand U4875 (N_4875,N_4719,N_4799);
nand U4876 (N_4876,N_4737,N_4734);
and U4877 (N_4877,N_4722,N_4741);
or U4878 (N_4878,N_4784,N_4766);
or U4879 (N_4879,N_4760,N_4701);
or U4880 (N_4880,N_4773,N_4799);
nor U4881 (N_4881,N_4705,N_4748);
and U4882 (N_4882,N_4778,N_4753);
and U4883 (N_4883,N_4740,N_4714);
nand U4884 (N_4884,N_4722,N_4723);
nand U4885 (N_4885,N_4785,N_4793);
or U4886 (N_4886,N_4702,N_4778);
or U4887 (N_4887,N_4750,N_4744);
and U4888 (N_4888,N_4759,N_4758);
nor U4889 (N_4889,N_4740,N_4760);
nand U4890 (N_4890,N_4765,N_4776);
and U4891 (N_4891,N_4732,N_4755);
or U4892 (N_4892,N_4761,N_4765);
nor U4893 (N_4893,N_4770,N_4726);
and U4894 (N_4894,N_4799,N_4726);
and U4895 (N_4895,N_4722,N_4724);
or U4896 (N_4896,N_4781,N_4753);
and U4897 (N_4897,N_4720,N_4723);
or U4898 (N_4898,N_4777,N_4711);
nand U4899 (N_4899,N_4763,N_4756);
or U4900 (N_4900,N_4841,N_4853);
xor U4901 (N_4901,N_4885,N_4875);
nand U4902 (N_4902,N_4840,N_4834);
or U4903 (N_4903,N_4827,N_4874);
xor U4904 (N_4904,N_4835,N_4807);
or U4905 (N_4905,N_4802,N_4871);
or U4906 (N_4906,N_4829,N_4845);
and U4907 (N_4907,N_4878,N_4861);
and U4908 (N_4908,N_4877,N_4839);
nor U4909 (N_4909,N_4806,N_4820);
nor U4910 (N_4910,N_4867,N_4837);
nor U4911 (N_4911,N_4855,N_4823);
nor U4912 (N_4912,N_4844,N_4838);
and U4913 (N_4913,N_4860,N_4880);
nand U4914 (N_4914,N_4819,N_4882);
and U4915 (N_4915,N_4825,N_4826);
nor U4916 (N_4916,N_4887,N_4873);
nand U4917 (N_4917,N_4881,N_4863);
nand U4918 (N_4918,N_4811,N_4824);
and U4919 (N_4919,N_4857,N_4865);
nor U4920 (N_4920,N_4894,N_4864);
and U4921 (N_4921,N_4862,N_4804);
nor U4922 (N_4922,N_4868,N_4859);
nand U4923 (N_4923,N_4801,N_4828);
nor U4924 (N_4924,N_4870,N_4879);
nor U4925 (N_4925,N_4842,N_4850);
xnor U4926 (N_4926,N_4832,N_4890);
and U4927 (N_4927,N_4833,N_4866);
and U4928 (N_4928,N_4897,N_4893);
and U4929 (N_4929,N_4852,N_4815);
nand U4930 (N_4930,N_4883,N_4872);
and U4931 (N_4931,N_4822,N_4803);
nand U4932 (N_4932,N_4817,N_4814);
nand U4933 (N_4933,N_4847,N_4813);
nand U4934 (N_4934,N_4895,N_4896);
or U4935 (N_4935,N_4800,N_4869);
nand U4936 (N_4936,N_4899,N_4898);
nor U4937 (N_4937,N_4821,N_4884);
and U4938 (N_4938,N_4831,N_4808);
nand U4939 (N_4939,N_4889,N_4854);
and U4940 (N_4940,N_4810,N_4848);
nor U4941 (N_4941,N_4858,N_4886);
and U4942 (N_4942,N_4816,N_4818);
or U4943 (N_4943,N_4846,N_4888);
nand U4944 (N_4944,N_4843,N_4892);
xnor U4945 (N_4945,N_4812,N_4830);
and U4946 (N_4946,N_4891,N_4856);
and U4947 (N_4947,N_4876,N_4809);
and U4948 (N_4948,N_4805,N_4849);
xor U4949 (N_4949,N_4836,N_4851);
and U4950 (N_4950,N_4864,N_4842);
nand U4951 (N_4951,N_4807,N_4810);
nor U4952 (N_4952,N_4867,N_4808);
and U4953 (N_4953,N_4891,N_4885);
nand U4954 (N_4954,N_4890,N_4852);
or U4955 (N_4955,N_4830,N_4821);
nand U4956 (N_4956,N_4899,N_4808);
xor U4957 (N_4957,N_4871,N_4833);
or U4958 (N_4958,N_4808,N_4827);
and U4959 (N_4959,N_4847,N_4854);
nor U4960 (N_4960,N_4894,N_4813);
or U4961 (N_4961,N_4876,N_4823);
nand U4962 (N_4962,N_4868,N_4805);
nand U4963 (N_4963,N_4870,N_4855);
nor U4964 (N_4964,N_4897,N_4869);
nand U4965 (N_4965,N_4823,N_4800);
xnor U4966 (N_4966,N_4834,N_4895);
nand U4967 (N_4967,N_4830,N_4850);
xor U4968 (N_4968,N_4895,N_4810);
nand U4969 (N_4969,N_4806,N_4815);
nand U4970 (N_4970,N_4820,N_4815);
nor U4971 (N_4971,N_4895,N_4815);
nor U4972 (N_4972,N_4889,N_4801);
nor U4973 (N_4973,N_4817,N_4873);
nand U4974 (N_4974,N_4843,N_4823);
or U4975 (N_4975,N_4844,N_4894);
nor U4976 (N_4976,N_4827,N_4837);
nor U4977 (N_4977,N_4881,N_4823);
nand U4978 (N_4978,N_4878,N_4847);
nor U4979 (N_4979,N_4810,N_4872);
and U4980 (N_4980,N_4837,N_4895);
nand U4981 (N_4981,N_4819,N_4875);
nor U4982 (N_4982,N_4826,N_4831);
and U4983 (N_4983,N_4835,N_4819);
or U4984 (N_4984,N_4827,N_4840);
and U4985 (N_4985,N_4877,N_4808);
nand U4986 (N_4986,N_4803,N_4809);
xor U4987 (N_4987,N_4873,N_4862);
or U4988 (N_4988,N_4855,N_4858);
nor U4989 (N_4989,N_4829,N_4858);
and U4990 (N_4990,N_4869,N_4856);
and U4991 (N_4991,N_4844,N_4878);
or U4992 (N_4992,N_4812,N_4860);
nand U4993 (N_4993,N_4808,N_4848);
and U4994 (N_4994,N_4830,N_4819);
and U4995 (N_4995,N_4885,N_4890);
and U4996 (N_4996,N_4880,N_4893);
nor U4997 (N_4997,N_4835,N_4849);
and U4998 (N_4998,N_4857,N_4869);
xor U4999 (N_4999,N_4856,N_4893);
and UO_0 (O_0,N_4996,N_4952);
and UO_1 (O_1,N_4964,N_4966);
xor UO_2 (O_2,N_4905,N_4965);
nand UO_3 (O_3,N_4981,N_4992);
and UO_4 (O_4,N_4971,N_4994);
nand UO_5 (O_5,N_4954,N_4987);
nand UO_6 (O_6,N_4917,N_4972);
or UO_7 (O_7,N_4922,N_4923);
or UO_8 (O_8,N_4913,N_4989);
nand UO_9 (O_9,N_4931,N_4961);
nand UO_10 (O_10,N_4963,N_4962);
and UO_11 (O_11,N_4948,N_4937);
or UO_12 (O_12,N_4943,N_4924);
nand UO_13 (O_13,N_4990,N_4951);
or UO_14 (O_14,N_4983,N_4984);
nor UO_15 (O_15,N_4955,N_4926);
or UO_16 (O_16,N_4918,N_4998);
nand UO_17 (O_17,N_4950,N_4995);
nand UO_18 (O_18,N_4925,N_4945);
nand UO_19 (O_19,N_4970,N_4977);
nor UO_20 (O_20,N_4919,N_4932);
and UO_21 (O_21,N_4974,N_4973);
nand UO_22 (O_22,N_4959,N_4921);
and UO_23 (O_23,N_4979,N_4910);
nor UO_24 (O_24,N_4929,N_4982);
nor UO_25 (O_25,N_4942,N_4988);
and UO_26 (O_26,N_4911,N_4960);
nand UO_27 (O_27,N_4900,N_4933);
or UO_28 (O_28,N_4935,N_4993);
nor UO_29 (O_29,N_4944,N_4916);
and UO_30 (O_30,N_4901,N_4914);
nand UO_31 (O_31,N_4907,N_4949);
and UO_32 (O_32,N_4938,N_4978);
and UO_33 (O_33,N_4956,N_4991);
xor UO_34 (O_34,N_4947,N_4928);
nand UO_35 (O_35,N_4934,N_4909);
nand UO_36 (O_36,N_4906,N_4969);
nor UO_37 (O_37,N_4980,N_4912);
nand UO_38 (O_38,N_4936,N_4908);
or UO_39 (O_39,N_4903,N_4986);
and UO_40 (O_40,N_4975,N_4939);
nor UO_41 (O_41,N_4927,N_4941);
or UO_42 (O_42,N_4999,N_4930);
or UO_43 (O_43,N_4985,N_4976);
and UO_44 (O_44,N_4968,N_4958);
xor UO_45 (O_45,N_4902,N_4953);
nor UO_46 (O_46,N_4957,N_4915);
nor UO_47 (O_47,N_4920,N_4997);
and UO_48 (O_48,N_4946,N_4940);
or UO_49 (O_49,N_4904,N_4967);
nand UO_50 (O_50,N_4966,N_4949);
nor UO_51 (O_51,N_4996,N_4927);
nor UO_52 (O_52,N_4969,N_4965);
nand UO_53 (O_53,N_4962,N_4965);
and UO_54 (O_54,N_4994,N_4978);
and UO_55 (O_55,N_4938,N_4944);
nor UO_56 (O_56,N_4915,N_4924);
or UO_57 (O_57,N_4999,N_4949);
nand UO_58 (O_58,N_4933,N_4978);
and UO_59 (O_59,N_4989,N_4974);
and UO_60 (O_60,N_4912,N_4956);
nor UO_61 (O_61,N_4900,N_4968);
or UO_62 (O_62,N_4912,N_4954);
nor UO_63 (O_63,N_4911,N_4981);
nand UO_64 (O_64,N_4958,N_4967);
nand UO_65 (O_65,N_4923,N_4979);
nand UO_66 (O_66,N_4969,N_4985);
or UO_67 (O_67,N_4918,N_4936);
xnor UO_68 (O_68,N_4964,N_4935);
nor UO_69 (O_69,N_4923,N_4936);
xor UO_70 (O_70,N_4934,N_4977);
or UO_71 (O_71,N_4962,N_4905);
xor UO_72 (O_72,N_4990,N_4927);
or UO_73 (O_73,N_4939,N_4927);
nor UO_74 (O_74,N_4948,N_4908);
and UO_75 (O_75,N_4975,N_4925);
and UO_76 (O_76,N_4994,N_4950);
nand UO_77 (O_77,N_4991,N_4927);
nor UO_78 (O_78,N_4954,N_4915);
and UO_79 (O_79,N_4931,N_4971);
nor UO_80 (O_80,N_4906,N_4983);
and UO_81 (O_81,N_4979,N_4986);
xnor UO_82 (O_82,N_4952,N_4975);
nor UO_83 (O_83,N_4940,N_4958);
and UO_84 (O_84,N_4956,N_4985);
nand UO_85 (O_85,N_4926,N_4957);
nand UO_86 (O_86,N_4976,N_4949);
nor UO_87 (O_87,N_4965,N_4904);
or UO_88 (O_88,N_4962,N_4945);
and UO_89 (O_89,N_4929,N_4964);
and UO_90 (O_90,N_4940,N_4982);
nand UO_91 (O_91,N_4973,N_4988);
nor UO_92 (O_92,N_4915,N_4953);
or UO_93 (O_93,N_4999,N_4981);
and UO_94 (O_94,N_4907,N_4917);
and UO_95 (O_95,N_4941,N_4980);
nand UO_96 (O_96,N_4974,N_4924);
or UO_97 (O_97,N_4901,N_4968);
and UO_98 (O_98,N_4972,N_4979);
xnor UO_99 (O_99,N_4972,N_4944);
nand UO_100 (O_100,N_4960,N_4992);
nor UO_101 (O_101,N_4923,N_4928);
nand UO_102 (O_102,N_4968,N_4936);
nand UO_103 (O_103,N_4958,N_4965);
nand UO_104 (O_104,N_4990,N_4993);
nand UO_105 (O_105,N_4949,N_4935);
or UO_106 (O_106,N_4923,N_4977);
nand UO_107 (O_107,N_4909,N_4925);
nor UO_108 (O_108,N_4986,N_4938);
and UO_109 (O_109,N_4943,N_4900);
or UO_110 (O_110,N_4945,N_4978);
or UO_111 (O_111,N_4977,N_4927);
nor UO_112 (O_112,N_4908,N_4974);
and UO_113 (O_113,N_4994,N_4949);
and UO_114 (O_114,N_4908,N_4921);
nor UO_115 (O_115,N_4917,N_4989);
nor UO_116 (O_116,N_4979,N_4975);
xor UO_117 (O_117,N_4977,N_4947);
nor UO_118 (O_118,N_4964,N_4994);
nor UO_119 (O_119,N_4973,N_4976);
nand UO_120 (O_120,N_4952,N_4930);
nor UO_121 (O_121,N_4976,N_4953);
and UO_122 (O_122,N_4956,N_4978);
nand UO_123 (O_123,N_4980,N_4950);
and UO_124 (O_124,N_4957,N_4954);
or UO_125 (O_125,N_4941,N_4912);
nand UO_126 (O_126,N_4973,N_4949);
nor UO_127 (O_127,N_4902,N_4959);
and UO_128 (O_128,N_4926,N_4923);
nor UO_129 (O_129,N_4916,N_4967);
xor UO_130 (O_130,N_4989,N_4997);
and UO_131 (O_131,N_4934,N_4920);
nand UO_132 (O_132,N_4939,N_4999);
and UO_133 (O_133,N_4965,N_4985);
nor UO_134 (O_134,N_4926,N_4968);
nor UO_135 (O_135,N_4931,N_4933);
nor UO_136 (O_136,N_4948,N_4934);
nor UO_137 (O_137,N_4920,N_4933);
and UO_138 (O_138,N_4988,N_4919);
nand UO_139 (O_139,N_4970,N_4953);
nand UO_140 (O_140,N_4981,N_4958);
nor UO_141 (O_141,N_4999,N_4970);
nand UO_142 (O_142,N_4933,N_4922);
nor UO_143 (O_143,N_4921,N_4965);
and UO_144 (O_144,N_4920,N_4987);
nand UO_145 (O_145,N_4904,N_4995);
nor UO_146 (O_146,N_4922,N_4911);
or UO_147 (O_147,N_4903,N_4973);
and UO_148 (O_148,N_4945,N_4975);
nor UO_149 (O_149,N_4990,N_4923);
nand UO_150 (O_150,N_4949,N_4928);
and UO_151 (O_151,N_4926,N_4918);
nor UO_152 (O_152,N_4983,N_4997);
nor UO_153 (O_153,N_4934,N_4966);
nand UO_154 (O_154,N_4930,N_4971);
or UO_155 (O_155,N_4901,N_4959);
nor UO_156 (O_156,N_4995,N_4911);
or UO_157 (O_157,N_4913,N_4973);
and UO_158 (O_158,N_4933,N_4964);
and UO_159 (O_159,N_4911,N_4985);
and UO_160 (O_160,N_4981,N_4918);
xnor UO_161 (O_161,N_4921,N_4968);
and UO_162 (O_162,N_4961,N_4928);
or UO_163 (O_163,N_4983,N_4977);
or UO_164 (O_164,N_4929,N_4905);
nand UO_165 (O_165,N_4916,N_4927);
or UO_166 (O_166,N_4987,N_4979);
nand UO_167 (O_167,N_4972,N_4989);
nor UO_168 (O_168,N_4913,N_4958);
and UO_169 (O_169,N_4934,N_4931);
nand UO_170 (O_170,N_4946,N_4926);
nor UO_171 (O_171,N_4955,N_4949);
or UO_172 (O_172,N_4956,N_4929);
and UO_173 (O_173,N_4989,N_4984);
and UO_174 (O_174,N_4952,N_4969);
and UO_175 (O_175,N_4962,N_4991);
and UO_176 (O_176,N_4961,N_4936);
and UO_177 (O_177,N_4977,N_4942);
nand UO_178 (O_178,N_4925,N_4929);
and UO_179 (O_179,N_4936,N_4937);
nor UO_180 (O_180,N_4955,N_4992);
or UO_181 (O_181,N_4984,N_4963);
nor UO_182 (O_182,N_4900,N_4916);
and UO_183 (O_183,N_4962,N_4967);
or UO_184 (O_184,N_4949,N_4904);
nor UO_185 (O_185,N_4931,N_4920);
nand UO_186 (O_186,N_4939,N_4950);
or UO_187 (O_187,N_4979,N_4941);
xnor UO_188 (O_188,N_4965,N_4937);
or UO_189 (O_189,N_4909,N_4913);
or UO_190 (O_190,N_4983,N_4902);
and UO_191 (O_191,N_4954,N_4918);
or UO_192 (O_192,N_4975,N_4967);
nor UO_193 (O_193,N_4970,N_4966);
or UO_194 (O_194,N_4944,N_4943);
nand UO_195 (O_195,N_4991,N_4928);
xor UO_196 (O_196,N_4949,N_4940);
nand UO_197 (O_197,N_4918,N_4940);
or UO_198 (O_198,N_4931,N_4990);
or UO_199 (O_199,N_4954,N_4936);
and UO_200 (O_200,N_4974,N_4980);
and UO_201 (O_201,N_4923,N_4905);
and UO_202 (O_202,N_4906,N_4929);
and UO_203 (O_203,N_4913,N_4904);
nor UO_204 (O_204,N_4916,N_4964);
nand UO_205 (O_205,N_4959,N_4948);
or UO_206 (O_206,N_4994,N_4944);
xor UO_207 (O_207,N_4920,N_4927);
and UO_208 (O_208,N_4916,N_4904);
and UO_209 (O_209,N_4966,N_4936);
or UO_210 (O_210,N_4999,N_4915);
nor UO_211 (O_211,N_4961,N_4971);
or UO_212 (O_212,N_4991,N_4935);
and UO_213 (O_213,N_4979,N_4983);
or UO_214 (O_214,N_4979,N_4962);
nor UO_215 (O_215,N_4931,N_4941);
and UO_216 (O_216,N_4917,N_4927);
or UO_217 (O_217,N_4995,N_4915);
nand UO_218 (O_218,N_4913,N_4947);
nand UO_219 (O_219,N_4919,N_4925);
nor UO_220 (O_220,N_4998,N_4966);
or UO_221 (O_221,N_4941,N_4937);
or UO_222 (O_222,N_4933,N_4974);
nand UO_223 (O_223,N_4995,N_4951);
nor UO_224 (O_224,N_4955,N_4909);
and UO_225 (O_225,N_4971,N_4984);
or UO_226 (O_226,N_4945,N_4911);
nand UO_227 (O_227,N_4931,N_4925);
and UO_228 (O_228,N_4905,N_4988);
nor UO_229 (O_229,N_4938,N_4993);
nand UO_230 (O_230,N_4941,N_4999);
nor UO_231 (O_231,N_4936,N_4958);
or UO_232 (O_232,N_4907,N_4965);
or UO_233 (O_233,N_4994,N_4983);
or UO_234 (O_234,N_4986,N_4943);
and UO_235 (O_235,N_4900,N_4961);
nor UO_236 (O_236,N_4982,N_4911);
nor UO_237 (O_237,N_4935,N_4950);
or UO_238 (O_238,N_4919,N_4997);
or UO_239 (O_239,N_4915,N_4937);
nor UO_240 (O_240,N_4980,N_4949);
nor UO_241 (O_241,N_4978,N_4905);
or UO_242 (O_242,N_4935,N_4941);
nor UO_243 (O_243,N_4942,N_4987);
or UO_244 (O_244,N_4940,N_4931);
or UO_245 (O_245,N_4970,N_4994);
or UO_246 (O_246,N_4989,N_4947);
nand UO_247 (O_247,N_4976,N_4948);
or UO_248 (O_248,N_4981,N_4943);
nor UO_249 (O_249,N_4910,N_4988);
nor UO_250 (O_250,N_4901,N_4956);
nor UO_251 (O_251,N_4984,N_4958);
and UO_252 (O_252,N_4965,N_4976);
or UO_253 (O_253,N_4949,N_4974);
nand UO_254 (O_254,N_4986,N_4914);
or UO_255 (O_255,N_4919,N_4907);
nor UO_256 (O_256,N_4951,N_4968);
nand UO_257 (O_257,N_4993,N_4997);
nand UO_258 (O_258,N_4904,N_4922);
or UO_259 (O_259,N_4955,N_4994);
xor UO_260 (O_260,N_4988,N_4994);
or UO_261 (O_261,N_4901,N_4979);
and UO_262 (O_262,N_4947,N_4934);
or UO_263 (O_263,N_4934,N_4983);
nand UO_264 (O_264,N_4945,N_4993);
xor UO_265 (O_265,N_4989,N_4980);
or UO_266 (O_266,N_4960,N_4916);
nor UO_267 (O_267,N_4990,N_4991);
nor UO_268 (O_268,N_4961,N_4956);
and UO_269 (O_269,N_4980,N_4904);
or UO_270 (O_270,N_4909,N_4933);
and UO_271 (O_271,N_4968,N_4994);
nand UO_272 (O_272,N_4976,N_4950);
or UO_273 (O_273,N_4962,N_4996);
and UO_274 (O_274,N_4912,N_4900);
nand UO_275 (O_275,N_4987,N_4934);
nor UO_276 (O_276,N_4944,N_4950);
nand UO_277 (O_277,N_4976,N_4931);
and UO_278 (O_278,N_4986,N_4961);
and UO_279 (O_279,N_4906,N_4935);
nor UO_280 (O_280,N_4993,N_4934);
xnor UO_281 (O_281,N_4990,N_4941);
xor UO_282 (O_282,N_4908,N_4990);
and UO_283 (O_283,N_4937,N_4966);
or UO_284 (O_284,N_4975,N_4993);
or UO_285 (O_285,N_4922,N_4948);
and UO_286 (O_286,N_4955,N_4914);
and UO_287 (O_287,N_4985,N_4954);
and UO_288 (O_288,N_4927,N_4929);
nand UO_289 (O_289,N_4920,N_4906);
nor UO_290 (O_290,N_4933,N_4934);
nor UO_291 (O_291,N_4977,N_4999);
and UO_292 (O_292,N_4979,N_4982);
nand UO_293 (O_293,N_4987,N_4913);
nor UO_294 (O_294,N_4996,N_4956);
and UO_295 (O_295,N_4992,N_4998);
nand UO_296 (O_296,N_4921,N_4981);
nor UO_297 (O_297,N_4911,N_4994);
or UO_298 (O_298,N_4991,N_4918);
nor UO_299 (O_299,N_4946,N_4913);
and UO_300 (O_300,N_4952,N_4932);
nor UO_301 (O_301,N_4989,N_4946);
and UO_302 (O_302,N_4966,N_4959);
or UO_303 (O_303,N_4956,N_4977);
nand UO_304 (O_304,N_4947,N_4946);
xnor UO_305 (O_305,N_4980,N_4935);
or UO_306 (O_306,N_4901,N_4902);
nor UO_307 (O_307,N_4996,N_4926);
nand UO_308 (O_308,N_4966,N_4972);
nand UO_309 (O_309,N_4903,N_4962);
nor UO_310 (O_310,N_4994,N_4907);
nor UO_311 (O_311,N_4945,N_4955);
or UO_312 (O_312,N_4910,N_4975);
or UO_313 (O_313,N_4907,N_4925);
and UO_314 (O_314,N_4964,N_4902);
nor UO_315 (O_315,N_4976,N_4916);
and UO_316 (O_316,N_4926,N_4983);
or UO_317 (O_317,N_4968,N_4957);
nor UO_318 (O_318,N_4903,N_4961);
nand UO_319 (O_319,N_4958,N_4921);
and UO_320 (O_320,N_4911,N_4944);
nor UO_321 (O_321,N_4953,N_4938);
nor UO_322 (O_322,N_4969,N_4942);
and UO_323 (O_323,N_4912,N_4948);
or UO_324 (O_324,N_4935,N_4924);
or UO_325 (O_325,N_4936,N_4969);
and UO_326 (O_326,N_4937,N_4921);
and UO_327 (O_327,N_4958,N_4973);
or UO_328 (O_328,N_4982,N_4966);
or UO_329 (O_329,N_4919,N_4924);
and UO_330 (O_330,N_4928,N_4942);
nor UO_331 (O_331,N_4918,N_4935);
xnor UO_332 (O_332,N_4916,N_4931);
or UO_333 (O_333,N_4927,N_4905);
and UO_334 (O_334,N_4908,N_4983);
nand UO_335 (O_335,N_4921,N_4962);
nand UO_336 (O_336,N_4967,N_4955);
and UO_337 (O_337,N_4949,N_4919);
nor UO_338 (O_338,N_4997,N_4908);
nor UO_339 (O_339,N_4974,N_4981);
nand UO_340 (O_340,N_4930,N_4920);
nand UO_341 (O_341,N_4965,N_4961);
nand UO_342 (O_342,N_4996,N_4988);
and UO_343 (O_343,N_4916,N_4989);
and UO_344 (O_344,N_4918,N_4979);
or UO_345 (O_345,N_4996,N_4905);
and UO_346 (O_346,N_4992,N_4940);
nor UO_347 (O_347,N_4999,N_4971);
or UO_348 (O_348,N_4984,N_4920);
nand UO_349 (O_349,N_4986,N_4998);
nor UO_350 (O_350,N_4972,N_4938);
nand UO_351 (O_351,N_4998,N_4977);
and UO_352 (O_352,N_4929,N_4970);
nand UO_353 (O_353,N_4902,N_4954);
and UO_354 (O_354,N_4989,N_4970);
nand UO_355 (O_355,N_4905,N_4926);
nand UO_356 (O_356,N_4930,N_4961);
or UO_357 (O_357,N_4942,N_4964);
or UO_358 (O_358,N_4985,N_4966);
or UO_359 (O_359,N_4987,N_4909);
or UO_360 (O_360,N_4962,N_4928);
xor UO_361 (O_361,N_4952,N_4980);
or UO_362 (O_362,N_4978,N_4913);
nand UO_363 (O_363,N_4930,N_4902);
or UO_364 (O_364,N_4951,N_4930);
nor UO_365 (O_365,N_4955,N_4939);
or UO_366 (O_366,N_4987,N_4921);
nand UO_367 (O_367,N_4905,N_4989);
xor UO_368 (O_368,N_4998,N_4979);
or UO_369 (O_369,N_4949,N_4932);
nand UO_370 (O_370,N_4998,N_4970);
or UO_371 (O_371,N_4915,N_4926);
nor UO_372 (O_372,N_4946,N_4962);
or UO_373 (O_373,N_4915,N_4942);
nand UO_374 (O_374,N_4930,N_4918);
nor UO_375 (O_375,N_4925,N_4986);
nor UO_376 (O_376,N_4973,N_4924);
nand UO_377 (O_377,N_4958,N_4908);
nor UO_378 (O_378,N_4989,N_4990);
or UO_379 (O_379,N_4973,N_4983);
and UO_380 (O_380,N_4931,N_4988);
nor UO_381 (O_381,N_4955,N_4981);
nor UO_382 (O_382,N_4906,N_4957);
or UO_383 (O_383,N_4952,N_4971);
and UO_384 (O_384,N_4902,N_4989);
nand UO_385 (O_385,N_4996,N_4974);
nand UO_386 (O_386,N_4980,N_4936);
or UO_387 (O_387,N_4942,N_4930);
or UO_388 (O_388,N_4971,N_4900);
or UO_389 (O_389,N_4937,N_4913);
or UO_390 (O_390,N_4914,N_4959);
or UO_391 (O_391,N_4968,N_4910);
or UO_392 (O_392,N_4989,N_4981);
or UO_393 (O_393,N_4925,N_4992);
or UO_394 (O_394,N_4943,N_4983);
nor UO_395 (O_395,N_4931,N_4972);
or UO_396 (O_396,N_4998,N_4942);
nor UO_397 (O_397,N_4966,N_4987);
or UO_398 (O_398,N_4930,N_4933);
nand UO_399 (O_399,N_4967,N_4906);
nand UO_400 (O_400,N_4958,N_4950);
nor UO_401 (O_401,N_4980,N_4993);
nand UO_402 (O_402,N_4960,N_4953);
nor UO_403 (O_403,N_4913,N_4967);
nand UO_404 (O_404,N_4926,N_4935);
and UO_405 (O_405,N_4930,N_4985);
and UO_406 (O_406,N_4907,N_4910);
and UO_407 (O_407,N_4963,N_4939);
or UO_408 (O_408,N_4993,N_4952);
or UO_409 (O_409,N_4924,N_4996);
or UO_410 (O_410,N_4933,N_4963);
nor UO_411 (O_411,N_4916,N_4918);
or UO_412 (O_412,N_4975,N_4962);
and UO_413 (O_413,N_4995,N_4960);
or UO_414 (O_414,N_4959,N_4977);
xnor UO_415 (O_415,N_4927,N_4973);
nand UO_416 (O_416,N_4961,N_4996);
and UO_417 (O_417,N_4926,N_4965);
nor UO_418 (O_418,N_4975,N_4966);
nor UO_419 (O_419,N_4904,N_4999);
nand UO_420 (O_420,N_4964,N_4921);
nand UO_421 (O_421,N_4951,N_4935);
nand UO_422 (O_422,N_4903,N_4970);
nor UO_423 (O_423,N_4975,N_4919);
and UO_424 (O_424,N_4932,N_4928);
or UO_425 (O_425,N_4969,N_4902);
nand UO_426 (O_426,N_4902,N_4956);
nor UO_427 (O_427,N_4954,N_4988);
and UO_428 (O_428,N_4973,N_4932);
or UO_429 (O_429,N_4930,N_4965);
nor UO_430 (O_430,N_4956,N_4906);
and UO_431 (O_431,N_4934,N_4992);
or UO_432 (O_432,N_4952,N_4908);
and UO_433 (O_433,N_4909,N_4906);
xor UO_434 (O_434,N_4970,N_4963);
and UO_435 (O_435,N_4906,N_4992);
and UO_436 (O_436,N_4974,N_4959);
nor UO_437 (O_437,N_4969,N_4923);
or UO_438 (O_438,N_4939,N_4936);
nand UO_439 (O_439,N_4957,N_4928);
nor UO_440 (O_440,N_4999,N_4967);
or UO_441 (O_441,N_4923,N_4938);
nand UO_442 (O_442,N_4935,N_4983);
nand UO_443 (O_443,N_4959,N_4985);
xnor UO_444 (O_444,N_4959,N_4961);
nand UO_445 (O_445,N_4983,N_4970);
and UO_446 (O_446,N_4950,N_4932);
or UO_447 (O_447,N_4925,N_4995);
nand UO_448 (O_448,N_4931,N_4901);
nor UO_449 (O_449,N_4926,N_4974);
nor UO_450 (O_450,N_4904,N_4997);
nor UO_451 (O_451,N_4907,N_4909);
nor UO_452 (O_452,N_4981,N_4987);
nor UO_453 (O_453,N_4973,N_4935);
nand UO_454 (O_454,N_4911,N_4932);
or UO_455 (O_455,N_4960,N_4950);
and UO_456 (O_456,N_4932,N_4967);
or UO_457 (O_457,N_4984,N_4951);
nor UO_458 (O_458,N_4903,N_4921);
nor UO_459 (O_459,N_4997,N_4951);
nand UO_460 (O_460,N_4942,N_4996);
nand UO_461 (O_461,N_4930,N_4909);
nand UO_462 (O_462,N_4978,N_4927);
nand UO_463 (O_463,N_4919,N_4916);
and UO_464 (O_464,N_4936,N_4947);
or UO_465 (O_465,N_4904,N_4941);
or UO_466 (O_466,N_4903,N_4933);
nand UO_467 (O_467,N_4971,N_4989);
and UO_468 (O_468,N_4907,N_4976);
and UO_469 (O_469,N_4909,N_4924);
nand UO_470 (O_470,N_4959,N_4952);
nand UO_471 (O_471,N_4931,N_4935);
and UO_472 (O_472,N_4904,N_4959);
and UO_473 (O_473,N_4907,N_4972);
or UO_474 (O_474,N_4906,N_4926);
nand UO_475 (O_475,N_4908,N_4957);
and UO_476 (O_476,N_4933,N_4913);
nor UO_477 (O_477,N_4942,N_4947);
and UO_478 (O_478,N_4906,N_4918);
nand UO_479 (O_479,N_4939,N_4956);
and UO_480 (O_480,N_4973,N_4972);
and UO_481 (O_481,N_4973,N_4963);
or UO_482 (O_482,N_4904,N_4945);
nor UO_483 (O_483,N_4932,N_4995);
nor UO_484 (O_484,N_4972,N_4915);
nor UO_485 (O_485,N_4922,N_4943);
nor UO_486 (O_486,N_4907,N_4989);
nand UO_487 (O_487,N_4960,N_4904);
nand UO_488 (O_488,N_4995,N_4961);
nor UO_489 (O_489,N_4998,N_4994);
and UO_490 (O_490,N_4998,N_4980);
xor UO_491 (O_491,N_4959,N_4957);
or UO_492 (O_492,N_4948,N_4957);
and UO_493 (O_493,N_4918,N_4939);
or UO_494 (O_494,N_4906,N_4936);
nor UO_495 (O_495,N_4991,N_4915);
nor UO_496 (O_496,N_4966,N_4906);
or UO_497 (O_497,N_4950,N_4948);
nand UO_498 (O_498,N_4925,N_4963);
and UO_499 (O_499,N_4953,N_4926);
or UO_500 (O_500,N_4965,N_4952);
nand UO_501 (O_501,N_4959,N_4949);
nor UO_502 (O_502,N_4957,N_4900);
nor UO_503 (O_503,N_4912,N_4981);
xor UO_504 (O_504,N_4968,N_4915);
and UO_505 (O_505,N_4965,N_4986);
or UO_506 (O_506,N_4944,N_4988);
nand UO_507 (O_507,N_4911,N_4964);
nor UO_508 (O_508,N_4945,N_4947);
or UO_509 (O_509,N_4988,N_4985);
nor UO_510 (O_510,N_4957,N_4973);
nand UO_511 (O_511,N_4950,N_4938);
nand UO_512 (O_512,N_4992,N_4911);
nand UO_513 (O_513,N_4906,N_4916);
nor UO_514 (O_514,N_4958,N_4938);
nor UO_515 (O_515,N_4905,N_4919);
nor UO_516 (O_516,N_4988,N_4981);
nor UO_517 (O_517,N_4942,N_4939);
nor UO_518 (O_518,N_4914,N_4934);
or UO_519 (O_519,N_4991,N_4964);
nor UO_520 (O_520,N_4960,N_4926);
or UO_521 (O_521,N_4970,N_4975);
nand UO_522 (O_522,N_4955,N_4956);
or UO_523 (O_523,N_4994,N_4986);
or UO_524 (O_524,N_4906,N_4924);
or UO_525 (O_525,N_4929,N_4961);
nor UO_526 (O_526,N_4969,N_4981);
or UO_527 (O_527,N_4990,N_4948);
or UO_528 (O_528,N_4908,N_4959);
or UO_529 (O_529,N_4937,N_4907);
nand UO_530 (O_530,N_4957,N_4977);
nor UO_531 (O_531,N_4922,N_4983);
nor UO_532 (O_532,N_4964,N_4993);
nand UO_533 (O_533,N_4984,N_4927);
nand UO_534 (O_534,N_4917,N_4921);
nand UO_535 (O_535,N_4988,N_4979);
nand UO_536 (O_536,N_4974,N_4992);
nor UO_537 (O_537,N_4996,N_4918);
nand UO_538 (O_538,N_4978,N_4998);
or UO_539 (O_539,N_4927,N_4949);
nand UO_540 (O_540,N_4912,N_4903);
and UO_541 (O_541,N_4905,N_4979);
nor UO_542 (O_542,N_4971,N_4934);
nand UO_543 (O_543,N_4949,N_4992);
nor UO_544 (O_544,N_4974,N_4928);
and UO_545 (O_545,N_4947,N_4998);
or UO_546 (O_546,N_4933,N_4942);
or UO_547 (O_547,N_4927,N_4901);
nand UO_548 (O_548,N_4903,N_4972);
nor UO_549 (O_549,N_4971,N_4972);
nor UO_550 (O_550,N_4962,N_4900);
and UO_551 (O_551,N_4999,N_4990);
nand UO_552 (O_552,N_4927,N_4960);
nor UO_553 (O_553,N_4950,N_4982);
and UO_554 (O_554,N_4936,N_4907);
and UO_555 (O_555,N_4990,N_4937);
nor UO_556 (O_556,N_4960,N_4913);
or UO_557 (O_557,N_4999,N_4927);
nand UO_558 (O_558,N_4984,N_4923);
nor UO_559 (O_559,N_4961,N_4922);
or UO_560 (O_560,N_4917,N_4935);
and UO_561 (O_561,N_4982,N_4957);
or UO_562 (O_562,N_4924,N_4972);
and UO_563 (O_563,N_4959,N_4939);
or UO_564 (O_564,N_4996,N_4953);
or UO_565 (O_565,N_4999,N_4925);
xnor UO_566 (O_566,N_4911,N_4908);
nand UO_567 (O_567,N_4956,N_4988);
nand UO_568 (O_568,N_4967,N_4942);
nor UO_569 (O_569,N_4968,N_4903);
nor UO_570 (O_570,N_4932,N_4990);
or UO_571 (O_571,N_4974,N_4967);
nor UO_572 (O_572,N_4905,N_4982);
and UO_573 (O_573,N_4905,N_4947);
nand UO_574 (O_574,N_4966,N_4917);
nand UO_575 (O_575,N_4974,N_4923);
and UO_576 (O_576,N_4960,N_4986);
nor UO_577 (O_577,N_4919,N_4994);
nor UO_578 (O_578,N_4909,N_4927);
nor UO_579 (O_579,N_4931,N_4982);
and UO_580 (O_580,N_4984,N_4996);
nor UO_581 (O_581,N_4962,N_4971);
and UO_582 (O_582,N_4957,N_4980);
nor UO_583 (O_583,N_4995,N_4956);
or UO_584 (O_584,N_4998,N_4972);
nor UO_585 (O_585,N_4910,N_4976);
nor UO_586 (O_586,N_4936,N_4992);
and UO_587 (O_587,N_4904,N_4989);
or UO_588 (O_588,N_4966,N_4944);
and UO_589 (O_589,N_4909,N_4931);
nand UO_590 (O_590,N_4972,N_4912);
or UO_591 (O_591,N_4978,N_4900);
nor UO_592 (O_592,N_4998,N_4922);
nand UO_593 (O_593,N_4906,N_4917);
or UO_594 (O_594,N_4943,N_4976);
nand UO_595 (O_595,N_4991,N_4929);
or UO_596 (O_596,N_4927,N_4948);
or UO_597 (O_597,N_4941,N_4960);
and UO_598 (O_598,N_4919,N_4951);
nand UO_599 (O_599,N_4907,N_4970);
or UO_600 (O_600,N_4905,N_4970);
nor UO_601 (O_601,N_4901,N_4967);
xnor UO_602 (O_602,N_4915,N_4979);
and UO_603 (O_603,N_4922,N_4945);
nor UO_604 (O_604,N_4990,N_4912);
nor UO_605 (O_605,N_4999,N_4929);
nand UO_606 (O_606,N_4903,N_4910);
and UO_607 (O_607,N_4989,N_4908);
or UO_608 (O_608,N_4924,N_4952);
or UO_609 (O_609,N_4972,N_4993);
and UO_610 (O_610,N_4918,N_4900);
nor UO_611 (O_611,N_4920,N_4978);
and UO_612 (O_612,N_4950,N_4922);
and UO_613 (O_613,N_4945,N_4949);
nor UO_614 (O_614,N_4909,N_4996);
and UO_615 (O_615,N_4954,N_4943);
nor UO_616 (O_616,N_4909,N_4965);
or UO_617 (O_617,N_4997,N_4928);
or UO_618 (O_618,N_4932,N_4918);
and UO_619 (O_619,N_4985,N_4931);
and UO_620 (O_620,N_4941,N_4962);
nand UO_621 (O_621,N_4907,N_4973);
nand UO_622 (O_622,N_4998,N_4940);
nor UO_623 (O_623,N_4964,N_4987);
nand UO_624 (O_624,N_4967,N_4924);
nor UO_625 (O_625,N_4941,N_4940);
nor UO_626 (O_626,N_4978,N_4974);
and UO_627 (O_627,N_4969,N_4944);
nand UO_628 (O_628,N_4907,N_4991);
nor UO_629 (O_629,N_4919,N_4937);
and UO_630 (O_630,N_4985,N_4939);
nand UO_631 (O_631,N_4953,N_4981);
or UO_632 (O_632,N_4915,N_4992);
and UO_633 (O_633,N_4925,N_4989);
xnor UO_634 (O_634,N_4902,N_4921);
or UO_635 (O_635,N_4990,N_4997);
and UO_636 (O_636,N_4954,N_4948);
and UO_637 (O_637,N_4900,N_4977);
or UO_638 (O_638,N_4905,N_4976);
and UO_639 (O_639,N_4934,N_4989);
nor UO_640 (O_640,N_4961,N_4901);
nand UO_641 (O_641,N_4947,N_4974);
or UO_642 (O_642,N_4939,N_4922);
nand UO_643 (O_643,N_4918,N_4990);
and UO_644 (O_644,N_4936,N_4964);
and UO_645 (O_645,N_4971,N_4901);
nand UO_646 (O_646,N_4976,N_4968);
and UO_647 (O_647,N_4997,N_4974);
or UO_648 (O_648,N_4971,N_4979);
and UO_649 (O_649,N_4981,N_4939);
and UO_650 (O_650,N_4979,N_4999);
nor UO_651 (O_651,N_4948,N_4923);
and UO_652 (O_652,N_4925,N_4900);
and UO_653 (O_653,N_4981,N_4961);
nand UO_654 (O_654,N_4914,N_4992);
nand UO_655 (O_655,N_4922,N_4946);
or UO_656 (O_656,N_4999,N_4966);
nand UO_657 (O_657,N_4993,N_4989);
nor UO_658 (O_658,N_4983,N_4928);
nand UO_659 (O_659,N_4975,N_4943);
and UO_660 (O_660,N_4952,N_4961);
nor UO_661 (O_661,N_4988,N_4983);
nand UO_662 (O_662,N_4921,N_4915);
or UO_663 (O_663,N_4957,N_4952);
or UO_664 (O_664,N_4920,N_4982);
nor UO_665 (O_665,N_4971,N_4946);
nor UO_666 (O_666,N_4954,N_4910);
and UO_667 (O_667,N_4905,N_4902);
and UO_668 (O_668,N_4949,N_4987);
nand UO_669 (O_669,N_4903,N_4925);
or UO_670 (O_670,N_4950,N_4988);
nor UO_671 (O_671,N_4952,N_4995);
nand UO_672 (O_672,N_4995,N_4971);
nand UO_673 (O_673,N_4980,N_4996);
nand UO_674 (O_674,N_4910,N_4987);
nand UO_675 (O_675,N_4974,N_4956);
or UO_676 (O_676,N_4956,N_4921);
and UO_677 (O_677,N_4946,N_4935);
nor UO_678 (O_678,N_4941,N_4967);
or UO_679 (O_679,N_4900,N_4908);
nand UO_680 (O_680,N_4906,N_4908);
or UO_681 (O_681,N_4922,N_4980);
or UO_682 (O_682,N_4957,N_4981);
and UO_683 (O_683,N_4957,N_4913);
and UO_684 (O_684,N_4943,N_4903);
xnor UO_685 (O_685,N_4903,N_4965);
or UO_686 (O_686,N_4961,N_4932);
or UO_687 (O_687,N_4940,N_4969);
or UO_688 (O_688,N_4980,N_4945);
nor UO_689 (O_689,N_4925,N_4952);
nor UO_690 (O_690,N_4932,N_4936);
nor UO_691 (O_691,N_4937,N_4986);
and UO_692 (O_692,N_4987,N_4976);
nand UO_693 (O_693,N_4938,N_4930);
nand UO_694 (O_694,N_4947,N_4914);
or UO_695 (O_695,N_4947,N_4919);
or UO_696 (O_696,N_4937,N_4906);
or UO_697 (O_697,N_4940,N_4916);
or UO_698 (O_698,N_4964,N_4904);
nand UO_699 (O_699,N_4998,N_4927);
nor UO_700 (O_700,N_4995,N_4930);
and UO_701 (O_701,N_4977,N_4935);
nand UO_702 (O_702,N_4976,N_4983);
or UO_703 (O_703,N_4947,N_4930);
xnor UO_704 (O_704,N_4927,N_4915);
xor UO_705 (O_705,N_4922,N_4947);
nand UO_706 (O_706,N_4944,N_4917);
nor UO_707 (O_707,N_4922,N_4930);
nor UO_708 (O_708,N_4919,N_4914);
and UO_709 (O_709,N_4930,N_4967);
or UO_710 (O_710,N_4955,N_4952);
nor UO_711 (O_711,N_4944,N_4999);
and UO_712 (O_712,N_4914,N_4980);
or UO_713 (O_713,N_4925,N_4974);
or UO_714 (O_714,N_4945,N_4995);
xnor UO_715 (O_715,N_4990,N_4992);
nand UO_716 (O_716,N_4910,N_4935);
nand UO_717 (O_717,N_4973,N_4959);
xor UO_718 (O_718,N_4989,N_4957);
nand UO_719 (O_719,N_4981,N_4949);
nand UO_720 (O_720,N_4928,N_4985);
xor UO_721 (O_721,N_4975,N_4902);
xnor UO_722 (O_722,N_4999,N_4973);
and UO_723 (O_723,N_4934,N_4960);
and UO_724 (O_724,N_4917,N_4957);
nand UO_725 (O_725,N_4940,N_4961);
nor UO_726 (O_726,N_4991,N_4909);
or UO_727 (O_727,N_4908,N_4950);
and UO_728 (O_728,N_4937,N_4964);
nor UO_729 (O_729,N_4920,N_4962);
nand UO_730 (O_730,N_4916,N_4924);
and UO_731 (O_731,N_4960,N_4920);
or UO_732 (O_732,N_4982,N_4969);
nand UO_733 (O_733,N_4998,N_4916);
nand UO_734 (O_734,N_4970,N_4984);
or UO_735 (O_735,N_4927,N_4923);
nor UO_736 (O_736,N_4953,N_4954);
nand UO_737 (O_737,N_4909,N_4932);
nand UO_738 (O_738,N_4997,N_4991);
and UO_739 (O_739,N_4925,N_4927);
nand UO_740 (O_740,N_4978,N_4941);
nor UO_741 (O_741,N_4920,N_4916);
nand UO_742 (O_742,N_4971,N_4990);
or UO_743 (O_743,N_4920,N_4950);
or UO_744 (O_744,N_4969,N_4996);
nor UO_745 (O_745,N_4947,N_4975);
or UO_746 (O_746,N_4924,N_4923);
or UO_747 (O_747,N_4919,N_4960);
nor UO_748 (O_748,N_4972,N_4962);
or UO_749 (O_749,N_4959,N_4953);
or UO_750 (O_750,N_4993,N_4923);
nor UO_751 (O_751,N_4990,N_4900);
nand UO_752 (O_752,N_4992,N_4902);
nand UO_753 (O_753,N_4989,N_4987);
nor UO_754 (O_754,N_4942,N_4917);
and UO_755 (O_755,N_4950,N_4914);
nand UO_756 (O_756,N_4976,N_4937);
or UO_757 (O_757,N_4907,N_4911);
and UO_758 (O_758,N_4941,N_4998);
and UO_759 (O_759,N_4976,N_4959);
and UO_760 (O_760,N_4937,N_4922);
or UO_761 (O_761,N_4930,N_4973);
xor UO_762 (O_762,N_4945,N_4919);
nand UO_763 (O_763,N_4967,N_4969);
nor UO_764 (O_764,N_4954,N_4986);
nor UO_765 (O_765,N_4915,N_4946);
and UO_766 (O_766,N_4993,N_4995);
and UO_767 (O_767,N_4942,N_4994);
and UO_768 (O_768,N_4918,N_4978);
and UO_769 (O_769,N_4968,N_4956);
and UO_770 (O_770,N_4958,N_4988);
nand UO_771 (O_771,N_4989,N_4918);
and UO_772 (O_772,N_4958,N_4944);
nor UO_773 (O_773,N_4970,N_4937);
nor UO_774 (O_774,N_4940,N_4911);
nand UO_775 (O_775,N_4914,N_4999);
nor UO_776 (O_776,N_4997,N_4956);
nor UO_777 (O_777,N_4940,N_4924);
nor UO_778 (O_778,N_4960,N_4936);
nand UO_779 (O_779,N_4944,N_4970);
nand UO_780 (O_780,N_4998,N_4911);
or UO_781 (O_781,N_4905,N_4930);
or UO_782 (O_782,N_4941,N_4951);
and UO_783 (O_783,N_4906,N_4999);
nor UO_784 (O_784,N_4940,N_4903);
nand UO_785 (O_785,N_4904,N_4912);
xor UO_786 (O_786,N_4999,N_4980);
or UO_787 (O_787,N_4945,N_4902);
nor UO_788 (O_788,N_4939,N_4977);
and UO_789 (O_789,N_4905,N_4949);
or UO_790 (O_790,N_4966,N_4979);
xor UO_791 (O_791,N_4951,N_4932);
or UO_792 (O_792,N_4920,N_4948);
or UO_793 (O_793,N_4984,N_4979);
nand UO_794 (O_794,N_4936,N_4959);
or UO_795 (O_795,N_4983,N_4927);
nor UO_796 (O_796,N_4965,N_4953);
nor UO_797 (O_797,N_4923,N_4917);
and UO_798 (O_798,N_4933,N_4984);
nand UO_799 (O_799,N_4948,N_4984);
nor UO_800 (O_800,N_4996,N_4922);
nor UO_801 (O_801,N_4906,N_4950);
or UO_802 (O_802,N_4979,N_4989);
and UO_803 (O_803,N_4925,N_4982);
and UO_804 (O_804,N_4981,N_4998);
and UO_805 (O_805,N_4959,N_4931);
or UO_806 (O_806,N_4901,N_4925);
or UO_807 (O_807,N_4918,N_4904);
or UO_808 (O_808,N_4911,N_4910);
nand UO_809 (O_809,N_4995,N_4983);
and UO_810 (O_810,N_4998,N_4955);
nand UO_811 (O_811,N_4904,N_4969);
nor UO_812 (O_812,N_4989,N_4983);
nor UO_813 (O_813,N_4962,N_4955);
and UO_814 (O_814,N_4962,N_4951);
and UO_815 (O_815,N_4970,N_4938);
and UO_816 (O_816,N_4948,N_4998);
nor UO_817 (O_817,N_4983,N_4971);
nand UO_818 (O_818,N_4922,N_4991);
or UO_819 (O_819,N_4972,N_4951);
nand UO_820 (O_820,N_4986,N_4931);
nand UO_821 (O_821,N_4983,N_4993);
and UO_822 (O_822,N_4989,N_4965);
or UO_823 (O_823,N_4964,N_4968);
or UO_824 (O_824,N_4964,N_4913);
and UO_825 (O_825,N_4977,N_4905);
and UO_826 (O_826,N_4950,N_4924);
or UO_827 (O_827,N_4939,N_4988);
nand UO_828 (O_828,N_4938,N_4998);
xnor UO_829 (O_829,N_4908,N_4994);
and UO_830 (O_830,N_4909,N_4942);
nor UO_831 (O_831,N_4985,N_4924);
or UO_832 (O_832,N_4940,N_4930);
nor UO_833 (O_833,N_4967,N_4915);
or UO_834 (O_834,N_4973,N_4967);
nor UO_835 (O_835,N_4984,N_4956);
nor UO_836 (O_836,N_4913,N_4944);
and UO_837 (O_837,N_4991,N_4972);
or UO_838 (O_838,N_4910,N_4956);
nor UO_839 (O_839,N_4907,N_4926);
or UO_840 (O_840,N_4991,N_4936);
xor UO_841 (O_841,N_4982,N_4910);
nand UO_842 (O_842,N_4931,N_4915);
or UO_843 (O_843,N_4938,N_4999);
or UO_844 (O_844,N_4987,N_4927);
nor UO_845 (O_845,N_4934,N_4907);
xnor UO_846 (O_846,N_4942,N_4956);
nor UO_847 (O_847,N_4931,N_4997);
and UO_848 (O_848,N_4920,N_4971);
xor UO_849 (O_849,N_4986,N_4980);
or UO_850 (O_850,N_4977,N_4926);
nand UO_851 (O_851,N_4918,N_4919);
nand UO_852 (O_852,N_4923,N_4904);
nand UO_853 (O_853,N_4923,N_4918);
nand UO_854 (O_854,N_4968,N_4943);
nor UO_855 (O_855,N_4988,N_4959);
nor UO_856 (O_856,N_4958,N_4939);
and UO_857 (O_857,N_4919,N_4986);
nor UO_858 (O_858,N_4997,N_4937);
or UO_859 (O_859,N_4992,N_4978);
nand UO_860 (O_860,N_4913,N_4929);
or UO_861 (O_861,N_4965,N_4923);
or UO_862 (O_862,N_4982,N_4958);
and UO_863 (O_863,N_4963,N_4987);
nor UO_864 (O_864,N_4992,N_4968);
or UO_865 (O_865,N_4979,N_4961);
nand UO_866 (O_866,N_4903,N_4947);
or UO_867 (O_867,N_4904,N_4981);
nor UO_868 (O_868,N_4909,N_4995);
nor UO_869 (O_869,N_4980,N_4959);
nand UO_870 (O_870,N_4960,N_4999);
nor UO_871 (O_871,N_4923,N_4906);
nor UO_872 (O_872,N_4972,N_4982);
nor UO_873 (O_873,N_4990,N_4982);
and UO_874 (O_874,N_4959,N_4960);
nand UO_875 (O_875,N_4903,N_4984);
or UO_876 (O_876,N_4911,N_4933);
nand UO_877 (O_877,N_4993,N_4973);
or UO_878 (O_878,N_4913,N_4953);
and UO_879 (O_879,N_4995,N_4939);
and UO_880 (O_880,N_4902,N_4994);
nor UO_881 (O_881,N_4978,N_4962);
or UO_882 (O_882,N_4933,N_4969);
or UO_883 (O_883,N_4913,N_4910);
nor UO_884 (O_884,N_4918,N_4980);
or UO_885 (O_885,N_4905,N_4904);
nand UO_886 (O_886,N_4989,N_4969);
and UO_887 (O_887,N_4918,N_4947);
and UO_888 (O_888,N_4938,N_4926);
nor UO_889 (O_889,N_4956,N_4934);
nand UO_890 (O_890,N_4973,N_4970);
or UO_891 (O_891,N_4908,N_4962);
xor UO_892 (O_892,N_4922,N_4907);
xor UO_893 (O_893,N_4956,N_4969);
and UO_894 (O_894,N_4936,N_4903);
nor UO_895 (O_895,N_4989,N_4930);
nor UO_896 (O_896,N_4984,N_4998);
and UO_897 (O_897,N_4992,N_4922);
nand UO_898 (O_898,N_4906,N_4987);
and UO_899 (O_899,N_4936,N_4965);
or UO_900 (O_900,N_4939,N_4933);
or UO_901 (O_901,N_4932,N_4922);
nor UO_902 (O_902,N_4925,N_4978);
or UO_903 (O_903,N_4978,N_4932);
nor UO_904 (O_904,N_4987,N_4926);
or UO_905 (O_905,N_4974,N_4918);
or UO_906 (O_906,N_4949,N_4937);
nand UO_907 (O_907,N_4952,N_4920);
nor UO_908 (O_908,N_4992,N_4999);
and UO_909 (O_909,N_4908,N_4939);
or UO_910 (O_910,N_4928,N_4936);
or UO_911 (O_911,N_4957,N_4956);
and UO_912 (O_912,N_4955,N_4913);
nor UO_913 (O_913,N_4942,N_4952);
and UO_914 (O_914,N_4914,N_4917);
nor UO_915 (O_915,N_4971,N_4942);
or UO_916 (O_916,N_4986,N_4912);
and UO_917 (O_917,N_4944,N_4993);
nor UO_918 (O_918,N_4943,N_4974);
or UO_919 (O_919,N_4901,N_4978);
nor UO_920 (O_920,N_4972,N_4999);
and UO_921 (O_921,N_4981,N_4982);
nor UO_922 (O_922,N_4917,N_4955);
nor UO_923 (O_923,N_4935,N_4961);
and UO_924 (O_924,N_4939,N_4994);
or UO_925 (O_925,N_4932,N_4955);
nor UO_926 (O_926,N_4919,N_4929);
nor UO_927 (O_927,N_4926,N_4994);
or UO_928 (O_928,N_4924,N_4912);
or UO_929 (O_929,N_4921,N_4945);
nand UO_930 (O_930,N_4907,N_4962);
and UO_931 (O_931,N_4909,N_4977);
xnor UO_932 (O_932,N_4926,N_4961);
nor UO_933 (O_933,N_4959,N_4915);
nor UO_934 (O_934,N_4985,N_4943);
nor UO_935 (O_935,N_4990,N_4936);
and UO_936 (O_936,N_4992,N_4932);
nor UO_937 (O_937,N_4929,N_4995);
or UO_938 (O_938,N_4947,N_4929);
and UO_939 (O_939,N_4948,N_4900);
or UO_940 (O_940,N_4903,N_4914);
and UO_941 (O_941,N_4953,N_4972);
and UO_942 (O_942,N_4907,N_4908);
nand UO_943 (O_943,N_4936,N_4938);
and UO_944 (O_944,N_4944,N_4908);
xnor UO_945 (O_945,N_4936,N_4984);
nor UO_946 (O_946,N_4901,N_4949);
xor UO_947 (O_947,N_4972,N_4949);
xor UO_948 (O_948,N_4980,N_4909);
nor UO_949 (O_949,N_4900,N_4937);
and UO_950 (O_950,N_4943,N_4960);
nand UO_951 (O_951,N_4939,N_4954);
or UO_952 (O_952,N_4963,N_4991);
nand UO_953 (O_953,N_4929,N_4968);
xnor UO_954 (O_954,N_4925,N_4923);
nand UO_955 (O_955,N_4972,N_4919);
or UO_956 (O_956,N_4971,N_4948);
nor UO_957 (O_957,N_4901,N_4934);
or UO_958 (O_958,N_4961,N_4974);
and UO_959 (O_959,N_4930,N_4948);
and UO_960 (O_960,N_4901,N_4938);
or UO_961 (O_961,N_4976,N_4957);
or UO_962 (O_962,N_4980,N_4985);
nand UO_963 (O_963,N_4931,N_4927);
and UO_964 (O_964,N_4972,N_4910);
and UO_965 (O_965,N_4981,N_4967);
or UO_966 (O_966,N_4952,N_4906);
and UO_967 (O_967,N_4912,N_4982);
nand UO_968 (O_968,N_4919,N_4993);
and UO_969 (O_969,N_4961,N_4912);
or UO_970 (O_970,N_4929,N_4950);
nand UO_971 (O_971,N_4906,N_4959);
nand UO_972 (O_972,N_4936,N_4982);
or UO_973 (O_973,N_4988,N_4949);
and UO_974 (O_974,N_4956,N_4953);
nand UO_975 (O_975,N_4908,N_4985);
nor UO_976 (O_976,N_4949,N_4961);
or UO_977 (O_977,N_4988,N_4968);
and UO_978 (O_978,N_4904,N_4979);
and UO_979 (O_979,N_4905,N_4975);
nand UO_980 (O_980,N_4945,N_4987);
nor UO_981 (O_981,N_4995,N_4959);
nand UO_982 (O_982,N_4908,N_4902);
nor UO_983 (O_983,N_4974,N_4911);
and UO_984 (O_984,N_4926,N_4954);
nor UO_985 (O_985,N_4931,N_4958);
nor UO_986 (O_986,N_4915,N_4900);
nor UO_987 (O_987,N_4906,N_4944);
and UO_988 (O_988,N_4991,N_4959);
or UO_989 (O_989,N_4962,N_4976);
and UO_990 (O_990,N_4986,N_4946);
and UO_991 (O_991,N_4948,N_4967);
and UO_992 (O_992,N_4928,N_4970);
nor UO_993 (O_993,N_4979,N_4992);
nor UO_994 (O_994,N_4926,N_4970);
nand UO_995 (O_995,N_4902,N_4946);
or UO_996 (O_996,N_4989,N_4903);
nand UO_997 (O_997,N_4951,N_4945);
nor UO_998 (O_998,N_4905,N_4972);
nand UO_999 (O_999,N_4910,N_4965);
endmodule