module basic_1000_10000_1500_4_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_957,In_646);
or U1 (N_1,In_881,In_629);
nor U2 (N_2,In_870,In_27);
or U3 (N_3,In_645,In_638);
nand U4 (N_4,In_947,In_916);
or U5 (N_5,In_586,In_833);
nor U6 (N_6,In_852,In_404);
and U7 (N_7,In_501,In_329);
or U8 (N_8,In_22,In_878);
or U9 (N_9,In_68,In_677);
or U10 (N_10,In_1,In_908);
nor U11 (N_11,In_372,In_396);
or U12 (N_12,In_258,In_488);
and U13 (N_13,In_814,In_340);
nor U14 (N_14,In_699,In_477);
nor U15 (N_15,In_845,In_216);
and U16 (N_16,In_171,In_377);
nor U17 (N_17,In_652,In_331);
and U18 (N_18,In_587,In_619);
nand U19 (N_19,In_735,In_758);
and U20 (N_20,In_668,In_342);
or U21 (N_21,In_548,In_525);
or U22 (N_22,In_764,In_61);
and U23 (N_23,In_254,In_263);
and U24 (N_24,In_755,In_28);
xnor U25 (N_25,In_681,In_352);
nand U26 (N_26,In_598,In_973);
nand U27 (N_27,In_999,In_392);
nor U28 (N_28,In_489,In_439);
xnor U29 (N_29,In_937,In_235);
and U30 (N_30,In_534,In_760);
or U31 (N_31,In_268,In_911);
and U32 (N_32,In_286,In_820);
or U33 (N_33,In_12,In_389);
nand U34 (N_34,In_982,In_436);
and U35 (N_35,In_790,In_2);
or U36 (N_36,In_444,In_185);
xor U37 (N_37,In_669,In_513);
or U38 (N_38,In_615,In_219);
nand U39 (N_39,In_335,In_0);
xnor U40 (N_40,In_754,In_294);
and U41 (N_41,In_129,In_327);
nand U42 (N_42,In_38,In_529);
and U43 (N_43,In_97,In_133);
nor U44 (N_44,In_673,In_147);
and U45 (N_45,In_935,In_802);
nand U46 (N_46,In_332,In_927);
nand U47 (N_47,In_157,In_694);
and U48 (N_48,In_901,In_160);
nand U49 (N_49,In_320,In_19);
nor U50 (N_50,In_691,In_544);
xnor U51 (N_51,In_300,In_430);
nand U52 (N_52,In_960,In_549);
or U53 (N_53,In_307,In_302);
or U54 (N_54,In_648,In_791);
nand U55 (N_55,In_610,In_511);
or U56 (N_56,In_884,In_785);
nand U57 (N_57,In_596,In_528);
nand U58 (N_58,In_745,In_136);
and U59 (N_59,In_228,In_657);
nand U60 (N_60,In_486,In_653);
nand U61 (N_61,In_104,In_249);
and U62 (N_62,In_174,In_350);
nor U63 (N_63,In_551,In_631);
or U64 (N_64,In_153,In_364);
nand U65 (N_65,In_312,In_406);
or U66 (N_66,In_582,In_950);
or U67 (N_67,In_266,In_30);
and U68 (N_68,In_289,In_40);
or U69 (N_69,In_81,In_943);
nand U70 (N_70,In_48,In_236);
and U71 (N_71,In_162,In_39);
xor U72 (N_72,In_568,In_301);
or U73 (N_73,In_116,In_72);
nand U74 (N_74,In_799,In_209);
or U75 (N_75,In_401,In_290);
and U76 (N_76,In_376,In_445);
nand U77 (N_77,In_92,In_964);
or U78 (N_78,In_592,In_463);
nor U79 (N_79,In_283,In_435);
and U80 (N_80,In_491,In_590);
and U81 (N_81,In_930,In_409);
nand U82 (N_82,In_193,In_841);
nand U83 (N_83,In_580,In_484);
and U84 (N_84,In_780,In_732);
or U85 (N_85,In_736,In_541);
nor U86 (N_86,In_925,In_661);
xnor U87 (N_87,In_561,In_713);
and U88 (N_88,In_252,In_373);
nor U89 (N_89,In_80,In_88);
nor U90 (N_90,In_448,In_73);
and U91 (N_91,In_634,In_9);
nor U92 (N_92,In_784,In_163);
and U93 (N_93,In_966,In_811);
or U94 (N_94,In_569,In_468);
nand U95 (N_95,In_381,In_778);
or U96 (N_96,In_837,In_397);
or U97 (N_97,In_469,In_743);
nand U98 (N_98,In_860,In_853);
or U99 (N_99,In_206,In_494);
nand U100 (N_100,In_442,In_410);
xnor U101 (N_101,In_684,In_285);
nor U102 (N_102,In_261,In_42);
or U103 (N_103,In_667,In_959);
or U104 (N_104,In_623,In_708);
nor U105 (N_105,In_287,In_308);
or U106 (N_106,In_761,In_356);
and U107 (N_107,In_51,In_924);
or U108 (N_108,In_44,In_512);
and U109 (N_109,In_979,In_919);
nand U110 (N_110,In_433,In_992);
or U111 (N_111,In_946,In_208);
nand U112 (N_112,In_798,In_385);
or U113 (N_113,In_751,In_255);
xor U114 (N_114,In_744,In_282);
nand U115 (N_115,In_125,In_461);
nor U116 (N_116,In_59,In_917);
nand U117 (N_117,In_835,In_573);
and U118 (N_118,In_237,In_17);
and U119 (N_119,In_720,In_63);
or U120 (N_120,In_972,In_523);
nor U121 (N_121,In_807,In_326);
nand U122 (N_122,In_706,In_535);
and U123 (N_123,In_889,In_613);
and U124 (N_124,In_138,In_422);
nor U125 (N_125,In_666,In_557);
or U126 (N_126,In_462,In_159);
and U127 (N_127,In_981,In_990);
nor U128 (N_128,In_131,In_759);
nor U129 (N_129,In_82,In_909);
nand U130 (N_130,In_299,In_186);
xnor U131 (N_131,In_432,In_793);
nand U132 (N_132,In_274,In_29);
xnor U133 (N_133,In_812,In_188);
nor U134 (N_134,In_650,In_358);
or U135 (N_135,In_231,In_180);
or U136 (N_136,In_4,In_707);
nand U137 (N_137,In_284,In_750);
nor U138 (N_138,In_637,In_939);
and U139 (N_139,In_505,In_822);
and U140 (N_140,In_633,In_245);
xnor U141 (N_141,In_702,In_37);
nor U142 (N_142,In_656,In_337);
and U143 (N_143,In_387,In_612);
xor U144 (N_144,In_609,In_295);
nor U145 (N_145,In_602,In_627);
nand U146 (N_146,In_495,In_118);
or U147 (N_147,In_330,In_746);
and U148 (N_148,In_213,In_67);
nor U149 (N_149,In_108,In_933);
and U150 (N_150,In_408,In_374);
or U151 (N_151,In_310,In_278);
nor U152 (N_152,In_556,In_52);
and U153 (N_153,In_378,In_796);
or U154 (N_154,In_164,In_693);
and U155 (N_155,In_229,In_277);
nand U156 (N_156,In_844,In_265);
and U157 (N_157,In_168,In_687);
xor U158 (N_158,In_597,In_942);
and U159 (N_159,In_543,In_829);
nor U160 (N_160,In_975,In_210);
xor U161 (N_161,In_156,In_774);
nand U162 (N_162,In_905,In_124);
nand U163 (N_163,In_450,In_492);
and U164 (N_164,In_989,In_956);
nor U165 (N_165,In_487,In_453);
nor U166 (N_166,In_894,In_899);
and U167 (N_167,In_275,In_663);
or U168 (N_168,In_762,In_718);
nor U169 (N_169,In_731,In_660);
and U170 (N_170,In_10,In_234);
nor U171 (N_171,In_69,In_722);
or U172 (N_172,In_730,In_647);
nand U173 (N_173,In_649,In_578);
xor U174 (N_174,In_572,In_842);
and U175 (N_175,In_969,In_143);
nor U176 (N_176,In_898,In_194);
and U177 (N_177,In_620,In_338);
nor U178 (N_178,In_149,In_536);
nor U179 (N_179,In_665,In_483);
nor U180 (N_180,In_58,In_948);
or U181 (N_181,In_293,In_55);
and U182 (N_182,In_34,In_875);
nor U183 (N_183,In_3,In_757);
nor U184 (N_184,In_874,In_53);
nor U185 (N_185,In_426,In_414);
or U186 (N_186,In_742,In_184);
or U187 (N_187,In_144,In_922);
or U188 (N_188,In_111,In_542);
nor U189 (N_189,In_565,In_384);
xnor U190 (N_190,In_70,In_482);
and U191 (N_191,In_782,In_411);
and U192 (N_192,In_360,In_84);
and U193 (N_193,In_831,In_876);
nand U194 (N_194,In_716,In_574);
nand U195 (N_195,In_178,In_161);
nand U196 (N_196,In_388,In_695);
and U197 (N_197,In_768,In_246);
nand U198 (N_198,In_662,In_522);
nand U199 (N_199,In_719,In_165);
and U200 (N_200,In_527,In_242);
nand U201 (N_201,In_739,In_787);
nor U202 (N_202,In_303,In_365);
or U203 (N_203,In_298,In_955);
and U204 (N_204,In_56,In_704);
nor U205 (N_205,In_819,In_386);
xnor U206 (N_206,In_882,In_437);
nand U207 (N_207,In_983,In_747);
nand U208 (N_208,In_15,In_50);
or U209 (N_209,In_250,In_117);
nor U210 (N_210,In_963,In_204);
nand U211 (N_211,In_890,In_804);
nor U212 (N_212,In_714,In_741);
nor U213 (N_213,In_651,In_521);
or U214 (N_214,In_766,In_788);
nor U215 (N_215,In_577,In_325);
or U216 (N_216,In_106,In_509);
xnor U217 (N_217,In_251,In_517);
or U218 (N_218,In_836,In_697);
nand U219 (N_219,In_13,In_120);
and U220 (N_220,In_221,In_203);
and U221 (N_221,In_421,In_207);
nor U222 (N_222,In_336,In_135);
or U223 (N_223,In_628,In_317);
nor U224 (N_224,In_239,In_167);
or U225 (N_225,In_296,In_644);
and U226 (N_226,In_109,In_90);
nand U227 (N_227,In_570,In_398);
nor U228 (N_228,In_847,In_98);
nand U229 (N_229,In_481,In_929);
xnor U230 (N_230,In_407,In_451);
xnor U231 (N_231,In_686,In_247);
and U232 (N_232,In_480,In_65);
and U233 (N_233,In_233,In_457);
xnor U234 (N_234,In_458,In_191);
nand U235 (N_235,In_832,In_546);
nand U236 (N_236,In_363,In_794);
nand U237 (N_237,In_828,In_850);
nand U238 (N_238,In_446,In_608);
nand U239 (N_239,In_672,In_334);
nor U240 (N_240,In_846,In_532);
and U241 (N_241,In_78,In_139);
nand U242 (N_242,In_36,In_201);
and U243 (N_243,In_31,In_271);
and U244 (N_244,In_781,In_225);
and U245 (N_245,In_16,In_455);
or U246 (N_246,In_351,In_599);
or U247 (N_247,In_75,In_141);
nand U248 (N_248,In_197,In_253);
and U249 (N_249,In_826,In_825);
xnor U250 (N_250,In_626,In_641);
or U251 (N_251,In_539,In_506);
nand U252 (N_252,In_128,In_443);
and U253 (N_253,In_855,In_954);
nand U254 (N_254,In_906,In_962);
nor U255 (N_255,In_618,In_988);
and U256 (N_256,In_215,In_721);
or U257 (N_257,In_370,In_941);
nor U258 (N_258,In_926,In_395);
and U259 (N_259,In_914,In_83);
or U260 (N_260,In_823,In_617);
xnor U261 (N_261,In_915,In_493);
nor U262 (N_262,In_438,In_526);
or U263 (N_263,In_273,In_8);
nand U264 (N_264,In_447,In_47);
and U265 (N_265,In_238,In_767);
and U266 (N_266,In_622,In_974);
and U267 (N_267,In_636,In_607);
or U268 (N_268,In_728,In_211);
nor U269 (N_269,In_777,In_856);
nand U270 (N_270,In_464,In_471);
and U271 (N_271,In_579,In_770);
nor U272 (N_272,In_861,In_840);
xor U273 (N_273,In_918,In_545);
nand U274 (N_274,In_474,In_454);
or U275 (N_275,In_262,In_466);
and U276 (N_276,In_868,In_808);
nor U277 (N_277,In_357,In_934);
or U278 (N_278,In_353,In_400);
xnor U279 (N_279,In_816,In_476);
or U280 (N_280,In_858,In_997);
nor U281 (N_281,In_41,In_140);
nand U282 (N_282,In_859,In_187);
nand U283 (N_283,In_698,In_412);
nand U284 (N_284,In_394,In_86);
nor U285 (N_285,In_503,In_148);
or U286 (N_286,In_232,In_520);
and U287 (N_287,In_998,In_115);
nor U288 (N_288,In_643,In_102);
and U289 (N_289,In_260,In_897);
nand U290 (N_290,In_405,In_490);
or U291 (N_291,In_107,In_961);
and U292 (N_292,In_883,In_220);
or U293 (N_293,In_904,In_313);
or U294 (N_294,In_869,In_57);
nor U295 (N_295,In_729,In_560);
or U296 (N_296,In_383,In_676);
and U297 (N_297,In_256,In_459);
nand U298 (N_298,In_420,In_839);
nand U299 (N_299,In_813,In_817);
xnor U300 (N_300,In_671,In_49);
nand U301 (N_301,In_871,In_333);
and U302 (N_302,In_786,In_431);
nand U303 (N_303,In_257,In_967);
nor U304 (N_304,In_348,In_427);
nand U305 (N_305,In_413,In_391);
and U306 (N_306,In_126,In_753);
xor U307 (N_307,In_712,In_315);
xnor U308 (N_308,In_95,In_566);
nor U309 (N_309,In_775,In_524);
and U310 (N_310,In_33,In_272);
xnor U311 (N_311,In_715,In_563);
nand U312 (N_312,In_752,In_103);
nor U313 (N_313,In_584,In_809);
nor U314 (N_314,In_863,In_900);
or U315 (N_315,In_280,In_214);
and U316 (N_316,In_680,In_177);
nand U317 (N_317,In_339,In_43);
or U318 (N_318,In_485,In_46);
nand U319 (N_319,In_675,In_276);
or U320 (N_320,In_150,In_26);
nor U321 (N_321,In_267,In_738);
or U322 (N_322,In_259,In_71);
or U323 (N_323,In_99,In_949);
and U324 (N_324,In_601,In_984);
or U325 (N_325,In_472,In_769);
xor U326 (N_326,In_606,In_200);
nand U327 (N_327,In_182,In_328);
and U328 (N_328,In_604,In_18);
or U329 (N_329,In_311,In_585);
nor U330 (N_330,In_244,In_429);
and U331 (N_331,In_849,In_25);
nor U332 (N_332,In_815,In_371);
nand U333 (N_333,In_217,In_895);
and U334 (N_334,In_701,In_155);
and U335 (N_335,In_60,In_553);
xor U336 (N_336,In_418,In_230);
or U337 (N_337,In_576,In_940);
and U338 (N_338,In_519,In_611);
xor U339 (N_339,In_54,In_945);
and U340 (N_340,In_417,In_223);
nor U341 (N_341,In_345,In_733);
nor U342 (N_342,In_765,In_449);
or U343 (N_343,In_709,In_416);
nand U344 (N_344,In_688,In_690);
or U345 (N_345,In_803,In_625);
nand U346 (N_346,In_323,In_783);
or U347 (N_347,In_571,In_240);
and U348 (N_348,In_425,In_291);
and U349 (N_349,In_5,In_952);
and U350 (N_350,In_196,In_66);
or U351 (N_351,In_20,In_419);
xor U352 (N_352,In_362,In_62);
and U353 (N_353,In_564,In_862);
or U354 (N_354,In_297,In_314);
and U355 (N_355,In_91,In_896);
or U356 (N_356,In_540,In_470);
or U357 (N_357,In_772,In_976);
and U358 (N_358,In_591,In_114);
nand U359 (N_359,In_172,In_595);
and U360 (N_360,In_887,In_987);
or U361 (N_361,In_467,In_797);
or U362 (N_362,In_740,In_380);
or U363 (N_363,In_885,In_995);
or U364 (N_364,In_674,In_134);
and U365 (N_365,In_864,In_248);
or U366 (N_366,In_478,In_936);
xnor U367 (N_367,In_45,In_122);
or U368 (N_368,In_857,In_403);
nor U369 (N_369,In_367,In_879);
or U370 (N_370,In_100,In_994);
and U371 (N_371,In_834,In_85);
nand U372 (N_372,In_851,In_763);
nand U373 (N_373,In_269,In_792);
nand U374 (N_374,In_821,In_89);
and U375 (N_375,In_843,In_877);
nor U376 (N_376,In_205,In_175);
and U377 (N_377,In_723,In_77);
and U378 (N_378,In_324,In_496);
and U379 (N_379,In_192,In_169);
and U380 (N_380,In_375,In_771);
and U381 (N_381,In_827,In_605);
or U382 (N_382,In_304,In_390);
xnor U383 (N_383,In_944,In_359);
and U384 (N_384,In_190,In_530);
and U385 (N_385,In_913,In_552);
nand U386 (N_386,In_224,In_281);
and U387 (N_387,In_382,In_270);
and U388 (N_388,In_154,In_119);
and U389 (N_389,In_902,In_953);
and U390 (N_390,In_555,In_514);
or U391 (N_391,In_621,In_538);
xor U392 (N_392,In_212,In_399);
nand U393 (N_393,In_393,In_241);
xnor U394 (N_394,In_243,In_932);
nor U395 (N_395,In_11,In_977);
xnor U396 (N_396,In_655,In_931);
nand U397 (N_397,In_830,In_748);
nor U398 (N_398,In_891,In_951);
and U399 (N_399,In_344,In_309);
xnor U400 (N_400,In_498,In_880);
or U401 (N_401,In_146,In_642);
and U402 (N_402,In_428,In_810);
nor U403 (N_403,In_465,In_199);
nor U404 (N_404,In_773,In_776);
nand U405 (N_405,In_434,In_910);
nand U406 (N_406,In_112,In_756);
or U407 (N_407,In_630,In_635);
or U408 (N_408,In_94,In_292);
nand U409 (N_409,In_189,In_516);
nor U410 (N_410,In_554,In_379);
and U411 (N_411,In_24,In_152);
or U412 (N_412,In_993,In_537);
or U413 (N_413,In_550,In_179);
or U414 (N_414,In_920,In_64);
nor U415 (N_415,In_659,In_679);
nand U416 (N_416,In_508,In_978);
or U417 (N_417,In_479,In_137);
nor U418 (N_418,In_23,In_678);
nand U419 (N_419,In_907,In_21);
nand U420 (N_420,In_658,In_873);
or U421 (N_421,In_670,In_692);
or U422 (N_422,In_355,In_616);
or U423 (N_423,In_173,In_76);
xnor U424 (N_424,In_664,In_181);
and U425 (N_425,In_319,In_347);
and U426 (N_426,In_958,In_318);
nor U427 (N_427,In_306,In_639);
or U428 (N_428,In_504,In_113);
or U429 (N_429,In_725,In_921);
or U430 (N_430,In_806,In_288);
or U431 (N_431,In_575,In_886);
or U432 (N_432,In_6,In_888);
or U433 (N_433,In_101,In_183);
and U434 (N_434,In_166,In_198);
or U435 (N_435,In_562,In_264);
nand U436 (N_436,In_226,In_145);
or U437 (N_437,In_749,In_499);
or U438 (N_438,In_683,In_369);
nor U439 (N_439,In_158,In_14);
nand U440 (N_440,In_475,In_402);
or U441 (N_441,In_703,In_567);
nor U442 (N_442,In_700,In_581);
or U443 (N_443,In_971,In_600);
nor U444 (N_444,In_132,In_121);
or U445 (N_445,In_361,In_801);
nor U446 (N_446,In_473,In_170);
or U447 (N_447,In_603,In_717);
nand U448 (N_448,In_903,In_986);
and U449 (N_449,In_452,In_151);
and U450 (N_450,In_805,In_515);
nand U451 (N_451,In_74,In_510);
nand U452 (N_452,In_456,In_724);
nand U453 (N_453,In_980,In_867);
or U454 (N_454,In_93,In_354);
xnor U455 (N_455,In_865,In_368);
nor U456 (N_456,In_321,In_912);
nor U457 (N_457,In_866,In_779);
nor U458 (N_458,In_727,In_559);
and U459 (N_459,In_96,In_343);
or U460 (N_460,In_32,In_593);
and U461 (N_461,In_583,In_985);
xor U462 (N_462,In_654,In_497);
and U463 (N_463,In_35,In_531);
nand U464 (N_464,In_996,In_110);
and U465 (N_465,In_689,In_558);
and U466 (N_466,In_460,In_824);
nor U467 (N_467,In_279,In_624);
nand U468 (N_468,In_79,In_423);
xnor U469 (N_469,In_341,In_7);
or U470 (N_470,In_789,In_127);
nand U471 (N_471,In_854,In_227);
or U472 (N_472,In_441,In_589);
xor U473 (N_473,In_928,In_588);
or U474 (N_474,In_222,In_518);
and U475 (N_475,In_346,In_502);
nand U476 (N_476,In_632,In_130);
xnor U477 (N_477,In_970,In_737);
or U478 (N_478,In_872,In_968);
nand U479 (N_479,In_938,In_696);
or U480 (N_480,In_685,In_734);
and U481 (N_481,In_142,In_594);
nor U482 (N_482,In_682,In_848);
nor U483 (N_483,In_349,In_218);
nand U484 (N_484,In_176,In_533);
or U485 (N_485,In_500,In_711);
nor U486 (N_486,In_105,In_818);
or U487 (N_487,In_87,In_705);
nand U488 (N_488,In_800,In_710);
and U489 (N_489,In_838,In_965);
nand U490 (N_490,In_923,In_892);
or U491 (N_491,In_415,In_123);
nor U492 (N_492,In_424,In_893);
or U493 (N_493,In_305,In_366);
and U494 (N_494,In_195,In_507);
or U495 (N_495,In_795,In_991);
nand U496 (N_496,In_614,In_440);
or U497 (N_497,In_640,In_726);
nor U498 (N_498,In_547,In_202);
or U499 (N_499,In_316,In_322);
nor U500 (N_500,In_750,In_714);
nor U501 (N_501,In_634,In_988);
xnor U502 (N_502,In_448,In_26);
nand U503 (N_503,In_342,In_913);
nand U504 (N_504,In_695,In_896);
nor U505 (N_505,In_903,In_376);
nor U506 (N_506,In_357,In_957);
xnor U507 (N_507,In_362,In_871);
and U508 (N_508,In_63,In_537);
and U509 (N_509,In_806,In_257);
and U510 (N_510,In_750,In_997);
or U511 (N_511,In_337,In_764);
nor U512 (N_512,In_966,In_151);
nor U513 (N_513,In_99,In_495);
nor U514 (N_514,In_287,In_314);
and U515 (N_515,In_948,In_690);
nor U516 (N_516,In_139,In_510);
and U517 (N_517,In_304,In_604);
and U518 (N_518,In_774,In_319);
and U519 (N_519,In_681,In_874);
nor U520 (N_520,In_957,In_112);
or U521 (N_521,In_952,In_616);
and U522 (N_522,In_915,In_693);
xnor U523 (N_523,In_241,In_918);
and U524 (N_524,In_667,In_508);
xor U525 (N_525,In_13,In_144);
nor U526 (N_526,In_573,In_207);
or U527 (N_527,In_628,In_428);
or U528 (N_528,In_637,In_884);
nand U529 (N_529,In_166,In_407);
or U530 (N_530,In_303,In_858);
or U531 (N_531,In_365,In_575);
xnor U532 (N_532,In_229,In_115);
or U533 (N_533,In_761,In_420);
nand U534 (N_534,In_599,In_706);
nor U535 (N_535,In_477,In_862);
xnor U536 (N_536,In_921,In_650);
nand U537 (N_537,In_538,In_167);
and U538 (N_538,In_830,In_651);
and U539 (N_539,In_922,In_573);
or U540 (N_540,In_816,In_849);
nand U541 (N_541,In_992,In_236);
nand U542 (N_542,In_761,In_49);
nor U543 (N_543,In_406,In_828);
nand U544 (N_544,In_685,In_746);
or U545 (N_545,In_285,In_425);
nor U546 (N_546,In_584,In_275);
and U547 (N_547,In_777,In_631);
and U548 (N_548,In_49,In_314);
nor U549 (N_549,In_169,In_15);
and U550 (N_550,In_767,In_135);
nor U551 (N_551,In_308,In_18);
nor U552 (N_552,In_779,In_342);
and U553 (N_553,In_663,In_317);
or U554 (N_554,In_629,In_425);
nor U555 (N_555,In_801,In_123);
nor U556 (N_556,In_554,In_527);
nor U557 (N_557,In_239,In_421);
and U558 (N_558,In_284,In_476);
and U559 (N_559,In_491,In_519);
and U560 (N_560,In_719,In_72);
or U561 (N_561,In_593,In_685);
and U562 (N_562,In_708,In_840);
nor U563 (N_563,In_824,In_270);
or U564 (N_564,In_264,In_205);
or U565 (N_565,In_605,In_164);
nor U566 (N_566,In_344,In_885);
xor U567 (N_567,In_221,In_304);
and U568 (N_568,In_126,In_216);
or U569 (N_569,In_215,In_314);
and U570 (N_570,In_593,In_473);
and U571 (N_571,In_944,In_629);
nand U572 (N_572,In_929,In_515);
and U573 (N_573,In_639,In_186);
or U574 (N_574,In_378,In_969);
nand U575 (N_575,In_795,In_738);
nor U576 (N_576,In_258,In_445);
nand U577 (N_577,In_249,In_278);
nand U578 (N_578,In_509,In_259);
nor U579 (N_579,In_301,In_736);
nand U580 (N_580,In_486,In_441);
and U581 (N_581,In_666,In_821);
or U582 (N_582,In_380,In_707);
nand U583 (N_583,In_305,In_90);
nand U584 (N_584,In_962,In_958);
xor U585 (N_585,In_829,In_128);
xor U586 (N_586,In_395,In_604);
nor U587 (N_587,In_872,In_869);
and U588 (N_588,In_622,In_40);
or U589 (N_589,In_291,In_436);
nand U590 (N_590,In_461,In_579);
or U591 (N_591,In_674,In_368);
or U592 (N_592,In_618,In_262);
and U593 (N_593,In_600,In_924);
xor U594 (N_594,In_5,In_187);
nand U595 (N_595,In_122,In_824);
xnor U596 (N_596,In_56,In_302);
and U597 (N_597,In_23,In_133);
nor U598 (N_598,In_735,In_686);
nor U599 (N_599,In_939,In_116);
nand U600 (N_600,In_15,In_957);
and U601 (N_601,In_346,In_370);
or U602 (N_602,In_538,In_290);
nor U603 (N_603,In_802,In_900);
and U604 (N_604,In_865,In_132);
nand U605 (N_605,In_152,In_325);
and U606 (N_606,In_888,In_39);
or U607 (N_607,In_245,In_204);
nor U608 (N_608,In_809,In_806);
nand U609 (N_609,In_134,In_484);
xnor U610 (N_610,In_879,In_996);
nand U611 (N_611,In_134,In_630);
or U612 (N_612,In_681,In_314);
nor U613 (N_613,In_459,In_352);
nor U614 (N_614,In_658,In_553);
nor U615 (N_615,In_461,In_931);
nor U616 (N_616,In_419,In_302);
xnor U617 (N_617,In_400,In_956);
xor U618 (N_618,In_448,In_706);
nand U619 (N_619,In_350,In_240);
nand U620 (N_620,In_460,In_507);
nand U621 (N_621,In_963,In_289);
or U622 (N_622,In_542,In_987);
nand U623 (N_623,In_183,In_749);
xnor U624 (N_624,In_96,In_570);
or U625 (N_625,In_724,In_214);
and U626 (N_626,In_928,In_209);
nor U627 (N_627,In_287,In_322);
nand U628 (N_628,In_326,In_529);
and U629 (N_629,In_850,In_711);
nor U630 (N_630,In_572,In_110);
or U631 (N_631,In_753,In_927);
and U632 (N_632,In_882,In_550);
nor U633 (N_633,In_83,In_469);
nor U634 (N_634,In_879,In_954);
nor U635 (N_635,In_170,In_126);
or U636 (N_636,In_553,In_370);
xnor U637 (N_637,In_332,In_555);
or U638 (N_638,In_806,In_463);
nand U639 (N_639,In_791,In_723);
xor U640 (N_640,In_381,In_550);
nor U641 (N_641,In_917,In_93);
and U642 (N_642,In_79,In_990);
or U643 (N_643,In_648,In_592);
nor U644 (N_644,In_907,In_94);
and U645 (N_645,In_497,In_21);
and U646 (N_646,In_798,In_962);
and U647 (N_647,In_164,In_219);
nor U648 (N_648,In_723,In_44);
nor U649 (N_649,In_397,In_296);
nor U650 (N_650,In_486,In_564);
nand U651 (N_651,In_575,In_297);
xor U652 (N_652,In_389,In_832);
or U653 (N_653,In_838,In_991);
or U654 (N_654,In_554,In_125);
nand U655 (N_655,In_323,In_356);
xnor U656 (N_656,In_354,In_374);
or U657 (N_657,In_586,In_442);
or U658 (N_658,In_108,In_134);
and U659 (N_659,In_209,In_159);
nand U660 (N_660,In_623,In_926);
and U661 (N_661,In_571,In_280);
or U662 (N_662,In_417,In_714);
and U663 (N_663,In_184,In_270);
nand U664 (N_664,In_689,In_374);
or U665 (N_665,In_385,In_227);
nand U666 (N_666,In_423,In_408);
nand U667 (N_667,In_961,In_702);
xnor U668 (N_668,In_465,In_929);
nor U669 (N_669,In_318,In_531);
xor U670 (N_670,In_247,In_383);
nor U671 (N_671,In_218,In_296);
and U672 (N_672,In_300,In_979);
and U673 (N_673,In_609,In_866);
nand U674 (N_674,In_721,In_419);
or U675 (N_675,In_887,In_836);
or U676 (N_676,In_770,In_479);
and U677 (N_677,In_695,In_677);
and U678 (N_678,In_691,In_593);
nor U679 (N_679,In_396,In_851);
or U680 (N_680,In_792,In_796);
nor U681 (N_681,In_588,In_346);
and U682 (N_682,In_8,In_356);
or U683 (N_683,In_127,In_126);
nor U684 (N_684,In_638,In_364);
nor U685 (N_685,In_101,In_747);
nand U686 (N_686,In_96,In_476);
xnor U687 (N_687,In_311,In_115);
nor U688 (N_688,In_644,In_196);
or U689 (N_689,In_276,In_844);
or U690 (N_690,In_853,In_336);
nor U691 (N_691,In_300,In_80);
and U692 (N_692,In_655,In_779);
xnor U693 (N_693,In_55,In_182);
nand U694 (N_694,In_290,In_607);
or U695 (N_695,In_215,In_503);
xor U696 (N_696,In_754,In_344);
nor U697 (N_697,In_447,In_158);
nor U698 (N_698,In_765,In_23);
and U699 (N_699,In_393,In_495);
nor U700 (N_700,In_94,In_970);
nand U701 (N_701,In_578,In_542);
nand U702 (N_702,In_41,In_665);
or U703 (N_703,In_504,In_672);
and U704 (N_704,In_739,In_548);
or U705 (N_705,In_522,In_839);
nor U706 (N_706,In_959,In_344);
nand U707 (N_707,In_98,In_57);
nand U708 (N_708,In_480,In_246);
nand U709 (N_709,In_784,In_67);
xor U710 (N_710,In_888,In_219);
and U711 (N_711,In_541,In_733);
nand U712 (N_712,In_608,In_184);
xor U713 (N_713,In_71,In_202);
xor U714 (N_714,In_86,In_441);
or U715 (N_715,In_343,In_203);
or U716 (N_716,In_916,In_949);
and U717 (N_717,In_787,In_681);
or U718 (N_718,In_61,In_662);
and U719 (N_719,In_523,In_401);
xnor U720 (N_720,In_914,In_904);
nor U721 (N_721,In_992,In_257);
nor U722 (N_722,In_246,In_61);
nor U723 (N_723,In_702,In_753);
nor U724 (N_724,In_518,In_191);
xnor U725 (N_725,In_126,In_536);
nand U726 (N_726,In_827,In_708);
nand U727 (N_727,In_305,In_153);
or U728 (N_728,In_933,In_418);
nand U729 (N_729,In_125,In_764);
nand U730 (N_730,In_455,In_833);
nor U731 (N_731,In_504,In_227);
nor U732 (N_732,In_583,In_556);
and U733 (N_733,In_771,In_9);
nor U734 (N_734,In_325,In_905);
and U735 (N_735,In_575,In_521);
or U736 (N_736,In_255,In_509);
nand U737 (N_737,In_317,In_982);
nand U738 (N_738,In_774,In_583);
nor U739 (N_739,In_496,In_650);
xor U740 (N_740,In_997,In_531);
and U741 (N_741,In_403,In_56);
or U742 (N_742,In_221,In_938);
nor U743 (N_743,In_431,In_915);
nand U744 (N_744,In_582,In_169);
nand U745 (N_745,In_566,In_472);
nor U746 (N_746,In_223,In_460);
nand U747 (N_747,In_439,In_524);
nor U748 (N_748,In_457,In_747);
nor U749 (N_749,In_956,In_344);
and U750 (N_750,In_55,In_112);
nand U751 (N_751,In_125,In_968);
xor U752 (N_752,In_808,In_693);
and U753 (N_753,In_654,In_385);
or U754 (N_754,In_51,In_81);
or U755 (N_755,In_135,In_312);
nand U756 (N_756,In_708,In_104);
and U757 (N_757,In_682,In_216);
nand U758 (N_758,In_908,In_267);
xnor U759 (N_759,In_5,In_327);
and U760 (N_760,In_344,In_825);
nand U761 (N_761,In_650,In_601);
nand U762 (N_762,In_183,In_600);
xor U763 (N_763,In_276,In_579);
nand U764 (N_764,In_703,In_825);
or U765 (N_765,In_661,In_114);
nand U766 (N_766,In_242,In_949);
xnor U767 (N_767,In_504,In_418);
nor U768 (N_768,In_836,In_523);
or U769 (N_769,In_649,In_61);
and U770 (N_770,In_745,In_73);
or U771 (N_771,In_556,In_228);
xor U772 (N_772,In_872,In_691);
or U773 (N_773,In_533,In_917);
and U774 (N_774,In_629,In_784);
nor U775 (N_775,In_766,In_100);
and U776 (N_776,In_246,In_786);
xnor U777 (N_777,In_494,In_170);
nand U778 (N_778,In_555,In_270);
or U779 (N_779,In_225,In_714);
nor U780 (N_780,In_676,In_867);
or U781 (N_781,In_574,In_226);
or U782 (N_782,In_625,In_400);
or U783 (N_783,In_332,In_483);
nor U784 (N_784,In_714,In_664);
nor U785 (N_785,In_317,In_76);
nand U786 (N_786,In_615,In_91);
nor U787 (N_787,In_588,In_775);
nand U788 (N_788,In_151,In_327);
nor U789 (N_789,In_235,In_184);
and U790 (N_790,In_876,In_477);
nand U791 (N_791,In_696,In_917);
nor U792 (N_792,In_772,In_29);
and U793 (N_793,In_990,In_746);
nand U794 (N_794,In_332,In_885);
nand U795 (N_795,In_646,In_189);
xnor U796 (N_796,In_300,In_48);
or U797 (N_797,In_713,In_999);
or U798 (N_798,In_69,In_699);
nand U799 (N_799,In_97,In_616);
or U800 (N_800,In_402,In_340);
and U801 (N_801,In_595,In_405);
and U802 (N_802,In_970,In_920);
or U803 (N_803,In_402,In_47);
nand U804 (N_804,In_219,In_638);
and U805 (N_805,In_99,In_854);
nand U806 (N_806,In_318,In_492);
and U807 (N_807,In_979,In_48);
and U808 (N_808,In_420,In_742);
xnor U809 (N_809,In_953,In_918);
nor U810 (N_810,In_966,In_312);
or U811 (N_811,In_272,In_702);
nand U812 (N_812,In_282,In_756);
or U813 (N_813,In_740,In_165);
or U814 (N_814,In_167,In_126);
nor U815 (N_815,In_988,In_911);
or U816 (N_816,In_788,In_724);
or U817 (N_817,In_808,In_584);
nor U818 (N_818,In_651,In_223);
and U819 (N_819,In_648,In_364);
or U820 (N_820,In_21,In_789);
or U821 (N_821,In_667,In_431);
or U822 (N_822,In_249,In_927);
nor U823 (N_823,In_122,In_808);
or U824 (N_824,In_598,In_860);
nand U825 (N_825,In_308,In_862);
nor U826 (N_826,In_672,In_233);
and U827 (N_827,In_910,In_538);
nor U828 (N_828,In_343,In_523);
nand U829 (N_829,In_329,In_54);
or U830 (N_830,In_887,In_206);
or U831 (N_831,In_673,In_931);
nand U832 (N_832,In_390,In_449);
or U833 (N_833,In_375,In_804);
and U834 (N_834,In_200,In_823);
nor U835 (N_835,In_820,In_994);
and U836 (N_836,In_447,In_198);
xor U837 (N_837,In_638,In_850);
xor U838 (N_838,In_53,In_229);
nor U839 (N_839,In_870,In_87);
nor U840 (N_840,In_92,In_745);
nand U841 (N_841,In_62,In_786);
nor U842 (N_842,In_247,In_216);
nor U843 (N_843,In_854,In_398);
and U844 (N_844,In_43,In_531);
nand U845 (N_845,In_248,In_204);
and U846 (N_846,In_521,In_171);
or U847 (N_847,In_858,In_262);
or U848 (N_848,In_811,In_705);
nand U849 (N_849,In_418,In_155);
xor U850 (N_850,In_343,In_556);
nor U851 (N_851,In_744,In_545);
nand U852 (N_852,In_334,In_193);
and U853 (N_853,In_558,In_799);
nor U854 (N_854,In_658,In_480);
nand U855 (N_855,In_687,In_684);
nor U856 (N_856,In_510,In_116);
nand U857 (N_857,In_873,In_729);
nor U858 (N_858,In_520,In_450);
and U859 (N_859,In_989,In_51);
or U860 (N_860,In_986,In_798);
or U861 (N_861,In_751,In_781);
nor U862 (N_862,In_536,In_389);
and U863 (N_863,In_721,In_514);
nor U864 (N_864,In_780,In_637);
and U865 (N_865,In_746,In_821);
or U866 (N_866,In_280,In_694);
nand U867 (N_867,In_837,In_881);
and U868 (N_868,In_334,In_357);
xor U869 (N_869,In_898,In_874);
xnor U870 (N_870,In_601,In_971);
xnor U871 (N_871,In_390,In_410);
or U872 (N_872,In_4,In_776);
nor U873 (N_873,In_521,In_950);
or U874 (N_874,In_712,In_771);
and U875 (N_875,In_310,In_317);
and U876 (N_876,In_51,In_258);
nor U877 (N_877,In_757,In_556);
or U878 (N_878,In_976,In_176);
and U879 (N_879,In_938,In_271);
and U880 (N_880,In_941,In_265);
or U881 (N_881,In_256,In_104);
or U882 (N_882,In_56,In_792);
xor U883 (N_883,In_110,In_132);
nor U884 (N_884,In_453,In_422);
and U885 (N_885,In_222,In_369);
nor U886 (N_886,In_493,In_829);
nand U887 (N_887,In_426,In_235);
nand U888 (N_888,In_213,In_263);
or U889 (N_889,In_898,In_262);
or U890 (N_890,In_604,In_891);
or U891 (N_891,In_299,In_238);
xnor U892 (N_892,In_643,In_962);
and U893 (N_893,In_413,In_562);
nor U894 (N_894,In_750,In_440);
xnor U895 (N_895,In_862,In_27);
or U896 (N_896,In_755,In_173);
nor U897 (N_897,In_812,In_915);
nor U898 (N_898,In_543,In_981);
and U899 (N_899,In_207,In_898);
nand U900 (N_900,In_67,In_770);
and U901 (N_901,In_200,In_672);
nor U902 (N_902,In_836,In_442);
or U903 (N_903,In_30,In_750);
or U904 (N_904,In_587,In_52);
or U905 (N_905,In_143,In_729);
nor U906 (N_906,In_531,In_499);
and U907 (N_907,In_688,In_542);
nand U908 (N_908,In_261,In_501);
nand U909 (N_909,In_901,In_356);
nand U910 (N_910,In_135,In_601);
nand U911 (N_911,In_549,In_309);
and U912 (N_912,In_628,In_281);
nor U913 (N_913,In_844,In_11);
or U914 (N_914,In_963,In_2);
or U915 (N_915,In_264,In_424);
or U916 (N_916,In_252,In_406);
or U917 (N_917,In_967,In_392);
nand U918 (N_918,In_963,In_463);
xnor U919 (N_919,In_136,In_675);
nor U920 (N_920,In_87,In_729);
and U921 (N_921,In_115,In_638);
and U922 (N_922,In_990,In_303);
or U923 (N_923,In_795,In_756);
and U924 (N_924,In_541,In_948);
or U925 (N_925,In_714,In_897);
and U926 (N_926,In_824,In_289);
nor U927 (N_927,In_264,In_505);
nor U928 (N_928,In_902,In_128);
xnor U929 (N_929,In_536,In_521);
and U930 (N_930,In_189,In_208);
nand U931 (N_931,In_959,In_571);
and U932 (N_932,In_381,In_210);
xnor U933 (N_933,In_921,In_478);
nand U934 (N_934,In_115,In_804);
or U935 (N_935,In_521,In_547);
nand U936 (N_936,In_447,In_372);
nor U937 (N_937,In_774,In_673);
nor U938 (N_938,In_660,In_869);
nor U939 (N_939,In_206,In_711);
nand U940 (N_940,In_991,In_43);
nand U941 (N_941,In_568,In_539);
xnor U942 (N_942,In_704,In_541);
xnor U943 (N_943,In_27,In_513);
and U944 (N_944,In_208,In_766);
nor U945 (N_945,In_444,In_786);
nand U946 (N_946,In_716,In_318);
nor U947 (N_947,In_264,In_96);
nand U948 (N_948,In_776,In_769);
and U949 (N_949,In_795,In_371);
nor U950 (N_950,In_931,In_515);
nand U951 (N_951,In_215,In_937);
nand U952 (N_952,In_912,In_144);
nor U953 (N_953,In_431,In_106);
nor U954 (N_954,In_564,In_105);
nor U955 (N_955,In_302,In_305);
nand U956 (N_956,In_278,In_662);
nor U957 (N_957,In_791,In_98);
and U958 (N_958,In_456,In_37);
and U959 (N_959,In_218,In_944);
and U960 (N_960,In_780,In_974);
xnor U961 (N_961,In_112,In_999);
or U962 (N_962,In_628,In_374);
xor U963 (N_963,In_180,In_3);
and U964 (N_964,In_61,In_198);
and U965 (N_965,In_409,In_825);
xor U966 (N_966,In_91,In_876);
or U967 (N_967,In_296,In_436);
or U968 (N_968,In_134,In_560);
nor U969 (N_969,In_708,In_241);
nand U970 (N_970,In_295,In_903);
and U971 (N_971,In_801,In_628);
and U972 (N_972,In_94,In_826);
or U973 (N_973,In_448,In_112);
nor U974 (N_974,In_232,In_754);
or U975 (N_975,In_125,In_923);
nand U976 (N_976,In_782,In_969);
and U977 (N_977,In_144,In_498);
nand U978 (N_978,In_457,In_49);
or U979 (N_979,In_454,In_252);
or U980 (N_980,In_382,In_105);
nor U981 (N_981,In_864,In_371);
or U982 (N_982,In_131,In_648);
nand U983 (N_983,In_346,In_684);
or U984 (N_984,In_234,In_761);
and U985 (N_985,In_781,In_638);
xor U986 (N_986,In_857,In_36);
and U987 (N_987,In_393,In_695);
nand U988 (N_988,In_305,In_133);
and U989 (N_989,In_5,In_753);
or U990 (N_990,In_129,In_104);
and U991 (N_991,In_494,In_886);
and U992 (N_992,In_281,In_66);
and U993 (N_993,In_818,In_61);
nand U994 (N_994,In_0,In_152);
nor U995 (N_995,In_669,In_909);
or U996 (N_996,In_70,In_34);
or U997 (N_997,In_563,In_694);
nor U998 (N_998,In_795,In_158);
nand U999 (N_999,In_383,In_639);
nand U1000 (N_1000,In_824,In_24);
and U1001 (N_1001,In_962,In_441);
nor U1002 (N_1002,In_304,In_845);
xor U1003 (N_1003,In_165,In_242);
nand U1004 (N_1004,In_189,In_577);
or U1005 (N_1005,In_740,In_392);
and U1006 (N_1006,In_62,In_991);
nor U1007 (N_1007,In_636,In_913);
nand U1008 (N_1008,In_235,In_143);
nand U1009 (N_1009,In_589,In_925);
nand U1010 (N_1010,In_114,In_796);
and U1011 (N_1011,In_142,In_330);
and U1012 (N_1012,In_763,In_379);
nand U1013 (N_1013,In_456,In_484);
nor U1014 (N_1014,In_325,In_225);
and U1015 (N_1015,In_839,In_348);
xor U1016 (N_1016,In_549,In_332);
and U1017 (N_1017,In_396,In_715);
or U1018 (N_1018,In_651,In_646);
nor U1019 (N_1019,In_823,In_73);
nand U1020 (N_1020,In_707,In_752);
nor U1021 (N_1021,In_781,In_804);
or U1022 (N_1022,In_868,In_198);
and U1023 (N_1023,In_998,In_198);
or U1024 (N_1024,In_603,In_708);
and U1025 (N_1025,In_107,In_422);
xor U1026 (N_1026,In_578,In_902);
xor U1027 (N_1027,In_369,In_157);
xnor U1028 (N_1028,In_52,In_817);
xor U1029 (N_1029,In_140,In_172);
nand U1030 (N_1030,In_423,In_654);
nor U1031 (N_1031,In_718,In_936);
nor U1032 (N_1032,In_95,In_694);
or U1033 (N_1033,In_431,In_2);
or U1034 (N_1034,In_737,In_255);
xor U1035 (N_1035,In_604,In_330);
nor U1036 (N_1036,In_543,In_510);
or U1037 (N_1037,In_822,In_586);
or U1038 (N_1038,In_619,In_398);
and U1039 (N_1039,In_207,In_152);
and U1040 (N_1040,In_703,In_895);
or U1041 (N_1041,In_694,In_657);
or U1042 (N_1042,In_377,In_442);
or U1043 (N_1043,In_796,In_875);
nand U1044 (N_1044,In_953,In_230);
and U1045 (N_1045,In_684,In_771);
nand U1046 (N_1046,In_269,In_387);
and U1047 (N_1047,In_39,In_926);
or U1048 (N_1048,In_177,In_476);
nor U1049 (N_1049,In_94,In_137);
nand U1050 (N_1050,In_871,In_962);
or U1051 (N_1051,In_260,In_676);
and U1052 (N_1052,In_292,In_610);
or U1053 (N_1053,In_305,In_854);
or U1054 (N_1054,In_816,In_956);
or U1055 (N_1055,In_518,In_418);
nand U1056 (N_1056,In_762,In_261);
xor U1057 (N_1057,In_76,In_683);
nand U1058 (N_1058,In_111,In_963);
nand U1059 (N_1059,In_404,In_963);
and U1060 (N_1060,In_767,In_667);
nor U1061 (N_1061,In_163,In_278);
nor U1062 (N_1062,In_571,In_480);
and U1063 (N_1063,In_581,In_347);
nand U1064 (N_1064,In_600,In_800);
nor U1065 (N_1065,In_258,In_0);
or U1066 (N_1066,In_201,In_413);
nor U1067 (N_1067,In_155,In_961);
nand U1068 (N_1068,In_91,In_987);
nor U1069 (N_1069,In_728,In_533);
nand U1070 (N_1070,In_577,In_552);
and U1071 (N_1071,In_707,In_828);
nor U1072 (N_1072,In_785,In_672);
nor U1073 (N_1073,In_611,In_637);
and U1074 (N_1074,In_147,In_723);
and U1075 (N_1075,In_661,In_636);
nand U1076 (N_1076,In_333,In_311);
and U1077 (N_1077,In_911,In_515);
nand U1078 (N_1078,In_162,In_313);
nor U1079 (N_1079,In_162,In_625);
and U1080 (N_1080,In_887,In_402);
or U1081 (N_1081,In_487,In_976);
xnor U1082 (N_1082,In_789,In_22);
nand U1083 (N_1083,In_276,In_422);
and U1084 (N_1084,In_638,In_396);
nor U1085 (N_1085,In_661,In_532);
nand U1086 (N_1086,In_284,In_883);
or U1087 (N_1087,In_931,In_243);
or U1088 (N_1088,In_691,In_166);
nand U1089 (N_1089,In_784,In_929);
or U1090 (N_1090,In_465,In_734);
xnor U1091 (N_1091,In_363,In_76);
nand U1092 (N_1092,In_605,In_851);
nand U1093 (N_1093,In_576,In_523);
nand U1094 (N_1094,In_5,In_776);
nand U1095 (N_1095,In_260,In_288);
and U1096 (N_1096,In_171,In_163);
and U1097 (N_1097,In_563,In_925);
nor U1098 (N_1098,In_541,In_950);
nand U1099 (N_1099,In_836,In_920);
nor U1100 (N_1100,In_147,In_805);
nand U1101 (N_1101,In_97,In_18);
nor U1102 (N_1102,In_315,In_655);
and U1103 (N_1103,In_190,In_309);
nor U1104 (N_1104,In_34,In_493);
and U1105 (N_1105,In_433,In_880);
nor U1106 (N_1106,In_863,In_256);
xnor U1107 (N_1107,In_840,In_398);
and U1108 (N_1108,In_461,In_605);
and U1109 (N_1109,In_735,In_79);
and U1110 (N_1110,In_145,In_875);
and U1111 (N_1111,In_124,In_37);
or U1112 (N_1112,In_186,In_752);
xor U1113 (N_1113,In_48,In_257);
nor U1114 (N_1114,In_72,In_920);
xnor U1115 (N_1115,In_536,In_600);
or U1116 (N_1116,In_404,In_733);
xor U1117 (N_1117,In_718,In_663);
or U1118 (N_1118,In_743,In_346);
or U1119 (N_1119,In_942,In_433);
or U1120 (N_1120,In_268,In_940);
or U1121 (N_1121,In_75,In_4);
and U1122 (N_1122,In_477,In_457);
nor U1123 (N_1123,In_512,In_991);
nand U1124 (N_1124,In_636,In_922);
or U1125 (N_1125,In_972,In_893);
xor U1126 (N_1126,In_857,In_414);
nor U1127 (N_1127,In_417,In_176);
nand U1128 (N_1128,In_183,In_737);
nand U1129 (N_1129,In_265,In_435);
nor U1130 (N_1130,In_842,In_392);
nor U1131 (N_1131,In_14,In_401);
nand U1132 (N_1132,In_853,In_388);
nand U1133 (N_1133,In_94,In_707);
xor U1134 (N_1134,In_635,In_629);
nand U1135 (N_1135,In_41,In_236);
or U1136 (N_1136,In_27,In_679);
or U1137 (N_1137,In_781,In_125);
and U1138 (N_1138,In_920,In_647);
nor U1139 (N_1139,In_157,In_481);
xor U1140 (N_1140,In_356,In_594);
xor U1141 (N_1141,In_946,In_91);
nand U1142 (N_1142,In_270,In_185);
xnor U1143 (N_1143,In_732,In_926);
nor U1144 (N_1144,In_243,In_981);
nor U1145 (N_1145,In_119,In_814);
and U1146 (N_1146,In_77,In_441);
nand U1147 (N_1147,In_19,In_300);
nor U1148 (N_1148,In_767,In_35);
nor U1149 (N_1149,In_731,In_177);
or U1150 (N_1150,In_897,In_215);
or U1151 (N_1151,In_877,In_868);
nand U1152 (N_1152,In_537,In_580);
nand U1153 (N_1153,In_728,In_566);
xnor U1154 (N_1154,In_295,In_168);
nand U1155 (N_1155,In_232,In_844);
and U1156 (N_1156,In_6,In_934);
xnor U1157 (N_1157,In_777,In_281);
nand U1158 (N_1158,In_102,In_757);
nor U1159 (N_1159,In_263,In_903);
nand U1160 (N_1160,In_463,In_575);
and U1161 (N_1161,In_600,In_996);
nor U1162 (N_1162,In_496,In_639);
or U1163 (N_1163,In_172,In_243);
nand U1164 (N_1164,In_925,In_962);
nor U1165 (N_1165,In_810,In_744);
or U1166 (N_1166,In_382,In_522);
xor U1167 (N_1167,In_24,In_88);
xor U1168 (N_1168,In_197,In_508);
or U1169 (N_1169,In_221,In_957);
or U1170 (N_1170,In_65,In_730);
and U1171 (N_1171,In_459,In_638);
and U1172 (N_1172,In_253,In_367);
nor U1173 (N_1173,In_388,In_228);
or U1174 (N_1174,In_702,In_329);
xnor U1175 (N_1175,In_553,In_176);
nor U1176 (N_1176,In_199,In_194);
nor U1177 (N_1177,In_357,In_538);
or U1178 (N_1178,In_832,In_786);
nor U1179 (N_1179,In_691,In_226);
or U1180 (N_1180,In_490,In_721);
nor U1181 (N_1181,In_664,In_651);
xnor U1182 (N_1182,In_147,In_152);
and U1183 (N_1183,In_717,In_35);
nand U1184 (N_1184,In_235,In_849);
nor U1185 (N_1185,In_304,In_206);
and U1186 (N_1186,In_730,In_551);
or U1187 (N_1187,In_255,In_918);
nand U1188 (N_1188,In_562,In_848);
nor U1189 (N_1189,In_24,In_447);
nor U1190 (N_1190,In_781,In_260);
or U1191 (N_1191,In_664,In_703);
and U1192 (N_1192,In_811,In_803);
and U1193 (N_1193,In_459,In_41);
nand U1194 (N_1194,In_14,In_428);
and U1195 (N_1195,In_142,In_291);
and U1196 (N_1196,In_727,In_820);
and U1197 (N_1197,In_337,In_673);
or U1198 (N_1198,In_683,In_342);
xor U1199 (N_1199,In_671,In_390);
nand U1200 (N_1200,In_509,In_847);
nand U1201 (N_1201,In_983,In_363);
nand U1202 (N_1202,In_366,In_789);
and U1203 (N_1203,In_921,In_948);
or U1204 (N_1204,In_787,In_56);
nor U1205 (N_1205,In_94,In_917);
or U1206 (N_1206,In_900,In_541);
or U1207 (N_1207,In_288,In_920);
nand U1208 (N_1208,In_439,In_930);
nand U1209 (N_1209,In_241,In_795);
nand U1210 (N_1210,In_480,In_302);
and U1211 (N_1211,In_442,In_72);
xnor U1212 (N_1212,In_223,In_689);
and U1213 (N_1213,In_189,In_272);
nand U1214 (N_1214,In_319,In_742);
nor U1215 (N_1215,In_451,In_781);
xnor U1216 (N_1216,In_528,In_987);
or U1217 (N_1217,In_821,In_740);
or U1218 (N_1218,In_192,In_61);
xor U1219 (N_1219,In_948,In_674);
xnor U1220 (N_1220,In_349,In_922);
xor U1221 (N_1221,In_632,In_374);
or U1222 (N_1222,In_417,In_5);
nand U1223 (N_1223,In_819,In_67);
and U1224 (N_1224,In_800,In_510);
or U1225 (N_1225,In_271,In_620);
nor U1226 (N_1226,In_221,In_904);
nand U1227 (N_1227,In_431,In_366);
or U1228 (N_1228,In_166,In_750);
nor U1229 (N_1229,In_537,In_66);
nor U1230 (N_1230,In_84,In_642);
nor U1231 (N_1231,In_957,In_459);
nor U1232 (N_1232,In_814,In_893);
nand U1233 (N_1233,In_958,In_272);
and U1234 (N_1234,In_260,In_592);
or U1235 (N_1235,In_888,In_208);
xnor U1236 (N_1236,In_430,In_997);
and U1237 (N_1237,In_512,In_683);
nand U1238 (N_1238,In_573,In_762);
or U1239 (N_1239,In_254,In_94);
and U1240 (N_1240,In_926,In_441);
or U1241 (N_1241,In_475,In_771);
or U1242 (N_1242,In_162,In_978);
nor U1243 (N_1243,In_383,In_974);
and U1244 (N_1244,In_302,In_289);
and U1245 (N_1245,In_338,In_385);
and U1246 (N_1246,In_486,In_841);
or U1247 (N_1247,In_723,In_892);
nor U1248 (N_1248,In_522,In_492);
nor U1249 (N_1249,In_436,In_644);
or U1250 (N_1250,In_454,In_10);
nor U1251 (N_1251,In_169,In_663);
or U1252 (N_1252,In_88,In_222);
or U1253 (N_1253,In_890,In_380);
nor U1254 (N_1254,In_191,In_77);
nand U1255 (N_1255,In_991,In_76);
nand U1256 (N_1256,In_685,In_999);
and U1257 (N_1257,In_975,In_36);
or U1258 (N_1258,In_51,In_489);
nor U1259 (N_1259,In_738,In_481);
xor U1260 (N_1260,In_296,In_109);
nor U1261 (N_1261,In_299,In_472);
xor U1262 (N_1262,In_896,In_581);
xor U1263 (N_1263,In_315,In_991);
and U1264 (N_1264,In_53,In_894);
nor U1265 (N_1265,In_290,In_408);
or U1266 (N_1266,In_3,In_946);
or U1267 (N_1267,In_140,In_213);
and U1268 (N_1268,In_579,In_398);
nor U1269 (N_1269,In_386,In_181);
and U1270 (N_1270,In_463,In_765);
nor U1271 (N_1271,In_63,In_640);
and U1272 (N_1272,In_810,In_311);
xor U1273 (N_1273,In_948,In_83);
or U1274 (N_1274,In_980,In_592);
nor U1275 (N_1275,In_101,In_190);
nor U1276 (N_1276,In_389,In_810);
or U1277 (N_1277,In_223,In_730);
nand U1278 (N_1278,In_782,In_7);
or U1279 (N_1279,In_55,In_881);
or U1280 (N_1280,In_896,In_100);
and U1281 (N_1281,In_567,In_316);
or U1282 (N_1282,In_872,In_721);
or U1283 (N_1283,In_961,In_990);
and U1284 (N_1284,In_236,In_817);
and U1285 (N_1285,In_536,In_345);
and U1286 (N_1286,In_268,In_987);
and U1287 (N_1287,In_393,In_113);
nand U1288 (N_1288,In_457,In_405);
nor U1289 (N_1289,In_851,In_473);
and U1290 (N_1290,In_354,In_586);
or U1291 (N_1291,In_900,In_360);
and U1292 (N_1292,In_967,In_919);
or U1293 (N_1293,In_9,In_756);
and U1294 (N_1294,In_929,In_362);
nand U1295 (N_1295,In_935,In_87);
or U1296 (N_1296,In_35,In_744);
xnor U1297 (N_1297,In_25,In_362);
and U1298 (N_1298,In_272,In_95);
nand U1299 (N_1299,In_475,In_518);
nor U1300 (N_1300,In_570,In_378);
nor U1301 (N_1301,In_397,In_613);
or U1302 (N_1302,In_86,In_699);
nand U1303 (N_1303,In_977,In_967);
nand U1304 (N_1304,In_954,In_17);
or U1305 (N_1305,In_722,In_541);
nor U1306 (N_1306,In_179,In_783);
nand U1307 (N_1307,In_580,In_162);
nor U1308 (N_1308,In_178,In_230);
and U1309 (N_1309,In_450,In_853);
and U1310 (N_1310,In_89,In_860);
or U1311 (N_1311,In_629,In_282);
and U1312 (N_1312,In_845,In_376);
and U1313 (N_1313,In_734,In_255);
xor U1314 (N_1314,In_359,In_556);
and U1315 (N_1315,In_960,In_707);
or U1316 (N_1316,In_201,In_946);
nand U1317 (N_1317,In_228,In_216);
nor U1318 (N_1318,In_712,In_583);
nand U1319 (N_1319,In_101,In_213);
nand U1320 (N_1320,In_493,In_410);
nor U1321 (N_1321,In_838,In_911);
and U1322 (N_1322,In_207,In_399);
and U1323 (N_1323,In_346,In_471);
or U1324 (N_1324,In_69,In_788);
or U1325 (N_1325,In_363,In_346);
and U1326 (N_1326,In_82,In_128);
nor U1327 (N_1327,In_13,In_107);
nor U1328 (N_1328,In_973,In_413);
or U1329 (N_1329,In_769,In_296);
xor U1330 (N_1330,In_538,In_256);
nor U1331 (N_1331,In_816,In_950);
or U1332 (N_1332,In_455,In_475);
or U1333 (N_1333,In_653,In_64);
and U1334 (N_1334,In_839,In_84);
and U1335 (N_1335,In_836,In_346);
nand U1336 (N_1336,In_575,In_545);
or U1337 (N_1337,In_340,In_951);
nor U1338 (N_1338,In_612,In_144);
nor U1339 (N_1339,In_373,In_198);
and U1340 (N_1340,In_108,In_17);
or U1341 (N_1341,In_667,In_386);
nand U1342 (N_1342,In_420,In_325);
or U1343 (N_1343,In_641,In_813);
and U1344 (N_1344,In_108,In_556);
nand U1345 (N_1345,In_159,In_293);
nor U1346 (N_1346,In_608,In_237);
nor U1347 (N_1347,In_59,In_233);
and U1348 (N_1348,In_146,In_148);
or U1349 (N_1349,In_405,In_89);
xor U1350 (N_1350,In_837,In_726);
and U1351 (N_1351,In_777,In_564);
or U1352 (N_1352,In_737,In_859);
or U1353 (N_1353,In_224,In_207);
and U1354 (N_1354,In_301,In_54);
or U1355 (N_1355,In_164,In_864);
and U1356 (N_1356,In_858,In_645);
and U1357 (N_1357,In_564,In_635);
nor U1358 (N_1358,In_39,In_118);
and U1359 (N_1359,In_296,In_569);
nor U1360 (N_1360,In_385,In_870);
and U1361 (N_1361,In_528,In_128);
nand U1362 (N_1362,In_794,In_950);
nand U1363 (N_1363,In_666,In_449);
nor U1364 (N_1364,In_523,In_642);
and U1365 (N_1365,In_317,In_74);
or U1366 (N_1366,In_92,In_909);
xor U1367 (N_1367,In_748,In_245);
nor U1368 (N_1368,In_520,In_528);
or U1369 (N_1369,In_7,In_499);
or U1370 (N_1370,In_597,In_240);
or U1371 (N_1371,In_565,In_541);
and U1372 (N_1372,In_941,In_93);
and U1373 (N_1373,In_554,In_563);
or U1374 (N_1374,In_38,In_948);
nand U1375 (N_1375,In_612,In_254);
nor U1376 (N_1376,In_12,In_618);
nor U1377 (N_1377,In_620,In_66);
nand U1378 (N_1378,In_486,In_552);
or U1379 (N_1379,In_795,In_582);
or U1380 (N_1380,In_859,In_305);
nand U1381 (N_1381,In_821,In_591);
and U1382 (N_1382,In_533,In_739);
or U1383 (N_1383,In_784,In_185);
xnor U1384 (N_1384,In_693,In_996);
nor U1385 (N_1385,In_378,In_670);
and U1386 (N_1386,In_967,In_528);
nor U1387 (N_1387,In_816,In_87);
nor U1388 (N_1388,In_483,In_682);
nor U1389 (N_1389,In_804,In_711);
and U1390 (N_1390,In_528,In_345);
xnor U1391 (N_1391,In_149,In_301);
or U1392 (N_1392,In_568,In_922);
or U1393 (N_1393,In_90,In_33);
nor U1394 (N_1394,In_712,In_201);
or U1395 (N_1395,In_62,In_943);
and U1396 (N_1396,In_308,In_954);
or U1397 (N_1397,In_231,In_151);
nand U1398 (N_1398,In_963,In_449);
nand U1399 (N_1399,In_850,In_988);
nand U1400 (N_1400,In_456,In_626);
nor U1401 (N_1401,In_375,In_544);
and U1402 (N_1402,In_902,In_991);
nand U1403 (N_1403,In_515,In_77);
and U1404 (N_1404,In_163,In_537);
or U1405 (N_1405,In_309,In_506);
nor U1406 (N_1406,In_93,In_845);
nor U1407 (N_1407,In_956,In_978);
nand U1408 (N_1408,In_818,In_847);
nand U1409 (N_1409,In_216,In_870);
xnor U1410 (N_1410,In_613,In_906);
xor U1411 (N_1411,In_677,In_184);
or U1412 (N_1412,In_771,In_897);
nor U1413 (N_1413,In_404,In_713);
nand U1414 (N_1414,In_858,In_800);
nand U1415 (N_1415,In_990,In_945);
or U1416 (N_1416,In_182,In_574);
nor U1417 (N_1417,In_228,In_184);
and U1418 (N_1418,In_82,In_847);
nor U1419 (N_1419,In_101,In_310);
or U1420 (N_1420,In_791,In_86);
nand U1421 (N_1421,In_68,In_904);
or U1422 (N_1422,In_855,In_225);
nor U1423 (N_1423,In_166,In_223);
or U1424 (N_1424,In_329,In_335);
nor U1425 (N_1425,In_329,In_856);
nor U1426 (N_1426,In_478,In_271);
nand U1427 (N_1427,In_702,In_506);
xnor U1428 (N_1428,In_388,In_639);
nand U1429 (N_1429,In_970,In_990);
nor U1430 (N_1430,In_791,In_166);
or U1431 (N_1431,In_714,In_673);
nand U1432 (N_1432,In_969,In_399);
or U1433 (N_1433,In_353,In_424);
xor U1434 (N_1434,In_26,In_382);
and U1435 (N_1435,In_900,In_870);
and U1436 (N_1436,In_529,In_483);
nor U1437 (N_1437,In_58,In_271);
and U1438 (N_1438,In_375,In_184);
nor U1439 (N_1439,In_882,In_355);
nor U1440 (N_1440,In_372,In_233);
nor U1441 (N_1441,In_650,In_301);
nor U1442 (N_1442,In_248,In_376);
or U1443 (N_1443,In_333,In_10);
and U1444 (N_1444,In_478,In_858);
nor U1445 (N_1445,In_134,In_421);
and U1446 (N_1446,In_283,In_746);
xor U1447 (N_1447,In_600,In_812);
or U1448 (N_1448,In_160,In_159);
or U1449 (N_1449,In_55,In_811);
nand U1450 (N_1450,In_774,In_814);
or U1451 (N_1451,In_87,In_687);
nand U1452 (N_1452,In_469,In_865);
nand U1453 (N_1453,In_994,In_428);
or U1454 (N_1454,In_76,In_303);
nand U1455 (N_1455,In_754,In_104);
nand U1456 (N_1456,In_610,In_265);
and U1457 (N_1457,In_447,In_282);
nand U1458 (N_1458,In_137,In_134);
nand U1459 (N_1459,In_286,In_810);
nor U1460 (N_1460,In_545,In_356);
and U1461 (N_1461,In_232,In_578);
nor U1462 (N_1462,In_260,In_833);
xor U1463 (N_1463,In_409,In_141);
and U1464 (N_1464,In_662,In_910);
xor U1465 (N_1465,In_363,In_124);
and U1466 (N_1466,In_815,In_278);
nand U1467 (N_1467,In_425,In_993);
nand U1468 (N_1468,In_750,In_798);
or U1469 (N_1469,In_221,In_325);
or U1470 (N_1470,In_959,In_141);
and U1471 (N_1471,In_669,In_889);
or U1472 (N_1472,In_114,In_56);
and U1473 (N_1473,In_506,In_88);
nor U1474 (N_1474,In_605,In_515);
and U1475 (N_1475,In_574,In_477);
nor U1476 (N_1476,In_295,In_604);
nor U1477 (N_1477,In_160,In_86);
or U1478 (N_1478,In_760,In_819);
xor U1479 (N_1479,In_719,In_81);
nor U1480 (N_1480,In_818,In_257);
xnor U1481 (N_1481,In_176,In_507);
nand U1482 (N_1482,In_921,In_993);
and U1483 (N_1483,In_0,In_808);
and U1484 (N_1484,In_373,In_205);
xnor U1485 (N_1485,In_923,In_68);
or U1486 (N_1486,In_732,In_349);
nand U1487 (N_1487,In_169,In_768);
nand U1488 (N_1488,In_534,In_831);
xor U1489 (N_1489,In_316,In_917);
nand U1490 (N_1490,In_115,In_20);
and U1491 (N_1491,In_710,In_5);
or U1492 (N_1492,In_404,In_743);
xor U1493 (N_1493,In_361,In_158);
and U1494 (N_1494,In_263,In_323);
and U1495 (N_1495,In_315,In_137);
nor U1496 (N_1496,In_799,In_636);
nand U1497 (N_1497,In_382,In_578);
nand U1498 (N_1498,In_825,In_36);
nor U1499 (N_1499,In_707,In_159);
nor U1500 (N_1500,In_252,In_249);
and U1501 (N_1501,In_10,In_792);
or U1502 (N_1502,In_264,In_751);
or U1503 (N_1503,In_596,In_784);
nand U1504 (N_1504,In_585,In_245);
nor U1505 (N_1505,In_749,In_24);
and U1506 (N_1506,In_772,In_647);
nand U1507 (N_1507,In_302,In_971);
or U1508 (N_1508,In_954,In_288);
and U1509 (N_1509,In_418,In_873);
xor U1510 (N_1510,In_304,In_195);
and U1511 (N_1511,In_109,In_892);
or U1512 (N_1512,In_69,In_583);
nor U1513 (N_1513,In_689,In_941);
nor U1514 (N_1514,In_31,In_132);
or U1515 (N_1515,In_830,In_544);
nand U1516 (N_1516,In_938,In_700);
nor U1517 (N_1517,In_866,In_148);
nor U1518 (N_1518,In_533,In_42);
and U1519 (N_1519,In_996,In_360);
nand U1520 (N_1520,In_855,In_245);
and U1521 (N_1521,In_650,In_682);
nand U1522 (N_1522,In_922,In_528);
xor U1523 (N_1523,In_294,In_28);
nand U1524 (N_1524,In_723,In_926);
nand U1525 (N_1525,In_554,In_943);
and U1526 (N_1526,In_563,In_47);
and U1527 (N_1527,In_469,In_368);
nor U1528 (N_1528,In_752,In_278);
xnor U1529 (N_1529,In_837,In_684);
and U1530 (N_1530,In_512,In_325);
xnor U1531 (N_1531,In_647,In_19);
or U1532 (N_1532,In_538,In_307);
and U1533 (N_1533,In_563,In_155);
and U1534 (N_1534,In_75,In_769);
nand U1535 (N_1535,In_775,In_654);
nand U1536 (N_1536,In_937,In_585);
xnor U1537 (N_1537,In_113,In_114);
and U1538 (N_1538,In_80,In_287);
or U1539 (N_1539,In_139,In_282);
nor U1540 (N_1540,In_241,In_146);
nor U1541 (N_1541,In_329,In_795);
or U1542 (N_1542,In_971,In_932);
and U1543 (N_1543,In_450,In_193);
nand U1544 (N_1544,In_256,In_302);
xnor U1545 (N_1545,In_593,In_188);
nor U1546 (N_1546,In_603,In_701);
or U1547 (N_1547,In_899,In_150);
nand U1548 (N_1548,In_764,In_84);
nand U1549 (N_1549,In_239,In_298);
or U1550 (N_1550,In_961,In_881);
or U1551 (N_1551,In_426,In_200);
nand U1552 (N_1552,In_163,In_21);
nor U1553 (N_1553,In_985,In_523);
or U1554 (N_1554,In_680,In_849);
or U1555 (N_1555,In_955,In_567);
nand U1556 (N_1556,In_56,In_27);
and U1557 (N_1557,In_604,In_947);
nor U1558 (N_1558,In_154,In_560);
xor U1559 (N_1559,In_194,In_756);
and U1560 (N_1560,In_552,In_905);
nand U1561 (N_1561,In_209,In_795);
and U1562 (N_1562,In_311,In_425);
nand U1563 (N_1563,In_850,In_634);
nor U1564 (N_1564,In_630,In_127);
nand U1565 (N_1565,In_590,In_213);
and U1566 (N_1566,In_940,In_411);
nor U1567 (N_1567,In_534,In_280);
xnor U1568 (N_1568,In_509,In_298);
nand U1569 (N_1569,In_471,In_852);
or U1570 (N_1570,In_122,In_912);
xnor U1571 (N_1571,In_536,In_683);
nor U1572 (N_1572,In_40,In_597);
and U1573 (N_1573,In_202,In_812);
and U1574 (N_1574,In_830,In_846);
and U1575 (N_1575,In_224,In_140);
or U1576 (N_1576,In_924,In_541);
or U1577 (N_1577,In_380,In_50);
or U1578 (N_1578,In_486,In_983);
nor U1579 (N_1579,In_439,In_775);
nor U1580 (N_1580,In_947,In_575);
or U1581 (N_1581,In_932,In_514);
nor U1582 (N_1582,In_708,In_193);
nand U1583 (N_1583,In_878,In_547);
nor U1584 (N_1584,In_375,In_517);
or U1585 (N_1585,In_275,In_279);
or U1586 (N_1586,In_128,In_808);
and U1587 (N_1587,In_266,In_525);
nand U1588 (N_1588,In_653,In_265);
nand U1589 (N_1589,In_467,In_258);
and U1590 (N_1590,In_105,In_322);
nor U1591 (N_1591,In_113,In_16);
nand U1592 (N_1592,In_206,In_664);
xor U1593 (N_1593,In_677,In_278);
nand U1594 (N_1594,In_71,In_753);
nor U1595 (N_1595,In_272,In_303);
or U1596 (N_1596,In_725,In_358);
or U1597 (N_1597,In_263,In_162);
or U1598 (N_1598,In_698,In_600);
or U1599 (N_1599,In_582,In_955);
and U1600 (N_1600,In_466,In_739);
nor U1601 (N_1601,In_626,In_844);
or U1602 (N_1602,In_891,In_344);
or U1603 (N_1603,In_639,In_776);
nand U1604 (N_1604,In_86,In_836);
nor U1605 (N_1605,In_366,In_86);
and U1606 (N_1606,In_968,In_976);
and U1607 (N_1607,In_638,In_21);
nand U1608 (N_1608,In_631,In_211);
or U1609 (N_1609,In_232,In_353);
xor U1610 (N_1610,In_977,In_135);
and U1611 (N_1611,In_186,In_944);
nor U1612 (N_1612,In_976,In_549);
nand U1613 (N_1613,In_170,In_830);
or U1614 (N_1614,In_271,In_929);
and U1615 (N_1615,In_329,In_880);
and U1616 (N_1616,In_377,In_974);
and U1617 (N_1617,In_495,In_465);
nand U1618 (N_1618,In_912,In_865);
nor U1619 (N_1619,In_493,In_28);
nor U1620 (N_1620,In_211,In_925);
or U1621 (N_1621,In_309,In_139);
or U1622 (N_1622,In_113,In_640);
xnor U1623 (N_1623,In_2,In_853);
nor U1624 (N_1624,In_615,In_114);
xor U1625 (N_1625,In_879,In_855);
and U1626 (N_1626,In_511,In_939);
nor U1627 (N_1627,In_343,In_993);
nor U1628 (N_1628,In_31,In_446);
nor U1629 (N_1629,In_623,In_879);
nand U1630 (N_1630,In_654,In_534);
nor U1631 (N_1631,In_218,In_993);
xor U1632 (N_1632,In_117,In_930);
nor U1633 (N_1633,In_455,In_952);
nor U1634 (N_1634,In_208,In_343);
nor U1635 (N_1635,In_744,In_169);
nor U1636 (N_1636,In_696,In_12);
and U1637 (N_1637,In_803,In_82);
nor U1638 (N_1638,In_994,In_470);
or U1639 (N_1639,In_711,In_126);
and U1640 (N_1640,In_538,In_768);
xnor U1641 (N_1641,In_679,In_431);
nor U1642 (N_1642,In_265,In_45);
nand U1643 (N_1643,In_609,In_645);
nand U1644 (N_1644,In_508,In_558);
nand U1645 (N_1645,In_239,In_837);
nand U1646 (N_1646,In_652,In_579);
xnor U1647 (N_1647,In_20,In_232);
nand U1648 (N_1648,In_260,In_745);
nor U1649 (N_1649,In_511,In_551);
or U1650 (N_1650,In_403,In_397);
nand U1651 (N_1651,In_884,In_449);
nand U1652 (N_1652,In_588,In_170);
nand U1653 (N_1653,In_357,In_567);
nor U1654 (N_1654,In_230,In_747);
or U1655 (N_1655,In_545,In_428);
xor U1656 (N_1656,In_350,In_920);
nor U1657 (N_1657,In_710,In_812);
xor U1658 (N_1658,In_282,In_111);
nor U1659 (N_1659,In_295,In_850);
or U1660 (N_1660,In_360,In_407);
nand U1661 (N_1661,In_203,In_730);
or U1662 (N_1662,In_221,In_202);
nand U1663 (N_1663,In_891,In_296);
nand U1664 (N_1664,In_243,In_190);
nand U1665 (N_1665,In_679,In_960);
nor U1666 (N_1666,In_527,In_951);
nor U1667 (N_1667,In_941,In_577);
nand U1668 (N_1668,In_48,In_114);
nor U1669 (N_1669,In_251,In_227);
and U1670 (N_1670,In_93,In_208);
nand U1671 (N_1671,In_132,In_144);
nand U1672 (N_1672,In_687,In_649);
and U1673 (N_1673,In_325,In_410);
and U1674 (N_1674,In_579,In_83);
nor U1675 (N_1675,In_648,In_790);
and U1676 (N_1676,In_3,In_24);
nand U1677 (N_1677,In_865,In_162);
nand U1678 (N_1678,In_796,In_151);
and U1679 (N_1679,In_279,In_29);
nor U1680 (N_1680,In_530,In_907);
nor U1681 (N_1681,In_830,In_315);
and U1682 (N_1682,In_406,In_668);
and U1683 (N_1683,In_581,In_377);
and U1684 (N_1684,In_328,In_822);
nand U1685 (N_1685,In_606,In_337);
or U1686 (N_1686,In_392,In_939);
nand U1687 (N_1687,In_523,In_50);
or U1688 (N_1688,In_411,In_211);
nand U1689 (N_1689,In_732,In_607);
and U1690 (N_1690,In_436,In_807);
nor U1691 (N_1691,In_993,In_631);
xnor U1692 (N_1692,In_229,In_109);
nor U1693 (N_1693,In_711,In_940);
and U1694 (N_1694,In_261,In_67);
nand U1695 (N_1695,In_640,In_797);
or U1696 (N_1696,In_591,In_617);
nor U1697 (N_1697,In_251,In_163);
nand U1698 (N_1698,In_396,In_261);
and U1699 (N_1699,In_604,In_575);
and U1700 (N_1700,In_502,In_105);
or U1701 (N_1701,In_823,In_381);
and U1702 (N_1702,In_183,In_913);
nand U1703 (N_1703,In_893,In_940);
nor U1704 (N_1704,In_144,In_627);
and U1705 (N_1705,In_73,In_18);
nand U1706 (N_1706,In_703,In_953);
nor U1707 (N_1707,In_817,In_152);
or U1708 (N_1708,In_892,In_990);
nand U1709 (N_1709,In_267,In_4);
nor U1710 (N_1710,In_11,In_897);
nand U1711 (N_1711,In_778,In_329);
xnor U1712 (N_1712,In_528,In_165);
nor U1713 (N_1713,In_894,In_457);
or U1714 (N_1714,In_299,In_989);
and U1715 (N_1715,In_849,In_803);
or U1716 (N_1716,In_774,In_937);
xnor U1717 (N_1717,In_400,In_484);
or U1718 (N_1718,In_646,In_770);
or U1719 (N_1719,In_949,In_277);
nor U1720 (N_1720,In_279,In_111);
xnor U1721 (N_1721,In_502,In_773);
or U1722 (N_1722,In_449,In_5);
and U1723 (N_1723,In_853,In_886);
and U1724 (N_1724,In_621,In_924);
or U1725 (N_1725,In_19,In_534);
nand U1726 (N_1726,In_816,In_44);
and U1727 (N_1727,In_721,In_832);
and U1728 (N_1728,In_876,In_53);
or U1729 (N_1729,In_148,In_514);
and U1730 (N_1730,In_141,In_607);
and U1731 (N_1731,In_436,In_143);
and U1732 (N_1732,In_515,In_106);
and U1733 (N_1733,In_798,In_533);
or U1734 (N_1734,In_579,In_945);
nor U1735 (N_1735,In_279,In_508);
nand U1736 (N_1736,In_876,In_460);
nand U1737 (N_1737,In_252,In_516);
or U1738 (N_1738,In_749,In_335);
nor U1739 (N_1739,In_961,In_353);
xor U1740 (N_1740,In_14,In_807);
nor U1741 (N_1741,In_153,In_572);
or U1742 (N_1742,In_971,In_612);
xor U1743 (N_1743,In_894,In_282);
or U1744 (N_1744,In_234,In_59);
or U1745 (N_1745,In_20,In_834);
nand U1746 (N_1746,In_371,In_301);
nor U1747 (N_1747,In_208,In_539);
or U1748 (N_1748,In_403,In_805);
nor U1749 (N_1749,In_852,In_352);
xor U1750 (N_1750,In_131,In_427);
nand U1751 (N_1751,In_160,In_146);
nand U1752 (N_1752,In_507,In_101);
or U1753 (N_1753,In_803,In_346);
nand U1754 (N_1754,In_21,In_621);
nor U1755 (N_1755,In_15,In_654);
nand U1756 (N_1756,In_212,In_657);
and U1757 (N_1757,In_425,In_251);
nor U1758 (N_1758,In_240,In_252);
xnor U1759 (N_1759,In_843,In_615);
nor U1760 (N_1760,In_368,In_924);
and U1761 (N_1761,In_575,In_417);
nor U1762 (N_1762,In_17,In_873);
xor U1763 (N_1763,In_873,In_519);
and U1764 (N_1764,In_345,In_182);
or U1765 (N_1765,In_658,In_793);
and U1766 (N_1766,In_834,In_442);
nor U1767 (N_1767,In_587,In_676);
nor U1768 (N_1768,In_294,In_44);
nand U1769 (N_1769,In_225,In_820);
and U1770 (N_1770,In_970,In_413);
nor U1771 (N_1771,In_818,In_4);
nand U1772 (N_1772,In_227,In_805);
or U1773 (N_1773,In_375,In_393);
nor U1774 (N_1774,In_759,In_187);
nor U1775 (N_1775,In_546,In_521);
xnor U1776 (N_1776,In_37,In_40);
or U1777 (N_1777,In_506,In_908);
nor U1778 (N_1778,In_681,In_835);
nand U1779 (N_1779,In_31,In_495);
nor U1780 (N_1780,In_777,In_306);
nor U1781 (N_1781,In_855,In_559);
nor U1782 (N_1782,In_182,In_53);
and U1783 (N_1783,In_965,In_698);
nor U1784 (N_1784,In_494,In_304);
or U1785 (N_1785,In_882,In_153);
or U1786 (N_1786,In_105,In_312);
nand U1787 (N_1787,In_376,In_200);
nor U1788 (N_1788,In_140,In_786);
and U1789 (N_1789,In_843,In_988);
and U1790 (N_1790,In_212,In_331);
nor U1791 (N_1791,In_567,In_891);
nor U1792 (N_1792,In_666,In_656);
or U1793 (N_1793,In_777,In_447);
nor U1794 (N_1794,In_569,In_464);
and U1795 (N_1795,In_362,In_718);
and U1796 (N_1796,In_280,In_853);
xnor U1797 (N_1797,In_456,In_330);
nand U1798 (N_1798,In_955,In_125);
nand U1799 (N_1799,In_651,In_295);
nor U1800 (N_1800,In_158,In_446);
nor U1801 (N_1801,In_197,In_289);
and U1802 (N_1802,In_729,In_430);
nand U1803 (N_1803,In_601,In_78);
xnor U1804 (N_1804,In_401,In_105);
nand U1805 (N_1805,In_941,In_897);
nor U1806 (N_1806,In_593,In_62);
nor U1807 (N_1807,In_479,In_901);
or U1808 (N_1808,In_426,In_743);
nand U1809 (N_1809,In_472,In_150);
and U1810 (N_1810,In_809,In_68);
and U1811 (N_1811,In_48,In_716);
nand U1812 (N_1812,In_327,In_754);
or U1813 (N_1813,In_338,In_605);
or U1814 (N_1814,In_583,In_222);
nor U1815 (N_1815,In_690,In_41);
nor U1816 (N_1816,In_47,In_614);
nor U1817 (N_1817,In_79,In_39);
xnor U1818 (N_1818,In_671,In_754);
nand U1819 (N_1819,In_602,In_396);
xor U1820 (N_1820,In_163,In_945);
xnor U1821 (N_1821,In_924,In_936);
and U1822 (N_1822,In_641,In_888);
and U1823 (N_1823,In_931,In_972);
and U1824 (N_1824,In_363,In_225);
nand U1825 (N_1825,In_641,In_909);
xor U1826 (N_1826,In_826,In_384);
or U1827 (N_1827,In_579,In_686);
nor U1828 (N_1828,In_327,In_577);
nand U1829 (N_1829,In_275,In_857);
nor U1830 (N_1830,In_269,In_493);
or U1831 (N_1831,In_36,In_643);
and U1832 (N_1832,In_568,In_938);
nor U1833 (N_1833,In_151,In_370);
nand U1834 (N_1834,In_342,In_893);
nand U1835 (N_1835,In_576,In_434);
and U1836 (N_1836,In_248,In_942);
nand U1837 (N_1837,In_724,In_567);
nor U1838 (N_1838,In_514,In_884);
xnor U1839 (N_1839,In_384,In_56);
nand U1840 (N_1840,In_172,In_15);
and U1841 (N_1841,In_97,In_768);
and U1842 (N_1842,In_243,In_117);
and U1843 (N_1843,In_596,In_443);
and U1844 (N_1844,In_740,In_488);
or U1845 (N_1845,In_45,In_851);
and U1846 (N_1846,In_952,In_917);
nor U1847 (N_1847,In_974,In_548);
or U1848 (N_1848,In_534,In_772);
or U1849 (N_1849,In_624,In_274);
xnor U1850 (N_1850,In_999,In_690);
nand U1851 (N_1851,In_871,In_571);
nand U1852 (N_1852,In_128,In_830);
and U1853 (N_1853,In_811,In_132);
nor U1854 (N_1854,In_465,In_988);
or U1855 (N_1855,In_43,In_583);
nand U1856 (N_1856,In_218,In_700);
nor U1857 (N_1857,In_701,In_821);
nand U1858 (N_1858,In_557,In_743);
xor U1859 (N_1859,In_831,In_145);
nor U1860 (N_1860,In_746,In_654);
nand U1861 (N_1861,In_142,In_369);
nand U1862 (N_1862,In_305,In_343);
or U1863 (N_1863,In_555,In_170);
or U1864 (N_1864,In_154,In_430);
nor U1865 (N_1865,In_427,In_966);
or U1866 (N_1866,In_423,In_123);
nand U1867 (N_1867,In_475,In_477);
nor U1868 (N_1868,In_244,In_670);
nor U1869 (N_1869,In_932,In_123);
nor U1870 (N_1870,In_208,In_128);
xor U1871 (N_1871,In_699,In_107);
nor U1872 (N_1872,In_177,In_117);
and U1873 (N_1873,In_156,In_488);
xnor U1874 (N_1874,In_206,In_440);
and U1875 (N_1875,In_427,In_51);
nor U1876 (N_1876,In_523,In_590);
nand U1877 (N_1877,In_574,In_515);
and U1878 (N_1878,In_393,In_654);
and U1879 (N_1879,In_681,In_526);
or U1880 (N_1880,In_532,In_219);
nand U1881 (N_1881,In_346,In_797);
nand U1882 (N_1882,In_407,In_584);
and U1883 (N_1883,In_56,In_978);
nor U1884 (N_1884,In_492,In_8);
nand U1885 (N_1885,In_664,In_129);
or U1886 (N_1886,In_207,In_735);
nand U1887 (N_1887,In_408,In_450);
nor U1888 (N_1888,In_317,In_473);
or U1889 (N_1889,In_685,In_510);
and U1890 (N_1890,In_559,In_430);
and U1891 (N_1891,In_405,In_389);
xor U1892 (N_1892,In_769,In_730);
and U1893 (N_1893,In_371,In_620);
nor U1894 (N_1894,In_732,In_852);
nor U1895 (N_1895,In_771,In_449);
and U1896 (N_1896,In_695,In_616);
xor U1897 (N_1897,In_339,In_431);
or U1898 (N_1898,In_826,In_907);
nor U1899 (N_1899,In_194,In_783);
nor U1900 (N_1900,In_66,In_650);
and U1901 (N_1901,In_930,In_186);
xnor U1902 (N_1902,In_553,In_378);
nor U1903 (N_1903,In_399,In_21);
nand U1904 (N_1904,In_701,In_912);
and U1905 (N_1905,In_540,In_805);
nand U1906 (N_1906,In_80,In_552);
xor U1907 (N_1907,In_874,In_767);
or U1908 (N_1908,In_54,In_418);
xor U1909 (N_1909,In_767,In_305);
nor U1910 (N_1910,In_394,In_875);
xor U1911 (N_1911,In_29,In_455);
nand U1912 (N_1912,In_477,In_325);
or U1913 (N_1913,In_432,In_874);
or U1914 (N_1914,In_111,In_548);
nand U1915 (N_1915,In_467,In_996);
or U1916 (N_1916,In_737,In_276);
or U1917 (N_1917,In_983,In_550);
nor U1918 (N_1918,In_178,In_49);
nand U1919 (N_1919,In_457,In_653);
and U1920 (N_1920,In_61,In_592);
xor U1921 (N_1921,In_853,In_711);
nor U1922 (N_1922,In_985,In_243);
nand U1923 (N_1923,In_802,In_907);
or U1924 (N_1924,In_147,In_102);
xnor U1925 (N_1925,In_88,In_568);
and U1926 (N_1926,In_114,In_212);
and U1927 (N_1927,In_168,In_844);
or U1928 (N_1928,In_679,In_523);
xor U1929 (N_1929,In_739,In_98);
xnor U1930 (N_1930,In_980,In_237);
or U1931 (N_1931,In_607,In_251);
and U1932 (N_1932,In_687,In_938);
nand U1933 (N_1933,In_637,In_514);
nand U1934 (N_1934,In_449,In_742);
or U1935 (N_1935,In_677,In_173);
nor U1936 (N_1936,In_270,In_126);
nand U1937 (N_1937,In_893,In_516);
and U1938 (N_1938,In_58,In_203);
nand U1939 (N_1939,In_483,In_222);
nor U1940 (N_1940,In_440,In_442);
nand U1941 (N_1941,In_655,In_105);
xnor U1942 (N_1942,In_93,In_885);
and U1943 (N_1943,In_282,In_260);
nor U1944 (N_1944,In_551,In_431);
nand U1945 (N_1945,In_6,In_574);
nand U1946 (N_1946,In_956,In_267);
nor U1947 (N_1947,In_868,In_455);
and U1948 (N_1948,In_699,In_65);
nor U1949 (N_1949,In_283,In_684);
and U1950 (N_1950,In_750,In_208);
or U1951 (N_1951,In_1,In_899);
nor U1952 (N_1952,In_688,In_330);
nand U1953 (N_1953,In_429,In_392);
or U1954 (N_1954,In_292,In_725);
and U1955 (N_1955,In_545,In_948);
nand U1956 (N_1956,In_460,In_894);
xor U1957 (N_1957,In_865,In_626);
or U1958 (N_1958,In_878,In_213);
nor U1959 (N_1959,In_401,In_520);
nor U1960 (N_1960,In_294,In_408);
nand U1961 (N_1961,In_741,In_77);
nand U1962 (N_1962,In_880,In_777);
nand U1963 (N_1963,In_241,In_286);
xor U1964 (N_1964,In_416,In_504);
nor U1965 (N_1965,In_883,In_56);
nor U1966 (N_1966,In_834,In_449);
and U1967 (N_1967,In_781,In_310);
nor U1968 (N_1968,In_815,In_523);
and U1969 (N_1969,In_139,In_355);
nor U1970 (N_1970,In_498,In_335);
nand U1971 (N_1971,In_303,In_44);
or U1972 (N_1972,In_387,In_705);
nand U1973 (N_1973,In_460,In_456);
nand U1974 (N_1974,In_388,In_918);
nand U1975 (N_1975,In_316,In_614);
and U1976 (N_1976,In_725,In_26);
nor U1977 (N_1977,In_303,In_254);
nor U1978 (N_1978,In_979,In_269);
and U1979 (N_1979,In_350,In_727);
nor U1980 (N_1980,In_995,In_216);
nor U1981 (N_1981,In_594,In_346);
or U1982 (N_1982,In_832,In_372);
or U1983 (N_1983,In_989,In_127);
nand U1984 (N_1984,In_966,In_931);
xnor U1985 (N_1985,In_794,In_680);
or U1986 (N_1986,In_975,In_15);
and U1987 (N_1987,In_748,In_871);
nor U1988 (N_1988,In_647,In_508);
and U1989 (N_1989,In_798,In_943);
nor U1990 (N_1990,In_337,In_635);
or U1991 (N_1991,In_268,In_197);
and U1992 (N_1992,In_851,In_654);
nand U1993 (N_1993,In_416,In_528);
or U1994 (N_1994,In_511,In_113);
and U1995 (N_1995,In_241,In_23);
nor U1996 (N_1996,In_224,In_911);
and U1997 (N_1997,In_914,In_348);
and U1998 (N_1998,In_764,In_478);
nand U1999 (N_1999,In_137,In_978);
xor U2000 (N_2000,In_910,In_181);
nand U2001 (N_2001,In_574,In_570);
nor U2002 (N_2002,In_533,In_268);
nand U2003 (N_2003,In_720,In_216);
xor U2004 (N_2004,In_371,In_630);
nor U2005 (N_2005,In_276,In_11);
xor U2006 (N_2006,In_196,In_927);
nor U2007 (N_2007,In_341,In_385);
nor U2008 (N_2008,In_727,In_861);
and U2009 (N_2009,In_99,In_894);
nor U2010 (N_2010,In_791,In_863);
and U2011 (N_2011,In_184,In_672);
and U2012 (N_2012,In_574,In_854);
and U2013 (N_2013,In_623,In_718);
nand U2014 (N_2014,In_684,In_401);
nor U2015 (N_2015,In_602,In_836);
nand U2016 (N_2016,In_283,In_875);
or U2017 (N_2017,In_276,In_180);
nor U2018 (N_2018,In_168,In_141);
nand U2019 (N_2019,In_302,In_867);
and U2020 (N_2020,In_791,In_543);
and U2021 (N_2021,In_866,In_853);
nor U2022 (N_2022,In_767,In_558);
or U2023 (N_2023,In_218,In_571);
or U2024 (N_2024,In_960,In_652);
or U2025 (N_2025,In_888,In_827);
and U2026 (N_2026,In_312,In_704);
nor U2027 (N_2027,In_461,In_301);
and U2028 (N_2028,In_294,In_632);
or U2029 (N_2029,In_760,In_489);
nand U2030 (N_2030,In_735,In_129);
nor U2031 (N_2031,In_258,In_985);
nor U2032 (N_2032,In_333,In_928);
and U2033 (N_2033,In_175,In_643);
nor U2034 (N_2034,In_406,In_288);
nand U2035 (N_2035,In_442,In_689);
or U2036 (N_2036,In_229,In_238);
or U2037 (N_2037,In_17,In_534);
or U2038 (N_2038,In_409,In_519);
and U2039 (N_2039,In_653,In_412);
or U2040 (N_2040,In_416,In_115);
or U2041 (N_2041,In_377,In_961);
xnor U2042 (N_2042,In_274,In_696);
or U2043 (N_2043,In_856,In_355);
and U2044 (N_2044,In_7,In_706);
nor U2045 (N_2045,In_298,In_3);
and U2046 (N_2046,In_655,In_451);
and U2047 (N_2047,In_935,In_673);
nor U2048 (N_2048,In_916,In_507);
nor U2049 (N_2049,In_584,In_350);
nor U2050 (N_2050,In_438,In_484);
nor U2051 (N_2051,In_468,In_763);
and U2052 (N_2052,In_386,In_836);
nand U2053 (N_2053,In_399,In_572);
and U2054 (N_2054,In_713,In_466);
nand U2055 (N_2055,In_944,In_895);
and U2056 (N_2056,In_644,In_29);
and U2057 (N_2057,In_117,In_773);
nor U2058 (N_2058,In_623,In_92);
or U2059 (N_2059,In_767,In_704);
and U2060 (N_2060,In_649,In_620);
nand U2061 (N_2061,In_333,In_317);
nor U2062 (N_2062,In_209,In_829);
nand U2063 (N_2063,In_574,In_681);
and U2064 (N_2064,In_694,In_916);
nand U2065 (N_2065,In_917,In_131);
or U2066 (N_2066,In_837,In_195);
nor U2067 (N_2067,In_135,In_212);
xnor U2068 (N_2068,In_868,In_306);
or U2069 (N_2069,In_621,In_737);
xor U2070 (N_2070,In_962,In_65);
xnor U2071 (N_2071,In_457,In_709);
and U2072 (N_2072,In_920,In_890);
xnor U2073 (N_2073,In_930,In_223);
xor U2074 (N_2074,In_243,In_46);
nor U2075 (N_2075,In_656,In_149);
nor U2076 (N_2076,In_613,In_967);
or U2077 (N_2077,In_176,In_615);
xnor U2078 (N_2078,In_214,In_99);
or U2079 (N_2079,In_991,In_515);
or U2080 (N_2080,In_243,In_440);
nor U2081 (N_2081,In_72,In_829);
or U2082 (N_2082,In_388,In_696);
nor U2083 (N_2083,In_283,In_422);
and U2084 (N_2084,In_331,In_862);
or U2085 (N_2085,In_666,In_863);
or U2086 (N_2086,In_789,In_183);
and U2087 (N_2087,In_162,In_648);
nor U2088 (N_2088,In_279,In_684);
nand U2089 (N_2089,In_221,In_580);
nor U2090 (N_2090,In_395,In_599);
or U2091 (N_2091,In_211,In_960);
nand U2092 (N_2092,In_388,In_704);
and U2093 (N_2093,In_560,In_671);
or U2094 (N_2094,In_513,In_26);
nand U2095 (N_2095,In_759,In_799);
or U2096 (N_2096,In_710,In_935);
and U2097 (N_2097,In_419,In_148);
nand U2098 (N_2098,In_740,In_618);
xor U2099 (N_2099,In_794,In_497);
or U2100 (N_2100,In_142,In_136);
nand U2101 (N_2101,In_239,In_322);
or U2102 (N_2102,In_807,In_16);
nor U2103 (N_2103,In_959,In_783);
nand U2104 (N_2104,In_863,In_618);
nand U2105 (N_2105,In_167,In_551);
nor U2106 (N_2106,In_394,In_786);
xnor U2107 (N_2107,In_307,In_246);
xnor U2108 (N_2108,In_75,In_148);
or U2109 (N_2109,In_246,In_160);
and U2110 (N_2110,In_674,In_34);
nor U2111 (N_2111,In_981,In_137);
and U2112 (N_2112,In_899,In_480);
nor U2113 (N_2113,In_48,In_726);
xor U2114 (N_2114,In_542,In_131);
nor U2115 (N_2115,In_159,In_183);
nor U2116 (N_2116,In_886,In_133);
and U2117 (N_2117,In_131,In_270);
nand U2118 (N_2118,In_164,In_538);
nor U2119 (N_2119,In_577,In_815);
nor U2120 (N_2120,In_640,In_642);
or U2121 (N_2121,In_59,In_975);
nor U2122 (N_2122,In_873,In_312);
nand U2123 (N_2123,In_922,In_255);
nor U2124 (N_2124,In_341,In_592);
and U2125 (N_2125,In_672,In_213);
nor U2126 (N_2126,In_22,In_873);
or U2127 (N_2127,In_282,In_337);
nor U2128 (N_2128,In_190,In_928);
nand U2129 (N_2129,In_64,In_924);
or U2130 (N_2130,In_329,In_871);
nor U2131 (N_2131,In_348,In_182);
nor U2132 (N_2132,In_428,In_489);
nor U2133 (N_2133,In_863,In_644);
nand U2134 (N_2134,In_970,In_118);
nor U2135 (N_2135,In_818,In_18);
xor U2136 (N_2136,In_7,In_518);
nand U2137 (N_2137,In_825,In_697);
and U2138 (N_2138,In_469,In_677);
nor U2139 (N_2139,In_932,In_315);
or U2140 (N_2140,In_44,In_54);
or U2141 (N_2141,In_703,In_768);
and U2142 (N_2142,In_508,In_781);
nor U2143 (N_2143,In_489,In_154);
nand U2144 (N_2144,In_721,In_970);
and U2145 (N_2145,In_720,In_163);
nor U2146 (N_2146,In_351,In_455);
nor U2147 (N_2147,In_840,In_35);
or U2148 (N_2148,In_896,In_221);
nand U2149 (N_2149,In_587,In_415);
nor U2150 (N_2150,In_364,In_531);
nand U2151 (N_2151,In_544,In_618);
nand U2152 (N_2152,In_878,In_875);
or U2153 (N_2153,In_811,In_39);
and U2154 (N_2154,In_337,In_820);
nand U2155 (N_2155,In_504,In_276);
or U2156 (N_2156,In_196,In_504);
and U2157 (N_2157,In_310,In_653);
and U2158 (N_2158,In_310,In_727);
nand U2159 (N_2159,In_209,In_941);
and U2160 (N_2160,In_539,In_708);
or U2161 (N_2161,In_688,In_528);
nand U2162 (N_2162,In_291,In_313);
and U2163 (N_2163,In_310,In_556);
and U2164 (N_2164,In_701,In_958);
or U2165 (N_2165,In_204,In_511);
or U2166 (N_2166,In_524,In_410);
xor U2167 (N_2167,In_126,In_539);
and U2168 (N_2168,In_4,In_214);
nand U2169 (N_2169,In_111,In_686);
nor U2170 (N_2170,In_632,In_164);
nand U2171 (N_2171,In_756,In_336);
nand U2172 (N_2172,In_850,In_877);
xor U2173 (N_2173,In_127,In_825);
nand U2174 (N_2174,In_177,In_162);
and U2175 (N_2175,In_397,In_314);
xor U2176 (N_2176,In_57,In_940);
nand U2177 (N_2177,In_117,In_835);
and U2178 (N_2178,In_103,In_240);
or U2179 (N_2179,In_682,In_303);
or U2180 (N_2180,In_28,In_605);
nand U2181 (N_2181,In_349,In_244);
and U2182 (N_2182,In_116,In_950);
and U2183 (N_2183,In_700,In_0);
xor U2184 (N_2184,In_979,In_949);
xnor U2185 (N_2185,In_635,In_100);
nor U2186 (N_2186,In_348,In_545);
or U2187 (N_2187,In_794,In_732);
and U2188 (N_2188,In_502,In_348);
and U2189 (N_2189,In_752,In_250);
xnor U2190 (N_2190,In_310,In_369);
nor U2191 (N_2191,In_688,In_863);
nor U2192 (N_2192,In_660,In_76);
nand U2193 (N_2193,In_799,In_25);
nor U2194 (N_2194,In_674,In_829);
and U2195 (N_2195,In_248,In_50);
nor U2196 (N_2196,In_477,In_20);
or U2197 (N_2197,In_253,In_128);
and U2198 (N_2198,In_250,In_714);
nand U2199 (N_2199,In_790,In_997);
nand U2200 (N_2200,In_234,In_437);
and U2201 (N_2201,In_816,In_406);
or U2202 (N_2202,In_635,In_529);
and U2203 (N_2203,In_455,In_626);
nand U2204 (N_2204,In_393,In_439);
nand U2205 (N_2205,In_824,In_209);
and U2206 (N_2206,In_339,In_743);
nand U2207 (N_2207,In_291,In_90);
nor U2208 (N_2208,In_479,In_634);
and U2209 (N_2209,In_499,In_665);
or U2210 (N_2210,In_257,In_126);
nor U2211 (N_2211,In_973,In_173);
and U2212 (N_2212,In_281,In_294);
nand U2213 (N_2213,In_936,In_422);
nand U2214 (N_2214,In_980,In_216);
nand U2215 (N_2215,In_602,In_674);
nand U2216 (N_2216,In_2,In_304);
nand U2217 (N_2217,In_498,In_653);
nand U2218 (N_2218,In_206,In_727);
nor U2219 (N_2219,In_760,In_716);
nor U2220 (N_2220,In_817,In_211);
nor U2221 (N_2221,In_64,In_660);
nor U2222 (N_2222,In_946,In_715);
nand U2223 (N_2223,In_19,In_726);
nand U2224 (N_2224,In_397,In_641);
or U2225 (N_2225,In_796,In_632);
nor U2226 (N_2226,In_435,In_993);
and U2227 (N_2227,In_879,In_370);
nand U2228 (N_2228,In_151,In_441);
and U2229 (N_2229,In_178,In_803);
or U2230 (N_2230,In_830,In_58);
nor U2231 (N_2231,In_979,In_239);
xor U2232 (N_2232,In_115,In_51);
nand U2233 (N_2233,In_38,In_778);
and U2234 (N_2234,In_731,In_481);
nand U2235 (N_2235,In_776,In_57);
and U2236 (N_2236,In_159,In_268);
or U2237 (N_2237,In_974,In_358);
or U2238 (N_2238,In_570,In_131);
and U2239 (N_2239,In_724,In_439);
or U2240 (N_2240,In_678,In_734);
and U2241 (N_2241,In_55,In_140);
nor U2242 (N_2242,In_516,In_691);
nor U2243 (N_2243,In_594,In_387);
and U2244 (N_2244,In_961,In_655);
and U2245 (N_2245,In_669,In_421);
nor U2246 (N_2246,In_807,In_810);
and U2247 (N_2247,In_279,In_748);
nor U2248 (N_2248,In_817,In_121);
and U2249 (N_2249,In_733,In_462);
nand U2250 (N_2250,In_57,In_235);
nor U2251 (N_2251,In_124,In_334);
or U2252 (N_2252,In_136,In_131);
and U2253 (N_2253,In_954,In_611);
or U2254 (N_2254,In_445,In_321);
or U2255 (N_2255,In_140,In_558);
and U2256 (N_2256,In_605,In_356);
and U2257 (N_2257,In_360,In_677);
xor U2258 (N_2258,In_70,In_623);
nor U2259 (N_2259,In_273,In_718);
and U2260 (N_2260,In_650,In_207);
xor U2261 (N_2261,In_627,In_43);
xor U2262 (N_2262,In_60,In_7);
xor U2263 (N_2263,In_687,In_771);
xor U2264 (N_2264,In_634,In_157);
or U2265 (N_2265,In_733,In_866);
nor U2266 (N_2266,In_526,In_315);
nor U2267 (N_2267,In_792,In_322);
nand U2268 (N_2268,In_977,In_729);
or U2269 (N_2269,In_603,In_879);
xor U2270 (N_2270,In_124,In_927);
and U2271 (N_2271,In_291,In_800);
nor U2272 (N_2272,In_447,In_897);
and U2273 (N_2273,In_918,In_446);
or U2274 (N_2274,In_40,In_654);
nor U2275 (N_2275,In_581,In_406);
nand U2276 (N_2276,In_42,In_115);
and U2277 (N_2277,In_712,In_666);
nor U2278 (N_2278,In_112,In_22);
nor U2279 (N_2279,In_387,In_763);
nor U2280 (N_2280,In_951,In_11);
nor U2281 (N_2281,In_278,In_705);
and U2282 (N_2282,In_537,In_240);
or U2283 (N_2283,In_425,In_267);
nor U2284 (N_2284,In_324,In_605);
nor U2285 (N_2285,In_934,In_401);
and U2286 (N_2286,In_413,In_435);
and U2287 (N_2287,In_988,In_44);
nand U2288 (N_2288,In_689,In_849);
nor U2289 (N_2289,In_921,In_44);
or U2290 (N_2290,In_41,In_64);
and U2291 (N_2291,In_506,In_937);
nor U2292 (N_2292,In_337,In_622);
nand U2293 (N_2293,In_427,In_298);
nand U2294 (N_2294,In_720,In_497);
nand U2295 (N_2295,In_588,In_318);
and U2296 (N_2296,In_930,In_870);
nor U2297 (N_2297,In_925,In_553);
nor U2298 (N_2298,In_437,In_341);
nand U2299 (N_2299,In_506,In_37);
nor U2300 (N_2300,In_890,In_452);
nand U2301 (N_2301,In_366,In_999);
or U2302 (N_2302,In_549,In_80);
or U2303 (N_2303,In_867,In_907);
nand U2304 (N_2304,In_789,In_757);
nand U2305 (N_2305,In_901,In_505);
or U2306 (N_2306,In_953,In_733);
and U2307 (N_2307,In_830,In_661);
and U2308 (N_2308,In_446,In_215);
nand U2309 (N_2309,In_790,In_497);
and U2310 (N_2310,In_995,In_642);
xnor U2311 (N_2311,In_746,In_545);
nor U2312 (N_2312,In_425,In_893);
nand U2313 (N_2313,In_851,In_791);
or U2314 (N_2314,In_822,In_176);
xor U2315 (N_2315,In_106,In_401);
nand U2316 (N_2316,In_548,In_922);
nand U2317 (N_2317,In_698,In_583);
and U2318 (N_2318,In_16,In_687);
xor U2319 (N_2319,In_627,In_628);
nand U2320 (N_2320,In_229,In_603);
or U2321 (N_2321,In_921,In_451);
xor U2322 (N_2322,In_455,In_939);
nor U2323 (N_2323,In_169,In_103);
and U2324 (N_2324,In_591,In_9);
nor U2325 (N_2325,In_116,In_765);
nand U2326 (N_2326,In_835,In_894);
nor U2327 (N_2327,In_246,In_120);
or U2328 (N_2328,In_834,In_807);
and U2329 (N_2329,In_946,In_524);
xor U2330 (N_2330,In_577,In_605);
xor U2331 (N_2331,In_177,In_206);
nor U2332 (N_2332,In_645,In_425);
xnor U2333 (N_2333,In_503,In_957);
nand U2334 (N_2334,In_610,In_42);
or U2335 (N_2335,In_565,In_379);
and U2336 (N_2336,In_44,In_356);
nand U2337 (N_2337,In_940,In_280);
and U2338 (N_2338,In_393,In_848);
and U2339 (N_2339,In_507,In_824);
and U2340 (N_2340,In_209,In_193);
nor U2341 (N_2341,In_760,In_787);
xor U2342 (N_2342,In_496,In_993);
nand U2343 (N_2343,In_939,In_387);
and U2344 (N_2344,In_531,In_783);
nand U2345 (N_2345,In_635,In_920);
nand U2346 (N_2346,In_82,In_968);
and U2347 (N_2347,In_893,In_580);
and U2348 (N_2348,In_687,In_488);
nor U2349 (N_2349,In_69,In_269);
nand U2350 (N_2350,In_48,In_354);
nor U2351 (N_2351,In_976,In_469);
and U2352 (N_2352,In_412,In_576);
or U2353 (N_2353,In_151,In_6);
and U2354 (N_2354,In_600,In_461);
nand U2355 (N_2355,In_211,In_174);
or U2356 (N_2356,In_979,In_920);
or U2357 (N_2357,In_763,In_808);
and U2358 (N_2358,In_44,In_757);
or U2359 (N_2359,In_434,In_366);
nor U2360 (N_2360,In_785,In_700);
or U2361 (N_2361,In_658,In_612);
nor U2362 (N_2362,In_108,In_319);
nand U2363 (N_2363,In_507,In_352);
nand U2364 (N_2364,In_847,In_539);
nand U2365 (N_2365,In_726,In_370);
nand U2366 (N_2366,In_242,In_401);
nor U2367 (N_2367,In_976,In_30);
nand U2368 (N_2368,In_497,In_441);
nand U2369 (N_2369,In_770,In_540);
nand U2370 (N_2370,In_695,In_555);
nand U2371 (N_2371,In_716,In_898);
nor U2372 (N_2372,In_308,In_917);
or U2373 (N_2373,In_764,In_829);
nand U2374 (N_2374,In_125,In_268);
or U2375 (N_2375,In_463,In_974);
xor U2376 (N_2376,In_381,In_764);
or U2377 (N_2377,In_144,In_231);
or U2378 (N_2378,In_243,In_819);
nand U2379 (N_2379,In_148,In_471);
and U2380 (N_2380,In_672,In_900);
or U2381 (N_2381,In_328,In_918);
nor U2382 (N_2382,In_259,In_28);
or U2383 (N_2383,In_783,In_591);
xnor U2384 (N_2384,In_812,In_774);
xnor U2385 (N_2385,In_36,In_144);
nor U2386 (N_2386,In_410,In_352);
nand U2387 (N_2387,In_218,In_434);
or U2388 (N_2388,In_280,In_844);
and U2389 (N_2389,In_457,In_939);
xnor U2390 (N_2390,In_756,In_944);
nor U2391 (N_2391,In_748,In_469);
or U2392 (N_2392,In_716,In_783);
nand U2393 (N_2393,In_814,In_973);
nand U2394 (N_2394,In_455,In_531);
nor U2395 (N_2395,In_216,In_310);
or U2396 (N_2396,In_494,In_143);
nand U2397 (N_2397,In_486,In_346);
xnor U2398 (N_2398,In_939,In_561);
xnor U2399 (N_2399,In_725,In_895);
or U2400 (N_2400,In_959,In_134);
xor U2401 (N_2401,In_164,In_711);
nor U2402 (N_2402,In_517,In_572);
and U2403 (N_2403,In_461,In_754);
xnor U2404 (N_2404,In_763,In_590);
nand U2405 (N_2405,In_366,In_487);
or U2406 (N_2406,In_938,In_133);
xor U2407 (N_2407,In_191,In_198);
nor U2408 (N_2408,In_250,In_813);
xnor U2409 (N_2409,In_616,In_867);
nand U2410 (N_2410,In_958,In_58);
or U2411 (N_2411,In_131,In_113);
or U2412 (N_2412,In_580,In_21);
and U2413 (N_2413,In_379,In_366);
and U2414 (N_2414,In_518,In_850);
or U2415 (N_2415,In_922,In_487);
and U2416 (N_2416,In_728,In_322);
and U2417 (N_2417,In_314,In_309);
nor U2418 (N_2418,In_135,In_484);
or U2419 (N_2419,In_299,In_779);
or U2420 (N_2420,In_840,In_796);
and U2421 (N_2421,In_369,In_926);
or U2422 (N_2422,In_558,In_590);
and U2423 (N_2423,In_545,In_728);
and U2424 (N_2424,In_596,In_567);
nand U2425 (N_2425,In_319,In_874);
or U2426 (N_2426,In_145,In_228);
or U2427 (N_2427,In_685,In_626);
nor U2428 (N_2428,In_26,In_842);
xnor U2429 (N_2429,In_971,In_817);
nor U2430 (N_2430,In_328,In_365);
and U2431 (N_2431,In_618,In_883);
nor U2432 (N_2432,In_738,In_710);
nor U2433 (N_2433,In_770,In_943);
or U2434 (N_2434,In_194,In_384);
or U2435 (N_2435,In_430,In_959);
xnor U2436 (N_2436,In_750,In_288);
and U2437 (N_2437,In_85,In_433);
nand U2438 (N_2438,In_719,In_665);
and U2439 (N_2439,In_523,In_541);
or U2440 (N_2440,In_384,In_255);
or U2441 (N_2441,In_142,In_292);
and U2442 (N_2442,In_460,In_952);
nand U2443 (N_2443,In_993,In_657);
and U2444 (N_2444,In_275,In_608);
xor U2445 (N_2445,In_574,In_528);
nand U2446 (N_2446,In_706,In_274);
and U2447 (N_2447,In_628,In_909);
or U2448 (N_2448,In_922,In_833);
nand U2449 (N_2449,In_484,In_83);
or U2450 (N_2450,In_235,In_526);
nor U2451 (N_2451,In_833,In_130);
or U2452 (N_2452,In_79,In_589);
and U2453 (N_2453,In_54,In_168);
or U2454 (N_2454,In_294,In_987);
nand U2455 (N_2455,In_957,In_894);
nor U2456 (N_2456,In_867,In_597);
xnor U2457 (N_2457,In_29,In_487);
or U2458 (N_2458,In_198,In_993);
nor U2459 (N_2459,In_57,In_498);
and U2460 (N_2460,In_676,In_483);
nand U2461 (N_2461,In_763,In_441);
nor U2462 (N_2462,In_478,In_443);
nor U2463 (N_2463,In_751,In_983);
and U2464 (N_2464,In_154,In_431);
nor U2465 (N_2465,In_69,In_742);
or U2466 (N_2466,In_167,In_522);
or U2467 (N_2467,In_970,In_606);
nor U2468 (N_2468,In_844,In_482);
and U2469 (N_2469,In_448,In_226);
nand U2470 (N_2470,In_925,In_649);
or U2471 (N_2471,In_298,In_8);
nor U2472 (N_2472,In_106,In_223);
nor U2473 (N_2473,In_943,In_136);
or U2474 (N_2474,In_649,In_102);
xnor U2475 (N_2475,In_914,In_818);
nor U2476 (N_2476,In_180,In_328);
and U2477 (N_2477,In_389,In_459);
or U2478 (N_2478,In_601,In_104);
and U2479 (N_2479,In_635,In_130);
and U2480 (N_2480,In_522,In_838);
nand U2481 (N_2481,In_236,In_285);
or U2482 (N_2482,In_752,In_712);
nand U2483 (N_2483,In_512,In_168);
or U2484 (N_2484,In_774,In_31);
nor U2485 (N_2485,In_258,In_289);
nand U2486 (N_2486,In_833,In_197);
and U2487 (N_2487,In_928,In_91);
and U2488 (N_2488,In_352,In_917);
xnor U2489 (N_2489,In_348,In_526);
or U2490 (N_2490,In_373,In_76);
xor U2491 (N_2491,In_293,In_752);
or U2492 (N_2492,In_443,In_780);
and U2493 (N_2493,In_388,In_583);
or U2494 (N_2494,In_266,In_606);
or U2495 (N_2495,In_835,In_565);
nor U2496 (N_2496,In_544,In_27);
and U2497 (N_2497,In_727,In_910);
nor U2498 (N_2498,In_231,In_966);
nand U2499 (N_2499,In_610,In_601);
nor U2500 (N_2500,N_1035,N_304);
and U2501 (N_2501,N_279,N_1551);
and U2502 (N_2502,N_1932,N_2231);
nand U2503 (N_2503,N_374,N_1131);
or U2504 (N_2504,N_765,N_1924);
or U2505 (N_2505,N_1639,N_2145);
nand U2506 (N_2506,N_1589,N_315);
and U2507 (N_2507,N_2134,N_121);
and U2508 (N_2508,N_174,N_1797);
and U2509 (N_2509,N_2194,N_2291);
nor U2510 (N_2510,N_1356,N_2156);
or U2511 (N_2511,N_836,N_2312);
xor U2512 (N_2512,N_2416,N_515);
nand U2513 (N_2513,N_1312,N_827);
nor U2514 (N_2514,N_1740,N_23);
and U2515 (N_2515,N_1898,N_2111);
nand U2516 (N_2516,N_2252,N_166);
or U2517 (N_2517,N_848,N_1439);
and U2518 (N_2518,N_2473,N_1960);
nor U2519 (N_2519,N_197,N_669);
or U2520 (N_2520,N_1665,N_777);
and U2521 (N_2521,N_118,N_1552);
or U2522 (N_2522,N_2214,N_2016);
and U2523 (N_2523,N_1805,N_1337);
nand U2524 (N_2524,N_957,N_668);
nand U2525 (N_2525,N_1204,N_821);
or U2526 (N_2526,N_1179,N_1223);
xnor U2527 (N_2527,N_2035,N_2201);
nand U2528 (N_2528,N_1994,N_400);
nor U2529 (N_2529,N_1432,N_794);
and U2530 (N_2530,N_1542,N_1486);
nand U2531 (N_2531,N_474,N_1592);
nand U2532 (N_2532,N_1902,N_1921);
xnor U2533 (N_2533,N_355,N_1111);
nand U2534 (N_2534,N_2485,N_226);
or U2535 (N_2535,N_1756,N_1662);
and U2536 (N_2536,N_2182,N_256);
nor U2537 (N_2537,N_886,N_1392);
nor U2538 (N_2538,N_1796,N_309);
and U2539 (N_2539,N_2043,N_2098);
or U2540 (N_2540,N_743,N_290);
or U2541 (N_2541,N_755,N_606);
or U2542 (N_2542,N_2386,N_1070);
and U2543 (N_2543,N_1858,N_543);
nor U2544 (N_2544,N_1832,N_787);
or U2545 (N_2545,N_1666,N_2398);
nand U2546 (N_2546,N_789,N_1144);
and U2547 (N_2547,N_806,N_181);
and U2548 (N_2548,N_225,N_776);
nand U2549 (N_2549,N_2345,N_1983);
or U2550 (N_2550,N_972,N_1352);
or U2551 (N_2551,N_641,N_2288);
nor U2552 (N_2552,N_2212,N_2074);
nand U2553 (N_2553,N_1955,N_237);
nor U2554 (N_2554,N_2334,N_546);
nor U2555 (N_2555,N_1928,N_522);
nand U2556 (N_2556,N_44,N_1804);
or U2557 (N_2557,N_1986,N_2122);
nand U2558 (N_2558,N_1140,N_1321);
nor U2559 (N_2559,N_1656,N_658);
nor U2560 (N_2560,N_2415,N_2441);
xnor U2561 (N_2561,N_343,N_2191);
nor U2562 (N_2562,N_215,N_1033);
xor U2563 (N_2563,N_1157,N_910);
xor U2564 (N_2564,N_2474,N_1807);
nor U2565 (N_2565,N_567,N_1276);
xnor U2566 (N_2566,N_754,N_1197);
or U2567 (N_2567,N_1692,N_357);
nor U2568 (N_2568,N_2299,N_407);
xor U2569 (N_2569,N_746,N_81);
and U2570 (N_2570,N_231,N_1774);
xnor U2571 (N_2571,N_1382,N_50);
nand U2572 (N_2572,N_1491,N_571);
nand U2573 (N_2573,N_2408,N_1930);
or U2574 (N_2574,N_459,N_1625);
xor U2575 (N_2575,N_2365,N_427);
and U2576 (N_2576,N_65,N_1926);
and U2577 (N_2577,N_1097,N_1202);
nand U2578 (N_2578,N_1121,N_2038);
and U2579 (N_2579,N_95,N_831);
nand U2580 (N_2580,N_1386,N_1046);
and U2581 (N_2581,N_2080,N_698);
and U2582 (N_2582,N_785,N_2263);
and U2583 (N_2583,N_1482,N_1596);
and U2584 (N_2584,N_1794,N_1091);
nor U2585 (N_2585,N_2301,N_490);
nor U2586 (N_2586,N_2149,N_2209);
or U2587 (N_2587,N_2010,N_2433);
nor U2588 (N_2588,N_2465,N_1430);
nor U2589 (N_2589,N_1328,N_1559);
or U2590 (N_2590,N_1823,N_1311);
or U2591 (N_2591,N_1350,N_2190);
and U2592 (N_2592,N_72,N_1273);
or U2593 (N_2593,N_704,N_1063);
or U2594 (N_2594,N_1998,N_69);
xor U2595 (N_2595,N_1168,N_1243);
or U2596 (N_2596,N_1113,N_987);
nand U2597 (N_2597,N_2259,N_507);
or U2598 (N_2598,N_1906,N_1899);
or U2599 (N_2599,N_501,N_1881);
nor U2600 (N_2600,N_210,N_291);
xor U2601 (N_2601,N_2014,N_274);
nor U2602 (N_2602,N_2118,N_707);
or U2603 (N_2603,N_676,N_112);
and U2604 (N_2604,N_2371,N_1484);
nor U2605 (N_2605,N_2022,N_1056);
xnor U2606 (N_2606,N_949,N_2174);
xor U2607 (N_2607,N_552,N_2113);
nor U2608 (N_2608,N_871,N_175);
nor U2609 (N_2609,N_1431,N_1198);
nor U2610 (N_2610,N_1762,N_563);
nor U2611 (N_2611,N_692,N_2112);
or U2612 (N_2612,N_865,N_298);
and U2613 (N_2613,N_1271,N_2409);
or U2614 (N_2614,N_113,N_127);
and U2615 (N_2615,N_1489,N_155);
nor U2616 (N_2616,N_1128,N_1866);
or U2617 (N_2617,N_598,N_832);
or U2618 (N_2618,N_1761,N_2);
nor U2619 (N_2619,N_2338,N_1241);
nor U2620 (N_2620,N_824,N_453);
nand U2621 (N_2621,N_1852,N_652);
or U2622 (N_2622,N_715,N_857);
nand U2623 (N_2623,N_570,N_240);
or U2624 (N_2624,N_450,N_2477);
nand U2625 (N_2625,N_491,N_2232);
and U2626 (N_2626,N_1323,N_2335);
nor U2627 (N_2627,N_1614,N_736);
xnor U2628 (N_2628,N_797,N_2105);
nand U2629 (N_2629,N_862,N_2411);
xnor U2630 (N_2630,N_2251,N_431);
or U2631 (N_2631,N_872,N_1057);
nor U2632 (N_2632,N_117,N_1936);
nand U2633 (N_2633,N_116,N_804);
nor U2634 (N_2634,N_1309,N_518);
or U2635 (N_2635,N_1478,N_275);
and U2636 (N_2636,N_2197,N_958);
and U2637 (N_2637,N_358,N_313);
nand U2638 (N_2638,N_1269,N_1218);
and U2639 (N_2639,N_2050,N_2308);
xnor U2640 (N_2640,N_2271,N_2225);
or U2641 (N_2641,N_1428,N_2123);
and U2642 (N_2642,N_426,N_1962);
nand U2643 (N_2643,N_1635,N_1836);
nor U2644 (N_2644,N_2330,N_554);
or U2645 (N_2645,N_247,N_205);
nor U2646 (N_2646,N_2213,N_741);
or U2647 (N_2647,N_901,N_1678);
nor U2648 (N_2648,N_2188,N_1905);
nand U2649 (N_2649,N_2374,N_1378);
and U2650 (N_2650,N_792,N_1690);
nand U2651 (N_2651,N_1909,N_525);
nor U2652 (N_2652,N_892,N_1401);
and U2653 (N_2653,N_1974,N_575);
and U2654 (N_2654,N_1588,N_2139);
and U2655 (N_2655,N_93,N_51);
nand U2656 (N_2656,N_1245,N_1904);
nor U2657 (N_2657,N_640,N_392);
or U2658 (N_2658,N_1353,N_1238);
nor U2659 (N_2659,N_869,N_1539);
nand U2660 (N_2660,N_562,N_389);
and U2661 (N_2661,N_2382,N_595);
xor U2662 (N_2662,N_1919,N_1730);
and U2663 (N_2663,N_1834,N_1498);
and U2664 (N_2664,N_145,N_2400);
or U2665 (N_2665,N_1845,N_967);
xnor U2666 (N_2666,N_941,N_1660);
nor U2667 (N_2667,N_1058,N_1525);
nand U2668 (N_2668,N_1390,N_1684);
and U2669 (N_2669,N_54,N_2006);
nand U2670 (N_2670,N_1615,N_721);
nor U2671 (N_2671,N_330,N_2119);
or U2672 (N_2672,N_1040,N_2096);
or U2673 (N_2673,N_2310,N_1739);
or U2674 (N_2674,N_1014,N_1863);
xnor U2675 (N_2675,N_216,N_1531);
and U2676 (N_2676,N_1536,N_2493);
and U2677 (N_2677,N_1800,N_608);
and U2678 (N_2678,N_504,N_1546);
and U2679 (N_2679,N_1130,N_904);
or U2680 (N_2680,N_2392,N_1059);
nand U2681 (N_2681,N_1585,N_1565);
or U2682 (N_2682,N_1791,N_1342);
and U2683 (N_2683,N_2205,N_691);
nor U2684 (N_2684,N_62,N_928);
and U2685 (N_2685,N_537,N_1150);
nor U2686 (N_2686,N_381,N_1544);
and U2687 (N_2687,N_284,N_73);
or U2688 (N_2688,N_1274,N_616);
nand U2689 (N_2689,N_918,N_295);
and U2690 (N_2690,N_2041,N_2053);
and U2691 (N_2691,N_1734,N_1122);
nand U2692 (N_2692,N_795,N_1013);
or U2693 (N_2693,N_913,N_206);
xor U2694 (N_2694,N_1418,N_2293);
nor U2695 (N_2695,N_1671,N_981);
nor U2696 (N_2696,N_1843,N_757);
and U2697 (N_2697,N_2475,N_2405);
or U2698 (N_2698,N_384,N_1997);
nor U2699 (N_2699,N_1383,N_2247);
and U2700 (N_2700,N_1976,N_218);
nand U2701 (N_2701,N_443,N_375);
nor U2702 (N_2702,N_276,N_961);
nor U2703 (N_2703,N_874,N_378);
or U2704 (N_2704,N_992,N_421);
and U2705 (N_2705,N_1950,N_14);
nor U2706 (N_2706,N_25,N_1492);
and U2707 (N_2707,N_1182,N_906);
xnor U2708 (N_2708,N_248,N_1951);
nand U2709 (N_2709,N_1763,N_1812);
xor U2710 (N_2710,N_633,N_1379);
nor U2711 (N_2711,N_1686,N_495);
nand U2712 (N_2712,N_2381,N_1853);
nand U2713 (N_2713,N_1532,N_194);
or U2714 (N_2714,N_611,N_1911);
and U2715 (N_2715,N_1084,N_2368);
nand U2716 (N_2716,N_2442,N_1860);
nor U2717 (N_2717,N_1148,N_147);
or U2718 (N_2718,N_725,N_1402);
or U2719 (N_2719,N_1340,N_1563);
nand U2720 (N_2720,N_939,N_1952);
nand U2721 (N_2721,N_406,N_1862);
nand U2722 (N_2722,N_609,N_436);
nor U2723 (N_2723,N_921,N_1365);
nand U2724 (N_2724,N_1261,N_1258);
nor U2725 (N_2725,N_1189,N_1847);
and U2726 (N_2726,N_1357,N_11);
and U2727 (N_2727,N_260,N_1861);
nand U2728 (N_2728,N_241,N_2264);
or U2729 (N_2729,N_199,N_1735);
and U2730 (N_2730,N_2203,N_532);
nor U2731 (N_2731,N_723,N_517);
and U2732 (N_2732,N_706,N_398);
nor U2733 (N_2733,N_2210,N_513);
nand U2734 (N_2734,N_2155,N_720);
and U2735 (N_2735,N_376,N_1288);
nand U2736 (N_2736,N_2032,N_1263);
and U2737 (N_2737,N_2181,N_371);
xor U2738 (N_2738,N_2423,N_1510);
or U2739 (N_2739,N_1842,N_1147);
nor U2740 (N_2740,N_631,N_78);
nor U2741 (N_2741,N_1989,N_1134);
nand U2742 (N_2742,N_472,N_583);
and U2743 (N_2743,N_657,N_2341);
nor U2744 (N_2744,N_45,N_134);
and U2745 (N_2745,N_512,N_163);
nor U2746 (N_2746,N_2151,N_2195);
and U2747 (N_2747,N_1008,N_2045);
nor U2748 (N_2748,N_1023,N_1108);
and U2749 (N_2749,N_1727,N_2023);
xor U2750 (N_2750,N_1123,N_520);
nand U2751 (N_2751,N_1088,N_1825);
or U2752 (N_2752,N_1327,N_487);
or U2753 (N_2753,N_1162,N_839);
nor U2754 (N_2754,N_319,N_1581);
and U2755 (N_2755,N_419,N_224);
or U2756 (N_2756,N_1803,N_2306);
and U2757 (N_2757,N_895,N_2221);
nor U2758 (N_2758,N_601,N_1272);
and U2759 (N_2759,N_592,N_867);
or U2760 (N_2760,N_346,N_1895);
xnor U2761 (N_2761,N_1914,N_861);
and U2762 (N_2762,N_87,N_1641);
and U2763 (N_2763,N_680,N_2440);
xnor U2764 (N_2764,N_752,N_2404);
nor U2765 (N_2765,N_1782,N_1381);
and U2766 (N_2766,N_1330,N_1587);
or U2767 (N_2767,N_629,N_342);
or U2768 (N_2768,N_335,N_1579);
nand U2769 (N_2769,N_2296,N_2066);
or U2770 (N_2770,N_2164,N_182);
or U2771 (N_2771,N_1235,N_962);
or U2772 (N_2772,N_1129,N_1687);
and U2773 (N_2773,N_2140,N_2091);
xnor U2774 (N_2774,N_21,N_2124);
or U2775 (N_2775,N_2448,N_236);
nand U2776 (N_2776,N_128,N_418);
nor U2777 (N_2777,N_1672,N_1374);
and U2778 (N_2778,N_586,N_2036);
and U2779 (N_2779,N_1281,N_969);
and U2780 (N_2780,N_833,N_482);
nand U2781 (N_2781,N_2175,N_1138);
nand U2782 (N_2782,N_2393,N_430);
or U2783 (N_2783,N_524,N_1125);
xor U2784 (N_2784,N_2383,N_458);
or U2785 (N_2785,N_1784,N_273);
nor U2786 (N_2786,N_758,N_2460);
nand U2787 (N_2787,N_1933,N_2378);
nand U2788 (N_2788,N_1995,N_26);
xnor U2789 (N_2789,N_359,N_1160);
and U2790 (N_2790,N_484,N_1028);
nand U2791 (N_2791,N_727,N_980);
nor U2792 (N_2792,N_1467,N_327);
and U2793 (N_2793,N_894,N_1116);
nor U2794 (N_2794,N_457,N_348);
nand U2795 (N_2795,N_1133,N_2260);
or U2796 (N_2796,N_306,N_565);
nand U2797 (N_2797,N_12,N_1717);
xor U2798 (N_2798,N_452,N_251);
nand U2799 (N_2799,N_2417,N_807);
and U2800 (N_2800,N_661,N_445);
xnor U2801 (N_2801,N_989,N_549);
or U2802 (N_2802,N_2418,N_106);
or U2803 (N_2803,N_2314,N_349);
nand U2804 (N_2804,N_506,N_1572);
nor U2805 (N_2805,N_1500,N_2226);
and U2806 (N_2806,N_528,N_77);
nor U2807 (N_2807,N_2033,N_1900);
nor U2808 (N_2808,N_1344,N_2461);
nand U2809 (N_2809,N_1716,N_1640);
nand U2810 (N_2810,N_2402,N_96);
nand U2811 (N_2811,N_39,N_2107);
nand U2812 (N_2812,N_1869,N_1104);
or U2813 (N_2813,N_508,N_1267);
nor U2814 (N_2814,N_1436,N_1470);
or U2815 (N_2815,N_207,N_1226);
or U2816 (N_2816,N_2062,N_1815);
nand U2817 (N_2817,N_1433,N_1854);
and U2818 (N_2818,N_340,N_1561);
nor U2819 (N_2819,N_5,N_2246);
and U2820 (N_2820,N_1371,N_1788);
nor U2821 (N_2821,N_2236,N_33);
nand U2822 (N_2822,N_1445,N_228);
or U2823 (N_2823,N_2339,N_2025);
xnor U2824 (N_2824,N_1151,N_223);
nand U2825 (N_2825,N_1260,N_1499);
and U2826 (N_2826,N_1634,N_1554);
nor U2827 (N_2827,N_402,N_1607);
or U2828 (N_2828,N_614,N_446);
xor U2829 (N_2829,N_2240,N_1188);
and U2830 (N_2830,N_2327,N_1757);
nand U2831 (N_2831,N_318,N_1521);
and U2832 (N_2832,N_1027,N_28);
or U2833 (N_2833,N_1954,N_1452);
nand U2834 (N_2834,N_2026,N_238);
nor U2835 (N_2835,N_1193,N_1917);
nor U2836 (N_2836,N_1957,N_2425);
nor U2837 (N_2837,N_2084,N_410);
nor U2838 (N_2838,N_816,N_461);
nor U2839 (N_2839,N_534,N_943);
nand U2840 (N_2840,N_1367,N_2362);
and U2841 (N_2841,N_740,N_1620);
xor U2842 (N_2842,N_1022,N_107);
or U2843 (N_2843,N_424,N_1576);
or U2844 (N_2844,N_1710,N_1265);
or U2845 (N_2845,N_1002,N_2482);
and U2846 (N_2846,N_143,N_133);
nand U2847 (N_2847,N_1929,N_1137);
nor U2848 (N_2848,N_168,N_1840);
nor U2849 (N_2849,N_2165,N_529);
and U2850 (N_2850,N_779,N_1166);
or U2851 (N_2851,N_734,N_1819);
nand U2852 (N_2852,N_1586,N_801);
and U2853 (N_2853,N_1231,N_257);
or U2854 (N_2854,N_778,N_627);
nor U2855 (N_2855,N_1871,N_756);
or U2856 (N_2856,N_1017,N_863);
nor U2857 (N_2857,N_841,N_300);
xnor U2858 (N_2858,N_1878,N_139);
or U2859 (N_2859,N_638,N_413);
and U2860 (N_2860,N_1548,N_176);
nor U2861 (N_2861,N_864,N_1465);
or U2862 (N_2862,N_1809,N_1912);
or U2863 (N_2863,N_1829,N_15);
nor U2864 (N_2864,N_2358,N_333);
and U2865 (N_2865,N_1018,N_1669);
nand U2866 (N_2866,N_1802,N_997);
nor U2867 (N_2867,N_924,N_2072);
xor U2868 (N_2868,N_367,N_2283);
or U2869 (N_2869,N_844,N_509);
nand U2870 (N_2870,N_411,N_670);
and U2871 (N_2871,N_1783,N_1206);
and U2872 (N_2872,N_1443,N_1674);
nand U2873 (N_2873,N_1711,N_656);
nor U2874 (N_2874,N_2034,N_2357);
nor U2875 (N_2875,N_417,N_724);
and U2876 (N_2876,N_57,N_1714);
nand U2877 (N_2877,N_1345,N_931);
nor U2878 (N_2878,N_322,N_373);
nor U2879 (N_2879,N_17,N_1517);
nor U2880 (N_2880,N_186,N_1738);
and U2881 (N_2881,N_1250,N_64);
nand U2882 (N_2882,N_2087,N_1481);
nor U2883 (N_2883,N_885,N_2196);
or U2884 (N_2884,N_86,N_1550);
nand U2885 (N_2885,N_718,N_2487);
and U2886 (N_2886,N_1488,N_2311);
nor U2887 (N_2887,N_280,N_1988);
and U2888 (N_2888,N_2057,N_1844);
and U2889 (N_2889,N_1463,N_1000);
nor U2890 (N_2890,N_578,N_881);
and U2891 (N_2891,N_1742,N_2462);
and U2892 (N_2892,N_790,N_336);
nand U2893 (N_2893,N_714,N_1143);
nand U2894 (N_2894,N_933,N_2200);
xnor U2895 (N_2895,N_860,N_998);
nor U2896 (N_2896,N_2177,N_829);
nor U2897 (N_2897,N_954,N_317);
nand U2898 (N_2898,N_2239,N_1435);
xnor U2899 (N_2899,N_2077,N_1074);
xnor U2900 (N_2900,N_2258,N_1778);
or U2901 (N_2901,N_2410,N_1732);
nand U2902 (N_2902,N_2219,N_1349);
and U2903 (N_2903,N_1232,N_1959);
nor U2904 (N_2904,N_2204,N_952);
or U2905 (N_2905,N_798,N_1520);
nor U2906 (N_2906,N_1255,N_184);
nand U2907 (N_2907,N_544,N_2224);
nor U2908 (N_2908,N_1295,N_557);
nor U2909 (N_2909,N_1915,N_2248);
and U2910 (N_2910,N_2432,N_1174);
nor U2911 (N_2911,N_126,N_200);
nor U2912 (N_2912,N_1045,N_1076);
xor U2913 (N_2913,N_82,N_19);
nor U2914 (N_2914,N_1385,N_2459);
or U2915 (N_2915,N_884,N_1090);
nor U2916 (N_2916,N_1212,N_123);
xor U2917 (N_2917,N_465,N_1984);
or U2918 (N_2918,N_2108,N_982);
nand U2919 (N_2919,N_618,N_283);
or U2920 (N_2920,N_2391,N_1429);
xor U2921 (N_2921,N_1616,N_1225);
xnor U2922 (N_2922,N_185,N_2396);
xor U2923 (N_2923,N_2085,N_1042);
and U2924 (N_2924,N_1141,N_2012);
and U2925 (N_2925,N_1442,N_1705);
and U2926 (N_2926,N_2354,N_1302);
or U2927 (N_2927,N_1657,N_2268);
and U2928 (N_2928,N_1748,N_1173);
nand U2929 (N_2929,N_742,N_2300);
or U2930 (N_2930,N_1903,N_292);
nor U2931 (N_2931,N_2017,N_242);
xor U2932 (N_2932,N_79,N_751);
or U2933 (N_2933,N_662,N_1913);
nand U2934 (N_2934,N_2115,N_1109);
and U2935 (N_2935,N_281,N_1833);
or U2936 (N_2936,N_1533,N_523);
and U2937 (N_2937,N_1857,N_2384);
nand U2938 (N_2938,N_1752,N_2466);
nand U2939 (N_2939,N_1598,N_1721);
and U2940 (N_2940,N_2444,N_912);
nor U2941 (N_2941,N_157,N_1780);
xor U2942 (N_2942,N_191,N_217);
nor U2943 (N_2943,N_1668,N_621);
xor U2944 (N_2944,N_187,N_561);
and U2945 (N_2945,N_703,N_1677);
or U2946 (N_2946,N_1702,N_362);
nor U2947 (N_2947,N_500,N_930);
nand U2948 (N_2948,N_2261,N_350);
or U2949 (N_2949,N_1718,N_329);
or U2950 (N_2950,N_1230,N_1398);
and U2951 (N_2951,N_814,N_2456);
and U2952 (N_2952,N_1153,N_855);
and U2953 (N_2953,N_682,N_908);
or U2954 (N_2954,N_1165,N_763);
and U2955 (N_2955,N_761,N_950);
and U2956 (N_2956,N_808,N_854);
nand U2957 (N_2957,N_619,N_1629);
nor U2958 (N_2958,N_1642,N_666);
and U2959 (N_2959,N_1534,N_1200);
nor U2960 (N_2960,N_1645,N_1112);
or U2961 (N_2961,N_566,N_1313);
nand U2962 (N_2962,N_976,N_539);
xor U2963 (N_2963,N_1069,N_266);
and U2964 (N_2964,N_882,N_2127);
nand U2965 (N_2965,N_2486,N_1683);
and U2966 (N_2966,N_1252,N_1848);
nor U2967 (N_2967,N_2211,N_1817);
or U2968 (N_2968,N_574,N_244);
nand U2969 (N_2969,N_61,N_1694);
nor U2970 (N_2970,N_1476,N_2430);
nand U2971 (N_2971,N_301,N_1972);
or U2972 (N_2972,N_481,N_2355);
nand U2973 (N_2973,N_1766,N_1685);
nand U2974 (N_2974,N_360,N_1758);
and U2975 (N_2975,N_42,N_772);
nor U2976 (N_2976,N_2379,N_1971);
and U2977 (N_2977,N_2147,N_122);
nand U2978 (N_2978,N_2007,N_678);
nor U2979 (N_2979,N_956,N_212);
and U2980 (N_2980,N_1172,N_314);
xor U2981 (N_2981,N_2090,N_569);
nand U2982 (N_2982,N_935,N_1583);
nand U2983 (N_2983,N_766,N_1320);
nand U2984 (N_2984,N_2292,N_1889);
and U2985 (N_2985,N_316,N_1613);
nor U2986 (N_2986,N_285,N_594);
nor U2987 (N_2987,N_996,N_1264);
or U2988 (N_2988,N_2303,N_1518);
xnor U2989 (N_2989,N_959,N_485);
nand U2990 (N_2990,N_377,N_1726);
nor U2991 (N_2991,N_1556,N_843);
nor U2992 (N_2992,N_890,N_542);
nand U2993 (N_2993,N_1075,N_365);
nor U2994 (N_2994,N_2295,N_2317);
and U2995 (N_2995,N_2001,N_2234);
and U2996 (N_2996,N_1649,N_979);
or U2997 (N_2997,N_270,N_1787);
nor U2998 (N_2998,N_1980,N_1759);
xor U2999 (N_2999,N_250,N_382);
nand U3000 (N_3000,N_2348,N_2297);
or U3001 (N_3001,N_2039,N_2102);
and U3002 (N_3002,N_2492,N_167);
or U3003 (N_3003,N_1700,N_1460);
nand U3004 (N_3004,N_1291,N_920);
xor U3005 (N_3005,N_828,N_1894);
or U3006 (N_3006,N_2468,N_1209);
nor U3007 (N_3007,N_1464,N_852);
nor U3008 (N_3008,N_760,N_2245);
nor U3009 (N_3009,N_2347,N_2008);
nor U3010 (N_3010,N_909,N_53);
nand U3011 (N_3011,N_1526,N_560);
and U3012 (N_3012,N_1105,N_2290);
or U3013 (N_3013,N_395,N_1704);
nand U3014 (N_3014,N_1991,N_202);
nor U3015 (N_3015,N_1632,N_2215);
and U3016 (N_3016,N_1126,N_219);
xor U3017 (N_3017,N_2309,N_579);
nor U3018 (N_3018,N_1183,N_252);
xnor U3019 (N_3019,N_345,N_1205);
nor U3020 (N_3020,N_278,N_1728);
nor U3021 (N_3021,N_2126,N_289);
nand U3022 (N_3022,N_840,N_2336);
or U3023 (N_3023,N_2166,N_1567);
nand U3024 (N_3024,N_1603,N_699);
and U3025 (N_3025,N_1159,N_1171);
or U3026 (N_3026,N_2399,N_388);
nor U3027 (N_3027,N_230,N_1953);
and U3028 (N_3028,N_2143,N_9);
or U3029 (N_3029,N_255,N_1336);
nor U3030 (N_3030,N_2159,N_635);
and U3031 (N_3031,N_425,N_438);
nand U3032 (N_3032,N_1893,N_325);
and U3033 (N_3033,N_2067,N_0);
or U3034 (N_3034,N_135,N_2132);
and U3035 (N_3035,N_2135,N_1190);
or U3036 (N_3036,N_1947,N_2367);
or U3037 (N_3037,N_2325,N_489);
and U3038 (N_3038,N_94,N_713);
and U3039 (N_3039,N_385,N_1999);
nand U3040 (N_3040,N_1136,N_326);
nor U3041 (N_3041,N_294,N_915);
nor U3042 (N_3042,N_1324,N_2095);
nor U3043 (N_3043,N_1421,N_2060);
or U3044 (N_3044,N_2097,N_462);
or U3045 (N_3045,N_737,N_2435);
and U3046 (N_3046,N_1038,N_2326);
nor U3047 (N_3047,N_415,N_46);
nand U3048 (N_3048,N_1358,N_974);
or U3049 (N_3049,N_22,N_2385);
and U3050 (N_3050,N_1754,N_499);
nor U3051 (N_3051,N_2049,N_2332);
or U3052 (N_3052,N_1211,N_1360);
nor U3053 (N_3053,N_412,N_1831);
or U3054 (N_3054,N_1555,N_2279);
nor U3055 (N_3055,N_1931,N_826);
nand U3056 (N_3056,N_1712,N_1106);
and U3057 (N_3057,N_2420,N_851);
nand U3058 (N_3058,N_83,N_1347);
or U3059 (N_3059,N_1354,N_2024);
and U3060 (N_3060,N_762,N_2394);
xor U3061 (N_3061,N_288,N_690);
xor U3062 (N_3062,N_1410,N_1622);
and U3063 (N_3063,N_1420,N_1300);
and U3064 (N_3064,N_31,N_2052);
nor U3065 (N_3065,N_2267,N_927);
and U3066 (N_3066,N_2162,N_2047);
or U3067 (N_3067,N_1359,N_2037);
and U3068 (N_3068,N_1731,N_2167);
nor U3069 (N_3069,N_922,N_1152);
and U3070 (N_3070,N_1664,N_2436);
nor U3071 (N_3071,N_1304,N_2170);
and U3072 (N_3072,N_810,N_2481);
nor U3073 (N_3073,N_262,N_2238);
or U3074 (N_3074,N_2454,N_1095);
and U3075 (N_3075,N_722,N_1425);
or U3076 (N_3076,N_1573,N_2081);
or U3077 (N_3077,N_1099,N_1689);
nor U3078 (N_3078,N_494,N_1262);
nor U3079 (N_3079,N_68,N_177);
and U3080 (N_3080,N_1600,N_404);
or U3081 (N_3081,N_590,N_1631);
and U3082 (N_3082,N_2443,N_1590);
and U3083 (N_3083,N_2152,N_120);
nand U3084 (N_3084,N_1305,N_1195);
nor U3085 (N_3085,N_764,N_1818);
and U3086 (N_3086,N_1808,N_942);
nor U3087 (N_3087,N_1897,N_1187);
nand U3088 (N_3088,N_1471,N_1944);
xnor U3089 (N_3089,N_29,N_2437);
and U3090 (N_3090,N_1987,N_492);
or U3091 (N_3091,N_1557,N_1036);
and U3092 (N_3092,N_1679,N_1795);
nand U3093 (N_3093,N_209,N_142);
xor U3094 (N_3094,N_2284,N_1278);
nor U3095 (N_3095,N_269,N_2104);
nor U3096 (N_3096,N_2453,N_1628);
or U3097 (N_3097,N_770,N_624);
nor U3098 (N_3098,N_7,N_2315);
nand U3099 (N_3099,N_1156,N_1118);
and U3100 (N_3100,N_2262,N_1707);
nand U3101 (N_3101,N_1453,N_1127);
or U3102 (N_3102,N_1297,N_1455);
and U3103 (N_3103,N_1538,N_1713);
nor U3104 (N_3104,N_1081,N_985);
or U3105 (N_3105,N_966,N_1965);
and U3106 (N_3106,N_1100,N_1394);
or U3107 (N_3107,N_401,N_1060);
nor U3108 (N_3108,N_1941,N_531);
xnor U3109 (N_3109,N_100,N_1419);
and U3110 (N_3110,N_13,N_1892);
and U3111 (N_3111,N_702,N_898);
or U3112 (N_3112,N_1880,N_1885);
nor U3113 (N_3113,N_391,N_1981);
xnor U3114 (N_3114,N_623,N_1703);
and U3115 (N_3115,N_204,N_2192);
and U3116 (N_3116,N_27,N_6);
nor U3117 (N_3117,N_2015,N_47);
or U3118 (N_3118,N_1466,N_889);
and U3119 (N_3119,N_2364,N_2028);
nor U3120 (N_3120,N_1207,N_1751);
nor U3121 (N_3121,N_1937,N_677);
or U3122 (N_3122,N_2089,N_1722);
nand U3123 (N_3123,N_1266,N_393);
nor U3124 (N_3124,N_2241,N_2030);
nand U3125 (N_3125,N_2005,N_1875);
xnor U3126 (N_3126,N_502,N_1821);
or U3127 (N_3127,N_1178,N_838);
or U3128 (N_3128,N_2137,N_667);
xor U3129 (N_3129,N_409,N_2099);
nor U3130 (N_3130,N_1768,N_796);
xnor U3131 (N_3131,N_1507,N_1169);
nand U3132 (N_3132,N_2020,N_1873);
or U3133 (N_3133,N_331,N_1301);
nand U3134 (N_3134,N_1610,N_405);
or U3135 (N_3135,N_911,N_705);
nor U3136 (N_3136,N_2042,N_220);
or U3137 (N_3137,N_846,N_2031);
or U3138 (N_3138,N_696,N_917);
nand U3139 (N_3139,N_40,N_2463);
or U3140 (N_3140,N_1967,N_664);
nor U3141 (N_3141,N_1368,N_1102);
xor U3142 (N_3142,N_2044,N_1124);
or U3143 (N_3143,N_822,N_441);
nand U3144 (N_3144,N_604,N_1720);
xor U3145 (N_3145,N_820,N_2313);
nor U3146 (N_3146,N_497,N_1196);
nand U3147 (N_3147,N_334,N_1275);
or U3148 (N_3148,N_1477,N_2154);
and U3149 (N_3149,N_550,N_399);
and U3150 (N_3150,N_916,N_999);
xnor U3151 (N_3151,N_2086,N_2490);
and U3152 (N_3152,N_645,N_1216);
and U3153 (N_3153,N_2009,N_243);
and U3154 (N_3154,N_1186,N_1279);
and U3155 (N_3155,N_261,N_85);
nand U3156 (N_3156,N_471,N_1497);
nor U3157 (N_3157,N_2235,N_907);
and U3158 (N_3158,N_1777,N_963);
xor U3159 (N_3159,N_1268,N_1939);
nand U3160 (N_3160,N_2206,N_2479);
or U3161 (N_3161,N_192,N_2496);
and U3162 (N_3162,N_18,N_1448);
nand U3163 (N_3163,N_572,N_1569);
nor U3164 (N_3164,N_1637,N_1229);
and U3165 (N_3165,N_1745,N_1380);
or U3166 (N_3166,N_1814,N_681);
and U3167 (N_3167,N_153,N_447);
and U3168 (N_3168,N_1943,N_994);
nor U3169 (N_3169,N_1888,N_1234);
and U3170 (N_3170,N_510,N_1982);
or U3171 (N_3171,N_2457,N_1661);
xor U3172 (N_3172,N_433,N_2478);
or U3173 (N_3173,N_856,N_455);
nor U3174 (N_3174,N_468,N_414);
or U3175 (N_3175,N_92,N_2471);
and U3176 (N_3176,N_464,N_2051);
xnor U3177 (N_3177,N_1370,N_659);
xor U3178 (N_3178,N_1085,N_1870);
or U3179 (N_3179,N_1019,N_679);
nand U3180 (N_3180,N_154,N_947);
and U3181 (N_3181,N_582,N_179);
or U3182 (N_3182,N_2429,N_1562);
nor U3183 (N_3183,N_800,N_2389);
and U3184 (N_3184,N_1695,N_1872);
nor U3185 (N_3185,N_600,N_303);
nand U3186 (N_3186,N_2227,N_1693);
and U3187 (N_3187,N_1372,N_55);
xor U3188 (N_3188,N_1338,N_1308);
nor U3189 (N_3189,N_221,N_2103);
or U3190 (N_3190,N_2287,N_1653);
nor U3191 (N_3191,N_1219,N_265);
nor U3192 (N_3192,N_973,N_84);
or U3193 (N_3193,N_2449,N_1624);
nand U3194 (N_3194,N_171,N_1366);
nor U3195 (N_3195,N_2048,N_2186);
or U3196 (N_3196,N_971,N_478);
and U3197 (N_3197,N_338,N_1031);
or U3198 (N_3198,N_1458,N_1050);
or U3199 (N_3199,N_2121,N_1375);
nor U3200 (N_3200,N_597,N_1461);
nand U3201 (N_3201,N_558,N_617);
or U3202 (N_3202,N_1456,N_983);
or U3203 (N_3203,N_847,N_2286);
or U3204 (N_3204,N_233,N_1222);
nor U3205 (N_3205,N_2128,N_665);
nor U3206 (N_3206,N_1393,N_1837);
nand U3207 (N_3207,N_1257,N_977);
and U3208 (N_3208,N_339,N_946);
or U3209 (N_3209,N_2422,N_893);
nand U3210 (N_3210,N_1654,N_2353);
nor U3211 (N_3211,N_873,N_960);
or U3212 (N_3212,N_1811,N_1901);
nor U3213 (N_3213,N_2266,N_1568);
nand U3214 (N_3214,N_2272,N_1098);
or U3215 (N_3215,N_626,N_926);
xnor U3216 (N_3216,N_310,N_548);
and U3217 (N_3217,N_1149,N_1348);
xnor U3218 (N_3218,N_2488,N_1767);
nand U3219 (N_3219,N_637,N_1606);
and U3220 (N_3220,N_1322,N_470);
nor U3221 (N_3221,N_576,N_493);
nand U3222 (N_3222,N_1335,N_1867);
nor U3223 (N_3223,N_1523,N_439);
xnor U3224 (N_3224,N_1376,N_1908);
nand U3225 (N_3225,N_2289,N_607);
and U3226 (N_3226,N_258,N_2058);
nor U3227 (N_3227,N_1487,N_1101);
nor U3228 (N_3228,N_673,N_253);
and U3229 (N_3229,N_2100,N_1623);
or U3230 (N_3230,N_1948,N_1170);
or U3231 (N_3231,N_1850,N_2125);
nor U3232 (N_3232,N_1985,N_902);
xor U3233 (N_3233,N_2343,N_1034);
or U3234 (N_3234,N_2141,N_1364);
nand U3235 (N_3235,N_2321,N_246);
nand U3236 (N_3236,N_2499,N_1650);
xnor U3237 (N_3237,N_1495,N_229);
nand U3238 (N_3238,N_2217,N_781);
and U3239 (N_3239,N_1029,N_1427);
nor U3240 (N_3240,N_434,N_1923);
or U3241 (N_3241,N_1696,N_1827);
nor U3242 (N_3242,N_817,N_2387);
and U3243 (N_3243,N_1916,N_1388);
nand U3244 (N_3244,N_1770,N_1208);
nand U3245 (N_3245,N_297,N_818);
and U3246 (N_3246,N_1092,N_1293);
or U3247 (N_3247,N_953,N_305);
or U3248 (N_3248,N_2438,N_2450);
nand U3249 (N_3249,N_1412,N_1404);
or U3250 (N_3250,N_308,N_1062);
or U3251 (N_3251,N_80,N_773);
or U3252 (N_3252,N_151,N_1009);
nand U3253 (N_3253,N_1975,N_2027);
nand U3254 (N_3254,N_1373,N_2380);
nand U3255 (N_3255,N_1882,N_1969);
and U3256 (N_3256,N_1423,N_1647);
nor U3257 (N_3257,N_1530,N_2011);
or U3258 (N_3258,N_2269,N_1294);
and U3259 (N_3259,N_1181,N_991);
and U3260 (N_3260,N_1769,N_589);
or U3261 (N_3261,N_2073,N_2363);
or U3262 (N_3262,N_89,N_2346);
and U3263 (N_3263,N_4,N_1334);
nor U3264 (N_3264,N_2352,N_1547);
and U3265 (N_3265,N_1935,N_1054);
and U3266 (N_3266,N_2249,N_1922);
and U3267 (N_3267,N_2063,N_2183);
or U3268 (N_3268,N_1608,N_2199);
or U3269 (N_3269,N_1363,N_2421);
or U3270 (N_3270,N_671,N_1775);
nand U3271 (N_3271,N_361,N_2202);
nor U3272 (N_3272,N_2483,N_71);
and U3273 (N_3273,N_1089,N_2094);
nand U3274 (N_3274,N_1723,N_1601);
nand U3275 (N_3275,N_830,N_919);
or U3276 (N_3276,N_1454,N_710);
nand U3277 (N_3277,N_1314,N_1280);
and U3278 (N_3278,N_1719,N_479);
nor U3279 (N_3279,N_1341,N_1384);
nor U3280 (N_3280,N_2342,N_75);
nor U3281 (N_3281,N_2307,N_1781);
nor U3282 (N_3282,N_1549,N_320);
or U3283 (N_3283,N_1515,N_745);
and U3284 (N_3284,N_2497,N_136);
or U3285 (N_3285,N_2434,N_1449);
nor U3286 (N_3286,N_2055,N_1886);
and U3287 (N_3287,N_141,N_1799);
nand U3288 (N_3288,N_1541,N_1813);
or U3289 (N_3289,N_1830,N_1043);
or U3290 (N_3290,N_1403,N_2285);
and U3291 (N_3291,N_774,N_587);
or U3292 (N_3292,N_2244,N_2318);
nor U3293 (N_3293,N_1771,N_538);
nor U3294 (N_3294,N_287,N_2013);
nand U3295 (N_3295,N_988,N_2304);
nand U3296 (N_3296,N_568,N_719);
nand U3297 (N_3297,N_1773,N_1001);
or U3298 (N_3298,N_1175,N_834);
and U3299 (N_3299,N_613,N_1945);
xor U3300 (N_3300,N_1012,N_2412);
nor U3301 (N_3301,N_337,N_1438);
nand U3302 (N_3302,N_1619,N_835);
nand U3303 (N_3303,N_110,N_1287);
or U3304 (N_3304,N_535,N_2390);
or U3305 (N_3305,N_2138,N_1450);
nand U3306 (N_3306,N_1306,N_1409);
nand U3307 (N_3307,N_2157,N_1110);
or U3308 (N_3308,N_1224,N_694);
nor U3309 (N_3309,N_1516,N_1874);
and U3310 (N_3310,N_581,N_2257);
nor U3311 (N_3311,N_1079,N_880);
nor U3312 (N_3312,N_2220,N_311);
or U3313 (N_3313,N_984,N_1514);
nand U3314 (N_3314,N_435,N_2150);
nor U3315 (N_3315,N_130,N_1503);
nand U3316 (N_3316,N_2109,N_769);
and U3317 (N_3317,N_2403,N_651);
or U3318 (N_3318,N_1822,N_1627);
and U3319 (N_3319,N_1729,N_1715);
and U3320 (N_3320,N_2189,N_2163);
or U3321 (N_3321,N_245,N_738);
nand U3322 (N_3322,N_1240,N_1626);
nand U3323 (N_3323,N_978,N_296);
or U3324 (N_3324,N_1644,N_188);
or U3325 (N_3325,N_1333,N_423);
nand U3326 (N_3326,N_1835,N_380);
and U3327 (N_3327,N_1785,N_685);
or U3328 (N_3328,N_1071,N_1277);
or U3329 (N_3329,N_299,N_2270);
and U3330 (N_3330,N_48,N_1228);
or U3331 (N_3331,N_2254,N_488);
or U3332 (N_3332,N_577,N_1992);
or U3333 (N_3333,N_1096,N_1318);
and U3334 (N_3334,N_2255,N_164);
nand U3335 (N_3335,N_1578,N_688);
xor U3336 (N_3336,N_540,N_955);
xnor U3337 (N_3337,N_467,N_1746);
nand U3338 (N_3338,N_2397,N_1362);
and U3339 (N_3339,N_1391,N_1638);
nand U3340 (N_3340,N_2495,N_483);
or U3341 (N_3341,N_1519,N_396);
or U3342 (N_3342,N_1407,N_551);
xnor U3343 (N_3343,N_1502,N_2316);
nor U3344 (N_3344,N_137,N_1682);
or U3345 (N_3345,N_473,N_341);
nand U3346 (N_3346,N_2451,N_1977);
nor U3347 (N_3347,N_2388,N_1676);
nor U3348 (N_3348,N_1698,N_2184);
or U3349 (N_3349,N_2208,N_1810);
nor U3350 (N_3350,N_968,N_1284);
or U3351 (N_3351,N_1332,N_1236);
nand U3352 (N_3352,N_1571,N_2171);
nand U3353 (N_3353,N_20,N_390);
xnor U3354 (N_3354,N_1061,N_1643);
xnor U3355 (N_3355,N_1039,N_899);
xor U3356 (N_3356,N_1080,N_602);
nor U3357 (N_3357,N_2065,N_1564);
or U3358 (N_3358,N_1457,N_2426);
nand U3359 (N_3359,N_183,N_2198);
nand U3360 (N_3360,N_654,N_1927);
nor U3361 (N_3361,N_559,N_2004);
nor U3362 (N_3362,N_347,N_2281);
and U3363 (N_3363,N_2427,N_1424);
nand U3364 (N_3364,N_1087,N_870);
nand U3365 (N_3365,N_1553,N_172);
or U3366 (N_3366,N_1741,N_663);
nand U3367 (N_3367,N_91,N_1066);
or U3368 (N_3368,N_878,N_1239);
or U3369 (N_3369,N_307,N_97);
nor U3370 (N_3370,N_731,N_585);
nor U3371 (N_3371,N_695,N_2130);
and U3372 (N_3372,N_1736,N_1907);
or U3373 (N_3373,N_448,N_1217);
or U3374 (N_3374,N_573,N_1996);
or U3375 (N_3375,N_1298,N_936);
or U3376 (N_3376,N_2351,N_277);
and U3377 (N_3377,N_612,N_2401);
and U3378 (N_3378,N_1609,N_456);
and U3379 (N_3379,N_1253,N_2146);
nand U3380 (N_3380,N_647,N_195);
and U3381 (N_3381,N_748,N_2040);
nor U3382 (N_3382,N_1792,N_24);
nor U3383 (N_3383,N_203,N_2230);
nand U3384 (N_3384,N_1249,N_932);
and U3385 (N_3385,N_1329,N_271);
nand U3386 (N_3386,N_837,N_1529);
nand U3387 (N_3387,N_2377,N_1446);
nand U3388 (N_3388,N_1528,N_115);
and U3389 (N_3389,N_2445,N_109);
nand U3390 (N_3390,N_1411,N_2019);
nand U3391 (N_3391,N_282,N_1706);
xor U3392 (N_3392,N_2216,N_254);
and U3393 (N_3393,N_545,N_1879);
xnor U3394 (N_3394,N_170,N_328);
or U3395 (N_3395,N_2333,N_1254);
or U3396 (N_3396,N_625,N_780);
and U3397 (N_3397,N_2114,N_521);
nor U3398 (N_3398,N_2161,N_687);
nor U3399 (N_3399,N_1292,N_1934);
and U3400 (N_3400,N_1760,N_1979);
and U3401 (N_3401,N_1078,N_131);
or U3402 (N_3402,N_970,N_1724);
or U3403 (N_3403,N_76,N_408);
or U3404 (N_3404,N_1750,N_2133);
nand U3405 (N_3405,N_1176,N_1599);
nand U3406 (N_3406,N_541,N_1490);
xnor U3407 (N_3407,N_2360,N_138);
and U3408 (N_3408,N_2328,N_1633);
nor U3409 (N_3409,N_1180,N_208);
nor U3410 (N_3410,N_2046,N_387);
nor U3411 (N_3411,N_934,N_1493);
nand U3412 (N_3412,N_150,N_286);
or U3413 (N_3413,N_900,N_2282);
nor U3414 (N_3414,N_2223,N_1237);
and U3415 (N_3415,N_1618,N_1772);
and U3416 (N_3416,N_1790,N_2322);
xnor U3417 (N_3417,N_2029,N_1524);
nand U3418 (N_3418,N_1164,N_1699);
nand U3419 (N_3419,N_2406,N_1779);
nand U3420 (N_3420,N_2370,N_1582);
and U3421 (N_3421,N_1475,N_2446);
or U3422 (N_3422,N_1346,N_466);
nor U3423 (N_3423,N_2131,N_990);
or U3424 (N_3424,N_1966,N_1115);
or U3425 (N_3425,N_2110,N_1636);
nor U3426 (N_3426,N_369,N_1049);
nand U3427 (N_3427,N_1968,N_1942);
or U3428 (N_3428,N_1511,N_2000);
nor U3429 (N_3429,N_2018,N_2075);
nor U3430 (N_3430,N_2467,N_1841);
nand U3431 (N_3431,N_697,N_2265);
nand U3432 (N_3432,N_2359,N_1697);
or U3433 (N_3433,N_268,N_1285);
nand U3434 (N_3434,N_2242,N_2116);
or U3435 (N_3435,N_103,N_897);
nor U3436 (N_3436,N_791,N_180);
or U3437 (N_3437,N_1290,N_813);
nor U3438 (N_3438,N_213,N_1413);
xor U3439 (N_3439,N_1011,N_1142);
and U3440 (N_3440,N_1494,N_370);
xor U3441 (N_3441,N_198,N_2071);
and U3442 (N_3442,N_2173,N_2484);
nand U3443 (N_3443,N_1978,N_1513);
nand U3444 (N_3444,N_793,N_1161);
and U3445 (N_3445,N_263,N_352);
xor U3446 (N_3446,N_2068,N_717);
nand U3447 (N_3447,N_74,N_1566);
nand U3448 (N_3448,N_1584,N_1472);
and U3449 (N_3449,N_1053,N_2373);
nand U3450 (N_3450,N_1743,N_653);
nand U3451 (N_3451,N_1820,N_1194);
nand U3452 (N_3452,N_1918,N_2356);
nor U3453 (N_3453,N_1612,N_1248);
nor U3454 (N_3454,N_1003,N_1282);
and U3455 (N_3455,N_2169,N_2129);
nand U3456 (N_3456,N_1326,N_2480);
and U3457 (N_3457,N_858,N_302);
and U3458 (N_3458,N_944,N_929);
nand U3459 (N_3459,N_925,N_700);
nor U3460 (N_3460,N_2277,N_2491);
nor U3461 (N_3461,N_41,N_239);
and U3462 (N_3462,N_610,N_469);
nor U3463 (N_3463,N_511,N_975);
nor U3464 (N_3464,N_189,N_35);
xnor U3465 (N_3465,N_2168,N_1065);
nand U3466 (N_3466,N_729,N_2228);
and U3467 (N_3467,N_1395,N_211);
nand U3468 (N_3468,N_1213,N_1753);
and U3469 (N_3469,N_1296,N_32);
nor U3470 (N_3470,N_675,N_1158);
and U3471 (N_3471,N_1220,N_1824);
and U3472 (N_3472,N_1199,N_730);
or U3473 (N_3473,N_1201,N_536);
nand U3474 (N_3474,N_1047,N_938);
and U3475 (N_3475,N_1242,N_649);
or U3476 (N_3476,N_2464,N_2092);
nor U3477 (N_3477,N_2455,N_1733);
or U3478 (N_3478,N_739,N_744);
nor U3479 (N_3479,N_503,N_1233);
and U3480 (N_3480,N_1405,N_8);
and U3481 (N_3481,N_38,N_1073);
nor U3482 (N_3482,N_905,N_1611);
nor U3483 (N_3483,N_620,N_36);
nor U3484 (N_3484,N_1055,N_476);
or U3485 (N_3485,N_2458,N_312);
and U3486 (N_3486,N_1145,N_437);
or U3487 (N_3487,N_1973,N_403);
nor U3488 (N_3488,N_1437,N_119);
nand U3489 (N_3489,N_1708,N_555);
nand U3490 (N_3490,N_1469,N_323);
or U3491 (N_3491,N_948,N_2088);
nand U3492 (N_3492,N_1325,N_1658);
nor U3493 (N_3493,N_442,N_2185);
or U3494 (N_3494,N_1005,N_2233);
or U3495 (N_3495,N_655,N_1067);
nand U3496 (N_3496,N_1964,N_945);
and U3497 (N_3497,N_264,N_1630);
nand U3498 (N_3498,N_505,N_1574);
nor U3499 (N_3499,N_2002,N_712);
nand U3500 (N_3500,N_1444,N_940);
or U3501 (N_3501,N_1891,N_1399);
nand U3502 (N_3502,N_2207,N_2187);
and U3503 (N_3503,N_803,N_811);
nand U3504 (N_3504,N_1351,N_1316);
or U3505 (N_3505,N_1361,N_1910);
nor U3506 (N_3506,N_1422,N_1227);
nand U3507 (N_3507,N_1310,N_272);
nand U3508 (N_3508,N_99,N_526);
and U3509 (N_3509,N_1283,N_684);
nor U3510 (N_3510,N_1839,N_1993);
nor U3511 (N_3511,N_1744,N_2179);
or U3512 (N_3512,N_1163,N_1331);
or U3513 (N_3513,N_43,N_1479);
or U3514 (N_3514,N_1414,N_2218);
and U3515 (N_3515,N_672,N_599);
and U3516 (N_3516,N_1828,N_903);
nand U3517 (N_3517,N_1868,N_173);
or U3518 (N_3518,N_819,N_1480);
nand U3519 (N_3519,N_2431,N_2337);
nand U3520 (N_3520,N_888,N_165);
nor U3521 (N_3521,N_1286,N_1765);
nor U3522 (N_3522,N_1120,N_2101);
nor U3523 (N_3523,N_190,N_1826);
or U3524 (N_3524,N_2142,N_630);
and U3525 (N_3525,N_1025,N_1016);
and U3526 (N_3526,N_477,N_850);
nor U3527 (N_3527,N_650,N_1851);
nor U3528 (N_3528,N_2275,N_1940);
or U3529 (N_3529,N_451,N_1315);
nand U3530 (N_3530,N_1648,N_708);
or U3531 (N_3531,N_144,N_1203);
and U3532 (N_3532,N_2376,N_480);
nand U3533 (N_3533,N_2056,N_2120);
and U3534 (N_3534,N_783,N_1139);
and U3535 (N_3535,N_1010,N_1652);
and U3536 (N_3536,N_877,N_1426);
and U3537 (N_3537,N_711,N_642);
and U3538 (N_3538,N_2180,N_859);
nor U3539 (N_3539,N_356,N_1072);
or U3540 (N_3540,N_432,N_235);
or U3541 (N_3541,N_995,N_584);
nor U3542 (N_3542,N_2350,N_768);
and U3543 (N_3543,N_2319,N_553);
nand U3544 (N_3544,N_1303,N_449);
xnor U3545 (N_3545,N_2428,N_1474);
or U3546 (N_3546,N_527,N_1675);
nand U3547 (N_3547,N_1864,N_460);
nor U3548 (N_3548,N_1185,N_1855);
and U3549 (N_3549,N_759,N_486);
or U3550 (N_3550,N_1339,N_2093);
xor U3551 (N_3551,N_1655,N_2148);
nand U3552 (N_3552,N_428,N_636);
nor U3553 (N_3553,N_2472,N_1776);
nand U3554 (N_3554,N_2178,N_169);
nor U3555 (N_3555,N_1621,N_1816);
nor U3556 (N_3556,N_1044,N_2160);
or U3557 (N_3557,N_1396,N_249);
or U3558 (N_3558,N_2106,N_1605);
xnor U3559 (N_3559,N_1543,N_556);
or U3560 (N_3560,N_530,N_2273);
nand U3561 (N_3561,N_1946,N_1896);
nand U3562 (N_3562,N_845,N_2470);
nor U3563 (N_3563,N_519,N_1041);
and U3564 (N_3564,N_1015,N_1177);
nand U3565 (N_3565,N_1244,N_1441);
or U3566 (N_3566,N_1859,N_1593);
or U3567 (N_3567,N_1030,N_2407);
or U3568 (N_3568,N_2366,N_683);
nand U3569 (N_3569,N_753,N_63);
or U3570 (N_3570,N_420,N_1192);
and U3571 (N_3571,N_1406,N_1747);
and U3572 (N_3572,N_1026,N_2294);
nor U3573 (N_3573,N_88,N_1210);
nand U3574 (N_3574,N_1114,N_1389);
and U3575 (N_3575,N_1970,N_2375);
or U3576 (N_3576,N_161,N_149);
xor U3577 (N_3577,N_1506,N_383);
or U3578 (N_3578,N_2003,N_1299);
or U3579 (N_3579,N_1307,N_2256);
and U3580 (N_3580,N_259,N_444);
xnor U3581 (N_3581,N_879,N_1887);
nand U3582 (N_3582,N_2229,N_2280);
and U3583 (N_3583,N_1447,N_1504);
xnor U3584 (N_3584,N_1673,N_1865);
nor U3585 (N_3585,N_227,N_214);
or U3586 (N_3586,N_1938,N_1462);
xnor U3587 (N_3587,N_1215,N_1680);
and U3588 (N_3588,N_883,N_1068);
or U3589 (N_3589,N_37,N_709);
nand U3590 (N_3590,N_1214,N_1604);
nand U3591 (N_3591,N_2079,N_1270);
or U3592 (N_3592,N_1246,N_815);
or U3593 (N_3593,N_750,N_1725);
and U3594 (N_3594,N_2237,N_379);
nand U3595 (N_3595,N_775,N_156);
or U3596 (N_3596,N_66,N_2447);
and U3597 (N_3597,N_2144,N_784);
nor U3598 (N_3598,N_747,N_2078);
nor U3599 (N_3599,N_1558,N_2082);
or U3600 (N_3600,N_2021,N_1167);
and U3601 (N_3601,N_2136,N_321);
and U3602 (N_3602,N_812,N_726);
nand U3603 (N_3603,N_1451,N_1256);
or U3604 (N_3604,N_564,N_1007);
or U3605 (N_3605,N_1135,N_152);
nor U3606 (N_3606,N_728,N_108);
xor U3607 (N_3607,N_293,N_2117);
xor U3608 (N_3608,N_363,N_1801);
nor U3609 (N_3609,N_580,N_496);
nand U3610 (N_3610,N_160,N_2320);
and U3611 (N_3611,N_440,N_782);
nand U3612 (N_3612,N_1024,N_1020);
nand U3613 (N_3613,N_1154,N_809);
or U3614 (N_3614,N_603,N_749);
or U3615 (N_3615,N_1037,N_234);
nand U3616 (N_3616,N_876,N_1786);
nor U3617 (N_3617,N_159,N_1317);
nor U3618 (N_3618,N_1883,N_1806);
and U3619 (N_3619,N_102,N_1103);
or U3620 (N_3620,N_1132,N_849);
and U3621 (N_3621,N_622,N_2298);
xnor U3622 (N_3622,N_735,N_60);
nor U3623 (N_3623,N_1595,N_1749);
nand U3624 (N_3624,N_2172,N_615);
or U3625 (N_3625,N_1051,N_1107);
nand U3626 (N_3626,N_1191,N_1004);
and U3627 (N_3627,N_1434,N_2414);
xnor U3628 (N_3628,N_475,N_1961);
nand U3629 (N_3629,N_923,N_1594);
nand U3630 (N_3630,N_49,N_2153);
nor U3631 (N_3631,N_162,N_887);
or U3632 (N_3632,N_498,N_2369);
xnor U3633 (N_3633,N_2469,N_1483);
nand U3634 (N_3634,N_788,N_591);
or U3635 (N_3635,N_1155,N_1570);
nor U3636 (N_3636,N_964,N_98);
nor U3637 (N_3637,N_596,N_30);
nand U3638 (N_3638,N_1094,N_1737);
or U3639 (N_3639,N_386,N_993);
or U3640 (N_3640,N_693,N_1508);
nand U3641 (N_3641,N_114,N_201);
nor U3642 (N_3642,N_1670,N_648);
nor U3643 (N_3643,N_2494,N_10);
and U3644 (N_3644,N_1798,N_1667);
nor U3645 (N_3645,N_1,N_1468);
xnor U3646 (N_3646,N_158,N_368);
nor U3647 (N_3647,N_1052,N_353);
and U3648 (N_3648,N_364,N_1184);
nor U3649 (N_3649,N_1221,N_1709);
and U3650 (N_3650,N_891,N_1289);
or U3651 (N_3651,N_516,N_2274);
or U3652 (N_3652,N_463,N_689);
and U3653 (N_3653,N_1701,N_1117);
nand U3654 (N_3654,N_1485,N_222);
or U3655 (N_3655,N_1597,N_1681);
and U3656 (N_3656,N_1400,N_59);
and U3657 (N_3657,N_132,N_1408);
nor U3658 (N_3658,N_646,N_1956);
nor U3659 (N_3659,N_1963,N_2176);
nor U3660 (N_3660,N_397,N_2158);
and U3661 (N_3661,N_2054,N_354);
and U3662 (N_3662,N_1884,N_786);
nor U3663 (N_3663,N_1659,N_1083);
and U3664 (N_3664,N_875,N_2253);
or U3665 (N_3665,N_1856,N_634);
or U3666 (N_3666,N_1877,N_429);
nor U3667 (N_3667,N_2344,N_2222);
nor U3668 (N_3668,N_1343,N_533);
nand U3669 (N_3669,N_104,N_196);
nand U3670 (N_3670,N_1846,N_2413);
nor U3671 (N_3671,N_1575,N_16);
and U3672 (N_3672,N_1387,N_1651);
nor U3673 (N_3673,N_1509,N_2419);
or U3674 (N_3674,N_2059,N_3);
nand U3675 (N_3675,N_422,N_1990);
nor U3676 (N_3676,N_802,N_1764);
nor U3677 (N_3677,N_701,N_1793);
or U3678 (N_3678,N_632,N_2083);
nor U3679 (N_3679,N_101,N_372);
nor U3680 (N_3680,N_628,N_394);
or U3681 (N_3681,N_823,N_2331);
or U3682 (N_3682,N_1890,N_1925);
xnor U3683 (N_3683,N_1838,N_1021);
xnor U3684 (N_3684,N_767,N_1082);
or U3685 (N_3685,N_1247,N_366);
and U3686 (N_3686,N_1646,N_853);
or U3687 (N_3687,N_1417,N_2489);
nand U3688 (N_3688,N_1949,N_1259);
nand U3689 (N_3689,N_805,N_2372);
or U3690 (N_3690,N_1876,N_1691);
or U3691 (N_3691,N_965,N_2243);
and U3692 (N_3692,N_67,N_514);
and U3693 (N_3693,N_1789,N_2070);
nor U3694 (N_3694,N_686,N_799);
and U3695 (N_3695,N_588,N_1440);
and U3696 (N_3696,N_1369,N_2324);
nand U3697 (N_3697,N_1415,N_1416);
or U3698 (N_3698,N_52,N_148);
nand U3699 (N_3699,N_1617,N_146);
and U3700 (N_3700,N_1086,N_178);
or U3701 (N_3701,N_1377,N_842);
or U3702 (N_3702,N_267,N_1958);
xnor U3703 (N_3703,N_2329,N_1032);
nor U3704 (N_3704,N_1251,N_125);
nand U3705 (N_3705,N_2276,N_1663);
and U3706 (N_3706,N_868,N_1505);
nor U3707 (N_3707,N_1355,N_1527);
or U3708 (N_3708,N_129,N_1512);
or U3709 (N_3709,N_896,N_1537);
nor U3710 (N_3710,N_1755,N_1319);
and U3711 (N_3711,N_866,N_2395);
or U3712 (N_3712,N_140,N_232);
nand U3713 (N_3713,N_2193,N_1397);
or U3714 (N_3714,N_660,N_1006);
nand U3715 (N_3715,N_1920,N_1688);
or U3716 (N_3716,N_2069,N_1119);
nor U3717 (N_3717,N_643,N_639);
and U3718 (N_3718,N_416,N_1048);
and U3719 (N_3719,N_1501,N_105);
xor U3720 (N_3720,N_2340,N_1459);
or U3721 (N_3721,N_332,N_733);
nor U3722 (N_3722,N_1093,N_593);
nor U3723 (N_3723,N_1591,N_825);
nor U3724 (N_3724,N_2424,N_2250);
or U3725 (N_3725,N_1602,N_324);
xor U3726 (N_3726,N_2349,N_454);
nor U3727 (N_3727,N_2061,N_1540);
xnor U3728 (N_3728,N_2361,N_90);
and U3729 (N_3729,N_56,N_1560);
or U3730 (N_3730,N_547,N_1849);
nor U3731 (N_3731,N_771,N_951);
nor U3732 (N_3732,N_2302,N_2452);
nand U3733 (N_3733,N_674,N_2476);
nor U3734 (N_3734,N_111,N_34);
xor U3735 (N_3735,N_2439,N_70);
or U3736 (N_3736,N_351,N_344);
or U3737 (N_3737,N_986,N_1535);
and U3738 (N_3738,N_1545,N_2305);
nand U3739 (N_3739,N_2278,N_58);
nand U3740 (N_3740,N_2064,N_937);
or U3741 (N_3741,N_1064,N_1577);
or U3742 (N_3742,N_914,N_1496);
or U3743 (N_3743,N_1580,N_193);
nand U3744 (N_3744,N_1473,N_1146);
or U3745 (N_3745,N_124,N_2323);
or U3746 (N_3746,N_1522,N_644);
and U3747 (N_3747,N_2076,N_716);
nor U3748 (N_3748,N_1077,N_605);
or U3749 (N_3749,N_732,N_2498);
nor U3750 (N_3750,N_96,N_1203);
and U3751 (N_3751,N_2148,N_2475);
or U3752 (N_3752,N_1457,N_2272);
nor U3753 (N_3753,N_1328,N_1352);
and U3754 (N_3754,N_687,N_1037);
nand U3755 (N_3755,N_1222,N_492);
nor U3756 (N_3756,N_379,N_1575);
and U3757 (N_3757,N_801,N_2461);
nor U3758 (N_3758,N_1719,N_1276);
and U3759 (N_3759,N_2489,N_1996);
and U3760 (N_3760,N_2270,N_2311);
or U3761 (N_3761,N_170,N_1900);
nor U3762 (N_3762,N_1044,N_1455);
nand U3763 (N_3763,N_1961,N_1504);
nand U3764 (N_3764,N_2075,N_160);
nand U3765 (N_3765,N_1415,N_1353);
nand U3766 (N_3766,N_2270,N_888);
nand U3767 (N_3767,N_950,N_2287);
or U3768 (N_3768,N_1264,N_1227);
and U3769 (N_3769,N_429,N_1194);
or U3770 (N_3770,N_2000,N_1227);
or U3771 (N_3771,N_1969,N_1914);
and U3772 (N_3772,N_1466,N_1379);
or U3773 (N_3773,N_1050,N_1435);
nand U3774 (N_3774,N_1272,N_941);
nor U3775 (N_3775,N_1970,N_75);
nand U3776 (N_3776,N_2386,N_1211);
nor U3777 (N_3777,N_2230,N_2460);
or U3778 (N_3778,N_1815,N_437);
and U3779 (N_3779,N_1642,N_1559);
nor U3780 (N_3780,N_546,N_1146);
and U3781 (N_3781,N_2477,N_2120);
or U3782 (N_3782,N_65,N_1653);
and U3783 (N_3783,N_1482,N_1058);
xor U3784 (N_3784,N_893,N_2259);
and U3785 (N_3785,N_281,N_1663);
nor U3786 (N_3786,N_751,N_2440);
or U3787 (N_3787,N_1094,N_609);
xnor U3788 (N_3788,N_2155,N_1650);
or U3789 (N_3789,N_1886,N_1707);
or U3790 (N_3790,N_67,N_1978);
and U3791 (N_3791,N_339,N_2054);
xor U3792 (N_3792,N_1676,N_426);
or U3793 (N_3793,N_1865,N_1331);
and U3794 (N_3794,N_1496,N_501);
and U3795 (N_3795,N_1259,N_156);
xnor U3796 (N_3796,N_249,N_2480);
and U3797 (N_3797,N_1348,N_2058);
or U3798 (N_3798,N_660,N_2438);
nand U3799 (N_3799,N_1080,N_529);
nand U3800 (N_3800,N_2222,N_1689);
or U3801 (N_3801,N_1403,N_1151);
and U3802 (N_3802,N_958,N_2222);
xor U3803 (N_3803,N_909,N_1823);
or U3804 (N_3804,N_1477,N_829);
nor U3805 (N_3805,N_1423,N_1372);
nor U3806 (N_3806,N_1119,N_1056);
nand U3807 (N_3807,N_1404,N_267);
nand U3808 (N_3808,N_1248,N_2198);
nand U3809 (N_3809,N_1246,N_2387);
xnor U3810 (N_3810,N_1288,N_177);
nand U3811 (N_3811,N_2134,N_446);
and U3812 (N_3812,N_811,N_2163);
or U3813 (N_3813,N_2384,N_1087);
nor U3814 (N_3814,N_820,N_292);
and U3815 (N_3815,N_1164,N_1041);
xnor U3816 (N_3816,N_77,N_1695);
xor U3817 (N_3817,N_1588,N_1574);
and U3818 (N_3818,N_1893,N_1961);
or U3819 (N_3819,N_1185,N_2320);
or U3820 (N_3820,N_367,N_1243);
nand U3821 (N_3821,N_1788,N_1087);
nand U3822 (N_3822,N_1746,N_2276);
xnor U3823 (N_3823,N_1847,N_2201);
and U3824 (N_3824,N_1151,N_33);
nand U3825 (N_3825,N_497,N_97);
nand U3826 (N_3826,N_699,N_1498);
nand U3827 (N_3827,N_1537,N_1800);
nor U3828 (N_3828,N_2206,N_504);
or U3829 (N_3829,N_2165,N_1560);
or U3830 (N_3830,N_1949,N_717);
or U3831 (N_3831,N_2148,N_2047);
and U3832 (N_3832,N_222,N_1413);
xor U3833 (N_3833,N_1120,N_133);
nor U3834 (N_3834,N_2330,N_1320);
nand U3835 (N_3835,N_353,N_85);
nor U3836 (N_3836,N_2003,N_142);
nor U3837 (N_3837,N_1837,N_902);
and U3838 (N_3838,N_842,N_24);
nand U3839 (N_3839,N_1838,N_307);
nand U3840 (N_3840,N_1945,N_1020);
nor U3841 (N_3841,N_825,N_337);
nor U3842 (N_3842,N_1838,N_43);
nor U3843 (N_3843,N_1725,N_1395);
nand U3844 (N_3844,N_324,N_656);
nor U3845 (N_3845,N_434,N_1427);
nor U3846 (N_3846,N_2202,N_1382);
nor U3847 (N_3847,N_2036,N_795);
nor U3848 (N_3848,N_1772,N_1293);
nor U3849 (N_3849,N_521,N_1939);
and U3850 (N_3850,N_182,N_1418);
nor U3851 (N_3851,N_1524,N_2314);
and U3852 (N_3852,N_101,N_1033);
and U3853 (N_3853,N_1152,N_441);
nor U3854 (N_3854,N_1161,N_1094);
nand U3855 (N_3855,N_44,N_1827);
and U3856 (N_3856,N_10,N_212);
or U3857 (N_3857,N_444,N_721);
nor U3858 (N_3858,N_1290,N_201);
nand U3859 (N_3859,N_1673,N_1285);
and U3860 (N_3860,N_1713,N_1925);
nand U3861 (N_3861,N_2052,N_1337);
nand U3862 (N_3862,N_1609,N_691);
or U3863 (N_3863,N_1061,N_1687);
nand U3864 (N_3864,N_926,N_1677);
nand U3865 (N_3865,N_1179,N_1427);
or U3866 (N_3866,N_2285,N_989);
xor U3867 (N_3867,N_276,N_1360);
and U3868 (N_3868,N_1301,N_478);
nand U3869 (N_3869,N_144,N_2383);
nor U3870 (N_3870,N_1000,N_1636);
nand U3871 (N_3871,N_524,N_1437);
xor U3872 (N_3872,N_1379,N_51);
nand U3873 (N_3873,N_1830,N_59);
nand U3874 (N_3874,N_1125,N_97);
or U3875 (N_3875,N_2218,N_1893);
or U3876 (N_3876,N_2364,N_631);
and U3877 (N_3877,N_288,N_919);
and U3878 (N_3878,N_403,N_1492);
nor U3879 (N_3879,N_296,N_1425);
nor U3880 (N_3880,N_1261,N_897);
nand U3881 (N_3881,N_1821,N_427);
and U3882 (N_3882,N_570,N_43);
nand U3883 (N_3883,N_825,N_1945);
nand U3884 (N_3884,N_401,N_705);
nand U3885 (N_3885,N_1020,N_1485);
and U3886 (N_3886,N_1160,N_258);
nand U3887 (N_3887,N_384,N_2453);
nor U3888 (N_3888,N_1453,N_1713);
xor U3889 (N_3889,N_2165,N_1295);
nand U3890 (N_3890,N_2332,N_1351);
or U3891 (N_3891,N_1256,N_286);
xnor U3892 (N_3892,N_1622,N_931);
nor U3893 (N_3893,N_2114,N_1144);
nor U3894 (N_3894,N_141,N_1717);
and U3895 (N_3895,N_251,N_50);
nand U3896 (N_3896,N_585,N_102);
nor U3897 (N_3897,N_2379,N_2457);
xnor U3898 (N_3898,N_757,N_1866);
and U3899 (N_3899,N_2096,N_672);
or U3900 (N_3900,N_1879,N_1028);
nand U3901 (N_3901,N_579,N_1977);
nor U3902 (N_3902,N_2437,N_247);
and U3903 (N_3903,N_2147,N_2278);
nor U3904 (N_3904,N_1182,N_352);
or U3905 (N_3905,N_2424,N_852);
nand U3906 (N_3906,N_2351,N_2169);
or U3907 (N_3907,N_2149,N_1151);
or U3908 (N_3908,N_319,N_1305);
or U3909 (N_3909,N_1556,N_2301);
or U3910 (N_3910,N_1854,N_1577);
nand U3911 (N_3911,N_253,N_818);
and U3912 (N_3912,N_1318,N_631);
nor U3913 (N_3913,N_2358,N_1719);
nand U3914 (N_3914,N_202,N_291);
and U3915 (N_3915,N_984,N_1708);
or U3916 (N_3916,N_136,N_927);
nand U3917 (N_3917,N_1822,N_2253);
xor U3918 (N_3918,N_816,N_1079);
nand U3919 (N_3919,N_2225,N_346);
or U3920 (N_3920,N_1586,N_1276);
or U3921 (N_3921,N_473,N_2187);
or U3922 (N_3922,N_517,N_816);
xor U3923 (N_3923,N_2324,N_225);
nand U3924 (N_3924,N_1056,N_28);
nand U3925 (N_3925,N_2444,N_2158);
or U3926 (N_3926,N_522,N_1809);
nand U3927 (N_3927,N_1625,N_1566);
and U3928 (N_3928,N_2059,N_265);
and U3929 (N_3929,N_1391,N_1203);
nand U3930 (N_3930,N_1218,N_321);
and U3931 (N_3931,N_2291,N_1725);
nor U3932 (N_3932,N_36,N_1617);
or U3933 (N_3933,N_1401,N_599);
nand U3934 (N_3934,N_1472,N_999);
and U3935 (N_3935,N_317,N_2383);
nor U3936 (N_3936,N_2034,N_1766);
and U3937 (N_3937,N_1159,N_1178);
nor U3938 (N_3938,N_581,N_656);
nand U3939 (N_3939,N_958,N_1878);
and U3940 (N_3940,N_1939,N_268);
or U3941 (N_3941,N_173,N_2021);
nor U3942 (N_3942,N_2437,N_407);
nand U3943 (N_3943,N_2273,N_1238);
nand U3944 (N_3944,N_808,N_41);
nand U3945 (N_3945,N_117,N_1601);
and U3946 (N_3946,N_1239,N_1139);
nor U3947 (N_3947,N_1773,N_1892);
nor U3948 (N_3948,N_1679,N_857);
or U3949 (N_3949,N_1862,N_598);
or U3950 (N_3950,N_827,N_1859);
nor U3951 (N_3951,N_686,N_529);
and U3952 (N_3952,N_1298,N_2347);
or U3953 (N_3953,N_1164,N_1174);
nand U3954 (N_3954,N_740,N_270);
nand U3955 (N_3955,N_2260,N_1820);
nor U3956 (N_3956,N_336,N_531);
xnor U3957 (N_3957,N_594,N_863);
xnor U3958 (N_3958,N_1332,N_2317);
or U3959 (N_3959,N_235,N_108);
and U3960 (N_3960,N_2033,N_28);
and U3961 (N_3961,N_2395,N_345);
xor U3962 (N_3962,N_705,N_1662);
nand U3963 (N_3963,N_33,N_2104);
and U3964 (N_3964,N_1601,N_608);
and U3965 (N_3965,N_708,N_661);
nand U3966 (N_3966,N_1782,N_2312);
and U3967 (N_3967,N_828,N_1433);
and U3968 (N_3968,N_1031,N_2118);
nor U3969 (N_3969,N_417,N_1108);
or U3970 (N_3970,N_1768,N_1774);
or U3971 (N_3971,N_1667,N_110);
nor U3972 (N_3972,N_1885,N_411);
or U3973 (N_3973,N_931,N_29);
nor U3974 (N_3974,N_1465,N_2091);
xnor U3975 (N_3975,N_294,N_2334);
xnor U3976 (N_3976,N_1901,N_1098);
or U3977 (N_3977,N_1774,N_1913);
and U3978 (N_3978,N_510,N_183);
xnor U3979 (N_3979,N_1872,N_525);
and U3980 (N_3980,N_2372,N_1530);
and U3981 (N_3981,N_1692,N_1240);
nand U3982 (N_3982,N_398,N_1);
nand U3983 (N_3983,N_1875,N_2052);
xor U3984 (N_3984,N_2351,N_2467);
or U3985 (N_3985,N_2146,N_2050);
nor U3986 (N_3986,N_960,N_171);
nand U3987 (N_3987,N_2295,N_1322);
nand U3988 (N_3988,N_1221,N_348);
nand U3989 (N_3989,N_870,N_1461);
nand U3990 (N_3990,N_2412,N_1802);
nand U3991 (N_3991,N_2,N_1022);
or U3992 (N_3992,N_2068,N_2165);
and U3993 (N_3993,N_202,N_1048);
or U3994 (N_3994,N_1694,N_497);
and U3995 (N_3995,N_1441,N_532);
or U3996 (N_3996,N_471,N_1744);
nor U3997 (N_3997,N_1500,N_2224);
nand U3998 (N_3998,N_923,N_1818);
and U3999 (N_3999,N_1050,N_1457);
nand U4000 (N_4000,N_368,N_1894);
and U4001 (N_4001,N_1241,N_1130);
nor U4002 (N_4002,N_2273,N_1747);
xnor U4003 (N_4003,N_657,N_292);
nand U4004 (N_4004,N_5,N_1625);
nor U4005 (N_4005,N_1039,N_290);
and U4006 (N_4006,N_467,N_1748);
nand U4007 (N_4007,N_2264,N_702);
and U4008 (N_4008,N_1801,N_2320);
nand U4009 (N_4009,N_836,N_2210);
and U4010 (N_4010,N_2070,N_233);
and U4011 (N_4011,N_315,N_454);
and U4012 (N_4012,N_1285,N_1712);
and U4013 (N_4013,N_1381,N_1491);
and U4014 (N_4014,N_1336,N_333);
and U4015 (N_4015,N_1957,N_2004);
or U4016 (N_4016,N_437,N_1363);
xor U4017 (N_4017,N_1226,N_148);
nand U4018 (N_4018,N_150,N_1745);
or U4019 (N_4019,N_872,N_2446);
nor U4020 (N_4020,N_477,N_826);
nor U4021 (N_4021,N_1309,N_2426);
nand U4022 (N_4022,N_1886,N_881);
or U4023 (N_4023,N_271,N_2264);
nor U4024 (N_4024,N_2008,N_439);
and U4025 (N_4025,N_2126,N_131);
and U4026 (N_4026,N_1097,N_199);
nor U4027 (N_4027,N_1653,N_2007);
xnor U4028 (N_4028,N_221,N_318);
and U4029 (N_4029,N_1336,N_1606);
or U4030 (N_4030,N_1632,N_764);
nor U4031 (N_4031,N_1057,N_1245);
nand U4032 (N_4032,N_1269,N_1569);
and U4033 (N_4033,N_2396,N_2053);
xnor U4034 (N_4034,N_528,N_2440);
or U4035 (N_4035,N_474,N_1172);
or U4036 (N_4036,N_307,N_808);
and U4037 (N_4037,N_1030,N_1884);
nand U4038 (N_4038,N_1146,N_2091);
nand U4039 (N_4039,N_470,N_378);
or U4040 (N_4040,N_2254,N_102);
nand U4041 (N_4041,N_694,N_1643);
xor U4042 (N_4042,N_297,N_512);
nand U4043 (N_4043,N_544,N_242);
or U4044 (N_4044,N_2488,N_2426);
and U4045 (N_4045,N_2249,N_552);
and U4046 (N_4046,N_2402,N_335);
and U4047 (N_4047,N_2180,N_1687);
or U4048 (N_4048,N_1098,N_680);
and U4049 (N_4049,N_294,N_772);
xnor U4050 (N_4050,N_1371,N_37);
nand U4051 (N_4051,N_328,N_1684);
nand U4052 (N_4052,N_2390,N_1783);
xor U4053 (N_4053,N_559,N_576);
nand U4054 (N_4054,N_1242,N_2199);
xor U4055 (N_4055,N_791,N_1369);
nor U4056 (N_4056,N_2420,N_661);
nor U4057 (N_4057,N_2088,N_1519);
nand U4058 (N_4058,N_243,N_2489);
or U4059 (N_4059,N_2482,N_79);
and U4060 (N_4060,N_1853,N_430);
nor U4061 (N_4061,N_2043,N_2025);
or U4062 (N_4062,N_785,N_2272);
and U4063 (N_4063,N_2200,N_565);
xor U4064 (N_4064,N_2451,N_1398);
nand U4065 (N_4065,N_1909,N_105);
nand U4066 (N_4066,N_1462,N_1840);
or U4067 (N_4067,N_522,N_90);
nand U4068 (N_4068,N_1981,N_2109);
and U4069 (N_4069,N_801,N_663);
nor U4070 (N_4070,N_1489,N_1249);
nand U4071 (N_4071,N_4,N_1520);
nor U4072 (N_4072,N_1767,N_2329);
nor U4073 (N_4073,N_452,N_261);
or U4074 (N_4074,N_1062,N_2151);
or U4075 (N_4075,N_1195,N_476);
nor U4076 (N_4076,N_2150,N_1685);
and U4077 (N_4077,N_933,N_360);
nand U4078 (N_4078,N_1773,N_1335);
nor U4079 (N_4079,N_1794,N_6);
nor U4080 (N_4080,N_1735,N_978);
and U4081 (N_4081,N_1763,N_2230);
nand U4082 (N_4082,N_1229,N_1568);
and U4083 (N_4083,N_1376,N_811);
and U4084 (N_4084,N_1701,N_162);
or U4085 (N_4085,N_1640,N_1739);
nor U4086 (N_4086,N_2275,N_1524);
and U4087 (N_4087,N_1381,N_989);
nor U4088 (N_4088,N_1702,N_2244);
and U4089 (N_4089,N_1188,N_1417);
and U4090 (N_4090,N_1297,N_2209);
nor U4091 (N_4091,N_179,N_1310);
nand U4092 (N_4092,N_2060,N_81);
xor U4093 (N_4093,N_1892,N_1578);
nand U4094 (N_4094,N_725,N_1725);
nand U4095 (N_4095,N_141,N_118);
and U4096 (N_4096,N_2030,N_1862);
nand U4097 (N_4097,N_2188,N_1724);
and U4098 (N_4098,N_608,N_73);
and U4099 (N_4099,N_2022,N_2494);
nor U4100 (N_4100,N_753,N_1879);
nor U4101 (N_4101,N_2107,N_56);
and U4102 (N_4102,N_759,N_2455);
xnor U4103 (N_4103,N_1146,N_1675);
nor U4104 (N_4104,N_1268,N_2204);
nor U4105 (N_4105,N_1997,N_798);
and U4106 (N_4106,N_24,N_1531);
and U4107 (N_4107,N_644,N_1657);
or U4108 (N_4108,N_290,N_842);
nor U4109 (N_4109,N_2175,N_1305);
nand U4110 (N_4110,N_949,N_1580);
nor U4111 (N_4111,N_449,N_892);
nand U4112 (N_4112,N_215,N_1643);
and U4113 (N_4113,N_294,N_2340);
nand U4114 (N_4114,N_737,N_333);
nand U4115 (N_4115,N_102,N_463);
nand U4116 (N_4116,N_15,N_1563);
nor U4117 (N_4117,N_712,N_454);
and U4118 (N_4118,N_1629,N_386);
or U4119 (N_4119,N_1575,N_2451);
nand U4120 (N_4120,N_673,N_2374);
or U4121 (N_4121,N_1452,N_772);
or U4122 (N_4122,N_2126,N_414);
nor U4123 (N_4123,N_1489,N_325);
nor U4124 (N_4124,N_2151,N_934);
nor U4125 (N_4125,N_45,N_227);
nand U4126 (N_4126,N_1021,N_137);
nand U4127 (N_4127,N_2095,N_1950);
nand U4128 (N_4128,N_731,N_1024);
nand U4129 (N_4129,N_1475,N_1783);
xor U4130 (N_4130,N_675,N_904);
nor U4131 (N_4131,N_1906,N_953);
nor U4132 (N_4132,N_556,N_1099);
nand U4133 (N_4133,N_1767,N_1452);
nor U4134 (N_4134,N_357,N_1476);
or U4135 (N_4135,N_1284,N_518);
and U4136 (N_4136,N_1015,N_2326);
nand U4137 (N_4137,N_1415,N_1024);
nor U4138 (N_4138,N_1667,N_1214);
and U4139 (N_4139,N_2085,N_1482);
or U4140 (N_4140,N_865,N_2376);
xor U4141 (N_4141,N_870,N_1918);
nand U4142 (N_4142,N_2330,N_842);
nand U4143 (N_4143,N_377,N_721);
and U4144 (N_4144,N_1797,N_1354);
nand U4145 (N_4145,N_2495,N_2463);
and U4146 (N_4146,N_2205,N_708);
nor U4147 (N_4147,N_140,N_801);
nor U4148 (N_4148,N_660,N_411);
or U4149 (N_4149,N_1588,N_1828);
or U4150 (N_4150,N_1561,N_786);
nand U4151 (N_4151,N_2185,N_521);
nor U4152 (N_4152,N_532,N_2168);
nand U4153 (N_4153,N_1316,N_1293);
xor U4154 (N_4154,N_2374,N_1859);
nor U4155 (N_4155,N_1077,N_2267);
or U4156 (N_4156,N_57,N_679);
nor U4157 (N_4157,N_2,N_181);
or U4158 (N_4158,N_1226,N_1090);
and U4159 (N_4159,N_967,N_350);
nor U4160 (N_4160,N_2058,N_166);
or U4161 (N_4161,N_2381,N_1794);
xnor U4162 (N_4162,N_492,N_840);
or U4163 (N_4163,N_106,N_1469);
and U4164 (N_4164,N_1573,N_2044);
nor U4165 (N_4165,N_289,N_1320);
xor U4166 (N_4166,N_847,N_1381);
nand U4167 (N_4167,N_1589,N_1959);
nand U4168 (N_4168,N_46,N_2181);
nand U4169 (N_4169,N_57,N_1343);
nand U4170 (N_4170,N_2480,N_1430);
or U4171 (N_4171,N_700,N_154);
nor U4172 (N_4172,N_1672,N_1009);
nand U4173 (N_4173,N_160,N_1207);
or U4174 (N_4174,N_943,N_113);
or U4175 (N_4175,N_1788,N_28);
and U4176 (N_4176,N_2306,N_2459);
and U4177 (N_4177,N_1077,N_1510);
or U4178 (N_4178,N_2042,N_1696);
nor U4179 (N_4179,N_1712,N_1617);
or U4180 (N_4180,N_533,N_2108);
nor U4181 (N_4181,N_1569,N_729);
or U4182 (N_4182,N_275,N_2064);
xnor U4183 (N_4183,N_1488,N_1583);
or U4184 (N_4184,N_903,N_1240);
or U4185 (N_4185,N_1269,N_1967);
and U4186 (N_4186,N_1836,N_258);
nand U4187 (N_4187,N_825,N_2023);
nand U4188 (N_4188,N_658,N_1715);
and U4189 (N_4189,N_1806,N_2195);
xor U4190 (N_4190,N_1106,N_724);
nor U4191 (N_4191,N_2359,N_1242);
and U4192 (N_4192,N_2461,N_722);
and U4193 (N_4193,N_1060,N_357);
and U4194 (N_4194,N_571,N_1342);
nor U4195 (N_4195,N_1933,N_1385);
nor U4196 (N_4196,N_2018,N_1525);
or U4197 (N_4197,N_875,N_2414);
nand U4198 (N_4198,N_1732,N_1173);
nand U4199 (N_4199,N_2327,N_2384);
and U4200 (N_4200,N_2201,N_1580);
nand U4201 (N_4201,N_244,N_1870);
or U4202 (N_4202,N_783,N_1137);
nand U4203 (N_4203,N_846,N_1265);
nand U4204 (N_4204,N_508,N_1710);
and U4205 (N_4205,N_2294,N_1218);
nand U4206 (N_4206,N_319,N_1148);
or U4207 (N_4207,N_771,N_1169);
nor U4208 (N_4208,N_572,N_762);
and U4209 (N_4209,N_2390,N_899);
nor U4210 (N_4210,N_467,N_1980);
nor U4211 (N_4211,N_116,N_2479);
nand U4212 (N_4212,N_1344,N_2005);
and U4213 (N_4213,N_2078,N_724);
and U4214 (N_4214,N_1340,N_419);
or U4215 (N_4215,N_2077,N_13);
and U4216 (N_4216,N_604,N_1871);
and U4217 (N_4217,N_1550,N_1618);
nor U4218 (N_4218,N_2106,N_498);
nor U4219 (N_4219,N_828,N_497);
or U4220 (N_4220,N_49,N_2350);
or U4221 (N_4221,N_1060,N_1336);
nor U4222 (N_4222,N_1263,N_2271);
xnor U4223 (N_4223,N_155,N_1537);
nand U4224 (N_4224,N_2412,N_852);
nor U4225 (N_4225,N_992,N_1502);
xnor U4226 (N_4226,N_548,N_2493);
nor U4227 (N_4227,N_603,N_2447);
and U4228 (N_4228,N_2343,N_841);
and U4229 (N_4229,N_625,N_413);
and U4230 (N_4230,N_277,N_2462);
nor U4231 (N_4231,N_2076,N_1395);
nand U4232 (N_4232,N_942,N_2068);
or U4233 (N_4233,N_125,N_194);
nand U4234 (N_4234,N_2342,N_1581);
nor U4235 (N_4235,N_336,N_1408);
and U4236 (N_4236,N_1785,N_617);
or U4237 (N_4237,N_683,N_1863);
or U4238 (N_4238,N_1408,N_344);
and U4239 (N_4239,N_1212,N_1771);
or U4240 (N_4240,N_2205,N_78);
or U4241 (N_4241,N_2061,N_1622);
xor U4242 (N_4242,N_2051,N_2466);
nand U4243 (N_4243,N_1579,N_582);
or U4244 (N_4244,N_933,N_1020);
nor U4245 (N_4245,N_2401,N_378);
or U4246 (N_4246,N_1082,N_327);
nor U4247 (N_4247,N_2384,N_897);
nor U4248 (N_4248,N_1093,N_222);
nor U4249 (N_4249,N_1539,N_1364);
nor U4250 (N_4250,N_1324,N_2370);
and U4251 (N_4251,N_2046,N_1433);
xnor U4252 (N_4252,N_1818,N_2068);
nand U4253 (N_4253,N_1306,N_954);
and U4254 (N_4254,N_380,N_1425);
nand U4255 (N_4255,N_1248,N_1691);
xor U4256 (N_4256,N_379,N_233);
or U4257 (N_4257,N_2122,N_1271);
nor U4258 (N_4258,N_1252,N_691);
nand U4259 (N_4259,N_1840,N_1275);
nand U4260 (N_4260,N_364,N_2362);
nand U4261 (N_4261,N_177,N_2388);
nor U4262 (N_4262,N_744,N_1668);
and U4263 (N_4263,N_176,N_1699);
nor U4264 (N_4264,N_2355,N_2135);
xor U4265 (N_4265,N_1675,N_95);
and U4266 (N_4266,N_1042,N_113);
or U4267 (N_4267,N_1250,N_142);
or U4268 (N_4268,N_570,N_1980);
or U4269 (N_4269,N_770,N_791);
or U4270 (N_4270,N_1654,N_2065);
and U4271 (N_4271,N_767,N_844);
nand U4272 (N_4272,N_1110,N_742);
and U4273 (N_4273,N_67,N_2343);
or U4274 (N_4274,N_1975,N_2286);
nor U4275 (N_4275,N_1192,N_1478);
xnor U4276 (N_4276,N_291,N_1501);
and U4277 (N_4277,N_531,N_1646);
nand U4278 (N_4278,N_647,N_1642);
nand U4279 (N_4279,N_666,N_2363);
nand U4280 (N_4280,N_2115,N_1276);
nand U4281 (N_4281,N_1571,N_1498);
or U4282 (N_4282,N_1658,N_1774);
or U4283 (N_4283,N_775,N_683);
and U4284 (N_4284,N_1720,N_1983);
or U4285 (N_4285,N_1592,N_837);
and U4286 (N_4286,N_169,N_2376);
and U4287 (N_4287,N_2290,N_713);
nand U4288 (N_4288,N_2227,N_952);
nor U4289 (N_4289,N_1897,N_376);
xor U4290 (N_4290,N_1805,N_1519);
nand U4291 (N_4291,N_2396,N_1555);
nor U4292 (N_4292,N_1779,N_2360);
nand U4293 (N_4293,N_533,N_1055);
or U4294 (N_4294,N_1333,N_1860);
or U4295 (N_4295,N_2171,N_2425);
nor U4296 (N_4296,N_1872,N_207);
xor U4297 (N_4297,N_1753,N_1146);
nor U4298 (N_4298,N_1060,N_2011);
and U4299 (N_4299,N_1821,N_1233);
nor U4300 (N_4300,N_1178,N_837);
and U4301 (N_4301,N_2297,N_2131);
nor U4302 (N_4302,N_2235,N_335);
or U4303 (N_4303,N_790,N_960);
or U4304 (N_4304,N_410,N_2059);
and U4305 (N_4305,N_1837,N_1204);
and U4306 (N_4306,N_1125,N_1844);
and U4307 (N_4307,N_715,N_1730);
and U4308 (N_4308,N_1098,N_1432);
nand U4309 (N_4309,N_1547,N_1149);
or U4310 (N_4310,N_2429,N_1151);
nor U4311 (N_4311,N_1747,N_2206);
nor U4312 (N_4312,N_550,N_978);
nor U4313 (N_4313,N_34,N_2122);
or U4314 (N_4314,N_254,N_1811);
nor U4315 (N_4315,N_2494,N_1805);
and U4316 (N_4316,N_1343,N_689);
nand U4317 (N_4317,N_2424,N_1613);
or U4318 (N_4318,N_338,N_1625);
xor U4319 (N_4319,N_2168,N_1190);
xor U4320 (N_4320,N_527,N_1823);
xnor U4321 (N_4321,N_622,N_244);
and U4322 (N_4322,N_95,N_568);
nor U4323 (N_4323,N_295,N_503);
or U4324 (N_4324,N_600,N_1050);
nand U4325 (N_4325,N_1475,N_1115);
nand U4326 (N_4326,N_1699,N_795);
or U4327 (N_4327,N_1200,N_1309);
and U4328 (N_4328,N_1154,N_244);
nor U4329 (N_4329,N_1779,N_1180);
nor U4330 (N_4330,N_1631,N_2411);
nor U4331 (N_4331,N_1366,N_2490);
nor U4332 (N_4332,N_1253,N_1871);
or U4333 (N_4333,N_2452,N_107);
and U4334 (N_4334,N_2089,N_741);
nor U4335 (N_4335,N_1153,N_2335);
nor U4336 (N_4336,N_1511,N_1385);
nor U4337 (N_4337,N_1808,N_1557);
xor U4338 (N_4338,N_1842,N_170);
nor U4339 (N_4339,N_1064,N_1420);
nor U4340 (N_4340,N_1120,N_1574);
and U4341 (N_4341,N_1719,N_2279);
nand U4342 (N_4342,N_1072,N_1122);
nor U4343 (N_4343,N_2030,N_1131);
or U4344 (N_4344,N_2497,N_1150);
or U4345 (N_4345,N_2278,N_1999);
nand U4346 (N_4346,N_966,N_317);
and U4347 (N_4347,N_1915,N_2142);
nor U4348 (N_4348,N_1564,N_1457);
nor U4349 (N_4349,N_715,N_1866);
nor U4350 (N_4350,N_2187,N_1331);
nor U4351 (N_4351,N_1577,N_1725);
nor U4352 (N_4352,N_83,N_2163);
and U4353 (N_4353,N_1664,N_1501);
or U4354 (N_4354,N_780,N_567);
and U4355 (N_4355,N_76,N_1057);
xnor U4356 (N_4356,N_2489,N_2030);
nand U4357 (N_4357,N_1406,N_2383);
nand U4358 (N_4358,N_742,N_2347);
or U4359 (N_4359,N_1573,N_1862);
nor U4360 (N_4360,N_953,N_611);
or U4361 (N_4361,N_2242,N_40);
nor U4362 (N_4362,N_1386,N_1110);
nand U4363 (N_4363,N_484,N_1606);
xnor U4364 (N_4364,N_151,N_2191);
xnor U4365 (N_4365,N_93,N_351);
or U4366 (N_4366,N_1394,N_1907);
or U4367 (N_4367,N_1065,N_113);
or U4368 (N_4368,N_742,N_93);
nand U4369 (N_4369,N_1555,N_1493);
nor U4370 (N_4370,N_1,N_1856);
nand U4371 (N_4371,N_1126,N_2273);
nor U4372 (N_4372,N_1838,N_2013);
nand U4373 (N_4373,N_2172,N_2460);
nor U4374 (N_4374,N_62,N_466);
or U4375 (N_4375,N_489,N_580);
nand U4376 (N_4376,N_1460,N_1744);
and U4377 (N_4377,N_1700,N_1813);
and U4378 (N_4378,N_1286,N_2153);
or U4379 (N_4379,N_187,N_1696);
nand U4380 (N_4380,N_16,N_883);
or U4381 (N_4381,N_1951,N_1892);
or U4382 (N_4382,N_816,N_83);
and U4383 (N_4383,N_2025,N_63);
or U4384 (N_4384,N_1296,N_1782);
nand U4385 (N_4385,N_1501,N_2380);
nand U4386 (N_4386,N_2434,N_677);
nor U4387 (N_4387,N_944,N_2111);
xor U4388 (N_4388,N_984,N_360);
or U4389 (N_4389,N_656,N_2174);
and U4390 (N_4390,N_1957,N_386);
nand U4391 (N_4391,N_1847,N_1437);
and U4392 (N_4392,N_667,N_2219);
nor U4393 (N_4393,N_338,N_1955);
xor U4394 (N_4394,N_2383,N_1320);
nand U4395 (N_4395,N_83,N_1972);
nor U4396 (N_4396,N_1570,N_427);
xnor U4397 (N_4397,N_1264,N_2227);
or U4398 (N_4398,N_1846,N_2095);
and U4399 (N_4399,N_1099,N_2196);
and U4400 (N_4400,N_163,N_381);
nand U4401 (N_4401,N_1527,N_1016);
and U4402 (N_4402,N_1261,N_2194);
and U4403 (N_4403,N_279,N_1107);
nor U4404 (N_4404,N_1473,N_1863);
nor U4405 (N_4405,N_2067,N_2358);
nand U4406 (N_4406,N_1176,N_2046);
and U4407 (N_4407,N_2037,N_1114);
nand U4408 (N_4408,N_1386,N_1633);
nand U4409 (N_4409,N_396,N_1811);
or U4410 (N_4410,N_2104,N_2331);
or U4411 (N_4411,N_1096,N_1073);
or U4412 (N_4412,N_2075,N_965);
or U4413 (N_4413,N_1142,N_59);
or U4414 (N_4414,N_264,N_2321);
nor U4415 (N_4415,N_493,N_749);
xnor U4416 (N_4416,N_855,N_2494);
or U4417 (N_4417,N_552,N_14);
or U4418 (N_4418,N_1994,N_899);
nor U4419 (N_4419,N_1862,N_2094);
nor U4420 (N_4420,N_2493,N_296);
and U4421 (N_4421,N_1712,N_1964);
and U4422 (N_4422,N_1879,N_734);
xor U4423 (N_4423,N_1292,N_1072);
nand U4424 (N_4424,N_1204,N_286);
nor U4425 (N_4425,N_1227,N_964);
and U4426 (N_4426,N_1410,N_788);
and U4427 (N_4427,N_1213,N_1293);
nand U4428 (N_4428,N_1818,N_1903);
and U4429 (N_4429,N_601,N_2325);
nor U4430 (N_4430,N_726,N_113);
nor U4431 (N_4431,N_642,N_1698);
and U4432 (N_4432,N_1418,N_1534);
or U4433 (N_4433,N_119,N_1408);
and U4434 (N_4434,N_44,N_964);
nand U4435 (N_4435,N_1092,N_1428);
xnor U4436 (N_4436,N_2259,N_1593);
nand U4437 (N_4437,N_2024,N_405);
or U4438 (N_4438,N_765,N_435);
nand U4439 (N_4439,N_1634,N_1927);
xor U4440 (N_4440,N_1894,N_2126);
xnor U4441 (N_4441,N_1206,N_2039);
and U4442 (N_4442,N_1023,N_2231);
and U4443 (N_4443,N_1953,N_2240);
nor U4444 (N_4444,N_13,N_38);
xor U4445 (N_4445,N_2042,N_67);
and U4446 (N_4446,N_1438,N_171);
xor U4447 (N_4447,N_2101,N_2264);
and U4448 (N_4448,N_1545,N_1503);
and U4449 (N_4449,N_1848,N_2179);
or U4450 (N_4450,N_465,N_140);
or U4451 (N_4451,N_1058,N_476);
nand U4452 (N_4452,N_1275,N_1375);
nand U4453 (N_4453,N_929,N_1726);
nor U4454 (N_4454,N_810,N_352);
or U4455 (N_4455,N_451,N_1274);
and U4456 (N_4456,N_1625,N_1016);
and U4457 (N_4457,N_1946,N_1088);
nand U4458 (N_4458,N_2031,N_95);
or U4459 (N_4459,N_2120,N_2417);
xor U4460 (N_4460,N_2379,N_324);
xnor U4461 (N_4461,N_1226,N_1696);
nand U4462 (N_4462,N_1318,N_2372);
nand U4463 (N_4463,N_1033,N_1524);
or U4464 (N_4464,N_305,N_1602);
xnor U4465 (N_4465,N_1231,N_1901);
nand U4466 (N_4466,N_1933,N_937);
nor U4467 (N_4467,N_673,N_2464);
xnor U4468 (N_4468,N_467,N_2248);
and U4469 (N_4469,N_1186,N_609);
nor U4470 (N_4470,N_1585,N_240);
or U4471 (N_4471,N_714,N_349);
xor U4472 (N_4472,N_2430,N_536);
and U4473 (N_4473,N_415,N_2365);
and U4474 (N_4474,N_543,N_807);
or U4475 (N_4475,N_1003,N_204);
nor U4476 (N_4476,N_639,N_1542);
nor U4477 (N_4477,N_388,N_1213);
nor U4478 (N_4478,N_545,N_666);
nand U4479 (N_4479,N_2419,N_641);
nand U4480 (N_4480,N_886,N_887);
xor U4481 (N_4481,N_2138,N_1282);
and U4482 (N_4482,N_2203,N_922);
or U4483 (N_4483,N_462,N_1056);
and U4484 (N_4484,N_137,N_319);
xnor U4485 (N_4485,N_1120,N_1213);
nand U4486 (N_4486,N_1307,N_2167);
xnor U4487 (N_4487,N_785,N_1013);
nor U4488 (N_4488,N_1193,N_1234);
or U4489 (N_4489,N_75,N_386);
nand U4490 (N_4490,N_1279,N_1685);
nor U4491 (N_4491,N_745,N_1943);
nor U4492 (N_4492,N_2182,N_2073);
or U4493 (N_4493,N_62,N_1684);
nor U4494 (N_4494,N_1599,N_1630);
or U4495 (N_4495,N_2486,N_503);
nor U4496 (N_4496,N_1195,N_13);
or U4497 (N_4497,N_2103,N_210);
and U4498 (N_4498,N_2319,N_1322);
or U4499 (N_4499,N_1546,N_1866);
or U4500 (N_4500,N_2096,N_1676);
nor U4501 (N_4501,N_313,N_1611);
nor U4502 (N_4502,N_895,N_16);
or U4503 (N_4503,N_171,N_1555);
xor U4504 (N_4504,N_262,N_967);
nand U4505 (N_4505,N_1011,N_490);
or U4506 (N_4506,N_824,N_2437);
or U4507 (N_4507,N_1402,N_1867);
xnor U4508 (N_4508,N_1861,N_1849);
nor U4509 (N_4509,N_1160,N_467);
xnor U4510 (N_4510,N_852,N_1010);
and U4511 (N_4511,N_2499,N_1657);
or U4512 (N_4512,N_1050,N_1261);
or U4513 (N_4513,N_1995,N_1662);
nor U4514 (N_4514,N_1548,N_194);
nor U4515 (N_4515,N_1739,N_970);
xor U4516 (N_4516,N_216,N_1967);
nor U4517 (N_4517,N_2199,N_1556);
nor U4518 (N_4518,N_961,N_822);
or U4519 (N_4519,N_640,N_962);
nand U4520 (N_4520,N_393,N_2057);
nor U4521 (N_4521,N_1803,N_599);
nand U4522 (N_4522,N_440,N_343);
nor U4523 (N_4523,N_1457,N_1188);
and U4524 (N_4524,N_1562,N_2201);
and U4525 (N_4525,N_176,N_593);
and U4526 (N_4526,N_1882,N_2376);
nand U4527 (N_4527,N_1183,N_579);
xor U4528 (N_4528,N_595,N_1073);
and U4529 (N_4529,N_669,N_1558);
nand U4530 (N_4530,N_1755,N_1426);
and U4531 (N_4531,N_537,N_2416);
nor U4532 (N_4532,N_2092,N_1094);
and U4533 (N_4533,N_1995,N_1298);
nor U4534 (N_4534,N_1008,N_1862);
and U4535 (N_4535,N_95,N_1574);
or U4536 (N_4536,N_2381,N_1622);
nor U4537 (N_4537,N_199,N_2082);
nor U4538 (N_4538,N_2446,N_2433);
xnor U4539 (N_4539,N_1607,N_1920);
or U4540 (N_4540,N_1503,N_1888);
xor U4541 (N_4541,N_1160,N_2308);
or U4542 (N_4542,N_2310,N_1356);
nand U4543 (N_4543,N_1645,N_100);
nand U4544 (N_4544,N_321,N_310);
xnor U4545 (N_4545,N_339,N_2138);
xnor U4546 (N_4546,N_1927,N_1683);
nor U4547 (N_4547,N_992,N_1981);
or U4548 (N_4548,N_161,N_1352);
or U4549 (N_4549,N_350,N_69);
and U4550 (N_4550,N_1646,N_1294);
nor U4551 (N_4551,N_1654,N_497);
nor U4552 (N_4552,N_2299,N_1625);
or U4553 (N_4553,N_2354,N_208);
nand U4554 (N_4554,N_636,N_1069);
and U4555 (N_4555,N_2104,N_1243);
or U4556 (N_4556,N_1382,N_2411);
nand U4557 (N_4557,N_1188,N_2477);
nand U4558 (N_4558,N_1890,N_960);
and U4559 (N_4559,N_1948,N_51);
nor U4560 (N_4560,N_1067,N_2247);
nor U4561 (N_4561,N_295,N_1957);
or U4562 (N_4562,N_2476,N_988);
nor U4563 (N_4563,N_255,N_2085);
nor U4564 (N_4564,N_704,N_1301);
nor U4565 (N_4565,N_628,N_791);
nor U4566 (N_4566,N_1264,N_840);
and U4567 (N_4567,N_1178,N_2169);
and U4568 (N_4568,N_583,N_1977);
or U4569 (N_4569,N_1111,N_1416);
nand U4570 (N_4570,N_883,N_1721);
and U4571 (N_4571,N_452,N_1031);
nor U4572 (N_4572,N_1868,N_814);
or U4573 (N_4573,N_2250,N_1438);
or U4574 (N_4574,N_1331,N_185);
nor U4575 (N_4575,N_2003,N_2430);
and U4576 (N_4576,N_2241,N_1025);
nand U4577 (N_4577,N_421,N_1088);
and U4578 (N_4578,N_764,N_116);
or U4579 (N_4579,N_1983,N_2483);
xor U4580 (N_4580,N_610,N_1071);
and U4581 (N_4581,N_1336,N_1485);
and U4582 (N_4582,N_2278,N_1094);
nor U4583 (N_4583,N_1025,N_1127);
and U4584 (N_4584,N_2495,N_2285);
nor U4585 (N_4585,N_2455,N_2287);
or U4586 (N_4586,N_1437,N_1058);
and U4587 (N_4587,N_1072,N_1715);
and U4588 (N_4588,N_937,N_1195);
or U4589 (N_4589,N_1960,N_1415);
and U4590 (N_4590,N_2150,N_1192);
and U4591 (N_4591,N_1308,N_1197);
nand U4592 (N_4592,N_2074,N_159);
or U4593 (N_4593,N_125,N_1467);
nand U4594 (N_4594,N_277,N_1261);
and U4595 (N_4595,N_1558,N_413);
nor U4596 (N_4596,N_1048,N_166);
or U4597 (N_4597,N_2417,N_271);
nor U4598 (N_4598,N_2422,N_1713);
nand U4599 (N_4599,N_1937,N_1079);
xnor U4600 (N_4600,N_154,N_1763);
nand U4601 (N_4601,N_381,N_1303);
and U4602 (N_4602,N_770,N_1660);
xnor U4603 (N_4603,N_1978,N_2043);
nand U4604 (N_4604,N_1439,N_373);
nand U4605 (N_4605,N_274,N_1424);
and U4606 (N_4606,N_1564,N_2073);
nand U4607 (N_4607,N_2230,N_120);
nand U4608 (N_4608,N_1867,N_1244);
nor U4609 (N_4609,N_1609,N_2003);
nand U4610 (N_4610,N_1770,N_792);
or U4611 (N_4611,N_822,N_308);
nor U4612 (N_4612,N_2398,N_2001);
nor U4613 (N_4613,N_842,N_2393);
and U4614 (N_4614,N_2440,N_462);
or U4615 (N_4615,N_593,N_947);
and U4616 (N_4616,N_105,N_1453);
or U4617 (N_4617,N_2205,N_1528);
or U4618 (N_4618,N_1502,N_1398);
and U4619 (N_4619,N_450,N_1278);
or U4620 (N_4620,N_2395,N_1662);
nor U4621 (N_4621,N_761,N_1785);
nand U4622 (N_4622,N_2269,N_27);
or U4623 (N_4623,N_2165,N_1734);
and U4624 (N_4624,N_939,N_1732);
or U4625 (N_4625,N_2284,N_2358);
or U4626 (N_4626,N_1242,N_4);
xor U4627 (N_4627,N_247,N_296);
nand U4628 (N_4628,N_1592,N_725);
xor U4629 (N_4629,N_1502,N_2222);
nand U4630 (N_4630,N_2231,N_1951);
and U4631 (N_4631,N_480,N_1379);
and U4632 (N_4632,N_1485,N_2432);
nand U4633 (N_4633,N_371,N_1099);
and U4634 (N_4634,N_1590,N_1386);
or U4635 (N_4635,N_1596,N_954);
and U4636 (N_4636,N_1260,N_2431);
nand U4637 (N_4637,N_1348,N_1499);
nand U4638 (N_4638,N_841,N_2296);
nand U4639 (N_4639,N_1231,N_2390);
or U4640 (N_4640,N_655,N_902);
or U4641 (N_4641,N_1134,N_514);
xnor U4642 (N_4642,N_1352,N_320);
xor U4643 (N_4643,N_1664,N_633);
nor U4644 (N_4644,N_2030,N_250);
or U4645 (N_4645,N_1569,N_2102);
nand U4646 (N_4646,N_1292,N_2112);
nor U4647 (N_4647,N_1484,N_650);
nand U4648 (N_4648,N_162,N_608);
or U4649 (N_4649,N_1495,N_1259);
and U4650 (N_4650,N_358,N_2305);
or U4651 (N_4651,N_432,N_815);
and U4652 (N_4652,N_496,N_873);
and U4653 (N_4653,N_137,N_93);
or U4654 (N_4654,N_8,N_1121);
or U4655 (N_4655,N_1997,N_1771);
and U4656 (N_4656,N_656,N_1229);
and U4657 (N_4657,N_93,N_1513);
and U4658 (N_4658,N_2365,N_1258);
and U4659 (N_4659,N_1486,N_1991);
xor U4660 (N_4660,N_375,N_264);
nand U4661 (N_4661,N_704,N_375);
and U4662 (N_4662,N_102,N_1723);
and U4663 (N_4663,N_1184,N_599);
and U4664 (N_4664,N_906,N_2282);
nor U4665 (N_4665,N_876,N_1635);
nand U4666 (N_4666,N_691,N_1760);
nor U4667 (N_4667,N_2346,N_2360);
or U4668 (N_4668,N_58,N_1240);
nand U4669 (N_4669,N_1244,N_2361);
nand U4670 (N_4670,N_408,N_678);
nand U4671 (N_4671,N_1044,N_1227);
xor U4672 (N_4672,N_12,N_1594);
and U4673 (N_4673,N_1526,N_408);
or U4674 (N_4674,N_1668,N_1597);
and U4675 (N_4675,N_1047,N_1190);
or U4676 (N_4676,N_1606,N_1936);
and U4677 (N_4677,N_1638,N_1681);
and U4678 (N_4678,N_933,N_1245);
and U4679 (N_4679,N_732,N_1812);
and U4680 (N_4680,N_517,N_1307);
or U4681 (N_4681,N_2241,N_2347);
nand U4682 (N_4682,N_609,N_365);
and U4683 (N_4683,N_2130,N_2084);
or U4684 (N_4684,N_2242,N_1586);
and U4685 (N_4685,N_2237,N_1846);
and U4686 (N_4686,N_91,N_533);
and U4687 (N_4687,N_126,N_866);
xnor U4688 (N_4688,N_1228,N_781);
or U4689 (N_4689,N_234,N_2228);
or U4690 (N_4690,N_1383,N_1230);
or U4691 (N_4691,N_1906,N_735);
and U4692 (N_4692,N_1717,N_1852);
or U4693 (N_4693,N_1522,N_942);
nor U4694 (N_4694,N_577,N_918);
and U4695 (N_4695,N_2243,N_2311);
and U4696 (N_4696,N_2488,N_2164);
nor U4697 (N_4697,N_1737,N_1523);
nand U4698 (N_4698,N_151,N_1770);
or U4699 (N_4699,N_2178,N_529);
nor U4700 (N_4700,N_1251,N_386);
or U4701 (N_4701,N_1338,N_1865);
or U4702 (N_4702,N_845,N_1731);
and U4703 (N_4703,N_124,N_1138);
nand U4704 (N_4704,N_2039,N_496);
or U4705 (N_4705,N_350,N_347);
or U4706 (N_4706,N_1481,N_1103);
and U4707 (N_4707,N_1129,N_2039);
xnor U4708 (N_4708,N_2484,N_273);
nand U4709 (N_4709,N_1704,N_2417);
or U4710 (N_4710,N_144,N_2268);
nand U4711 (N_4711,N_107,N_2273);
nor U4712 (N_4712,N_1473,N_317);
nor U4713 (N_4713,N_632,N_1206);
nand U4714 (N_4714,N_216,N_1387);
nor U4715 (N_4715,N_1300,N_330);
nand U4716 (N_4716,N_1368,N_1899);
or U4717 (N_4717,N_535,N_1883);
and U4718 (N_4718,N_1946,N_1260);
nand U4719 (N_4719,N_106,N_2411);
nand U4720 (N_4720,N_61,N_2115);
or U4721 (N_4721,N_1521,N_106);
nor U4722 (N_4722,N_506,N_643);
nand U4723 (N_4723,N_2020,N_1664);
and U4724 (N_4724,N_2168,N_866);
nand U4725 (N_4725,N_1424,N_1960);
nand U4726 (N_4726,N_1193,N_1667);
xnor U4727 (N_4727,N_110,N_804);
or U4728 (N_4728,N_415,N_2136);
and U4729 (N_4729,N_2083,N_523);
and U4730 (N_4730,N_1475,N_140);
nand U4731 (N_4731,N_1173,N_1936);
nor U4732 (N_4732,N_1572,N_2388);
and U4733 (N_4733,N_178,N_2072);
or U4734 (N_4734,N_1288,N_1242);
nor U4735 (N_4735,N_966,N_226);
or U4736 (N_4736,N_1933,N_1150);
or U4737 (N_4737,N_1767,N_1230);
nor U4738 (N_4738,N_498,N_1078);
nor U4739 (N_4739,N_255,N_1271);
and U4740 (N_4740,N_288,N_193);
nand U4741 (N_4741,N_1953,N_613);
nand U4742 (N_4742,N_1836,N_1965);
and U4743 (N_4743,N_1628,N_752);
nor U4744 (N_4744,N_814,N_1254);
nor U4745 (N_4745,N_2496,N_2427);
nand U4746 (N_4746,N_690,N_377);
nor U4747 (N_4747,N_1310,N_313);
and U4748 (N_4748,N_1612,N_522);
and U4749 (N_4749,N_1095,N_1384);
nand U4750 (N_4750,N_1440,N_199);
nand U4751 (N_4751,N_55,N_1157);
nor U4752 (N_4752,N_1471,N_351);
or U4753 (N_4753,N_1148,N_1716);
nand U4754 (N_4754,N_144,N_123);
or U4755 (N_4755,N_429,N_1529);
and U4756 (N_4756,N_720,N_1289);
or U4757 (N_4757,N_1659,N_1804);
or U4758 (N_4758,N_917,N_2036);
xor U4759 (N_4759,N_2129,N_25);
nor U4760 (N_4760,N_989,N_542);
nor U4761 (N_4761,N_2384,N_2074);
nand U4762 (N_4762,N_331,N_320);
nand U4763 (N_4763,N_1045,N_2418);
nand U4764 (N_4764,N_2240,N_1344);
or U4765 (N_4765,N_1729,N_1167);
nand U4766 (N_4766,N_1036,N_1740);
nand U4767 (N_4767,N_712,N_1796);
nand U4768 (N_4768,N_1955,N_638);
and U4769 (N_4769,N_269,N_405);
or U4770 (N_4770,N_766,N_590);
xnor U4771 (N_4771,N_1306,N_1);
or U4772 (N_4772,N_1499,N_545);
or U4773 (N_4773,N_1850,N_2445);
nor U4774 (N_4774,N_635,N_81);
or U4775 (N_4775,N_402,N_1799);
or U4776 (N_4776,N_164,N_1364);
or U4777 (N_4777,N_846,N_1364);
or U4778 (N_4778,N_429,N_915);
and U4779 (N_4779,N_205,N_1541);
xnor U4780 (N_4780,N_1717,N_487);
xor U4781 (N_4781,N_494,N_159);
nor U4782 (N_4782,N_2172,N_1971);
or U4783 (N_4783,N_1196,N_1835);
or U4784 (N_4784,N_2377,N_2222);
nand U4785 (N_4785,N_803,N_105);
nor U4786 (N_4786,N_758,N_145);
nor U4787 (N_4787,N_1711,N_2195);
xor U4788 (N_4788,N_410,N_1038);
nor U4789 (N_4789,N_1598,N_2372);
and U4790 (N_4790,N_1732,N_869);
or U4791 (N_4791,N_1439,N_2471);
or U4792 (N_4792,N_403,N_138);
nand U4793 (N_4793,N_2076,N_512);
nor U4794 (N_4794,N_2199,N_1880);
nand U4795 (N_4795,N_1126,N_1091);
or U4796 (N_4796,N_1494,N_2354);
nor U4797 (N_4797,N_1349,N_1627);
or U4798 (N_4798,N_1524,N_2048);
xnor U4799 (N_4799,N_851,N_1724);
xor U4800 (N_4800,N_1842,N_945);
or U4801 (N_4801,N_1152,N_1800);
nand U4802 (N_4802,N_412,N_2490);
xor U4803 (N_4803,N_1625,N_329);
nand U4804 (N_4804,N_530,N_1900);
or U4805 (N_4805,N_1780,N_836);
and U4806 (N_4806,N_2397,N_386);
xor U4807 (N_4807,N_603,N_725);
or U4808 (N_4808,N_990,N_1634);
or U4809 (N_4809,N_2466,N_967);
and U4810 (N_4810,N_403,N_2297);
or U4811 (N_4811,N_115,N_184);
or U4812 (N_4812,N_1008,N_268);
and U4813 (N_4813,N_2447,N_1305);
nand U4814 (N_4814,N_2243,N_932);
or U4815 (N_4815,N_1098,N_1021);
or U4816 (N_4816,N_2268,N_2096);
nand U4817 (N_4817,N_1617,N_554);
and U4818 (N_4818,N_1697,N_304);
nand U4819 (N_4819,N_1927,N_32);
nand U4820 (N_4820,N_2448,N_2236);
or U4821 (N_4821,N_1718,N_2272);
nand U4822 (N_4822,N_1470,N_2051);
and U4823 (N_4823,N_2432,N_2135);
nand U4824 (N_4824,N_1627,N_2453);
nor U4825 (N_4825,N_13,N_2267);
or U4826 (N_4826,N_2120,N_417);
or U4827 (N_4827,N_2498,N_1148);
nor U4828 (N_4828,N_1677,N_1093);
and U4829 (N_4829,N_317,N_99);
nand U4830 (N_4830,N_251,N_1366);
nor U4831 (N_4831,N_1895,N_1473);
or U4832 (N_4832,N_2475,N_1888);
or U4833 (N_4833,N_2112,N_1396);
and U4834 (N_4834,N_623,N_982);
nor U4835 (N_4835,N_1150,N_777);
nor U4836 (N_4836,N_1142,N_291);
nor U4837 (N_4837,N_575,N_939);
or U4838 (N_4838,N_276,N_165);
and U4839 (N_4839,N_590,N_1033);
and U4840 (N_4840,N_1555,N_2295);
nor U4841 (N_4841,N_974,N_141);
nand U4842 (N_4842,N_2485,N_1589);
or U4843 (N_4843,N_2225,N_1007);
xor U4844 (N_4844,N_2373,N_807);
nor U4845 (N_4845,N_85,N_1031);
nand U4846 (N_4846,N_1594,N_140);
or U4847 (N_4847,N_2481,N_1268);
nor U4848 (N_4848,N_1085,N_2431);
nor U4849 (N_4849,N_1250,N_1635);
nand U4850 (N_4850,N_245,N_597);
and U4851 (N_4851,N_87,N_471);
nand U4852 (N_4852,N_1884,N_2303);
xnor U4853 (N_4853,N_19,N_1567);
xor U4854 (N_4854,N_1665,N_1482);
nand U4855 (N_4855,N_2044,N_677);
nand U4856 (N_4856,N_2243,N_255);
nand U4857 (N_4857,N_1480,N_1982);
or U4858 (N_4858,N_1152,N_1472);
nand U4859 (N_4859,N_1386,N_1347);
xor U4860 (N_4860,N_453,N_2341);
or U4861 (N_4861,N_926,N_2408);
and U4862 (N_4862,N_309,N_2402);
nand U4863 (N_4863,N_1822,N_1299);
nand U4864 (N_4864,N_2302,N_851);
nand U4865 (N_4865,N_986,N_1593);
and U4866 (N_4866,N_224,N_158);
nor U4867 (N_4867,N_621,N_305);
nor U4868 (N_4868,N_440,N_2202);
xnor U4869 (N_4869,N_771,N_276);
nand U4870 (N_4870,N_1559,N_1319);
nor U4871 (N_4871,N_147,N_1674);
nor U4872 (N_4872,N_574,N_2179);
or U4873 (N_4873,N_1706,N_1827);
nor U4874 (N_4874,N_882,N_1586);
or U4875 (N_4875,N_888,N_716);
nor U4876 (N_4876,N_1847,N_537);
and U4877 (N_4877,N_904,N_785);
xor U4878 (N_4878,N_1138,N_1893);
nand U4879 (N_4879,N_449,N_863);
nor U4880 (N_4880,N_1922,N_245);
nor U4881 (N_4881,N_988,N_757);
and U4882 (N_4882,N_2230,N_525);
nor U4883 (N_4883,N_730,N_2316);
nand U4884 (N_4884,N_628,N_1743);
and U4885 (N_4885,N_196,N_1905);
nor U4886 (N_4886,N_1780,N_1674);
nor U4887 (N_4887,N_2309,N_1735);
and U4888 (N_4888,N_1438,N_1687);
nand U4889 (N_4889,N_957,N_1187);
nor U4890 (N_4890,N_318,N_2119);
and U4891 (N_4891,N_960,N_770);
and U4892 (N_4892,N_1844,N_816);
and U4893 (N_4893,N_1230,N_534);
or U4894 (N_4894,N_1608,N_240);
and U4895 (N_4895,N_849,N_2298);
xnor U4896 (N_4896,N_1149,N_164);
and U4897 (N_4897,N_1545,N_332);
nor U4898 (N_4898,N_2285,N_1763);
nand U4899 (N_4899,N_802,N_2332);
xor U4900 (N_4900,N_365,N_1775);
nor U4901 (N_4901,N_359,N_2082);
and U4902 (N_4902,N_472,N_2431);
nand U4903 (N_4903,N_1335,N_575);
nor U4904 (N_4904,N_1072,N_1253);
nand U4905 (N_4905,N_2277,N_1096);
or U4906 (N_4906,N_1328,N_1820);
xor U4907 (N_4907,N_1828,N_988);
xor U4908 (N_4908,N_2246,N_1055);
and U4909 (N_4909,N_2060,N_2493);
nand U4910 (N_4910,N_1309,N_406);
and U4911 (N_4911,N_773,N_1844);
and U4912 (N_4912,N_255,N_1669);
and U4913 (N_4913,N_1532,N_1658);
nand U4914 (N_4914,N_631,N_1824);
xnor U4915 (N_4915,N_2088,N_1116);
or U4916 (N_4916,N_1481,N_2161);
or U4917 (N_4917,N_1009,N_1334);
and U4918 (N_4918,N_1803,N_455);
or U4919 (N_4919,N_52,N_864);
xnor U4920 (N_4920,N_194,N_327);
or U4921 (N_4921,N_2281,N_283);
nand U4922 (N_4922,N_353,N_2220);
nor U4923 (N_4923,N_2447,N_212);
or U4924 (N_4924,N_1016,N_1949);
nand U4925 (N_4925,N_2438,N_547);
nor U4926 (N_4926,N_2103,N_953);
nand U4927 (N_4927,N_453,N_2031);
nand U4928 (N_4928,N_923,N_2042);
nand U4929 (N_4929,N_1704,N_2211);
nand U4930 (N_4930,N_686,N_1953);
xnor U4931 (N_4931,N_714,N_1299);
nor U4932 (N_4932,N_1695,N_1998);
or U4933 (N_4933,N_2165,N_220);
nand U4934 (N_4934,N_837,N_2182);
nand U4935 (N_4935,N_1010,N_2227);
or U4936 (N_4936,N_2018,N_2414);
and U4937 (N_4937,N_100,N_1063);
nand U4938 (N_4938,N_446,N_1818);
and U4939 (N_4939,N_475,N_215);
nand U4940 (N_4940,N_1703,N_317);
and U4941 (N_4941,N_471,N_1643);
nor U4942 (N_4942,N_529,N_997);
and U4943 (N_4943,N_2302,N_1813);
nor U4944 (N_4944,N_1522,N_1342);
nor U4945 (N_4945,N_2020,N_1652);
and U4946 (N_4946,N_2043,N_197);
nor U4947 (N_4947,N_1683,N_2048);
or U4948 (N_4948,N_1487,N_614);
nand U4949 (N_4949,N_311,N_1163);
nor U4950 (N_4950,N_1337,N_1226);
xor U4951 (N_4951,N_805,N_1230);
and U4952 (N_4952,N_200,N_2295);
nand U4953 (N_4953,N_629,N_340);
nand U4954 (N_4954,N_219,N_323);
and U4955 (N_4955,N_1611,N_466);
xor U4956 (N_4956,N_883,N_389);
nor U4957 (N_4957,N_1780,N_400);
or U4958 (N_4958,N_2469,N_2373);
or U4959 (N_4959,N_1434,N_984);
and U4960 (N_4960,N_2137,N_23);
xnor U4961 (N_4961,N_386,N_906);
nand U4962 (N_4962,N_37,N_75);
xor U4963 (N_4963,N_2141,N_267);
or U4964 (N_4964,N_1337,N_617);
and U4965 (N_4965,N_1615,N_192);
or U4966 (N_4966,N_1464,N_947);
nor U4967 (N_4967,N_1222,N_116);
nand U4968 (N_4968,N_1675,N_1245);
nand U4969 (N_4969,N_1623,N_1779);
nor U4970 (N_4970,N_1654,N_1371);
nor U4971 (N_4971,N_1348,N_2175);
or U4972 (N_4972,N_706,N_2183);
nor U4973 (N_4973,N_1519,N_2188);
or U4974 (N_4974,N_1856,N_1811);
nand U4975 (N_4975,N_599,N_13);
nor U4976 (N_4976,N_1308,N_1998);
nand U4977 (N_4977,N_1732,N_1998);
xor U4978 (N_4978,N_1816,N_1897);
and U4979 (N_4979,N_430,N_2388);
or U4980 (N_4980,N_2162,N_906);
and U4981 (N_4981,N_317,N_817);
and U4982 (N_4982,N_1847,N_436);
and U4983 (N_4983,N_931,N_2288);
and U4984 (N_4984,N_2166,N_406);
xor U4985 (N_4985,N_601,N_1663);
and U4986 (N_4986,N_941,N_1393);
nor U4987 (N_4987,N_576,N_281);
nand U4988 (N_4988,N_2303,N_80);
and U4989 (N_4989,N_1961,N_2203);
and U4990 (N_4990,N_693,N_49);
or U4991 (N_4991,N_1311,N_178);
or U4992 (N_4992,N_2466,N_1234);
nand U4993 (N_4993,N_1982,N_256);
or U4994 (N_4994,N_599,N_919);
nand U4995 (N_4995,N_236,N_36);
nor U4996 (N_4996,N_1510,N_1853);
and U4997 (N_4997,N_616,N_2139);
nor U4998 (N_4998,N_411,N_420);
or U4999 (N_4999,N_1066,N_2167);
and U5000 (N_5000,N_3132,N_3719);
nor U5001 (N_5001,N_4019,N_3105);
or U5002 (N_5002,N_4403,N_3302);
nor U5003 (N_5003,N_3768,N_2914);
nor U5004 (N_5004,N_4379,N_4923);
nand U5005 (N_5005,N_4995,N_4469);
nand U5006 (N_5006,N_4078,N_3597);
nand U5007 (N_5007,N_3200,N_3339);
nor U5008 (N_5008,N_3535,N_2823);
nand U5009 (N_5009,N_4641,N_4620);
nand U5010 (N_5010,N_4960,N_2655);
and U5011 (N_5011,N_2532,N_3253);
nor U5012 (N_5012,N_2929,N_3359);
nor U5013 (N_5013,N_3179,N_2697);
nor U5014 (N_5014,N_4030,N_3990);
nor U5015 (N_5015,N_3757,N_4767);
and U5016 (N_5016,N_3075,N_2972);
nor U5017 (N_5017,N_2692,N_4291);
or U5018 (N_5018,N_3497,N_3322);
and U5019 (N_5019,N_3084,N_4413);
nor U5020 (N_5020,N_3934,N_3584);
nand U5021 (N_5021,N_3961,N_2676);
or U5022 (N_5022,N_2699,N_3162);
nand U5023 (N_5023,N_3493,N_4417);
nor U5024 (N_5024,N_3430,N_2940);
or U5025 (N_5025,N_2641,N_4587);
xnor U5026 (N_5026,N_3752,N_2746);
nand U5027 (N_5027,N_4332,N_3031);
and U5028 (N_5028,N_2984,N_3405);
or U5029 (N_5029,N_2985,N_4146);
and U5030 (N_5030,N_3946,N_2616);
or U5031 (N_5031,N_2881,N_4730);
or U5032 (N_5032,N_4026,N_4474);
or U5033 (N_5033,N_4476,N_3996);
or U5034 (N_5034,N_4732,N_3107);
xnor U5035 (N_5035,N_3674,N_3228);
or U5036 (N_5036,N_4447,N_3547);
xor U5037 (N_5037,N_2729,N_2853);
nor U5038 (N_5038,N_3877,N_4201);
nor U5039 (N_5039,N_3008,N_3890);
nand U5040 (N_5040,N_2667,N_2948);
nor U5041 (N_5041,N_3263,N_3551);
nand U5042 (N_5042,N_2975,N_2609);
xor U5043 (N_5043,N_3303,N_2836);
nand U5044 (N_5044,N_3541,N_4288);
nor U5045 (N_5045,N_2950,N_2679);
nor U5046 (N_5046,N_4583,N_3879);
or U5047 (N_5047,N_3619,N_4986);
and U5048 (N_5048,N_4346,N_3478);
nand U5049 (N_5049,N_4451,N_3867);
or U5050 (N_5050,N_4126,N_4112);
nand U5051 (N_5051,N_3842,N_2748);
xor U5052 (N_5052,N_3203,N_3400);
and U5053 (N_5053,N_3706,N_3317);
xnor U5054 (N_5054,N_4245,N_2727);
or U5055 (N_5055,N_3505,N_4860);
nand U5056 (N_5056,N_2612,N_2859);
or U5057 (N_5057,N_3533,N_4193);
or U5058 (N_5058,N_4044,N_4788);
or U5059 (N_5059,N_4557,N_3281);
or U5060 (N_5060,N_2968,N_3503);
or U5061 (N_5061,N_4998,N_3506);
nor U5062 (N_5062,N_3720,N_2856);
or U5063 (N_5063,N_2526,N_2514);
xor U5064 (N_5064,N_2625,N_3110);
or U5065 (N_5065,N_4881,N_2730);
nand U5066 (N_5066,N_2931,N_2787);
nor U5067 (N_5067,N_4434,N_4615);
xnor U5068 (N_5068,N_3894,N_2894);
or U5069 (N_5069,N_2804,N_3728);
and U5070 (N_5070,N_3680,N_3734);
and U5071 (N_5071,N_3169,N_3664);
or U5072 (N_5072,N_3417,N_4950);
or U5073 (N_5073,N_3868,N_3518);
or U5074 (N_5074,N_3237,N_4808);
nand U5075 (N_5075,N_4852,N_2918);
and U5076 (N_5076,N_3278,N_4856);
and U5077 (N_5077,N_4264,N_3294);
nand U5078 (N_5078,N_4436,N_4147);
or U5079 (N_5079,N_3920,N_2789);
or U5080 (N_5080,N_2848,N_2539);
and U5081 (N_5081,N_3001,N_3765);
xnor U5082 (N_5082,N_4760,N_4188);
nor U5083 (N_5083,N_4187,N_4070);
nand U5084 (N_5084,N_3896,N_4214);
xor U5085 (N_5085,N_2769,N_4952);
or U5086 (N_5086,N_4034,N_4603);
nand U5087 (N_5087,N_3861,N_4235);
nand U5088 (N_5088,N_4203,N_3870);
nor U5089 (N_5089,N_4978,N_3436);
and U5090 (N_5090,N_3191,N_4638);
or U5091 (N_5091,N_3611,N_3862);
nor U5092 (N_5092,N_2973,N_4783);
nor U5093 (N_5093,N_3225,N_3065);
nor U5094 (N_5094,N_4505,N_4576);
nor U5095 (N_5095,N_3211,N_2688);
and U5096 (N_5096,N_2902,N_3422);
nor U5097 (N_5097,N_3045,N_3349);
nor U5098 (N_5098,N_3609,N_2621);
nand U5099 (N_5099,N_3058,N_3499);
or U5100 (N_5100,N_3793,N_2610);
or U5101 (N_5101,N_2669,N_4478);
nand U5102 (N_5102,N_4239,N_3018);
nand U5103 (N_5103,N_3968,N_3631);
nand U5104 (N_5104,N_2772,N_4920);
nor U5105 (N_5105,N_4406,N_4786);
or U5106 (N_5106,N_3052,N_2543);
and U5107 (N_5107,N_4739,N_4254);
nor U5108 (N_5108,N_3285,N_3764);
nor U5109 (N_5109,N_4903,N_3994);
xor U5110 (N_5110,N_4566,N_4278);
and U5111 (N_5111,N_3628,N_2978);
nor U5112 (N_5112,N_2648,N_3908);
and U5113 (N_5113,N_3563,N_3012);
xnor U5114 (N_5114,N_3826,N_4316);
nor U5115 (N_5115,N_3883,N_3427);
nor U5116 (N_5116,N_4409,N_2980);
nor U5117 (N_5117,N_4580,N_4608);
or U5118 (N_5118,N_4516,N_4547);
and U5119 (N_5119,N_2599,N_4311);
xnor U5120 (N_5120,N_3672,N_3582);
and U5121 (N_5121,N_2888,N_3139);
and U5122 (N_5122,N_4368,N_2777);
or U5123 (N_5123,N_4969,N_4072);
nand U5124 (N_5124,N_4851,N_3942);
nand U5125 (N_5125,N_3027,N_3447);
and U5126 (N_5126,N_2759,N_3135);
or U5127 (N_5127,N_2969,N_4339);
nand U5128 (N_5128,N_2687,N_4232);
nor U5129 (N_5129,N_4449,N_2762);
nand U5130 (N_5130,N_4705,N_3494);
xnor U5131 (N_5131,N_3472,N_2521);
and U5132 (N_5132,N_4675,N_4817);
nor U5133 (N_5133,N_2831,N_2845);
and U5134 (N_5134,N_3025,N_4305);
or U5135 (N_5135,N_4828,N_3217);
or U5136 (N_5136,N_3823,N_2611);
or U5137 (N_5137,N_4604,N_2710);
and U5138 (N_5138,N_4962,N_3014);
or U5139 (N_5139,N_4586,N_4521);
nor U5140 (N_5140,N_4052,N_3694);
nand U5141 (N_5141,N_2878,N_3475);
nand U5142 (N_5142,N_2910,N_2898);
or U5143 (N_5143,N_3779,N_3820);
nand U5144 (N_5144,N_3227,N_3519);
and U5145 (N_5145,N_4518,N_3893);
or U5146 (N_5146,N_4156,N_4884);
or U5147 (N_5147,N_3881,N_2749);
nor U5148 (N_5148,N_3548,N_4691);
and U5149 (N_5149,N_2562,N_4205);
or U5150 (N_5150,N_3553,N_2587);
nand U5151 (N_5151,N_3755,N_4749);
or U5152 (N_5152,N_4191,N_3435);
nand U5153 (N_5153,N_3980,N_3164);
nand U5154 (N_5154,N_4271,N_4227);
and U5155 (N_5155,N_4257,N_4894);
nand U5156 (N_5156,N_4999,N_2722);
nand U5157 (N_5157,N_4829,N_4504);
nand U5158 (N_5158,N_2880,N_2889);
or U5159 (N_5159,N_3639,N_3749);
or U5160 (N_5160,N_4161,N_3232);
or U5161 (N_5161,N_3288,N_4766);
or U5162 (N_5162,N_3386,N_4513);
nor U5163 (N_5163,N_2788,N_4865);
xnor U5164 (N_5164,N_3158,N_2714);
nor U5165 (N_5165,N_3011,N_3956);
nand U5166 (N_5166,N_3299,N_4342);
xor U5167 (N_5167,N_3072,N_4177);
nor U5168 (N_5168,N_4882,N_3258);
nor U5169 (N_5169,N_3246,N_4990);
xor U5170 (N_5170,N_4333,N_3212);
nor U5171 (N_5171,N_2650,N_2752);
or U5172 (N_5172,N_3688,N_2732);
or U5173 (N_5173,N_4519,N_4728);
or U5174 (N_5174,N_4563,N_2583);
nor U5175 (N_5175,N_3292,N_2840);
nand U5176 (N_5176,N_4821,N_3856);
nor U5177 (N_5177,N_4128,N_2541);
nand U5178 (N_5178,N_3420,N_4934);
or U5179 (N_5179,N_3906,N_4165);
nor U5180 (N_5180,N_3751,N_3635);
nor U5181 (N_5181,N_3666,N_4537);
nand U5182 (N_5182,N_4209,N_3204);
or U5183 (N_5183,N_3426,N_2593);
xor U5184 (N_5184,N_4080,N_4462);
nand U5185 (N_5185,N_2837,N_3959);
and U5186 (N_5186,N_3773,N_4336);
or U5187 (N_5187,N_3971,N_2753);
nand U5188 (N_5188,N_2673,N_2670);
xor U5189 (N_5189,N_3131,N_4769);
or U5190 (N_5190,N_4867,N_4699);
nor U5191 (N_5191,N_2799,N_3248);
nor U5192 (N_5192,N_4507,N_4915);
and U5193 (N_5193,N_4415,N_3707);
nand U5194 (N_5194,N_2865,N_4768);
or U5195 (N_5195,N_3822,N_3182);
nor U5196 (N_5196,N_4763,N_2807);
and U5197 (N_5197,N_2510,N_4051);
nand U5198 (N_5198,N_3526,N_3767);
xnor U5199 (N_5199,N_3352,N_4972);
and U5200 (N_5200,N_4129,N_3161);
xnor U5201 (N_5201,N_3723,N_4400);
nand U5202 (N_5202,N_4989,N_2668);
nor U5203 (N_5203,N_4579,N_3256);
nor U5204 (N_5204,N_4470,N_2996);
nand U5205 (N_5205,N_2717,N_4125);
or U5206 (N_5206,N_4012,N_3252);
nor U5207 (N_5207,N_4858,N_4480);
nor U5208 (N_5208,N_4384,N_2890);
nand U5209 (N_5209,N_2505,N_4377);
and U5210 (N_5210,N_3652,N_3944);
and U5211 (N_5211,N_4646,N_3766);
and U5212 (N_5212,N_2995,N_3301);
nand U5213 (N_5213,N_4197,N_4155);
nor U5214 (N_5214,N_4086,N_4779);
nand U5215 (N_5215,N_2813,N_3198);
or U5216 (N_5216,N_3009,N_4486);
or U5217 (N_5217,N_3163,N_4911);
or U5218 (N_5218,N_3486,N_4243);
nand U5219 (N_5219,N_4676,N_4991);
or U5220 (N_5220,N_3513,N_2545);
nand U5221 (N_5221,N_2857,N_2872);
and U5222 (N_5222,N_2594,N_3995);
xor U5223 (N_5223,N_3119,N_3904);
nand U5224 (N_5224,N_4532,N_3583);
nand U5225 (N_5225,N_2842,N_4785);
or U5226 (N_5226,N_3991,N_3887);
or U5227 (N_5227,N_4724,N_3095);
nor U5228 (N_5228,N_3341,N_3943);
and U5229 (N_5229,N_3905,N_4929);
or U5230 (N_5230,N_2988,N_3026);
nor U5231 (N_5231,N_4900,N_3094);
nor U5232 (N_5232,N_3627,N_3891);
nand U5233 (N_5233,N_4906,N_3446);
nand U5234 (N_5234,N_3230,N_3098);
or U5235 (N_5235,N_4976,N_4636);
nand U5236 (N_5236,N_4250,N_3771);
nand U5237 (N_5237,N_4649,N_3721);
or U5238 (N_5238,N_3869,N_3196);
and U5239 (N_5239,N_3595,N_3633);
xor U5240 (N_5240,N_4226,N_2815);
nand U5241 (N_5241,N_4747,N_2660);
and U5242 (N_5242,N_4647,N_2803);
nand U5243 (N_5243,N_4565,N_4622);
xor U5244 (N_5244,N_3006,N_3214);
or U5245 (N_5245,N_4120,N_4048);
nand U5246 (N_5246,N_3327,N_4115);
and U5247 (N_5247,N_3395,N_3019);
xnor U5248 (N_5248,N_3849,N_4375);
nor U5249 (N_5249,N_4922,N_4351);
and U5250 (N_5250,N_4325,N_4266);
or U5251 (N_5251,N_4787,N_3261);
and U5252 (N_5252,N_4025,N_2512);
nor U5253 (N_5253,N_4558,N_3712);
nor U5254 (N_5254,N_2633,N_2951);
nor U5255 (N_5255,N_3251,N_2838);
or U5256 (N_5256,N_4401,N_4733);
nand U5257 (N_5257,N_2513,N_2809);
xnor U5258 (N_5258,N_2690,N_3283);
xnor U5259 (N_5259,N_3264,N_3986);
or U5260 (N_5260,N_2570,N_2953);
or U5261 (N_5261,N_2944,N_4632);
nand U5262 (N_5262,N_3282,N_4694);
nor U5263 (N_5263,N_3554,N_4634);
or U5264 (N_5264,N_3013,N_4249);
nor U5265 (N_5265,N_3832,N_3142);
or U5266 (N_5266,N_3268,N_4941);
nand U5267 (N_5267,N_4596,N_4875);
nor U5268 (N_5268,N_3035,N_3007);
xnor U5269 (N_5269,N_4574,N_4643);
or U5270 (N_5270,N_4578,N_4600);
nand U5271 (N_5271,N_4772,N_3489);
nor U5272 (N_5272,N_2764,N_3310);
nor U5273 (N_5273,N_3096,N_2963);
or U5274 (N_5274,N_3235,N_2586);
and U5275 (N_5275,N_4588,N_4623);
and U5276 (N_5276,N_3314,N_3402);
nand U5277 (N_5277,N_4689,N_4715);
nor U5278 (N_5278,N_4742,N_3809);
nor U5279 (N_5279,N_4425,N_3088);
nand U5280 (N_5280,N_2602,N_4195);
and U5281 (N_5281,N_4844,N_3209);
nand U5282 (N_5282,N_2938,N_4688);
nand U5283 (N_5283,N_4198,N_4223);
nand U5284 (N_5284,N_3411,N_4420);
nor U5285 (N_5285,N_4392,N_4711);
and U5286 (N_5286,N_2579,N_4130);
nor U5287 (N_5287,N_3234,N_2866);
nand U5288 (N_5288,N_4697,N_4422);
xor U5289 (N_5289,N_4360,N_4473);
nor U5290 (N_5290,N_2644,N_3592);
nand U5291 (N_5291,N_3074,N_3950);
and U5292 (N_5292,N_2983,N_2850);
and U5293 (N_5293,N_3882,N_3482);
or U5294 (N_5294,N_3120,N_2954);
nand U5295 (N_5295,N_4764,N_4897);
and U5296 (N_5296,N_4179,N_2805);
and U5297 (N_5297,N_3484,N_4369);
or U5298 (N_5298,N_4550,N_4317);
nor U5299 (N_5299,N_4877,N_4221);
nand U5300 (N_5300,N_4166,N_4135);
nor U5301 (N_5301,N_4217,N_2955);
and U5302 (N_5302,N_3743,N_2582);
and U5303 (N_5303,N_3469,N_4095);
or U5304 (N_5304,N_3407,N_4762);
or U5305 (N_5305,N_4277,N_4815);
and U5306 (N_5306,N_4544,N_3922);
and U5307 (N_5307,N_4714,N_3201);
or U5308 (N_5308,N_3442,N_2999);
and U5309 (N_5309,N_3824,N_3585);
and U5310 (N_5310,N_4863,N_3173);
or U5311 (N_5311,N_4483,N_4612);
and U5312 (N_5312,N_4741,N_4490);
nor U5313 (N_5313,N_4531,N_4402);
nand U5314 (N_5314,N_3085,N_3912);
nor U5315 (N_5315,N_4846,N_2656);
and U5316 (N_5316,N_4506,N_3509);
or U5317 (N_5317,N_2675,N_2811);
or U5318 (N_5318,N_2645,N_4987);
xor U5319 (N_5319,N_4255,N_4873);
nor U5320 (N_5320,N_4562,N_2504);
nor U5321 (N_5321,N_4966,N_3586);
or U5322 (N_5322,N_2715,N_4488);
or U5323 (N_5323,N_4984,N_4716);
nor U5324 (N_5324,N_2870,N_3607);
nand U5325 (N_5325,N_3988,N_2651);
and U5326 (N_5326,N_4114,N_4211);
and U5327 (N_5327,N_3865,N_3969);
nand U5328 (N_5328,N_3960,N_3276);
nor U5329 (N_5329,N_2998,N_4753);
and U5330 (N_5330,N_2916,N_2515);
or U5331 (N_5331,N_2793,N_4213);
and U5332 (N_5332,N_3337,N_3587);
and U5333 (N_5333,N_3514,N_3938);
nand U5334 (N_5334,N_3655,N_3542);
nand U5335 (N_5335,N_3703,N_3559);
nor U5336 (N_5336,N_3815,N_4816);
nand U5337 (N_5337,N_3747,N_3853);
nand U5338 (N_5338,N_4605,N_4833);
and U5339 (N_5339,N_3731,N_4681);
nor U5340 (N_5340,N_3092,N_2604);
or U5341 (N_5341,N_4938,N_3250);
xor U5342 (N_5342,N_2751,N_3661);
nor U5343 (N_5343,N_4848,N_4445);
and U5344 (N_5344,N_2824,N_3847);
or U5345 (N_5345,N_2832,N_3955);
or U5346 (N_5346,N_2643,N_3255);
nand U5347 (N_5347,N_4010,N_2623);
xor U5348 (N_5348,N_4594,N_4614);
xor U5349 (N_5349,N_4940,N_3056);
or U5350 (N_5350,N_3852,N_4079);
or U5351 (N_5351,N_2994,N_4859);
or U5352 (N_5352,N_3388,N_2942);
and U5353 (N_5353,N_4349,N_4994);
nand U5354 (N_5354,N_3070,N_2816);
nor U5355 (N_5355,N_3277,N_2993);
nor U5356 (N_5356,N_2663,N_4082);
nor U5357 (N_5357,N_3623,N_4357);
nor U5358 (N_5358,N_3023,N_3677);
and U5359 (N_5359,N_4642,N_2775);
nor U5360 (N_5360,N_2786,N_3077);
nand U5361 (N_5361,N_3599,N_2529);
or U5362 (N_5362,N_2970,N_3698);
nand U5363 (N_5363,N_3210,N_4465);
nor U5364 (N_5364,N_3468,N_3321);
or U5365 (N_5365,N_2626,N_4348);
or U5366 (N_5366,N_3638,N_2581);
and U5367 (N_5367,N_4713,N_4301);
and U5368 (N_5368,N_3498,N_3774);
or U5369 (N_5369,N_4467,N_4055);
nand U5370 (N_5370,N_2891,N_2884);
nand U5371 (N_5371,N_2720,N_3297);
nor U5372 (N_5372,N_3454,N_4395);
or U5373 (N_5373,N_3632,N_2770);
and U5374 (N_5374,N_4610,N_4459);
or U5375 (N_5375,N_2672,N_3236);
xnor U5376 (N_5376,N_2658,N_4098);
nor U5377 (N_5377,N_4570,N_4811);
and U5378 (N_5378,N_3540,N_3108);
or U5379 (N_5379,N_4870,N_2897);
nand U5380 (N_5380,N_3644,N_2851);
or U5381 (N_5381,N_4207,N_2964);
xor U5382 (N_5382,N_2934,N_4660);
nor U5383 (N_5383,N_4031,N_4390);
nor U5384 (N_5384,N_4123,N_2588);
nor U5385 (N_5385,N_4542,N_3183);
nor U5386 (N_5386,N_3239,N_3187);
and U5387 (N_5387,N_2737,N_4463);
and U5388 (N_5388,N_4439,N_3517);
or U5389 (N_5389,N_4977,N_4391);
or U5390 (N_5390,N_4892,N_2558);
xnor U5391 (N_5391,N_3280,N_4290);
and U5392 (N_5392,N_2522,N_3385);
nand U5393 (N_5393,N_4294,N_4830);
nand U5394 (N_5394,N_3115,N_3176);
and U5395 (N_5395,N_4874,N_4359);
and U5396 (N_5396,N_3936,N_3848);
and U5397 (N_5397,N_3409,N_3434);
nor U5398 (N_5398,N_4560,N_2517);
or U5399 (N_5399,N_3821,N_3641);
nand U5400 (N_5400,N_4789,N_3401);
nand U5401 (N_5401,N_3345,N_3932);
and U5402 (N_5402,N_4347,N_3002);
nand U5403 (N_5403,N_3704,N_2571);
or U5404 (N_5404,N_3662,N_3103);
nor U5405 (N_5405,N_4602,N_4891);
nand U5406 (N_5406,N_2719,N_2523);
and U5407 (N_5407,N_4139,N_2949);
nand U5408 (N_5408,N_4868,N_4210);
or U5409 (N_5409,N_4598,N_4016);
nor U5410 (N_5410,N_2511,N_3081);
or U5411 (N_5411,N_3152,N_3937);
nand U5412 (N_5412,N_3671,N_3534);
nand U5413 (N_5413,N_4692,N_4393);
or U5414 (N_5414,N_2566,N_4782);
or U5415 (N_5415,N_2576,N_4831);
xor U5416 (N_5416,N_3485,N_3166);
and U5417 (N_5417,N_3202,N_3355);
or U5418 (N_5418,N_4101,N_3978);
nand U5419 (N_5419,N_4708,N_3590);
xor U5420 (N_5420,N_4773,N_2654);
and U5421 (N_5421,N_3690,N_3722);
nand U5422 (N_5422,N_3799,N_3199);
nand U5423 (N_5423,N_3827,N_2637);
nor U5424 (N_5424,N_4280,N_4035);
nand U5425 (N_5425,N_3589,N_4584);
or U5426 (N_5426,N_4710,N_2686);
nand U5427 (N_5427,N_3304,N_4606);
nor U5428 (N_5428,N_4168,N_3213);
and U5429 (N_5429,N_3348,N_4200);
nand U5430 (N_5430,N_2761,N_3384);
and U5431 (N_5431,N_4430,N_4062);
or U5432 (N_5432,N_3884,N_4836);
or U5433 (N_5433,N_4312,N_3039);
or U5434 (N_5434,N_2618,N_2551);
or U5435 (N_5435,N_3149,N_3814);
xnor U5436 (N_5436,N_3983,N_2783);
or U5437 (N_5437,N_2774,N_3404);
and U5438 (N_5438,N_2731,N_4320);
or U5439 (N_5439,N_3354,N_4354);
nor U5440 (N_5440,N_3886,N_4526);
xor U5441 (N_5441,N_3818,N_4066);
nor U5442 (N_5442,N_4380,N_4286);
xnor U5443 (N_5443,N_3568,N_3508);
nand U5444 (N_5444,N_4279,N_4282);
xor U5445 (N_5445,N_3458,N_4388);
and U5446 (N_5446,N_4119,N_4485);
and U5447 (N_5447,N_3496,N_3933);
nand U5448 (N_5448,N_3606,N_4064);
and U5449 (N_5449,N_4927,N_3759);
nor U5450 (N_5450,N_4803,N_2671);
and U5451 (N_5451,N_4672,N_4458);
and U5452 (N_5452,N_3715,N_3783);
nor U5453 (N_5453,N_4242,N_3642);
or U5454 (N_5454,N_3305,N_3374);
or U5455 (N_5455,N_3835,N_3566);
or U5456 (N_5456,N_3421,N_4840);
and U5457 (N_5457,N_3829,N_4635);
xor U5458 (N_5458,N_3876,N_4158);
nand U5459 (N_5459,N_2653,N_4790);
nand U5460 (N_5460,N_2711,N_4667);
nand U5461 (N_5461,N_3086,N_3803);
nor U5462 (N_5462,N_3254,N_4032);
or U5463 (N_5463,N_3308,N_2546);
nor U5464 (N_5464,N_3265,N_3373);
nor U5465 (N_5465,N_2858,N_3155);
nand U5466 (N_5466,N_2875,N_3190);
xnor U5467 (N_5467,N_3802,N_3948);
or U5468 (N_5468,N_4387,N_3432);
or U5469 (N_5469,N_4720,N_4942);
nand U5470 (N_5470,N_4398,N_3732);
nor U5471 (N_5471,N_2613,N_4795);
xor U5472 (N_5472,N_4225,N_3444);
and U5473 (N_5473,N_3247,N_3653);
xnor U5474 (N_5474,N_4104,N_2615);
or U5475 (N_5475,N_3490,N_3624);
xor U5476 (N_5476,N_4341,N_4755);
nand U5477 (N_5477,N_2819,N_3350);
xnor U5478 (N_5478,N_4424,N_4778);
or U5479 (N_5479,N_2661,N_4650);
nor U5480 (N_5480,N_4818,N_2818);
nor U5481 (N_5481,N_2795,N_4440);
nand U5482 (N_5482,N_4745,N_3329);
nor U5483 (N_5483,N_3062,N_3394);
or U5484 (N_5484,N_4524,N_3923);
or U5485 (N_5485,N_4813,N_4930);
nor U5486 (N_5486,N_3917,N_4110);
nand U5487 (N_5487,N_3387,N_2605);
and U5488 (N_5488,N_4220,N_2622);
xor U5489 (N_5489,N_3622,N_4985);
nand U5490 (N_5490,N_4050,N_4238);
or U5491 (N_5491,N_4613,N_4535);
nor U5492 (N_5492,N_2619,N_4366);
and U5493 (N_5493,N_3392,N_2703);
nor U5494 (N_5494,N_4310,N_4298);
or U5495 (N_5495,N_2724,N_4085);
nand U5496 (N_5496,N_3379,N_3973);
or U5497 (N_5497,N_3501,N_2598);
xnor U5498 (N_5498,N_2627,N_4798);
xor U5499 (N_5499,N_4276,N_3681);
or U5500 (N_5500,N_3796,N_3574);
or U5501 (N_5501,N_4408,N_4269);
nor U5502 (N_5502,N_3043,N_4965);
and U5503 (N_5503,N_4639,N_4807);
and U5504 (N_5504,N_4182,N_3361);
nand U5505 (N_5505,N_2728,N_2886);
nor U5506 (N_5506,N_4740,N_4842);
or U5507 (N_5507,N_4907,N_4945);
nand U5508 (N_5508,N_3748,N_3910);
nand U5509 (N_5509,N_3479,N_2561);
or U5510 (N_5510,N_4407,N_3193);
nor U5511 (N_5511,N_4796,N_2548);
and U5512 (N_5512,N_4528,N_4530);
and U5513 (N_5513,N_2763,N_2747);
or U5514 (N_5514,N_4003,N_2524);
or U5515 (N_5515,N_3874,N_4108);
nand U5516 (N_5516,N_2509,N_2585);
xor U5517 (N_5517,N_2830,N_3491);
nor U5518 (N_5518,N_3224,N_3289);
xnor U5519 (N_5519,N_2885,N_3965);
and U5520 (N_5520,N_2961,N_3760);
and U5521 (N_5521,N_3682,N_3323);
or U5522 (N_5522,N_3958,N_3104);
nor U5523 (N_5523,N_2806,N_3602);
and U5524 (N_5524,N_3356,N_3197);
nand U5525 (N_5525,N_4047,N_4967);
xor U5526 (N_5526,N_4835,N_4373);
nand U5527 (N_5527,N_3985,N_4864);
nand U5528 (N_5528,N_3925,N_2962);
xnor U5529 (N_5529,N_4411,N_4054);
nand U5530 (N_5530,N_3903,N_4499);
and U5531 (N_5531,N_4702,N_3596);
and U5532 (N_5532,N_3073,N_3834);
nor U5533 (N_5533,N_3730,N_3577);
nor U5534 (N_5534,N_4394,N_2528);
and U5535 (N_5535,N_4997,N_3015);
xnor U5536 (N_5536,N_3679,N_4138);
xor U5537 (N_5537,N_4781,N_2740);
or U5538 (N_5538,N_3579,N_2925);
or U5539 (N_5539,N_4855,N_3691);
or U5540 (N_5540,N_4185,N_2826);
nand U5541 (N_5541,N_4230,N_2614);
nand U5542 (N_5542,N_4673,N_3038);
nand U5543 (N_5543,N_2642,N_3555);
or U5544 (N_5544,N_3911,N_4124);
or U5545 (N_5545,N_3931,N_3398);
or U5546 (N_5546,N_3940,N_4825);
xnor U5547 (N_5547,N_3030,N_3046);
nor U5548 (N_5548,N_4533,N_3953);
nor U5549 (N_5549,N_3029,N_3414);
nor U5550 (N_5550,N_3741,N_3137);
nand U5551 (N_5551,N_4498,N_2628);
nand U5552 (N_5552,N_3445,N_4696);
nand U5553 (N_5553,N_4592,N_3460);
nor U5554 (N_5554,N_2674,N_4553);
and U5555 (N_5555,N_3331,N_3569);
and U5556 (N_5556,N_4759,N_4539);
nand U5557 (N_5557,N_3249,N_4902);
and U5558 (N_5558,N_4106,N_4805);
xnor U5559 (N_5559,N_3470,N_4495);
or U5560 (N_5560,N_3047,N_3892);
and U5561 (N_5561,N_4068,N_3116);
or U5562 (N_5562,N_4917,N_3811);
nand U5563 (N_5563,N_2506,N_4208);
or U5564 (N_5564,N_3243,N_3524);
nor U5565 (N_5565,N_3003,N_4640);
or U5566 (N_5566,N_4037,N_3516);
nor U5567 (N_5567,N_2895,N_3369);
nand U5568 (N_5568,N_3974,N_4418);
and U5569 (N_5569,N_4352,N_3957);
nor U5570 (N_5570,N_3122,N_4827);
nand U5571 (N_5571,N_2755,N_4703);
nand U5572 (N_5572,N_2846,N_3069);
xnor U5573 (N_5573,N_3219,N_4511);
and U5574 (N_5574,N_2577,N_4683);
nand U5575 (N_5575,N_3713,N_2708);
nor U5576 (N_5576,N_3878,N_3502);
nor U5577 (N_5577,N_3567,N_3620);
nor U5578 (N_5578,N_4042,N_4625);
or U5579 (N_5579,N_4204,N_4655);
and U5580 (N_5580,N_3068,N_2952);
nor U5581 (N_5581,N_2765,N_2976);
nand U5582 (N_5582,N_4585,N_4656);
xnor U5583 (N_5583,N_3476,N_3593);
or U5584 (N_5584,N_4162,N_4089);
xor U5585 (N_5585,N_3186,N_3451);
xnor U5586 (N_5586,N_4087,N_3082);
and U5587 (N_5587,N_2796,N_4717);
nand U5588 (N_5588,N_2828,N_3330);
and U5589 (N_5589,N_3165,N_4121);
xnor U5590 (N_5590,N_4231,N_3223);
or U5591 (N_5591,N_4284,N_3604);
and U5592 (N_5592,N_4063,N_4572);
and U5593 (N_5593,N_3787,N_3954);
nor U5594 (N_5594,N_3184,N_4918);
xor U5595 (N_5595,N_3406,N_4627);
or U5596 (N_5596,N_3170,N_4241);
nand U5597 (N_5597,N_3456,N_2896);
nand U5598 (N_5598,N_3761,N_2966);
nor U5599 (N_5599,N_4222,N_3206);
or U5600 (N_5600,N_3702,N_3871);
nor U5601 (N_5601,N_4429,N_3054);
and U5602 (N_5602,N_3670,N_4300);
nor U5603 (N_5603,N_3836,N_4581);
nand U5604 (N_5604,N_4094,N_3306);
and U5605 (N_5605,N_3143,N_4259);
nor U5606 (N_5606,N_4015,N_3840);
nor U5607 (N_5607,N_3174,N_3067);
nor U5608 (N_5608,N_4194,N_2901);
nand U5609 (N_5609,N_4275,N_3238);
or U5610 (N_5610,N_3845,N_3807);
nor U5611 (N_5611,N_2591,N_4883);
and U5612 (N_5612,N_4319,N_2790);
nor U5613 (N_5613,N_3262,N_4652);
nand U5614 (N_5614,N_4854,N_3780);
and U5615 (N_5615,N_2735,N_3488);
xnor U5616 (N_5616,N_3172,N_4904);
nor U5617 (N_5617,N_4889,N_4431);
or U5618 (N_5618,N_3838,N_2817);
xor U5619 (N_5619,N_4843,N_2695);
nand U5620 (N_5620,N_3382,N_3320);
or U5621 (N_5621,N_3271,N_2572);
nand U5622 (N_5622,N_3977,N_2563);
or U5623 (N_5623,N_4886,N_3381);
nand U5624 (N_5624,N_2920,N_4734);
xor U5625 (N_5625,N_4039,N_4099);
xnor U5626 (N_5626,N_3902,N_2767);
nor U5627 (N_5627,N_4564,N_3726);
xnor U5628 (N_5628,N_4822,N_3326);
and U5629 (N_5629,N_3557,N_4545);
and U5630 (N_5630,N_4979,N_3561);
nor U5631 (N_5631,N_3036,N_4957);
or U5632 (N_5632,N_4693,N_2726);
xor U5633 (N_5633,N_4364,N_3195);
or U5634 (N_5634,N_4329,N_3159);
and U5635 (N_5635,N_2990,N_2527);
nand U5636 (N_5636,N_4363,N_3909);
and U5637 (N_5637,N_4331,N_2704);
nand U5638 (N_5638,N_4053,N_2629);
or U5639 (N_5639,N_4736,N_3428);
nor U5640 (N_5640,N_4433,N_2538);
nor U5641 (N_5641,N_4471,N_3080);
nand U5642 (N_5642,N_3781,N_3689);
xor U5643 (N_5643,N_2589,N_2863);
or U5644 (N_5644,N_4142,N_4296);
nand U5645 (N_5645,N_2941,N_4664);
nor U5646 (N_5646,N_4944,N_3270);
nand U5647 (N_5647,N_4421,N_2712);
or U5648 (N_5648,N_4926,N_3778);
and U5649 (N_5649,N_2833,N_2649);
or U5650 (N_5650,N_4880,N_2684);
nor U5651 (N_5651,N_3309,N_2810);
or U5652 (N_5652,N_4682,N_3466);
nand U5653 (N_5653,N_4928,N_4554);
or U5654 (N_5654,N_4706,N_4396);
and U5655 (N_5655,N_4905,N_4236);
or U5656 (N_5656,N_2792,N_3578);
nand U5657 (N_5657,N_2659,N_4726);
nand U5658 (N_5658,N_3443,N_3530);
nand U5659 (N_5659,N_3613,N_4097);
nor U5660 (N_5660,N_4160,N_3177);
nor U5661 (N_5661,N_4370,N_4181);
or U5662 (N_5662,N_4921,N_4935);
nor U5663 (N_5663,N_2861,N_3138);
and U5664 (N_5664,N_4725,N_3181);
or U5665 (N_5665,N_4644,N_3913);
nand U5666 (N_5666,N_3857,N_2932);
and U5667 (N_5667,N_4687,N_3123);
nor U5668 (N_5668,N_4630,N_3291);
nor U5669 (N_5669,N_2631,N_3351);
and U5670 (N_5670,N_4774,N_4541);
nor U5671 (N_5671,N_4405,N_3650);
or U5672 (N_5672,N_3570,N_3636);
nor U5673 (N_5673,N_4247,N_3693);
nand U5674 (N_5674,N_4427,N_2689);
or U5675 (N_5675,N_3367,N_3634);
and U5676 (N_5676,N_3797,N_4666);
and U5677 (N_5677,N_4229,N_2555);
nand U5678 (N_5678,N_3375,N_4045);
nor U5679 (N_5679,N_2500,N_4297);
and U5680 (N_5680,N_3510,N_2691);
nor U5681 (N_5681,N_3573,N_2781);
nor U5682 (N_5682,N_3335,N_2797);
or U5683 (N_5683,N_3898,N_4452);
nor U5684 (N_5684,N_3477,N_4503);
nand U5685 (N_5685,N_3915,N_3625);
nand U5686 (N_5686,N_3614,N_2868);
or U5687 (N_5687,N_3873,N_4939);
nand U5688 (N_5688,N_4216,N_3926);
nand U5689 (N_5689,N_3939,N_4913);
and U5690 (N_5690,N_3572,N_4001);
or U5691 (N_5691,N_3378,N_3128);
nand U5692 (N_5692,N_4381,N_3129);
and U5693 (N_5693,N_3050,N_4059);
nand U5694 (N_5694,N_4132,N_4060);
nand U5695 (N_5695,N_3810,N_4548);
nand U5696 (N_5696,N_4731,N_3949);
or U5697 (N_5697,N_3880,N_3360);
and U5698 (N_5698,N_3049,N_4154);
or U5699 (N_5699,N_3997,N_3366);
nand U5700 (N_5700,N_3140,N_2776);
or U5701 (N_5701,N_3078,N_3180);
or U5702 (N_5702,N_4727,N_4670);
nor U5703 (N_5703,N_3192,N_4314);
nand U5704 (N_5704,N_4169,N_3629);
and U5705 (N_5705,N_2559,N_4879);
or U5706 (N_5706,N_4024,N_3284);
nand U5707 (N_5707,N_2862,N_2754);
or U5708 (N_5708,N_4441,N_3733);
nor U5709 (N_5709,N_2960,N_4058);
nand U5710 (N_5710,N_4040,N_3032);
nor U5711 (N_5711,N_3118,N_3575);
nand U5712 (N_5712,N_4281,N_3028);
xor U5713 (N_5713,N_2946,N_3817);
nand U5714 (N_5714,N_3692,N_3286);
and U5715 (N_5715,N_3746,N_3380);
or U5716 (N_5716,N_3695,N_4924);
nor U5717 (N_5717,N_4482,N_2578);
nor U5718 (N_5718,N_2893,N_3296);
nand U5719 (N_5719,N_3916,N_2822);
nand U5720 (N_5720,N_3649,N_4721);
nand U5721 (N_5721,N_4794,N_3626);
nand U5722 (N_5722,N_3951,N_4552);
or U5723 (N_5723,N_2820,N_4841);
nand U5724 (N_5724,N_2974,N_4980);
nor U5725 (N_5725,N_2989,N_3124);
xor U5726 (N_5726,N_4515,N_4389);
xnor U5727 (N_5727,N_3389,N_3591);
nand U5728 (N_5728,N_4758,N_3560);
and U5729 (N_5729,N_3318,N_3160);
or U5730 (N_5730,N_3017,N_4192);
xor U5731 (N_5731,N_2943,N_4618);
xor U5732 (N_5732,N_4568,N_3543);
and U5733 (N_5733,N_4164,N_3828);
xor U5734 (N_5734,N_4455,N_4599);
or U5735 (N_5735,N_3207,N_4215);
nor U5736 (N_5736,N_4959,N_4857);
nor U5737 (N_5737,N_4096,N_4750);
nand U5738 (N_5738,N_4908,N_4228);
xor U5739 (N_5739,N_3725,N_3372);
and U5740 (N_5740,N_2516,N_3736);
nand U5741 (N_5741,N_3408,N_3724);
and U5742 (N_5742,N_2997,N_4399);
nand U5743 (N_5743,N_2852,N_4662);
or U5744 (N_5744,N_2982,N_2744);
and U5745 (N_5745,N_3616,N_3257);
nand U5746 (N_5746,N_2912,N_3101);
and U5747 (N_5747,N_2827,N_4307);
or U5748 (N_5748,N_4374,N_4273);
and U5749 (N_5749,N_4362,N_3640);
and U5750 (N_5750,N_4218,N_4358);
nor U5751 (N_5751,N_4869,N_3205);
nor U5752 (N_5752,N_3918,N_3663);
nand U5753 (N_5753,N_4090,N_4679);
and U5754 (N_5754,N_3467,N_4260);
xnor U5755 (N_5755,N_2812,N_3133);
or U5756 (N_5756,N_3071,N_2947);
nand U5757 (N_5757,N_3544,N_3564);
and U5758 (N_5758,N_3549,N_3146);
xnor U5759 (N_5759,N_4137,N_4628);
nand U5760 (N_5760,N_3945,N_2639);
xnor U5761 (N_5761,N_3357,N_2716);
and U5762 (N_5762,N_4102,N_3789);
or U5763 (N_5763,N_4084,N_3063);
or U5764 (N_5764,N_4466,N_4274);
nand U5765 (N_5765,N_3004,N_4046);
xor U5766 (N_5766,N_2844,N_4057);
or U5767 (N_5767,N_4963,N_3928);
xnor U5768 (N_5768,N_2519,N_2738);
nand U5769 (N_5769,N_2718,N_4262);
or U5770 (N_5770,N_4497,N_4536);
nor U5771 (N_5771,N_3964,N_2677);
xnor U5772 (N_5772,N_3492,N_4933);
and U5773 (N_5773,N_4771,N_3410);
or U5774 (N_5774,N_2839,N_3825);
nor U5775 (N_5775,N_3233,N_3455);
nand U5776 (N_5776,N_3929,N_3231);
xor U5777 (N_5777,N_2864,N_3079);
and U5778 (N_5778,N_4122,N_2584);
nor U5779 (N_5779,N_4327,N_2620);
nand U5780 (N_5780,N_3527,N_3097);
and U5781 (N_5781,N_4252,N_3005);
nor U5782 (N_5782,N_4428,N_3109);
nor U5783 (N_5783,N_4792,N_2959);
or U5784 (N_5784,N_2939,N_3112);
and U5785 (N_5785,N_4083,N_2608);
nor U5786 (N_5786,N_4543,N_4776);
or U5787 (N_5787,N_4799,N_3683);
nor U5788 (N_5788,N_4916,N_3999);
or U5789 (N_5789,N_3368,N_3245);
or U5790 (N_5790,N_4258,N_4041);
xnor U5791 (N_5791,N_3076,N_2601);
and U5792 (N_5792,N_4668,N_3437);
nand U5793 (N_5793,N_3851,N_4631);
nor U5794 (N_5794,N_4525,N_3833);
nor U5795 (N_5795,N_4426,N_2508);
nand U5796 (N_5796,N_4328,N_4983);
xor U5797 (N_5797,N_3397,N_3010);
or U5798 (N_5798,N_3798,N_3512);
nor U5799 (N_5799,N_4270,N_4414);
or U5800 (N_5800,N_3711,N_3782);
nor U5801 (N_5801,N_4109,N_3738);
nand U5802 (N_5802,N_2518,N_4233);
xnor U5803 (N_5803,N_4701,N_3795);
xor U5804 (N_5804,N_4157,N_4475);
xor U5805 (N_5805,N_3338,N_4065);
nand U5806 (N_5806,N_4657,N_2557);
xnor U5807 (N_5807,N_3952,N_3393);
nor U5808 (N_5808,N_2829,N_4573);
or U5809 (N_5809,N_3148,N_4951);
and U5810 (N_5810,N_2905,N_4671);
nand U5811 (N_5811,N_2600,N_2678);
nor U5812 (N_5812,N_4509,N_3546);
and U5813 (N_5813,N_4306,N_4819);
and U5814 (N_5814,N_3024,N_2569);
and U5815 (N_5815,N_3739,N_4283);
nor U5816 (N_5816,N_4337,N_4496);
and U5817 (N_5817,N_4791,N_4540);
nor U5818 (N_5818,N_4202,N_3500);
nand U5819 (N_5819,N_4321,N_4416);
nand U5820 (N_5820,N_3433,N_3813);
or U5821 (N_5821,N_4589,N_4492);
nand U5822 (N_5822,N_3189,N_3042);
nand U5823 (N_5823,N_4709,N_4450);
and U5824 (N_5824,N_2936,N_4633);
xnor U5825 (N_5825,N_4948,N_2802);
and U5826 (N_5826,N_3218,N_4253);
and U5827 (N_5827,N_4186,N_2919);
nor U5828 (N_5828,N_4116,N_3066);
nand U5829 (N_5829,N_3665,N_3336);
or U5830 (N_5830,N_3740,N_4595);
nand U5831 (N_5831,N_3850,N_3093);
nand U5832 (N_5832,N_2909,N_4481);
nor U5833 (N_5833,N_4265,N_4383);
xnor U5834 (N_5834,N_4017,N_3675);
or U5835 (N_5835,N_4690,N_3371);
nand U5836 (N_5836,N_4523,N_3935);
or U5837 (N_5837,N_4982,N_3647);
nand U5838 (N_5838,N_3989,N_4559);
and U5839 (N_5839,N_3328,N_3588);
nand U5840 (N_5840,N_3889,N_4315);
and U5841 (N_5841,N_4878,N_3040);
or U5842 (N_5842,N_3895,N_3000);
nand U5843 (N_5843,N_4793,N_3717);
and U5844 (N_5844,N_2883,N_3800);
nand U5845 (N_5845,N_3901,N_4775);
nand U5846 (N_5846,N_3770,N_4159);
or U5847 (N_5847,N_4077,N_3090);
xor U5848 (N_5848,N_2766,N_4567);
or U5849 (N_5849,N_3020,N_4961);
nand U5850 (N_5850,N_4748,N_4973);
nor U5851 (N_5851,N_3875,N_3272);
and U5852 (N_5852,N_3794,N_3696);
or U5853 (N_5853,N_3144,N_2564);
nand U5854 (N_5854,N_4448,N_4853);
nand U5855 (N_5855,N_4111,N_4534);
and U5856 (N_5856,N_3522,N_2554);
xnor U5857 (N_5857,N_4723,N_3907);
nor U5858 (N_5858,N_2542,N_3269);
nor U5859 (N_5859,N_3295,N_3343);
nor U5860 (N_5860,N_3462,N_3843);
or U5861 (N_5861,N_3819,N_3854);
nand U5862 (N_5862,N_4005,N_3053);
or U5863 (N_5863,N_3727,N_4479);
nand U5864 (N_5864,N_3453,N_4183);
or U5865 (N_5865,N_4677,N_4493);
nand U5866 (N_5866,N_3888,N_2696);
and U5867 (N_5867,N_4974,N_2855);
and U5868 (N_5868,N_3685,N_4133);
or U5869 (N_5869,N_4172,N_4624);
nor U5870 (N_5870,N_4134,N_2741);
or U5871 (N_5871,N_4131,N_4272);
nor U5872 (N_5872,N_4707,N_4092);
nor U5873 (N_5873,N_3792,N_2553);
or U5874 (N_5874,N_3041,N_4000);
nand U5875 (N_5875,N_4353,N_4569);
nand U5876 (N_5876,N_4324,N_4678);
nand U5877 (N_5877,N_3089,N_3975);
nor U5878 (N_5878,N_4178,N_2507);
or U5879 (N_5879,N_4953,N_2981);
and U5880 (N_5880,N_3424,N_2635);
nand U5881 (N_5881,N_3416,N_2535);
or U5882 (N_5882,N_4036,N_4512);
nand U5883 (N_5883,N_4937,N_3171);
and U5884 (N_5884,N_2756,N_4765);
and U5885 (N_5885,N_4832,N_3637);
and U5886 (N_5886,N_3449,N_4502);
or U5887 (N_5887,N_4367,N_3742);
nand U5888 (N_5888,N_4629,N_4170);
or U5889 (N_5889,N_4171,N_3538);
nand U5890 (N_5890,N_2911,N_4442);
and U5891 (N_5891,N_3684,N_4372);
or U5892 (N_5892,N_2849,N_4645);
nand U5893 (N_5893,N_4338,N_3208);
and U5894 (N_5894,N_3156,N_2867);
nand U5895 (N_5895,N_4412,N_2800);
nand U5896 (N_5896,N_4140,N_4237);
nor U5897 (N_5897,N_3370,N_3154);
nand U5898 (N_5898,N_4461,N_4663);
nor U5899 (N_5899,N_2595,N_4076);
and U5900 (N_5900,N_4477,N_3353);
and U5901 (N_5901,N_4801,N_4658);
and U5902 (N_5902,N_3390,N_4571);
and U5903 (N_5903,N_2757,N_3900);
xor U5904 (N_5904,N_4946,N_3364);
nor U5905 (N_5905,N_3127,N_2632);
or U5906 (N_5906,N_2879,N_3659);
nor U5907 (N_5907,N_4680,N_4323);
and U5908 (N_5908,N_3608,N_3927);
nand U5909 (N_5909,N_2742,N_2977);
nand U5910 (N_5910,N_3756,N_4754);
and U5911 (N_5911,N_2567,N_4263);
or U5912 (N_5912,N_3536,N_3839);
and U5913 (N_5913,N_3511,N_2580);
or U5914 (N_5914,N_4464,N_3229);
nor U5915 (N_5915,N_2869,N_3412);
and U5916 (N_5916,N_2784,N_4022);
nand U5917 (N_5917,N_4577,N_3178);
nor U5918 (N_5918,N_4308,N_4410);
or U5919 (N_5919,N_3830,N_3175);
xnor U5920 (N_5920,N_4073,N_3525);
or U5921 (N_5921,N_3860,N_3537);
nor U5922 (N_5922,N_4871,N_4607);
xor U5923 (N_5923,N_4698,N_4735);
or U5924 (N_5924,N_3763,N_2798);
nor U5925 (N_5925,N_3844,N_2779);
nor U5926 (N_5926,N_2782,N_4555);
nor U5927 (N_5927,N_2745,N_4861);
nor U5928 (N_5928,N_3293,N_2536);
xor U5929 (N_5929,N_2502,N_4248);
and U5930 (N_5930,N_2657,N_3423);
and U5931 (N_5931,N_4893,N_3784);
and U5932 (N_5932,N_2725,N_2525);
nand U5933 (N_5933,N_2636,N_4152);
and U5934 (N_5934,N_4520,N_4556);
nand U5935 (N_5935,N_3457,N_4199);
and U5936 (N_5936,N_4382,N_3654);
nor U5937 (N_5937,N_2937,N_2904);
nand U5938 (N_5938,N_3660,N_2520);
nor U5939 (N_5939,N_3481,N_3083);
nor U5940 (N_5940,N_4719,N_2917);
nand U5941 (N_5941,N_2922,N_2924);
or U5942 (N_5942,N_3668,N_3298);
xnor U5943 (N_5943,N_3147,N_4489);
or U5944 (N_5944,N_3087,N_4113);
nor U5945 (N_5945,N_3718,N_3242);
xor U5946 (N_5946,N_4180,N_2560);
and U5947 (N_5947,N_2760,N_3311);
and U5948 (N_5948,N_4023,N_3523);
or U5949 (N_5949,N_4163,N_2854);
and U5950 (N_5950,N_4074,N_2568);
nor U5951 (N_5951,N_4996,N_3266);
nand U5952 (N_5952,N_3984,N_4196);
nand U5953 (N_5953,N_4510,N_4964);
nand U5954 (N_5954,N_3576,N_3772);
or U5955 (N_5955,N_4397,N_2693);
nor U5956 (N_5956,N_4234,N_2778);
or U5957 (N_5957,N_3667,N_3859);
or U5958 (N_5958,N_4295,N_2537);
nor U5959 (N_5959,N_4167,N_4839);
nand U5960 (N_5960,N_4018,N_4432);
and U5961 (N_5961,N_4756,N_2662);
nor U5962 (N_5962,N_3941,N_4350);
and U5963 (N_5963,N_3998,N_4876);
nor U5964 (N_5964,N_4491,N_2638);
or U5965 (N_5965,N_3520,N_3111);
or U5966 (N_5966,N_2640,N_2926);
xor U5967 (N_5967,N_3552,N_4700);
nor U5968 (N_5968,N_3064,N_3565);
nand U5969 (N_5969,N_4033,N_4145);
nand U5970 (N_5970,N_4872,N_4071);
xor U5971 (N_5971,N_4925,N_2682);
nor U5972 (N_5972,N_3777,N_2556);
xor U5973 (N_5973,N_4517,N_3837);
nor U5974 (N_5974,N_4437,N_3686);
and U5975 (N_5975,N_2733,N_4757);
or U5976 (N_5976,N_4056,N_4385);
nand U5977 (N_5977,N_3708,N_3605);
nor U5978 (N_5978,N_4212,N_4729);
or U5979 (N_5979,N_3226,N_4784);
nand U5980 (N_5980,N_3801,N_3897);
xor U5981 (N_5981,N_4970,N_4814);
or U5982 (N_5982,N_3658,N_4810);
nor U5983 (N_5983,N_3273,N_3924);
or U5984 (N_5984,N_3630,N_2835);
nor U5985 (N_5985,N_3791,N_3914);
nand U5986 (N_5986,N_3812,N_4896);
xnor U5987 (N_5987,N_4932,N_3979);
nand U5988 (N_5988,N_2771,N_3464);
and U5989 (N_5989,N_3921,N_4751);
nand U5990 (N_5990,N_4743,N_2533);
nand U5991 (N_5991,N_3325,N_2921);
nand U5992 (N_5992,N_4043,N_4013);
nand U5993 (N_5993,N_4189,N_2531);
nor U5994 (N_5994,N_3415,N_3167);
nor U5995 (N_5995,N_4206,N_3391);
and U5996 (N_5996,N_3287,N_3396);
and U5997 (N_5997,N_3244,N_4004);
nor U5998 (N_5998,N_4802,N_4661);
or U5999 (N_5999,N_4712,N_4069);
nor U6000 (N_6000,N_4335,N_4975);
or U6001 (N_6001,N_3617,N_3221);
or U6002 (N_6002,N_4601,N_4423);
and U6003 (N_6003,N_4088,N_3487);
nor U6004 (N_6004,N_3358,N_3377);
xor U6005 (N_6005,N_4849,N_2707);
nand U6006 (N_6006,N_2847,N_2913);
and U6007 (N_6007,N_4529,N_3776);
nor U6008 (N_6008,N_3022,N_4943);
xnor U6009 (N_6009,N_3117,N_2834);
xor U6010 (N_6010,N_2700,N_4617);
nand U6011 (N_6011,N_3055,N_2927);
nor U6012 (N_6012,N_3947,N_4824);
nand U6013 (N_6013,N_2821,N_4289);
or U6014 (N_6014,N_4862,N_3754);
and U6015 (N_6015,N_4500,N_3057);
and U6016 (N_6016,N_3459,N_2617);
or U6017 (N_6017,N_3507,N_4355);
nand U6018 (N_6018,N_4322,N_2721);
and U6019 (N_6019,N_2877,N_3967);
nor U6020 (N_6020,N_4651,N_4912);
xnor U6021 (N_6021,N_4292,N_4143);
or U6022 (N_6022,N_4117,N_3037);
nand U6023 (N_6023,N_2956,N_4888);
or U6024 (N_6024,N_3697,N_3504);
nor U6025 (N_6025,N_3705,N_2882);
nand U6026 (N_6026,N_3333,N_4303);
nand U6027 (N_6027,N_4318,N_2750);
or U6028 (N_6028,N_3515,N_3762);
nor U6029 (N_6029,N_4219,N_3279);
or U6030 (N_6030,N_2794,N_3474);
or U6031 (N_6031,N_3646,N_4472);
xnor U6032 (N_6032,N_2501,N_4027);
and U6033 (N_6033,N_3598,N_4549);
or U6034 (N_6034,N_3188,N_3556);
or U6035 (N_6035,N_4648,N_3899);
and U6036 (N_6036,N_4008,N_2871);
and U6037 (N_6037,N_3439,N_3615);
nand U6038 (N_6038,N_2773,N_3993);
xnor U6039 (N_6039,N_3528,N_3806);
and U6040 (N_6040,N_4446,N_3785);
or U6041 (N_6041,N_3676,N_3753);
nor U6042 (N_6042,N_2549,N_4806);
xor U6043 (N_6043,N_2544,N_2873);
nand U6044 (N_6044,N_3714,N_4674);
nand U6045 (N_6045,N_3091,N_2785);
xnor U6046 (N_6046,N_4780,N_4514);
and U6047 (N_6047,N_3480,N_2723);
nand U6048 (N_6048,N_4931,N_4685);
and U6049 (N_6049,N_3855,N_4340);
nor U6050 (N_6050,N_4609,N_3919);
nand U6051 (N_6051,N_4686,N_2991);
nor U6052 (N_6052,N_2630,N_2971);
nor U6053 (N_6053,N_3450,N_4718);
and U6054 (N_6054,N_4546,N_3194);
or U6055 (N_6055,N_2843,N_3863);
and U6056 (N_6056,N_3259,N_4293);
and U6057 (N_6057,N_4637,N_3102);
or U6058 (N_6058,N_2647,N_2965);
or U6059 (N_6059,N_3716,N_2957);
nor U6060 (N_6060,N_4174,N_2574);
and U6061 (N_6061,N_4141,N_4105);
or U6062 (N_6062,N_3347,N_2624);
and U6063 (N_6063,N_2899,N_3463);
nand U6064 (N_6064,N_4029,N_4885);
nor U6065 (N_6065,N_4261,N_2590);
nor U6066 (N_6066,N_2685,N_4593);
nor U6067 (N_6067,N_2923,N_3710);
nor U6068 (N_6068,N_4175,N_3700);
nor U6069 (N_6069,N_3648,N_4453);
nor U6070 (N_6070,N_4823,N_4256);
and U6071 (N_6071,N_4845,N_3970);
and U6072 (N_6072,N_3735,N_3315);
and U6073 (N_6073,N_4190,N_3864);
nand U6074 (N_6074,N_4621,N_3790);
or U6075 (N_6075,N_4240,N_4330);
nor U6076 (N_6076,N_4136,N_4299);
or U6077 (N_6077,N_4992,N_4011);
nand U6078 (N_6078,N_4127,N_4067);
or U6079 (N_6079,N_4501,N_3121);
and U6080 (N_6080,N_4826,N_3114);
or U6081 (N_6081,N_2530,N_4590);
or U6082 (N_6082,N_2825,N_3438);
nand U6083 (N_6083,N_4538,N_3151);
nor U6084 (N_6084,N_3033,N_4914);
and U6085 (N_6085,N_3594,N_3126);
and U6086 (N_6086,N_3319,N_4285);
or U6087 (N_6087,N_4669,N_3403);
xor U6088 (N_6088,N_4007,N_2906);
xnor U6089 (N_6089,N_2992,N_4988);
xor U6090 (N_6090,N_3363,N_3440);
and U6091 (N_6091,N_3150,N_4487);
and U6092 (N_6092,N_4591,N_4684);
nor U6093 (N_6093,N_4704,N_3866);
and U6094 (N_6094,N_2652,N_3441);
and U6095 (N_6095,N_4508,N_3216);
nor U6096 (N_6096,N_3610,N_4695);
nand U6097 (N_6097,N_4268,N_3044);
nor U6098 (N_6098,N_4457,N_2874);
or U6099 (N_6099,N_2540,N_4958);
or U6100 (N_6100,N_2606,N_4049);
nor U6101 (N_6101,N_4287,N_4309);
and U6102 (N_6102,N_2987,N_2597);
nor U6103 (N_6103,N_3113,N_2565);
nor U6104 (N_6104,N_2664,N_4746);
or U6105 (N_6105,N_3562,N_3982);
and U6106 (N_6106,N_4456,N_3758);
nand U6107 (N_6107,N_3831,N_2930);
nor U6108 (N_6108,N_3621,N_3618);
nand U6109 (N_6109,N_4081,N_4665);
nand U6110 (N_6110,N_4527,N_4378);
or U6111 (N_6111,N_4361,N_3846);
and U6112 (N_6112,N_4344,N_4251);
or U6113 (N_6113,N_4993,N_4561);
nand U6114 (N_6114,N_4002,N_3657);
and U6115 (N_6115,N_3465,N_3737);
or U6116 (N_6116,N_3168,N_4582);
xor U6117 (N_6117,N_3745,N_2933);
or U6118 (N_6118,N_3383,N_2607);
nand U6119 (N_6119,N_2908,N_3581);
or U6120 (N_6120,N_4890,N_3558);
or U6121 (N_6121,N_3344,N_3612);
nand U6122 (N_6122,N_3656,N_4834);
and U6123 (N_6123,N_3334,N_3342);
nor U6124 (N_6124,N_2887,N_4454);
nand U6125 (N_6125,N_3550,N_2665);
nor U6126 (N_6126,N_3841,N_2935);
xor U6127 (N_6127,N_4654,N_2768);
xor U6128 (N_6128,N_3669,N_4722);
xnor U6129 (N_6129,N_3963,N_3687);
or U6130 (N_6130,N_3145,N_3651);
and U6131 (N_6131,N_2979,N_2573);
nor U6132 (N_6132,N_4075,N_2903);
nand U6133 (N_6133,N_4009,N_3521);
xor U6134 (N_6134,N_4777,N_3603);
or U6135 (N_6135,N_4038,N_3240);
nor U6136 (N_6136,N_4820,N_3461);
and U6137 (N_6137,N_4468,N_4100);
or U6138 (N_6138,N_2680,N_4770);
nand U6139 (N_6139,N_2860,N_3431);
xnor U6140 (N_6140,N_3786,N_2892);
nor U6141 (N_6141,N_4744,N_3290);
and U6142 (N_6142,N_3729,N_4014);
nand U6143 (N_6143,N_3539,N_3275);
nor U6144 (N_6144,N_3788,N_3376);
nor U6145 (N_6145,N_3034,N_2986);
nor U6146 (N_6146,N_4028,N_4020);
and U6147 (N_6147,N_3153,N_4444);
and U6148 (N_6148,N_4376,N_4910);
nand U6149 (N_6149,N_3452,N_4304);
and U6150 (N_6150,N_4144,N_4460);
nor U6151 (N_6151,N_4176,N_3419);
and U6152 (N_6152,N_4267,N_2734);
nand U6153 (N_6153,N_4887,N_3222);
nand U6154 (N_6154,N_4797,N_2739);
nand U6155 (N_6155,N_2758,N_4494);
nor U6156 (N_6156,N_4107,N_4021);
and U6157 (N_6157,N_4093,N_4850);
and U6158 (N_6158,N_4981,N_2814);
nor U6159 (N_6159,N_3709,N_2945);
nand U6160 (N_6160,N_4838,N_3769);
nor U6161 (N_6161,N_4659,N_3805);
and U6162 (N_6162,N_4246,N_4419);
and U6163 (N_6163,N_3100,N_3600);
nand U6164 (N_6164,N_2666,N_3346);
or U6165 (N_6165,N_2743,N_2780);
and U6166 (N_6166,N_3972,N_4386);
xnor U6167 (N_6167,N_2575,N_2681);
or U6168 (N_6168,N_4404,N_2683);
nor U6169 (N_6169,N_4949,N_3215);
and U6170 (N_6170,N_4919,N_3061);
nor U6171 (N_6171,N_4365,N_4326);
and U6172 (N_6172,N_2928,N_3016);
nand U6173 (N_6173,N_4091,N_4313);
and U6174 (N_6174,N_2958,N_2876);
and U6175 (N_6175,N_2709,N_3473);
nor U6176 (N_6176,N_2596,N_4954);
and U6177 (N_6177,N_3976,N_3099);
and U6178 (N_6178,N_2705,N_3930);
and U6179 (N_6179,N_2694,N_4955);
or U6180 (N_6180,N_2706,N_3966);
nand U6181 (N_6181,N_4184,N_3340);
nand U6182 (N_6182,N_4484,N_4356);
nor U6183 (N_6183,N_4800,N_3529);
and U6184 (N_6184,N_3313,N_4761);
and U6185 (N_6185,N_3106,N_3399);
nor U6186 (N_6186,N_4619,N_3495);
and U6187 (N_6187,N_3060,N_4148);
nand U6188 (N_6188,N_3059,N_4898);
and U6189 (N_6189,N_3365,N_4345);
nor U6190 (N_6190,N_2702,N_4899);
and U6191 (N_6191,N_3413,N_4752);
nand U6192 (N_6192,N_3048,N_3645);
xor U6193 (N_6193,N_4061,N_4837);
nand U6194 (N_6194,N_3312,N_3267);
nor U6195 (N_6195,N_4812,N_2547);
nor U6196 (N_6196,N_4334,N_2900);
and U6197 (N_6197,N_4443,N_4909);
nand U6198 (N_6198,N_3678,N_4438);
nor U6199 (N_6199,N_3021,N_3141);
or U6200 (N_6200,N_2552,N_4809);
or U6201 (N_6201,N_2801,N_2967);
xnor U6202 (N_6202,N_4006,N_4302);
and U6203 (N_6203,N_2808,N_3981);
xor U6204 (N_6204,N_4804,N_3643);
or U6205 (N_6205,N_4343,N_2907);
or U6206 (N_6206,N_3362,N_4901);
nor U6207 (N_6207,N_4738,N_3744);
xor U6208 (N_6208,N_3701,N_4626);
nor U6209 (N_6209,N_4149,N_4947);
nor U6210 (N_6210,N_4151,N_3332);
nand U6211 (N_6211,N_3992,N_3418);
or U6212 (N_6212,N_3316,N_2791);
nand U6213 (N_6213,N_4371,N_3601);
or U6214 (N_6214,N_3885,N_3699);
or U6215 (N_6215,N_2592,N_3130);
nand U6216 (N_6216,N_3307,N_3300);
or U6217 (N_6217,N_2646,N_3532);
xnor U6218 (N_6218,N_4616,N_3580);
and U6219 (N_6219,N_3425,N_2534);
and U6220 (N_6220,N_4153,N_4522);
and U6221 (N_6221,N_2603,N_3274);
or U6222 (N_6222,N_2698,N_3804);
xnor U6223 (N_6223,N_2503,N_2736);
or U6224 (N_6224,N_3471,N_3858);
or U6225 (N_6225,N_2634,N_2550);
nand U6226 (N_6226,N_4971,N_3483);
nor U6227 (N_6227,N_4847,N_4224);
or U6228 (N_6228,N_4118,N_4103);
or U6229 (N_6229,N_4597,N_4936);
and U6230 (N_6230,N_3134,N_3750);
nor U6231 (N_6231,N_3241,N_3962);
nand U6232 (N_6232,N_4150,N_4895);
xor U6233 (N_6233,N_4737,N_2915);
nand U6234 (N_6234,N_3571,N_3136);
or U6235 (N_6235,N_4956,N_3816);
and U6236 (N_6236,N_3808,N_3987);
nor U6237 (N_6237,N_4968,N_3448);
or U6238 (N_6238,N_2841,N_3545);
xnor U6239 (N_6239,N_3220,N_3429);
nor U6240 (N_6240,N_3872,N_3051);
or U6241 (N_6241,N_2701,N_3157);
or U6242 (N_6242,N_3531,N_4551);
or U6243 (N_6243,N_3673,N_4244);
and U6244 (N_6244,N_3260,N_3324);
or U6245 (N_6245,N_4611,N_4653);
nor U6246 (N_6246,N_3775,N_3185);
nor U6247 (N_6247,N_4173,N_2713);
and U6248 (N_6248,N_3125,N_4575);
nor U6249 (N_6249,N_4435,N_4866);
and U6250 (N_6250,N_2611,N_4453);
or U6251 (N_6251,N_4896,N_3315);
and U6252 (N_6252,N_4666,N_3271);
or U6253 (N_6253,N_3467,N_3583);
nand U6254 (N_6254,N_4357,N_4499);
and U6255 (N_6255,N_2582,N_4690);
or U6256 (N_6256,N_4472,N_2948);
nand U6257 (N_6257,N_4527,N_2527);
or U6258 (N_6258,N_3659,N_3840);
nand U6259 (N_6259,N_4177,N_4460);
nand U6260 (N_6260,N_2819,N_3985);
and U6261 (N_6261,N_4880,N_2794);
and U6262 (N_6262,N_4522,N_4298);
and U6263 (N_6263,N_4807,N_3545);
or U6264 (N_6264,N_2563,N_4736);
nand U6265 (N_6265,N_4227,N_3069);
or U6266 (N_6266,N_3160,N_4156);
nand U6267 (N_6267,N_3362,N_4037);
or U6268 (N_6268,N_3425,N_3108);
nor U6269 (N_6269,N_3113,N_3803);
or U6270 (N_6270,N_2629,N_3089);
or U6271 (N_6271,N_3229,N_2528);
or U6272 (N_6272,N_3792,N_4093);
and U6273 (N_6273,N_4560,N_2810);
and U6274 (N_6274,N_3786,N_2624);
nand U6275 (N_6275,N_3067,N_3099);
or U6276 (N_6276,N_4871,N_4316);
or U6277 (N_6277,N_3578,N_3586);
and U6278 (N_6278,N_2898,N_4163);
or U6279 (N_6279,N_3478,N_4954);
nor U6280 (N_6280,N_2581,N_4112);
nand U6281 (N_6281,N_2646,N_3234);
nor U6282 (N_6282,N_4687,N_3864);
or U6283 (N_6283,N_4814,N_4702);
nor U6284 (N_6284,N_3395,N_3171);
nor U6285 (N_6285,N_4885,N_4095);
nand U6286 (N_6286,N_2800,N_3957);
nor U6287 (N_6287,N_3541,N_2873);
xor U6288 (N_6288,N_4709,N_4814);
nor U6289 (N_6289,N_3480,N_2847);
or U6290 (N_6290,N_3157,N_3115);
or U6291 (N_6291,N_4182,N_3577);
or U6292 (N_6292,N_3283,N_4373);
or U6293 (N_6293,N_4541,N_2918);
nor U6294 (N_6294,N_2812,N_3412);
nor U6295 (N_6295,N_4403,N_4170);
or U6296 (N_6296,N_4792,N_3973);
and U6297 (N_6297,N_3246,N_3367);
nor U6298 (N_6298,N_3649,N_4944);
or U6299 (N_6299,N_4572,N_4628);
or U6300 (N_6300,N_4811,N_3420);
nor U6301 (N_6301,N_4772,N_4620);
or U6302 (N_6302,N_3436,N_3836);
nand U6303 (N_6303,N_3961,N_2599);
nand U6304 (N_6304,N_2846,N_3073);
and U6305 (N_6305,N_2811,N_2783);
nor U6306 (N_6306,N_4906,N_3215);
nand U6307 (N_6307,N_4961,N_2948);
and U6308 (N_6308,N_4088,N_4577);
and U6309 (N_6309,N_2923,N_3280);
nor U6310 (N_6310,N_3589,N_3563);
nor U6311 (N_6311,N_4582,N_4213);
xnor U6312 (N_6312,N_4467,N_4746);
and U6313 (N_6313,N_4112,N_2513);
nor U6314 (N_6314,N_3091,N_3899);
and U6315 (N_6315,N_4041,N_3001);
and U6316 (N_6316,N_3115,N_4568);
and U6317 (N_6317,N_4519,N_3869);
or U6318 (N_6318,N_2616,N_3611);
and U6319 (N_6319,N_3876,N_3079);
nand U6320 (N_6320,N_3085,N_4103);
or U6321 (N_6321,N_4294,N_2619);
nor U6322 (N_6322,N_3429,N_4494);
nand U6323 (N_6323,N_3924,N_2960);
or U6324 (N_6324,N_4884,N_3184);
and U6325 (N_6325,N_4762,N_2777);
and U6326 (N_6326,N_4411,N_4441);
and U6327 (N_6327,N_4877,N_3330);
nor U6328 (N_6328,N_4414,N_3288);
or U6329 (N_6329,N_2654,N_3391);
xnor U6330 (N_6330,N_3076,N_3843);
and U6331 (N_6331,N_4964,N_3030);
nor U6332 (N_6332,N_2602,N_3397);
nand U6333 (N_6333,N_3165,N_4203);
nor U6334 (N_6334,N_3069,N_4504);
nor U6335 (N_6335,N_4837,N_2807);
and U6336 (N_6336,N_4862,N_3693);
nor U6337 (N_6337,N_4477,N_4772);
nand U6338 (N_6338,N_4123,N_3879);
nor U6339 (N_6339,N_3992,N_4022);
and U6340 (N_6340,N_2941,N_3932);
or U6341 (N_6341,N_3849,N_4925);
nand U6342 (N_6342,N_4149,N_2875);
and U6343 (N_6343,N_3599,N_2894);
xor U6344 (N_6344,N_4886,N_2681);
nand U6345 (N_6345,N_4789,N_3697);
nor U6346 (N_6346,N_2629,N_4612);
or U6347 (N_6347,N_3863,N_2779);
nor U6348 (N_6348,N_4862,N_4795);
nor U6349 (N_6349,N_3429,N_4833);
nor U6350 (N_6350,N_4475,N_4969);
xor U6351 (N_6351,N_3494,N_3082);
and U6352 (N_6352,N_2857,N_3004);
nand U6353 (N_6353,N_4074,N_2964);
or U6354 (N_6354,N_3037,N_3637);
or U6355 (N_6355,N_4284,N_4698);
nor U6356 (N_6356,N_3168,N_4000);
nand U6357 (N_6357,N_3246,N_4658);
or U6358 (N_6358,N_2715,N_4912);
or U6359 (N_6359,N_3470,N_3409);
or U6360 (N_6360,N_4127,N_2757);
nor U6361 (N_6361,N_4996,N_3851);
nor U6362 (N_6362,N_2666,N_2927);
or U6363 (N_6363,N_2639,N_4838);
or U6364 (N_6364,N_3924,N_4613);
nor U6365 (N_6365,N_4064,N_3740);
nand U6366 (N_6366,N_3035,N_3767);
or U6367 (N_6367,N_3129,N_3627);
xor U6368 (N_6368,N_4650,N_2647);
nand U6369 (N_6369,N_4957,N_4961);
and U6370 (N_6370,N_4979,N_4411);
nor U6371 (N_6371,N_4419,N_4752);
or U6372 (N_6372,N_2803,N_3863);
or U6373 (N_6373,N_4640,N_2795);
and U6374 (N_6374,N_4644,N_3018);
or U6375 (N_6375,N_2881,N_4652);
and U6376 (N_6376,N_3508,N_2535);
and U6377 (N_6377,N_4437,N_4191);
nor U6378 (N_6378,N_4832,N_4885);
and U6379 (N_6379,N_3976,N_4635);
and U6380 (N_6380,N_4439,N_2683);
nand U6381 (N_6381,N_2841,N_4445);
and U6382 (N_6382,N_4013,N_3608);
nor U6383 (N_6383,N_3376,N_2833);
nand U6384 (N_6384,N_3660,N_4921);
nand U6385 (N_6385,N_2857,N_3328);
and U6386 (N_6386,N_4232,N_4872);
nor U6387 (N_6387,N_2969,N_4632);
nor U6388 (N_6388,N_2964,N_2984);
or U6389 (N_6389,N_3608,N_4570);
nand U6390 (N_6390,N_2697,N_2907);
and U6391 (N_6391,N_4913,N_4666);
nand U6392 (N_6392,N_4207,N_3170);
or U6393 (N_6393,N_3013,N_3094);
xnor U6394 (N_6394,N_2915,N_3051);
and U6395 (N_6395,N_3320,N_3932);
or U6396 (N_6396,N_4115,N_2994);
nand U6397 (N_6397,N_3045,N_4070);
nor U6398 (N_6398,N_2817,N_4125);
nor U6399 (N_6399,N_2886,N_3919);
and U6400 (N_6400,N_2780,N_4054);
and U6401 (N_6401,N_3217,N_2634);
xnor U6402 (N_6402,N_4349,N_4307);
nor U6403 (N_6403,N_3988,N_4625);
and U6404 (N_6404,N_3729,N_4552);
nand U6405 (N_6405,N_3129,N_3043);
nor U6406 (N_6406,N_4904,N_3943);
or U6407 (N_6407,N_2657,N_3844);
or U6408 (N_6408,N_4503,N_3631);
or U6409 (N_6409,N_4502,N_4120);
nor U6410 (N_6410,N_4496,N_4906);
nand U6411 (N_6411,N_2675,N_3570);
and U6412 (N_6412,N_2718,N_4084);
nand U6413 (N_6413,N_2905,N_3053);
or U6414 (N_6414,N_4545,N_3988);
or U6415 (N_6415,N_2839,N_3639);
nand U6416 (N_6416,N_3117,N_3559);
nor U6417 (N_6417,N_3365,N_2681);
xnor U6418 (N_6418,N_3619,N_2546);
xor U6419 (N_6419,N_4225,N_4813);
nor U6420 (N_6420,N_3271,N_3996);
or U6421 (N_6421,N_3216,N_4100);
nor U6422 (N_6422,N_4368,N_4928);
nor U6423 (N_6423,N_4689,N_3512);
and U6424 (N_6424,N_2675,N_4163);
xnor U6425 (N_6425,N_2516,N_3321);
and U6426 (N_6426,N_2989,N_4744);
or U6427 (N_6427,N_2688,N_4439);
nand U6428 (N_6428,N_3968,N_4884);
nand U6429 (N_6429,N_2600,N_4318);
and U6430 (N_6430,N_3535,N_3737);
nor U6431 (N_6431,N_4859,N_3334);
nor U6432 (N_6432,N_3973,N_4464);
nor U6433 (N_6433,N_4251,N_3581);
or U6434 (N_6434,N_4993,N_2911);
or U6435 (N_6435,N_3224,N_2867);
or U6436 (N_6436,N_2911,N_3139);
and U6437 (N_6437,N_4754,N_3708);
xnor U6438 (N_6438,N_3904,N_3708);
nor U6439 (N_6439,N_3410,N_2609);
nand U6440 (N_6440,N_4964,N_4466);
nor U6441 (N_6441,N_3689,N_4591);
and U6442 (N_6442,N_3668,N_4808);
and U6443 (N_6443,N_2958,N_3826);
xnor U6444 (N_6444,N_2961,N_3519);
or U6445 (N_6445,N_3317,N_3973);
nand U6446 (N_6446,N_2894,N_2545);
and U6447 (N_6447,N_2656,N_3842);
or U6448 (N_6448,N_3016,N_2526);
xor U6449 (N_6449,N_3313,N_3304);
nand U6450 (N_6450,N_3369,N_4952);
or U6451 (N_6451,N_3285,N_4088);
nor U6452 (N_6452,N_2708,N_4174);
xnor U6453 (N_6453,N_2814,N_3726);
nand U6454 (N_6454,N_3288,N_2652);
or U6455 (N_6455,N_4357,N_3876);
nor U6456 (N_6456,N_2976,N_2556);
or U6457 (N_6457,N_2750,N_2748);
nor U6458 (N_6458,N_4458,N_4265);
nand U6459 (N_6459,N_4742,N_3853);
or U6460 (N_6460,N_2651,N_2843);
and U6461 (N_6461,N_3705,N_4498);
nand U6462 (N_6462,N_3038,N_3210);
nor U6463 (N_6463,N_2998,N_4620);
or U6464 (N_6464,N_3835,N_4298);
and U6465 (N_6465,N_4245,N_3621);
nand U6466 (N_6466,N_3431,N_4058);
and U6467 (N_6467,N_4021,N_3764);
nor U6468 (N_6468,N_2673,N_3756);
and U6469 (N_6469,N_2952,N_3601);
or U6470 (N_6470,N_4696,N_3737);
or U6471 (N_6471,N_3277,N_3857);
or U6472 (N_6472,N_4342,N_4753);
nand U6473 (N_6473,N_2926,N_2801);
or U6474 (N_6474,N_3525,N_2926);
nand U6475 (N_6475,N_3585,N_3987);
nand U6476 (N_6476,N_3016,N_4501);
nand U6477 (N_6477,N_2999,N_2719);
and U6478 (N_6478,N_2675,N_4092);
or U6479 (N_6479,N_2511,N_4479);
and U6480 (N_6480,N_3332,N_2807);
nand U6481 (N_6481,N_4213,N_4957);
nor U6482 (N_6482,N_3251,N_4742);
nor U6483 (N_6483,N_3980,N_3632);
or U6484 (N_6484,N_3235,N_3512);
or U6485 (N_6485,N_4025,N_4149);
nor U6486 (N_6486,N_4671,N_3974);
nor U6487 (N_6487,N_4018,N_4194);
and U6488 (N_6488,N_4494,N_4619);
nor U6489 (N_6489,N_3018,N_4383);
nor U6490 (N_6490,N_4562,N_4813);
or U6491 (N_6491,N_3260,N_3909);
or U6492 (N_6492,N_4423,N_2974);
or U6493 (N_6493,N_3370,N_2879);
nor U6494 (N_6494,N_4678,N_4939);
nor U6495 (N_6495,N_2966,N_3539);
and U6496 (N_6496,N_2867,N_3400);
and U6497 (N_6497,N_3564,N_4011);
and U6498 (N_6498,N_2864,N_3492);
or U6499 (N_6499,N_3240,N_2804);
or U6500 (N_6500,N_3339,N_2724);
nor U6501 (N_6501,N_4030,N_4885);
and U6502 (N_6502,N_3214,N_2673);
nand U6503 (N_6503,N_4063,N_2976);
nand U6504 (N_6504,N_4923,N_3135);
nand U6505 (N_6505,N_3450,N_3638);
or U6506 (N_6506,N_3703,N_4126);
or U6507 (N_6507,N_2678,N_3297);
nand U6508 (N_6508,N_3465,N_3570);
and U6509 (N_6509,N_3901,N_2827);
nor U6510 (N_6510,N_4493,N_4739);
nor U6511 (N_6511,N_3321,N_3036);
nand U6512 (N_6512,N_3294,N_4934);
or U6513 (N_6513,N_3448,N_4528);
nand U6514 (N_6514,N_4004,N_2768);
nor U6515 (N_6515,N_3754,N_2653);
or U6516 (N_6516,N_4198,N_3646);
nand U6517 (N_6517,N_4770,N_3240);
or U6518 (N_6518,N_4489,N_4346);
or U6519 (N_6519,N_3888,N_4301);
xnor U6520 (N_6520,N_3797,N_4651);
or U6521 (N_6521,N_3464,N_2996);
or U6522 (N_6522,N_4638,N_3864);
and U6523 (N_6523,N_3608,N_4347);
nand U6524 (N_6524,N_4309,N_3861);
nand U6525 (N_6525,N_2662,N_3701);
nand U6526 (N_6526,N_3955,N_4313);
nor U6527 (N_6527,N_3457,N_2745);
nand U6528 (N_6528,N_2733,N_3529);
and U6529 (N_6529,N_3318,N_3253);
or U6530 (N_6530,N_3370,N_4682);
nor U6531 (N_6531,N_4776,N_2550);
nor U6532 (N_6532,N_3818,N_3151);
and U6533 (N_6533,N_4684,N_3128);
nand U6534 (N_6534,N_2956,N_3989);
and U6535 (N_6535,N_3948,N_2792);
and U6536 (N_6536,N_4765,N_3624);
and U6537 (N_6537,N_3036,N_3992);
nor U6538 (N_6538,N_3247,N_2520);
nor U6539 (N_6539,N_4057,N_3542);
or U6540 (N_6540,N_3836,N_2641);
or U6541 (N_6541,N_4585,N_4324);
nor U6542 (N_6542,N_3299,N_3043);
xor U6543 (N_6543,N_3381,N_4114);
nor U6544 (N_6544,N_4727,N_4524);
nand U6545 (N_6545,N_3585,N_4440);
or U6546 (N_6546,N_3479,N_4383);
nor U6547 (N_6547,N_3262,N_2614);
nand U6548 (N_6548,N_3624,N_2632);
or U6549 (N_6549,N_4202,N_3358);
nand U6550 (N_6550,N_3933,N_4042);
and U6551 (N_6551,N_3164,N_3272);
and U6552 (N_6552,N_3299,N_4076);
nor U6553 (N_6553,N_2957,N_4282);
nand U6554 (N_6554,N_3062,N_2780);
nor U6555 (N_6555,N_3231,N_3081);
or U6556 (N_6556,N_3732,N_2694);
and U6557 (N_6557,N_2548,N_3990);
nand U6558 (N_6558,N_3370,N_2902);
or U6559 (N_6559,N_2829,N_3459);
nand U6560 (N_6560,N_3835,N_2703);
and U6561 (N_6561,N_4934,N_3098);
nand U6562 (N_6562,N_3685,N_2794);
nand U6563 (N_6563,N_3182,N_3399);
nand U6564 (N_6564,N_4557,N_2859);
nand U6565 (N_6565,N_4997,N_3769);
xnor U6566 (N_6566,N_4263,N_2511);
xnor U6567 (N_6567,N_3930,N_3472);
nor U6568 (N_6568,N_2973,N_4963);
and U6569 (N_6569,N_3579,N_4870);
and U6570 (N_6570,N_2775,N_4042);
or U6571 (N_6571,N_2636,N_4139);
and U6572 (N_6572,N_3698,N_3019);
nand U6573 (N_6573,N_2735,N_3731);
nor U6574 (N_6574,N_2553,N_4680);
nand U6575 (N_6575,N_4522,N_4481);
and U6576 (N_6576,N_4732,N_3930);
and U6577 (N_6577,N_4424,N_2780);
xnor U6578 (N_6578,N_2961,N_4965);
and U6579 (N_6579,N_3706,N_4972);
and U6580 (N_6580,N_3822,N_4103);
xor U6581 (N_6581,N_3778,N_2688);
nand U6582 (N_6582,N_4696,N_4438);
nand U6583 (N_6583,N_2821,N_4209);
nand U6584 (N_6584,N_2936,N_2752);
xnor U6585 (N_6585,N_3381,N_4541);
nor U6586 (N_6586,N_2785,N_4578);
or U6587 (N_6587,N_3616,N_4098);
nor U6588 (N_6588,N_4917,N_3776);
nor U6589 (N_6589,N_4740,N_3970);
or U6590 (N_6590,N_2625,N_4631);
or U6591 (N_6591,N_4643,N_4518);
xnor U6592 (N_6592,N_3535,N_3516);
nand U6593 (N_6593,N_3630,N_3600);
nand U6594 (N_6594,N_4924,N_4315);
nand U6595 (N_6595,N_4832,N_3930);
and U6596 (N_6596,N_2700,N_3799);
nand U6597 (N_6597,N_4597,N_4270);
and U6598 (N_6598,N_3089,N_3177);
nand U6599 (N_6599,N_4227,N_2820);
nand U6600 (N_6600,N_3249,N_4262);
xor U6601 (N_6601,N_4992,N_3435);
or U6602 (N_6602,N_4262,N_4258);
and U6603 (N_6603,N_4187,N_4115);
nand U6604 (N_6604,N_3359,N_3763);
and U6605 (N_6605,N_4508,N_3797);
or U6606 (N_6606,N_4312,N_3893);
xor U6607 (N_6607,N_2618,N_3436);
and U6608 (N_6608,N_3187,N_3629);
nand U6609 (N_6609,N_3987,N_3250);
nand U6610 (N_6610,N_3293,N_4754);
nor U6611 (N_6611,N_3649,N_3723);
nor U6612 (N_6612,N_4514,N_3101);
nand U6613 (N_6613,N_3536,N_2835);
or U6614 (N_6614,N_2892,N_3438);
xnor U6615 (N_6615,N_2950,N_3868);
nor U6616 (N_6616,N_3016,N_4749);
xor U6617 (N_6617,N_4304,N_2780);
or U6618 (N_6618,N_3538,N_3261);
nand U6619 (N_6619,N_3161,N_2623);
or U6620 (N_6620,N_4673,N_4634);
nand U6621 (N_6621,N_2645,N_2940);
nor U6622 (N_6622,N_2698,N_4059);
nor U6623 (N_6623,N_3810,N_3584);
or U6624 (N_6624,N_4530,N_4366);
nor U6625 (N_6625,N_4278,N_3958);
nor U6626 (N_6626,N_4270,N_3248);
nor U6627 (N_6627,N_3073,N_4816);
nand U6628 (N_6628,N_3822,N_4272);
nor U6629 (N_6629,N_4239,N_4695);
and U6630 (N_6630,N_3802,N_2859);
nand U6631 (N_6631,N_4268,N_4835);
nor U6632 (N_6632,N_4646,N_3532);
xnor U6633 (N_6633,N_4090,N_4513);
or U6634 (N_6634,N_3479,N_4333);
nand U6635 (N_6635,N_4494,N_2874);
nand U6636 (N_6636,N_4912,N_3816);
and U6637 (N_6637,N_4193,N_2764);
and U6638 (N_6638,N_4880,N_3258);
and U6639 (N_6639,N_3993,N_3296);
nand U6640 (N_6640,N_3794,N_2628);
and U6641 (N_6641,N_4385,N_4554);
nand U6642 (N_6642,N_4606,N_4409);
and U6643 (N_6643,N_4900,N_3891);
nor U6644 (N_6644,N_3622,N_3886);
xnor U6645 (N_6645,N_3906,N_4454);
xnor U6646 (N_6646,N_4937,N_2553);
nand U6647 (N_6647,N_4512,N_3814);
and U6648 (N_6648,N_3330,N_4046);
nand U6649 (N_6649,N_4249,N_4102);
xor U6650 (N_6650,N_4081,N_3028);
or U6651 (N_6651,N_4540,N_3200);
or U6652 (N_6652,N_4844,N_4236);
xor U6653 (N_6653,N_4017,N_4748);
xnor U6654 (N_6654,N_2661,N_3250);
and U6655 (N_6655,N_3376,N_4422);
and U6656 (N_6656,N_3883,N_3655);
or U6657 (N_6657,N_3635,N_3433);
nor U6658 (N_6658,N_4113,N_3663);
and U6659 (N_6659,N_4369,N_3551);
nor U6660 (N_6660,N_4393,N_2953);
nand U6661 (N_6661,N_2540,N_2570);
nand U6662 (N_6662,N_3203,N_2643);
nor U6663 (N_6663,N_2894,N_4600);
nor U6664 (N_6664,N_2594,N_4649);
and U6665 (N_6665,N_3466,N_2674);
and U6666 (N_6666,N_3515,N_2682);
nand U6667 (N_6667,N_4599,N_2533);
xnor U6668 (N_6668,N_2539,N_4808);
or U6669 (N_6669,N_4717,N_2644);
or U6670 (N_6670,N_4034,N_2631);
and U6671 (N_6671,N_4398,N_3071);
nor U6672 (N_6672,N_3683,N_3579);
or U6673 (N_6673,N_3264,N_3759);
and U6674 (N_6674,N_2606,N_3830);
nor U6675 (N_6675,N_3819,N_4795);
nor U6676 (N_6676,N_4606,N_4279);
or U6677 (N_6677,N_4862,N_3162);
or U6678 (N_6678,N_4971,N_3989);
and U6679 (N_6679,N_3375,N_2895);
nand U6680 (N_6680,N_3995,N_3493);
nand U6681 (N_6681,N_3685,N_4412);
and U6682 (N_6682,N_2555,N_4977);
nand U6683 (N_6683,N_4177,N_3227);
nand U6684 (N_6684,N_4279,N_4628);
or U6685 (N_6685,N_2613,N_4219);
or U6686 (N_6686,N_4118,N_4000);
nor U6687 (N_6687,N_4211,N_4806);
or U6688 (N_6688,N_4820,N_3910);
nor U6689 (N_6689,N_4187,N_4325);
nand U6690 (N_6690,N_4131,N_3580);
or U6691 (N_6691,N_3972,N_3429);
nor U6692 (N_6692,N_4214,N_3899);
nand U6693 (N_6693,N_2823,N_4264);
nand U6694 (N_6694,N_3533,N_3473);
nor U6695 (N_6695,N_4819,N_3013);
nor U6696 (N_6696,N_4287,N_4915);
nor U6697 (N_6697,N_3566,N_4152);
and U6698 (N_6698,N_4887,N_2696);
nand U6699 (N_6699,N_4073,N_4524);
nor U6700 (N_6700,N_2681,N_4198);
and U6701 (N_6701,N_4763,N_4305);
or U6702 (N_6702,N_2913,N_4210);
nor U6703 (N_6703,N_3724,N_3775);
nand U6704 (N_6704,N_3086,N_4696);
nand U6705 (N_6705,N_4756,N_3347);
nor U6706 (N_6706,N_3134,N_3287);
nand U6707 (N_6707,N_4850,N_2522);
nand U6708 (N_6708,N_3443,N_3153);
xor U6709 (N_6709,N_2577,N_3526);
nor U6710 (N_6710,N_4076,N_3846);
nor U6711 (N_6711,N_3289,N_2906);
nor U6712 (N_6712,N_2739,N_4740);
nand U6713 (N_6713,N_2762,N_4520);
nand U6714 (N_6714,N_3374,N_4904);
nand U6715 (N_6715,N_4350,N_3702);
nand U6716 (N_6716,N_4077,N_2861);
nor U6717 (N_6717,N_2679,N_4459);
or U6718 (N_6718,N_4815,N_3099);
or U6719 (N_6719,N_3336,N_3446);
nor U6720 (N_6720,N_3058,N_3786);
or U6721 (N_6721,N_2818,N_3205);
nand U6722 (N_6722,N_2976,N_4871);
or U6723 (N_6723,N_4003,N_4873);
nand U6724 (N_6724,N_3070,N_4354);
nand U6725 (N_6725,N_3074,N_3470);
and U6726 (N_6726,N_4066,N_3901);
nand U6727 (N_6727,N_4300,N_3041);
and U6728 (N_6728,N_3422,N_4068);
nand U6729 (N_6729,N_4577,N_3475);
xor U6730 (N_6730,N_2555,N_3249);
xor U6731 (N_6731,N_3520,N_4893);
nand U6732 (N_6732,N_3886,N_2595);
or U6733 (N_6733,N_2982,N_2693);
nor U6734 (N_6734,N_2876,N_3973);
nor U6735 (N_6735,N_3228,N_2537);
nor U6736 (N_6736,N_3231,N_3356);
and U6737 (N_6737,N_4187,N_3729);
and U6738 (N_6738,N_2541,N_2858);
and U6739 (N_6739,N_3823,N_4304);
or U6740 (N_6740,N_4245,N_3663);
nor U6741 (N_6741,N_4693,N_3711);
and U6742 (N_6742,N_3771,N_4989);
nor U6743 (N_6743,N_4425,N_2682);
nand U6744 (N_6744,N_4840,N_4688);
or U6745 (N_6745,N_3756,N_3299);
or U6746 (N_6746,N_3546,N_4894);
or U6747 (N_6747,N_2792,N_2612);
nor U6748 (N_6748,N_4050,N_3604);
xor U6749 (N_6749,N_4690,N_3777);
or U6750 (N_6750,N_3847,N_4781);
nand U6751 (N_6751,N_3552,N_4239);
and U6752 (N_6752,N_3533,N_2910);
and U6753 (N_6753,N_2620,N_4297);
and U6754 (N_6754,N_3884,N_2556);
nand U6755 (N_6755,N_4426,N_3358);
xnor U6756 (N_6756,N_3952,N_3388);
and U6757 (N_6757,N_3876,N_3878);
or U6758 (N_6758,N_4296,N_4619);
nand U6759 (N_6759,N_4570,N_3652);
or U6760 (N_6760,N_2744,N_3232);
nand U6761 (N_6761,N_2528,N_3227);
nor U6762 (N_6762,N_4024,N_4246);
and U6763 (N_6763,N_2708,N_3553);
or U6764 (N_6764,N_4270,N_4546);
nor U6765 (N_6765,N_3624,N_4811);
nor U6766 (N_6766,N_4494,N_2990);
nand U6767 (N_6767,N_3890,N_2625);
nor U6768 (N_6768,N_2795,N_3655);
or U6769 (N_6769,N_3421,N_3221);
and U6770 (N_6770,N_3082,N_4274);
and U6771 (N_6771,N_3698,N_4693);
or U6772 (N_6772,N_4534,N_3557);
or U6773 (N_6773,N_4258,N_4661);
nor U6774 (N_6774,N_3695,N_3800);
and U6775 (N_6775,N_2811,N_3628);
and U6776 (N_6776,N_3774,N_3419);
xnor U6777 (N_6777,N_4177,N_4796);
xnor U6778 (N_6778,N_4543,N_4205);
and U6779 (N_6779,N_3518,N_2605);
nor U6780 (N_6780,N_4985,N_4817);
xnor U6781 (N_6781,N_3681,N_2912);
xnor U6782 (N_6782,N_3545,N_3662);
or U6783 (N_6783,N_2634,N_3410);
nand U6784 (N_6784,N_4054,N_3008);
xnor U6785 (N_6785,N_3148,N_3678);
and U6786 (N_6786,N_4366,N_4785);
or U6787 (N_6787,N_4343,N_3428);
nand U6788 (N_6788,N_3500,N_3559);
nand U6789 (N_6789,N_4984,N_4741);
nand U6790 (N_6790,N_3805,N_4550);
nand U6791 (N_6791,N_4793,N_4977);
nor U6792 (N_6792,N_4396,N_4268);
nand U6793 (N_6793,N_3835,N_4479);
nor U6794 (N_6794,N_3361,N_4474);
and U6795 (N_6795,N_4891,N_4759);
nand U6796 (N_6796,N_2903,N_4619);
xor U6797 (N_6797,N_2628,N_2601);
nor U6798 (N_6798,N_2888,N_4712);
nor U6799 (N_6799,N_3825,N_4169);
nor U6800 (N_6800,N_2754,N_4233);
nand U6801 (N_6801,N_3679,N_3410);
or U6802 (N_6802,N_3706,N_3734);
or U6803 (N_6803,N_3622,N_3289);
and U6804 (N_6804,N_2802,N_4387);
or U6805 (N_6805,N_3862,N_3433);
or U6806 (N_6806,N_4829,N_2800);
nor U6807 (N_6807,N_2627,N_4153);
and U6808 (N_6808,N_3903,N_3512);
or U6809 (N_6809,N_3796,N_2871);
nand U6810 (N_6810,N_2773,N_3147);
or U6811 (N_6811,N_3710,N_4930);
or U6812 (N_6812,N_3462,N_4468);
and U6813 (N_6813,N_2790,N_4900);
and U6814 (N_6814,N_3120,N_3410);
nand U6815 (N_6815,N_3534,N_3689);
nand U6816 (N_6816,N_4066,N_2586);
nand U6817 (N_6817,N_3552,N_2889);
or U6818 (N_6818,N_4101,N_4011);
xnor U6819 (N_6819,N_4271,N_2507);
nor U6820 (N_6820,N_3338,N_3272);
or U6821 (N_6821,N_2656,N_2559);
and U6822 (N_6822,N_3891,N_3505);
nor U6823 (N_6823,N_3220,N_4483);
or U6824 (N_6824,N_3077,N_2835);
nand U6825 (N_6825,N_3779,N_3701);
and U6826 (N_6826,N_4843,N_4917);
and U6827 (N_6827,N_2820,N_4415);
nor U6828 (N_6828,N_4313,N_3182);
nand U6829 (N_6829,N_2630,N_2586);
nand U6830 (N_6830,N_2833,N_4133);
xor U6831 (N_6831,N_4711,N_3439);
or U6832 (N_6832,N_3032,N_3315);
nand U6833 (N_6833,N_3419,N_2517);
nor U6834 (N_6834,N_4159,N_3908);
or U6835 (N_6835,N_3579,N_4068);
and U6836 (N_6836,N_4542,N_4342);
nand U6837 (N_6837,N_4512,N_2539);
or U6838 (N_6838,N_3573,N_3195);
nor U6839 (N_6839,N_4620,N_3524);
nand U6840 (N_6840,N_3836,N_2640);
nand U6841 (N_6841,N_3741,N_4743);
nor U6842 (N_6842,N_4709,N_2601);
nand U6843 (N_6843,N_4654,N_2921);
nand U6844 (N_6844,N_4061,N_2605);
xor U6845 (N_6845,N_2827,N_4386);
xor U6846 (N_6846,N_3171,N_2965);
xnor U6847 (N_6847,N_2537,N_4101);
and U6848 (N_6848,N_4070,N_4964);
nor U6849 (N_6849,N_4883,N_4957);
nand U6850 (N_6850,N_3263,N_3218);
and U6851 (N_6851,N_4006,N_2534);
or U6852 (N_6852,N_2548,N_3110);
nor U6853 (N_6853,N_3406,N_4807);
nand U6854 (N_6854,N_3719,N_4743);
nand U6855 (N_6855,N_3063,N_4092);
and U6856 (N_6856,N_3523,N_4039);
and U6857 (N_6857,N_4467,N_4837);
nand U6858 (N_6858,N_2978,N_4927);
or U6859 (N_6859,N_3051,N_2828);
and U6860 (N_6860,N_3174,N_3894);
or U6861 (N_6861,N_4080,N_2591);
nor U6862 (N_6862,N_3011,N_4277);
nand U6863 (N_6863,N_3995,N_4065);
nand U6864 (N_6864,N_2930,N_3423);
nor U6865 (N_6865,N_3265,N_2961);
nand U6866 (N_6866,N_2813,N_3640);
nand U6867 (N_6867,N_3255,N_3616);
nor U6868 (N_6868,N_3799,N_4525);
nor U6869 (N_6869,N_3490,N_2681);
or U6870 (N_6870,N_3007,N_3238);
and U6871 (N_6871,N_4134,N_3745);
or U6872 (N_6872,N_3577,N_4906);
nand U6873 (N_6873,N_3362,N_2896);
nand U6874 (N_6874,N_2995,N_3303);
or U6875 (N_6875,N_4301,N_4256);
nand U6876 (N_6876,N_4967,N_2898);
nor U6877 (N_6877,N_2513,N_3916);
nand U6878 (N_6878,N_4830,N_3002);
and U6879 (N_6879,N_3377,N_2577);
nor U6880 (N_6880,N_4895,N_4338);
or U6881 (N_6881,N_4870,N_4355);
and U6882 (N_6882,N_3835,N_2680);
or U6883 (N_6883,N_3787,N_4160);
and U6884 (N_6884,N_3941,N_3034);
and U6885 (N_6885,N_4069,N_4953);
nor U6886 (N_6886,N_2947,N_3210);
or U6887 (N_6887,N_3636,N_3056);
xor U6888 (N_6888,N_3163,N_3396);
nand U6889 (N_6889,N_2717,N_4503);
or U6890 (N_6890,N_3181,N_4248);
nor U6891 (N_6891,N_2689,N_3393);
nor U6892 (N_6892,N_3648,N_3846);
and U6893 (N_6893,N_3099,N_3602);
and U6894 (N_6894,N_4366,N_4045);
nand U6895 (N_6895,N_4742,N_2913);
xor U6896 (N_6896,N_4978,N_4933);
or U6897 (N_6897,N_4546,N_3283);
nor U6898 (N_6898,N_4202,N_3227);
or U6899 (N_6899,N_3538,N_3403);
nor U6900 (N_6900,N_3485,N_3107);
and U6901 (N_6901,N_3430,N_3096);
nor U6902 (N_6902,N_3393,N_3781);
and U6903 (N_6903,N_4343,N_3699);
or U6904 (N_6904,N_4740,N_3262);
or U6905 (N_6905,N_2825,N_3690);
nor U6906 (N_6906,N_4169,N_3385);
xor U6907 (N_6907,N_3211,N_4400);
nor U6908 (N_6908,N_4265,N_3172);
and U6909 (N_6909,N_2575,N_4700);
or U6910 (N_6910,N_2793,N_4663);
nand U6911 (N_6911,N_4387,N_3554);
or U6912 (N_6912,N_4471,N_4668);
nand U6913 (N_6913,N_4180,N_3202);
nor U6914 (N_6914,N_3870,N_4683);
or U6915 (N_6915,N_4578,N_4832);
or U6916 (N_6916,N_4369,N_3960);
nor U6917 (N_6917,N_4093,N_2851);
nand U6918 (N_6918,N_3397,N_2592);
nor U6919 (N_6919,N_4974,N_3633);
nor U6920 (N_6920,N_4209,N_3943);
and U6921 (N_6921,N_2998,N_4347);
or U6922 (N_6922,N_2867,N_4197);
and U6923 (N_6923,N_2932,N_3165);
or U6924 (N_6924,N_4315,N_4110);
and U6925 (N_6925,N_2666,N_3232);
nor U6926 (N_6926,N_4047,N_4277);
or U6927 (N_6927,N_4313,N_3181);
xnor U6928 (N_6928,N_3235,N_4269);
nand U6929 (N_6929,N_3325,N_4866);
and U6930 (N_6930,N_4300,N_4577);
nor U6931 (N_6931,N_3793,N_4820);
or U6932 (N_6932,N_4320,N_3678);
nor U6933 (N_6933,N_4896,N_3890);
nor U6934 (N_6934,N_4653,N_3987);
or U6935 (N_6935,N_3452,N_4737);
and U6936 (N_6936,N_2857,N_4599);
nand U6937 (N_6937,N_3733,N_3906);
nor U6938 (N_6938,N_2788,N_2611);
nor U6939 (N_6939,N_3814,N_2691);
nand U6940 (N_6940,N_4412,N_3796);
or U6941 (N_6941,N_3941,N_3235);
nand U6942 (N_6942,N_4558,N_3372);
nand U6943 (N_6943,N_4683,N_3597);
and U6944 (N_6944,N_4673,N_3954);
xor U6945 (N_6945,N_4648,N_4468);
or U6946 (N_6946,N_3093,N_3782);
or U6947 (N_6947,N_4081,N_3003);
nand U6948 (N_6948,N_3609,N_2653);
and U6949 (N_6949,N_4303,N_2696);
or U6950 (N_6950,N_4205,N_4078);
nor U6951 (N_6951,N_2516,N_3747);
and U6952 (N_6952,N_2547,N_3747);
or U6953 (N_6953,N_3754,N_2834);
or U6954 (N_6954,N_2897,N_3840);
and U6955 (N_6955,N_4897,N_3346);
and U6956 (N_6956,N_3447,N_4284);
and U6957 (N_6957,N_4525,N_2526);
or U6958 (N_6958,N_3172,N_3022);
and U6959 (N_6959,N_4767,N_3940);
nor U6960 (N_6960,N_4721,N_3412);
nor U6961 (N_6961,N_3075,N_4602);
nand U6962 (N_6962,N_4285,N_3420);
and U6963 (N_6963,N_3912,N_4388);
nor U6964 (N_6964,N_2509,N_2877);
or U6965 (N_6965,N_3647,N_4560);
nand U6966 (N_6966,N_3676,N_2848);
or U6967 (N_6967,N_4826,N_3970);
nand U6968 (N_6968,N_3076,N_3358);
nand U6969 (N_6969,N_3055,N_4791);
nor U6970 (N_6970,N_4678,N_4374);
nand U6971 (N_6971,N_2681,N_3496);
and U6972 (N_6972,N_3313,N_2925);
or U6973 (N_6973,N_4127,N_3887);
nor U6974 (N_6974,N_3143,N_3031);
nand U6975 (N_6975,N_3608,N_3196);
nor U6976 (N_6976,N_2886,N_3580);
or U6977 (N_6977,N_3086,N_4171);
and U6978 (N_6978,N_4928,N_3074);
or U6979 (N_6979,N_2935,N_2834);
and U6980 (N_6980,N_2944,N_3389);
nor U6981 (N_6981,N_4303,N_2968);
nand U6982 (N_6982,N_3756,N_4292);
and U6983 (N_6983,N_4733,N_3750);
nor U6984 (N_6984,N_3488,N_4683);
nor U6985 (N_6985,N_3373,N_3531);
nor U6986 (N_6986,N_4438,N_4909);
or U6987 (N_6987,N_3108,N_4626);
nand U6988 (N_6988,N_2707,N_4459);
and U6989 (N_6989,N_3515,N_3421);
nor U6990 (N_6990,N_2852,N_4141);
xnor U6991 (N_6991,N_4830,N_3329);
nand U6992 (N_6992,N_3204,N_3084);
or U6993 (N_6993,N_3314,N_3545);
or U6994 (N_6994,N_4451,N_3938);
and U6995 (N_6995,N_3898,N_4225);
or U6996 (N_6996,N_3392,N_4058);
or U6997 (N_6997,N_3518,N_3534);
or U6998 (N_6998,N_2583,N_3408);
xnor U6999 (N_6999,N_3057,N_2627);
and U7000 (N_7000,N_3944,N_4933);
nor U7001 (N_7001,N_3926,N_2992);
and U7002 (N_7002,N_3374,N_2887);
nand U7003 (N_7003,N_3193,N_4940);
or U7004 (N_7004,N_4608,N_4958);
and U7005 (N_7005,N_2651,N_2545);
or U7006 (N_7006,N_3567,N_3128);
or U7007 (N_7007,N_3690,N_4735);
or U7008 (N_7008,N_3524,N_4271);
and U7009 (N_7009,N_4113,N_4980);
xnor U7010 (N_7010,N_4858,N_4268);
nor U7011 (N_7011,N_3527,N_4048);
or U7012 (N_7012,N_4812,N_3021);
xor U7013 (N_7013,N_2697,N_3702);
xor U7014 (N_7014,N_4486,N_3968);
xor U7015 (N_7015,N_4620,N_3628);
and U7016 (N_7016,N_3589,N_2607);
or U7017 (N_7017,N_3415,N_4206);
nor U7018 (N_7018,N_3174,N_3321);
or U7019 (N_7019,N_3985,N_4955);
nand U7020 (N_7020,N_4734,N_3775);
nand U7021 (N_7021,N_3820,N_3859);
nand U7022 (N_7022,N_4497,N_4416);
nor U7023 (N_7023,N_2909,N_4015);
or U7024 (N_7024,N_4338,N_3143);
and U7025 (N_7025,N_3949,N_4773);
and U7026 (N_7026,N_3734,N_3256);
nand U7027 (N_7027,N_4958,N_2729);
or U7028 (N_7028,N_4943,N_3522);
nor U7029 (N_7029,N_3983,N_3380);
nor U7030 (N_7030,N_4334,N_2892);
or U7031 (N_7031,N_3014,N_4402);
xnor U7032 (N_7032,N_4789,N_4350);
xnor U7033 (N_7033,N_3008,N_3409);
xnor U7034 (N_7034,N_4035,N_3614);
or U7035 (N_7035,N_4253,N_3156);
or U7036 (N_7036,N_3160,N_3444);
nand U7037 (N_7037,N_4443,N_3736);
nand U7038 (N_7038,N_2902,N_2575);
xor U7039 (N_7039,N_3558,N_4208);
nor U7040 (N_7040,N_2543,N_4973);
or U7041 (N_7041,N_2724,N_4467);
and U7042 (N_7042,N_2971,N_3385);
and U7043 (N_7043,N_4079,N_4257);
xnor U7044 (N_7044,N_3005,N_2871);
nor U7045 (N_7045,N_4173,N_3671);
xor U7046 (N_7046,N_2923,N_2552);
and U7047 (N_7047,N_4200,N_3156);
nor U7048 (N_7048,N_3434,N_2636);
xnor U7049 (N_7049,N_2861,N_2983);
and U7050 (N_7050,N_2616,N_2533);
nand U7051 (N_7051,N_3413,N_2825);
and U7052 (N_7052,N_3028,N_3634);
and U7053 (N_7053,N_3028,N_3598);
nand U7054 (N_7054,N_2853,N_3660);
nor U7055 (N_7055,N_2607,N_4701);
nor U7056 (N_7056,N_3122,N_4590);
and U7057 (N_7057,N_4994,N_3392);
nor U7058 (N_7058,N_2778,N_2767);
and U7059 (N_7059,N_3990,N_4425);
nor U7060 (N_7060,N_2765,N_4188);
and U7061 (N_7061,N_3139,N_3470);
nand U7062 (N_7062,N_3775,N_4177);
nor U7063 (N_7063,N_4908,N_3027);
or U7064 (N_7064,N_3862,N_3268);
or U7065 (N_7065,N_3010,N_3244);
nor U7066 (N_7066,N_4781,N_3595);
nand U7067 (N_7067,N_3451,N_3899);
and U7068 (N_7068,N_4693,N_2508);
or U7069 (N_7069,N_4207,N_2981);
xor U7070 (N_7070,N_4342,N_2727);
or U7071 (N_7071,N_4367,N_3203);
or U7072 (N_7072,N_3015,N_2748);
or U7073 (N_7073,N_2671,N_4387);
xor U7074 (N_7074,N_4132,N_3412);
nor U7075 (N_7075,N_4238,N_3108);
or U7076 (N_7076,N_3617,N_3891);
nor U7077 (N_7077,N_4506,N_4853);
or U7078 (N_7078,N_2573,N_2957);
or U7079 (N_7079,N_4159,N_4300);
or U7080 (N_7080,N_2566,N_4047);
or U7081 (N_7081,N_2928,N_4828);
nor U7082 (N_7082,N_4980,N_4566);
nor U7083 (N_7083,N_4495,N_4144);
and U7084 (N_7084,N_2946,N_4260);
and U7085 (N_7085,N_2568,N_3864);
or U7086 (N_7086,N_3605,N_4013);
and U7087 (N_7087,N_3532,N_3551);
nand U7088 (N_7088,N_3600,N_2749);
or U7089 (N_7089,N_3782,N_3271);
nor U7090 (N_7090,N_4058,N_3169);
nand U7091 (N_7091,N_4333,N_4726);
and U7092 (N_7092,N_4540,N_3730);
nand U7093 (N_7093,N_3692,N_3346);
xor U7094 (N_7094,N_3750,N_3708);
xor U7095 (N_7095,N_4926,N_3899);
nor U7096 (N_7096,N_2911,N_4217);
nor U7097 (N_7097,N_3990,N_2522);
or U7098 (N_7098,N_4012,N_3071);
nor U7099 (N_7099,N_3608,N_3118);
or U7100 (N_7100,N_3298,N_3168);
nand U7101 (N_7101,N_2934,N_3364);
and U7102 (N_7102,N_4916,N_3651);
nand U7103 (N_7103,N_3148,N_2648);
nand U7104 (N_7104,N_3099,N_2686);
nor U7105 (N_7105,N_3162,N_2760);
and U7106 (N_7106,N_2959,N_4823);
nor U7107 (N_7107,N_3542,N_3006);
and U7108 (N_7108,N_3221,N_3601);
nand U7109 (N_7109,N_3677,N_2765);
and U7110 (N_7110,N_2979,N_2855);
and U7111 (N_7111,N_3306,N_4781);
and U7112 (N_7112,N_3846,N_4844);
and U7113 (N_7113,N_4957,N_2673);
and U7114 (N_7114,N_2563,N_3362);
nand U7115 (N_7115,N_3626,N_4481);
nor U7116 (N_7116,N_2741,N_3109);
and U7117 (N_7117,N_4032,N_4696);
and U7118 (N_7118,N_3267,N_3036);
nor U7119 (N_7119,N_4792,N_3787);
nor U7120 (N_7120,N_3845,N_4379);
nand U7121 (N_7121,N_3755,N_3783);
and U7122 (N_7122,N_3809,N_3026);
and U7123 (N_7123,N_4854,N_3821);
nand U7124 (N_7124,N_4044,N_4536);
xnor U7125 (N_7125,N_3215,N_3538);
nand U7126 (N_7126,N_4932,N_4999);
or U7127 (N_7127,N_3854,N_3583);
xnor U7128 (N_7128,N_3022,N_4523);
and U7129 (N_7129,N_4303,N_2758);
or U7130 (N_7130,N_2524,N_3148);
nor U7131 (N_7131,N_4480,N_3105);
xor U7132 (N_7132,N_3299,N_3347);
nor U7133 (N_7133,N_4327,N_4113);
and U7134 (N_7134,N_3324,N_3226);
nand U7135 (N_7135,N_3537,N_2826);
and U7136 (N_7136,N_2587,N_2766);
nand U7137 (N_7137,N_4137,N_2597);
and U7138 (N_7138,N_2550,N_3671);
or U7139 (N_7139,N_2596,N_2890);
or U7140 (N_7140,N_3984,N_3326);
and U7141 (N_7141,N_4744,N_2709);
nor U7142 (N_7142,N_4366,N_2570);
or U7143 (N_7143,N_4998,N_4937);
nand U7144 (N_7144,N_4152,N_3553);
xnor U7145 (N_7145,N_3845,N_3606);
nor U7146 (N_7146,N_3627,N_3385);
or U7147 (N_7147,N_2536,N_2818);
or U7148 (N_7148,N_3479,N_4551);
nand U7149 (N_7149,N_3971,N_3325);
nor U7150 (N_7150,N_3571,N_4911);
nand U7151 (N_7151,N_4722,N_4274);
xnor U7152 (N_7152,N_3442,N_4596);
nand U7153 (N_7153,N_4586,N_2703);
or U7154 (N_7154,N_4349,N_4666);
nor U7155 (N_7155,N_4792,N_4100);
xor U7156 (N_7156,N_3540,N_2517);
nor U7157 (N_7157,N_4003,N_4554);
or U7158 (N_7158,N_4780,N_4960);
nor U7159 (N_7159,N_4158,N_2881);
nand U7160 (N_7160,N_4151,N_3253);
nor U7161 (N_7161,N_3987,N_2935);
xnor U7162 (N_7162,N_2971,N_3108);
nand U7163 (N_7163,N_3658,N_4304);
or U7164 (N_7164,N_2813,N_3628);
nand U7165 (N_7165,N_3152,N_3902);
or U7166 (N_7166,N_2911,N_4349);
or U7167 (N_7167,N_4889,N_2562);
and U7168 (N_7168,N_4836,N_2855);
xor U7169 (N_7169,N_4953,N_2690);
nor U7170 (N_7170,N_4586,N_3573);
nor U7171 (N_7171,N_4125,N_3316);
nor U7172 (N_7172,N_2771,N_3964);
nor U7173 (N_7173,N_2967,N_4863);
nand U7174 (N_7174,N_3194,N_4572);
xnor U7175 (N_7175,N_4501,N_4168);
or U7176 (N_7176,N_3854,N_3807);
nand U7177 (N_7177,N_3145,N_2544);
and U7178 (N_7178,N_4838,N_2900);
or U7179 (N_7179,N_2940,N_3993);
and U7180 (N_7180,N_3174,N_3448);
and U7181 (N_7181,N_2507,N_3794);
nand U7182 (N_7182,N_3369,N_3404);
nand U7183 (N_7183,N_4927,N_3952);
and U7184 (N_7184,N_4788,N_4236);
xor U7185 (N_7185,N_4391,N_3140);
or U7186 (N_7186,N_4993,N_4092);
or U7187 (N_7187,N_3107,N_3826);
or U7188 (N_7188,N_3629,N_2603);
or U7189 (N_7189,N_4733,N_3914);
and U7190 (N_7190,N_2519,N_4535);
nand U7191 (N_7191,N_4209,N_3508);
xor U7192 (N_7192,N_4944,N_3306);
nand U7193 (N_7193,N_4259,N_4844);
nand U7194 (N_7194,N_4736,N_3889);
nand U7195 (N_7195,N_3491,N_3680);
nor U7196 (N_7196,N_4725,N_4042);
or U7197 (N_7197,N_2668,N_2823);
or U7198 (N_7198,N_4548,N_4436);
and U7199 (N_7199,N_3509,N_4055);
and U7200 (N_7200,N_2909,N_3753);
nor U7201 (N_7201,N_3183,N_4208);
nor U7202 (N_7202,N_4025,N_3683);
nand U7203 (N_7203,N_4437,N_3004);
nand U7204 (N_7204,N_4917,N_2713);
or U7205 (N_7205,N_4240,N_3254);
nand U7206 (N_7206,N_2605,N_4899);
nor U7207 (N_7207,N_3289,N_4719);
xor U7208 (N_7208,N_3068,N_4372);
nor U7209 (N_7209,N_4809,N_4452);
nor U7210 (N_7210,N_3881,N_2856);
and U7211 (N_7211,N_4217,N_3286);
or U7212 (N_7212,N_3324,N_3649);
and U7213 (N_7213,N_4809,N_4906);
nor U7214 (N_7214,N_3759,N_2894);
nor U7215 (N_7215,N_4312,N_3799);
nor U7216 (N_7216,N_2782,N_3456);
or U7217 (N_7217,N_4490,N_3555);
and U7218 (N_7218,N_3067,N_2787);
and U7219 (N_7219,N_4173,N_4972);
nor U7220 (N_7220,N_3441,N_4900);
or U7221 (N_7221,N_4291,N_2636);
nand U7222 (N_7222,N_4274,N_2715);
nor U7223 (N_7223,N_3400,N_2704);
and U7224 (N_7224,N_4070,N_4230);
nand U7225 (N_7225,N_3988,N_4812);
nor U7226 (N_7226,N_2880,N_2987);
nor U7227 (N_7227,N_3841,N_2764);
nor U7228 (N_7228,N_4828,N_4183);
xor U7229 (N_7229,N_2689,N_4742);
nand U7230 (N_7230,N_2842,N_3424);
and U7231 (N_7231,N_3940,N_3227);
xor U7232 (N_7232,N_3514,N_3320);
and U7233 (N_7233,N_3346,N_4383);
or U7234 (N_7234,N_3062,N_4055);
or U7235 (N_7235,N_4871,N_3760);
xor U7236 (N_7236,N_3944,N_3423);
nor U7237 (N_7237,N_3215,N_4135);
nor U7238 (N_7238,N_3696,N_2706);
nand U7239 (N_7239,N_4158,N_3351);
or U7240 (N_7240,N_4818,N_3027);
and U7241 (N_7241,N_3376,N_3296);
or U7242 (N_7242,N_4833,N_2637);
nor U7243 (N_7243,N_3230,N_3516);
or U7244 (N_7244,N_3194,N_4637);
or U7245 (N_7245,N_3459,N_3779);
nor U7246 (N_7246,N_3234,N_4498);
and U7247 (N_7247,N_4267,N_3555);
xnor U7248 (N_7248,N_4092,N_4652);
xnor U7249 (N_7249,N_3928,N_2539);
or U7250 (N_7250,N_4679,N_3927);
nor U7251 (N_7251,N_2793,N_4844);
xor U7252 (N_7252,N_4229,N_2788);
and U7253 (N_7253,N_3841,N_3570);
or U7254 (N_7254,N_3647,N_4353);
xnor U7255 (N_7255,N_3516,N_3953);
and U7256 (N_7256,N_3332,N_4817);
or U7257 (N_7257,N_2966,N_3056);
nand U7258 (N_7258,N_3694,N_3262);
nand U7259 (N_7259,N_3330,N_4659);
xor U7260 (N_7260,N_4711,N_3378);
and U7261 (N_7261,N_4717,N_3704);
or U7262 (N_7262,N_3708,N_3702);
or U7263 (N_7263,N_3492,N_4977);
nand U7264 (N_7264,N_4656,N_2685);
xnor U7265 (N_7265,N_4848,N_2975);
or U7266 (N_7266,N_2800,N_3116);
nand U7267 (N_7267,N_4091,N_4586);
nor U7268 (N_7268,N_4888,N_4132);
and U7269 (N_7269,N_2639,N_3193);
and U7270 (N_7270,N_3922,N_2823);
nand U7271 (N_7271,N_4717,N_4565);
xnor U7272 (N_7272,N_2890,N_3388);
nand U7273 (N_7273,N_4072,N_2905);
nand U7274 (N_7274,N_3888,N_4364);
nor U7275 (N_7275,N_2751,N_3209);
xnor U7276 (N_7276,N_3810,N_4918);
and U7277 (N_7277,N_4300,N_4108);
or U7278 (N_7278,N_4814,N_4043);
and U7279 (N_7279,N_4420,N_4211);
or U7280 (N_7280,N_4806,N_3829);
and U7281 (N_7281,N_3603,N_2610);
nand U7282 (N_7282,N_4365,N_4198);
or U7283 (N_7283,N_2845,N_2936);
and U7284 (N_7284,N_4216,N_3429);
and U7285 (N_7285,N_3971,N_2677);
and U7286 (N_7286,N_3576,N_4944);
and U7287 (N_7287,N_3793,N_2520);
or U7288 (N_7288,N_4732,N_3846);
nand U7289 (N_7289,N_3688,N_3256);
nand U7290 (N_7290,N_2960,N_4587);
or U7291 (N_7291,N_3998,N_3865);
xor U7292 (N_7292,N_4670,N_3099);
nand U7293 (N_7293,N_4475,N_2996);
or U7294 (N_7294,N_3770,N_2628);
xor U7295 (N_7295,N_2916,N_4954);
nor U7296 (N_7296,N_3350,N_2804);
nor U7297 (N_7297,N_3967,N_3361);
or U7298 (N_7298,N_2912,N_4166);
and U7299 (N_7299,N_2768,N_4687);
nor U7300 (N_7300,N_2557,N_2607);
nor U7301 (N_7301,N_4635,N_3031);
nor U7302 (N_7302,N_3800,N_2647);
xnor U7303 (N_7303,N_2884,N_4523);
nand U7304 (N_7304,N_2532,N_3311);
nor U7305 (N_7305,N_3114,N_4438);
or U7306 (N_7306,N_4180,N_4580);
xnor U7307 (N_7307,N_2832,N_4751);
xnor U7308 (N_7308,N_4791,N_4348);
and U7309 (N_7309,N_4110,N_4175);
and U7310 (N_7310,N_4013,N_3631);
nor U7311 (N_7311,N_2942,N_3242);
or U7312 (N_7312,N_3397,N_3393);
and U7313 (N_7313,N_4678,N_2810);
and U7314 (N_7314,N_3737,N_3567);
or U7315 (N_7315,N_3314,N_3430);
and U7316 (N_7316,N_2725,N_3585);
nand U7317 (N_7317,N_3943,N_4228);
and U7318 (N_7318,N_3356,N_4649);
nor U7319 (N_7319,N_4508,N_4100);
and U7320 (N_7320,N_3604,N_3778);
nand U7321 (N_7321,N_4341,N_4768);
and U7322 (N_7322,N_3295,N_3519);
nand U7323 (N_7323,N_3917,N_4040);
xor U7324 (N_7324,N_2606,N_2522);
xor U7325 (N_7325,N_4727,N_3290);
or U7326 (N_7326,N_4471,N_3944);
nand U7327 (N_7327,N_2703,N_4287);
nor U7328 (N_7328,N_3485,N_3938);
or U7329 (N_7329,N_2981,N_2899);
nand U7330 (N_7330,N_3857,N_4857);
nand U7331 (N_7331,N_4590,N_3676);
or U7332 (N_7332,N_3976,N_3255);
nor U7333 (N_7333,N_4260,N_3278);
nand U7334 (N_7334,N_3412,N_4030);
nor U7335 (N_7335,N_2677,N_3351);
and U7336 (N_7336,N_4639,N_2644);
or U7337 (N_7337,N_4168,N_4975);
nand U7338 (N_7338,N_3600,N_3533);
nand U7339 (N_7339,N_3591,N_2973);
and U7340 (N_7340,N_2867,N_2653);
nor U7341 (N_7341,N_4817,N_4279);
nor U7342 (N_7342,N_3783,N_4330);
nand U7343 (N_7343,N_4633,N_2776);
xor U7344 (N_7344,N_4214,N_4582);
xor U7345 (N_7345,N_3390,N_2995);
and U7346 (N_7346,N_4045,N_4563);
and U7347 (N_7347,N_3531,N_4994);
and U7348 (N_7348,N_4905,N_3101);
nor U7349 (N_7349,N_3808,N_4203);
or U7350 (N_7350,N_3266,N_4178);
xnor U7351 (N_7351,N_3878,N_4359);
nand U7352 (N_7352,N_3000,N_3538);
nand U7353 (N_7353,N_2903,N_3140);
nor U7354 (N_7354,N_3633,N_4068);
nor U7355 (N_7355,N_2654,N_4799);
nor U7356 (N_7356,N_2660,N_4417);
nand U7357 (N_7357,N_3685,N_3711);
xnor U7358 (N_7358,N_4629,N_3467);
nor U7359 (N_7359,N_4598,N_4184);
or U7360 (N_7360,N_4281,N_4289);
or U7361 (N_7361,N_3975,N_4017);
or U7362 (N_7362,N_4283,N_3688);
nand U7363 (N_7363,N_3838,N_3359);
nand U7364 (N_7364,N_4905,N_2651);
nand U7365 (N_7365,N_4099,N_3038);
nand U7366 (N_7366,N_2963,N_4460);
or U7367 (N_7367,N_4671,N_3920);
or U7368 (N_7368,N_2537,N_4439);
or U7369 (N_7369,N_3719,N_2876);
or U7370 (N_7370,N_4733,N_4391);
nand U7371 (N_7371,N_3121,N_4410);
nand U7372 (N_7372,N_3392,N_2651);
and U7373 (N_7373,N_3244,N_3691);
xor U7374 (N_7374,N_2662,N_3918);
xnor U7375 (N_7375,N_2912,N_4009);
nand U7376 (N_7376,N_3008,N_3054);
and U7377 (N_7377,N_2522,N_3826);
nand U7378 (N_7378,N_3716,N_4612);
nand U7379 (N_7379,N_3302,N_2979);
xor U7380 (N_7380,N_4841,N_2832);
or U7381 (N_7381,N_3818,N_3605);
and U7382 (N_7382,N_2977,N_3275);
nor U7383 (N_7383,N_3940,N_3865);
or U7384 (N_7384,N_2875,N_4880);
nand U7385 (N_7385,N_3300,N_4376);
nor U7386 (N_7386,N_4797,N_4644);
xor U7387 (N_7387,N_3650,N_3390);
nor U7388 (N_7388,N_3498,N_4902);
and U7389 (N_7389,N_4111,N_4512);
nor U7390 (N_7390,N_4065,N_2698);
nand U7391 (N_7391,N_3237,N_4259);
or U7392 (N_7392,N_3374,N_3027);
xor U7393 (N_7393,N_4066,N_4179);
or U7394 (N_7394,N_4160,N_3352);
nor U7395 (N_7395,N_4225,N_3973);
and U7396 (N_7396,N_4310,N_4723);
or U7397 (N_7397,N_4523,N_3268);
or U7398 (N_7398,N_2710,N_2505);
xor U7399 (N_7399,N_4651,N_4593);
nor U7400 (N_7400,N_3427,N_3361);
nor U7401 (N_7401,N_3695,N_3821);
nor U7402 (N_7402,N_2660,N_3801);
and U7403 (N_7403,N_4866,N_4788);
nor U7404 (N_7404,N_4121,N_2708);
nor U7405 (N_7405,N_4678,N_3007);
xor U7406 (N_7406,N_4741,N_2756);
or U7407 (N_7407,N_4678,N_4950);
or U7408 (N_7408,N_4339,N_2615);
or U7409 (N_7409,N_4734,N_4752);
nand U7410 (N_7410,N_4748,N_4337);
nor U7411 (N_7411,N_3663,N_3103);
or U7412 (N_7412,N_3224,N_2584);
or U7413 (N_7413,N_2586,N_3030);
and U7414 (N_7414,N_4523,N_3535);
or U7415 (N_7415,N_3898,N_3660);
and U7416 (N_7416,N_4967,N_3425);
and U7417 (N_7417,N_3190,N_3135);
or U7418 (N_7418,N_2818,N_4620);
nand U7419 (N_7419,N_2899,N_3791);
nor U7420 (N_7420,N_4454,N_4602);
xor U7421 (N_7421,N_3754,N_3518);
and U7422 (N_7422,N_4038,N_3686);
nand U7423 (N_7423,N_3319,N_3533);
nor U7424 (N_7424,N_3103,N_2577);
and U7425 (N_7425,N_3156,N_2914);
or U7426 (N_7426,N_4974,N_3178);
and U7427 (N_7427,N_4121,N_3444);
or U7428 (N_7428,N_4798,N_2633);
and U7429 (N_7429,N_4810,N_2942);
nand U7430 (N_7430,N_3097,N_3752);
xnor U7431 (N_7431,N_3285,N_4275);
xor U7432 (N_7432,N_4732,N_3146);
nand U7433 (N_7433,N_4068,N_3211);
nand U7434 (N_7434,N_3906,N_3177);
and U7435 (N_7435,N_4477,N_4715);
and U7436 (N_7436,N_3173,N_3904);
and U7437 (N_7437,N_3083,N_4248);
and U7438 (N_7438,N_4949,N_4986);
nor U7439 (N_7439,N_2908,N_4679);
or U7440 (N_7440,N_4003,N_3700);
and U7441 (N_7441,N_3890,N_3188);
and U7442 (N_7442,N_3991,N_2643);
nand U7443 (N_7443,N_3348,N_4689);
nand U7444 (N_7444,N_4362,N_3253);
nand U7445 (N_7445,N_2565,N_4842);
or U7446 (N_7446,N_3446,N_3832);
and U7447 (N_7447,N_3160,N_4357);
and U7448 (N_7448,N_3797,N_2700);
and U7449 (N_7449,N_3137,N_4456);
or U7450 (N_7450,N_3704,N_3195);
xor U7451 (N_7451,N_4137,N_3753);
or U7452 (N_7452,N_4884,N_3059);
and U7453 (N_7453,N_3244,N_4086);
nor U7454 (N_7454,N_3024,N_4370);
or U7455 (N_7455,N_4559,N_4960);
nor U7456 (N_7456,N_4644,N_4361);
nor U7457 (N_7457,N_3569,N_3520);
nand U7458 (N_7458,N_3748,N_4317);
nand U7459 (N_7459,N_2855,N_4584);
and U7460 (N_7460,N_3049,N_4115);
nor U7461 (N_7461,N_2719,N_3391);
and U7462 (N_7462,N_4304,N_4224);
xnor U7463 (N_7463,N_4519,N_3573);
nand U7464 (N_7464,N_4920,N_2824);
and U7465 (N_7465,N_4460,N_3969);
nand U7466 (N_7466,N_4061,N_3558);
and U7467 (N_7467,N_2960,N_2691);
and U7468 (N_7468,N_3285,N_4094);
or U7469 (N_7469,N_3543,N_3277);
nor U7470 (N_7470,N_3437,N_3388);
or U7471 (N_7471,N_3848,N_4723);
xor U7472 (N_7472,N_4460,N_4057);
and U7473 (N_7473,N_4527,N_3763);
or U7474 (N_7474,N_3608,N_4758);
or U7475 (N_7475,N_3960,N_3963);
or U7476 (N_7476,N_2786,N_2813);
nand U7477 (N_7477,N_3228,N_3805);
xor U7478 (N_7478,N_3437,N_3871);
and U7479 (N_7479,N_2552,N_3207);
nand U7480 (N_7480,N_3787,N_2960);
nand U7481 (N_7481,N_4769,N_3288);
and U7482 (N_7482,N_3304,N_3393);
and U7483 (N_7483,N_3721,N_4912);
nand U7484 (N_7484,N_3347,N_4122);
xnor U7485 (N_7485,N_4337,N_2515);
nand U7486 (N_7486,N_3403,N_4262);
nor U7487 (N_7487,N_4537,N_4966);
and U7488 (N_7488,N_3065,N_3841);
nand U7489 (N_7489,N_4830,N_3179);
nor U7490 (N_7490,N_2949,N_4049);
and U7491 (N_7491,N_4522,N_4570);
nand U7492 (N_7492,N_3165,N_4368);
nor U7493 (N_7493,N_3823,N_3442);
nor U7494 (N_7494,N_3693,N_3603);
xnor U7495 (N_7495,N_4316,N_3855);
xor U7496 (N_7496,N_2930,N_4839);
and U7497 (N_7497,N_4501,N_3486);
nand U7498 (N_7498,N_3393,N_2589);
nor U7499 (N_7499,N_2717,N_4942);
nor U7500 (N_7500,N_7432,N_5011);
nor U7501 (N_7501,N_6302,N_6733);
and U7502 (N_7502,N_5898,N_7103);
and U7503 (N_7503,N_7008,N_5467);
nor U7504 (N_7504,N_5888,N_6319);
nand U7505 (N_7505,N_5503,N_5872);
nor U7506 (N_7506,N_6178,N_6249);
nand U7507 (N_7507,N_6150,N_6274);
and U7508 (N_7508,N_6576,N_5222);
or U7509 (N_7509,N_6650,N_5165);
and U7510 (N_7510,N_6663,N_5370);
nand U7511 (N_7511,N_5936,N_6024);
nor U7512 (N_7512,N_6337,N_5951);
nand U7513 (N_7513,N_5233,N_5306);
and U7514 (N_7514,N_7063,N_5963);
and U7515 (N_7515,N_6635,N_5982);
and U7516 (N_7516,N_6995,N_5482);
nand U7517 (N_7517,N_5298,N_6193);
nand U7518 (N_7518,N_6767,N_6124);
and U7519 (N_7519,N_5088,N_6043);
nor U7520 (N_7520,N_5847,N_5707);
xnor U7521 (N_7521,N_7411,N_5236);
nor U7522 (N_7522,N_6952,N_5556);
nand U7523 (N_7523,N_5713,N_7175);
nor U7524 (N_7524,N_7195,N_6180);
nand U7525 (N_7525,N_6657,N_5302);
or U7526 (N_7526,N_6745,N_5044);
nor U7527 (N_7527,N_5020,N_7304);
xor U7528 (N_7528,N_6688,N_5309);
xor U7529 (N_7529,N_6342,N_5822);
nand U7530 (N_7530,N_5369,N_5228);
xor U7531 (N_7531,N_5993,N_6002);
nor U7532 (N_7532,N_7346,N_6447);
nor U7533 (N_7533,N_6777,N_6729);
or U7534 (N_7534,N_5667,N_6452);
and U7535 (N_7535,N_5381,N_5045);
nor U7536 (N_7536,N_5288,N_6738);
and U7537 (N_7537,N_7424,N_5489);
nor U7538 (N_7538,N_6838,N_7107);
and U7539 (N_7539,N_5386,N_6308);
nand U7540 (N_7540,N_6255,N_6503);
and U7541 (N_7541,N_6469,N_6485);
or U7542 (N_7542,N_6393,N_6106);
nand U7543 (N_7543,N_5411,N_6779);
and U7544 (N_7544,N_7287,N_7388);
nor U7545 (N_7545,N_5692,N_5462);
or U7546 (N_7546,N_7119,N_5798);
and U7547 (N_7547,N_5238,N_5647);
and U7548 (N_7548,N_6913,N_6912);
nand U7549 (N_7549,N_5785,N_6459);
nor U7550 (N_7550,N_5491,N_7430);
and U7551 (N_7551,N_6118,N_5094);
or U7552 (N_7552,N_7339,N_7193);
or U7553 (N_7553,N_6895,N_7487);
and U7554 (N_7554,N_6800,N_7074);
nand U7555 (N_7555,N_6722,N_6453);
nand U7556 (N_7556,N_7456,N_6827);
or U7557 (N_7557,N_5379,N_5634);
nor U7558 (N_7558,N_5355,N_6048);
nand U7559 (N_7559,N_6202,N_5835);
nor U7560 (N_7560,N_5345,N_7344);
xor U7561 (N_7561,N_6347,N_5916);
or U7562 (N_7562,N_6539,N_6637);
and U7563 (N_7563,N_7232,N_6338);
nor U7564 (N_7564,N_5706,N_5552);
xnor U7565 (N_7565,N_7222,N_5065);
and U7566 (N_7566,N_6102,N_7459);
or U7567 (N_7567,N_5112,N_6015);
nor U7568 (N_7568,N_7375,N_6289);
or U7569 (N_7569,N_5249,N_6413);
or U7570 (N_7570,N_6051,N_6488);
nor U7571 (N_7571,N_6534,N_6837);
nor U7572 (N_7572,N_7147,N_5476);
nor U7573 (N_7573,N_7178,N_5547);
and U7574 (N_7574,N_5447,N_7039);
and U7575 (N_7575,N_6325,N_6680);
nor U7576 (N_7576,N_5277,N_5725);
nand U7577 (N_7577,N_7386,N_6335);
or U7578 (N_7578,N_7099,N_6173);
nor U7579 (N_7579,N_5892,N_7263);
and U7580 (N_7580,N_5002,N_5864);
nand U7581 (N_7581,N_6559,N_6731);
or U7582 (N_7582,N_7405,N_6125);
nor U7583 (N_7583,N_7091,N_5895);
nand U7584 (N_7584,N_6804,N_6501);
nor U7585 (N_7585,N_6080,N_5600);
xor U7586 (N_7586,N_7262,N_6348);
and U7587 (N_7587,N_5187,N_6862);
or U7588 (N_7588,N_5842,N_6009);
and U7589 (N_7589,N_6824,N_6889);
and U7590 (N_7590,N_6753,N_6599);
or U7591 (N_7591,N_7224,N_7217);
or U7592 (N_7592,N_5732,N_5627);
nor U7593 (N_7593,N_7241,N_6197);
and U7594 (N_7594,N_6153,N_6605);
nand U7595 (N_7595,N_6419,N_6471);
nor U7596 (N_7596,N_6196,N_6281);
nor U7597 (N_7597,N_6557,N_5127);
nand U7598 (N_7598,N_6283,N_6326);
nand U7599 (N_7599,N_5434,N_7324);
and U7600 (N_7600,N_5367,N_5340);
xor U7601 (N_7601,N_6865,N_5365);
or U7602 (N_7602,N_6328,N_5069);
xor U7603 (N_7603,N_6649,N_6911);
nand U7604 (N_7604,N_6304,N_6735);
nor U7605 (N_7605,N_6100,N_5068);
nand U7606 (N_7606,N_7403,N_6414);
and U7607 (N_7607,N_7289,N_5965);
and U7608 (N_7608,N_6290,N_6363);
xor U7609 (N_7609,N_7188,N_7394);
and U7610 (N_7610,N_7427,N_6896);
nand U7611 (N_7611,N_7154,N_5296);
nand U7612 (N_7612,N_6771,N_5224);
and U7613 (N_7613,N_5909,N_6754);
nand U7614 (N_7614,N_7000,N_6914);
nand U7615 (N_7615,N_5854,N_6336);
or U7616 (N_7616,N_5147,N_5279);
or U7617 (N_7617,N_5320,N_7401);
and U7618 (N_7618,N_7264,N_6127);
nor U7619 (N_7619,N_7228,N_5745);
and U7620 (N_7620,N_5805,N_6147);
nor U7621 (N_7621,N_7235,N_7413);
or U7622 (N_7622,N_6233,N_5189);
nand U7623 (N_7623,N_6636,N_5404);
nor U7624 (N_7624,N_7055,N_5117);
and U7625 (N_7625,N_5661,N_6714);
nor U7626 (N_7626,N_6016,N_6245);
nor U7627 (N_7627,N_7485,N_5658);
nor U7628 (N_7628,N_5354,N_7182);
nand U7629 (N_7629,N_5014,N_7292);
nor U7630 (N_7630,N_7070,N_6358);
or U7631 (N_7631,N_5517,N_6404);
or U7632 (N_7632,N_7204,N_7001);
nand U7633 (N_7633,N_5940,N_5158);
or U7634 (N_7634,N_6765,N_5597);
xnor U7635 (N_7635,N_7135,N_6993);
and U7636 (N_7636,N_6828,N_5263);
or U7637 (N_7637,N_6466,N_5535);
or U7638 (N_7638,N_5608,N_5268);
and U7639 (N_7639,N_5304,N_7471);
and U7640 (N_7640,N_5034,N_6789);
or U7641 (N_7641,N_6985,N_6305);
nor U7642 (N_7642,N_6634,N_6686);
nand U7643 (N_7643,N_5680,N_5651);
nand U7644 (N_7644,N_6848,N_5414);
or U7645 (N_7645,N_6491,N_5943);
or U7646 (N_7646,N_6061,N_6899);
xnor U7647 (N_7647,N_6221,N_5495);
xor U7648 (N_7648,N_6306,N_6670);
xnor U7649 (N_7649,N_6448,N_6518);
nor U7650 (N_7650,N_5148,N_5646);
nand U7651 (N_7651,N_5954,N_6619);
nor U7652 (N_7652,N_6318,N_5811);
nor U7653 (N_7653,N_6201,N_5793);
nand U7654 (N_7654,N_5962,N_5625);
nor U7655 (N_7655,N_5698,N_5032);
or U7656 (N_7656,N_5172,N_6246);
nor U7657 (N_7657,N_5933,N_5823);
xnor U7658 (N_7658,N_7391,N_5097);
nand U7659 (N_7659,N_5229,N_6710);
and U7660 (N_7660,N_5669,N_5609);
nor U7661 (N_7661,N_5999,N_5972);
nand U7662 (N_7662,N_5214,N_6979);
nand U7663 (N_7663,N_6543,N_6756);
and U7664 (N_7664,N_6160,N_6785);
nand U7665 (N_7665,N_5699,N_6186);
nand U7666 (N_7666,N_6408,N_7492);
and U7667 (N_7667,N_5440,N_7057);
nand U7668 (N_7668,N_6470,N_6536);
or U7669 (N_7669,N_6372,N_7283);
or U7670 (N_7670,N_6473,N_6062);
nand U7671 (N_7671,N_7296,N_6384);
nor U7672 (N_7672,N_5358,N_6316);
nor U7673 (N_7673,N_5194,N_5806);
and U7674 (N_7674,N_5937,N_5944);
nand U7675 (N_7675,N_5644,N_7059);
or U7676 (N_7676,N_5153,N_5300);
or U7677 (N_7677,N_6874,N_5144);
or U7678 (N_7678,N_6700,N_6692);
xor U7679 (N_7679,N_6996,N_5013);
xnor U7680 (N_7680,N_6967,N_7073);
and U7681 (N_7681,N_6887,N_5246);
or U7682 (N_7682,N_6239,N_5998);
or U7683 (N_7683,N_6935,N_6926);
nor U7684 (N_7684,N_5889,N_7088);
nand U7685 (N_7685,N_5635,N_5461);
nand U7686 (N_7686,N_5168,N_5110);
nor U7687 (N_7687,N_5576,N_6535);
or U7688 (N_7688,N_7376,N_5104);
xor U7689 (N_7689,N_5432,N_6880);
nand U7690 (N_7690,N_6299,N_5039);
or U7691 (N_7691,N_6421,N_6278);
xor U7692 (N_7692,N_5865,N_6642);
nor U7693 (N_7693,N_5218,N_6742);
nor U7694 (N_7694,N_5396,N_6973);
or U7695 (N_7695,N_7279,N_6088);
and U7696 (N_7696,N_7172,N_5463);
nand U7697 (N_7697,N_6240,N_6451);
and U7698 (N_7698,N_5791,N_6128);
and U7699 (N_7699,N_6928,N_7408);
xor U7700 (N_7700,N_5058,N_6608);
and U7701 (N_7701,N_6146,N_7179);
nand U7702 (N_7702,N_7362,N_5726);
or U7703 (N_7703,N_6875,N_7024);
xor U7704 (N_7704,N_6528,N_5109);
and U7705 (N_7705,N_5848,N_7229);
nand U7706 (N_7706,N_7393,N_5717);
nor U7707 (N_7707,N_6676,N_5009);
nand U7708 (N_7708,N_6029,N_6437);
nor U7709 (N_7709,N_6888,N_5468);
or U7710 (N_7710,N_6091,N_7083);
and U7711 (N_7711,N_5991,N_6718);
nor U7712 (N_7712,N_6067,N_5286);
and U7713 (N_7713,N_6620,N_5986);
or U7714 (N_7714,N_7349,N_5728);
nand U7715 (N_7715,N_7072,N_5073);
and U7716 (N_7716,N_7280,N_5210);
nand U7717 (N_7717,N_7331,N_5507);
nand U7718 (N_7718,N_6740,N_7341);
xor U7719 (N_7719,N_6360,N_6774);
xor U7720 (N_7720,N_7406,N_5884);
nand U7721 (N_7721,N_6724,N_5677);
or U7722 (N_7722,N_6431,N_6959);
nor U7723 (N_7723,N_6660,N_5555);
and U7724 (N_7724,N_6181,N_6440);
nor U7725 (N_7725,N_7042,N_6823);
and U7726 (N_7726,N_6276,N_5668);
nor U7727 (N_7727,N_5182,N_6486);
and U7728 (N_7728,N_5359,N_6727);
and U7729 (N_7729,N_5603,N_5352);
and U7730 (N_7730,N_7461,N_6861);
nor U7731 (N_7731,N_7298,N_5970);
nor U7732 (N_7732,N_6517,N_6027);
nor U7733 (N_7733,N_7399,N_5676);
or U7734 (N_7734,N_7020,N_6708);
nand U7735 (N_7735,N_6078,N_6641);
or U7736 (N_7736,N_7177,N_7373);
nor U7737 (N_7737,N_5211,N_7437);
and U7738 (N_7738,N_6898,N_5024);
and U7739 (N_7739,N_5385,N_5176);
and U7740 (N_7740,N_5128,N_5615);
or U7741 (N_7741,N_5612,N_6168);
nand U7742 (N_7742,N_5265,N_6931);
or U7743 (N_7743,N_5893,N_5037);
nor U7744 (N_7744,N_6939,N_5235);
nand U7745 (N_7745,N_5469,N_6286);
or U7746 (N_7746,N_6937,N_7017);
or U7747 (N_7747,N_6904,N_6585);
xnor U7748 (N_7748,N_7221,N_7276);
or U7749 (N_7749,N_5227,N_5018);
and U7750 (N_7750,N_6402,N_6007);
and U7751 (N_7751,N_5927,N_5093);
or U7752 (N_7752,N_5729,N_7248);
xor U7753 (N_7753,N_6174,N_5656);
and U7754 (N_7754,N_5995,N_6901);
or U7755 (N_7755,N_5038,N_6721);
nand U7756 (N_7756,N_7265,N_7442);
or U7757 (N_7757,N_5366,N_6600);
or U7758 (N_7758,N_7161,N_6624);
or U7759 (N_7759,N_5048,N_6312);
or U7760 (N_7760,N_6726,N_6117);
nor U7761 (N_7761,N_5643,N_6445);
and U7762 (N_7762,N_5178,N_5558);
nand U7763 (N_7763,N_5885,N_5742);
nand U7764 (N_7764,N_6120,N_6796);
or U7765 (N_7765,N_7431,N_7335);
and U7766 (N_7766,N_5531,N_5107);
or U7767 (N_7767,N_5186,N_5377);
nor U7768 (N_7768,N_7170,N_6251);
nor U7769 (N_7769,N_6136,N_6017);
or U7770 (N_7770,N_5861,N_6023);
and U7771 (N_7771,N_5741,N_7367);
or U7772 (N_7772,N_5425,N_5493);
or U7773 (N_7773,N_6579,N_5212);
and U7774 (N_7774,N_5666,N_6370);
and U7775 (N_7775,N_5314,N_6213);
or U7776 (N_7776,N_5833,N_5958);
and U7777 (N_7777,N_5201,N_7479);
nand U7778 (N_7778,N_5920,N_7309);
and U7779 (N_7779,N_5490,N_6036);
xnor U7780 (N_7780,N_5990,N_6275);
or U7781 (N_7781,N_6092,N_5383);
nor U7782 (N_7782,N_5510,N_7358);
and U7783 (N_7783,N_5957,N_6142);
xnor U7784 (N_7784,N_7272,N_6294);
nor U7785 (N_7785,N_6791,N_5449);
nand U7786 (N_7786,N_5311,N_5353);
nor U7787 (N_7787,N_5239,N_5159);
nor U7788 (N_7788,N_6032,N_6712);
nor U7789 (N_7789,N_5479,N_5284);
nand U7790 (N_7790,N_5593,N_5619);
or U7791 (N_7791,N_6678,N_6034);
nand U7792 (N_7792,N_5525,N_5869);
nand U7793 (N_7793,N_6520,N_7452);
and U7794 (N_7794,N_7082,N_5620);
and U7795 (N_7795,N_6463,N_6732);
or U7796 (N_7796,N_7480,N_6607);
nand U7797 (N_7797,N_6577,N_5701);
nor U7798 (N_7798,N_5511,N_7140);
xnor U7799 (N_7799,N_5915,N_7332);
and U7800 (N_7800,N_6151,N_6940);
nor U7801 (N_7801,N_6065,N_6332);
or U7802 (N_7802,N_5223,N_7223);
and U7803 (N_7803,N_5537,N_7495);
nand U7804 (N_7804,N_7164,N_7102);
or U7805 (N_7805,N_5271,N_5981);
nor U7806 (N_7806,N_6610,N_6545);
nand U7807 (N_7807,N_5342,N_5921);
and U7808 (N_7808,N_7149,N_5106);
or U7809 (N_7809,N_6130,N_5071);
nor U7810 (N_7810,N_6411,N_6521);
and U7811 (N_7811,N_6556,N_5336);
and U7812 (N_7812,N_6664,N_6439);
and U7813 (N_7813,N_6671,N_5195);
xor U7814 (N_7814,N_7348,N_6375);
or U7815 (N_7815,N_5825,N_6698);
nor U7816 (N_7816,N_7313,N_6184);
xnor U7817 (N_7817,N_6008,N_6825);
nor U7818 (N_7818,N_7269,N_6905);
nor U7819 (N_7819,N_5587,N_5611);
or U7820 (N_7820,N_6857,N_5906);
and U7821 (N_7821,N_5204,N_6685);
nor U7822 (N_7822,N_5459,N_7120);
nor U7823 (N_7823,N_6544,N_5989);
nor U7824 (N_7824,N_7104,N_6443);
nor U7825 (N_7825,N_6999,N_7286);
nor U7826 (N_7826,N_6050,N_6182);
or U7827 (N_7827,N_5772,N_6005);
and U7828 (N_7828,N_6192,N_5569);
nor U7829 (N_7829,N_5278,N_6205);
nor U7830 (N_7830,N_5456,N_7036);
and U7831 (N_7831,N_7166,N_6357);
nor U7832 (N_7832,N_6177,N_6910);
or U7833 (N_7833,N_5083,N_6046);
xnor U7834 (N_7834,N_7407,N_7462);
xnor U7835 (N_7835,N_5527,N_5481);
or U7836 (N_7836,N_6787,N_6695);
nor U7837 (N_7837,N_6717,N_5022);
nand U7838 (N_7838,N_5554,N_5640);
or U7839 (N_7839,N_5193,N_7054);
and U7840 (N_7840,N_5166,N_6341);
and U7841 (N_7841,N_6749,N_6238);
or U7842 (N_7842,N_5975,N_7301);
nor U7843 (N_7843,N_5057,N_5051);
and U7844 (N_7844,N_6334,N_5673);
nand U7845 (N_7845,N_6962,N_6883);
nor U7846 (N_7846,N_6492,N_5544);
nor U7847 (N_7847,N_5140,N_5886);
xnor U7848 (N_7848,N_6262,N_5697);
or U7849 (N_7849,N_5992,N_6815);
nand U7850 (N_7850,N_5606,N_6230);
and U7851 (N_7851,N_6793,N_7278);
or U7852 (N_7852,N_5581,N_7203);
and U7853 (N_7853,N_6612,N_5549);
or U7854 (N_7854,N_6941,N_5623);
nor U7855 (N_7855,N_5007,N_6524);
nor U7856 (N_7856,N_7151,N_5475);
or U7857 (N_7857,N_6021,N_6723);
or U7858 (N_7858,N_6747,N_5394);
or U7859 (N_7859,N_6583,N_6339);
nor U7860 (N_7860,N_6589,N_5264);
nor U7861 (N_7861,N_6506,N_5904);
nand U7862 (N_7862,N_5136,N_7111);
and U7863 (N_7863,N_6256,N_6482);
nor U7864 (N_7864,N_6075,N_6683);
and U7865 (N_7865,N_5457,N_6068);
or U7866 (N_7866,N_6906,N_6667);
or U7867 (N_7867,N_6398,N_5451);
and U7868 (N_7868,N_5041,N_7300);
nor U7869 (N_7869,N_5023,N_6522);
xor U7870 (N_7870,N_7029,N_6775);
nor U7871 (N_7871,N_5252,N_6587);
nand U7872 (N_7872,N_7090,N_5711);
or U7873 (N_7873,N_5063,N_6766);
and U7874 (N_7874,N_5444,N_6609);
nand U7875 (N_7875,N_6540,N_6509);
and U7876 (N_7876,N_7414,N_7384);
nor U7877 (N_7877,N_5322,N_5551);
or U7878 (N_7878,N_6322,N_6943);
nor U7879 (N_7879,N_6854,N_5005);
xnor U7880 (N_7880,N_6949,N_6707);
nand U7881 (N_7881,N_7062,N_5733);
nor U7882 (N_7882,N_7435,N_5375);
xnor U7883 (N_7883,N_6387,N_6260);
nor U7884 (N_7884,N_6126,N_6161);
and U7885 (N_7885,N_7037,N_7429);
nand U7886 (N_7886,N_6936,N_6878);
xnor U7887 (N_7887,N_6222,N_6755);
or U7888 (N_7888,N_6541,N_7330);
nor U7889 (N_7889,N_6198,N_6814);
nand U7890 (N_7890,N_5035,N_6119);
nand U7891 (N_7891,N_6715,N_7096);
nor U7892 (N_7892,N_7199,N_6855);
and U7893 (N_7893,N_5143,N_5338);
nand U7894 (N_7894,N_5371,N_5494);
or U7895 (N_7895,N_5770,N_6868);
or U7896 (N_7896,N_5090,N_5033);
or U7897 (N_7897,N_6643,N_6548);
or U7898 (N_7898,N_7048,N_6379);
or U7899 (N_7899,N_7234,N_5773);
xnor U7900 (N_7900,N_5372,N_5310);
nor U7901 (N_7901,N_5070,N_6798);
nand U7902 (N_7902,N_6764,N_6070);
nand U7903 (N_7903,N_7499,N_6455);
and U7904 (N_7904,N_6257,N_6042);
nand U7905 (N_7905,N_5179,N_6762);
or U7906 (N_7906,N_6041,N_5704);
nand U7907 (N_7907,N_5727,N_7069);
and U7908 (N_7908,N_5540,N_6303);
or U7909 (N_7909,N_6069,N_6992);
nand U7910 (N_7910,N_5696,N_7052);
nor U7911 (N_7911,N_5720,N_7288);
or U7912 (N_7912,N_5081,N_7089);
xor U7913 (N_7913,N_5942,N_6494);
nand U7914 (N_7914,N_5708,N_5514);
nor U7915 (N_7915,N_6369,N_7100);
nand U7916 (N_7916,N_6018,N_5877);
nor U7917 (N_7917,N_5580,N_5781);
nand U7918 (N_7918,N_5253,N_5546);
or U7919 (N_7919,N_5938,N_6971);
and U7920 (N_7920,N_7398,N_6551);
nor U7921 (N_7921,N_6300,N_5205);
nor U7922 (N_7922,N_5519,N_7115);
or U7923 (N_7923,N_6432,N_6190);
nor U7924 (N_7924,N_5133,N_7385);
nand U7925 (N_7925,N_6652,N_6309);
nor U7926 (N_7926,N_6225,N_7246);
and U7927 (N_7927,N_5430,N_5301);
nand U7928 (N_7928,N_6675,N_7006);
nand U7929 (N_7929,N_5429,N_5583);
or U7930 (N_7930,N_6594,N_6961);
nand U7931 (N_7931,N_7418,N_6954);
xor U7932 (N_7932,N_5096,N_5907);
and U7933 (N_7933,N_5971,N_6618);
and U7934 (N_7934,N_6554,N_5575);
nor U7935 (N_7935,N_7066,N_5797);
and U7936 (N_7936,N_6921,N_6981);
and U7937 (N_7937,N_6866,N_6415);
and U7938 (N_7938,N_6821,N_6661);
and U7939 (N_7939,N_5170,N_5843);
nand U7940 (N_7940,N_6340,N_7122);
or U7941 (N_7941,N_6493,N_6014);
and U7942 (N_7942,N_6640,N_5826);
or U7943 (N_7943,N_5062,N_5231);
nor U7944 (N_7944,N_5775,N_6138);
nor U7945 (N_7945,N_5219,N_6438);
nor U7946 (N_7946,N_6809,N_5631);
and U7947 (N_7947,N_6832,N_5181);
xnor U7948 (N_7948,N_6071,N_6656);
or U7949 (N_7949,N_5795,N_7340);
nor U7950 (N_7950,N_6420,N_6456);
or U7951 (N_7951,N_5715,N_5767);
nand U7952 (N_7952,N_6930,N_6792);
or U7953 (N_7953,N_5559,N_5557);
nand U7954 (N_7954,N_5908,N_6978);
nand U7955 (N_7955,N_6542,N_5874);
nor U7956 (N_7956,N_7013,N_5466);
nor U7957 (N_7957,N_7259,N_5074);
and U7958 (N_7958,N_6076,N_5431);
or U7959 (N_7959,N_5637,N_5591);
xnor U7960 (N_7960,N_5538,N_5348);
nand U7961 (N_7961,N_5010,N_6394);
or U7962 (N_7962,N_5512,N_7325);
or U7963 (N_7963,N_5845,N_5376);
nand U7964 (N_7964,N_5776,N_6812);
nor U7965 (N_7965,N_6842,N_7114);
xnor U7966 (N_7966,N_6575,N_7118);
and U7967 (N_7967,N_5473,N_6945);
xor U7968 (N_7968,N_6659,N_5234);
or U7969 (N_7969,N_6550,N_5384);
nand U7970 (N_7970,N_5454,N_6442);
nor U7971 (N_7971,N_5934,N_7440);
nor U7972 (N_7972,N_5832,N_7284);
and U7973 (N_7973,N_6907,N_6179);
nor U7974 (N_7974,N_5064,N_5207);
nor U7975 (N_7975,N_6519,N_7302);
or U7976 (N_7976,N_5948,N_6813);
xnor U7977 (N_7977,N_6533,N_6366);
and U7978 (N_7978,N_5712,N_7379);
or U7979 (N_7979,N_7132,N_6739);
and U7980 (N_7980,N_5543,N_6552);
nor U7981 (N_7981,N_6873,N_6244);
and U7982 (N_7982,N_5924,N_6362);
or U7983 (N_7983,N_6799,N_5021);
or U7984 (N_7984,N_5118,N_6523);
and U7985 (N_7985,N_7488,N_5327);
nand U7986 (N_7986,N_5137,N_7117);
or U7987 (N_7987,N_6314,N_5163);
or U7988 (N_7988,N_6165,N_5164);
nand U7989 (N_7989,N_7148,N_5003);
and U7990 (N_7990,N_6558,N_5111);
and U7991 (N_7991,N_5856,N_7453);
and U7992 (N_7992,N_7004,N_6460);
and U7993 (N_7993,N_5419,N_6925);
and U7994 (N_7994,N_6401,N_6131);
nor U7995 (N_7995,N_5131,N_5562);
or U7996 (N_7996,N_5135,N_7035);
nor U7997 (N_7997,N_6356,N_5536);
or U7998 (N_7998,N_7047,N_6291);
xor U7999 (N_7999,N_5901,N_7053);
and U8000 (N_8000,N_6383,N_5653);
and U8001 (N_8001,N_6948,N_5483);
or U8002 (N_8002,N_7470,N_5758);
or U8003 (N_8003,N_7143,N_5961);
xor U8004 (N_8004,N_6422,N_6863);
nand U8005 (N_8005,N_7273,N_7023);
or U8006 (N_8006,N_6831,N_5734);
or U8007 (N_8007,N_6039,N_6565);
or U8008 (N_8008,N_6220,N_6321);
nor U8009 (N_8009,N_6129,N_5332);
xnor U8010 (N_8010,N_7212,N_5043);
nand U8011 (N_8011,N_5967,N_6218);
or U8012 (N_8012,N_5059,N_7455);
or U8013 (N_8013,N_5794,N_7422);
and U8014 (N_8014,N_6313,N_5817);
and U8015 (N_8015,N_5761,N_6655);
nor U8016 (N_8016,N_6805,N_5448);
or U8017 (N_8017,N_6472,N_6085);
nor U8018 (N_8018,N_6497,N_6392);
nor U8019 (N_8019,N_5217,N_5700);
or U8020 (N_8020,N_5855,N_6324);
nand U8021 (N_8021,N_5796,N_5244);
nand U8022 (N_8022,N_5679,N_6020);
xnor U8023 (N_8023,N_6604,N_6574);
nand U8024 (N_8024,N_7294,N_6301);
nor U8025 (N_8025,N_5804,N_5830);
or U8026 (N_8026,N_7176,N_6242);
or U8027 (N_8027,N_5220,N_7450);
nand U8028 (N_8028,N_6056,N_6511);
and U8029 (N_8029,N_5801,N_7377);
and U8030 (N_8030,N_5424,N_5484);
xor U8031 (N_8031,N_5683,N_5955);
nand U8032 (N_8032,N_5883,N_7359);
nor U8033 (N_8033,N_5180,N_6677);
nand U8034 (N_8034,N_7257,N_7127);
nor U8035 (N_8035,N_5800,N_7295);
nand U8036 (N_8036,N_7327,N_7019);
nand U8037 (N_8037,N_6613,N_7383);
xnor U8038 (N_8038,N_6788,N_5584);
and U8039 (N_8039,N_7124,N_6135);
nand U8040 (N_8040,N_6833,N_6329);
or U8041 (N_8041,N_6269,N_5266);
and U8042 (N_8042,N_5245,N_5760);
and U8043 (N_8043,N_6696,N_5076);
nor U8044 (N_8044,N_6298,N_5628);
and U8045 (N_8045,N_6975,N_5067);
nand U8046 (N_8046,N_7061,N_5652);
or U8047 (N_8047,N_7167,N_5397);
xor U8048 (N_8048,N_6886,N_6011);
nor U8049 (N_8049,N_5077,N_5149);
nand U8050 (N_8050,N_5052,N_6586);
xor U8051 (N_8051,N_6516,N_5395);
or U8052 (N_8052,N_5724,N_6713);
or U8053 (N_8053,N_5108,N_6323);
xnor U8054 (N_8054,N_6860,N_6354);
and U8055 (N_8055,N_5138,N_5156);
and U8056 (N_8056,N_6288,N_7420);
and U8057 (N_8057,N_6441,N_5303);
nor U8058 (N_8058,N_7293,N_5198);
and U8059 (N_8059,N_5532,N_6350);
and U8060 (N_8060,N_5663,N_5087);
nor U8061 (N_8061,N_7109,N_6094);
and U8062 (N_8062,N_5026,N_5025);
xnor U8063 (N_8063,N_5878,N_6057);
or U8064 (N_8064,N_7356,N_5784);
nand U8065 (N_8065,N_6424,N_5814);
and U8066 (N_8066,N_6156,N_7160);
nor U8067 (N_8067,N_7336,N_6134);
xnor U8068 (N_8068,N_6287,N_7159);
nand U8069 (N_8069,N_6436,N_7395);
xor U8070 (N_8070,N_5506,N_5417);
and U8071 (N_8071,N_7094,N_5247);
or U8072 (N_8072,N_7436,N_5738);
nor U8073 (N_8073,N_5821,N_5686);
or U8074 (N_8074,N_5573,N_7285);
nor U8075 (N_8075,N_5325,N_5122);
and U8076 (N_8076,N_7417,N_6248);
nor U8077 (N_8077,N_5488,N_7190);
xnor U8078 (N_8078,N_7144,N_5530);
nand U8079 (N_8079,N_5542,N_5616);
xor U8080 (N_8080,N_5988,N_5752);
nand U8081 (N_8081,N_5870,N_6744);
or U8082 (N_8082,N_6674,N_7274);
xnor U8083 (N_8083,N_6279,N_6951);
or U8084 (N_8084,N_6297,N_5850);
or U8085 (N_8085,N_5755,N_7473);
and U8086 (N_8086,N_5840,N_5313);
or U8087 (N_8087,N_5334,N_5743);
or U8088 (N_8088,N_5150,N_6955);
nand U8089 (N_8089,N_7139,N_5577);
or U8090 (N_8090,N_5935,N_5504);
nor U8091 (N_8091,N_7423,N_6417);
and U8092 (N_8092,N_6803,N_6897);
xor U8093 (N_8093,N_7308,N_6343);
and U8094 (N_8094,N_5592,N_7491);
xor U8095 (N_8095,N_5578,N_5678);
and U8096 (N_8096,N_7180,N_5947);
nand U8097 (N_8097,N_7323,N_5486);
nand U8098 (N_8098,N_7322,N_6639);
xnor U8099 (N_8099,N_5171,N_5523);
nor U8100 (N_8100,N_7181,N_6498);
or U8101 (N_8101,N_6790,N_6876);
nor U8102 (N_8102,N_6982,N_6141);
nor U8103 (N_8103,N_5739,N_7498);
or U8104 (N_8104,N_7361,N_6709);
nor U8105 (N_8105,N_5123,N_6572);
or U8106 (N_8106,N_5317,N_5571);
nand U8107 (N_8107,N_7240,N_7189);
nand U8108 (N_8108,N_6512,N_6381);
xor U8109 (N_8109,N_5197,N_5120);
and U8110 (N_8110,N_7380,N_7354);
or U8111 (N_8111,N_5875,N_6990);
nand U8112 (N_8112,N_6734,N_5046);
nand U8113 (N_8113,N_5570,N_5694);
and U8114 (N_8114,N_5155,N_5868);
and U8115 (N_8115,N_5987,N_5939);
or U8116 (N_8116,N_6782,N_6209);
and U8117 (N_8117,N_6480,N_6818);
and U8118 (N_8118,N_5349,N_7247);
xor U8119 (N_8119,N_7200,N_7171);
or U8120 (N_8120,N_6157,N_6426);
and U8121 (N_8121,N_5790,N_7347);
or U8122 (N_8122,N_6741,N_6019);
and U8123 (N_8123,N_7360,N_5930);
or U8124 (N_8124,N_5762,N_6847);
nor U8125 (N_8125,N_6001,N_5453);
or U8126 (N_8126,N_5061,N_6684);
nor U8127 (N_8127,N_5818,N_5803);
and U8128 (N_8128,N_6780,N_5498);
nor U8129 (N_8129,N_7071,N_6808);
nand U8130 (N_8130,N_6217,N_6826);
and U8131 (N_8131,N_5084,N_5196);
or U8132 (N_8132,N_5289,N_7447);
and U8133 (N_8133,N_7351,N_5598);
and U8134 (N_8134,N_5436,N_6423);
and U8135 (N_8135,N_5116,N_7382);
or U8136 (N_8136,N_5896,N_7174);
and U8137 (N_8137,N_6345,N_6617);
nand U8138 (N_8138,N_6228,N_5029);
nor U8139 (N_8139,N_6349,N_5813);
or U8140 (N_8140,N_5202,N_6646);
or U8141 (N_8141,N_6651,N_6615);
and U8142 (N_8142,N_5860,N_6025);
nor U8143 (N_8143,N_5632,N_5442);
nand U8144 (N_8144,N_6648,N_5403);
or U8145 (N_8145,N_7486,N_7416);
or U8146 (N_8146,N_7163,N_6997);
and U8147 (N_8147,N_7466,N_5226);
or U8148 (N_8148,N_6399,N_7112);
nand U8149 (N_8149,N_5256,N_6079);
and U8150 (N_8150,N_6527,N_7075);
nor U8151 (N_8151,N_7205,N_5516);
xnor U8152 (N_8152,N_5956,N_6946);
nand U8153 (N_8153,N_6215,N_5487);
nor U8154 (N_8154,N_5911,N_7002);
and U8155 (N_8155,N_6364,N_7243);
xor U8156 (N_8156,N_6371,N_5905);
nand U8157 (N_8157,N_6730,N_5873);
xor U8158 (N_8158,N_5852,N_7303);
nand U8159 (N_8159,N_7400,N_6560);
or U8160 (N_8160,N_6746,N_7369);
nor U8161 (N_8161,N_6690,N_7329);
and U8162 (N_8162,N_5091,N_5031);
nand U8163 (N_8163,N_5674,N_6879);
nor U8164 (N_8164,N_5650,N_5307);
nand U8165 (N_8165,N_7026,N_5326);
or U8166 (N_8166,N_5968,N_5390);
nor U8167 (N_8167,N_5664,N_5250);
nor U8168 (N_8168,N_6388,N_7152);
nand U8169 (N_8169,N_7097,N_6047);
nand U8170 (N_8170,N_7010,N_6737);
nand U8171 (N_8171,N_7249,N_5019);
or U8172 (N_8172,N_6924,N_6743);
and U8173 (N_8173,N_5027,N_5787);
nand U8174 (N_8174,N_6820,N_7044);
or U8175 (N_8175,N_5879,N_5882);
or U8176 (N_8176,N_5269,N_5000);
nor U8177 (N_8177,N_5605,N_6702);
nor U8178 (N_8178,N_5588,N_5524);
and U8179 (N_8179,N_5691,N_5659);
and U8180 (N_8180,N_6189,N_6212);
nor U8181 (N_8181,N_6917,N_5098);
nor U8182 (N_8182,N_6169,N_6852);
and U8183 (N_8183,N_5505,N_5515);
or U8184 (N_8184,N_6631,N_5902);
and U8185 (N_8185,N_5312,N_6998);
xor U8186 (N_8186,N_6932,N_7129);
nand U8187 (N_8187,N_7194,N_7378);
nand U8188 (N_8188,N_6502,N_6004);
and U8189 (N_8189,N_6368,N_5645);
or U8190 (N_8190,N_5655,N_7350);
or U8191 (N_8191,N_5765,N_5736);
or U8192 (N_8192,N_5445,N_6327);
or U8193 (N_8193,N_7142,N_6507);
and U8194 (N_8194,N_5913,N_7009);
xor U8195 (N_8195,N_6705,N_7081);
and U8196 (N_8196,N_7267,N_7078);
and U8197 (N_8197,N_7368,N_5040);
nand U8198 (N_8198,N_7033,N_7056);
and U8199 (N_8199,N_5703,N_5199);
nor U8200 (N_8200,N_7311,N_5626);
and U8201 (N_8201,N_7261,N_6703);
or U8202 (N_8202,N_7493,N_5427);
or U8203 (N_8203,N_5949,N_5789);
and U8204 (N_8204,N_6012,N_6802);
xnor U8205 (N_8205,N_5997,N_6869);
nand U8206 (N_8206,N_7186,N_6066);
and U8207 (N_8207,N_6877,N_5400);
and U8208 (N_8208,N_5914,N_5161);
nor U8209 (N_8209,N_5175,N_6315);
nand U8210 (N_8210,N_5114,N_6103);
xor U8211 (N_8211,N_7372,N_5343);
nor U8212 (N_8212,N_6320,N_7049);
and U8213 (N_8213,N_6621,N_5528);
nand U8214 (N_8214,N_5594,N_6701);
nand U8215 (N_8215,N_7497,N_6638);
nand U8216 (N_8216,N_6908,N_5521);
or U8217 (N_8217,N_5260,N_5030);
and U8218 (N_8218,N_5748,N_6529);
nand U8219 (N_8219,N_5125,N_6628);
nor U8220 (N_8220,N_6110,N_6477);
xor U8221 (N_8221,N_6531,N_6614);
nor U8222 (N_8222,N_6444,N_7092);
nor U8223 (N_8223,N_5834,N_7067);
xor U8224 (N_8224,N_6496,N_6835);
nand U8225 (N_8225,N_7187,N_5816);
or U8226 (N_8226,N_6530,N_6231);
or U8227 (N_8227,N_5363,N_6778);
nand U8228 (N_8228,N_5518,N_5167);
and U8229 (N_8229,N_5747,N_6194);
and U8230 (N_8230,N_6693,N_6987);
nor U8231 (N_8231,N_6185,N_5350);
nand U8232 (N_8232,N_5339,N_7446);
nand U8233 (N_8233,N_7084,N_5500);
and U8234 (N_8234,N_6204,N_5867);
xnor U8235 (N_8235,N_6022,N_5929);
or U8236 (N_8236,N_5331,N_6947);
nor U8237 (N_8237,N_5401,N_7277);
xor U8238 (N_8238,N_7305,N_7011);
nor U8239 (N_8239,N_5928,N_5124);
nand U8240 (N_8240,N_6284,N_5200);
and U8241 (N_8241,N_5894,N_6794);
or U8242 (N_8242,N_6464,N_5926);
nand U8243 (N_8243,N_6567,N_6206);
nor U8244 (N_8244,N_7060,N_6719);
or U8245 (N_8245,N_6243,N_5464);
or U8246 (N_8246,N_5422,N_6259);
nor U8247 (N_8247,N_7475,N_6236);
nor U8248 (N_8248,N_5778,N_6407);
and U8249 (N_8249,N_6187,N_6697);
or U8250 (N_8250,N_7012,N_5055);
or U8251 (N_8251,N_5572,N_5347);
xor U8252 (N_8252,N_6155,N_6630);
nor U8253 (N_8253,N_5132,N_6429);
nand U8254 (N_8254,N_5862,N_6839);
xnor U8255 (N_8255,N_6694,N_6644);
or U8256 (N_8256,N_7169,N_5413);
and U8257 (N_8257,N_5257,N_7219);
or U8258 (N_8258,N_5480,N_5714);
or U8259 (N_8259,N_7252,N_5173);
nor U8260 (N_8260,N_6468,N_7145);
nand U8261 (N_8261,N_6584,N_7374);
nand U8262 (N_8262,N_7312,N_5857);
xnor U8263 (N_8263,N_5085,N_6784);
nand U8264 (N_8264,N_7366,N_5757);
nor U8265 (N_8265,N_6980,N_5685);
nor U8266 (N_8266,N_6953,N_6977);
nor U8267 (N_8267,N_5730,N_5446);
or U8268 (N_8268,N_6410,N_5783);
and U8269 (N_8269,N_7387,N_5478);
nor U8270 (N_8270,N_7025,N_6089);
or U8271 (N_8271,N_6964,N_7255);
nor U8272 (N_8272,N_5006,N_5185);
xor U8273 (N_8273,N_5660,N_6073);
or U8274 (N_8274,N_7472,N_6446);
and U8275 (N_8275,N_7185,N_6900);
nand U8276 (N_8276,N_6758,N_5812);
or U8277 (N_8277,N_5599,N_6475);
and U8278 (N_8278,N_6264,N_6199);
xor U8279 (N_8279,N_6400,N_6633);
or U8280 (N_8280,N_5485,N_6768);
nand U8281 (N_8281,N_7268,N_7468);
nor U8282 (N_8282,N_6296,N_7404);
and U8283 (N_8283,N_5437,N_6891);
and U8284 (N_8284,N_7027,N_5718);
and U8285 (N_8285,N_5617,N_7426);
nand U8286 (N_8286,N_5292,N_5287);
and U8287 (N_8287,N_6317,N_5251);
nor U8288 (N_8288,N_5295,N_6121);
nand U8289 (N_8289,N_6035,N_6107);
and U8290 (N_8290,N_5450,N_5952);
nor U8291 (N_8291,N_5082,N_6427);
nor U8292 (N_8292,N_5237,N_6273);
and U8293 (N_8293,N_6458,N_5820);
and U8294 (N_8294,N_5744,N_5008);
nor U8295 (N_8295,N_5319,N_5092);
or U8296 (N_8296,N_5851,N_5262);
and U8297 (N_8297,N_5567,N_5802);
or U8298 (N_8298,N_5984,N_6890);
and U8299 (N_8299,N_5838,N_5346);
and U8300 (N_8300,N_5740,N_6830);
xor U8301 (N_8301,N_6285,N_6211);
xor U8302 (N_8302,N_6603,N_5282);
and U8303 (N_8303,N_5017,N_6819);
or U8304 (N_8304,N_6669,N_6769);
nand U8305 (N_8305,N_5766,N_7196);
nand U8306 (N_8306,N_6006,N_6892);
and U8307 (N_8307,N_5184,N_6139);
or U8308 (N_8308,N_7291,N_6934);
nand U8309 (N_8309,N_5054,N_5308);
xnor U8310 (N_8310,N_5923,N_5344);
nand U8311 (N_8311,N_5735,N_7209);
or U8312 (N_8312,N_7251,N_5771);
nor U8313 (N_8313,N_5275,N_5782);
nor U8314 (N_8314,N_6082,N_6479);
nand U8315 (N_8315,N_5435,N_6525);
xor U8316 (N_8316,N_6390,N_7434);
nand U8317 (N_8317,N_5722,N_6270);
xor U8318 (N_8318,N_7282,N_7477);
nand U8319 (N_8319,N_6625,N_7321);
nor U8320 (N_8320,N_5582,N_5426);
nand U8321 (N_8321,N_6207,N_6461);
nor U8322 (N_8322,N_5078,N_7363);
xor U8323 (N_8323,N_6159,N_7441);
nor U8324 (N_8324,N_6549,N_7157);
and U8325 (N_8325,N_6920,N_7106);
and U8326 (N_8326,N_6172,N_6632);
xor U8327 (N_8327,N_5492,N_7271);
and U8328 (N_8328,N_5769,N_6716);
nor U8329 (N_8329,N_5604,N_5418);
nor U8330 (N_8330,N_7371,N_6829);
and U8331 (N_8331,N_6720,N_5272);
and U8332 (N_8332,N_6991,N_5357);
nand U8333 (N_8333,N_5539,N_5387);
or U8334 (N_8334,N_6810,N_7034);
and U8335 (N_8335,N_6894,N_6111);
nand U8336 (N_8336,N_6137,N_5080);
or U8337 (N_8337,N_5243,N_6919);
nor U8338 (N_8338,N_5513,N_5060);
nand U8339 (N_8339,N_6330,N_6561);
nand U8340 (N_8340,N_6505,N_6247);
nor U8341 (N_8341,N_6537,N_5897);
nand U8342 (N_8342,N_5853,N_5750);
xor U8343 (N_8343,N_5977,N_7392);
and U8344 (N_8344,N_6616,N_5684);
and U8345 (N_8345,N_5012,N_6033);
and U8346 (N_8346,N_7065,N_5545);
xor U8347 (N_8347,N_6736,N_5328);
and U8348 (N_8348,N_5183,N_6929);
and U8349 (N_8349,N_5474,N_6474);
and U8350 (N_8350,N_6028,N_5994);
and U8351 (N_8351,N_5721,N_5844);
nor U8352 (N_8352,N_6538,N_7306);
or U8353 (N_8353,N_5996,N_6870);
nor U8354 (N_8354,N_5682,N_7245);
xor U8355 (N_8355,N_5946,N_6353);
and U8356 (N_8356,N_5433,N_5931);
nor U8357 (N_8357,N_6510,N_6167);
or U8358 (N_8358,N_6772,N_6844);
nand U8359 (N_8359,N_6495,N_5258);
nor U8360 (N_8360,N_7465,N_5458);
and U8361 (N_8361,N_6581,N_5985);
and U8362 (N_8362,N_5809,N_5146);
and U8363 (N_8363,N_5723,N_7121);
and U8364 (N_8364,N_6467,N_5941);
or U8365 (N_8365,N_7334,N_5622);
xor U8366 (N_8366,N_5630,N_7214);
and U8367 (N_8367,N_6546,N_6418);
xor U8368 (N_8368,N_6406,N_7489);
nand U8369 (N_8369,N_7451,N_6188);
nor U8370 (N_8370,N_5409,N_5808);
nor U8371 (N_8371,N_6588,N_5585);
nor U8372 (N_8372,N_7165,N_6817);
or U8373 (N_8373,N_5047,N_5188);
nor U8374 (N_8374,N_6216,N_5174);
nor U8375 (N_8375,N_5642,N_7490);
nor U8376 (N_8376,N_5416,N_7079);
nor U8377 (N_8377,N_6836,N_5828);
or U8378 (N_8378,N_7058,N_6237);
or U8379 (N_8379,N_6602,N_5863);
nor U8380 (N_8380,N_7448,N_5360);
and U8381 (N_8381,N_7275,N_5807);
nand U8382 (N_8382,N_6465,N_6569);
or U8383 (N_8383,N_7326,N_6916);
or U8384 (N_8384,N_5402,N_5629);
xor U8385 (N_8385,N_6481,N_7231);
or U8386 (N_8386,N_5695,N_5912);
or U8387 (N_8387,N_7015,N_6310);
nand U8388 (N_8388,N_5075,N_6133);
nand U8389 (N_8389,N_5903,N_5560);
nand U8390 (N_8390,N_5113,N_6112);
and U8391 (N_8391,N_5254,N_7003);
nand U8392 (N_8392,N_6158,N_5315);
nor U8393 (N_8393,N_6881,N_6099);
nand U8394 (N_8394,N_6083,N_5509);
and U8395 (N_8395,N_5392,N_7068);
nand U8396 (N_8396,N_5382,N_7281);
and U8397 (N_8397,N_7236,N_6909);
or U8398 (N_8398,N_5103,N_5654);
nor U8399 (N_8399,N_7433,N_7041);
or U8400 (N_8400,N_7428,N_6054);
or U8401 (N_8401,N_7141,N_5533);
nand U8402 (N_8402,N_7412,N_6884);
or U8403 (N_8403,N_6942,N_5441);
or U8404 (N_8404,N_5267,N_6654);
or U8405 (N_8405,N_7220,N_5102);
nor U8406 (N_8406,N_6902,N_5471);
nand U8407 (N_8407,N_7410,N_7425);
nor U8408 (N_8408,N_5299,N_5380);
or U8409 (N_8409,N_5618,N_5979);
nand U8410 (N_8410,N_5053,N_6385);
xnor U8411 (N_8411,N_5373,N_6346);
xor U8412 (N_8412,N_6763,N_5681);
xor U8413 (N_8413,N_5341,N_6627);
nand U8414 (N_8414,N_5160,N_6093);
xor U8415 (N_8415,N_6152,N_6116);
or U8416 (N_8416,N_6532,N_7226);
or U8417 (N_8417,N_5438,N_5134);
nand U8418 (N_8418,N_7317,N_7421);
xor U8419 (N_8419,N_6430,N_5330);
nand U8420 (N_8420,N_6344,N_5919);
nand U8421 (N_8421,N_7481,N_6840);
or U8422 (N_8422,N_6547,N_6797);
and U8423 (N_8423,N_7230,N_7238);
and U8424 (N_8424,N_6647,N_7467);
or U8425 (N_8425,N_5596,N_5455);
and U8426 (N_8426,N_7197,N_6597);
nand U8427 (N_8427,N_6965,N_7454);
nand U8428 (N_8428,N_6267,N_5980);
nor U8429 (N_8429,N_7050,N_6938);
nand U8430 (N_8430,N_6555,N_7202);
and U8431 (N_8431,N_5405,N_6226);
and U8432 (N_8432,N_5601,N_5917);
xnor U8433 (N_8433,N_5815,N_7201);
and U8434 (N_8434,N_5819,N_5526);
or U8435 (N_8435,N_5329,N_5754);
and U8436 (N_8436,N_6200,N_7005);
or U8437 (N_8437,N_5648,N_5049);
and U8438 (N_8438,N_5276,N_5255);
nor U8439 (N_8439,N_6265,N_7254);
nand U8440 (N_8440,N_7443,N_6359);
or U8441 (N_8441,N_5079,N_6096);
nand U8442 (N_8442,N_6049,N_5779);
and U8443 (N_8443,N_5590,N_6662);
nand U8444 (N_8444,N_7355,N_5232);
or U8445 (N_8445,N_7085,N_5285);
nand U8446 (N_8446,N_6307,N_6154);
and U8447 (N_8447,N_7253,N_6960);
xnor U8448 (N_8448,N_6859,N_7007);
and U8449 (N_8449,N_6090,N_6331);
nand U8450 (N_8450,N_5240,N_5881);
or U8451 (N_8451,N_5192,N_5922);
nand U8452 (N_8452,N_5280,N_6582);
and U8453 (N_8453,N_6026,N_5297);
nor U8454 (N_8454,N_5259,N_5151);
and U8455 (N_8455,N_7116,N_6040);
xor U8456 (N_8456,N_5829,N_5764);
or U8457 (N_8457,N_6972,N_6811);
and U8458 (N_8458,N_5675,N_5472);
and U8459 (N_8459,N_6679,N_7045);
nor U8460 (N_8460,N_5215,N_7476);
nand U8461 (N_8461,N_6903,N_6974);
or U8462 (N_8462,N_5983,N_7098);
or U8463 (N_8463,N_7131,N_5399);
and U8464 (N_8464,N_6858,N_6351);
nand U8465 (N_8465,N_6922,N_5162);
nor U8466 (N_8466,N_7457,N_6031);
nand U8467 (N_8467,N_6224,N_6476);
and U8468 (N_8468,N_5641,N_6699);
or U8469 (N_8469,N_5976,N_6864);
nand U8470 (N_8470,N_6773,N_6807);
and U8471 (N_8471,N_5751,N_6770);
or U8472 (N_8472,N_7138,N_6373);
or U8473 (N_8473,N_6957,N_6389);
and U8474 (N_8474,N_5746,N_5191);
nand U8475 (N_8475,N_5871,N_5115);
nand U8476 (N_8476,N_6108,N_5470);
nand U8477 (N_8477,N_5670,N_6689);
nand U8478 (N_8478,N_5203,N_5089);
nand U8479 (N_8479,N_7299,N_5281);
nor U8480 (N_8480,N_5502,N_7168);
and U8481 (N_8481,N_6101,N_7469);
nor U8482 (N_8482,N_7250,N_5230);
nor U8483 (N_8483,N_6573,N_5415);
nor U8484 (N_8484,N_5788,N_6052);
or U8485 (N_8485,N_6801,N_5139);
or U8486 (N_8486,N_5129,N_5831);
or U8487 (N_8487,N_5564,N_6113);
and U8488 (N_8488,N_7260,N_7483);
xor U8489 (N_8489,N_6234,N_6053);
or U8490 (N_8490,N_6918,N_6374);
or U8491 (N_8491,N_6166,N_6272);
or U8492 (N_8492,N_6109,N_7464);
nand U8493 (N_8493,N_5636,N_5858);
nand U8494 (N_8494,N_5294,N_5925);
nor U8495 (N_8495,N_6311,N_7080);
or U8496 (N_8496,N_7087,N_5508);
or U8497 (N_8497,N_5649,N_7381);
or U8498 (N_8498,N_6183,N_6944);
nor U8499 (N_8499,N_5141,N_7210);
or U8500 (N_8500,N_7215,N_7319);
or U8501 (N_8501,N_6757,N_6252);
nand U8502 (N_8502,N_7150,N_5614);
or U8503 (N_8503,N_6986,N_6263);
and U8504 (N_8504,N_7153,N_6489);
nand U8505 (N_8505,N_6365,N_6750);
or U8506 (N_8506,N_6175,N_6526);
and U8507 (N_8507,N_6915,N_6132);
nor U8508 (N_8508,N_7439,N_6391);
or U8509 (N_8509,N_7218,N_6235);
or U8510 (N_8510,N_6653,N_7233);
and U8511 (N_8511,N_6994,N_6984);
nor U8512 (N_8512,N_7494,N_6013);
and U8513 (N_8513,N_6598,N_5248);
nor U8514 (N_8514,N_5393,N_6030);
nor U8515 (N_8515,N_6629,N_6386);
nand U8516 (N_8516,N_6380,N_5274);
or U8517 (N_8517,N_5824,N_6081);
nor U8518 (N_8518,N_5610,N_5154);
nand U8519 (N_8519,N_6454,N_5142);
nand U8520 (N_8520,N_6595,N_6989);
nand U8521 (N_8521,N_6114,N_6760);
nand U8522 (N_8522,N_5119,N_6208);
nand U8523 (N_8523,N_5579,N_5768);
and U8524 (N_8524,N_6578,N_5209);
and U8525 (N_8525,N_5225,N_6645);
xor U8526 (N_8526,N_5499,N_5550);
xnor U8527 (N_8527,N_7123,N_6176);
nand U8528 (N_8528,N_7338,N_5841);
xor U8529 (N_8529,N_5553,N_6403);
or U8530 (N_8530,N_6254,N_6776);
and U8531 (N_8531,N_6055,N_5452);
nor U8532 (N_8532,N_5305,N_7482);
nand U8533 (N_8533,N_7183,N_7016);
or U8534 (N_8534,N_6382,N_7242);
nand U8535 (N_8535,N_6087,N_5324);
nand U8536 (N_8536,N_5318,N_7318);
nand U8537 (N_8537,N_5837,N_5378);
nand U8538 (N_8538,N_6850,N_6843);
nor U8539 (N_8539,N_6711,N_6822);
or U8540 (N_8540,N_7198,N_7415);
and U8541 (N_8541,N_6867,N_5333);
or U8542 (N_8542,N_6592,N_6433);
xnor U8543 (N_8543,N_7396,N_5974);
or U8544 (N_8544,N_5548,N_6219);
nand U8545 (N_8545,N_7126,N_6095);
nand U8546 (N_8546,N_7365,N_6483);
nor U8547 (N_8547,N_5099,N_6806);
and U8548 (N_8548,N_7445,N_5763);
or U8549 (N_8549,N_5522,N_5501);
nor U8550 (N_8550,N_5004,N_5407);
and U8551 (N_8551,N_6144,N_6412);
nor U8552 (N_8552,N_6845,N_5016);
or U8553 (N_8553,N_6214,N_6728);
or U8554 (N_8554,N_6626,N_5953);
xnor U8555 (N_8555,N_5388,N_5105);
or U8556 (N_8556,N_7086,N_7108);
nor U8557 (N_8557,N_6761,N_6590);
and U8558 (N_8558,N_7256,N_6434);
nor U8559 (N_8559,N_7038,N_6611);
nand U8560 (N_8560,N_6658,N_5589);
or U8561 (N_8561,N_6355,N_6266);
xnor U8562 (N_8562,N_7031,N_6223);
or U8563 (N_8563,N_6923,N_6377);
and U8564 (N_8564,N_7389,N_5130);
or U8565 (N_8565,N_6148,N_7460);
xor U8566 (N_8566,N_6232,N_5028);
nand U8567 (N_8567,N_7173,N_6515);
and U8568 (N_8568,N_6499,N_7314);
nor U8569 (N_8569,N_6691,N_6591);
or U8570 (N_8570,N_6725,N_6593);
or U8571 (N_8571,N_6963,N_5095);
xor U8572 (N_8572,N_7028,N_5177);
and U8573 (N_8573,N_5169,N_5337);
and U8574 (N_8574,N_6783,N_7018);
nor U8575 (N_8575,N_5665,N_5072);
and U8576 (N_8576,N_6063,N_5566);
nand U8577 (N_8577,N_5290,N_7290);
or U8578 (N_8578,N_5206,N_7134);
or U8579 (N_8579,N_6258,N_6074);
nand U8580 (N_8580,N_5497,N_5001);
and U8581 (N_8581,N_5241,N_7191);
or U8582 (N_8582,N_6045,N_7496);
and U8583 (N_8583,N_5688,N_5799);
and U8584 (N_8584,N_5859,N_6668);
xor U8585 (N_8585,N_7337,N_6003);
and U8586 (N_8586,N_6781,N_5100);
and U8587 (N_8587,N_6622,N_6361);
xor U8588 (N_8588,N_5368,N_5460);
nor U8589 (N_8589,N_7046,N_6570);
nor U8590 (N_8590,N_6077,N_5086);
or U8591 (N_8591,N_7156,N_5900);
and U8592 (N_8592,N_6563,N_6580);
or U8593 (N_8593,N_7316,N_6171);
nand U8594 (N_8594,N_6704,N_7244);
xor U8595 (N_8595,N_6490,N_5849);
nor U8596 (N_8596,N_6405,N_5918);
nor U8597 (N_8597,N_6759,N_6149);
and U8598 (N_8598,N_5056,N_6268);
nor U8599 (N_8599,N_6333,N_7077);
and U8600 (N_8600,N_6748,N_5890);
or U8601 (N_8601,N_5145,N_7211);
nor U8602 (N_8602,N_5716,N_6105);
or U8603 (N_8603,N_7458,N_5973);
nand U8604 (N_8604,N_6933,N_5323);
and U8605 (N_8605,N_5887,N_5015);
xor U8606 (N_8606,N_5563,N_7438);
nor U8607 (N_8607,N_5693,N_6514);
nand U8608 (N_8608,N_5759,N_7397);
and U8609 (N_8609,N_7357,N_7402);
xor U8610 (N_8610,N_5428,N_6059);
nand U8611 (N_8611,N_7333,N_7213);
nand U8612 (N_8612,N_5945,N_5978);
nor U8613 (N_8613,N_6098,N_6145);
nand U8614 (N_8614,N_6253,N_6927);
or U8615 (N_8615,N_5335,N_6163);
or U8616 (N_8616,N_5876,N_5960);
nor U8617 (N_8617,N_5966,N_6969);
and U8618 (N_8618,N_5121,N_5891);
nand U8619 (N_8619,N_5410,N_6795);
and U8620 (N_8620,N_6508,N_5361);
nand U8621 (N_8621,N_5910,N_6623);
nor U8622 (N_8622,N_7370,N_5291);
xnor U8623 (N_8623,N_7158,N_6395);
nand U8624 (N_8624,N_7130,N_5443);
nor U8625 (N_8625,N_5672,N_5880);
nor U8626 (N_8626,N_5152,N_6816);
and U8627 (N_8627,N_7192,N_5351);
nor U8628 (N_8628,N_5283,N_6484);
and U8629 (N_8629,N_7128,N_7342);
nor U8630 (N_8630,N_6435,N_6250);
nor U8631 (N_8631,N_7484,N_7328);
nand U8632 (N_8632,N_6500,N_5273);
and U8633 (N_8633,N_6872,N_6681);
or U8634 (N_8634,N_5362,N_5270);
xor U8635 (N_8635,N_6893,N_5439);
nand U8636 (N_8636,N_6849,N_6665);
xor U8637 (N_8637,N_5356,N_5565);
and U8638 (N_8638,N_6277,N_6970);
nand U8639 (N_8639,N_5621,N_5613);
and U8640 (N_8640,N_7478,N_6295);
nor U8641 (N_8641,N_6871,N_6352);
or U8642 (N_8642,N_7146,N_6261);
nand U8643 (N_8643,N_7207,N_5190);
nand U8644 (N_8644,N_6425,N_6010);
or U8645 (N_8645,N_6950,N_5731);
nand U8646 (N_8646,N_6976,N_6428);
and U8647 (N_8647,N_6885,N_7133);
and U8648 (N_8648,N_7064,N_6115);
or U8649 (N_8649,N_7345,N_6086);
nand U8650 (N_8650,N_7136,N_5465);
and U8651 (N_8651,N_7239,N_7364);
xor U8652 (N_8652,N_5777,N_6853);
and U8653 (N_8653,N_7227,N_7162);
or U8654 (N_8654,N_5406,N_6958);
and U8655 (N_8655,N_6060,N_6280);
or U8656 (N_8656,N_6097,N_7095);
nand U8657 (N_8657,N_6752,N_5101);
nand U8658 (N_8658,N_6123,N_5950);
xor U8659 (N_8659,N_6606,N_6449);
and U8660 (N_8660,N_6000,N_6378);
or U8661 (N_8661,N_5586,N_6882);
and U8662 (N_8662,N_6851,N_7206);
and U8663 (N_8663,N_6227,N_7307);
or U8664 (N_8664,N_7051,N_5932);
and U8665 (N_8665,N_6571,N_5709);
nor U8666 (N_8666,N_7474,N_6988);
and U8667 (N_8667,N_6140,N_6084);
and U8668 (N_8668,N_5756,N_6564);
and U8669 (N_8669,N_5689,N_5792);
nand U8670 (N_8670,N_6397,N_6162);
nor U8671 (N_8671,N_6164,N_5705);
and U8672 (N_8672,N_6786,N_7266);
and U8673 (N_8673,N_5520,N_5737);
nand U8674 (N_8674,N_6553,N_7076);
nand U8675 (N_8675,N_6672,N_7208);
nor U8676 (N_8676,N_7032,N_7270);
or U8677 (N_8677,N_5702,N_5534);
or U8678 (N_8678,N_5639,N_5364);
and U8679 (N_8679,N_5036,N_7184);
and U8680 (N_8680,N_6203,N_6834);
nand U8681 (N_8681,N_5293,N_6856);
xnor U8682 (N_8682,N_5421,N_7155);
nor U8683 (N_8683,N_6396,N_7449);
or U8684 (N_8684,N_6409,N_6968);
and U8685 (N_8685,N_7110,N_7040);
nor U8686 (N_8686,N_7105,N_5042);
nand U8687 (N_8687,N_5624,N_6673);
or U8688 (N_8688,N_5836,N_6450);
or U8689 (N_8689,N_5827,N_6058);
nor U8690 (N_8690,N_6143,N_5657);
xor U8691 (N_8691,N_7021,N_6562);
or U8692 (N_8692,N_7297,N_7216);
and U8693 (N_8693,N_6064,N_5126);
nand U8694 (N_8694,N_6271,N_6596);
xor U8695 (N_8695,N_6241,N_7030);
and U8696 (N_8696,N_6566,N_7343);
and U8697 (N_8697,N_7352,N_5221);
nand U8698 (N_8698,N_5568,N_5561);
or U8699 (N_8699,N_6367,N_7014);
or U8700 (N_8700,N_6666,N_5208);
and U8701 (N_8701,N_5261,N_5529);
or U8702 (N_8702,N_7310,N_5690);
or U8703 (N_8703,N_6457,N_6966);
and U8704 (N_8704,N_5398,N_6706);
or U8705 (N_8705,N_6229,N_5964);
xor U8706 (N_8706,N_5866,N_5477);
nand U8707 (N_8707,N_7113,N_6478);
and U8708 (N_8708,N_5213,N_5216);
nand U8709 (N_8709,N_7093,N_6983);
and U8710 (N_8710,N_5810,N_5899);
or U8711 (N_8711,N_5157,N_7237);
and U8712 (N_8712,N_5753,N_5710);
nand U8713 (N_8713,N_7101,N_6568);
or U8714 (N_8714,N_5242,N_5638);
and U8715 (N_8715,N_7258,N_5066);
nor U8716 (N_8716,N_6462,N_7419);
and U8717 (N_8717,N_6293,N_5846);
nor U8718 (N_8718,N_7353,N_5671);
or U8719 (N_8719,N_7125,N_6170);
or U8720 (N_8720,N_7390,N_6682);
nor U8721 (N_8721,N_6513,N_5786);
and U8722 (N_8722,N_5541,N_5749);
xnor U8723 (N_8723,N_6504,N_5719);
or U8724 (N_8724,N_6601,N_5602);
or U8725 (N_8725,N_5607,N_5423);
and U8726 (N_8726,N_5412,N_6104);
nand U8727 (N_8727,N_5959,N_6037);
xnor U8728 (N_8728,N_5574,N_6376);
and U8729 (N_8729,N_6282,N_6416);
and U8730 (N_8730,N_6751,N_5595);
or U8731 (N_8731,N_7137,N_7409);
or U8732 (N_8732,N_6072,N_7444);
nor U8733 (N_8733,N_5662,N_5420);
nand U8734 (N_8734,N_5633,N_6292);
or U8735 (N_8735,N_6210,N_5050);
nor U8736 (N_8736,N_7320,N_5321);
and U8737 (N_8737,N_5780,N_7225);
or U8738 (N_8738,N_6044,N_5496);
or U8739 (N_8739,N_5391,N_7022);
nor U8740 (N_8740,N_5389,N_6195);
nand U8741 (N_8741,N_5316,N_7463);
nand U8742 (N_8742,N_5374,N_6956);
xnor U8743 (N_8743,N_7315,N_6038);
nor U8744 (N_8744,N_5408,N_6487);
nor U8745 (N_8745,N_5774,N_5969);
nor U8746 (N_8746,N_6191,N_5839);
or U8747 (N_8747,N_7043,N_6687);
and U8748 (N_8748,N_6122,N_5687);
and U8749 (N_8749,N_6846,N_6841);
nor U8750 (N_8750,N_5514,N_6058);
nor U8751 (N_8751,N_7442,N_6564);
or U8752 (N_8752,N_7087,N_6058);
nor U8753 (N_8753,N_7347,N_6535);
nand U8754 (N_8754,N_6682,N_6598);
or U8755 (N_8755,N_6692,N_6589);
xnor U8756 (N_8756,N_5337,N_5728);
and U8757 (N_8757,N_6758,N_6196);
or U8758 (N_8758,N_7254,N_6979);
or U8759 (N_8759,N_5234,N_6568);
nor U8760 (N_8760,N_5373,N_7177);
nor U8761 (N_8761,N_6626,N_6407);
xor U8762 (N_8762,N_5966,N_7032);
nand U8763 (N_8763,N_7098,N_6410);
and U8764 (N_8764,N_5087,N_6682);
nor U8765 (N_8765,N_6846,N_6875);
nor U8766 (N_8766,N_5377,N_7385);
nand U8767 (N_8767,N_5782,N_7024);
or U8768 (N_8768,N_7301,N_5691);
and U8769 (N_8769,N_5681,N_6990);
or U8770 (N_8770,N_5107,N_7068);
and U8771 (N_8771,N_7118,N_6344);
or U8772 (N_8772,N_7436,N_7495);
nand U8773 (N_8773,N_6828,N_5541);
nor U8774 (N_8774,N_7431,N_5489);
nand U8775 (N_8775,N_5374,N_5599);
nand U8776 (N_8776,N_5791,N_6971);
or U8777 (N_8777,N_5287,N_5994);
nand U8778 (N_8778,N_6455,N_5024);
or U8779 (N_8779,N_5252,N_5396);
nand U8780 (N_8780,N_5991,N_5622);
and U8781 (N_8781,N_5659,N_5841);
and U8782 (N_8782,N_5392,N_5009);
or U8783 (N_8783,N_5156,N_6231);
nand U8784 (N_8784,N_5958,N_6727);
or U8785 (N_8785,N_5594,N_5986);
nand U8786 (N_8786,N_7094,N_5798);
or U8787 (N_8787,N_5034,N_6228);
xnor U8788 (N_8788,N_5569,N_7245);
nor U8789 (N_8789,N_5554,N_5341);
and U8790 (N_8790,N_6212,N_5618);
or U8791 (N_8791,N_5510,N_5722);
xnor U8792 (N_8792,N_6150,N_7398);
or U8793 (N_8793,N_6245,N_6681);
nand U8794 (N_8794,N_5100,N_5707);
or U8795 (N_8795,N_6825,N_6189);
or U8796 (N_8796,N_5808,N_6143);
and U8797 (N_8797,N_7313,N_5382);
nand U8798 (N_8798,N_5160,N_5022);
and U8799 (N_8799,N_5778,N_5048);
nor U8800 (N_8800,N_5222,N_7043);
nand U8801 (N_8801,N_7476,N_7387);
nor U8802 (N_8802,N_6439,N_5735);
or U8803 (N_8803,N_6423,N_6712);
or U8804 (N_8804,N_6024,N_6262);
nor U8805 (N_8805,N_6818,N_7036);
nand U8806 (N_8806,N_6834,N_6430);
or U8807 (N_8807,N_7469,N_5149);
and U8808 (N_8808,N_6063,N_6081);
xor U8809 (N_8809,N_5238,N_7194);
and U8810 (N_8810,N_6670,N_5069);
or U8811 (N_8811,N_6831,N_5491);
nor U8812 (N_8812,N_7232,N_6633);
nor U8813 (N_8813,N_5567,N_5336);
nor U8814 (N_8814,N_5304,N_6539);
or U8815 (N_8815,N_5321,N_6135);
and U8816 (N_8816,N_7015,N_5173);
and U8817 (N_8817,N_5807,N_6600);
nand U8818 (N_8818,N_5163,N_7215);
or U8819 (N_8819,N_5232,N_5370);
or U8820 (N_8820,N_5696,N_7497);
or U8821 (N_8821,N_7165,N_5762);
and U8822 (N_8822,N_6271,N_7083);
nor U8823 (N_8823,N_5872,N_5662);
nor U8824 (N_8824,N_6763,N_6249);
or U8825 (N_8825,N_6326,N_7097);
nand U8826 (N_8826,N_5862,N_7198);
nand U8827 (N_8827,N_5525,N_5591);
and U8828 (N_8828,N_6521,N_6861);
xnor U8829 (N_8829,N_5042,N_7400);
and U8830 (N_8830,N_6055,N_6145);
nand U8831 (N_8831,N_6600,N_6191);
nand U8832 (N_8832,N_5400,N_6443);
nand U8833 (N_8833,N_7314,N_7433);
xnor U8834 (N_8834,N_5246,N_6557);
or U8835 (N_8835,N_5101,N_5142);
or U8836 (N_8836,N_6754,N_5406);
nand U8837 (N_8837,N_5661,N_6027);
and U8838 (N_8838,N_6059,N_6373);
nor U8839 (N_8839,N_7194,N_6816);
nand U8840 (N_8840,N_5252,N_7327);
nand U8841 (N_8841,N_5715,N_5433);
or U8842 (N_8842,N_6769,N_5668);
or U8843 (N_8843,N_5370,N_7359);
or U8844 (N_8844,N_7146,N_5411);
nor U8845 (N_8845,N_6452,N_7362);
and U8846 (N_8846,N_6494,N_6221);
and U8847 (N_8847,N_6569,N_6269);
or U8848 (N_8848,N_5625,N_5622);
nor U8849 (N_8849,N_6233,N_6500);
and U8850 (N_8850,N_7105,N_5169);
and U8851 (N_8851,N_6576,N_7188);
xnor U8852 (N_8852,N_7493,N_6176);
nor U8853 (N_8853,N_5383,N_5809);
xor U8854 (N_8854,N_5876,N_5669);
or U8855 (N_8855,N_6138,N_7230);
xor U8856 (N_8856,N_5048,N_6477);
or U8857 (N_8857,N_7145,N_5536);
nand U8858 (N_8858,N_5708,N_5915);
and U8859 (N_8859,N_6082,N_7133);
xor U8860 (N_8860,N_6974,N_5592);
nor U8861 (N_8861,N_7000,N_5834);
and U8862 (N_8862,N_6794,N_5981);
nand U8863 (N_8863,N_5007,N_6158);
xnor U8864 (N_8864,N_6902,N_5055);
and U8865 (N_8865,N_5716,N_5959);
and U8866 (N_8866,N_6514,N_5928);
xor U8867 (N_8867,N_7264,N_5123);
xor U8868 (N_8868,N_5067,N_6252);
nor U8869 (N_8869,N_7488,N_7396);
or U8870 (N_8870,N_6336,N_5843);
nor U8871 (N_8871,N_5486,N_5312);
nand U8872 (N_8872,N_7342,N_6003);
nor U8873 (N_8873,N_6242,N_6305);
and U8874 (N_8874,N_6209,N_6337);
nand U8875 (N_8875,N_7225,N_7058);
and U8876 (N_8876,N_5980,N_6855);
nor U8877 (N_8877,N_6769,N_6723);
or U8878 (N_8878,N_6716,N_5365);
nand U8879 (N_8879,N_7008,N_6809);
nor U8880 (N_8880,N_6902,N_5380);
nor U8881 (N_8881,N_5971,N_5395);
and U8882 (N_8882,N_7092,N_5106);
and U8883 (N_8883,N_6601,N_6305);
or U8884 (N_8884,N_6025,N_5239);
nor U8885 (N_8885,N_6347,N_5787);
xor U8886 (N_8886,N_7010,N_6504);
or U8887 (N_8887,N_6907,N_6971);
or U8888 (N_8888,N_7371,N_5957);
and U8889 (N_8889,N_5321,N_6830);
or U8890 (N_8890,N_5862,N_6080);
or U8891 (N_8891,N_5729,N_5378);
nor U8892 (N_8892,N_5995,N_5773);
or U8893 (N_8893,N_5683,N_6142);
and U8894 (N_8894,N_6790,N_5849);
nor U8895 (N_8895,N_5964,N_6715);
and U8896 (N_8896,N_5670,N_7492);
and U8897 (N_8897,N_6741,N_6374);
and U8898 (N_8898,N_6885,N_5075);
or U8899 (N_8899,N_5745,N_5487);
or U8900 (N_8900,N_6926,N_6409);
and U8901 (N_8901,N_5466,N_5686);
nand U8902 (N_8902,N_5157,N_6299);
or U8903 (N_8903,N_7492,N_5777);
nand U8904 (N_8904,N_5311,N_7219);
and U8905 (N_8905,N_6312,N_6820);
nand U8906 (N_8906,N_7481,N_6988);
nand U8907 (N_8907,N_6099,N_7303);
and U8908 (N_8908,N_6883,N_7336);
xor U8909 (N_8909,N_7204,N_6925);
nand U8910 (N_8910,N_6253,N_5445);
nand U8911 (N_8911,N_6079,N_7166);
xnor U8912 (N_8912,N_6041,N_6253);
nand U8913 (N_8913,N_5721,N_6182);
nand U8914 (N_8914,N_6533,N_5920);
and U8915 (N_8915,N_6625,N_5298);
and U8916 (N_8916,N_5023,N_5826);
and U8917 (N_8917,N_6671,N_5033);
nor U8918 (N_8918,N_5785,N_5199);
and U8919 (N_8919,N_6247,N_5708);
and U8920 (N_8920,N_6025,N_5520);
xnor U8921 (N_8921,N_5014,N_6898);
nor U8922 (N_8922,N_6575,N_7427);
nor U8923 (N_8923,N_6439,N_6301);
xnor U8924 (N_8924,N_6246,N_6349);
and U8925 (N_8925,N_7136,N_5032);
nor U8926 (N_8926,N_5703,N_6257);
nand U8927 (N_8927,N_5461,N_6801);
nand U8928 (N_8928,N_6077,N_5459);
or U8929 (N_8929,N_5562,N_6131);
and U8930 (N_8930,N_7359,N_5929);
xnor U8931 (N_8931,N_6571,N_7044);
or U8932 (N_8932,N_5911,N_5447);
nor U8933 (N_8933,N_6007,N_6881);
xnor U8934 (N_8934,N_5418,N_7431);
xor U8935 (N_8935,N_5468,N_6173);
or U8936 (N_8936,N_5420,N_6389);
or U8937 (N_8937,N_6719,N_5063);
and U8938 (N_8938,N_5853,N_7369);
nand U8939 (N_8939,N_5660,N_7018);
nor U8940 (N_8940,N_5911,N_5908);
nor U8941 (N_8941,N_5649,N_6109);
or U8942 (N_8942,N_6682,N_5230);
and U8943 (N_8943,N_7028,N_7286);
nand U8944 (N_8944,N_5590,N_5747);
xor U8945 (N_8945,N_5452,N_6513);
xnor U8946 (N_8946,N_5426,N_5497);
nand U8947 (N_8947,N_5662,N_5811);
or U8948 (N_8948,N_6624,N_5548);
nor U8949 (N_8949,N_6379,N_5875);
nand U8950 (N_8950,N_5034,N_5230);
or U8951 (N_8951,N_5919,N_6055);
nor U8952 (N_8952,N_6110,N_5683);
or U8953 (N_8953,N_6943,N_6708);
nor U8954 (N_8954,N_5234,N_5681);
and U8955 (N_8955,N_6096,N_5755);
and U8956 (N_8956,N_5897,N_6955);
nand U8957 (N_8957,N_6099,N_6220);
nor U8958 (N_8958,N_5239,N_7112);
xor U8959 (N_8959,N_5586,N_5173);
xnor U8960 (N_8960,N_6342,N_5210);
nand U8961 (N_8961,N_7266,N_5178);
or U8962 (N_8962,N_7094,N_7134);
nand U8963 (N_8963,N_7064,N_5164);
nand U8964 (N_8964,N_5096,N_5734);
nor U8965 (N_8965,N_6947,N_6990);
nand U8966 (N_8966,N_5767,N_5750);
nor U8967 (N_8967,N_6496,N_6277);
nor U8968 (N_8968,N_7002,N_5665);
nor U8969 (N_8969,N_5397,N_5272);
xor U8970 (N_8970,N_6004,N_5193);
or U8971 (N_8971,N_5772,N_6318);
nor U8972 (N_8972,N_5693,N_5183);
and U8973 (N_8973,N_6199,N_6345);
nor U8974 (N_8974,N_5653,N_6273);
nor U8975 (N_8975,N_7135,N_5282);
or U8976 (N_8976,N_7222,N_7291);
nand U8977 (N_8977,N_5028,N_7345);
or U8978 (N_8978,N_7099,N_7068);
nand U8979 (N_8979,N_6024,N_6243);
nand U8980 (N_8980,N_7284,N_5355);
or U8981 (N_8981,N_5800,N_5534);
and U8982 (N_8982,N_6006,N_6810);
nand U8983 (N_8983,N_6671,N_6153);
and U8984 (N_8984,N_6516,N_5827);
and U8985 (N_8985,N_7202,N_7252);
xnor U8986 (N_8986,N_6168,N_7406);
or U8987 (N_8987,N_7091,N_5675);
nor U8988 (N_8988,N_6400,N_7199);
xor U8989 (N_8989,N_5848,N_7425);
nand U8990 (N_8990,N_5007,N_5725);
or U8991 (N_8991,N_6723,N_5385);
nor U8992 (N_8992,N_6530,N_5107);
nor U8993 (N_8993,N_6424,N_5596);
xnor U8994 (N_8994,N_5974,N_5836);
nand U8995 (N_8995,N_6280,N_5920);
nor U8996 (N_8996,N_5520,N_5874);
nand U8997 (N_8997,N_7403,N_6750);
or U8998 (N_8998,N_7026,N_6493);
and U8999 (N_8999,N_6244,N_5793);
nand U9000 (N_9000,N_7408,N_5616);
and U9001 (N_9001,N_5761,N_5574);
nand U9002 (N_9002,N_5318,N_5719);
nand U9003 (N_9003,N_5886,N_6864);
and U9004 (N_9004,N_5819,N_5773);
and U9005 (N_9005,N_7292,N_6384);
xor U9006 (N_9006,N_6529,N_5063);
nor U9007 (N_9007,N_5212,N_7010);
nand U9008 (N_9008,N_5652,N_5624);
or U9009 (N_9009,N_6890,N_6813);
or U9010 (N_9010,N_5162,N_6790);
or U9011 (N_9011,N_5248,N_6323);
and U9012 (N_9012,N_6544,N_7023);
or U9013 (N_9013,N_6730,N_7073);
xnor U9014 (N_9014,N_6980,N_5709);
and U9015 (N_9015,N_6242,N_7229);
nor U9016 (N_9016,N_5688,N_7073);
xor U9017 (N_9017,N_5027,N_6887);
nor U9018 (N_9018,N_6706,N_7038);
or U9019 (N_9019,N_5183,N_6388);
nand U9020 (N_9020,N_7447,N_5341);
or U9021 (N_9021,N_6480,N_5491);
or U9022 (N_9022,N_6223,N_7321);
or U9023 (N_9023,N_7442,N_5220);
nor U9024 (N_9024,N_5514,N_5656);
or U9025 (N_9025,N_5727,N_5181);
and U9026 (N_9026,N_7419,N_5851);
nand U9027 (N_9027,N_7493,N_7342);
or U9028 (N_9028,N_5505,N_5331);
xnor U9029 (N_9029,N_7198,N_5713);
nor U9030 (N_9030,N_6908,N_5330);
nor U9031 (N_9031,N_7202,N_6605);
nor U9032 (N_9032,N_7428,N_5091);
and U9033 (N_9033,N_6733,N_5090);
and U9034 (N_9034,N_6269,N_7070);
and U9035 (N_9035,N_6377,N_7109);
nand U9036 (N_9036,N_6932,N_7436);
nand U9037 (N_9037,N_5032,N_6281);
and U9038 (N_9038,N_7259,N_7485);
nor U9039 (N_9039,N_7139,N_7454);
or U9040 (N_9040,N_6074,N_6505);
nor U9041 (N_9041,N_5084,N_6899);
or U9042 (N_9042,N_6539,N_6050);
or U9043 (N_9043,N_5441,N_5628);
nor U9044 (N_9044,N_6737,N_5847);
xnor U9045 (N_9045,N_5227,N_7409);
and U9046 (N_9046,N_6574,N_5679);
nor U9047 (N_9047,N_6163,N_6126);
or U9048 (N_9048,N_6759,N_7241);
and U9049 (N_9049,N_7102,N_5321);
and U9050 (N_9050,N_6277,N_7020);
nor U9051 (N_9051,N_6628,N_7018);
nor U9052 (N_9052,N_7184,N_6950);
and U9053 (N_9053,N_7429,N_6326);
nand U9054 (N_9054,N_7164,N_7369);
nor U9055 (N_9055,N_5445,N_5574);
nor U9056 (N_9056,N_7400,N_6262);
or U9057 (N_9057,N_6144,N_6746);
nor U9058 (N_9058,N_5326,N_5703);
xor U9059 (N_9059,N_6467,N_6983);
nor U9060 (N_9060,N_6017,N_5594);
and U9061 (N_9061,N_6773,N_6542);
and U9062 (N_9062,N_5218,N_6107);
nor U9063 (N_9063,N_5821,N_5945);
or U9064 (N_9064,N_7493,N_6469);
and U9065 (N_9065,N_7173,N_6471);
and U9066 (N_9066,N_5673,N_6247);
nor U9067 (N_9067,N_5726,N_7202);
nand U9068 (N_9068,N_5715,N_6316);
nand U9069 (N_9069,N_5810,N_6663);
xor U9070 (N_9070,N_6059,N_6493);
and U9071 (N_9071,N_6797,N_6376);
nand U9072 (N_9072,N_5668,N_6446);
or U9073 (N_9073,N_5883,N_6039);
or U9074 (N_9074,N_7188,N_6814);
nand U9075 (N_9075,N_6797,N_6295);
nor U9076 (N_9076,N_7302,N_7321);
nor U9077 (N_9077,N_6223,N_6506);
nor U9078 (N_9078,N_6631,N_7046);
and U9079 (N_9079,N_5354,N_5730);
or U9080 (N_9080,N_5894,N_6383);
nand U9081 (N_9081,N_5839,N_6295);
or U9082 (N_9082,N_5154,N_5511);
or U9083 (N_9083,N_6341,N_5930);
xor U9084 (N_9084,N_6442,N_5275);
and U9085 (N_9085,N_7158,N_5344);
or U9086 (N_9086,N_5251,N_6589);
and U9087 (N_9087,N_5412,N_6575);
or U9088 (N_9088,N_6146,N_6771);
nor U9089 (N_9089,N_5406,N_6994);
nor U9090 (N_9090,N_5807,N_5515);
nand U9091 (N_9091,N_6557,N_7389);
nand U9092 (N_9092,N_5567,N_7069);
and U9093 (N_9093,N_5058,N_5380);
nand U9094 (N_9094,N_6846,N_7078);
and U9095 (N_9095,N_5630,N_6405);
and U9096 (N_9096,N_5188,N_5610);
nor U9097 (N_9097,N_7102,N_6943);
xor U9098 (N_9098,N_6399,N_5576);
xor U9099 (N_9099,N_6772,N_6429);
nand U9100 (N_9100,N_5658,N_5925);
xnor U9101 (N_9101,N_6269,N_5507);
nand U9102 (N_9102,N_5125,N_6665);
nor U9103 (N_9103,N_6815,N_6337);
nor U9104 (N_9104,N_5734,N_6017);
xnor U9105 (N_9105,N_7091,N_6835);
and U9106 (N_9106,N_5511,N_6750);
or U9107 (N_9107,N_7489,N_7341);
nand U9108 (N_9108,N_6759,N_5997);
nand U9109 (N_9109,N_6516,N_7496);
or U9110 (N_9110,N_7067,N_6321);
nor U9111 (N_9111,N_6144,N_6324);
nor U9112 (N_9112,N_5059,N_6853);
and U9113 (N_9113,N_6239,N_6423);
nand U9114 (N_9114,N_5038,N_5443);
or U9115 (N_9115,N_7157,N_6927);
or U9116 (N_9116,N_5968,N_7268);
nor U9117 (N_9117,N_6962,N_6900);
nor U9118 (N_9118,N_5281,N_6048);
nor U9119 (N_9119,N_6370,N_5108);
and U9120 (N_9120,N_6659,N_6122);
nor U9121 (N_9121,N_6625,N_5793);
nand U9122 (N_9122,N_5699,N_5516);
and U9123 (N_9123,N_7188,N_6786);
nor U9124 (N_9124,N_7040,N_5986);
nor U9125 (N_9125,N_5055,N_7301);
xnor U9126 (N_9126,N_6881,N_7148);
and U9127 (N_9127,N_6957,N_5058);
or U9128 (N_9128,N_6729,N_5743);
nor U9129 (N_9129,N_5260,N_5493);
nor U9130 (N_9130,N_7181,N_7384);
nor U9131 (N_9131,N_5158,N_5434);
xor U9132 (N_9132,N_6679,N_6064);
nand U9133 (N_9133,N_5867,N_6555);
nand U9134 (N_9134,N_7380,N_6383);
and U9135 (N_9135,N_5023,N_5830);
nor U9136 (N_9136,N_5107,N_6283);
and U9137 (N_9137,N_5804,N_7085);
nor U9138 (N_9138,N_5103,N_6591);
or U9139 (N_9139,N_6265,N_5321);
nand U9140 (N_9140,N_5049,N_7353);
nand U9141 (N_9141,N_7331,N_5295);
or U9142 (N_9142,N_6803,N_5950);
nor U9143 (N_9143,N_6004,N_7126);
or U9144 (N_9144,N_7329,N_7363);
nor U9145 (N_9145,N_7009,N_5592);
or U9146 (N_9146,N_5675,N_7323);
nand U9147 (N_9147,N_5876,N_7235);
xnor U9148 (N_9148,N_6546,N_7136);
or U9149 (N_9149,N_7392,N_5580);
nand U9150 (N_9150,N_6093,N_5403);
and U9151 (N_9151,N_6056,N_6531);
and U9152 (N_9152,N_7496,N_5604);
and U9153 (N_9153,N_5096,N_6311);
or U9154 (N_9154,N_6026,N_5388);
nor U9155 (N_9155,N_6802,N_6885);
xnor U9156 (N_9156,N_5568,N_6630);
nor U9157 (N_9157,N_5161,N_7387);
nor U9158 (N_9158,N_5212,N_5265);
and U9159 (N_9159,N_6202,N_6063);
nor U9160 (N_9160,N_5942,N_6765);
nor U9161 (N_9161,N_5721,N_6537);
nor U9162 (N_9162,N_6823,N_5104);
nor U9163 (N_9163,N_5499,N_5837);
nand U9164 (N_9164,N_5012,N_7086);
and U9165 (N_9165,N_6763,N_5424);
or U9166 (N_9166,N_6884,N_5641);
nand U9167 (N_9167,N_6886,N_5163);
or U9168 (N_9168,N_7362,N_6779);
nor U9169 (N_9169,N_7218,N_7304);
nor U9170 (N_9170,N_7149,N_6823);
and U9171 (N_9171,N_6464,N_6364);
or U9172 (N_9172,N_6434,N_6441);
and U9173 (N_9173,N_5265,N_6841);
nor U9174 (N_9174,N_6430,N_7446);
and U9175 (N_9175,N_5699,N_6193);
and U9176 (N_9176,N_5054,N_5111);
or U9177 (N_9177,N_7276,N_7169);
nor U9178 (N_9178,N_5233,N_6230);
or U9179 (N_9179,N_5360,N_7452);
and U9180 (N_9180,N_5668,N_6892);
or U9181 (N_9181,N_6021,N_7325);
or U9182 (N_9182,N_5777,N_5445);
nor U9183 (N_9183,N_6419,N_6264);
or U9184 (N_9184,N_5573,N_5806);
or U9185 (N_9185,N_6364,N_6765);
nand U9186 (N_9186,N_7088,N_6303);
nor U9187 (N_9187,N_5316,N_5140);
and U9188 (N_9188,N_6855,N_5488);
or U9189 (N_9189,N_5328,N_6132);
and U9190 (N_9190,N_6572,N_7219);
nand U9191 (N_9191,N_5947,N_6510);
and U9192 (N_9192,N_6773,N_7340);
nor U9193 (N_9193,N_6497,N_6070);
or U9194 (N_9194,N_6748,N_6250);
and U9195 (N_9195,N_7298,N_5511);
and U9196 (N_9196,N_6526,N_7147);
xnor U9197 (N_9197,N_5239,N_5889);
nand U9198 (N_9198,N_6684,N_7378);
or U9199 (N_9199,N_5154,N_6064);
or U9200 (N_9200,N_6907,N_7497);
nor U9201 (N_9201,N_5923,N_6637);
nand U9202 (N_9202,N_6917,N_6256);
nor U9203 (N_9203,N_6614,N_7482);
or U9204 (N_9204,N_5318,N_6631);
and U9205 (N_9205,N_7325,N_7095);
nand U9206 (N_9206,N_6164,N_6836);
xor U9207 (N_9207,N_7374,N_7315);
or U9208 (N_9208,N_6076,N_5574);
and U9209 (N_9209,N_6232,N_6833);
and U9210 (N_9210,N_6727,N_7331);
nand U9211 (N_9211,N_5963,N_6904);
nand U9212 (N_9212,N_6722,N_7459);
nand U9213 (N_9213,N_6894,N_6474);
and U9214 (N_9214,N_5836,N_7201);
or U9215 (N_9215,N_7330,N_7004);
or U9216 (N_9216,N_5872,N_6334);
nand U9217 (N_9217,N_6878,N_5238);
and U9218 (N_9218,N_5450,N_6479);
and U9219 (N_9219,N_6274,N_6833);
and U9220 (N_9220,N_5483,N_5845);
or U9221 (N_9221,N_7214,N_7002);
and U9222 (N_9222,N_6657,N_6502);
or U9223 (N_9223,N_5663,N_6027);
xor U9224 (N_9224,N_6114,N_6716);
or U9225 (N_9225,N_5070,N_6764);
or U9226 (N_9226,N_6135,N_6284);
nand U9227 (N_9227,N_5878,N_7084);
nand U9228 (N_9228,N_5771,N_7141);
or U9229 (N_9229,N_6865,N_7483);
and U9230 (N_9230,N_7196,N_5064);
or U9231 (N_9231,N_5805,N_6577);
nor U9232 (N_9232,N_6278,N_6071);
or U9233 (N_9233,N_7054,N_5657);
and U9234 (N_9234,N_6988,N_6559);
nor U9235 (N_9235,N_5762,N_6844);
or U9236 (N_9236,N_5270,N_5698);
nor U9237 (N_9237,N_5578,N_7302);
nor U9238 (N_9238,N_7259,N_5974);
nand U9239 (N_9239,N_5030,N_5697);
or U9240 (N_9240,N_7315,N_6394);
and U9241 (N_9241,N_7333,N_7114);
or U9242 (N_9242,N_6964,N_5226);
nor U9243 (N_9243,N_6725,N_6996);
and U9244 (N_9244,N_6856,N_6832);
nor U9245 (N_9245,N_6593,N_7027);
or U9246 (N_9246,N_5651,N_6426);
or U9247 (N_9247,N_6074,N_7061);
nand U9248 (N_9248,N_7190,N_5775);
and U9249 (N_9249,N_6700,N_5915);
or U9250 (N_9250,N_6987,N_6086);
nand U9251 (N_9251,N_6032,N_7172);
nand U9252 (N_9252,N_6918,N_6467);
or U9253 (N_9253,N_5798,N_6584);
and U9254 (N_9254,N_5695,N_6515);
nor U9255 (N_9255,N_6994,N_6119);
nand U9256 (N_9256,N_6985,N_6514);
nand U9257 (N_9257,N_6557,N_7252);
nand U9258 (N_9258,N_7396,N_7331);
or U9259 (N_9259,N_5868,N_6592);
xor U9260 (N_9260,N_6494,N_6814);
and U9261 (N_9261,N_6999,N_6324);
or U9262 (N_9262,N_6038,N_5086);
and U9263 (N_9263,N_5089,N_7166);
and U9264 (N_9264,N_6650,N_5729);
or U9265 (N_9265,N_6917,N_5349);
and U9266 (N_9266,N_7242,N_6100);
or U9267 (N_9267,N_5749,N_6568);
nand U9268 (N_9268,N_6977,N_5643);
nand U9269 (N_9269,N_5316,N_6818);
and U9270 (N_9270,N_5289,N_5463);
and U9271 (N_9271,N_6103,N_6252);
or U9272 (N_9272,N_6162,N_5340);
nand U9273 (N_9273,N_5735,N_5818);
xor U9274 (N_9274,N_6686,N_6895);
and U9275 (N_9275,N_6701,N_5332);
or U9276 (N_9276,N_6610,N_5108);
xnor U9277 (N_9277,N_6360,N_5912);
nor U9278 (N_9278,N_5505,N_6782);
nor U9279 (N_9279,N_7421,N_6629);
nor U9280 (N_9280,N_6437,N_5183);
xnor U9281 (N_9281,N_7297,N_7409);
or U9282 (N_9282,N_5372,N_7444);
and U9283 (N_9283,N_5081,N_7470);
nor U9284 (N_9284,N_6714,N_6037);
xor U9285 (N_9285,N_5885,N_5339);
and U9286 (N_9286,N_6541,N_7093);
xor U9287 (N_9287,N_7048,N_5522);
nor U9288 (N_9288,N_5119,N_5555);
xor U9289 (N_9289,N_5408,N_5949);
and U9290 (N_9290,N_6145,N_5499);
and U9291 (N_9291,N_6795,N_5414);
or U9292 (N_9292,N_7285,N_5786);
nand U9293 (N_9293,N_5498,N_7072);
nand U9294 (N_9294,N_7086,N_6553);
and U9295 (N_9295,N_6652,N_5217);
or U9296 (N_9296,N_5873,N_6101);
nor U9297 (N_9297,N_6540,N_6561);
nand U9298 (N_9298,N_5330,N_6203);
xnor U9299 (N_9299,N_7304,N_6520);
nand U9300 (N_9300,N_5751,N_6365);
nand U9301 (N_9301,N_6757,N_5546);
and U9302 (N_9302,N_6650,N_5908);
nand U9303 (N_9303,N_5959,N_5938);
and U9304 (N_9304,N_5047,N_5864);
or U9305 (N_9305,N_5309,N_5174);
and U9306 (N_9306,N_5002,N_5911);
and U9307 (N_9307,N_6818,N_6390);
or U9308 (N_9308,N_5034,N_7442);
nor U9309 (N_9309,N_6525,N_7399);
nor U9310 (N_9310,N_5476,N_5956);
or U9311 (N_9311,N_5477,N_6321);
nand U9312 (N_9312,N_5763,N_6682);
and U9313 (N_9313,N_6029,N_6160);
or U9314 (N_9314,N_6768,N_6130);
nor U9315 (N_9315,N_5700,N_5318);
nor U9316 (N_9316,N_6467,N_6940);
and U9317 (N_9317,N_6211,N_6612);
and U9318 (N_9318,N_5892,N_5068);
nor U9319 (N_9319,N_6337,N_6982);
nand U9320 (N_9320,N_5759,N_7380);
or U9321 (N_9321,N_7492,N_5196);
nand U9322 (N_9322,N_5656,N_5585);
or U9323 (N_9323,N_7258,N_7314);
and U9324 (N_9324,N_7016,N_7288);
and U9325 (N_9325,N_6102,N_6680);
nor U9326 (N_9326,N_5234,N_6381);
nand U9327 (N_9327,N_7306,N_6803);
and U9328 (N_9328,N_7406,N_6163);
nand U9329 (N_9329,N_6849,N_5040);
or U9330 (N_9330,N_5495,N_7408);
nand U9331 (N_9331,N_5990,N_6920);
nor U9332 (N_9332,N_5255,N_6048);
or U9333 (N_9333,N_6246,N_6564);
and U9334 (N_9334,N_6203,N_7109);
or U9335 (N_9335,N_7481,N_6354);
nor U9336 (N_9336,N_6483,N_6297);
nand U9337 (N_9337,N_6206,N_5161);
nand U9338 (N_9338,N_5060,N_6047);
nor U9339 (N_9339,N_6212,N_5669);
nor U9340 (N_9340,N_7193,N_5570);
and U9341 (N_9341,N_7090,N_6233);
nand U9342 (N_9342,N_6555,N_5083);
nor U9343 (N_9343,N_5214,N_5267);
and U9344 (N_9344,N_5204,N_5734);
and U9345 (N_9345,N_6168,N_5526);
and U9346 (N_9346,N_6386,N_7134);
nor U9347 (N_9347,N_6628,N_5868);
nor U9348 (N_9348,N_5747,N_6333);
nand U9349 (N_9349,N_7080,N_6182);
or U9350 (N_9350,N_7309,N_7454);
and U9351 (N_9351,N_5702,N_7003);
and U9352 (N_9352,N_6521,N_7395);
or U9353 (N_9353,N_6023,N_6298);
and U9354 (N_9354,N_5195,N_5047);
nand U9355 (N_9355,N_5078,N_5385);
xnor U9356 (N_9356,N_7117,N_5767);
or U9357 (N_9357,N_5985,N_5526);
nor U9358 (N_9358,N_5716,N_6886);
xor U9359 (N_9359,N_6106,N_5079);
nor U9360 (N_9360,N_6573,N_6036);
and U9361 (N_9361,N_5977,N_7087);
xor U9362 (N_9362,N_5702,N_6865);
and U9363 (N_9363,N_6152,N_7295);
nor U9364 (N_9364,N_6689,N_6074);
and U9365 (N_9365,N_6105,N_7111);
nand U9366 (N_9366,N_6283,N_5953);
nor U9367 (N_9367,N_5367,N_6243);
and U9368 (N_9368,N_6931,N_6328);
and U9369 (N_9369,N_6000,N_6326);
nor U9370 (N_9370,N_7350,N_6809);
and U9371 (N_9371,N_5667,N_6555);
nand U9372 (N_9372,N_5050,N_5653);
or U9373 (N_9373,N_5919,N_5821);
nand U9374 (N_9374,N_5959,N_5076);
nand U9375 (N_9375,N_7281,N_6489);
nand U9376 (N_9376,N_6996,N_5721);
nor U9377 (N_9377,N_7210,N_6703);
xor U9378 (N_9378,N_7253,N_7270);
nor U9379 (N_9379,N_6847,N_6822);
or U9380 (N_9380,N_5106,N_5615);
and U9381 (N_9381,N_6872,N_7374);
xor U9382 (N_9382,N_6372,N_5302);
or U9383 (N_9383,N_7008,N_5599);
and U9384 (N_9384,N_5627,N_7206);
nor U9385 (N_9385,N_5015,N_6923);
or U9386 (N_9386,N_6382,N_6676);
xor U9387 (N_9387,N_5086,N_6284);
xor U9388 (N_9388,N_5252,N_5253);
or U9389 (N_9389,N_7067,N_5441);
and U9390 (N_9390,N_7180,N_7412);
or U9391 (N_9391,N_6777,N_7356);
or U9392 (N_9392,N_7042,N_6407);
and U9393 (N_9393,N_6464,N_6571);
and U9394 (N_9394,N_7030,N_5363);
or U9395 (N_9395,N_6679,N_7282);
nand U9396 (N_9396,N_7012,N_5797);
or U9397 (N_9397,N_6177,N_6216);
and U9398 (N_9398,N_7381,N_6545);
nor U9399 (N_9399,N_6248,N_5803);
nor U9400 (N_9400,N_5722,N_6037);
and U9401 (N_9401,N_5634,N_7435);
nand U9402 (N_9402,N_6557,N_5264);
or U9403 (N_9403,N_5354,N_7004);
or U9404 (N_9404,N_6096,N_5302);
or U9405 (N_9405,N_6320,N_5028);
or U9406 (N_9406,N_5734,N_6799);
nand U9407 (N_9407,N_5374,N_5063);
and U9408 (N_9408,N_6444,N_7402);
and U9409 (N_9409,N_5919,N_6500);
nor U9410 (N_9410,N_6032,N_5066);
or U9411 (N_9411,N_6843,N_6285);
and U9412 (N_9412,N_5643,N_6540);
or U9413 (N_9413,N_5919,N_5308);
nand U9414 (N_9414,N_7246,N_6143);
or U9415 (N_9415,N_7450,N_5532);
nor U9416 (N_9416,N_6808,N_5978);
nor U9417 (N_9417,N_7184,N_6188);
nand U9418 (N_9418,N_6370,N_6705);
nor U9419 (N_9419,N_6071,N_5487);
or U9420 (N_9420,N_6586,N_6990);
or U9421 (N_9421,N_6278,N_6102);
and U9422 (N_9422,N_6399,N_6481);
nand U9423 (N_9423,N_6765,N_6773);
nand U9424 (N_9424,N_5663,N_5755);
nand U9425 (N_9425,N_6914,N_7344);
or U9426 (N_9426,N_5407,N_6309);
and U9427 (N_9427,N_6379,N_6828);
or U9428 (N_9428,N_6021,N_5543);
and U9429 (N_9429,N_6682,N_5469);
nor U9430 (N_9430,N_5192,N_6112);
nor U9431 (N_9431,N_5906,N_5141);
nor U9432 (N_9432,N_5027,N_7403);
nand U9433 (N_9433,N_6604,N_7485);
nand U9434 (N_9434,N_6227,N_5223);
or U9435 (N_9435,N_5577,N_7371);
nand U9436 (N_9436,N_6477,N_6268);
nor U9437 (N_9437,N_7135,N_7281);
and U9438 (N_9438,N_6441,N_7210);
or U9439 (N_9439,N_5904,N_5609);
or U9440 (N_9440,N_5370,N_6418);
and U9441 (N_9441,N_6969,N_6701);
nand U9442 (N_9442,N_7348,N_6269);
or U9443 (N_9443,N_6937,N_5149);
or U9444 (N_9444,N_7410,N_5317);
nor U9445 (N_9445,N_6429,N_5672);
or U9446 (N_9446,N_5452,N_6629);
and U9447 (N_9447,N_7183,N_7362);
nand U9448 (N_9448,N_5826,N_5312);
and U9449 (N_9449,N_6552,N_7160);
and U9450 (N_9450,N_6550,N_6409);
or U9451 (N_9451,N_5396,N_5882);
or U9452 (N_9452,N_7481,N_6662);
and U9453 (N_9453,N_7433,N_7375);
nor U9454 (N_9454,N_7293,N_6323);
and U9455 (N_9455,N_6193,N_6288);
and U9456 (N_9456,N_5213,N_7439);
and U9457 (N_9457,N_6726,N_5241);
or U9458 (N_9458,N_7349,N_6378);
nor U9459 (N_9459,N_6980,N_6104);
or U9460 (N_9460,N_5408,N_7243);
nor U9461 (N_9461,N_5982,N_5184);
nor U9462 (N_9462,N_5121,N_5338);
xnor U9463 (N_9463,N_6612,N_6993);
nor U9464 (N_9464,N_7192,N_5667);
or U9465 (N_9465,N_5395,N_5343);
and U9466 (N_9466,N_5838,N_5135);
nand U9467 (N_9467,N_6190,N_6295);
nand U9468 (N_9468,N_5835,N_7441);
and U9469 (N_9469,N_6627,N_6066);
nand U9470 (N_9470,N_5854,N_7244);
xnor U9471 (N_9471,N_6364,N_5472);
nor U9472 (N_9472,N_6870,N_6752);
or U9473 (N_9473,N_6307,N_5561);
and U9474 (N_9474,N_6284,N_6775);
nand U9475 (N_9475,N_5078,N_7067);
nor U9476 (N_9476,N_5638,N_5467);
nand U9477 (N_9477,N_5279,N_7313);
nand U9478 (N_9478,N_6324,N_5682);
nor U9479 (N_9479,N_5285,N_7424);
xnor U9480 (N_9480,N_6334,N_7373);
xor U9481 (N_9481,N_5840,N_5405);
nor U9482 (N_9482,N_6476,N_6660);
nor U9483 (N_9483,N_7020,N_5430);
or U9484 (N_9484,N_7450,N_6922);
and U9485 (N_9485,N_5999,N_6113);
and U9486 (N_9486,N_6391,N_6396);
and U9487 (N_9487,N_7188,N_7465);
and U9488 (N_9488,N_6247,N_5691);
nand U9489 (N_9489,N_6950,N_5002);
xor U9490 (N_9490,N_5992,N_5194);
and U9491 (N_9491,N_7091,N_7452);
nand U9492 (N_9492,N_5709,N_5465);
and U9493 (N_9493,N_5964,N_6512);
nand U9494 (N_9494,N_5766,N_6320);
xor U9495 (N_9495,N_6291,N_5832);
and U9496 (N_9496,N_6862,N_7102);
nand U9497 (N_9497,N_7184,N_6612);
nor U9498 (N_9498,N_6861,N_7063);
nor U9499 (N_9499,N_7172,N_5407);
nand U9500 (N_9500,N_5711,N_7414);
or U9501 (N_9501,N_5697,N_7329);
or U9502 (N_9502,N_5198,N_5971);
or U9503 (N_9503,N_5575,N_6358);
or U9504 (N_9504,N_5018,N_7225);
nor U9505 (N_9505,N_6126,N_6204);
nor U9506 (N_9506,N_5480,N_7475);
nand U9507 (N_9507,N_5918,N_6801);
nand U9508 (N_9508,N_7015,N_7065);
and U9509 (N_9509,N_6353,N_6378);
and U9510 (N_9510,N_5015,N_6180);
nor U9511 (N_9511,N_7158,N_5177);
nand U9512 (N_9512,N_7269,N_5237);
and U9513 (N_9513,N_6341,N_6467);
and U9514 (N_9514,N_5864,N_6252);
nor U9515 (N_9515,N_7486,N_7039);
or U9516 (N_9516,N_5863,N_5308);
and U9517 (N_9517,N_6843,N_7355);
nand U9518 (N_9518,N_7417,N_5989);
and U9519 (N_9519,N_7348,N_7114);
nand U9520 (N_9520,N_7082,N_5076);
nand U9521 (N_9521,N_5169,N_7476);
nor U9522 (N_9522,N_6544,N_5698);
and U9523 (N_9523,N_6609,N_6258);
and U9524 (N_9524,N_5143,N_5460);
nand U9525 (N_9525,N_6285,N_5504);
or U9526 (N_9526,N_7405,N_7146);
nand U9527 (N_9527,N_6232,N_5683);
nor U9528 (N_9528,N_6577,N_6655);
or U9529 (N_9529,N_5587,N_5250);
nor U9530 (N_9530,N_6251,N_5442);
nor U9531 (N_9531,N_6271,N_6411);
nor U9532 (N_9532,N_5554,N_6812);
xor U9533 (N_9533,N_5988,N_6782);
nand U9534 (N_9534,N_6821,N_5508);
nor U9535 (N_9535,N_6570,N_7051);
or U9536 (N_9536,N_5815,N_5132);
xor U9537 (N_9537,N_6636,N_7362);
xnor U9538 (N_9538,N_7470,N_6138);
nand U9539 (N_9539,N_5600,N_6335);
or U9540 (N_9540,N_5700,N_5290);
or U9541 (N_9541,N_5222,N_7471);
nand U9542 (N_9542,N_5250,N_5330);
or U9543 (N_9543,N_6017,N_7491);
and U9544 (N_9544,N_6958,N_7332);
or U9545 (N_9545,N_6527,N_6707);
nor U9546 (N_9546,N_6781,N_7318);
xor U9547 (N_9547,N_7312,N_6409);
or U9548 (N_9548,N_6083,N_7198);
or U9549 (N_9549,N_5491,N_6486);
nor U9550 (N_9550,N_5251,N_7278);
or U9551 (N_9551,N_6065,N_6120);
and U9552 (N_9552,N_5919,N_6816);
nor U9553 (N_9553,N_6336,N_7378);
nand U9554 (N_9554,N_5706,N_6606);
nor U9555 (N_9555,N_7112,N_6683);
and U9556 (N_9556,N_7382,N_7490);
nor U9557 (N_9557,N_6600,N_7402);
or U9558 (N_9558,N_5876,N_6088);
nand U9559 (N_9559,N_6569,N_6434);
nand U9560 (N_9560,N_6599,N_5075);
or U9561 (N_9561,N_6852,N_6568);
nor U9562 (N_9562,N_5444,N_6413);
or U9563 (N_9563,N_5124,N_7290);
nand U9564 (N_9564,N_5726,N_7312);
nand U9565 (N_9565,N_6007,N_6002);
xor U9566 (N_9566,N_6162,N_5931);
or U9567 (N_9567,N_5987,N_7333);
nand U9568 (N_9568,N_6410,N_5737);
nand U9569 (N_9569,N_7172,N_5734);
or U9570 (N_9570,N_5359,N_5619);
nand U9571 (N_9571,N_5341,N_6421);
and U9572 (N_9572,N_6006,N_7092);
or U9573 (N_9573,N_7080,N_6149);
nor U9574 (N_9574,N_6810,N_6707);
nor U9575 (N_9575,N_6724,N_6866);
and U9576 (N_9576,N_5727,N_5342);
nand U9577 (N_9577,N_5456,N_5360);
and U9578 (N_9578,N_6617,N_6232);
or U9579 (N_9579,N_7494,N_6463);
nand U9580 (N_9580,N_6938,N_6469);
xnor U9581 (N_9581,N_7363,N_5388);
or U9582 (N_9582,N_5745,N_7226);
nand U9583 (N_9583,N_5700,N_5982);
or U9584 (N_9584,N_6765,N_6923);
and U9585 (N_9585,N_7130,N_5433);
xor U9586 (N_9586,N_6009,N_5972);
nand U9587 (N_9587,N_6356,N_6721);
xnor U9588 (N_9588,N_6320,N_7440);
nand U9589 (N_9589,N_6973,N_5492);
nor U9590 (N_9590,N_6386,N_7206);
nor U9591 (N_9591,N_6705,N_6859);
nor U9592 (N_9592,N_6933,N_6582);
nor U9593 (N_9593,N_6583,N_5663);
and U9594 (N_9594,N_5308,N_6123);
or U9595 (N_9595,N_5208,N_6139);
and U9596 (N_9596,N_6086,N_5467);
nor U9597 (N_9597,N_6264,N_5376);
nand U9598 (N_9598,N_5014,N_5896);
nand U9599 (N_9599,N_7495,N_5646);
nor U9600 (N_9600,N_7316,N_7229);
nand U9601 (N_9601,N_5457,N_5885);
and U9602 (N_9602,N_5340,N_7430);
nor U9603 (N_9603,N_5466,N_5256);
nor U9604 (N_9604,N_6106,N_5761);
xnor U9605 (N_9605,N_5120,N_7240);
or U9606 (N_9606,N_5127,N_5541);
nor U9607 (N_9607,N_7260,N_5679);
nor U9608 (N_9608,N_6030,N_5079);
or U9609 (N_9609,N_6975,N_5096);
nor U9610 (N_9610,N_7380,N_7166);
nand U9611 (N_9611,N_6912,N_5462);
and U9612 (N_9612,N_5371,N_7472);
or U9613 (N_9613,N_5830,N_6970);
nand U9614 (N_9614,N_5295,N_5537);
nand U9615 (N_9615,N_7168,N_7183);
or U9616 (N_9616,N_6834,N_7185);
and U9617 (N_9617,N_5809,N_5883);
and U9618 (N_9618,N_6713,N_6069);
or U9619 (N_9619,N_5125,N_7444);
nor U9620 (N_9620,N_5158,N_6602);
xor U9621 (N_9621,N_7056,N_7406);
nor U9622 (N_9622,N_6808,N_7095);
or U9623 (N_9623,N_6533,N_5390);
xor U9624 (N_9624,N_5042,N_7466);
nor U9625 (N_9625,N_5178,N_5188);
and U9626 (N_9626,N_5120,N_7319);
or U9627 (N_9627,N_5947,N_7040);
and U9628 (N_9628,N_7053,N_5946);
and U9629 (N_9629,N_5990,N_6770);
nand U9630 (N_9630,N_5725,N_5142);
nor U9631 (N_9631,N_7025,N_5444);
xnor U9632 (N_9632,N_5385,N_6452);
nor U9633 (N_9633,N_6406,N_5386);
nand U9634 (N_9634,N_5256,N_5126);
nor U9635 (N_9635,N_5313,N_6452);
nand U9636 (N_9636,N_7380,N_7125);
nand U9637 (N_9637,N_7365,N_7282);
nor U9638 (N_9638,N_7389,N_6898);
or U9639 (N_9639,N_5415,N_7191);
or U9640 (N_9640,N_7020,N_7151);
nand U9641 (N_9641,N_5575,N_5772);
or U9642 (N_9642,N_6605,N_7145);
and U9643 (N_9643,N_7340,N_7272);
xor U9644 (N_9644,N_5408,N_5393);
nor U9645 (N_9645,N_5006,N_5773);
and U9646 (N_9646,N_7351,N_7484);
nand U9647 (N_9647,N_7486,N_6285);
or U9648 (N_9648,N_7044,N_6256);
nor U9649 (N_9649,N_6853,N_5801);
or U9650 (N_9650,N_7247,N_5965);
and U9651 (N_9651,N_5344,N_5446);
nor U9652 (N_9652,N_7321,N_6697);
or U9653 (N_9653,N_5016,N_7177);
nand U9654 (N_9654,N_7376,N_5810);
nand U9655 (N_9655,N_5536,N_6441);
or U9656 (N_9656,N_6518,N_5177);
nand U9657 (N_9657,N_6282,N_6759);
or U9658 (N_9658,N_6286,N_7102);
or U9659 (N_9659,N_7206,N_6862);
and U9660 (N_9660,N_5656,N_6355);
and U9661 (N_9661,N_5188,N_6837);
and U9662 (N_9662,N_5906,N_6190);
or U9663 (N_9663,N_6416,N_7261);
or U9664 (N_9664,N_5159,N_6819);
and U9665 (N_9665,N_5654,N_7106);
and U9666 (N_9666,N_5464,N_6888);
nor U9667 (N_9667,N_7309,N_7427);
or U9668 (N_9668,N_6582,N_5759);
xnor U9669 (N_9669,N_5993,N_7064);
and U9670 (N_9670,N_5766,N_5150);
nor U9671 (N_9671,N_7485,N_6656);
nand U9672 (N_9672,N_6736,N_6945);
or U9673 (N_9673,N_6472,N_6864);
or U9674 (N_9674,N_7469,N_5292);
or U9675 (N_9675,N_6994,N_6211);
and U9676 (N_9676,N_6538,N_7375);
nand U9677 (N_9677,N_7421,N_6056);
or U9678 (N_9678,N_5837,N_5272);
and U9679 (N_9679,N_5127,N_5849);
or U9680 (N_9680,N_5143,N_6590);
nor U9681 (N_9681,N_5823,N_6676);
nand U9682 (N_9682,N_6163,N_5653);
nor U9683 (N_9683,N_7416,N_7271);
and U9684 (N_9684,N_6339,N_5435);
xor U9685 (N_9685,N_6220,N_5222);
nor U9686 (N_9686,N_5438,N_6140);
or U9687 (N_9687,N_7074,N_7070);
or U9688 (N_9688,N_7263,N_5569);
or U9689 (N_9689,N_5771,N_7369);
nor U9690 (N_9690,N_6807,N_5091);
or U9691 (N_9691,N_6547,N_6760);
xnor U9692 (N_9692,N_5551,N_7008);
or U9693 (N_9693,N_5478,N_5195);
xnor U9694 (N_9694,N_6843,N_5466);
nor U9695 (N_9695,N_5830,N_7101);
or U9696 (N_9696,N_5044,N_6063);
nor U9697 (N_9697,N_5634,N_5297);
or U9698 (N_9698,N_5026,N_6211);
nand U9699 (N_9699,N_6158,N_6217);
or U9700 (N_9700,N_6861,N_7065);
nand U9701 (N_9701,N_5659,N_7193);
and U9702 (N_9702,N_5805,N_6883);
and U9703 (N_9703,N_6737,N_5636);
xnor U9704 (N_9704,N_5619,N_5111);
or U9705 (N_9705,N_7375,N_7308);
xor U9706 (N_9706,N_5408,N_7145);
or U9707 (N_9707,N_5322,N_5246);
or U9708 (N_9708,N_6783,N_6929);
or U9709 (N_9709,N_6090,N_6951);
xor U9710 (N_9710,N_6758,N_6998);
or U9711 (N_9711,N_5958,N_6392);
or U9712 (N_9712,N_6437,N_6304);
nand U9713 (N_9713,N_6263,N_6441);
nor U9714 (N_9714,N_5488,N_6005);
and U9715 (N_9715,N_5601,N_6225);
and U9716 (N_9716,N_6744,N_6655);
and U9717 (N_9717,N_5677,N_7437);
and U9718 (N_9718,N_6610,N_5611);
nand U9719 (N_9719,N_6387,N_5288);
xor U9720 (N_9720,N_7088,N_6787);
or U9721 (N_9721,N_5559,N_7471);
nor U9722 (N_9722,N_5470,N_6986);
nand U9723 (N_9723,N_7052,N_6502);
nand U9724 (N_9724,N_7276,N_7386);
and U9725 (N_9725,N_5285,N_6114);
or U9726 (N_9726,N_6898,N_6006);
nand U9727 (N_9727,N_6150,N_6442);
nor U9728 (N_9728,N_6132,N_7127);
nand U9729 (N_9729,N_5543,N_7288);
and U9730 (N_9730,N_6919,N_5913);
nand U9731 (N_9731,N_6711,N_5231);
or U9732 (N_9732,N_5370,N_7364);
nor U9733 (N_9733,N_6968,N_5255);
nor U9734 (N_9734,N_7485,N_6919);
nand U9735 (N_9735,N_5058,N_6663);
nand U9736 (N_9736,N_6247,N_6322);
or U9737 (N_9737,N_7056,N_6447);
nand U9738 (N_9738,N_7465,N_7304);
and U9739 (N_9739,N_7108,N_5775);
and U9740 (N_9740,N_6385,N_5356);
nor U9741 (N_9741,N_5826,N_6652);
nor U9742 (N_9742,N_6396,N_6060);
nand U9743 (N_9743,N_6560,N_6746);
nand U9744 (N_9744,N_6962,N_7441);
nand U9745 (N_9745,N_6922,N_5420);
and U9746 (N_9746,N_5738,N_5384);
and U9747 (N_9747,N_5030,N_5601);
nand U9748 (N_9748,N_6659,N_6394);
nor U9749 (N_9749,N_5481,N_6982);
nor U9750 (N_9750,N_5722,N_5717);
nand U9751 (N_9751,N_5499,N_6172);
nand U9752 (N_9752,N_7072,N_6098);
nand U9753 (N_9753,N_6649,N_6129);
xnor U9754 (N_9754,N_6782,N_5865);
or U9755 (N_9755,N_5791,N_6382);
xor U9756 (N_9756,N_6013,N_7386);
nand U9757 (N_9757,N_7199,N_6754);
and U9758 (N_9758,N_5050,N_7369);
nand U9759 (N_9759,N_6886,N_7476);
nand U9760 (N_9760,N_7312,N_5714);
nand U9761 (N_9761,N_7353,N_6940);
or U9762 (N_9762,N_6675,N_6953);
nor U9763 (N_9763,N_7409,N_6527);
nand U9764 (N_9764,N_6425,N_6194);
nand U9765 (N_9765,N_6587,N_7224);
or U9766 (N_9766,N_6513,N_5892);
nor U9767 (N_9767,N_5313,N_5462);
nor U9768 (N_9768,N_6584,N_6170);
nor U9769 (N_9769,N_5592,N_5706);
nor U9770 (N_9770,N_6267,N_6946);
and U9771 (N_9771,N_7038,N_6031);
and U9772 (N_9772,N_6713,N_7241);
nor U9773 (N_9773,N_7487,N_5545);
or U9774 (N_9774,N_6427,N_7109);
or U9775 (N_9775,N_6763,N_5106);
and U9776 (N_9776,N_7053,N_7266);
xnor U9777 (N_9777,N_7235,N_6083);
and U9778 (N_9778,N_7303,N_5230);
and U9779 (N_9779,N_5084,N_6438);
nand U9780 (N_9780,N_6389,N_5677);
nor U9781 (N_9781,N_6744,N_5782);
or U9782 (N_9782,N_5219,N_5828);
or U9783 (N_9783,N_5111,N_5341);
or U9784 (N_9784,N_5637,N_6564);
and U9785 (N_9785,N_6596,N_6228);
or U9786 (N_9786,N_5978,N_5531);
and U9787 (N_9787,N_7407,N_6253);
nor U9788 (N_9788,N_6168,N_5222);
nor U9789 (N_9789,N_7049,N_7118);
nor U9790 (N_9790,N_5665,N_5256);
and U9791 (N_9791,N_7458,N_5063);
nor U9792 (N_9792,N_7426,N_5091);
and U9793 (N_9793,N_6632,N_6021);
and U9794 (N_9794,N_5541,N_7474);
nand U9795 (N_9795,N_6275,N_6198);
nor U9796 (N_9796,N_5796,N_5497);
nor U9797 (N_9797,N_5961,N_5000);
nand U9798 (N_9798,N_6411,N_7457);
nand U9799 (N_9799,N_5101,N_5159);
or U9800 (N_9800,N_6228,N_7182);
or U9801 (N_9801,N_6637,N_7186);
and U9802 (N_9802,N_6272,N_5815);
or U9803 (N_9803,N_5917,N_5768);
or U9804 (N_9804,N_5201,N_6717);
nor U9805 (N_9805,N_5762,N_6673);
and U9806 (N_9806,N_6278,N_6982);
or U9807 (N_9807,N_7495,N_7421);
or U9808 (N_9808,N_5647,N_7139);
and U9809 (N_9809,N_6310,N_5385);
nand U9810 (N_9810,N_6984,N_6432);
and U9811 (N_9811,N_7401,N_5534);
or U9812 (N_9812,N_5450,N_5889);
nand U9813 (N_9813,N_6976,N_6308);
and U9814 (N_9814,N_5702,N_6337);
nand U9815 (N_9815,N_6021,N_6116);
nor U9816 (N_9816,N_6715,N_7288);
or U9817 (N_9817,N_7385,N_6196);
nor U9818 (N_9818,N_7371,N_6801);
or U9819 (N_9819,N_5979,N_6664);
or U9820 (N_9820,N_6306,N_6055);
nand U9821 (N_9821,N_6833,N_5797);
or U9822 (N_9822,N_5197,N_7084);
or U9823 (N_9823,N_5217,N_6145);
nor U9824 (N_9824,N_5180,N_5560);
or U9825 (N_9825,N_6931,N_7395);
nor U9826 (N_9826,N_6027,N_6542);
and U9827 (N_9827,N_6140,N_5726);
and U9828 (N_9828,N_5957,N_5546);
and U9829 (N_9829,N_6353,N_5367);
or U9830 (N_9830,N_7276,N_6323);
nor U9831 (N_9831,N_6268,N_6141);
xnor U9832 (N_9832,N_6971,N_7312);
nand U9833 (N_9833,N_5675,N_6014);
and U9834 (N_9834,N_6613,N_7290);
xnor U9835 (N_9835,N_6021,N_5925);
or U9836 (N_9836,N_7320,N_5290);
xnor U9837 (N_9837,N_6027,N_7115);
nand U9838 (N_9838,N_6107,N_6456);
nand U9839 (N_9839,N_7074,N_5180);
nor U9840 (N_9840,N_6345,N_6526);
or U9841 (N_9841,N_6525,N_5914);
or U9842 (N_9842,N_6138,N_6713);
nand U9843 (N_9843,N_6984,N_7150);
nor U9844 (N_9844,N_6475,N_5711);
nor U9845 (N_9845,N_6027,N_5531);
nand U9846 (N_9846,N_6241,N_5019);
nor U9847 (N_9847,N_5101,N_5723);
nor U9848 (N_9848,N_6767,N_6777);
nand U9849 (N_9849,N_5467,N_7356);
nand U9850 (N_9850,N_7348,N_5843);
and U9851 (N_9851,N_6752,N_7269);
and U9852 (N_9852,N_5759,N_6074);
nand U9853 (N_9853,N_6639,N_6062);
nand U9854 (N_9854,N_6706,N_6051);
and U9855 (N_9855,N_7393,N_5494);
nor U9856 (N_9856,N_7270,N_5240);
nand U9857 (N_9857,N_5347,N_6877);
nand U9858 (N_9858,N_5734,N_5312);
nor U9859 (N_9859,N_7251,N_5187);
nand U9860 (N_9860,N_6119,N_7391);
nand U9861 (N_9861,N_5947,N_6191);
and U9862 (N_9862,N_5112,N_5790);
and U9863 (N_9863,N_5208,N_5606);
nand U9864 (N_9864,N_6927,N_7460);
nor U9865 (N_9865,N_5700,N_6641);
nor U9866 (N_9866,N_5355,N_5137);
and U9867 (N_9867,N_5601,N_6639);
nand U9868 (N_9868,N_6984,N_5225);
and U9869 (N_9869,N_5440,N_6939);
nand U9870 (N_9870,N_6093,N_6477);
and U9871 (N_9871,N_7158,N_5167);
or U9872 (N_9872,N_5133,N_6460);
and U9873 (N_9873,N_5712,N_6295);
xor U9874 (N_9874,N_5258,N_6821);
and U9875 (N_9875,N_5223,N_7074);
xnor U9876 (N_9876,N_6853,N_5881);
nor U9877 (N_9877,N_7084,N_5136);
nor U9878 (N_9878,N_7141,N_6987);
nor U9879 (N_9879,N_6000,N_7422);
and U9880 (N_9880,N_7211,N_6740);
nor U9881 (N_9881,N_5254,N_6909);
or U9882 (N_9882,N_7436,N_7004);
and U9883 (N_9883,N_6150,N_5461);
nand U9884 (N_9884,N_6199,N_5416);
xnor U9885 (N_9885,N_6893,N_6111);
and U9886 (N_9886,N_7132,N_5487);
xor U9887 (N_9887,N_6349,N_7246);
nand U9888 (N_9888,N_6578,N_7185);
nand U9889 (N_9889,N_6719,N_5992);
nor U9890 (N_9890,N_5965,N_6246);
and U9891 (N_9891,N_6637,N_5586);
nor U9892 (N_9892,N_6651,N_5579);
nor U9893 (N_9893,N_6447,N_7258);
or U9894 (N_9894,N_5548,N_6617);
nand U9895 (N_9895,N_5452,N_6707);
or U9896 (N_9896,N_7111,N_6298);
nor U9897 (N_9897,N_5541,N_5336);
nor U9898 (N_9898,N_7320,N_6769);
nand U9899 (N_9899,N_6916,N_6539);
nand U9900 (N_9900,N_6925,N_5196);
and U9901 (N_9901,N_6705,N_6547);
nor U9902 (N_9902,N_7382,N_5089);
nor U9903 (N_9903,N_5588,N_7266);
nor U9904 (N_9904,N_7285,N_7387);
nor U9905 (N_9905,N_5998,N_5193);
and U9906 (N_9906,N_7065,N_6680);
nor U9907 (N_9907,N_5775,N_5892);
nor U9908 (N_9908,N_7328,N_5035);
nand U9909 (N_9909,N_6107,N_5124);
and U9910 (N_9910,N_6608,N_5853);
or U9911 (N_9911,N_5085,N_5473);
nor U9912 (N_9912,N_5854,N_6972);
or U9913 (N_9913,N_6461,N_5664);
and U9914 (N_9914,N_5142,N_6482);
and U9915 (N_9915,N_6971,N_7406);
or U9916 (N_9916,N_6708,N_6239);
and U9917 (N_9917,N_6003,N_5238);
xnor U9918 (N_9918,N_6574,N_6986);
nand U9919 (N_9919,N_7461,N_5370);
nor U9920 (N_9920,N_6785,N_5258);
or U9921 (N_9921,N_6133,N_6534);
or U9922 (N_9922,N_6883,N_7317);
and U9923 (N_9923,N_7406,N_6438);
nand U9924 (N_9924,N_5197,N_7066);
nor U9925 (N_9925,N_6456,N_6049);
and U9926 (N_9926,N_5579,N_7266);
or U9927 (N_9927,N_5779,N_6508);
or U9928 (N_9928,N_5881,N_7304);
nor U9929 (N_9929,N_7365,N_7487);
and U9930 (N_9930,N_6361,N_5966);
and U9931 (N_9931,N_6331,N_5824);
or U9932 (N_9932,N_7434,N_5463);
or U9933 (N_9933,N_5432,N_5398);
or U9934 (N_9934,N_6429,N_7136);
and U9935 (N_9935,N_6609,N_5633);
nand U9936 (N_9936,N_6438,N_5817);
or U9937 (N_9937,N_5943,N_6964);
and U9938 (N_9938,N_6217,N_6078);
and U9939 (N_9939,N_5375,N_6697);
nor U9940 (N_9940,N_5382,N_5388);
nand U9941 (N_9941,N_7237,N_6788);
or U9942 (N_9942,N_5016,N_6675);
nand U9943 (N_9943,N_6454,N_7169);
nor U9944 (N_9944,N_7059,N_5903);
or U9945 (N_9945,N_7416,N_6283);
nand U9946 (N_9946,N_7120,N_5482);
nand U9947 (N_9947,N_6500,N_5386);
nor U9948 (N_9948,N_5576,N_6735);
xor U9949 (N_9949,N_5255,N_5974);
and U9950 (N_9950,N_5295,N_7131);
nor U9951 (N_9951,N_5453,N_5188);
xnor U9952 (N_9952,N_6483,N_6678);
nor U9953 (N_9953,N_6638,N_7408);
xor U9954 (N_9954,N_6686,N_7131);
nand U9955 (N_9955,N_6283,N_6158);
and U9956 (N_9956,N_6093,N_6713);
nand U9957 (N_9957,N_7422,N_7272);
nor U9958 (N_9958,N_6983,N_6192);
and U9959 (N_9959,N_5702,N_5419);
or U9960 (N_9960,N_5374,N_6412);
nand U9961 (N_9961,N_5613,N_5673);
or U9962 (N_9962,N_5517,N_7219);
nor U9963 (N_9963,N_7222,N_6682);
or U9964 (N_9964,N_7121,N_6350);
or U9965 (N_9965,N_6806,N_5479);
nor U9966 (N_9966,N_7182,N_7335);
nand U9967 (N_9967,N_5943,N_5704);
and U9968 (N_9968,N_7092,N_6103);
nor U9969 (N_9969,N_6409,N_5490);
or U9970 (N_9970,N_5134,N_6550);
nor U9971 (N_9971,N_6163,N_6751);
and U9972 (N_9972,N_6852,N_5328);
nand U9973 (N_9973,N_5111,N_7356);
nand U9974 (N_9974,N_5890,N_5927);
nor U9975 (N_9975,N_7492,N_6437);
xnor U9976 (N_9976,N_7163,N_7251);
nor U9977 (N_9977,N_6227,N_5906);
or U9978 (N_9978,N_7449,N_5465);
nand U9979 (N_9979,N_6520,N_5681);
and U9980 (N_9980,N_5214,N_6750);
and U9981 (N_9981,N_5195,N_5095);
or U9982 (N_9982,N_6625,N_6517);
nand U9983 (N_9983,N_5014,N_6937);
and U9984 (N_9984,N_6411,N_5327);
or U9985 (N_9985,N_5374,N_5456);
and U9986 (N_9986,N_6623,N_6505);
nor U9987 (N_9987,N_7141,N_6035);
xnor U9988 (N_9988,N_7172,N_6484);
and U9989 (N_9989,N_6421,N_7021);
and U9990 (N_9990,N_7114,N_6017);
or U9991 (N_9991,N_6836,N_7080);
nand U9992 (N_9992,N_7254,N_6585);
and U9993 (N_9993,N_7089,N_6276);
xnor U9994 (N_9994,N_5632,N_5962);
or U9995 (N_9995,N_5333,N_5250);
nand U9996 (N_9996,N_5269,N_5731);
nor U9997 (N_9997,N_5711,N_5871);
nand U9998 (N_9998,N_6800,N_7088);
xnor U9999 (N_9999,N_6809,N_6636);
nor UO_0 (O_0,N_8998,N_8647);
nand UO_1 (O_1,N_8704,N_9896);
and UO_2 (O_2,N_9579,N_9106);
or UO_3 (O_3,N_7584,N_9646);
and UO_4 (O_4,N_7927,N_8512);
and UO_5 (O_5,N_9396,N_7746);
or UO_6 (O_6,N_9758,N_9518);
nand UO_7 (O_7,N_7656,N_7840);
nand UO_8 (O_8,N_8706,N_9122);
and UO_9 (O_9,N_9252,N_7950);
nor UO_10 (O_10,N_9617,N_8525);
or UO_11 (O_11,N_9426,N_9733);
or UO_12 (O_12,N_9317,N_9371);
and UO_13 (O_13,N_9357,N_9353);
and UO_14 (O_14,N_9476,N_8827);
and UO_15 (O_15,N_9248,N_9922);
or UO_16 (O_16,N_9236,N_8792);
nor UO_17 (O_17,N_7504,N_8769);
and UO_18 (O_18,N_8528,N_8849);
nand UO_19 (O_19,N_9993,N_7754);
xor UO_20 (O_20,N_9759,N_9227);
or UO_21 (O_21,N_8441,N_7905);
nor UO_22 (O_22,N_8289,N_8178);
nand UO_23 (O_23,N_9451,N_8136);
nand UO_24 (O_24,N_9792,N_9727);
or UO_25 (O_25,N_7995,N_7909);
xor UO_26 (O_26,N_7668,N_9002);
and UO_27 (O_27,N_8170,N_8536);
or UO_28 (O_28,N_9626,N_9682);
nand UO_29 (O_29,N_7568,N_9302);
and UO_30 (O_30,N_9103,N_8714);
and UO_31 (O_31,N_8678,N_9416);
or UO_32 (O_32,N_9114,N_8995);
nor UO_33 (O_33,N_9823,N_9508);
or UO_34 (O_34,N_7908,N_8868);
nand UO_35 (O_35,N_9315,N_7784);
and UO_36 (O_36,N_9568,N_9105);
nand UO_37 (O_37,N_8328,N_8189);
or UO_38 (O_38,N_7736,N_8060);
nor UO_39 (O_39,N_9108,N_9323);
nor UO_40 (O_40,N_7541,N_9601);
nand UO_41 (O_41,N_8372,N_9224);
or UO_42 (O_42,N_9343,N_9716);
or UO_43 (O_43,N_9936,N_9597);
and UO_44 (O_44,N_7592,N_7721);
and UO_45 (O_45,N_8495,N_9745);
and UO_46 (O_46,N_9649,N_9949);
nor UO_47 (O_47,N_8099,N_9082);
nor UO_48 (O_48,N_8883,N_8805);
and UO_49 (O_49,N_8923,N_8763);
nor UO_50 (O_50,N_7875,N_8741);
or UO_51 (O_51,N_9872,N_8325);
nor UO_52 (O_52,N_9384,N_9032);
nor UO_53 (O_53,N_9347,N_7891);
nor UO_54 (O_54,N_7884,N_9174);
nand UO_55 (O_55,N_7790,N_9209);
or UO_56 (O_56,N_8848,N_7616);
nand UO_57 (O_57,N_8267,N_9713);
nor UO_58 (O_58,N_8947,N_8568);
or UO_59 (O_59,N_7526,N_7637);
nor UO_60 (O_60,N_9030,N_8760);
or UO_61 (O_61,N_9440,N_9552);
nand UO_62 (O_62,N_9256,N_9663);
or UO_63 (O_63,N_9613,N_8789);
or UO_64 (O_64,N_7712,N_9567);
nor UO_65 (O_65,N_9586,N_8213);
xnor UO_66 (O_66,N_7855,N_9378);
nor UO_67 (O_67,N_8301,N_9427);
nor UO_68 (O_68,N_7839,N_7633);
xor UO_69 (O_69,N_8479,N_8972);
or UO_70 (O_70,N_8544,N_8830);
and UO_71 (O_71,N_8881,N_7819);
nand UO_72 (O_72,N_9888,N_7557);
nand UO_73 (O_73,N_9324,N_8237);
xor UO_74 (O_74,N_8921,N_8553);
nand UO_75 (O_75,N_9536,N_8342);
xnor UO_76 (O_76,N_9621,N_8067);
nand UO_77 (O_77,N_9830,N_9254);
and UO_78 (O_78,N_9731,N_8806);
and UO_79 (O_79,N_8380,N_8684);
or UO_80 (O_80,N_8870,N_7734);
and UO_81 (O_81,N_8280,N_9214);
nand UO_82 (O_82,N_8221,N_9944);
and UO_83 (O_83,N_8516,N_9527);
nor UO_84 (O_84,N_8724,N_7589);
and UO_85 (O_85,N_9826,N_8208);
and UO_86 (O_86,N_8906,N_8837);
xnor UO_87 (O_87,N_9756,N_9517);
nand UO_88 (O_88,N_8541,N_8680);
nor UO_89 (O_89,N_8030,N_9433);
and UO_90 (O_90,N_8540,N_9898);
or UO_91 (O_91,N_8639,N_8964);
nand UO_92 (O_92,N_8955,N_8655);
nor UO_93 (O_93,N_8413,N_9467);
xnor UO_94 (O_94,N_9177,N_9041);
xnor UO_95 (O_95,N_8375,N_9056);
or UO_96 (O_96,N_9635,N_9878);
nor UO_97 (O_97,N_8748,N_8183);
or UO_98 (O_98,N_9829,N_8510);
nor UO_99 (O_99,N_8139,N_9084);
and UO_100 (O_100,N_9837,N_9901);
and UO_101 (O_101,N_9380,N_9955);
xnor UO_102 (O_102,N_9280,N_7823);
and UO_103 (O_103,N_8043,N_8638);
nand UO_104 (O_104,N_8521,N_8599);
and UO_105 (O_105,N_9895,N_8687);
and UO_106 (O_106,N_9804,N_9331);
xor UO_107 (O_107,N_9432,N_7893);
nor UO_108 (O_108,N_8448,N_8013);
or UO_109 (O_109,N_9839,N_8659);
nand UO_110 (O_110,N_9465,N_9924);
and UO_111 (O_111,N_8108,N_7586);
nor UO_112 (O_112,N_8798,N_9329);
nor UO_113 (O_113,N_8895,N_9781);
nand UO_114 (O_114,N_7998,N_9689);
nor UO_115 (O_115,N_8594,N_7545);
and UO_116 (O_116,N_8695,N_8415);
and UO_117 (O_117,N_7755,N_9711);
or UO_118 (O_118,N_9652,N_9857);
xnor UO_119 (O_119,N_9819,N_9962);
or UO_120 (O_120,N_9454,N_8693);
and UO_121 (O_121,N_7682,N_8123);
or UO_122 (O_122,N_9395,N_8429);
and UO_123 (O_123,N_9095,N_7506);
nand UO_124 (O_124,N_9471,N_8062);
nor UO_125 (O_125,N_8344,N_7932);
nor UO_126 (O_126,N_9514,N_8036);
or UO_127 (O_127,N_9183,N_9569);
and UO_128 (O_128,N_7732,N_9428);
xnor UO_129 (O_129,N_7759,N_8564);
nor UO_130 (O_130,N_9057,N_9695);
nor UO_131 (O_131,N_8385,N_8982);
or UO_132 (O_132,N_7537,N_8232);
or UO_133 (O_133,N_7867,N_7809);
and UO_134 (O_134,N_9403,N_8852);
nor UO_135 (O_135,N_8000,N_9399);
nor UO_136 (O_136,N_7947,N_7690);
nand UO_137 (O_137,N_9507,N_7781);
and UO_138 (O_138,N_9338,N_9398);
or UO_139 (O_139,N_7882,N_7536);
xnor UO_140 (O_140,N_7607,N_8713);
nand UO_141 (O_141,N_8231,N_9438);
xnor UO_142 (O_142,N_9630,N_9424);
nor UO_143 (O_143,N_9466,N_8316);
and UO_144 (O_144,N_9448,N_8869);
and UO_145 (O_145,N_8465,N_9726);
xor UO_146 (O_146,N_8345,N_7652);
nand UO_147 (O_147,N_9943,N_8975);
nand UO_148 (O_148,N_9442,N_7608);
nor UO_149 (O_149,N_8436,N_8166);
nand UO_150 (O_150,N_9952,N_9099);
nand UO_151 (O_151,N_8793,N_9840);
and UO_152 (O_152,N_9051,N_9939);
or UO_153 (O_153,N_7569,N_8885);
and UO_154 (O_154,N_8011,N_7779);
nor UO_155 (O_155,N_8373,N_7564);
nand UO_156 (O_156,N_9446,N_8212);
nand UO_157 (O_157,N_8399,N_7622);
and UO_158 (O_158,N_7868,N_9259);
or UO_159 (O_159,N_9593,N_9833);
and UO_160 (O_160,N_8660,N_8730);
nor UO_161 (O_161,N_7533,N_9683);
xor UO_162 (O_162,N_8922,N_8559);
nand UO_163 (O_163,N_8475,N_7636);
nor UO_164 (O_164,N_7518,N_9200);
nand UO_165 (O_165,N_8514,N_7820);
or UO_166 (O_166,N_8071,N_7812);
nand UO_167 (O_167,N_8871,N_9265);
and UO_168 (O_168,N_9887,N_8887);
nor UO_169 (O_169,N_8939,N_9916);
and UO_170 (O_170,N_9736,N_7705);
and UO_171 (O_171,N_8435,N_7673);
nor UO_172 (O_172,N_9881,N_7513);
or UO_173 (O_173,N_9836,N_9533);
nor UO_174 (O_174,N_9787,N_9489);
nand UO_175 (O_175,N_9349,N_8500);
xnor UO_176 (O_176,N_7688,N_8928);
or UO_177 (O_177,N_8523,N_7967);
or UO_178 (O_178,N_9957,N_9511);
or UO_179 (O_179,N_9856,N_8739);
xnor UO_180 (O_180,N_9575,N_9482);
or UO_181 (O_181,N_9954,N_7773);
nand UO_182 (O_182,N_8707,N_7698);
nand UO_183 (O_183,N_8586,N_9129);
nor UO_184 (O_184,N_8993,N_7554);
or UO_185 (O_185,N_9047,N_9871);
nand UO_186 (O_186,N_9144,N_8985);
xnor UO_187 (O_187,N_7544,N_8905);
nor UO_188 (O_188,N_9618,N_7565);
nand UO_189 (O_189,N_8158,N_9623);
and UO_190 (O_190,N_9495,N_9437);
nand UO_191 (O_191,N_8673,N_7877);
or UO_192 (O_192,N_8152,N_7583);
nand UO_193 (O_193,N_8692,N_9897);
nand UO_194 (O_194,N_8249,N_8031);
and UO_195 (O_195,N_7926,N_9505);
and UO_196 (O_196,N_7646,N_9019);
nor UO_197 (O_197,N_7801,N_9264);
xnor UO_198 (O_198,N_8725,N_9690);
or UO_199 (O_199,N_8620,N_9909);
and UO_200 (O_200,N_8530,N_8937);
nand UO_201 (O_201,N_9104,N_8863);
xor UO_202 (O_202,N_8129,N_8491);
and UO_203 (O_203,N_8818,N_9364);
and UO_204 (O_204,N_8233,N_9760);
or UO_205 (O_205,N_9267,N_9498);
nand UO_206 (O_206,N_9503,N_9691);
nor UO_207 (O_207,N_9052,N_8999);
nand UO_208 (O_208,N_8518,N_8276);
nor UO_209 (O_209,N_9948,N_9134);
nor UO_210 (O_210,N_9212,N_9033);
nor UO_211 (O_211,N_9170,N_8102);
nor UO_212 (O_212,N_7966,N_7859);
nand UO_213 (O_213,N_9592,N_8452);
nand UO_214 (O_214,N_8420,N_9239);
nor UO_215 (O_215,N_8624,N_8526);
nor UO_216 (O_216,N_7542,N_9257);
or UO_217 (O_217,N_9647,N_7802);
nand UO_218 (O_218,N_9602,N_9061);
nand UO_219 (O_219,N_8432,N_9054);
nor UO_220 (O_220,N_8338,N_8370);
nor UO_221 (O_221,N_9412,N_8990);
or UO_222 (O_222,N_9843,N_8778);
nand UO_223 (O_223,N_8560,N_8219);
nor UO_224 (O_224,N_7946,N_8744);
or UO_225 (O_225,N_8310,N_9217);
nor UO_226 (O_226,N_8391,N_8075);
or UO_227 (O_227,N_7810,N_9044);
or UO_228 (O_228,N_8520,N_8717);
xnor UO_229 (O_229,N_9947,N_9816);
nor UO_230 (O_230,N_7803,N_9761);
nor UO_231 (O_231,N_9876,N_9679);
and UO_232 (O_232,N_9607,N_8270);
nand UO_233 (O_233,N_8771,N_9735);
and UO_234 (O_234,N_8140,N_9802);
and UO_235 (O_235,N_8145,N_7922);
or UO_236 (O_236,N_8234,N_9540);
or UO_237 (O_237,N_8823,N_7540);
or UO_238 (O_238,N_7730,N_8841);
and UO_239 (O_239,N_9243,N_8073);
nand UO_240 (O_240,N_8260,N_9005);
or UO_241 (O_241,N_8845,N_9889);
or UO_242 (O_242,N_9284,N_8710);
nor UO_243 (O_243,N_9024,N_8142);
nand UO_244 (O_244,N_8349,N_8574);
and UO_245 (O_245,N_7697,N_7696);
xnor UO_246 (O_246,N_9994,N_9776);
xnor UO_247 (O_247,N_8164,N_7672);
or UO_248 (O_248,N_7610,N_9907);
nor UO_249 (O_249,N_9413,N_8122);
nor UO_250 (O_250,N_7982,N_9222);
and UO_251 (O_251,N_8098,N_8960);
or UO_252 (O_252,N_9846,N_8727);
nor UO_253 (O_253,N_7798,N_8236);
or UO_254 (O_254,N_8155,N_9671);
or UO_255 (O_255,N_7756,N_9408);
and UO_256 (O_256,N_8362,N_8271);
nand UO_257 (O_257,N_9484,N_9975);
or UO_258 (O_258,N_9908,N_8502);
and UO_259 (O_259,N_8651,N_8795);
nor UO_260 (O_260,N_8146,N_9705);
or UO_261 (O_261,N_9785,N_7772);
or UO_262 (O_262,N_8409,N_8854);
nor UO_263 (O_263,N_9298,N_7925);
nor UO_264 (O_264,N_7890,N_8915);
nor UO_265 (O_265,N_7737,N_8801);
or UO_266 (O_266,N_9449,N_9737);
nor UO_267 (O_267,N_8842,N_9917);
and UO_268 (O_268,N_8699,N_8309);
nor UO_269 (O_269,N_9258,N_8451);
nand UO_270 (O_270,N_9328,N_8055);
and UO_271 (O_271,N_9981,N_9132);
or UO_272 (O_272,N_8199,N_9612);
or UO_273 (O_273,N_8987,N_8573);
and UO_274 (O_274,N_9719,N_8114);
nand UO_275 (O_275,N_8312,N_8712);
and UO_276 (O_276,N_8578,N_8629);
nor UO_277 (O_277,N_8898,N_9886);
xnor UO_278 (O_278,N_9319,N_9101);
xor UO_279 (O_279,N_9806,N_7691);
nor UO_280 (O_280,N_9470,N_8320);
and UO_281 (O_281,N_9037,N_9670);
nor UO_282 (O_282,N_8902,N_8570);
or UO_283 (O_283,N_8296,N_8360);
nand UO_284 (O_284,N_9515,N_8216);
nand UO_285 (O_285,N_9542,N_8223);
nor UO_286 (O_286,N_9003,N_7965);
nand UO_287 (O_287,N_8708,N_9158);
nor UO_288 (O_288,N_7599,N_9450);
and UO_289 (O_289,N_8376,N_9039);
nor UO_290 (O_290,N_9491,N_9919);
xnor UO_291 (O_291,N_9867,N_8742);
or UO_292 (O_292,N_8767,N_9007);
or UO_293 (O_293,N_7930,N_7948);
and UO_294 (O_294,N_9891,N_7832);
nand UO_295 (O_295,N_8731,N_8804);
or UO_296 (O_296,N_9065,N_9182);
nor UO_297 (O_297,N_7917,N_8529);
nand UO_298 (O_298,N_7857,N_8449);
and UO_299 (O_299,N_9422,N_8471);
nor UO_300 (O_300,N_8899,N_9327);
nand UO_301 (O_301,N_7606,N_7864);
or UO_302 (O_302,N_9539,N_9832);
or UO_303 (O_303,N_8032,N_9241);
nor UO_304 (O_304,N_8253,N_8864);
nand UO_305 (O_305,N_8511,N_8839);
and UO_306 (O_306,N_8367,N_9064);
nor UO_307 (O_307,N_7870,N_9389);
or UO_308 (O_308,N_9763,N_9676);
or UO_309 (O_309,N_9220,N_9932);
or UO_310 (O_310,N_9494,N_8162);
or UO_311 (O_311,N_8949,N_9153);
nor UO_312 (O_312,N_8027,N_7625);
and UO_313 (O_313,N_8268,N_7761);
and UO_314 (O_314,N_9532,N_8897);
nor UO_315 (O_315,N_9615,N_8424);
nand UO_316 (O_316,N_7776,N_9194);
nand UO_317 (O_317,N_8548,N_9497);
and UO_318 (O_318,N_9873,N_7797);
and UO_319 (O_319,N_8621,N_9729);
xnor UO_320 (O_320,N_8867,N_8953);
and UO_321 (O_321,N_8263,N_7879);
nand UO_322 (O_322,N_8159,N_9121);
nor UO_323 (O_323,N_8390,N_9083);
nor UO_324 (O_324,N_9959,N_9847);
nor UO_325 (O_325,N_9724,N_8352);
nor UO_326 (O_326,N_8824,N_9381);
nand UO_327 (O_327,N_9530,N_7968);
nor UO_328 (O_328,N_9049,N_7510);
or UO_329 (O_329,N_9604,N_7630);
and UO_330 (O_330,N_9197,N_8141);
nand UO_331 (O_331,N_7817,N_7860);
nand UO_332 (O_332,N_8359,N_9864);
and UO_333 (O_333,N_9603,N_9606);
and UO_334 (O_334,N_8192,N_9700);
and UO_335 (O_335,N_8498,N_8242);
nand UO_336 (O_336,N_8917,N_8119);
nor UO_337 (O_337,N_7522,N_9199);
and UO_338 (O_338,N_8464,N_8259);
xor UO_339 (O_339,N_9697,N_8091);
or UO_340 (O_340,N_7814,N_9043);
nand UO_341 (O_341,N_8984,N_7714);
xor UO_342 (O_342,N_8616,N_9797);
xor UO_343 (O_343,N_7623,N_7530);
or UO_344 (O_344,N_8703,N_8239);
and UO_345 (O_345,N_8176,N_8229);
nand UO_346 (O_346,N_9654,N_8808);
or UO_347 (O_347,N_8977,N_8487);
nor UO_348 (O_348,N_8865,N_7738);
or UO_349 (O_349,N_8116,N_9143);
and UO_350 (O_350,N_9286,N_7643);
nand UO_351 (O_351,N_9693,N_7632);
nand UO_352 (O_352,N_7865,N_9928);
and UO_353 (O_353,N_8365,N_8324);
or UO_354 (O_354,N_7619,N_9046);
nand UO_355 (O_355,N_8054,N_9783);
and UO_356 (O_356,N_8992,N_7570);
xnor UO_357 (O_357,N_9557,N_8588);
and UO_358 (O_358,N_8455,N_9260);
and UO_359 (O_359,N_8001,N_8969);
nand UO_360 (O_360,N_9436,N_7900);
or UO_361 (O_361,N_9017,N_8535);
nand UO_362 (O_362,N_9390,N_9306);
xnor UO_363 (O_363,N_7951,N_9502);
and UO_364 (O_364,N_8097,N_7849);
xor UO_365 (O_365,N_9421,N_8579);
nor UO_366 (O_366,N_8545,N_9240);
nand UO_367 (O_367,N_8690,N_8374);
or UO_368 (O_368,N_8472,N_7524);
nand UO_369 (O_369,N_9588,N_9906);
or UO_370 (O_370,N_8843,N_8012);
nor UO_371 (O_371,N_8020,N_7594);
xor UO_372 (O_372,N_7969,N_9116);
nor UO_373 (O_373,N_8662,N_9513);
xor UO_374 (O_374,N_8278,N_7543);
nor UO_375 (O_375,N_9167,N_7984);
and UO_376 (O_376,N_8017,N_9685);
or UO_377 (O_377,N_8100,N_9565);
and UO_378 (O_378,N_8330,N_9192);
and UO_379 (O_379,N_8705,N_9556);
and UO_380 (O_380,N_9875,N_9696);
xnor UO_381 (O_381,N_8107,N_7878);
and UO_382 (O_382,N_8508,N_8674);
nor UO_383 (O_383,N_8938,N_7763);
nand UO_384 (O_384,N_9059,N_8026);
or UO_385 (O_385,N_7938,N_9834);
and UO_386 (O_386,N_8648,N_9581);
and UO_387 (O_387,N_9583,N_9577);
nand UO_388 (O_388,N_8138,N_8224);
or UO_389 (O_389,N_8504,N_9376);
or UO_390 (O_390,N_9316,N_9874);
or UO_391 (O_391,N_9367,N_9120);
or UO_392 (O_392,N_9855,N_8457);
nor UO_393 (O_393,N_9668,N_7683);
nor UO_394 (O_394,N_8218,N_8613);
and UO_395 (O_395,N_8762,N_7853);
or UO_396 (O_396,N_8716,N_7745);
or UO_397 (O_397,N_9340,N_8682);
and UO_398 (O_398,N_9665,N_7749);
nor UO_399 (O_399,N_8786,N_9660);
or UO_400 (O_400,N_9341,N_9266);
or UO_401 (O_401,N_9373,N_8968);
xor UO_402 (O_402,N_8790,N_8111);
nand UO_403 (O_403,N_8668,N_8049);
nor UO_404 (O_404,N_8623,N_9304);
nand UO_405 (O_405,N_9564,N_9000);
nor UO_406 (O_406,N_8758,N_8733);
and UO_407 (O_407,N_8404,N_9287);
or UO_408 (O_408,N_8115,N_7962);
xor UO_409 (O_409,N_8914,N_8770);
and UO_410 (O_410,N_7604,N_7588);
and UO_411 (O_411,N_8667,N_8774);
and UO_412 (O_412,N_9314,N_8524);
nand UO_413 (O_413,N_7873,N_9021);
or UO_414 (O_414,N_8794,N_9499);
or UO_415 (O_415,N_8294,N_8709);
or UO_416 (O_416,N_7992,N_9809);
nor UO_417 (O_417,N_8920,N_8440);
or UO_418 (O_418,N_7985,N_8205);
nor UO_419 (O_419,N_8109,N_8248);
nor UO_420 (O_420,N_9940,N_8406);
and UO_421 (O_421,N_9152,N_9998);
xnor UO_422 (O_422,N_8551,N_7548);
xor UO_423 (O_423,N_8833,N_9643);
or UO_424 (O_424,N_8095,N_8600);
nand UO_425 (O_425,N_9718,N_7631);
nand UO_426 (O_426,N_8635,N_9014);
nor UO_427 (O_427,N_8368,N_8198);
nand UO_428 (O_428,N_8041,N_9069);
nor UO_429 (O_429,N_8598,N_9018);
nor UO_430 (O_430,N_8182,N_7515);
or UO_431 (O_431,N_7710,N_9764);
and UO_432 (O_432,N_8168,N_8715);
and UO_433 (O_433,N_9544,N_8351);
or UO_434 (O_434,N_8505,N_8860);
or UO_435 (O_435,N_8936,N_8395);
and UO_436 (O_436,N_8008,N_9009);
nand UO_437 (O_437,N_7786,N_7828);
and UO_438 (O_438,N_9741,N_7923);
nand UO_439 (O_439,N_9425,N_8633);
nand UO_440 (O_440,N_7780,N_8596);
and UO_441 (O_441,N_8209,N_9958);
and UO_442 (O_442,N_8279,N_9510);
and UO_443 (O_443,N_9571,N_9475);
or UO_444 (O_444,N_7602,N_8482);
and UO_445 (O_445,N_8654,N_7808);
xor UO_446 (O_446,N_7914,N_8501);
or UO_447 (O_447,N_9087,N_9339);
or UO_448 (O_448,N_9815,N_9126);
nand UO_449 (O_449,N_9765,N_7675);
nor UO_450 (O_450,N_8488,N_9370);
nand UO_451 (O_451,N_7834,N_8246);
and UO_452 (O_452,N_9420,N_8206);
nand UO_453 (O_453,N_7609,N_8828);
and UO_454 (O_454,N_8909,N_8333);
nand UO_455 (O_455,N_9045,N_9325);
xor UO_456 (O_456,N_9342,N_8779);
nand UO_457 (O_457,N_8025,N_9702);
xor UO_458 (O_458,N_8561,N_8632);
and UO_459 (O_459,N_8187,N_7959);
and UO_460 (O_460,N_9397,N_9270);
nand UO_461 (O_461,N_8038,N_8861);
nand UO_462 (O_462,N_8812,N_9219);
nor UO_463 (O_463,N_9308,N_8124);
nand UO_464 (O_464,N_9927,N_8565);
nor UO_465 (O_465,N_9118,N_8003);
xor UO_466 (O_466,N_8235,N_8128);
xor UO_467 (O_467,N_9109,N_8967);
or UO_468 (O_468,N_8418,N_9172);
nor UO_469 (O_469,N_9020,N_8587);
and UO_470 (O_470,N_9960,N_8815);
nor UO_471 (O_471,N_9600,N_8096);
nand UO_472 (O_472,N_8477,N_9404);
nor UO_473 (O_473,N_7595,N_7918);
and UO_474 (O_474,N_8552,N_9225);
nand UO_475 (O_475,N_9487,N_9008);
and UO_476 (O_476,N_9811,N_8378);
and UO_477 (O_477,N_8533,N_9189);
nor UO_478 (O_478,N_8480,N_8611);
nand UO_479 (O_479,N_7503,N_8408);
or UO_480 (O_480,N_8509,N_8653);
nand UO_481 (O_481,N_8103,N_8569);
and UO_482 (O_482,N_8052,N_9249);
or UO_483 (O_483,N_9687,N_7804);
and UO_484 (O_484,N_8783,N_8628);
nor UO_485 (O_485,N_8799,N_9457);
and UO_486 (O_486,N_8009,N_9216);
and UO_487 (O_487,N_8004,N_9779);
nand UO_488 (O_488,N_8018,N_7852);
or UO_489 (O_489,N_9221,N_7898);
nor UO_490 (O_490,N_8076,N_7933);
and UO_491 (O_491,N_8834,N_9299);
or UO_492 (O_492,N_9464,N_8266);
and UO_493 (O_493,N_8846,N_8615);
and UO_494 (O_494,N_8781,N_8190);
nor UO_495 (O_495,N_9070,N_9486);
nand UO_496 (O_496,N_7963,N_8776);
nor UO_497 (O_497,N_8356,N_8603);
nor UO_498 (O_498,N_9075,N_8019);
and UO_499 (O_499,N_8257,N_8507);
or UO_500 (O_500,N_9031,N_8326);
or UO_501 (O_501,N_8859,N_9712);
and UO_502 (O_502,N_9882,N_9757);
nand UO_503 (O_503,N_8057,N_7556);
or UO_504 (O_504,N_9851,N_9157);
xor UO_505 (O_505,N_7792,N_7579);
and UO_506 (O_506,N_8445,N_8369);
nand UO_507 (O_507,N_9400,N_9276);
or UO_508 (O_508,N_9410,N_8156);
or UO_509 (O_509,N_7514,N_8550);
nand UO_510 (O_510,N_9206,N_7674);
and UO_511 (O_511,N_7818,N_9863);
or UO_512 (O_512,N_7915,N_9732);
nand UO_513 (O_513,N_7719,N_7717);
xnor UO_514 (O_514,N_8081,N_9963);
or UO_515 (O_515,N_7767,N_9485);
xor UO_516 (O_516,N_8607,N_7735);
nor UO_517 (O_517,N_9113,N_8930);
and UO_518 (O_518,N_9456,N_9110);
nor UO_519 (O_519,N_9933,N_9673);
and UO_520 (O_520,N_8908,N_9805);
xor UO_521 (O_521,N_8172,N_8419);
or UO_522 (O_522,N_9245,N_9411);
nand UO_523 (O_523,N_7593,N_8195);
nor UO_524 (O_524,N_9821,N_9973);
nand UO_525 (O_525,N_8996,N_9742);
or UO_526 (O_526,N_8609,N_9596);
and UO_527 (O_527,N_8132,N_9801);
or UO_528 (O_528,N_9078,N_9137);
or UO_529 (O_529,N_9996,N_8844);
or UO_530 (O_530,N_8531,N_8293);
and UO_531 (O_531,N_9755,N_7783);
nand UO_532 (O_532,N_7990,N_8220);
and UO_533 (O_533,N_9115,N_9822);
nor UO_534 (O_534,N_9242,N_9330);
nor UO_535 (O_535,N_8694,N_9006);
and UO_536 (O_536,N_8186,N_7896);
nor UO_537 (O_537,N_8946,N_7733);
or UO_538 (O_538,N_9619,N_9238);
or UO_539 (O_539,N_8558,N_8584);
and UO_540 (O_540,N_8971,N_8265);
xor UO_541 (O_541,N_9125,N_9201);
nand UO_542 (O_542,N_8387,N_9139);
nand UO_543 (O_543,N_7723,N_7641);
nand UO_544 (O_544,N_9296,N_7897);
nand UO_545 (O_545,N_8078,N_9290);
and UO_546 (O_546,N_9369,N_7885);
nor UO_547 (O_547,N_9004,N_9401);
nand UO_548 (O_548,N_7670,N_9394);
or UO_549 (O_549,N_7701,N_7535);
and UO_550 (O_550,N_9899,N_9053);
and UO_551 (O_551,N_9506,N_7949);
and UO_552 (O_552,N_7731,N_9156);
nor UO_553 (O_553,N_9995,N_9849);
nand UO_554 (O_554,N_7906,N_8252);
and UO_555 (O_555,N_9022,N_9013);
nor UO_556 (O_556,N_9148,N_9150);
xnor UO_557 (O_557,N_8101,N_7986);
and UO_558 (O_558,N_8230,N_8167);
nor UO_559 (O_559,N_9262,N_7999);
or UO_560 (O_560,N_9088,N_7547);
or UO_561 (O_561,N_8677,N_7987);
nand UO_562 (O_562,N_8288,N_8468);
or UO_563 (O_563,N_7601,N_7856);
nand UO_564 (O_564,N_9582,N_9181);
or UO_565 (O_565,N_8179,N_8113);
nand UO_566 (O_566,N_9291,N_9566);
and UO_567 (O_567,N_8393,N_7844);
and UO_568 (O_568,N_8446,N_9970);
and UO_569 (O_569,N_8450,N_8226);
or UO_570 (O_570,N_8582,N_7895);
and UO_571 (O_571,N_8723,N_9738);
or UO_572 (O_572,N_8672,N_9352);
or UO_573 (O_573,N_9858,N_9925);
nand UO_574 (O_574,N_9015,N_8127);
or UO_575 (O_575,N_9307,N_9336);
nand UO_576 (O_576,N_8254,N_9377);
or UO_577 (O_577,N_8966,N_9175);
or UO_578 (O_578,N_9534,N_8379);
nand UO_579 (O_579,N_9223,N_7708);
and UO_580 (O_580,N_9140,N_7978);
nand UO_581 (O_581,N_9638,N_9524);
nor UO_582 (O_582,N_8979,N_8765);
and UO_583 (O_583,N_8188,N_9098);
xor UO_584 (O_584,N_7728,N_9709);
and UO_585 (O_585,N_9525,N_7903);
and UO_586 (O_586,N_7980,N_8251);
nand UO_587 (O_587,N_9202,N_9281);
nor UO_588 (O_588,N_8912,N_9938);
xnor UO_589 (O_589,N_8597,N_8892);
and UO_590 (O_590,N_8649,N_9644);
or UO_591 (O_591,N_7720,N_8800);
and UO_592 (O_592,N_7657,N_9771);
nor UO_593 (O_593,N_8125,N_9812);
nor UO_594 (O_594,N_8347,N_9639);
nor UO_595 (O_595,N_9953,N_9850);
nand UO_596 (O_596,N_8143,N_7858);
nor UO_597 (O_597,N_7576,N_8606);
nand UO_598 (O_598,N_9165,N_7693);
and UO_599 (O_599,N_9976,N_9251);
nor UO_600 (O_600,N_8015,N_8458);
and UO_601 (O_601,N_8918,N_7861);
or UO_602 (O_602,N_8602,N_7709);
nor UO_603 (O_603,N_9230,N_9625);
nand UO_604 (O_604,N_9701,N_9042);
and UO_605 (O_605,N_8323,N_7627);
xor UO_606 (O_606,N_9885,N_9164);
or UO_607 (O_607,N_8386,N_7871);
nor UO_608 (O_608,N_9869,N_7611);
or UO_609 (O_609,N_8039,N_7680);
or UO_610 (O_610,N_9273,N_8297);
nand UO_611 (O_611,N_8959,N_7752);
and UO_612 (O_612,N_8469,N_9978);
and UO_613 (O_613,N_8644,N_9956);
nor UO_614 (O_614,N_8626,N_7685);
nand UO_615 (O_615,N_9559,N_7975);
or UO_616 (O_616,N_7919,N_9452);
xor UO_617 (O_617,N_8549,N_9750);
xor UO_618 (O_618,N_7613,N_8160);
nand UO_619 (O_619,N_7704,N_8983);
or UO_620 (O_620,N_9921,N_9393);
or UO_621 (O_621,N_8666,N_9097);
nor UO_622 (O_622,N_9368,N_8882);
nand UO_623 (O_623,N_8194,N_8747);
or UO_624 (O_624,N_9271,N_8277);
nor UO_625 (O_625,N_9149,N_9594);
xor UO_626 (O_626,N_8467,N_9434);
nor UO_627 (O_627,N_7559,N_7684);
nand UO_628 (O_628,N_8085,N_9161);
nand UO_629 (O_629,N_9163,N_8336);
or UO_630 (O_630,N_9541,N_9504);
nor UO_631 (O_631,N_8200,N_9294);
nand UO_632 (O_632,N_8154,N_9178);
nand UO_633 (O_633,N_9734,N_7807);
and UO_634 (O_634,N_9573,N_7800);
or UO_635 (O_635,N_9282,N_7911);
or UO_636 (O_636,N_9551,N_9723);
or UO_637 (O_637,N_8053,N_8701);
and UO_638 (O_638,N_7640,N_8082);
nand UO_639 (O_639,N_9092,N_9848);
or UO_640 (O_640,N_7574,N_9073);
nand UO_641 (O_641,N_9058,N_9715);
or UO_642 (O_642,N_9191,N_9678);
or UO_643 (O_643,N_9980,N_7634);
xor UO_644 (O_644,N_9708,N_7974);
and UO_645 (O_645,N_8063,N_8203);
or UO_646 (O_646,N_9155,N_9112);
or UO_647 (O_647,N_9318,N_8240);
xnor UO_648 (O_648,N_7835,N_9662);
nand UO_649 (O_649,N_9107,N_7770);
nand UO_650 (O_650,N_7572,N_8884);
or UO_651 (O_651,N_8104,N_8306);
and UO_652 (O_652,N_8042,N_7534);
and UO_653 (O_653,N_8046,N_8641);
or UO_654 (O_654,N_8978,N_9914);
xnor UO_655 (O_655,N_9554,N_8394);
xnor UO_656 (O_656,N_7687,N_8444);
nand UO_657 (O_657,N_8402,N_8601);
nor UO_658 (O_658,N_7566,N_9016);
and UO_659 (O_659,N_7713,N_9133);
nand UO_660 (O_660,N_7826,N_8604);
and UO_661 (O_661,N_9642,N_8007);
xor UO_662 (O_662,N_9704,N_8958);
nor UO_663 (O_663,N_9628,N_9831);
nor UO_664 (O_664,N_9877,N_9025);
xnor UO_665 (O_665,N_8303,N_9232);
or UO_666 (O_666,N_8428,N_9721);
or UO_667 (O_667,N_9633,N_9841);
nor UO_668 (O_668,N_7825,N_9431);
xor UO_669 (O_669,N_9538,N_8305);
xnor UO_670 (O_670,N_8658,N_7886);
xor UO_671 (O_671,N_8327,N_9951);
or UO_672 (O_672,N_9710,N_7508);
and UO_673 (O_673,N_8926,N_8483);
nand UO_674 (O_674,N_9142,N_8461);
xor UO_675 (O_675,N_9435,N_8752);
and UO_676 (O_676,N_9492,N_9124);
nand UO_677 (O_677,N_8817,N_8412);
nand UO_678 (O_678,N_9669,N_9605);
and UO_679 (O_679,N_7821,N_8734);
nor UO_680 (O_680,N_9430,N_7764);
or UO_681 (O_681,N_8608,N_7931);
nor UO_682 (O_682,N_9931,N_8663);
nand UO_683 (O_683,N_8728,N_8577);
nand UO_684 (O_684,N_8675,N_8047);
and UO_685 (O_685,N_9322,N_7977);
nor UO_686 (O_686,N_8227,N_7665);
or UO_687 (O_687,N_9166,N_9655);
or UO_688 (O_688,N_8910,N_9418);
or UO_689 (O_689,N_9406,N_8460);
nor UO_690 (O_690,N_8989,N_9253);
and UO_691 (O_691,N_8772,N_8077);
and UO_692 (O_692,N_7880,N_9321);
nor UO_693 (O_693,N_7663,N_9717);
nor UO_694 (O_694,N_8388,N_7943);
and UO_695 (O_695,N_9950,N_9520);
or UO_696 (O_696,N_9842,N_8281);
nor UO_697 (O_697,N_8554,N_8361);
and UO_698 (O_698,N_9674,N_9261);
or UO_699 (O_699,N_8400,N_8656);
nor UO_700 (O_700,N_7516,N_8718);
or UO_701 (O_701,N_8519,N_7970);
and UO_702 (O_702,N_8876,N_8965);
nor UO_703 (O_703,N_9990,N_8439);
or UO_704 (O_704,N_8006,N_9077);
or UO_705 (O_705,N_9190,N_7899);
nor UO_706 (O_706,N_8973,N_9146);
xor UO_707 (O_707,N_7811,N_9969);
nand UO_708 (O_708,N_7686,N_8056);
nand UO_709 (O_709,N_8997,N_8384);
nand UO_710 (O_710,N_9997,N_9941);
nor UO_711 (O_711,N_9942,N_9477);
or UO_712 (O_712,N_7635,N_8963);
nor UO_713 (O_713,N_8340,N_9985);
nor UO_714 (O_714,N_8721,N_9547);
and UO_715 (O_715,N_9694,N_8355);
xnor UO_716 (O_716,N_8766,N_8207);
and UO_717 (O_717,N_9102,N_9067);
and UO_718 (O_718,N_9196,N_8642);
nand UO_719 (O_719,N_9751,N_7833);
or UO_720 (O_720,N_7957,N_8272);
and UO_721 (O_721,N_8874,N_7778);
nand UO_722 (O_722,N_7907,N_7789);
nor UO_723 (O_723,N_8961,N_9415);
nand UO_724 (O_724,N_8433,N_8225);
and UO_725 (O_725,N_8274,N_7666);
nand UO_726 (O_726,N_7531,N_9423);
and UO_727 (O_727,N_8546,N_8147);
xnor UO_728 (O_728,N_9923,N_8957);
and UO_729 (O_729,N_8021,N_7921);
nor UO_730 (O_730,N_8048,N_7845);
or UO_731 (O_731,N_7934,N_9609);
and UO_732 (O_732,N_8447,N_8696);
and UO_733 (O_733,N_9279,N_9961);
nand UO_734 (O_734,N_7958,N_7902);
nor UO_735 (O_735,N_9179,N_8691);
xor UO_736 (O_736,N_8664,N_8120);
or UO_737 (O_737,N_8068,N_8506);
nand UO_738 (O_738,N_8149,N_8751);
or UO_739 (O_739,N_8175,N_8893);
and UO_740 (O_740,N_8261,N_8094);
nand UO_741 (O_741,N_9585,N_9766);
nor UO_742 (O_742,N_9233,N_9979);
or UO_743 (O_743,N_9062,N_7715);
nor UO_744 (O_744,N_9986,N_7796);
nor UO_745 (O_745,N_8924,N_9441);
nand UO_746 (O_746,N_9226,N_7961);
and UO_747 (O_747,N_8174,N_8919);
nor UO_748 (O_748,N_8431,N_7837);
and UO_749 (O_749,N_9365,N_9063);
nor UO_750 (O_750,N_7648,N_7863);
nor UO_751 (O_751,N_7561,N_8204);
xnor UO_752 (O_752,N_9516,N_9622);
nand UO_753 (O_753,N_7729,N_7769);
nor UO_754 (O_754,N_9359,N_7993);
or UO_755 (O_755,N_9992,N_8935);
nand UO_756 (O_756,N_8454,N_8334);
nor UO_757 (O_757,N_8322,N_9483);
and UO_758 (O_758,N_8029,N_7591);
and UO_759 (O_759,N_9545,N_7960);
or UO_760 (O_760,N_7651,N_7971);
nor UO_761 (O_761,N_9967,N_8749);
nand UO_762 (O_762,N_9068,N_8317);
nor UO_763 (O_763,N_8831,N_8891);
nor UO_764 (O_764,N_9447,N_9160);
and UO_765 (O_765,N_8614,N_9439);
nor UO_766 (O_766,N_8040,N_9827);
and UO_767 (O_767,N_8780,N_9168);
xor UO_768 (O_768,N_9740,N_9558);
and UO_769 (O_769,N_7936,N_9637);
and UO_770 (O_770,N_8286,N_8070);
or UO_771 (O_771,N_9012,N_9905);
nand UO_772 (O_772,N_8256,N_9752);
nand UO_773 (O_773,N_9500,N_9028);
nor UO_774 (O_774,N_7940,N_7913);
or UO_775 (O_775,N_9550,N_9854);
or UO_776 (O_776,N_9893,N_7702);
or UO_777 (O_777,N_7777,N_8022);
nand UO_778 (O_778,N_9023,N_8434);
nor UO_779 (O_779,N_8459,N_8411);
or UO_780 (O_780,N_9707,N_9136);
nand UO_781 (O_781,N_7577,N_7799);
or UO_782 (O_782,N_9912,N_9769);
nor UO_783 (O_783,N_9204,N_8738);
nand UO_784 (O_784,N_9354,N_9720);
or UO_785 (O_785,N_8931,N_8681);
nand UO_786 (O_786,N_9231,N_9730);
xor UO_787 (O_787,N_7739,N_8991);
nor UO_788 (O_788,N_9193,N_9055);
or UO_789 (O_789,N_9297,N_7681);
xnor UO_790 (O_790,N_9684,N_8746);
nand UO_791 (O_791,N_8153,N_8683);
nor UO_792 (O_792,N_7500,N_7529);
nor UO_793 (O_793,N_7843,N_9414);
nor UO_794 (O_794,N_9580,N_9127);
nor UO_795 (O_795,N_8250,N_8169);
nand UO_796 (O_796,N_9184,N_9493);
and UO_797 (O_797,N_8313,N_8689);
or UO_798 (O_798,N_9686,N_9681);
nor UO_799 (O_799,N_8425,N_9884);
nor UO_800 (O_800,N_8782,N_9176);
nor UO_801 (O_801,N_8069,N_7692);
xor UO_802 (O_802,N_7502,N_9860);
and UO_803 (O_803,N_8873,N_9835);
nand UO_804 (O_804,N_9272,N_8575);
nand UO_805 (O_805,N_8184,N_7953);
nand UO_806 (O_806,N_8543,N_9910);
nand UO_807 (O_807,N_8821,N_9640);
nor UO_808 (O_808,N_8238,N_8951);
nand UO_809 (O_809,N_9746,N_7869);
nor UO_810 (O_810,N_9048,N_9351);
nand UO_811 (O_811,N_8945,N_9548);
nand UO_812 (O_812,N_8567,N_8121);
nand UO_813 (O_813,N_8364,N_7546);
nor UO_814 (O_814,N_8426,N_7707);
nand UO_815 (O_815,N_9374,N_7874);
xnor UO_816 (O_816,N_8820,N_7795);
nor UO_817 (O_817,N_8222,N_7942);
nand UO_818 (O_818,N_8954,N_9034);
and UO_819 (O_819,N_8490,N_8366);
xor UO_820 (O_820,N_9205,N_7791);
and UO_821 (O_821,N_9937,N_9402);
xnor UO_822 (O_822,N_9578,N_8785);
nand UO_823 (O_823,N_9001,N_8088);
or UO_824 (O_824,N_7964,N_8350);
nand UO_825 (O_825,N_8745,N_8299);
xor UO_826 (O_826,N_9546,N_8637);
or UO_827 (O_827,N_7757,N_9090);
or UO_828 (O_828,N_9747,N_8646);
nand UO_829 (O_829,N_8851,N_9824);
xnor UO_830 (O_830,N_9094,N_9803);
and UO_831 (O_831,N_7620,N_9859);
or UO_832 (O_832,N_8423,N_9496);
and UO_833 (O_833,N_8150,N_7519);
and UO_834 (O_834,N_8377,N_9572);
or UO_835 (O_835,N_9455,N_8593);
nand UO_836 (O_836,N_7649,N_8619);
nor UO_837 (O_837,N_8580,N_9462);
and UO_838 (O_838,N_8816,N_9817);
xor UO_839 (O_839,N_9186,N_8976);
nor UO_840 (O_840,N_9474,N_9774);
xnor UO_841 (O_841,N_9269,N_9680);
nand UO_842 (O_842,N_8697,N_9419);
nor UO_843 (O_843,N_9714,N_8197);
or UO_844 (O_844,N_9333,N_9274);
nor UO_845 (O_845,N_9519,N_7578);
or UO_846 (O_846,N_8074,N_7580);
nand UO_847 (O_847,N_9460,N_9383);
nor UO_848 (O_848,N_8933,N_9521);
or UO_849 (O_849,N_8566,N_9355);
nand UO_850 (O_850,N_8084,N_9169);
or UO_851 (O_851,N_9195,N_7766);
nor UO_852 (O_852,N_8754,N_7892);
xnor UO_853 (O_853,N_8618,N_8840);
nand UO_854 (O_854,N_9828,N_7626);
and UO_855 (O_855,N_8679,N_9595);
and UO_856 (O_856,N_7727,N_7581);
xor UO_857 (O_857,N_9753,N_9813);
or UO_858 (O_858,N_9844,N_7590);
nor UO_859 (O_859,N_9661,N_9443);
nor UO_860 (O_860,N_9778,N_7782);
nand UO_861 (O_861,N_7771,N_8014);
nand UO_862 (O_862,N_8494,N_9632);
and UO_863 (O_863,N_8542,N_8879);
nand UO_864 (O_864,N_9334,N_9040);
and UO_865 (O_865,N_9862,N_7822);
nand UO_866 (O_866,N_8403,N_7629);
nor UO_867 (O_867,N_8290,N_9141);
nand UO_868 (O_868,N_8045,N_8665);
and UO_869 (O_869,N_7842,N_7910);
or UO_870 (O_870,N_9405,N_7894);
nor UO_871 (O_871,N_8210,N_9584);
nand UO_872 (O_872,N_7539,N_9210);
and UO_873 (O_873,N_8720,N_8339);
nor UO_874 (O_874,N_9072,N_7824);
and UO_875 (O_875,N_8262,N_9203);
nor UO_876 (O_876,N_9659,N_9293);
or UO_877 (O_877,N_8768,N_7550);
nor UO_878 (O_878,N_8726,N_9989);
nand UO_879 (O_879,N_7740,N_8437);
or UO_880 (O_880,N_8284,N_8788);
nand UO_881 (O_881,N_7846,N_9706);
nor UO_882 (O_882,N_7972,N_9145);
and UO_883 (O_883,N_8165,N_9479);
and UO_884 (O_884,N_8813,N_8855);
or UO_885 (O_885,N_8443,N_7793);
and UO_886 (O_886,N_9453,N_8466);
nor UO_887 (O_887,N_7836,N_7889);
nand UO_888 (O_888,N_8700,N_8878);
nor UO_889 (O_889,N_7664,N_8589);
or UO_890 (O_890,N_9598,N_9346);
or UO_891 (O_891,N_7644,N_8927);
nor UO_892 (O_892,N_7747,N_7654);
nand UO_893 (O_893,N_7525,N_9591);
xor UO_894 (O_894,N_9966,N_8066);
or UO_895 (O_895,N_8686,N_9076);
and UO_896 (O_896,N_8273,N_9417);
and UO_897 (O_897,N_8832,N_7955);
nor UO_898 (O_898,N_8023,N_9011);
nand UO_899 (O_899,N_8130,N_8307);
or UO_900 (O_900,N_8092,N_8630);
or UO_901 (O_901,N_9490,N_7743);
or UO_902 (O_902,N_8298,N_8470);
and UO_903 (O_903,N_8485,N_8201);
or UO_904 (O_904,N_9277,N_9645);
or UO_905 (O_905,N_7628,N_8736);
and UO_906 (O_906,N_9366,N_8650);
and UO_907 (O_907,N_7603,N_8590);
and UO_908 (O_908,N_7600,N_8131);
nand UO_909 (O_909,N_8757,N_8462);
and UO_910 (O_910,N_8836,N_9796);
nand UO_911 (O_911,N_8398,N_9010);
nor UO_912 (O_912,N_7711,N_7724);
nand UO_913 (O_913,N_9535,N_9562);
and UO_914 (O_914,N_7768,N_8148);
xor UO_915 (O_915,N_7532,N_7582);
nor UO_916 (O_916,N_8911,N_8534);
nor UO_917 (O_917,N_8777,N_9173);
or UO_918 (O_918,N_9292,N_9636);
or UO_919 (O_919,N_9866,N_7549);
nor UO_920 (O_920,N_9463,N_8974);
nand UO_921 (O_921,N_9807,N_7815);
nand UO_922 (O_922,N_7521,N_9892);
nor UO_923 (O_923,N_8981,N_8171);
nand UO_924 (O_924,N_8698,N_9512);
and UO_925 (O_925,N_7744,N_9444);
and UO_926 (O_926,N_9159,N_8329);
or UO_927 (O_927,N_8397,N_8422);
or UO_928 (O_928,N_9627,N_8735);
and UO_929 (O_929,N_8311,N_9629);
and UO_930 (O_930,N_9666,N_9608);
nor UO_931 (O_931,N_9865,N_8970);
xor UO_932 (O_932,N_9362,N_7571);
and UO_933 (O_933,N_7659,N_9692);
nand UO_934 (O_934,N_8478,N_8847);
nand UO_935 (O_935,N_9350,N_7785);
nand UO_936 (O_936,N_7831,N_9616);
nand UO_937 (O_937,N_9185,N_8105);
nand UO_938 (O_938,N_8243,N_9472);
xnor UO_939 (O_939,N_8346,N_9675);
or UO_940 (O_940,N_8211,N_8381);
and UO_941 (O_941,N_8517,N_8300);
or UO_942 (O_942,N_8557,N_8202);
or UO_943 (O_943,N_8463,N_8755);
xnor UO_944 (O_944,N_7703,N_8106);
nand UO_945 (O_945,N_8986,N_7650);
nand UO_946 (O_946,N_7653,N_9250);
nor UO_947 (O_947,N_8797,N_7658);
and UO_948 (O_948,N_8241,N_8264);
nor UO_949 (O_949,N_8807,N_7612);
xor UO_950 (O_950,N_8134,N_7551);
nand UO_951 (O_951,N_7573,N_9289);
or UO_952 (O_952,N_7614,N_7520);
xor UO_953 (O_953,N_8740,N_8016);
nand UO_954 (O_954,N_8877,N_9945);
nand UO_955 (O_955,N_8538,N_9386);
or UO_956 (O_956,N_9459,N_8072);
or UO_957 (O_957,N_7838,N_9537);
and UO_958 (O_958,N_9529,N_7850);
or UO_959 (O_959,N_9913,N_8117);
nand UO_960 (O_960,N_9656,N_8489);
nand UO_961 (O_961,N_9880,N_9614);
or UO_962 (O_962,N_9988,N_9522);
or UO_963 (O_963,N_9599,N_9553);
or UO_964 (O_964,N_8110,N_8438);
nand UO_965 (O_965,N_8940,N_9589);
nor UO_966 (O_966,N_7523,N_9093);
nor UO_967 (O_967,N_8090,N_8050);
and UO_968 (O_968,N_8058,N_9935);
or UO_969 (O_969,N_8215,N_9911);
or UO_970 (O_970,N_7555,N_7617);
nor UO_971 (O_971,N_7916,N_9974);
nand UO_972 (O_972,N_9348,N_8414);
xor UO_973 (O_973,N_8732,N_7621);
or UO_974 (O_974,N_8421,N_7598);
and UO_975 (O_975,N_8583,N_7883);
and UO_976 (O_976,N_7662,N_8382);
or UO_977 (O_977,N_9038,N_8486);
and UO_978 (O_978,N_9590,N_9667);
xnor UO_979 (O_979,N_9407,N_9187);
and UO_980 (O_980,N_9794,N_8901);
nand UO_981 (O_981,N_7699,N_8493);
and UO_982 (O_982,N_9066,N_8302);
and UO_983 (O_983,N_8245,N_8343);
xor UO_984 (O_984,N_9387,N_9770);
nor UO_985 (O_985,N_9300,N_9285);
and UO_986 (O_986,N_8083,N_8753);
nand UO_987 (O_987,N_7567,N_8392);
nor UO_988 (O_988,N_7996,N_9213);
or UO_989 (O_989,N_9372,N_7560);
xnor UO_990 (O_990,N_8605,N_9079);
nand UO_991 (O_991,N_8866,N_8944);
xnor UO_992 (O_992,N_8028,N_9946);
or UO_993 (O_993,N_9964,N_7655);
nand UO_994 (O_994,N_9725,N_9722);
or UO_995 (O_995,N_9356,N_8809);
and UO_996 (O_996,N_9968,N_7816);
nand UO_997 (O_997,N_9651,N_8228);
or UO_998 (O_998,N_8532,N_9188);
nand UO_999 (O_999,N_8676,N_9664);
and UO_1000 (O_1000,N_9147,N_7716);
and UO_1001 (O_1001,N_9526,N_8652);
nor UO_1002 (O_1002,N_9611,N_9983);
and UO_1003 (O_1003,N_7887,N_7851);
or UO_1004 (O_1004,N_8941,N_9501);
nand UO_1005 (O_1005,N_8456,N_9445);
nor UO_1006 (O_1006,N_8191,N_8151);
or UO_1007 (O_1007,N_8405,N_7750);
nand UO_1008 (O_1008,N_8759,N_8503);
and UO_1009 (O_1009,N_9965,N_8661);
or UO_1010 (O_1010,N_8610,N_7538);
and UO_1011 (O_1011,N_9883,N_8034);
nor UO_1012 (O_1012,N_9283,N_8196);
nor UO_1013 (O_1013,N_8576,N_8636);
and UO_1014 (O_1014,N_9982,N_8193);
nor UO_1015 (O_1015,N_7679,N_9345);
nor UO_1016 (O_1016,N_9748,N_7989);
nor UO_1017 (O_1017,N_9739,N_8453);
or UO_1018 (O_1018,N_8331,N_9820);
nor UO_1019 (O_1019,N_9100,N_9218);
nand UO_1020 (O_1020,N_9531,N_8711);
and UO_1021 (O_1021,N_7945,N_9800);
or UO_1022 (O_1022,N_8093,N_8829);
nor UO_1023 (O_1023,N_7615,N_9775);
or UO_1024 (O_1024,N_9360,N_7689);
and UO_1025 (O_1025,N_8645,N_7956);
or UO_1026 (O_1026,N_9162,N_9870);
nand UO_1027 (O_1027,N_8685,N_9698);
and UO_1028 (O_1028,N_7624,N_9894);
nand UO_1029 (O_1029,N_9312,N_8035);
and UO_1030 (O_1030,N_9570,N_9971);
nor UO_1031 (O_1031,N_8497,N_9657);
and UO_1032 (O_1032,N_9091,N_8592);
or UO_1033 (O_1033,N_9119,N_8033);
and UO_1034 (O_1034,N_9784,N_9036);
nand UO_1035 (O_1035,N_8773,N_9543);
xnor UO_1036 (O_1036,N_8002,N_9902);
nand UO_1037 (O_1037,N_8357,N_9027);
and UO_1038 (O_1038,N_8631,N_9480);
nor UO_1039 (O_1039,N_8934,N_8634);
nand UO_1040 (O_1040,N_9561,N_8622);
or UO_1041 (O_1041,N_9798,N_8669);
nand UO_1042 (O_1042,N_8907,N_9900);
nand UO_1043 (O_1043,N_7676,N_9029);
nand UO_1044 (O_1044,N_9228,N_9528);
nand UO_1045 (O_1045,N_9903,N_7512);
and UO_1046 (O_1046,N_8942,N_9268);
xnor UO_1047 (O_1047,N_9275,N_7952);
or UO_1048 (O_1048,N_9385,N_8643);
or UO_1049 (O_1049,N_8496,N_9929);
and UO_1050 (O_1050,N_9180,N_8137);
nor UO_1051 (O_1051,N_7904,N_9728);
nor UO_1052 (O_1052,N_8079,N_7642);
nand UO_1053 (O_1053,N_8722,N_9026);
xor UO_1054 (O_1054,N_9309,N_7939);
or UO_1055 (O_1055,N_9814,N_8522);
nand UO_1056 (O_1056,N_7605,N_7748);
nor UO_1057 (O_1057,N_8571,N_7983);
or UO_1058 (O_1058,N_9198,N_7647);
xnor UO_1059 (O_1059,N_8315,N_8994);
nand UO_1060 (O_1060,N_7558,N_8950);
and UO_1061 (O_1061,N_9703,N_9278);
and UO_1062 (O_1062,N_9135,N_9653);
and UO_1063 (O_1063,N_7669,N_7929);
nand UO_1064 (O_1064,N_9624,N_7937);
or UO_1065 (O_1065,N_8819,N_8775);
nand UO_1066 (O_1066,N_8308,N_9481);
nand UO_1067 (O_1067,N_9563,N_9861);
nand UO_1068 (O_1068,N_7806,N_8133);
nor UO_1069 (O_1069,N_9473,N_8556);
nor UO_1070 (O_1070,N_8283,N_8024);
or UO_1071 (O_1071,N_8537,N_9688);
or UO_1072 (O_1072,N_8473,N_9634);
or UO_1073 (O_1073,N_9458,N_7762);
and UO_1074 (O_1074,N_9247,N_9509);
nor UO_1075 (O_1075,N_8363,N_9171);
nor UO_1076 (O_1076,N_9852,N_9576);
nand UO_1077 (O_1077,N_8185,N_8318);
nor UO_1078 (O_1078,N_7700,N_9574);
nand UO_1079 (O_1079,N_8427,N_8826);
nor UO_1080 (O_1080,N_8481,N_8059);
and UO_1081 (O_1081,N_9288,N_8890);
and UO_1082 (O_1082,N_7597,N_9246);
nand UO_1083 (O_1083,N_8282,N_8247);
nand UO_1084 (O_1084,N_9672,N_8956);
or UO_1085 (O_1085,N_8617,N_9789);
or UO_1086 (O_1086,N_7741,N_7671);
and UO_1087 (O_1087,N_8850,N_7695);
nor UO_1088 (O_1088,N_9773,N_7694);
xnor UO_1089 (O_1089,N_7678,N_8810);
nand UO_1090 (O_1090,N_8988,N_9920);
nand UO_1091 (O_1091,N_8214,N_8796);
nor UO_1092 (O_1092,N_8811,N_8886);
nand UO_1093 (O_1093,N_7722,N_7944);
nor UO_1094 (O_1094,N_9631,N_8161);
and UO_1095 (O_1095,N_8255,N_9361);
nor UO_1096 (O_1096,N_8913,N_9035);
nand UO_1097 (O_1097,N_9138,N_8702);
xor UO_1098 (O_1098,N_9743,N_8925);
or UO_1099 (O_1099,N_9379,N_9131);
and UO_1100 (O_1100,N_7517,N_7553);
or UO_1101 (O_1101,N_7677,N_9128);
and UO_1102 (O_1102,N_8295,N_9337);
or UO_1103 (O_1103,N_8670,N_9313);
nand UO_1104 (O_1104,N_9791,N_8474);
or UO_1105 (O_1105,N_9332,N_8010);
and UO_1106 (O_1106,N_9310,N_9311);
and UO_1107 (O_1107,N_8163,N_9229);
nor UO_1108 (O_1108,N_9255,N_9234);
nand UO_1109 (O_1109,N_8401,N_8314);
or UO_1110 (O_1110,N_7928,N_9071);
or UO_1111 (O_1111,N_7726,N_9620);
nand UO_1112 (O_1112,N_9523,N_8080);
or UO_1113 (O_1113,N_9305,N_8173);
nor UO_1114 (O_1114,N_9244,N_8037);
nor UO_1115 (O_1115,N_7638,N_8353);
or UO_1116 (O_1116,N_8061,N_8856);
nand UO_1117 (O_1117,N_7667,N_9468);
and UO_1118 (O_1118,N_9918,N_7552);
or UO_1119 (O_1119,N_7829,N_8065);
and UO_1120 (O_1120,N_7991,N_8555);
or UO_1121 (O_1121,N_8627,N_7788);
or UO_1122 (O_1122,N_8857,N_9488);
nor UO_1123 (O_1123,N_8217,N_9699);
and UO_1124 (O_1124,N_9838,N_9295);
nand UO_1125 (O_1125,N_8591,N_8787);
and UO_1126 (O_1126,N_9972,N_8539);
and UO_1127 (O_1127,N_9890,N_8321);
and UO_1128 (O_1128,N_9762,N_7872);
and UO_1129 (O_1129,N_9658,N_8341);
nor UO_1130 (O_1130,N_9987,N_8858);
or UO_1131 (O_1131,N_9208,N_7501);
nor UO_1132 (O_1132,N_7805,N_9263);
and UO_1133 (O_1133,N_8671,N_8430);
nor UO_1134 (O_1134,N_9303,N_8750);
and UO_1135 (O_1135,N_8319,N_9799);
and UO_1136 (O_1136,N_8916,N_9081);
nand UO_1137 (O_1137,N_7813,N_9237);
nor UO_1138 (O_1138,N_9461,N_9409);
and UO_1139 (O_1139,N_7775,N_8563);
and UO_1140 (O_1140,N_8814,N_9744);
or UO_1141 (O_1141,N_9154,N_9772);
nor UO_1142 (O_1142,N_7742,N_9074);
nor UO_1143 (O_1143,N_7718,N_8258);
nand UO_1144 (O_1144,N_9810,N_8086);
and UO_1145 (O_1145,N_8657,N_9749);
xor UO_1146 (O_1146,N_7973,N_8761);
and UO_1147 (O_1147,N_9235,N_9926);
nand UO_1148 (O_1148,N_8838,N_7528);
and UO_1149 (O_1149,N_8822,N_7562);
nor UO_1150 (O_1150,N_9768,N_8005);
or UO_1151 (O_1151,N_9984,N_8275);
or UO_1152 (O_1152,N_7765,N_7758);
nor UO_1153 (O_1153,N_9795,N_8291);
and UO_1154 (O_1154,N_9845,N_7848);
nand UO_1155 (O_1155,N_8585,N_8416);
nand UO_1156 (O_1156,N_8417,N_7854);
or UO_1157 (O_1157,N_7876,N_7924);
and UO_1158 (O_1158,N_8784,N_9641);
and UO_1159 (O_1159,N_9782,N_7527);
xnor UO_1160 (O_1160,N_8135,N_9788);
nand UO_1161 (O_1161,N_7912,N_9080);
nor UO_1162 (O_1162,N_9904,N_8872);
nand UO_1163 (O_1163,N_7901,N_8089);
and UO_1164 (O_1164,N_8903,N_7706);
and UO_1165 (O_1165,N_9363,N_8051);
nor UO_1166 (O_1166,N_7774,N_7753);
nand UO_1167 (O_1167,N_8499,N_7645);
nand UO_1168 (O_1168,N_8562,N_8244);
and UO_1169 (O_1169,N_7639,N_8612);
nor UO_1170 (O_1170,N_8371,N_8888);
or UO_1171 (O_1171,N_9648,N_7787);
nor UO_1172 (O_1172,N_8688,N_8157);
or UO_1173 (O_1173,N_7507,N_9335);
and UO_1174 (O_1174,N_9999,N_9879);
nor UO_1175 (O_1175,N_7997,N_7941);
nand UO_1176 (O_1176,N_8269,N_9934);
nor UO_1177 (O_1177,N_7725,N_9549);
nand UO_1178 (O_1178,N_7954,N_7618);
nor UO_1179 (O_1179,N_9151,N_8894);
nor UO_1180 (O_1180,N_8943,N_9777);
nand UO_1181 (O_1181,N_8581,N_8547);
nand UO_1182 (O_1182,N_8572,N_8896);
nor UO_1183 (O_1183,N_8640,N_9060);
xor UO_1184 (O_1184,N_9930,N_8337);
nor UO_1185 (O_1185,N_9111,N_8335);
and UO_1186 (O_1186,N_8756,N_7862);
nand UO_1187 (O_1187,N_8625,N_8332);
nor UO_1188 (O_1188,N_8880,N_7981);
nor UO_1189 (O_1189,N_8118,N_9085);
nand UO_1190 (O_1190,N_9326,N_8948);
nand UO_1191 (O_1191,N_8595,N_7866);
and UO_1192 (O_1192,N_9429,N_8527);
xnor UO_1193 (O_1193,N_8791,N_9301);
nor UO_1194 (O_1194,N_9478,N_7660);
or UO_1195 (O_1195,N_7979,N_9207);
and UO_1196 (O_1196,N_9555,N_8719);
nor UO_1197 (O_1197,N_9853,N_8513);
or UO_1198 (O_1198,N_8492,N_8835);
or UO_1199 (O_1199,N_7751,N_8802);
and UO_1200 (O_1200,N_7563,N_8354);
or UO_1201 (O_1201,N_9610,N_8803);
or UO_1202 (O_1202,N_8476,N_7841);
or UO_1203 (O_1203,N_8442,N_9388);
xor UO_1204 (O_1204,N_8737,N_9786);
xnor UO_1205 (O_1205,N_7827,N_9469);
xor UO_1206 (O_1206,N_9215,N_9358);
nand UO_1207 (O_1207,N_9915,N_8932);
xor UO_1208 (O_1208,N_7920,N_9650);
and UO_1209 (O_1209,N_9780,N_8389);
xor UO_1210 (O_1210,N_7794,N_9382);
xnor UO_1211 (O_1211,N_7509,N_8889);
and UO_1212 (O_1212,N_9790,N_8515);
nor UO_1213 (O_1213,N_8980,N_8904);
nor UO_1214 (O_1214,N_7847,N_9754);
or UO_1215 (O_1215,N_9808,N_9086);
nand UO_1216 (O_1216,N_8410,N_9130);
nand UO_1217 (O_1217,N_9320,N_8484);
and UO_1218 (O_1218,N_7661,N_7760);
or UO_1219 (O_1219,N_9392,N_7585);
and UO_1220 (O_1220,N_8383,N_8396);
nand UO_1221 (O_1221,N_7511,N_8900);
and UO_1222 (O_1222,N_9211,N_9977);
xnor UO_1223 (O_1223,N_8875,N_8287);
or UO_1224 (O_1224,N_7888,N_8729);
and UO_1225 (O_1225,N_7596,N_7575);
or UO_1226 (O_1226,N_8853,N_8044);
and UO_1227 (O_1227,N_8358,N_9089);
xnor UO_1228 (O_1228,N_8862,N_8292);
nand UO_1229 (O_1229,N_7976,N_8952);
nand UO_1230 (O_1230,N_8764,N_8144);
nand UO_1231 (O_1231,N_9677,N_9991);
and UO_1232 (O_1232,N_9825,N_7830);
or UO_1233 (O_1233,N_7505,N_8407);
nand UO_1234 (O_1234,N_9096,N_9375);
and UO_1235 (O_1235,N_7988,N_7881);
or UO_1236 (O_1236,N_9818,N_9587);
xnor UO_1237 (O_1237,N_9050,N_8743);
nand UO_1238 (O_1238,N_8087,N_9391);
nor UO_1239 (O_1239,N_8929,N_7935);
nand UO_1240 (O_1240,N_8825,N_9560);
xor UO_1241 (O_1241,N_8064,N_9123);
xor UO_1242 (O_1242,N_9117,N_9767);
xor UO_1243 (O_1243,N_8126,N_8285);
nand UO_1244 (O_1244,N_8348,N_8180);
and UO_1245 (O_1245,N_8181,N_8304);
nor UO_1246 (O_1246,N_9793,N_8177);
nand UO_1247 (O_1247,N_7587,N_7994);
nand UO_1248 (O_1248,N_8962,N_9344);
nor UO_1249 (O_1249,N_8112,N_9868);
nand UO_1250 (O_1250,N_8812,N_9032);
or UO_1251 (O_1251,N_9053,N_8456);
nor UO_1252 (O_1252,N_7730,N_9857);
xor UO_1253 (O_1253,N_7694,N_9913);
nand UO_1254 (O_1254,N_8351,N_8227);
nor UO_1255 (O_1255,N_8098,N_7745);
or UO_1256 (O_1256,N_9550,N_8616);
and UO_1257 (O_1257,N_9376,N_9015);
and UO_1258 (O_1258,N_9080,N_8660);
xnor UO_1259 (O_1259,N_9243,N_8933);
or UO_1260 (O_1260,N_8750,N_8629);
or UO_1261 (O_1261,N_8155,N_8631);
nand UO_1262 (O_1262,N_8138,N_9139);
and UO_1263 (O_1263,N_9530,N_9492);
or UO_1264 (O_1264,N_9730,N_9620);
nand UO_1265 (O_1265,N_8932,N_9170);
or UO_1266 (O_1266,N_9652,N_9522);
and UO_1267 (O_1267,N_8903,N_9299);
xnor UO_1268 (O_1268,N_8961,N_9834);
or UO_1269 (O_1269,N_8517,N_8646);
or UO_1270 (O_1270,N_9595,N_9169);
and UO_1271 (O_1271,N_8293,N_8594);
nor UO_1272 (O_1272,N_8960,N_9133);
and UO_1273 (O_1273,N_9241,N_8745);
nand UO_1274 (O_1274,N_9492,N_7676);
and UO_1275 (O_1275,N_8913,N_8066);
or UO_1276 (O_1276,N_7790,N_8245);
and UO_1277 (O_1277,N_9789,N_9465);
or UO_1278 (O_1278,N_9015,N_8221);
xor UO_1279 (O_1279,N_9054,N_9127);
and UO_1280 (O_1280,N_9995,N_7964);
nand UO_1281 (O_1281,N_8665,N_9782);
and UO_1282 (O_1282,N_7670,N_7704);
and UO_1283 (O_1283,N_8257,N_9199);
nand UO_1284 (O_1284,N_9275,N_8662);
nor UO_1285 (O_1285,N_8060,N_8072);
nand UO_1286 (O_1286,N_8444,N_8848);
or UO_1287 (O_1287,N_7563,N_9575);
nor UO_1288 (O_1288,N_7636,N_7897);
and UO_1289 (O_1289,N_9984,N_9490);
and UO_1290 (O_1290,N_8790,N_8981);
or UO_1291 (O_1291,N_9641,N_7705);
and UO_1292 (O_1292,N_9235,N_8239);
xnor UO_1293 (O_1293,N_9946,N_8404);
or UO_1294 (O_1294,N_8543,N_8288);
or UO_1295 (O_1295,N_7851,N_8095);
and UO_1296 (O_1296,N_7754,N_9129);
nand UO_1297 (O_1297,N_8438,N_9294);
nand UO_1298 (O_1298,N_9702,N_9785);
and UO_1299 (O_1299,N_8659,N_9641);
xnor UO_1300 (O_1300,N_7551,N_8463);
or UO_1301 (O_1301,N_9939,N_7614);
nor UO_1302 (O_1302,N_9234,N_9559);
or UO_1303 (O_1303,N_7845,N_9973);
nor UO_1304 (O_1304,N_7659,N_7858);
nand UO_1305 (O_1305,N_9516,N_8806);
and UO_1306 (O_1306,N_9175,N_8087);
nand UO_1307 (O_1307,N_9598,N_8377);
xor UO_1308 (O_1308,N_7751,N_9029);
or UO_1309 (O_1309,N_8756,N_7619);
nor UO_1310 (O_1310,N_8146,N_7507);
and UO_1311 (O_1311,N_9472,N_8365);
and UO_1312 (O_1312,N_8679,N_8366);
or UO_1313 (O_1313,N_7533,N_8210);
xnor UO_1314 (O_1314,N_8210,N_9291);
or UO_1315 (O_1315,N_8616,N_8163);
xnor UO_1316 (O_1316,N_8694,N_9296);
nor UO_1317 (O_1317,N_9349,N_7821);
nor UO_1318 (O_1318,N_9310,N_8455);
and UO_1319 (O_1319,N_9838,N_9984);
nand UO_1320 (O_1320,N_9446,N_8430);
nor UO_1321 (O_1321,N_8725,N_9892);
and UO_1322 (O_1322,N_9162,N_7814);
nor UO_1323 (O_1323,N_7966,N_7642);
and UO_1324 (O_1324,N_8788,N_9399);
nor UO_1325 (O_1325,N_9193,N_8468);
and UO_1326 (O_1326,N_9498,N_9961);
xor UO_1327 (O_1327,N_9748,N_9251);
nor UO_1328 (O_1328,N_8766,N_7554);
and UO_1329 (O_1329,N_8000,N_9721);
nor UO_1330 (O_1330,N_7567,N_8425);
nor UO_1331 (O_1331,N_9733,N_9174);
nand UO_1332 (O_1332,N_7579,N_7634);
or UO_1333 (O_1333,N_8196,N_7977);
and UO_1334 (O_1334,N_9934,N_8181);
xnor UO_1335 (O_1335,N_9032,N_7889);
nand UO_1336 (O_1336,N_9215,N_8627);
nand UO_1337 (O_1337,N_7980,N_7755);
xor UO_1338 (O_1338,N_8165,N_9820);
and UO_1339 (O_1339,N_9964,N_7521);
nand UO_1340 (O_1340,N_8904,N_8347);
nand UO_1341 (O_1341,N_8507,N_9813);
and UO_1342 (O_1342,N_8959,N_8279);
and UO_1343 (O_1343,N_9117,N_9860);
and UO_1344 (O_1344,N_8200,N_7557);
or UO_1345 (O_1345,N_7896,N_9071);
nand UO_1346 (O_1346,N_9688,N_8328);
nand UO_1347 (O_1347,N_8028,N_9407);
or UO_1348 (O_1348,N_9822,N_9613);
xnor UO_1349 (O_1349,N_9811,N_9078);
or UO_1350 (O_1350,N_8018,N_9565);
or UO_1351 (O_1351,N_8530,N_8195);
nor UO_1352 (O_1352,N_8191,N_7721);
nand UO_1353 (O_1353,N_8160,N_7855);
nand UO_1354 (O_1354,N_8548,N_8321);
nand UO_1355 (O_1355,N_9818,N_8578);
xor UO_1356 (O_1356,N_8691,N_8148);
and UO_1357 (O_1357,N_9213,N_8460);
nor UO_1358 (O_1358,N_9457,N_8501);
or UO_1359 (O_1359,N_9780,N_9122);
and UO_1360 (O_1360,N_7833,N_7504);
or UO_1361 (O_1361,N_7776,N_8166);
or UO_1362 (O_1362,N_8459,N_8845);
and UO_1363 (O_1363,N_8516,N_9445);
nor UO_1364 (O_1364,N_8403,N_9248);
nor UO_1365 (O_1365,N_9089,N_9811);
or UO_1366 (O_1366,N_9179,N_9598);
and UO_1367 (O_1367,N_9716,N_7537);
and UO_1368 (O_1368,N_8007,N_8030);
nand UO_1369 (O_1369,N_8035,N_7969);
or UO_1370 (O_1370,N_8399,N_7664);
nor UO_1371 (O_1371,N_8853,N_9563);
or UO_1372 (O_1372,N_9630,N_9107);
or UO_1373 (O_1373,N_9316,N_9242);
nand UO_1374 (O_1374,N_8898,N_9558);
nand UO_1375 (O_1375,N_8180,N_8303);
nand UO_1376 (O_1376,N_9216,N_8574);
and UO_1377 (O_1377,N_7646,N_8976);
or UO_1378 (O_1378,N_9970,N_8597);
xnor UO_1379 (O_1379,N_7608,N_8763);
and UO_1380 (O_1380,N_8815,N_8803);
nor UO_1381 (O_1381,N_9106,N_7714);
nor UO_1382 (O_1382,N_7696,N_9937);
and UO_1383 (O_1383,N_8279,N_8488);
nor UO_1384 (O_1384,N_9255,N_9588);
and UO_1385 (O_1385,N_8469,N_8246);
nand UO_1386 (O_1386,N_9785,N_9225);
nor UO_1387 (O_1387,N_7900,N_8154);
nand UO_1388 (O_1388,N_8299,N_8327);
nor UO_1389 (O_1389,N_8441,N_8156);
nor UO_1390 (O_1390,N_8559,N_9511);
or UO_1391 (O_1391,N_9766,N_8277);
nand UO_1392 (O_1392,N_7959,N_8000);
or UO_1393 (O_1393,N_8728,N_8243);
nor UO_1394 (O_1394,N_8209,N_8003);
nand UO_1395 (O_1395,N_9684,N_8437);
xor UO_1396 (O_1396,N_8729,N_9888);
nand UO_1397 (O_1397,N_7959,N_7624);
and UO_1398 (O_1398,N_9822,N_9168);
nor UO_1399 (O_1399,N_8616,N_8061);
nor UO_1400 (O_1400,N_9512,N_9040);
or UO_1401 (O_1401,N_7568,N_8172);
nor UO_1402 (O_1402,N_9742,N_8241);
nor UO_1403 (O_1403,N_7752,N_8566);
and UO_1404 (O_1404,N_9152,N_9416);
or UO_1405 (O_1405,N_8567,N_9530);
nand UO_1406 (O_1406,N_9537,N_8450);
nor UO_1407 (O_1407,N_8078,N_9155);
or UO_1408 (O_1408,N_9750,N_9862);
nor UO_1409 (O_1409,N_9132,N_9250);
nor UO_1410 (O_1410,N_9988,N_9737);
nor UO_1411 (O_1411,N_9683,N_8338);
or UO_1412 (O_1412,N_9847,N_9265);
nor UO_1413 (O_1413,N_9131,N_9442);
nor UO_1414 (O_1414,N_8400,N_8767);
xor UO_1415 (O_1415,N_7522,N_8832);
or UO_1416 (O_1416,N_7848,N_8977);
and UO_1417 (O_1417,N_9530,N_8013);
nor UO_1418 (O_1418,N_9330,N_7788);
or UO_1419 (O_1419,N_8882,N_9537);
nor UO_1420 (O_1420,N_9662,N_7908);
or UO_1421 (O_1421,N_7671,N_9387);
and UO_1422 (O_1422,N_8329,N_9475);
nand UO_1423 (O_1423,N_8732,N_8218);
and UO_1424 (O_1424,N_8538,N_8151);
nor UO_1425 (O_1425,N_8041,N_8303);
nor UO_1426 (O_1426,N_8793,N_8611);
nand UO_1427 (O_1427,N_9460,N_9215);
and UO_1428 (O_1428,N_7887,N_9625);
nor UO_1429 (O_1429,N_8946,N_9179);
nand UO_1430 (O_1430,N_7997,N_9846);
xor UO_1431 (O_1431,N_8263,N_9434);
or UO_1432 (O_1432,N_9060,N_8923);
and UO_1433 (O_1433,N_8334,N_8808);
or UO_1434 (O_1434,N_8164,N_8660);
and UO_1435 (O_1435,N_7708,N_8523);
nand UO_1436 (O_1436,N_8309,N_8369);
and UO_1437 (O_1437,N_9807,N_9469);
or UO_1438 (O_1438,N_9031,N_7726);
nand UO_1439 (O_1439,N_9763,N_8752);
nor UO_1440 (O_1440,N_8497,N_9627);
and UO_1441 (O_1441,N_9185,N_8851);
nor UO_1442 (O_1442,N_8660,N_7646);
nand UO_1443 (O_1443,N_8621,N_7905);
or UO_1444 (O_1444,N_7652,N_7764);
nand UO_1445 (O_1445,N_8376,N_9330);
or UO_1446 (O_1446,N_9283,N_8939);
nand UO_1447 (O_1447,N_8978,N_9064);
xor UO_1448 (O_1448,N_8645,N_9737);
or UO_1449 (O_1449,N_9151,N_7539);
xnor UO_1450 (O_1450,N_9993,N_9634);
nand UO_1451 (O_1451,N_8372,N_9712);
or UO_1452 (O_1452,N_9362,N_7531);
or UO_1453 (O_1453,N_8338,N_7690);
nor UO_1454 (O_1454,N_9280,N_9264);
xor UO_1455 (O_1455,N_9979,N_7785);
or UO_1456 (O_1456,N_9166,N_9825);
nor UO_1457 (O_1457,N_7941,N_9750);
or UO_1458 (O_1458,N_9237,N_8140);
nand UO_1459 (O_1459,N_8268,N_7934);
nand UO_1460 (O_1460,N_7515,N_9295);
nand UO_1461 (O_1461,N_8298,N_7848);
nor UO_1462 (O_1462,N_7527,N_9593);
nand UO_1463 (O_1463,N_8239,N_7535);
xor UO_1464 (O_1464,N_9612,N_9998);
nand UO_1465 (O_1465,N_8867,N_9769);
nor UO_1466 (O_1466,N_7694,N_7898);
nand UO_1467 (O_1467,N_9592,N_8411);
or UO_1468 (O_1468,N_8617,N_8133);
nor UO_1469 (O_1469,N_8659,N_8558);
nor UO_1470 (O_1470,N_7887,N_7847);
xnor UO_1471 (O_1471,N_7722,N_8616);
and UO_1472 (O_1472,N_9822,N_7957);
nor UO_1473 (O_1473,N_8448,N_9711);
nor UO_1474 (O_1474,N_9652,N_9348);
and UO_1475 (O_1475,N_9054,N_7590);
nor UO_1476 (O_1476,N_7982,N_9396);
or UO_1477 (O_1477,N_7554,N_7677);
or UO_1478 (O_1478,N_8291,N_9880);
xnor UO_1479 (O_1479,N_8832,N_9379);
xnor UO_1480 (O_1480,N_9234,N_9912);
nand UO_1481 (O_1481,N_9614,N_8049);
and UO_1482 (O_1482,N_8772,N_9611);
xnor UO_1483 (O_1483,N_9794,N_9456);
and UO_1484 (O_1484,N_7573,N_9038);
nor UO_1485 (O_1485,N_8290,N_8882);
or UO_1486 (O_1486,N_8739,N_9875);
xor UO_1487 (O_1487,N_8253,N_9572);
or UO_1488 (O_1488,N_8797,N_8900);
and UO_1489 (O_1489,N_8182,N_8347);
nor UO_1490 (O_1490,N_7748,N_7939);
nor UO_1491 (O_1491,N_7639,N_9494);
or UO_1492 (O_1492,N_9777,N_8376);
xnor UO_1493 (O_1493,N_7802,N_7600);
nand UO_1494 (O_1494,N_7538,N_8048);
and UO_1495 (O_1495,N_8846,N_9986);
xnor UO_1496 (O_1496,N_9495,N_8356);
nor UO_1497 (O_1497,N_9343,N_7768);
nor UO_1498 (O_1498,N_9507,N_7964);
and UO_1499 (O_1499,N_9772,N_9296);
endmodule