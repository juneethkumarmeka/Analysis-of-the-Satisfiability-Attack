module basic_1000_10000_1500_100_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_23,In_325);
and U1 (N_1,In_778,In_27);
or U2 (N_2,In_434,In_558);
or U3 (N_3,In_285,In_368);
xor U4 (N_4,In_846,In_810);
or U5 (N_5,In_79,In_469);
xnor U6 (N_6,In_808,In_101);
or U7 (N_7,In_960,In_897);
nor U8 (N_8,In_315,In_196);
and U9 (N_9,In_605,In_984);
or U10 (N_10,In_94,In_68);
or U11 (N_11,In_208,In_979);
and U12 (N_12,In_474,In_87);
and U13 (N_13,In_35,In_338);
nand U14 (N_14,In_649,In_982);
nand U15 (N_15,In_924,In_981);
xnor U16 (N_16,In_277,In_383);
nand U17 (N_17,In_248,In_552);
and U18 (N_18,In_917,In_871);
xor U19 (N_19,In_115,In_849);
nand U20 (N_20,In_146,In_840);
nor U21 (N_21,In_36,In_843);
and U22 (N_22,In_501,In_63);
xor U23 (N_23,In_859,In_42);
nor U24 (N_24,In_75,In_936);
or U25 (N_25,In_668,In_420);
and U26 (N_26,In_58,In_449);
nor U27 (N_27,In_491,In_541);
or U28 (N_28,In_902,In_390);
nor U29 (N_29,In_529,In_784);
xnor U30 (N_30,In_166,In_522);
or U31 (N_31,In_956,In_402);
nor U32 (N_32,In_763,In_573);
xor U33 (N_33,In_895,In_354);
and U34 (N_34,In_701,In_143);
and U35 (N_35,In_953,In_199);
nor U36 (N_36,In_355,In_439);
or U37 (N_37,In_119,In_246);
or U38 (N_38,In_891,In_329);
nand U39 (N_39,In_811,In_665);
nand U40 (N_40,In_819,In_813);
xnor U41 (N_41,In_992,In_168);
and U42 (N_42,In_386,In_251);
and U43 (N_43,In_661,In_400);
or U44 (N_44,In_935,In_825);
xnor U45 (N_45,In_268,In_84);
or U46 (N_46,In_717,In_190);
xor U47 (N_47,In_603,In_412);
and U48 (N_48,In_393,In_272);
or U49 (N_49,In_644,In_705);
and U50 (N_50,In_687,In_607);
nand U51 (N_51,In_829,In_2);
and U52 (N_52,In_884,In_601);
nor U53 (N_53,In_582,In_271);
or U54 (N_54,In_318,In_815);
and U55 (N_55,In_954,In_711);
and U56 (N_56,In_985,In_228);
xnor U57 (N_57,In_316,In_215);
and U58 (N_58,In_577,In_653);
and U59 (N_59,In_957,In_540);
nor U60 (N_60,In_133,In_926);
and U61 (N_61,In_736,In_40);
or U62 (N_62,In_580,In_1);
or U63 (N_63,In_710,In_882);
and U64 (N_64,In_442,In_150);
nor U65 (N_65,In_578,In_759);
nand U66 (N_66,In_794,In_797);
or U67 (N_67,In_100,In_117);
nor U68 (N_68,In_500,In_174);
nor U69 (N_69,In_423,In_499);
nor U70 (N_70,In_457,In_131);
nand U71 (N_71,In_399,In_10);
or U72 (N_72,In_182,In_427);
xor U73 (N_73,In_546,In_265);
nand U74 (N_74,In_171,In_481);
or U75 (N_75,In_231,In_974);
nand U76 (N_76,In_562,In_911);
nand U77 (N_77,In_809,In_322);
and U78 (N_78,In_113,In_834);
or U79 (N_79,In_421,In_465);
xnor U80 (N_80,In_411,In_255);
and U81 (N_81,In_969,In_309);
nand U82 (N_82,In_323,In_132);
xnor U83 (N_83,In_147,In_127);
nor U84 (N_84,In_638,In_296);
nor U85 (N_85,In_618,In_769);
and U86 (N_86,In_586,In_373);
nor U87 (N_87,In_621,In_494);
nand U88 (N_88,In_302,In_803);
nand U89 (N_89,In_282,In_760);
or U90 (N_90,In_221,In_377);
and U91 (N_91,In_524,In_80);
nand U92 (N_92,In_567,In_581);
nor U93 (N_93,In_291,In_753);
nand U94 (N_94,In_771,In_867);
xnor U95 (N_95,In_996,In_555);
nor U96 (N_96,In_401,In_591);
and U97 (N_97,In_151,In_776);
xnor U98 (N_98,In_725,In_54);
or U99 (N_99,In_361,In_664);
nand U100 (N_100,In_447,In_791);
nand U101 (N_101,In_983,In_173);
xnor U102 (N_102,In_219,In_242);
xor U103 (N_103,In_801,In_209);
and U104 (N_104,In_213,In_340);
or U105 (N_105,In_735,In_631);
xnor U106 (N_106,In_925,In_875);
or U107 (N_107,In_528,In_972);
nor U108 (N_108,In_507,In_37);
or U109 (N_109,In_553,In_304);
or U110 (N_110,In_893,In_184);
or U111 (N_111,In_901,In_237);
or U112 (N_112,In_432,In_7);
and U113 (N_113,In_137,In_907);
and U114 (N_114,In_786,In_627);
xor U115 (N_115,In_415,N_84);
nand U116 (N_116,In_458,In_789);
and U117 (N_117,N_10,In_382);
nor U118 (N_118,In_448,N_93);
nand U119 (N_119,In_623,In_297);
nand U120 (N_120,In_124,In_994);
nand U121 (N_121,In_476,In_886);
nand U122 (N_122,In_545,In_50);
nor U123 (N_123,In_745,In_478);
or U124 (N_124,In_728,In_283);
and U125 (N_125,N_45,In_609);
nor U126 (N_126,In_916,N_4);
and U127 (N_127,In_389,In_772);
nand U128 (N_128,In_189,N_1);
xor U129 (N_129,N_70,In_428);
xor U130 (N_130,In_337,In_155);
nand U131 (N_131,In_977,In_806);
and U132 (N_132,In_21,In_396);
nand U133 (N_133,N_73,In_405);
nor U134 (N_134,In_286,In_645);
and U135 (N_135,N_49,In_874);
nand U136 (N_136,In_372,In_160);
xor U137 (N_137,In_57,In_308);
nand U138 (N_138,In_298,In_163);
xor U139 (N_139,In_986,In_836);
nor U140 (N_140,In_610,In_950);
nand U141 (N_141,In_636,In_656);
xnor U142 (N_142,In_938,In_947);
or U143 (N_143,In_937,In_326);
nor U144 (N_144,In_276,In_464);
nand U145 (N_145,In_12,In_353);
or U146 (N_146,In_556,N_87);
xor U147 (N_147,In_492,In_486);
and U148 (N_148,In_508,In_526);
xnor U149 (N_149,In_203,In_280);
or U150 (N_150,In_637,In_330);
or U151 (N_151,N_97,In_629);
nand U152 (N_152,In_716,In_239);
nor U153 (N_153,In_247,In_970);
and U154 (N_154,In_673,In_862);
and U155 (N_155,In_625,In_820);
xor U156 (N_156,In_165,In_530);
nor U157 (N_157,In_416,In_991);
nand U158 (N_158,In_224,In_669);
or U159 (N_159,In_39,N_88);
or U160 (N_160,N_69,N_55);
and U161 (N_161,In_685,In_112);
nand U162 (N_162,In_358,N_25);
or U163 (N_163,N_89,In_756);
xor U164 (N_164,In_24,In_306);
xor U165 (N_165,In_459,In_410);
nor U166 (N_166,In_134,In_666);
nor U167 (N_167,In_741,In_477);
nand U168 (N_168,In_369,In_520);
xor U169 (N_169,N_53,In_689);
nor U170 (N_170,In_738,N_59);
nand U171 (N_171,In_719,In_453);
and U172 (N_172,N_86,N_48);
nand U173 (N_173,In_480,In_816);
and U174 (N_174,In_890,In_38);
nor U175 (N_175,In_682,In_321);
and U176 (N_176,In_697,In_512);
xnor U177 (N_177,In_896,In_922);
xor U178 (N_178,In_91,In_195);
nand U179 (N_179,In_883,In_128);
or U180 (N_180,In_103,In_44);
xnor U181 (N_181,In_790,In_140);
nor U182 (N_182,In_301,In_903);
xnor U183 (N_183,N_47,In_48);
xnor U184 (N_184,In_595,In_216);
nor U185 (N_185,In_942,In_918);
xnor U186 (N_186,In_232,In_534);
nor U187 (N_187,In_214,In_76);
nand U188 (N_188,In_96,In_805);
and U189 (N_189,In_777,In_571);
nand U190 (N_190,In_225,N_0);
or U191 (N_191,N_51,In_651);
and U192 (N_192,In_273,In_90);
or U193 (N_193,In_192,In_479);
xnor U194 (N_194,In_352,N_39);
xnor U195 (N_195,In_648,In_130);
or U196 (N_196,In_779,N_14);
nor U197 (N_197,In_730,In_380);
nand U198 (N_198,In_443,N_63);
xor U199 (N_199,In_490,In_699);
nor U200 (N_200,In_873,In_718);
or U201 (N_201,In_89,In_948);
xnor U202 (N_202,In_740,N_189);
nand U203 (N_203,In_848,In_142);
nand U204 (N_204,In_197,In_574);
or U205 (N_205,In_906,N_150);
nand U206 (N_206,In_64,In_748);
nor U207 (N_207,N_177,In_927);
and U208 (N_208,In_126,In_109);
xor U209 (N_209,In_894,In_289);
or U210 (N_210,N_116,N_60);
nand U211 (N_211,In_932,In_376);
xnor U212 (N_212,N_151,In_995);
nor U213 (N_213,In_659,N_183);
xor U214 (N_214,In_792,In_519);
xnor U215 (N_215,In_74,In_737);
xnor U216 (N_216,N_2,In_25);
and U217 (N_217,N_129,In_868);
nand U218 (N_218,N_82,In_404);
or U219 (N_219,In_551,In_359);
and U220 (N_220,In_762,In_933);
or U221 (N_221,In_398,In_370);
nor U222 (N_222,In_702,In_498);
xor U223 (N_223,In_654,In_116);
and U224 (N_224,In_59,In_782);
nand U225 (N_225,N_170,In_841);
xor U226 (N_226,In_95,In_712);
nand U227 (N_227,N_126,In_46);
xor U228 (N_228,In_331,In_194);
nor U229 (N_229,In_347,In_920);
xor U230 (N_230,In_125,In_176);
xnor U231 (N_231,In_384,In_505);
nand U232 (N_232,N_43,N_138);
nor U233 (N_233,In_229,In_785);
nor U234 (N_234,In_588,In_915);
and U235 (N_235,In_764,In_278);
nor U236 (N_236,N_58,N_12);
xor U237 (N_237,N_160,In_292);
nand U238 (N_238,In_866,In_523);
xnor U239 (N_239,In_110,N_198);
nand U240 (N_240,In_460,N_147);
or U241 (N_241,In_904,In_709);
and U242 (N_242,In_966,In_622);
and U243 (N_243,In_31,In_341);
nand U244 (N_244,In_138,N_106);
nand U245 (N_245,In_451,In_861);
nand U246 (N_246,In_798,In_706);
xor U247 (N_247,In_345,In_880);
nor U248 (N_248,N_99,In_575);
or U249 (N_249,In_360,In_446);
or U250 (N_250,N_168,In_175);
and U251 (N_251,In_28,In_15);
xor U252 (N_252,In_374,In_830);
nor U253 (N_253,In_43,In_379);
and U254 (N_254,In_703,In_997);
xor U255 (N_255,In_750,In_241);
and U256 (N_256,N_22,N_143);
or U257 (N_257,In_319,In_156);
and U258 (N_258,In_139,In_557);
xor U259 (N_259,In_847,In_869);
or U260 (N_260,In_287,In_263);
and U261 (N_261,In_158,In_532);
nand U262 (N_262,In_4,In_364);
nand U263 (N_263,In_344,In_217);
and U264 (N_264,In_688,In_672);
xnor U265 (N_265,In_721,In_913);
nand U266 (N_266,In_258,In_495);
or U267 (N_267,In_826,In_941);
nor U268 (N_268,In_471,In_245);
and U269 (N_269,In_839,N_139);
nor U270 (N_270,N_104,In_187);
and U271 (N_271,In_842,In_989);
xor U272 (N_272,In_964,In_799);
nor U273 (N_273,In_720,In_889);
and U274 (N_274,In_980,N_64);
and U275 (N_275,In_853,In_732);
and U276 (N_276,In_684,In_441);
xor U277 (N_277,In_647,N_158);
or U278 (N_278,In_397,In_123);
and U279 (N_279,In_739,N_110);
and U280 (N_280,In_742,In_860);
xor U281 (N_281,In_837,In_99);
and U282 (N_282,In_513,In_566);
nand U283 (N_283,In_619,In_722);
and U284 (N_284,In_931,In_32);
nand U285 (N_285,In_250,In_149);
nor U286 (N_286,N_13,In_976);
xor U287 (N_287,In_332,N_9);
and U288 (N_288,In_963,In_34);
xnor U289 (N_289,In_821,In_945);
and U290 (N_290,In_787,In_342);
and U291 (N_291,N_62,In_406);
nor U292 (N_292,In_30,In_53);
nand U293 (N_293,In_41,In_136);
or U294 (N_294,In_657,In_632);
xor U295 (N_295,In_85,N_28);
and U296 (N_296,In_445,In_295);
and U297 (N_297,N_112,In_783);
nand U298 (N_298,In_488,In_559);
nor U299 (N_299,N_197,N_122);
or U300 (N_300,In_536,N_292);
nand U301 (N_301,N_227,In_554);
nand U302 (N_302,In_754,In_310);
xnor U303 (N_303,In_755,In_430);
and U304 (N_304,In_452,In_437);
nor U305 (N_305,N_34,In_456);
and U306 (N_306,N_125,N_258);
or U307 (N_307,N_278,N_268);
nand U308 (N_308,In_392,In_696);
xor U309 (N_309,In_356,In_462);
nor U310 (N_310,In_572,In_497);
or U311 (N_311,N_102,N_5);
and U312 (N_312,In_521,In_346);
nor U313 (N_313,N_295,In_788);
nor U314 (N_314,N_74,N_232);
and U315 (N_315,In_180,N_237);
and U316 (N_316,In_734,N_266);
nand U317 (N_317,In_993,N_15);
xnor U318 (N_318,N_111,In_419);
xnor U319 (N_319,N_220,In_9);
xnor U320 (N_320,N_117,In_371);
nor U321 (N_321,In_563,N_81);
or U322 (N_322,In_262,N_123);
or U323 (N_323,N_293,N_167);
or U324 (N_324,N_297,In_288);
and U325 (N_325,N_115,In_67);
xor U326 (N_326,In_222,N_140);
or U327 (N_327,In_640,In_751);
xor U328 (N_328,N_105,In_978);
or U329 (N_329,N_252,N_79);
or U330 (N_330,In_852,In_293);
xnor U331 (N_331,N_180,In_468);
or U332 (N_332,In_749,In_692);
xnor U333 (N_333,N_178,In_844);
or U334 (N_334,N_289,In_940);
or U335 (N_335,In_13,N_135);
nand U336 (N_336,In_608,N_20);
or U337 (N_337,In_204,N_265);
or U338 (N_338,In_8,In_857);
or U339 (N_339,In_81,N_207);
or U340 (N_340,In_202,N_256);
xor U341 (N_341,N_184,In_724);
xnor U342 (N_342,N_159,In_307);
nand U343 (N_343,In_624,N_272);
nor U344 (N_344,N_98,In_475);
nor U345 (N_345,In_281,In_205);
and U346 (N_346,N_54,In_923);
nor U347 (N_347,In_646,In_425);
xor U348 (N_348,In_333,N_57);
and U349 (N_349,In_865,N_263);
xnor U350 (N_350,In_952,In_678);
or U351 (N_351,In_435,In_570);
nand U352 (N_352,In_141,N_211);
or U353 (N_353,N_208,In_561);
or U354 (N_354,In_851,N_245);
nand U355 (N_355,In_822,In_655);
and U356 (N_356,N_249,N_171);
nand U357 (N_357,In_594,In_921);
xor U358 (N_358,N_222,In_193);
or U359 (N_359,In_19,In_365);
or U360 (N_360,In_450,N_236);
xor U361 (N_361,In_858,In_676);
xnor U362 (N_362,In_517,In_909);
nor U363 (N_363,In_5,N_72);
xnor U364 (N_364,In_29,N_101);
nor U365 (N_365,In_817,N_240);
nor U366 (N_366,In_616,In_814);
xnor U367 (N_367,In_431,N_38);
and U368 (N_368,In_294,In_780);
and U369 (N_369,N_35,N_196);
nand U370 (N_370,In_793,N_44);
or U371 (N_371,In_543,N_201);
nor U372 (N_372,In_157,N_205);
xnor U373 (N_373,In_45,N_66);
nor U374 (N_374,In_206,In_746);
xor U375 (N_375,In_888,In_910);
nand U376 (N_376,In_259,In_378);
xnor U377 (N_377,In_679,In_71);
nand U378 (N_378,In_120,In_872);
or U379 (N_379,In_426,In_877);
nor U380 (N_380,In_691,N_298);
xor U381 (N_381,N_225,N_31);
and U382 (N_382,N_200,In_518);
nand U383 (N_383,In_47,In_856);
and U384 (N_384,In_973,N_109);
nor U385 (N_385,N_223,In_16);
nor U386 (N_386,In_590,N_124);
or U387 (N_387,In_69,N_287);
or U388 (N_388,In_677,N_281);
nor U389 (N_389,In_73,In_261);
nand U390 (N_390,In_930,N_6);
xnor U391 (N_391,In_227,In_381);
nor U392 (N_392,In_284,N_41);
nand U393 (N_393,In_86,In_832);
nand U394 (N_394,N_275,N_192);
nor U395 (N_395,In_695,N_67);
and U396 (N_396,In_804,N_30);
nor U397 (N_397,In_951,In_587);
xor U398 (N_398,In_795,N_19);
or U399 (N_399,In_768,In_639);
and U400 (N_400,N_119,In_223);
nand U401 (N_401,In_823,In_313);
and U402 (N_402,N_359,N_283);
or U403 (N_403,N_257,In_169);
nand U404 (N_404,N_386,In_3);
xnor U405 (N_405,N_279,N_304);
or U406 (N_406,In_33,In_514);
and U407 (N_407,N_230,N_148);
nor U408 (N_408,In_164,In_807);
and U409 (N_409,In_349,N_157);
nor U410 (N_410,N_169,In_919);
nand U411 (N_411,N_288,In_211);
nor U412 (N_412,N_264,In_455);
and U413 (N_413,N_37,N_320);
nand U414 (N_414,In_569,N_203);
nor U415 (N_415,N_362,N_369);
and U416 (N_416,In_683,N_94);
or U417 (N_417,N_188,N_65);
xnor U418 (N_418,N_367,In_885);
or U419 (N_419,In_704,N_376);
or U420 (N_420,N_321,In_417);
nor U421 (N_421,In_114,N_337);
xor U422 (N_422,In_178,In_833);
and U423 (N_423,In_767,In_240);
and U424 (N_424,In_693,N_42);
nor U425 (N_425,In_949,In_968);
nand U426 (N_426,In_118,In_900);
or U427 (N_427,In_60,In_694);
nand U428 (N_428,In_987,In_387);
nor U429 (N_429,N_80,In_934);
or U430 (N_430,In_409,In_98);
and U431 (N_431,In_467,N_68);
nor U432 (N_432,N_92,In_876);
and U433 (N_433,N_343,In_413);
or U434 (N_434,In_312,N_319);
or U435 (N_435,In_348,N_52);
or U436 (N_436,N_233,In_267);
or U437 (N_437,In_958,In_244);
or U438 (N_438,In_599,N_341);
nand U439 (N_439,N_274,In_254);
nand U440 (N_440,N_329,In_105);
nand U441 (N_441,N_113,In_617);
nand U442 (N_442,In_800,N_267);
nor U443 (N_443,In_264,N_7);
and U444 (N_444,In_818,In_314);
nand U445 (N_445,N_389,N_361);
or U446 (N_446,N_399,In_482);
nor U447 (N_447,In_407,In_454);
nor U448 (N_448,N_242,N_378);
xnor U449 (N_449,In_774,N_351);
nand U450 (N_450,N_163,In_824);
nor U451 (N_451,In_812,N_96);
and U452 (N_452,In_320,In_870);
xor U453 (N_453,N_317,In_600);
or U454 (N_454,N_294,N_315);
xnor U455 (N_455,N_259,N_206);
nor U456 (N_456,In_210,N_379);
xnor U457 (N_457,N_149,N_316);
and U458 (N_458,In_388,In_473);
xnor U459 (N_459,N_327,In_614);
or U460 (N_460,In_335,N_356);
or U461 (N_461,In_626,In_510);
xnor U462 (N_462,In_744,N_179);
xnor U463 (N_463,In_106,In_674);
nor U464 (N_464,In_606,In_14);
or U465 (N_465,N_357,In_928);
xnor U466 (N_466,In_6,In_592);
nand U467 (N_467,In_327,N_194);
or U468 (N_468,N_244,In_55);
nand U469 (N_469,N_255,N_210);
xor U470 (N_470,N_365,In_172);
and U471 (N_471,In_233,In_802);
xnor U472 (N_472,N_385,In_878);
nand U473 (N_473,N_56,In_681);
nor U474 (N_474,N_330,In_547);
and U475 (N_475,N_347,In_367);
or U476 (N_476,In_300,In_463);
or U477 (N_477,In_503,In_729);
and U478 (N_478,N_229,N_164);
xnor U479 (N_479,N_366,In_496);
xor U480 (N_480,In_167,In_234);
nor U481 (N_481,In_835,N_243);
nand U482 (N_482,In_181,In_975);
xnor U483 (N_483,N_395,In_633);
or U484 (N_484,In_418,In_212);
or U485 (N_485,In_564,In_715);
xor U486 (N_486,In_568,In_362);
nor U487 (N_487,N_342,In_939);
nor U488 (N_488,In_324,In_667);
nor U489 (N_489,N_374,N_50);
nor U490 (N_490,N_371,In_72);
and U491 (N_491,N_204,In_275);
or U492 (N_492,In_828,In_429);
nand U493 (N_493,In_535,In_515);
nand U494 (N_494,In_864,N_32);
xnor U495 (N_495,N_155,In_88);
or U496 (N_496,N_216,In_727);
nand U497 (N_497,N_326,In_999);
and U498 (N_498,N_107,N_195);
or U499 (N_499,In_148,N_134);
and U500 (N_500,N_485,In_831);
nor U501 (N_501,In_731,In_511);
and U502 (N_502,In_257,In_61);
or U503 (N_503,In_752,In_299);
nor U504 (N_504,In_489,N_479);
nand U505 (N_505,In_611,In_757);
nor U506 (N_506,N_127,In_108);
nand U507 (N_507,In_17,N_146);
nand U508 (N_508,In_414,N_165);
nor U509 (N_509,In_290,N_403);
nand U510 (N_510,N_494,In_579);
nor U511 (N_511,In_576,N_27);
or U512 (N_512,N_120,N_483);
nor U513 (N_513,N_424,N_280);
or U514 (N_514,In_93,In_613);
nand U515 (N_515,N_166,In_177);
nor U516 (N_516,N_300,N_191);
and U517 (N_517,In_122,In_363);
nand U518 (N_518,In_145,N_18);
nor U519 (N_519,In_236,N_335);
nor U520 (N_520,In_854,N_348);
xnor U521 (N_521,N_402,N_85);
and U522 (N_522,N_425,In_733);
and U523 (N_523,N_383,In_218);
and U524 (N_524,In_18,N_473);
or U525 (N_525,N_458,In_170);
nor U526 (N_526,N_446,N_121);
xnor U527 (N_527,N_78,In_887);
nand U528 (N_528,In_726,N_352);
or U529 (N_529,In_403,N_199);
or U530 (N_530,N_380,In_670);
or U531 (N_531,In_690,N_423);
xor U532 (N_532,In_226,N_91);
xor U533 (N_533,In_758,N_349);
and U534 (N_534,N_261,N_33);
xor U535 (N_535,N_75,N_440);
xor U536 (N_536,In_394,N_488);
nor U537 (N_537,N_142,N_460);
and U538 (N_538,In_892,In_533);
xnor U539 (N_539,N_391,N_360);
nor U540 (N_540,N_451,In_107);
nor U541 (N_541,N_492,N_388);
nand U542 (N_542,N_447,In_899);
nand U543 (N_543,N_114,In_642);
and U544 (N_544,N_444,N_95);
nand U545 (N_545,In_97,In_198);
or U546 (N_546,N_273,N_302);
nor U547 (N_547,In_612,In_635);
nor U548 (N_548,N_334,N_482);
nor U549 (N_549,N_418,In_531);
or U550 (N_550,N_414,N_453);
nand U551 (N_551,In_504,In_339);
and U552 (N_552,In_761,N_470);
or U553 (N_553,N_416,N_239);
nand U554 (N_554,N_409,In_183);
nor U555 (N_555,N_152,N_392);
nor U556 (N_556,N_202,In_159);
nand U557 (N_557,N_234,In_351);
nor U558 (N_558,In_946,N_219);
or U559 (N_559,N_368,In_162);
and U560 (N_560,In_336,In_714);
nor U561 (N_561,In_22,In_11);
or U562 (N_562,N_301,N_456);
and U563 (N_563,N_186,In_775);
xnor U564 (N_564,In_845,N_172);
or U565 (N_565,In_484,In_959);
or U566 (N_566,N_382,N_21);
xor U567 (N_567,In_527,In_881);
xor U568 (N_568,N_269,In_444);
nand U569 (N_569,In_207,N_429);
nor U570 (N_570,N_358,N_407);
and U571 (N_571,N_328,N_397);
xor U572 (N_572,N_472,N_307);
nand U573 (N_573,N_305,In_634);
nand U574 (N_574,In_154,In_593);
nor U575 (N_575,In_0,In_83);
nor U576 (N_576,N_24,N_435);
and U577 (N_577,In_270,N_401);
or U578 (N_578,In_967,In_185);
nand U579 (N_579,N_173,In_311);
or U580 (N_580,N_71,In_62);
xor U581 (N_581,N_23,N_221);
or U582 (N_582,N_90,In_466);
and U583 (N_583,In_905,N_254);
nor U584 (N_584,In_585,N_284);
nor U585 (N_585,N_231,In_686);
nor U586 (N_586,N_332,In_509);
xnor U587 (N_587,N_375,N_271);
and U588 (N_588,N_411,N_497);
and U589 (N_589,In_179,In_965);
nor U590 (N_590,In_641,In_944);
and U591 (N_591,N_350,In_537);
nor U592 (N_592,N_285,In_269);
xnor U593 (N_593,N_308,N_226);
nor U594 (N_594,In_596,In_650);
nor U595 (N_595,N_421,N_212);
xnor U596 (N_596,N_214,In_675);
or U597 (N_597,In_20,In_111);
nand U598 (N_598,In_266,N_459);
nand U599 (N_599,N_487,N_465);
nor U600 (N_600,N_322,N_428);
nor U601 (N_601,N_469,N_538);
nor U602 (N_602,N_3,In_671);
or U603 (N_603,In_781,N_137);
and U604 (N_604,In_773,N_570);
nand U605 (N_605,N_8,N_100);
xor U606 (N_606,In_328,In_550);
and U607 (N_607,N_471,N_598);
and U608 (N_608,N_599,In_602);
or U609 (N_609,N_417,N_141);
and U610 (N_610,N_364,In_350);
nand U611 (N_611,N_585,N_291);
xor U612 (N_612,N_431,N_247);
nand U613 (N_613,In_630,In_929);
xor U614 (N_614,N_581,N_387);
or U615 (N_615,In_78,N_390);
or U616 (N_616,N_251,N_467);
nand U617 (N_617,N_16,N_420);
nand U618 (N_618,In_855,N_573);
xor U619 (N_619,N_432,N_248);
nand U620 (N_620,N_299,N_323);
or U621 (N_621,In_615,In_49);
xor U622 (N_622,N_587,In_385);
nand U623 (N_623,In_663,In_82);
nor U624 (N_624,N_346,N_533);
nor U625 (N_625,N_476,N_262);
nand U626 (N_626,N_528,N_503);
xnor U627 (N_627,N_564,N_539);
and U628 (N_628,N_535,N_521);
nand U629 (N_629,N_596,N_238);
nor U630 (N_630,N_597,In_470);
nand U631 (N_631,N_575,In_253);
nor U632 (N_632,In_990,N_185);
nand U633 (N_633,In_539,In_200);
or U634 (N_634,In_971,N_161);
nand U635 (N_635,N_532,N_496);
or U636 (N_636,N_448,In_549);
and U637 (N_637,In_658,N_452);
nand U638 (N_638,In_186,In_962);
nand U639 (N_639,N_540,N_250);
nand U640 (N_640,In_565,N_76);
xnor U641 (N_641,N_400,In_334);
xnor U642 (N_642,N_228,N_515);
xnor U643 (N_643,N_524,N_495);
xnor U644 (N_644,N_569,N_404);
and U645 (N_645,In_827,In_700);
xor U646 (N_646,N_558,N_514);
nand U647 (N_647,In_52,N_193);
and U648 (N_648,In_483,In_998);
and U649 (N_649,N_549,N_541);
nor U650 (N_650,N_209,N_579);
nand U651 (N_651,In_395,N_128);
nand U652 (N_652,N_588,N_118);
and U653 (N_653,In_144,N_235);
nor U654 (N_654,In_317,In_440);
or U655 (N_655,N_486,In_343);
nand U656 (N_656,N_333,N_512);
nand U657 (N_657,In_698,In_485);
nand U658 (N_658,N_11,In_589);
nand U659 (N_659,N_536,N_370);
xor U660 (N_660,In_249,N_354);
xor U661 (N_661,N_422,N_156);
and U662 (N_662,N_393,N_527);
nor U663 (N_663,In_560,In_135);
and U664 (N_664,N_153,N_520);
and U665 (N_665,N_557,In_643);
and U666 (N_666,In_525,In_961);
xnor U667 (N_667,N_439,N_436);
or U668 (N_668,N_270,N_190);
nand U669 (N_669,N_426,In_26);
nor U670 (N_670,In_660,N_176);
nor U671 (N_671,N_463,N_373);
xor U672 (N_672,N_433,N_519);
and U673 (N_673,In_472,N_438);
xor U674 (N_674,In_66,N_577);
xor U675 (N_675,N_490,In_620);
nand U676 (N_676,N_215,N_543);
nor U677 (N_677,N_108,In_102);
or U678 (N_678,N_583,N_449);
nor U679 (N_679,In_220,In_235);
xnor U680 (N_680,N_224,N_309);
nand U681 (N_681,N_545,N_508);
nand U682 (N_682,In_662,In_422);
xnor U683 (N_683,N_477,N_384);
and U684 (N_684,N_415,In_988);
nand U685 (N_685,N_396,In_487);
nor U686 (N_686,N_493,In_766);
and U687 (N_687,N_46,N_574);
nand U688 (N_688,N_312,N_145);
or U689 (N_689,N_518,In_680);
nand U690 (N_690,N_507,In_765);
nand U691 (N_691,N_572,In_628);
xnor U692 (N_692,N_475,N_461);
xor U693 (N_693,N_481,In_201);
nor U694 (N_694,In_230,N_555);
nor U695 (N_695,N_318,In_548);
nand U696 (N_696,N_466,In_912);
nand U697 (N_697,In_770,N_136);
or U698 (N_698,In_274,In_838);
nor U699 (N_699,In_65,N_175);
and U700 (N_700,N_679,In_243);
nand U701 (N_701,N_217,N_530);
nor U702 (N_702,N_614,N_313);
or U703 (N_703,N_688,N_282);
nor U704 (N_704,N_632,In_77);
nor U705 (N_705,N_544,In_70);
xor U706 (N_706,N_556,N_613);
xnor U707 (N_707,N_630,N_83);
nor U708 (N_708,N_562,In_188);
nor U709 (N_709,N_652,N_517);
nor U710 (N_710,N_686,N_260);
xor U711 (N_711,N_601,In_260);
or U712 (N_712,N_509,In_707);
or U713 (N_713,N_504,N_578);
nor U714 (N_714,N_666,N_698);
nand U715 (N_715,N_612,N_676);
nand U716 (N_716,N_670,N_602);
nor U717 (N_717,N_582,In_796);
nand U718 (N_718,N_130,N_408);
and U719 (N_719,In_303,N_568);
or U720 (N_720,N_525,N_668);
or U721 (N_721,N_450,N_639);
nor U722 (N_722,N_553,N_607);
xnor U723 (N_723,N_372,N_419);
or U724 (N_724,N_609,N_468);
xnor U725 (N_725,N_665,N_634);
nor U726 (N_726,N_661,N_547);
nand U727 (N_727,N_516,In_538);
nand U728 (N_728,N_218,In_391);
xor U729 (N_729,N_344,N_616);
xnor U730 (N_730,In_914,In_743);
nor U731 (N_731,N_692,N_590);
nor U732 (N_732,N_636,N_61);
nand U733 (N_733,N_454,N_649);
or U734 (N_734,N_324,N_691);
xor U735 (N_735,In_408,In_438);
nand U736 (N_736,N_484,N_604);
and U737 (N_737,N_241,In_493);
and U738 (N_738,N_561,N_600);
and U739 (N_739,In_747,N_537);
xnor U740 (N_740,N_213,N_611);
nor U741 (N_741,In_191,N_405);
nand U742 (N_742,N_441,N_489);
nor U743 (N_743,N_546,N_667);
xor U744 (N_744,N_394,N_646);
nand U745 (N_745,N_491,N_377);
xnor U746 (N_746,In_955,In_375);
nor U747 (N_747,N_17,N_412);
or U748 (N_748,N_398,In_908);
nand U749 (N_749,N_531,N_689);
nor U750 (N_750,N_606,N_311);
and U751 (N_751,N_656,N_584);
or U752 (N_752,N_336,N_406);
xnor U753 (N_753,N_478,N_499);
xor U754 (N_754,In_161,N_174);
and U755 (N_755,N_310,N_641);
xor U756 (N_756,In_104,In_583);
or U757 (N_757,In_713,In_92);
and U758 (N_758,N_633,In_879);
nand U759 (N_759,N_682,N_563);
nand U760 (N_760,N_353,N_591);
or U761 (N_761,N_621,N_26);
nor U762 (N_762,N_325,N_286);
xor U763 (N_763,N_542,N_339);
and U764 (N_764,N_133,N_510);
nor U765 (N_765,N_306,N_669);
nand U766 (N_766,N_246,N_363);
nand U767 (N_767,N_131,N_523);
xnor U768 (N_768,N_154,N_624);
or U769 (N_769,N_684,N_560);
nand U770 (N_770,In_56,In_305);
nand U771 (N_771,N_464,N_657);
nand U772 (N_772,N_615,In_129);
and U773 (N_773,N_586,N_660);
xnor U774 (N_774,N_511,N_608);
and U775 (N_775,N_655,N_480);
nand U776 (N_776,In_598,N_550);
xor U777 (N_777,N_505,N_434);
nor U778 (N_778,N_699,N_626);
nor U779 (N_779,N_559,N_690);
and U780 (N_780,In_516,N_697);
nand U781 (N_781,In_943,In_279);
xnor U782 (N_782,N_474,In_238);
or U783 (N_783,N_338,N_442);
or U784 (N_784,In_424,N_629);
and U785 (N_785,N_659,N_253);
and U786 (N_786,N_683,N_647);
and U787 (N_787,N_640,N_565);
or U788 (N_788,N_620,N_650);
or U789 (N_789,N_648,N_622);
nor U790 (N_790,N_644,N_455);
xor U791 (N_791,In_461,N_658);
nand U792 (N_792,N_662,In_584);
nor U793 (N_793,In_436,N_462);
or U794 (N_794,In_51,N_277);
or U795 (N_795,In_708,In_723);
nand U796 (N_796,N_355,N_695);
xnor U797 (N_797,N_651,In_152);
nand U798 (N_798,N_296,N_645);
xor U799 (N_799,N_276,N_181);
nor U800 (N_800,In_153,N_710);
or U801 (N_801,N_729,In_604);
xor U802 (N_802,N_642,N_664);
xnor U803 (N_803,N_768,N_747);
nor U804 (N_804,N_654,N_723);
or U805 (N_805,N_603,N_739);
or U806 (N_806,N_605,N_566);
nor U807 (N_807,In_433,In_357);
or U808 (N_808,N_726,N_742);
and U809 (N_809,N_777,N_529);
xnor U810 (N_810,N_303,N_733);
or U811 (N_811,N_671,N_795);
nand U812 (N_812,N_767,N_554);
nand U813 (N_813,N_756,N_314);
nor U814 (N_814,N_781,N_755);
nor U815 (N_815,In_121,N_445);
nor U816 (N_816,N_696,N_787);
xnor U817 (N_817,N_774,N_738);
and U818 (N_818,N_707,N_502);
and U819 (N_819,N_751,N_628);
xor U820 (N_820,N_724,N_498);
or U821 (N_821,N_759,N_782);
or U822 (N_822,N_571,N_430);
nand U823 (N_823,N_745,N_551);
nand U824 (N_824,N_720,N_29);
nor U825 (N_825,N_500,N_731);
nand U826 (N_826,N_773,N_592);
and U827 (N_827,N_427,N_693);
or U828 (N_828,N_716,N_754);
or U829 (N_829,N_182,N_674);
nand U830 (N_830,N_760,N_677);
or U831 (N_831,In_652,N_763);
nand U832 (N_832,N_703,N_706);
nor U833 (N_833,In_597,N_694);
and U834 (N_834,N_709,N_730);
and U835 (N_835,N_721,N_522);
nor U836 (N_836,N_766,N_792);
nand U837 (N_837,N_672,N_761);
and U838 (N_838,N_771,N_663);
or U839 (N_839,N_618,N_595);
xor U840 (N_840,N_701,N_673);
nor U841 (N_841,N_687,N_638);
nand U842 (N_842,N_713,N_758);
xnor U843 (N_843,N_797,N_345);
nand U844 (N_844,N_784,N_743);
nand U845 (N_845,N_714,N_785);
and U846 (N_846,N_750,In_542);
nand U847 (N_847,N_765,N_437);
xor U848 (N_848,N_775,N_788);
nor U849 (N_849,N_746,N_132);
nor U850 (N_850,In_898,N_526);
nor U851 (N_851,N_708,N_769);
nor U852 (N_852,N_741,N_653);
and U853 (N_853,N_552,N_780);
nor U854 (N_854,N_685,N_779);
xnor U855 (N_855,N_799,N_619);
xnor U856 (N_856,N_567,N_711);
and U857 (N_857,N_593,N_744);
and U858 (N_858,In_506,In_366);
or U859 (N_859,In_256,N_762);
nand U860 (N_860,N_790,N_631);
nor U861 (N_861,N_637,N_576);
nor U862 (N_862,N_617,N_625);
and U863 (N_863,N_783,N_681);
and U864 (N_864,N_635,N_36);
and U865 (N_865,N_40,N_798);
xnor U866 (N_866,N_513,N_589);
xnor U867 (N_867,N_700,N_705);
or U868 (N_868,N_702,N_772);
xnor U869 (N_869,N_410,N_725);
and U870 (N_870,N_580,In_502);
nor U871 (N_871,N_717,In_252);
nand U872 (N_872,N_290,N_675);
and U873 (N_873,N_678,N_752);
nor U874 (N_874,N_748,N_770);
and U875 (N_875,N_796,N_340);
nand U876 (N_876,N_753,N_381);
xor U877 (N_877,N_737,N_331);
xnor U878 (N_878,N_735,N_727);
and U879 (N_879,N_740,N_643);
nand U880 (N_880,N_457,N_791);
nand U881 (N_881,N_712,N_610);
and U882 (N_882,N_736,N_144);
and U883 (N_883,N_162,N_786);
or U884 (N_884,N_704,N_719);
and U885 (N_885,N_443,N_506);
xnor U886 (N_886,N_794,In_850);
nand U887 (N_887,N_789,N_793);
xnor U888 (N_888,N_501,N_103);
xor U889 (N_889,N_749,N_548);
and U890 (N_890,N_413,N_623);
or U891 (N_891,In_863,N_627);
or U892 (N_892,N_187,N_728);
or U893 (N_893,N_764,N_534);
nor U894 (N_894,N_594,N_776);
xor U895 (N_895,N_722,N_77);
xnor U896 (N_896,N_718,N_732);
nor U897 (N_897,N_734,N_757);
and U898 (N_898,N_778,N_715);
nand U899 (N_899,N_680,In_544);
and U900 (N_900,N_813,N_820);
and U901 (N_901,N_808,N_884);
xor U902 (N_902,N_860,N_878);
xnor U903 (N_903,N_836,N_814);
nor U904 (N_904,N_811,N_859);
or U905 (N_905,N_810,N_869);
and U906 (N_906,N_863,N_853);
or U907 (N_907,N_838,N_822);
or U908 (N_908,N_833,N_812);
nand U909 (N_909,N_800,N_877);
and U910 (N_910,N_850,N_827);
and U911 (N_911,N_807,N_840);
or U912 (N_912,N_809,N_893);
nor U913 (N_913,N_896,N_886);
and U914 (N_914,N_872,N_881);
or U915 (N_915,N_824,N_876);
nand U916 (N_916,N_879,N_894);
and U917 (N_917,N_899,N_837);
and U918 (N_918,N_830,N_817);
or U919 (N_919,N_870,N_871);
or U920 (N_920,N_851,N_803);
xor U921 (N_921,N_848,N_801);
xnor U922 (N_922,N_834,N_888);
nor U923 (N_923,N_867,N_825);
nor U924 (N_924,N_897,N_887);
nor U925 (N_925,N_818,N_885);
xor U926 (N_926,N_821,N_866);
or U927 (N_927,N_828,N_804);
xor U928 (N_928,N_856,N_835);
nor U929 (N_929,N_849,N_890);
nor U930 (N_930,N_823,N_880);
nor U931 (N_931,N_854,N_805);
nand U932 (N_932,N_815,N_868);
and U933 (N_933,N_839,N_826);
nand U934 (N_934,N_819,N_891);
xnor U935 (N_935,N_846,N_874);
nor U936 (N_936,N_895,N_841);
xnor U937 (N_937,N_882,N_829);
nor U938 (N_938,N_844,N_875);
xnor U939 (N_939,N_843,N_816);
nor U940 (N_940,N_857,N_847);
nor U941 (N_941,N_865,N_831);
nand U942 (N_942,N_845,N_862);
xor U943 (N_943,N_855,N_802);
nor U944 (N_944,N_852,N_889);
nand U945 (N_945,N_873,N_892);
and U946 (N_946,N_806,N_898);
xnor U947 (N_947,N_832,N_842);
nor U948 (N_948,N_861,N_864);
nor U949 (N_949,N_858,N_883);
xnor U950 (N_950,N_873,N_872);
nor U951 (N_951,N_840,N_813);
and U952 (N_952,N_867,N_801);
nand U953 (N_953,N_861,N_834);
nand U954 (N_954,N_854,N_837);
or U955 (N_955,N_851,N_895);
or U956 (N_956,N_829,N_822);
or U957 (N_957,N_857,N_898);
nand U958 (N_958,N_833,N_857);
and U959 (N_959,N_836,N_835);
nand U960 (N_960,N_821,N_889);
xor U961 (N_961,N_818,N_894);
nand U962 (N_962,N_847,N_803);
xor U963 (N_963,N_874,N_870);
or U964 (N_964,N_838,N_817);
nor U965 (N_965,N_870,N_847);
nand U966 (N_966,N_869,N_845);
and U967 (N_967,N_880,N_844);
nor U968 (N_968,N_856,N_861);
nand U969 (N_969,N_887,N_821);
or U970 (N_970,N_831,N_836);
and U971 (N_971,N_847,N_886);
and U972 (N_972,N_859,N_830);
nor U973 (N_973,N_834,N_877);
xnor U974 (N_974,N_863,N_835);
xor U975 (N_975,N_827,N_896);
nor U976 (N_976,N_817,N_842);
nand U977 (N_977,N_806,N_899);
nor U978 (N_978,N_882,N_822);
and U979 (N_979,N_879,N_848);
nor U980 (N_980,N_815,N_891);
xor U981 (N_981,N_889,N_809);
nand U982 (N_982,N_831,N_804);
xor U983 (N_983,N_857,N_854);
or U984 (N_984,N_802,N_848);
nand U985 (N_985,N_801,N_819);
nor U986 (N_986,N_829,N_808);
nand U987 (N_987,N_825,N_863);
nor U988 (N_988,N_868,N_888);
or U989 (N_989,N_830,N_826);
and U990 (N_990,N_825,N_850);
and U991 (N_991,N_863,N_852);
or U992 (N_992,N_899,N_844);
nor U993 (N_993,N_809,N_835);
or U994 (N_994,N_856,N_874);
and U995 (N_995,N_841,N_830);
and U996 (N_996,N_892,N_853);
xor U997 (N_997,N_882,N_849);
nor U998 (N_998,N_843,N_857);
nor U999 (N_999,N_888,N_882);
nand U1000 (N_1000,N_967,N_924);
nor U1001 (N_1001,N_903,N_987);
nor U1002 (N_1002,N_901,N_949);
nand U1003 (N_1003,N_907,N_966);
and U1004 (N_1004,N_995,N_928);
nand U1005 (N_1005,N_997,N_908);
xnor U1006 (N_1006,N_969,N_964);
nand U1007 (N_1007,N_976,N_951);
xnor U1008 (N_1008,N_915,N_905);
xor U1009 (N_1009,N_963,N_994);
xor U1010 (N_1010,N_921,N_932);
and U1011 (N_1011,N_927,N_941);
xnor U1012 (N_1012,N_902,N_913);
nor U1013 (N_1013,N_916,N_996);
xnor U1014 (N_1014,N_931,N_947);
or U1015 (N_1015,N_971,N_978);
or U1016 (N_1016,N_930,N_923);
nand U1017 (N_1017,N_943,N_939);
nand U1018 (N_1018,N_982,N_988);
nand U1019 (N_1019,N_925,N_942);
nor U1020 (N_1020,N_983,N_936);
or U1021 (N_1021,N_922,N_904);
nand U1022 (N_1022,N_998,N_985);
nor U1023 (N_1023,N_911,N_962);
nand U1024 (N_1024,N_929,N_933);
and U1025 (N_1025,N_955,N_918);
and U1026 (N_1026,N_965,N_981);
nand U1027 (N_1027,N_993,N_990);
nand U1028 (N_1028,N_946,N_917);
xor U1029 (N_1029,N_991,N_992);
or U1030 (N_1030,N_906,N_919);
xnor U1031 (N_1031,N_956,N_961);
and U1032 (N_1032,N_975,N_968);
nand U1033 (N_1033,N_953,N_958);
nand U1034 (N_1034,N_957,N_954);
nor U1035 (N_1035,N_986,N_940);
or U1036 (N_1036,N_979,N_999);
nor U1037 (N_1037,N_910,N_900);
nand U1038 (N_1038,N_959,N_950);
or U1039 (N_1039,N_945,N_974);
nand U1040 (N_1040,N_989,N_973);
or U1041 (N_1041,N_934,N_972);
nand U1042 (N_1042,N_914,N_970);
nand U1043 (N_1043,N_984,N_920);
nor U1044 (N_1044,N_935,N_912);
nor U1045 (N_1045,N_938,N_926);
or U1046 (N_1046,N_977,N_944);
xnor U1047 (N_1047,N_952,N_960);
xor U1048 (N_1048,N_980,N_909);
nor U1049 (N_1049,N_948,N_937);
nor U1050 (N_1050,N_987,N_941);
nor U1051 (N_1051,N_908,N_959);
or U1052 (N_1052,N_990,N_936);
or U1053 (N_1053,N_939,N_956);
nor U1054 (N_1054,N_938,N_957);
or U1055 (N_1055,N_950,N_945);
nand U1056 (N_1056,N_943,N_926);
or U1057 (N_1057,N_984,N_947);
xnor U1058 (N_1058,N_904,N_999);
nand U1059 (N_1059,N_989,N_947);
nor U1060 (N_1060,N_939,N_969);
or U1061 (N_1061,N_916,N_933);
and U1062 (N_1062,N_993,N_902);
nand U1063 (N_1063,N_949,N_966);
or U1064 (N_1064,N_901,N_938);
and U1065 (N_1065,N_941,N_978);
or U1066 (N_1066,N_924,N_989);
nor U1067 (N_1067,N_975,N_997);
nor U1068 (N_1068,N_975,N_915);
or U1069 (N_1069,N_974,N_932);
xnor U1070 (N_1070,N_910,N_984);
or U1071 (N_1071,N_965,N_932);
or U1072 (N_1072,N_980,N_964);
nor U1073 (N_1073,N_991,N_961);
xnor U1074 (N_1074,N_962,N_909);
nand U1075 (N_1075,N_955,N_906);
and U1076 (N_1076,N_946,N_936);
xor U1077 (N_1077,N_956,N_950);
nor U1078 (N_1078,N_925,N_998);
and U1079 (N_1079,N_998,N_965);
nand U1080 (N_1080,N_962,N_989);
xnor U1081 (N_1081,N_941,N_968);
and U1082 (N_1082,N_982,N_927);
nor U1083 (N_1083,N_944,N_935);
or U1084 (N_1084,N_940,N_916);
and U1085 (N_1085,N_957,N_921);
nor U1086 (N_1086,N_923,N_910);
and U1087 (N_1087,N_956,N_942);
nand U1088 (N_1088,N_981,N_904);
nand U1089 (N_1089,N_981,N_941);
nor U1090 (N_1090,N_956,N_904);
and U1091 (N_1091,N_999,N_933);
xnor U1092 (N_1092,N_921,N_905);
nor U1093 (N_1093,N_919,N_982);
nor U1094 (N_1094,N_935,N_900);
and U1095 (N_1095,N_937,N_965);
or U1096 (N_1096,N_958,N_920);
and U1097 (N_1097,N_903,N_907);
nand U1098 (N_1098,N_969,N_986);
nor U1099 (N_1099,N_934,N_994);
xnor U1100 (N_1100,N_1087,N_1089);
nand U1101 (N_1101,N_1048,N_1021);
or U1102 (N_1102,N_1033,N_1063);
xor U1103 (N_1103,N_1081,N_1078);
and U1104 (N_1104,N_1016,N_1009);
nand U1105 (N_1105,N_1075,N_1042);
and U1106 (N_1106,N_1030,N_1080);
nor U1107 (N_1107,N_1055,N_1057);
and U1108 (N_1108,N_1004,N_1059);
xor U1109 (N_1109,N_1071,N_1066);
nand U1110 (N_1110,N_1088,N_1037);
and U1111 (N_1111,N_1031,N_1090);
nor U1112 (N_1112,N_1005,N_1067);
nor U1113 (N_1113,N_1079,N_1069);
nor U1114 (N_1114,N_1058,N_1060);
and U1115 (N_1115,N_1093,N_1094);
nor U1116 (N_1116,N_1010,N_1034);
or U1117 (N_1117,N_1015,N_1032);
nor U1118 (N_1118,N_1013,N_1036);
nor U1119 (N_1119,N_1001,N_1050);
xor U1120 (N_1120,N_1028,N_1053);
nand U1121 (N_1121,N_1065,N_1092);
and U1122 (N_1122,N_1014,N_1018);
or U1123 (N_1123,N_1012,N_1040);
nor U1124 (N_1124,N_1061,N_1006);
nand U1125 (N_1125,N_1046,N_1022);
and U1126 (N_1126,N_1085,N_1025);
or U1127 (N_1127,N_1017,N_1064);
or U1128 (N_1128,N_1097,N_1086);
and U1129 (N_1129,N_1076,N_1073);
nand U1130 (N_1130,N_1082,N_1047);
or U1131 (N_1131,N_1074,N_1000);
or U1132 (N_1132,N_1054,N_1020);
or U1133 (N_1133,N_1024,N_1099);
xor U1134 (N_1134,N_1083,N_1056);
xnor U1135 (N_1135,N_1098,N_1039);
nand U1136 (N_1136,N_1027,N_1041);
or U1137 (N_1137,N_1019,N_1051);
and U1138 (N_1138,N_1095,N_1003);
xor U1139 (N_1139,N_1026,N_1096);
nand U1140 (N_1140,N_1044,N_1043);
or U1141 (N_1141,N_1038,N_1002);
xnor U1142 (N_1142,N_1052,N_1062);
nand U1143 (N_1143,N_1070,N_1029);
nor U1144 (N_1144,N_1011,N_1072);
nor U1145 (N_1145,N_1049,N_1035);
xnor U1146 (N_1146,N_1084,N_1023);
nor U1147 (N_1147,N_1007,N_1077);
or U1148 (N_1148,N_1045,N_1068);
and U1149 (N_1149,N_1008,N_1091);
xnor U1150 (N_1150,N_1088,N_1053);
xor U1151 (N_1151,N_1042,N_1067);
and U1152 (N_1152,N_1050,N_1037);
or U1153 (N_1153,N_1049,N_1071);
nand U1154 (N_1154,N_1079,N_1053);
nor U1155 (N_1155,N_1073,N_1011);
nor U1156 (N_1156,N_1005,N_1018);
nor U1157 (N_1157,N_1089,N_1060);
and U1158 (N_1158,N_1002,N_1007);
nand U1159 (N_1159,N_1079,N_1046);
xor U1160 (N_1160,N_1072,N_1045);
xor U1161 (N_1161,N_1030,N_1089);
nor U1162 (N_1162,N_1099,N_1020);
xnor U1163 (N_1163,N_1084,N_1087);
or U1164 (N_1164,N_1098,N_1043);
nor U1165 (N_1165,N_1085,N_1093);
or U1166 (N_1166,N_1020,N_1009);
nor U1167 (N_1167,N_1083,N_1015);
nand U1168 (N_1168,N_1062,N_1028);
nand U1169 (N_1169,N_1090,N_1067);
nor U1170 (N_1170,N_1050,N_1084);
and U1171 (N_1171,N_1026,N_1059);
or U1172 (N_1172,N_1036,N_1014);
nand U1173 (N_1173,N_1019,N_1038);
or U1174 (N_1174,N_1026,N_1069);
nor U1175 (N_1175,N_1045,N_1090);
nor U1176 (N_1176,N_1031,N_1024);
or U1177 (N_1177,N_1086,N_1055);
nor U1178 (N_1178,N_1087,N_1027);
and U1179 (N_1179,N_1014,N_1033);
xor U1180 (N_1180,N_1019,N_1026);
nor U1181 (N_1181,N_1060,N_1038);
xnor U1182 (N_1182,N_1056,N_1054);
xnor U1183 (N_1183,N_1013,N_1064);
nand U1184 (N_1184,N_1063,N_1056);
nor U1185 (N_1185,N_1056,N_1064);
nor U1186 (N_1186,N_1065,N_1019);
nor U1187 (N_1187,N_1068,N_1042);
xnor U1188 (N_1188,N_1083,N_1047);
nor U1189 (N_1189,N_1069,N_1062);
nor U1190 (N_1190,N_1021,N_1087);
and U1191 (N_1191,N_1051,N_1066);
and U1192 (N_1192,N_1029,N_1081);
nand U1193 (N_1193,N_1053,N_1032);
nor U1194 (N_1194,N_1095,N_1053);
xnor U1195 (N_1195,N_1029,N_1025);
nand U1196 (N_1196,N_1006,N_1092);
xnor U1197 (N_1197,N_1085,N_1038);
nor U1198 (N_1198,N_1041,N_1089);
xnor U1199 (N_1199,N_1093,N_1053);
nand U1200 (N_1200,N_1153,N_1189);
nor U1201 (N_1201,N_1190,N_1180);
or U1202 (N_1202,N_1127,N_1128);
or U1203 (N_1203,N_1177,N_1100);
xor U1204 (N_1204,N_1172,N_1152);
nor U1205 (N_1205,N_1121,N_1125);
nand U1206 (N_1206,N_1136,N_1111);
or U1207 (N_1207,N_1123,N_1129);
xnor U1208 (N_1208,N_1137,N_1175);
nand U1209 (N_1209,N_1120,N_1112);
xnor U1210 (N_1210,N_1101,N_1142);
nor U1211 (N_1211,N_1182,N_1109);
xor U1212 (N_1212,N_1124,N_1166);
xor U1213 (N_1213,N_1191,N_1154);
and U1214 (N_1214,N_1163,N_1132);
xnor U1215 (N_1215,N_1114,N_1176);
xnor U1216 (N_1216,N_1134,N_1181);
or U1217 (N_1217,N_1145,N_1179);
nor U1218 (N_1218,N_1118,N_1162);
nand U1219 (N_1219,N_1195,N_1161);
xnor U1220 (N_1220,N_1164,N_1196);
nand U1221 (N_1221,N_1108,N_1104);
xor U1222 (N_1222,N_1155,N_1116);
nand U1223 (N_1223,N_1115,N_1110);
nor U1224 (N_1224,N_1146,N_1188);
and U1225 (N_1225,N_1148,N_1119);
xnor U1226 (N_1226,N_1133,N_1107);
nor U1227 (N_1227,N_1158,N_1117);
xnor U1228 (N_1228,N_1149,N_1159);
or U1229 (N_1229,N_1169,N_1168);
and U1230 (N_1230,N_1199,N_1106);
or U1231 (N_1231,N_1102,N_1138);
nor U1232 (N_1232,N_1173,N_1140);
or U1233 (N_1233,N_1193,N_1144);
xor U1234 (N_1234,N_1197,N_1147);
xnor U1235 (N_1235,N_1151,N_1183);
nor U1236 (N_1236,N_1174,N_1103);
and U1237 (N_1237,N_1170,N_1192);
and U1238 (N_1238,N_1105,N_1198);
nor U1239 (N_1239,N_1122,N_1184);
and U1240 (N_1240,N_1130,N_1157);
xor U1241 (N_1241,N_1194,N_1135);
or U1242 (N_1242,N_1171,N_1167);
xnor U1243 (N_1243,N_1131,N_1185);
xor U1244 (N_1244,N_1187,N_1178);
nand U1245 (N_1245,N_1160,N_1186);
or U1246 (N_1246,N_1113,N_1143);
xor U1247 (N_1247,N_1150,N_1165);
nand U1248 (N_1248,N_1156,N_1139);
nand U1249 (N_1249,N_1141,N_1126);
nand U1250 (N_1250,N_1145,N_1108);
and U1251 (N_1251,N_1177,N_1134);
xnor U1252 (N_1252,N_1199,N_1138);
and U1253 (N_1253,N_1170,N_1135);
nand U1254 (N_1254,N_1150,N_1132);
or U1255 (N_1255,N_1132,N_1111);
or U1256 (N_1256,N_1192,N_1128);
or U1257 (N_1257,N_1194,N_1177);
and U1258 (N_1258,N_1131,N_1194);
xnor U1259 (N_1259,N_1164,N_1145);
and U1260 (N_1260,N_1121,N_1160);
xnor U1261 (N_1261,N_1128,N_1190);
nor U1262 (N_1262,N_1115,N_1137);
nand U1263 (N_1263,N_1193,N_1194);
and U1264 (N_1264,N_1198,N_1197);
and U1265 (N_1265,N_1145,N_1191);
or U1266 (N_1266,N_1193,N_1166);
nor U1267 (N_1267,N_1147,N_1172);
and U1268 (N_1268,N_1136,N_1127);
nor U1269 (N_1269,N_1186,N_1118);
xnor U1270 (N_1270,N_1121,N_1176);
nand U1271 (N_1271,N_1108,N_1147);
xnor U1272 (N_1272,N_1153,N_1121);
or U1273 (N_1273,N_1120,N_1181);
xor U1274 (N_1274,N_1195,N_1157);
nor U1275 (N_1275,N_1166,N_1189);
xor U1276 (N_1276,N_1138,N_1144);
or U1277 (N_1277,N_1161,N_1127);
xor U1278 (N_1278,N_1100,N_1191);
nor U1279 (N_1279,N_1169,N_1138);
xor U1280 (N_1280,N_1111,N_1160);
or U1281 (N_1281,N_1104,N_1183);
xor U1282 (N_1282,N_1140,N_1142);
and U1283 (N_1283,N_1161,N_1176);
xor U1284 (N_1284,N_1115,N_1147);
and U1285 (N_1285,N_1159,N_1183);
and U1286 (N_1286,N_1122,N_1188);
xnor U1287 (N_1287,N_1172,N_1117);
and U1288 (N_1288,N_1118,N_1190);
and U1289 (N_1289,N_1126,N_1124);
and U1290 (N_1290,N_1132,N_1159);
and U1291 (N_1291,N_1136,N_1181);
nand U1292 (N_1292,N_1159,N_1143);
and U1293 (N_1293,N_1144,N_1184);
and U1294 (N_1294,N_1170,N_1173);
nand U1295 (N_1295,N_1109,N_1157);
and U1296 (N_1296,N_1194,N_1132);
nand U1297 (N_1297,N_1135,N_1188);
or U1298 (N_1298,N_1175,N_1133);
nor U1299 (N_1299,N_1170,N_1140);
xnor U1300 (N_1300,N_1285,N_1262);
and U1301 (N_1301,N_1216,N_1267);
or U1302 (N_1302,N_1228,N_1207);
xnor U1303 (N_1303,N_1258,N_1241);
nand U1304 (N_1304,N_1223,N_1266);
nor U1305 (N_1305,N_1231,N_1261);
xor U1306 (N_1306,N_1201,N_1248);
nand U1307 (N_1307,N_1209,N_1239);
xor U1308 (N_1308,N_1210,N_1233);
or U1309 (N_1309,N_1269,N_1242);
and U1310 (N_1310,N_1294,N_1288);
xor U1311 (N_1311,N_1205,N_1278);
and U1312 (N_1312,N_1275,N_1283);
or U1313 (N_1313,N_1222,N_1206);
or U1314 (N_1314,N_1227,N_1244);
or U1315 (N_1315,N_1263,N_1286);
and U1316 (N_1316,N_1290,N_1282);
xor U1317 (N_1317,N_1254,N_1219);
and U1318 (N_1318,N_1264,N_1289);
or U1319 (N_1319,N_1214,N_1215);
and U1320 (N_1320,N_1213,N_1225);
nor U1321 (N_1321,N_1211,N_1240);
nor U1322 (N_1322,N_1238,N_1260);
nor U1323 (N_1323,N_1272,N_1247);
and U1324 (N_1324,N_1251,N_1243);
and U1325 (N_1325,N_1292,N_1252);
and U1326 (N_1326,N_1202,N_1268);
nand U1327 (N_1327,N_1277,N_1281);
and U1328 (N_1328,N_1291,N_1250);
or U1329 (N_1329,N_1274,N_1212);
and U1330 (N_1330,N_1203,N_1229);
nor U1331 (N_1331,N_1280,N_1232);
and U1332 (N_1332,N_1217,N_1235);
and U1333 (N_1333,N_1246,N_1220);
and U1334 (N_1334,N_1204,N_1256);
xor U1335 (N_1335,N_1236,N_1293);
and U1336 (N_1336,N_1253,N_1299);
and U1337 (N_1337,N_1279,N_1287);
and U1338 (N_1338,N_1249,N_1230);
or U1339 (N_1339,N_1273,N_1234);
or U1340 (N_1340,N_1270,N_1298);
and U1341 (N_1341,N_1200,N_1284);
or U1342 (N_1342,N_1276,N_1208);
and U1343 (N_1343,N_1226,N_1296);
and U1344 (N_1344,N_1271,N_1218);
nor U1345 (N_1345,N_1224,N_1255);
nand U1346 (N_1346,N_1245,N_1221);
nor U1347 (N_1347,N_1259,N_1265);
and U1348 (N_1348,N_1295,N_1237);
xnor U1349 (N_1349,N_1257,N_1297);
xor U1350 (N_1350,N_1244,N_1247);
and U1351 (N_1351,N_1267,N_1293);
nor U1352 (N_1352,N_1253,N_1251);
or U1353 (N_1353,N_1220,N_1206);
xnor U1354 (N_1354,N_1231,N_1247);
nor U1355 (N_1355,N_1212,N_1209);
xor U1356 (N_1356,N_1205,N_1201);
nand U1357 (N_1357,N_1229,N_1200);
nor U1358 (N_1358,N_1226,N_1267);
and U1359 (N_1359,N_1294,N_1297);
xor U1360 (N_1360,N_1299,N_1248);
and U1361 (N_1361,N_1236,N_1213);
or U1362 (N_1362,N_1266,N_1298);
nand U1363 (N_1363,N_1207,N_1247);
nand U1364 (N_1364,N_1201,N_1254);
nor U1365 (N_1365,N_1275,N_1297);
and U1366 (N_1366,N_1232,N_1293);
nor U1367 (N_1367,N_1258,N_1278);
nand U1368 (N_1368,N_1231,N_1258);
and U1369 (N_1369,N_1233,N_1207);
nand U1370 (N_1370,N_1208,N_1293);
and U1371 (N_1371,N_1229,N_1208);
or U1372 (N_1372,N_1222,N_1251);
nand U1373 (N_1373,N_1267,N_1201);
xnor U1374 (N_1374,N_1204,N_1298);
and U1375 (N_1375,N_1294,N_1235);
and U1376 (N_1376,N_1263,N_1290);
nor U1377 (N_1377,N_1242,N_1212);
and U1378 (N_1378,N_1205,N_1268);
and U1379 (N_1379,N_1244,N_1201);
nand U1380 (N_1380,N_1292,N_1269);
xor U1381 (N_1381,N_1236,N_1215);
nand U1382 (N_1382,N_1226,N_1284);
xnor U1383 (N_1383,N_1221,N_1222);
and U1384 (N_1384,N_1231,N_1234);
and U1385 (N_1385,N_1205,N_1272);
and U1386 (N_1386,N_1267,N_1274);
and U1387 (N_1387,N_1265,N_1274);
and U1388 (N_1388,N_1276,N_1269);
or U1389 (N_1389,N_1267,N_1206);
nor U1390 (N_1390,N_1290,N_1245);
or U1391 (N_1391,N_1232,N_1223);
nand U1392 (N_1392,N_1271,N_1253);
or U1393 (N_1393,N_1248,N_1293);
or U1394 (N_1394,N_1233,N_1216);
and U1395 (N_1395,N_1211,N_1260);
nand U1396 (N_1396,N_1289,N_1234);
xor U1397 (N_1397,N_1217,N_1295);
nand U1398 (N_1398,N_1251,N_1204);
or U1399 (N_1399,N_1296,N_1217);
or U1400 (N_1400,N_1314,N_1331);
or U1401 (N_1401,N_1340,N_1303);
nand U1402 (N_1402,N_1347,N_1359);
nand U1403 (N_1403,N_1352,N_1392);
nor U1404 (N_1404,N_1355,N_1354);
xnor U1405 (N_1405,N_1356,N_1316);
or U1406 (N_1406,N_1350,N_1388);
or U1407 (N_1407,N_1386,N_1368);
or U1408 (N_1408,N_1332,N_1345);
xor U1409 (N_1409,N_1397,N_1323);
nor U1410 (N_1410,N_1394,N_1334);
nor U1411 (N_1411,N_1390,N_1312);
nor U1412 (N_1412,N_1377,N_1361);
xor U1413 (N_1413,N_1358,N_1339);
and U1414 (N_1414,N_1343,N_1319);
and U1415 (N_1415,N_1328,N_1341);
or U1416 (N_1416,N_1369,N_1310);
or U1417 (N_1417,N_1395,N_1373);
xnor U1418 (N_1418,N_1384,N_1364);
xnor U1419 (N_1419,N_1333,N_1387);
or U1420 (N_1420,N_1348,N_1320);
and U1421 (N_1421,N_1338,N_1376);
or U1422 (N_1422,N_1324,N_1362);
or U1423 (N_1423,N_1302,N_1365);
nand U1424 (N_1424,N_1380,N_1383);
and U1425 (N_1425,N_1379,N_1344);
and U1426 (N_1426,N_1389,N_1307);
or U1427 (N_1427,N_1304,N_1318);
or U1428 (N_1428,N_1301,N_1335);
and U1429 (N_1429,N_1330,N_1393);
and U1430 (N_1430,N_1375,N_1357);
nor U1431 (N_1431,N_1315,N_1326);
or U1432 (N_1432,N_1329,N_1370);
and U1433 (N_1433,N_1367,N_1336);
or U1434 (N_1434,N_1325,N_1399);
or U1435 (N_1435,N_1363,N_1391);
or U1436 (N_1436,N_1308,N_1360);
nor U1437 (N_1437,N_1311,N_1374);
nand U1438 (N_1438,N_1305,N_1322);
nor U1439 (N_1439,N_1382,N_1371);
xor U1440 (N_1440,N_1366,N_1321);
nor U1441 (N_1441,N_1396,N_1385);
xnor U1442 (N_1442,N_1317,N_1378);
or U1443 (N_1443,N_1309,N_1327);
or U1444 (N_1444,N_1398,N_1349);
nand U1445 (N_1445,N_1300,N_1346);
nor U1446 (N_1446,N_1342,N_1381);
nand U1447 (N_1447,N_1306,N_1353);
xor U1448 (N_1448,N_1351,N_1372);
and U1449 (N_1449,N_1313,N_1337);
nor U1450 (N_1450,N_1332,N_1309);
or U1451 (N_1451,N_1339,N_1338);
or U1452 (N_1452,N_1385,N_1303);
xor U1453 (N_1453,N_1322,N_1373);
nand U1454 (N_1454,N_1380,N_1330);
nor U1455 (N_1455,N_1351,N_1349);
or U1456 (N_1456,N_1330,N_1386);
xor U1457 (N_1457,N_1332,N_1337);
or U1458 (N_1458,N_1321,N_1338);
nor U1459 (N_1459,N_1321,N_1311);
nand U1460 (N_1460,N_1382,N_1370);
or U1461 (N_1461,N_1353,N_1379);
nor U1462 (N_1462,N_1374,N_1347);
nand U1463 (N_1463,N_1345,N_1341);
or U1464 (N_1464,N_1377,N_1394);
nand U1465 (N_1465,N_1369,N_1360);
nor U1466 (N_1466,N_1336,N_1362);
nor U1467 (N_1467,N_1309,N_1319);
xnor U1468 (N_1468,N_1335,N_1353);
nand U1469 (N_1469,N_1340,N_1389);
or U1470 (N_1470,N_1358,N_1376);
xnor U1471 (N_1471,N_1370,N_1368);
nor U1472 (N_1472,N_1363,N_1386);
or U1473 (N_1473,N_1310,N_1341);
and U1474 (N_1474,N_1316,N_1307);
or U1475 (N_1475,N_1352,N_1310);
and U1476 (N_1476,N_1307,N_1321);
nor U1477 (N_1477,N_1319,N_1356);
xnor U1478 (N_1478,N_1380,N_1311);
and U1479 (N_1479,N_1398,N_1381);
xnor U1480 (N_1480,N_1318,N_1391);
nand U1481 (N_1481,N_1379,N_1376);
nor U1482 (N_1482,N_1373,N_1384);
xor U1483 (N_1483,N_1393,N_1397);
and U1484 (N_1484,N_1390,N_1323);
xor U1485 (N_1485,N_1397,N_1315);
nand U1486 (N_1486,N_1388,N_1387);
nor U1487 (N_1487,N_1352,N_1341);
nand U1488 (N_1488,N_1397,N_1339);
and U1489 (N_1489,N_1318,N_1374);
and U1490 (N_1490,N_1357,N_1314);
and U1491 (N_1491,N_1383,N_1356);
nor U1492 (N_1492,N_1369,N_1341);
or U1493 (N_1493,N_1389,N_1383);
xnor U1494 (N_1494,N_1363,N_1308);
nand U1495 (N_1495,N_1369,N_1361);
nor U1496 (N_1496,N_1389,N_1374);
and U1497 (N_1497,N_1347,N_1340);
nor U1498 (N_1498,N_1329,N_1346);
nor U1499 (N_1499,N_1356,N_1371);
or U1500 (N_1500,N_1495,N_1493);
xor U1501 (N_1501,N_1436,N_1474);
nor U1502 (N_1502,N_1434,N_1472);
nor U1503 (N_1503,N_1433,N_1448);
xnor U1504 (N_1504,N_1485,N_1446);
and U1505 (N_1505,N_1449,N_1425);
and U1506 (N_1506,N_1424,N_1460);
or U1507 (N_1507,N_1488,N_1465);
nor U1508 (N_1508,N_1471,N_1439);
nor U1509 (N_1509,N_1458,N_1438);
nor U1510 (N_1510,N_1475,N_1435);
or U1511 (N_1511,N_1453,N_1479);
or U1512 (N_1512,N_1402,N_1430);
and U1513 (N_1513,N_1432,N_1492);
nor U1514 (N_1514,N_1447,N_1410);
nand U1515 (N_1515,N_1409,N_1423);
and U1516 (N_1516,N_1412,N_1497);
nor U1517 (N_1517,N_1482,N_1431);
nor U1518 (N_1518,N_1417,N_1400);
xor U1519 (N_1519,N_1477,N_1455);
nand U1520 (N_1520,N_1422,N_1469);
and U1521 (N_1521,N_1442,N_1413);
or U1522 (N_1522,N_1428,N_1483);
nand U1523 (N_1523,N_1478,N_1407);
and U1524 (N_1524,N_1499,N_1440);
nand U1525 (N_1525,N_1451,N_1418);
xor U1526 (N_1526,N_1420,N_1456);
xnor U1527 (N_1527,N_1498,N_1415);
or U1528 (N_1528,N_1411,N_1414);
nand U1529 (N_1529,N_1487,N_1450);
nor U1530 (N_1530,N_1404,N_1480);
or U1531 (N_1531,N_1427,N_1426);
or U1532 (N_1532,N_1496,N_1416);
and U1533 (N_1533,N_1486,N_1494);
xnor U1534 (N_1534,N_1462,N_1464);
and U1535 (N_1535,N_1470,N_1489);
or U1536 (N_1536,N_1437,N_1401);
nand U1537 (N_1537,N_1461,N_1452);
and U1538 (N_1538,N_1421,N_1491);
nand U1539 (N_1539,N_1443,N_1403);
and U1540 (N_1540,N_1445,N_1463);
or U1541 (N_1541,N_1444,N_1473);
nand U1542 (N_1542,N_1419,N_1459);
nor U1543 (N_1543,N_1468,N_1484);
xnor U1544 (N_1544,N_1481,N_1467);
nor U1545 (N_1545,N_1441,N_1429);
and U1546 (N_1546,N_1408,N_1490);
nor U1547 (N_1547,N_1406,N_1454);
nand U1548 (N_1548,N_1457,N_1466);
or U1549 (N_1549,N_1405,N_1476);
nor U1550 (N_1550,N_1456,N_1408);
or U1551 (N_1551,N_1470,N_1479);
and U1552 (N_1552,N_1423,N_1475);
and U1553 (N_1553,N_1448,N_1462);
or U1554 (N_1554,N_1470,N_1412);
xor U1555 (N_1555,N_1416,N_1495);
nor U1556 (N_1556,N_1476,N_1466);
xnor U1557 (N_1557,N_1425,N_1472);
nand U1558 (N_1558,N_1431,N_1440);
xor U1559 (N_1559,N_1458,N_1457);
and U1560 (N_1560,N_1438,N_1469);
or U1561 (N_1561,N_1475,N_1434);
nand U1562 (N_1562,N_1431,N_1494);
nand U1563 (N_1563,N_1432,N_1419);
and U1564 (N_1564,N_1455,N_1442);
and U1565 (N_1565,N_1473,N_1405);
nand U1566 (N_1566,N_1444,N_1489);
nor U1567 (N_1567,N_1495,N_1428);
or U1568 (N_1568,N_1487,N_1476);
xnor U1569 (N_1569,N_1448,N_1494);
and U1570 (N_1570,N_1402,N_1457);
nand U1571 (N_1571,N_1453,N_1424);
xor U1572 (N_1572,N_1440,N_1456);
xor U1573 (N_1573,N_1467,N_1415);
or U1574 (N_1574,N_1489,N_1483);
nor U1575 (N_1575,N_1454,N_1430);
or U1576 (N_1576,N_1498,N_1472);
or U1577 (N_1577,N_1409,N_1460);
and U1578 (N_1578,N_1441,N_1451);
xor U1579 (N_1579,N_1484,N_1427);
and U1580 (N_1580,N_1444,N_1487);
and U1581 (N_1581,N_1400,N_1422);
or U1582 (N_1582,N_1479,N_1463);
nor U1583 (N_1583,N_1434,N_1430);
nand U1584 (N_1584,N_1453,N_1499);
or U1585 (N_1585,N_1430,N_1447);
or U1586 (N_1586,N_1474,N_1400);
nor U1587 (N_1587,N_1421,N_1448);
xor U1588 (N_1588,N_1419,N_1467);
nor U1589 (N_1589,N_1465,N_1426);
xnor U1590 (N_1590,N_1403,N_1438);
nor U1591 (N_1591,N_1439,N_1402);
nand U1592 (N_1592,N_1449,N_1443);
nand U1593 (N_1593,N_1406,N_1443);
xnor U1594 (N_1594,N_1439,N_1436);
nor U1595 (N_1595,N_1402,N_1465);
nand U1596 (N_1596,N_1440,N_1409);
nor U1597 (N_1597,N_1428,N_1423);
nand U1598 (N_1598,N_1478,N_1499);
and U1599 (N_1599,N_1438,N_1408);
and U1600 (N_1600,N_1509,N_1539);
nand U1601 (N_1601,N_1511,N_1578);
xor U1602 (N_1602,N_1591,N_1589);
and U1603 (N_1603,N_1581,N_1556);
and U1604 (N_1604,N_1513,N_1512);
xor U1605 (N_1605,N_1579,N_1557);
nand U1606 (N_1606,N_1598,N_1558);
and U1607 (N_1607,N_1569,N_1590);
xor U1608 (N_1608,N_1523,N_1501);
xor U1609 (N_1609,N_1516,N_1528);
and U1610 (N_1610,N_1505,N_1500);
or U1611 (N_1611,N_1510,N_1531);
and U1612 (N_1612,N_1560,N_1596);
nor U1613 (N_1613,N_1588,N_1533);
or U1614 (N_1614,N_1585,N_1526);
or U1615 (N_1615,N_1535,N_1503);
or U1616 (N_1616,N_1519,N_1553);
xor U1617 (N_1617,N_1575,N_1555);
or U1618 (N_1618,N_1532,N_1524);
nor U1619 (N_1619,N_1541,N_1561);
nor U1620 (N_1620,N_1599,N_1582);
xnor U1621 (N_1621,N_1522,N_1568);
or U1622 (N_1622,N_1594,N_1530);
nor U1623 (N_1623,N_1551,N_1549);
or U1624 (N_1624,N_1564,N_1507);
xor U1625 (N_1625,N_1543,N_1550);
and U1626 (N_1626,N_1515,N_1518);
nor U1627 (N_1627,N_1559,N_1504);
xnor U1628 (N_1628,N_1597,N_1573);
and U1629 (N_1629,N_1517,N_1565);
or U1630 (N_1630,N_1546,N_1593);
or U1631 (N_1631,N_1587,N_1548);
nor U1632 (N_1632,N_1563,N_1580);
or U1633 (N_1633,N_1572,N_1502);
and U1634 (N_1634,N_1538,N_1592);
or U1635 (N_1635,N_1547,N_1521);
or U1636 (N_1636,N_1567,N_1554);
xnor U1637 (N_1637,N_1562,N_1586);
nor U1638 (N_1638,N_1583,N_1506);
xnor U1639 (N_1639,N_1536,N_1527);
nor U1640 (N_1640,N_1542,N_1537);
and U1641 (N_1641,N_1545,N_1508);
nand U1642 (N_1642,N_1577,N_1520);
or U1643 (N_1643,N_1571,N_1552);
and U1644 (N_1644,N_1529,N_1570);
or U1645 (N_1645,N_1584,N_1514);
nand U1646 (N_1646,N_1595,N_1566);
and U1647 (N_1647,N_1576,N_1544);
and U1648 (N_1648,N_1525,N_1574);
xnor U1649 (N_1649,N_1540,N_1534);
xnor U1650 (N_1650,N_1585,N_1591);
xnor U1651 (N_1651,N_1590,N_1585);
xor U1652 (N_1652,N_1520,N_1521);
nor U1653 (N_1653,N_1556,N_1594);
and U1654 (N_1654,N_1520,N_1569);
or U1655 (N_1655,N_1543,N_1506);
or U1656 (N_1656,N_1573,N_1535);
nor U1657 (N_1657,N_1596,N_1583);
nand U1658 (N_1658,N_1561,N_1538);
nor U1659 (N_1659,N_1532,N_1536);
nand U1660 (N_1660,N_1510,N_1574);
and U1661 (N_1661,N_1560,N_1575);
xnor U1662 (N_1662,N_1548,N_1520);
and U1663 (N_1663,N_1517,N_1590);
or U1664 (N_1664,N_1538,N_1531);
nand U1665 (N_1665,N_1554,N_1536);
nor U1666 (N_1666,N_1527,N_1596);
or U1667 (N_1667,N_1579,N_1575);
and U1668 (N_1668,N_1527,N_1541);
nand U1669 (N_1669,N_1579,N_1564);
and U1670 (N_1670,N_1501,N_1500);
nor U1671 (N_1671,N_1518,N_1531);
nor U1672 (N_1672,N_1598,N_1547);
xor U1673 (N_1673,N_1566,N_1547);
nand U1674 (N_1674,N_1575,N_1532);
nor U1675 (N_1675,N_1515,N_1505);
or U1676 (N_1676,N_1526,N_1547);
or U1677 (N_1677,N_1533,N_1578);
or U1678 (N_1678,N_1596,N_1594);
nand U1679 (N_1679,N_1556,N_1507);
nand U1680 (N_1680,N_1589,N_1599);
nor U1681 (N_1681,N_1583,N_1537);
and U1682 (N_1682,N_1570,N_1598);
and U1683 (N_1683,N_1524,N_1507);
and U1684 (N_1684,N_1558,N_1559);
xor U1685 (N_1685,N_1518,N_1551);
xnor U1686 (N_1686,N_1541,N_1519);
or U1687 (N_1687,N_1523,N_1579);
nand U1688 (N_1688,N_1573,N_1569);
and U1689 (N_1689,N_1549,N_1578);
xor U1690 (N_1690,N_1589,N_1545);
or U1691 (N_1691,N_1528,N_1558);
xor U1692 (N_1692,N_1594,N_1515);
and U1693 (N_1693,N_1506,N_1589);
xnor U1694 (N_1694,N_1527,N_1592);
nand U1695 (N_1695,N_1551,N_1564);
or U1696 (N_1696,N_1536,N_1512);
nand U1697 (N_1697,N_1587,N_1509);
nand U1698 (N_1698,N_1548,N_1577);
and U1699 (N_1699,N_1507,N_1503);
xor U1700 (N_1700,N_1605,N_1668);
or U1701 (N_1701,N_1629,N_1674);
xor U1702 (N_1702,N_1687,N_1660);
nand U1703 (N_1703,N_1625,N_1665);
or U1704 (N_1704,N_1698,N_1686);
nand U1705 (N_1705,N_1615,N_1692);
nor U1706 (N_1706,N_1690,N_1663);
or U1707 (N_1707,N_1673,N_1627);
xor U1708 (N_1708,N_1643,N_1650);
or U1709 (N_1709,N_1677,N_1671);
nor U1710 (N_1710,N_1641,N_1658);
and U1711 (N_1711,N_1610,N_1657);
and U1712 (N_1712,N_1614,N_1685);
xnor U1713 (N_1713,N_1683,N_1634);
nor U1714 (N_1714,N_1631,N_1602);
or U1715 (N_1715,N_1682,N_1645);
nand U1716 (N_1716,N_1632,N_1633);
or U1717 (N_1717,N_1681,N_1616);
and U1718 (N_1718,N_1662,N_1624);
nand U1719 (N_1719,N_1679,N_1654);
nand U1720 (N_1720,N_1612,N_1667);
and U1721 (N_1721,N_1638,N_1604);
nor U1722 (N_1722,N_1618,N_1619);
nor U1723 (N_1723,N_1656,N_1695);
nand U1724 (N_1724,N_1623,N_1607);
and U1725 (N_1725,N_1651,N_1684);
xnor U1726 (N_1726,N_1649,N_1637);
xor U1727 (N_1727,N_1608,N_1600);
or U1728 (N_1728,N_1606,N_1689);
or U1729 (N_1729,N_1669,N_1630);
xnor U1730 (N_1730,N_1642,N_1680);
nand U1731 (N_1731,N_1697,N_1659);
nand U1732 (N_1732,N_1628,N_1603);
or U1733 (N_1733,N_1644,N_1611);
and U1734 (N_1734,N_1676,N_1613);
and U1735 (N_1735,N_1694,N_1647);
xor U1736 (N_1736,N_1666,N_1672);
xor U1737 (N_1737,N_1621,N_1675);
xnor U1738 (N_1738,N_1640,N_1696);
or U1739 (N_1739,N_1653,N_1617);
xnor U1740 (N_1740,N_1646,N_1693);
nand U1741 (N_1741,N_1652,N_1636);
and U1742 (N_1742,N_1670,N_1626);
nor U1743 (N_1743,N_1691,N_1664);
or U1744 (N_1744,N_1688,N_1678);
nor U1745 (N_1745,N_1609,N_1648);
nand U1746 (N_1746,N_1661,N_1699);
nor U1747 (N_1747,N_1601,N_1639);
nor U1748 (N_1748,N_1655,N_1622);
nand U1749 (N_1749,N_1635,N_1620);
xor U1750 (N_1750,N_1691,N_1653);
and U1751 (N_1751,N_1612,N_1694);
and U1752 (N_1752,N_1619,N_1676);
and U1753 (N_1753,N_1610,N_1663);
or U1754 (N_1754,N_1666,N_1643);
xor U1755 (N_1755,N_1657,N_1644);
nand U1756 (N_1756,N_1699,N_1672);
and U1757 (N_1757,N_1679,N_1615);
nand U1758 (N_1758,N_1690,N_1639);
and U1759 (N_1759,N_1600,N_1605);
nor U1760 (N_1760,N_1669,N_1628);
or U1761 (N_1761,N_1682,N_1603);
nor U1762 (N_1762,N_1629,N_1647);
nand U1763 (N_1763,N_1697,N_1694);
xnor U1764 (N_1764,N_1613,N_1648);
and U1765 (N_1765,N_1624,N_1677);
xor U1766 (N_1766,N_1656,N_1637);
xnor U1767 (N_1767,N_1645,N_1621);
nor U1768 (N_1768,N_1600,N_1685);
nor U1769 (N_1769,N_1660,N_1631);
or U1770 (N_1770,N_1643,N_1628);
nor U1771 (N_1771,N_1607,N_1690);
nand U1772 (N_1772,N_1689,N_1671);
and U1773 (N_1773,N_1607,N_1684);
nand U1774 (N_1774,N_1697,N_1636);
and U1775 (N_1775,N_1637,N_1640);
nand U1776 (N_1776,N_1636,N_1625);
and U1777 (N_1777,N_1650,N_1606);
and U1778 (N_1778,N_1643,N_1645);
nand U1779 (N_1779,N_1605,N_1647);
and U1780 (N_1780,N_1610,N_1695);
or U1781 (N_1781,N_1669,N_1673);
nor U1782 (N_1782,N_1695,N_1691);
nor U1783 (N_1783,N_1609,N_1630);
xor U1784 (N_1784,N_1697,N_1661);
nor U1785 (N_1785,N_1603,N_1685);
nor U1786 (N_1786,N_1692,N_1611);
xor U1787 (N_1787,N_1652,N_1612);
nand U1788 (N_1788,N_1648,N_1649);
xor U1789 (N_1789,N_1651,N_1614);
or U1790 (N_1790,N_1697,N_1663);
xnor U1791 (N_1791,N_1601,N_1606);
and U1792 (N_1792,N_1686,N_1630);
or U1793 (N_1793,N_1646,N_1699);
xnor U1794 (N_1794,N_1613,N_1611);
and U1795 (N_1795,N_1646,N_1637);
nor U1796 (N_1796,N_1607,N_1620);
or U1797 (N_1797,N_1679,N_1678);
nand U1798 (N_1798,N_1602,N_1617);
nor U1799 (N_1799,N_1681,N_1609);
nand U1800 (N_1800,N_1789,N_1736);
nand U1801 (N_1801,N_1762,N_1727);
nand U1802 (N_1802,N_1764,N_1744);
nand U1803 (N_1803,N_1739,N_1714);
nor U1804 (N_1804,N_1784,N_1756);
nor U1805 (N_1805,N_1751,N_1705);
nand U1806 (N_1806,N_1750,N_1708);
xnor U1807 (N_1807,N_1746,N_1729);
and U1808 (N_1808,N_1740,N_1783);
nor U1809 (N_1809,N_1735,N_1755);
nand U1810 (N_1810,N_1753,N_1765);
nand U1811 (N_1811,N_1713,N_1730);
xor U1812 (N_1812,N_1781,N_1718);
xor U1813 (N_1813,N_1754,N_1707);
nor U1814 (N_1814,N_1741,N_1770);
and U1815 (N_1815,N_1706,N_1763);
nand U1816 (N_1816,N_1722,N_1771);
or U1817 (N_1817,N_1712,N_1704);
or U1818 (N_1818,N_1772,N_1752);
nor U1819 (N_1819,N_1738,N_1798);
nor U1820 (N_1820,N_1702,N_1709);
xnor U1821 (N_1821,N_1728,N_1716);
or U1822 (N_1822,N_1792,N_1748);
xnor U1823 (N_1823,N_1757,N_1745);
nand U1824 (N_1824,N_1780,N_1785);
and U1825 (N_1825,N_1796,N_1723);
or U1826 (N_1826,N_1720,N_1700);
nor U1827 (N_1827,N_1788,N_1777);
and U1828 (N_1828,N_1797,N_1724);
nor U1829 (N_1829,N_1759,N_1768);
or U1830 (N_1830,N_1761,N_1775);
nor U1831 (N_1831,N_1773,N_1779);
or U1832 (N_1832,N_1737,N_1711);
or U1833 (N_1833,N_1742,N_1710);
xnor U1834 (N_1834,N_1733,N_1717);
or U1835 (N_1835,N_1731,N_1743);
nor U1836 (N_1836,N_1769,N_1747);
nand U1837 (N_1837,N_1786,N_1795);
xnor U1838 (N_1838,N_1790,N_1787);
nor U1839 (N_1839,N_1719,N_1715);
or U1840 (N_1840,N_1760,N_1766);
nand U1841 (N_1841,N_1734,N_1758);
or U1842 (N_1842,N_1774,N_1799);
nor U1843 (N_1843,N_1725,N_1701);
or U1844 (N_1844,N_1778,N_1791);
and U1845 (N_1845,N_1721,N_1726);
nor U1846 (N_1846,N_1749,N_1793);
and U1847 (N_1847,N_1732,N_1794);
nor U1848 (N_1848,N_1703,N_1767);
or U1849 (N_1849,N_1776,N_1782);
nand U1850 (N_1850,N_1726,N_1707);
xor U1851 (N_1851,N_1706,N_1758);
and U1852 (N_1852,N_1703,N_1706);
nand U1853 (N_1853,N_1759,N_1789);
xnor U1854 (N_1854,N_1731,N_1707);
xor U1855 (N_1855,N_1737,N_1789);
xnor U1856 (N_1856,N_1784,N_1791);
nor U1857 (N_1857,N_1777,N_1791);
nor U1858 (N_1858,N_1773,N_1760);
nor U1859 (N_1859,N_1757,N_1711);
and U1860 (N_1860,N_1741,N_1705);
nand U1861 (N_1861,N_1776,N_1700);
and U1862 (N_1862,N_1778,N_1704);
nand U1863 (N_1863,N_1718,N_1726);
nand U1864 (N_1864,N_1752,N_1791);
xor U1865 (N_1865,N_1722,N_1792);
and U1866 (N_1866,N_1707,N_1730);
xnor U1867 (N_1867,N_1754,N_1765);
xor U1868 (N_1868,N_1744,N_1701);
xor U1869 (N_1869,N_1740,N_1738);
nor U1870 (N_1870,N_1794,N_1707);
xor U1871 (N_1871,N_1718,N_1737);
nor U1872 (N_1872,N_1739,N_1782);
xnor U1873 (N_1873,N_1725,N_1731);
nand U1874 (N_1874,N_1757,N_1737);
or U1875 (N_1875,N_1717,N_1769);
or U1876 (N_1876,N_1799,N_1703);
nand U1877 (N_1877,N_1723,N_1763);
xnor U1878 (N_1878,N_1745,N_1728);
xor U1879 (N_1879,N_1754,N_1723);
xnor U1880 (N_1880,N_1726,N_1771);
and U1881 (N_1881,N_1724,N_1798);
nand U1882 (N_1882,N_1788,N_1779);
nor U1883 (N_1883,N_1748,N_1731);
nor U1884 (N_1884,N_1701,N_1723);
nand U1885 (N_1885,N_1751,N_1723);
nand U1886 (N_1886,N_1783,N_1765);
nor U1887 (N_1887,N_1748,N_1709);
and U1888 (N_1888,N_1796,N_1725);
or U1889 (N_1889,N_1780,N_1715);
and U1890 (N_1890,N_1782,N_1735);
nand U1891 (N_1891,N_1727,N_1779);
and U1892 (N_1892,N_1775,N_1758);
nor U1893 (N_1893,N_1753,N_1795);
or U1894 (N_1894,N_1773,N_1740);
or U1895 (N_1895,N_1782,N_1744);
and U1896 (N_1896,N_1768,N_1773);
or U1897 (N_1897,N_1798,N_1781);
nor U1898 (N_1898,N_1759,N_1703);
or U1899 (N_1899,N_1744,N_1795);
or U1900 (N_1900,N_1817,N_1865);
or U1901 (N_1901,N_1872,N_1836);
or U1902 (N_1902,N_1886,N_1853);
or U1903 (N_1903,N_1889,N_1876);
nor U1904 (N_1904,N_1880,N_1867);
and U1905 (N_1905,N_1845,N_1873);
nor U1906 (N_1906,N_1825,N_1859);
or U1907 (N_1907,N_1895,N_1899);
nand U1908 (N_1908,N_1801,N_1807);
and U1909 (N_1909,N_1811,N_1885);
and U1910 (N_1910,N_1860,N_1827);
xor U1911 (N_1911,N_1802,N_1887);
or U1912 (N_1912,N_1815,N_1881);
and U1913 (N_1913,N_1821,N_1823);
or U1914 (N_1914,N_1813,N_1839);
xor U1915 (N_1915,N_1803,N_1837);
nor U1916 (N_1916,N_1851,N_1809);
or U1917 (N_1917,N_1806,N_1864);
or U1918 (N_1918,N_1863,N_1849);
and U1919 (N_1919,N_1834,N_1822);
and U1920 (N_1920,N_1898,N_1844);
nand U1921 (N_1921,N_1894,N_1826);
and U1922 (N_1922,N_1866,N_1874);
nand U1923 (N_1923,N_1848,N_1818);
nand U1924 (N_1924,N_1862,N_1884);
xnor U1925 (N_1925,N_1878,N_1882);
nand U1926 (N_1926,N_1897,N_1838);
and U1927 (N_1927,N_1896,N_1800);
nor U1928 (N_1928,N_1870,N_1840);
xor U1929 (N_1929,N_1847,N_1868);
nand U1930 (N_1930,N_1824,N_1812);
xor U1931 (N_1931,N_1888,N_1816);
or U1932 (N_1932,N_1804,N_1820);
nand U1933 (N_1933,N_1879,N_1861);
and U1934 (N_1934,N_1850,N_1852);
xor U1935 (N_1935,N_1877,N_1819);
and U1936 (N_1936,N_1858,N_1814);
nor U1937 (N_1937,N_1841,N_1883);
nand U1938 (N_1938,N_1843,N_1832);
xnor U1939 (N_1939,N_1891,N_1892);
xnor U1940 (N_1940,N_1831,N_1871);
and U1941 (N_1941,N_1856,N_1829);
nor U1942 (N_1942,N_1828,N_1808);
and U1943 (N_1943,N_1805,N_1835);
nor U1944 (N_1944,N_1857,N_1842);
xnor U1945 (N_1945,N_1810,N_1893);
or U1946 (N_1946,N_1830,N_1869);
xnor U1947 (N_1947,N_1890,N_1875);
xor U1948 (N_1948,N_1855,N_1833);
or U1949 (N_1949,N_1854,N_1846);
xor U1950 (N_1950,N_1894,N_1886);
nand U1951 (N_1951,N_1842,N_1828);
nor U1952 (N_1952,N_1896,N_1831);
nand U1953 (N_1953,N_1837,N_1872);
and U1954 (N_1954,N_1852,N_1823);
nor U1955 (N_1955,N_1802,N_1884);
nor U1956 (N_1956,N_1824,N_1836);
xnor U1957 (N_1957,N_1837,N_1882);
or U1958 (N_1958,N_1868,N_1860);
xnor U1959 (N_1959,N_1818,N_1882);
xnor U1960 (N_1960,N_1892,N_1871);
or U1961 (N_1961,N_1890,N_1811);
xor U1962 (N_1962,N_1871,N_1842);
xnor U1963 (N_1963,N_1819,N_1896);
nand U1964 (N_1964,N_1832,N_1859);
and U1965 (N_1965,N_1849,N_1846);
xor U1966 (N_1966,N_1832,N_1800);
and U1967 (N_1967,N_1870,N_1898);
xnor U1968 (N_1968,N_1830,N_1877);
xor U1969 (N_1969,N_1896,N_1818);
and U1970 (N_1970,N_1870,N_1815);
or U1971 (N_1971,N_1802,N_1888);
nor U1972 (N_1972,N_1866,N_1849);
nand U1973 (N_1973,N_1819,N_1825);
and U1974 (N_1974,N_1885,N_1820);
nand U1975 (N_1975,N_1829,N_1899);
xor U1976 (N_1976,N_1868,N_1809);
nor U1977 (N_1977,N_1821,N_1866);
xnor U1978 (N_1978,N_1853,N_1879);
or U1979 (N_1979,N_1824,N_1862);
nand U1980 (N_1980,N_1828,N_1826);
nand U1981 (N_1981,N_1876,N_1824);
and U1982 (N_1982,N_1820,N_1861);
or U1983 (N_1983,N_1858,N_1810);
and U1984 (N_1984,N_1898,N_1862);
or U1985 (N_1985,N_1866,N_1857);
or U1986 (N_1986,N_1843,N_1854);
nor U1987 (N_1987,N_1819,N_1834);
and U1988 (N_1988,N_1893,N_1802);
and U1989 (N_1989,N_1875,N_1811);
nand U1990 (N_1990,N_1839,N_1853);
or U1991 (N_1991,N_1812,N_1846);
xnor U1992 (N_1992,N_1851,N_1836);
nor U1993 (N_1993,N_1858,N_1866);
nor U1994 (N_1994,N_1832,N_1831);
or U1995 (N_1995,N_1895,N_1846);
and U1996 (N_1996,N_1806,N_1820);
or U1997 (N_1997,N_1809,N_1818);
and U1998 (N_1998,N_1805,N_1859);
nand U1999 (N_1999,N_1898,N_1804);
nand U2000 (N_2000,N_1973,N_1981);
nor U2001 (N_2001,N_1901,N_1992);
nor U2002 (N_2002,N_1980,N_1913);
nor U2003 (N_2003,N_1945,N_1986);
nor U2004 (N_2004,N_1995,N_1947);
or U2005 (N_2005,N_1965,N_1934);
or U2006 (N_2006,N_1912,N_1921);
and U2007 (N_2007,N_1918,N_1906);
nand U2008 (N_2008,N_1940,N_1954);
nor U2009 (N_2009,N_1966,N_1955);
and U2010 (N_2010,N_1914,N_1923);
nand U2011 (N_2011,N_1926,N_1910);
xnor U2012 (N_2012,N_1988,N_1967);
or U2013 (N_2013,N_1904,N_1953);
nand U2014 (N_2014,N_1963,N_1975);
nor U2015 (N_2015,N_1939,N_1984);
nand U2016 (N_2016,N_1929,N_1970);
and U2017 (N_2017,N_1948,N_1961);
xor U2018 (N_2018,N_1942,N_1978);
xor U2019 (N_2019,N_1925,N_1977);
and U2020 (N_2020,N_1959,N_1997);
nand U2021 (N_2021,N_1958,N_1927);
nand U2022 (N_2022,N_1907,N_1938);
and U2023 (N_2023,N_1943,N_1911);
nor U2024 (N_2024,N_1998,N_1962);
xnor U2025 (N_2025,N_1909,N_1983);
xor U2026 (N_2026,N_1969,N_1944);
xnor U2027 (N_2027,N_1976,N_1941);
or U2028 (N_2028,N_1994,N_1968);
and U2029 (N_2029,N_1930,N_1900);
xnor U2030 (N_2030,N_1949,N_1971);
xor U2031 (N_2031,N_1951,N_1996);
xnor U2032 (N_2032,N_1982,N_1937);
and U2033 (N_2033,N_1999,N_1920);
xnor U2034 (N_2034,N_1924,N_1972);
and U2035 (N_2035,N_1908,N_1922);
xor U2036 (N_2036,N_1990,N_1952);
nor U2037 (N_2037,N_1979,N_1987);
or U2038 (N_2038,N_1915,N_1956);
nand U2039 (N_2039,N_1932,N_1919);
or U2040 (N_2040,N_1935,N_1964);
and U2041 (N_2041,N_1928,N_1916);
and U2042 (N_2042,N_1960,N_1931);
xor U2043 (N_2043,N_1903,N_1991);
or U2044 (N_2044,N_1902,N_1993);
xor U2045 (N_2045,N_1946,N_1985);
or U2046 (N_2046,N_1905,N_1936);
and U2047 (N_2047,N_1917,N_1957);
xnor U2048 (N_2048,N_1989,N_1974);
or U2049 (N_2049,N_1950,N_1933);
and U2050 (N_2050,N_1988,N_1963);
or U2051 (N_2051,N_1993,N_1916);
xnor U2052 (N_2052,N_1975,N_1935);
nor U2053 (N_2053,N_1915,N_1964);
and U2054 (N_2054,N_1914,N_1973);
nor U2055 (N_2055,N_1943,N_1984);
or U2056 (N_2056,N_1948,N_1974);
or U2057 (N_2057,N_1906,N_1970);
or U2058 (N_2058,N_1912,N_1939);
nand U2059 (N_2059,N_1996,N_1901);
or U2060 (N_2060,N_1905,N_1925);
nand U2061 (N_2061,N_1967,N_1952);
nand U2062 (N_2062,N_1902,N_1931);
nand U2063 (N_2063,N_1912,N_1935);
nor U2064 (N_2064,N_1953,N_1987);
xor U2065 (N_2065,N_1963,N_1912);
and U2066 (N_2066,N_1965,N_1986);
and U2067 (N_2067,N_1934,N_1963);
or U2068 (N_2068,N_1978,N_1949);
nor U2069 (N_2069,N_1946,N_1938);
and U2070 (N_2070,N_1994,N_1965);
and U2071 (N_2071,N_1979,N_1925);
nand U2072 (N_2072,N_1938,N_1936);
nand U2073 (N_2073,N_1985,N_1978);
nand U2074 (N_2074,N_1927,N_1957);
nor U2075 (N_2075,N_1908,N_1917);
and U2076 (N_2076,N_1969,N_1913);
xor U2077 (N_2077,N_1947,N_1918);
nand U2078 (N_2078,N_1961,N_1969);
and U2079 (N_2079,N_1989,N_1973);
and U2080 (N_2080,N_1991,N_1940);
nand U2081 (N_2081,N_1910,N_1971);
and U2082 (N_2082,N_1907,N_1984);
and U2083 (N_2083,N_1932,N_1960);
xor U2084 (N_2084,N_1957,N_1933);
and U2085 (N_2085,N_1966,N_1912);
and U2086 (N_2086,N_1965,N_1956);
nor U2087 (N_2087,N_1936,N_1942);
nand U2088 (N_2088,N_1985,N_1981);
nand U2089 (N_2089,N_1916,N_1992);
nor U2090 (N_2090,N_1985,N_1990);
xor U2091 (N_2091,N_1969,N_1925);
or U2092 (N_2092,N_1947,N_1973);
and U2093 (N_2093,N_1983,N_1921);
and U2094 (N_2094,N_1940,N_1918);
xor U2095 (N_2095,N_1909,N_1932);
nor U2096 (N_2096,N_1998,N_1926);
and U2097 (N_2097,N_1987,N_1933);
xnor U2098 (N_2098,N_1906,N_1974);
xnor U2099 (N_2099,N_1909,N_1903);
and U2100 (N_2100,N_2029,N_2015);
nand U2101 (N_2101,N_2066,N_2019);
nand U2102 (N_2102,N_2039,N_2060);
and U2103 (N_2103,N_2017,N_2054);
and U2104 (N_2104,N_2081,N_2071);
and U2105 (N_2105,N_2084,N_2085);
nor U2106 (N_2106,N_2063,N_2086);
and U2107 (N_2107,N_2043,N_2000);
nor U2108 (N_2108,N_2094,N_2013);
xnor U2109 (N_2109,N_2062,N_2074);
or U2110 (N_2110,N_2056,N_2027);
or U2111 (N_2111,N_2005,N_2046);
or U2112 (N_2112,N_2025,N_2055);
and U2113 (N_2113,N_2014,N_2048);
nor U2114 (N_2114,N_2057,N_2042);
nand U2115 (N_2115,N_2092,N_2036);
or U2116 (N_2116,N_2088,N_2068);
nor U2117 (N_2117,N_2041,N_2020);
and U2118 (N_2118,N_2012,N_2059);
or U2119 (N_2119,N_2058,N_2073);
and U2120 (N_2120,N_2098,N_2008);
xor U2121 (N_2121,N_2079,N_2028);
xnor U2122 (N_2122,N_2089,N_2099);
nor U2123 (N_2123,N_2075,N_2003);
nand U2124 (N_2124,N_2069,N_2023);
and U2125 (N_2125,N_2049,N_2052);
and U2126 (N_2126,N_2064,N_2006);
nor U2127 (N_2127,N_2009,N_2011);
xor U2128 (N_2128,N_2076,N_2072);
nor U2129 (N_2129,N_2090,N_2082);
nor U2130 (N_2130,N_2010,N_2097);
xnor U2131 (N_2131,N_2031,N_2050);
nand U2132 (N_2132,N_2007,N_2070);
nor U2133 (N_2133,N_2002,N_2026);
or U2134 (N_2134,N_2037,N_2065);
xor U2135 (N_2135,N_2038,N_2087);
and U2136 (N_2136,N_2033,N_2061);
nor U2137 (N_2137,N_2034,N_2083);
xnor U2138 (N_2138,N_2044,N_2051);
xnor U2139 (N_2139,N_2067,N_2040);
xnor U2140 (N_2140,N_2080,N_2053);
and U2141 (N_2141,N_2045,N_2030);
xnor U2142 (N_2142,N_2035,N_2091);
nor U2143 (N_2143,N_2077,N_2018);
xnor U2144 (N_2144,N_2024,N_2047);
and U2145 (N_2145,N_2021,N_2004);
nor U2146 (N_2146,N_2096,N_2022);
or U2147 (N_2147,N_2016,N_2095);
xnor U2148 (N_2148,N_2001,N_2078);
nor U2149 (N_2149,N_2032,N_2093);
nand U2150 (N_2150,N_2037,N_2033);
xnor U2151 (N_2151,N_2047,N_2083);
nor U2152 (N_2152,N_2035,N_2004);
nand U2153 (N_2153,N_2082,N_2023);
xor U2154 (N_2154,N_2051,N_2091);
nor U2155 (N_2155,N_2095,N_2056);
nand U2156 (N_2156,N_2047,N_2062);
nand U2157 (N_2157,N_2058,N_2023);
or U2158 (N_2158,N_2021,N_2086);
nand U2159 (N_2159,N_2061,N_2043);
nand U2160 (N_2160,N_2044,N_2073);
nand U2161 (N_2161,N_2078,N_2054);
and U2162 (N_2162,N_2091,N_2068);
xnor U2163 (N_2163,N_2009,N_2074);
nand U2164 (N_2164,N_2063,N_2048);
or U2165 (N_2165,N_2061,N_2016);
or U2166 (N_2166,N_2058,N_2016);
xor U2167 (N_2167,N_2037,N_2000);
nand U2168 (N_2168,N_2023,N_2073);
nand U2169 (N_2169,N_2096,N_2040);
nand U2170 (N_2170,N_2099,N_2058);
nand U2171 (N_2171,N_2080,N_2088);
nand U2172 (N_2172,N_2073,N_2036);
or U2173 (N_2173,N_2038,N_2054);
or U2174 (N_2174,N_2086,N_2067);
nand U2175 (N_2175,N_2049,N_2083);
and U2176 (N_2176,N_2072,N_2005);
and U2177 (N_2177,N_2088,N_2098);
and U2178 (N_2178,N_2010,N_2062);
nor U2179 (N_2179,N_2070,N_2053);
nand U2180 (N_2180,N_2060,N_2035);
and U2181 (N_2181,N_2075,N_2027);
and U2182 (N_2182,N_2041,N_2037);
nand U2183 (N_2183,N_2061,N_2080);
and U2184 (N_2184,N_2072,N_2028);
nand U2185 (N_2185,N_2056,N_2082);
or U2186 (N_2186,N_2041,N_2050);
nor U2187 (N_2187,N_2066,N_2099);
nor U2188 (N_2188,N_2028,N_2096);
nand U2189 (N_2189,N_2017,N_2026);
xnor U2190 (N_2190,N_2091,N_2007);
nor U2191 (N_2191,N_2023,N_2030);
and U2192 (N_2192,N_2059,N_2079);
nor U2193 (N_2193,N_2009,N_2092);
nand U2194 (N_2194,N_2002,N_2008);
nor U2195 (N_2195,N_2080,N_2051);
xor U2196 (N_2196,N_2090,N_2008);
or U2197 (N_2197,N_2006,N_2082);
nor U2198 (N_2198,N_2098,N_2062);
or U2199 (N_2199,N_2090,N_2097);
or U2200 (N_2200,N_2169,N_2143);
xor U2201 (N_2201,N_2157,N_2120);
xor U2202 (N_2202,N_2141,N_2110);
xnor U2203 (N_2203,N_2184,N_2182);
or U2204 (N_2204,N_2144,N_2163);
xnor U2205 (N_2205,N_2176,N_2183);
xnor U2206 (N_2206,N_2118,N_2116);
xor U2207 (N_2207,N_2185,N_2149);
nand U2208 (N_2208,N_2198,N_2191);
nand U2209 (N_2209,N_2190,N_2181);
and U2210 (N_2210,N_2146,N_2117);
or U2211 (N_2211,N_2102,N_2138);
or U2212 (N_2212,N_2113,N_2112);
nand U2213 (N_2213,N_2122,N_2159);
or U2214 (N_2214,N_2133,N_2187);
nor U2215 (N_2215,N_2114,N_2170);
or U2216 (N_2216,N_2145,N_2156);
and U2217 (N_2217,N_2128,N_2127);
and U2218 (N_2218,N_2167,N_2147);
and U2219 (N_2219,N_2161,N_2188);
and U2220 (N_2220,N_2197,N_2171);
nor U2221 (N_2221,N_2103,N_2104);
and U2222 (N_2222,N_2180,N_2140);
xnor U2223 (N_2223,N_2150,N_2177);
xnor U2224 (N_2224,N_2195,N_2142);
nor U2225 (N_2225,N_2173,N_2189);
xor U2226 (N_2226,N_2106,N_2139);
nor U2227 (N_2227,N_2165,N_2100);
nor U2228 (N_2228,N_2123,N_2155);
xnor U2229 (N_2229,N_2111,N_2178);
nor U2230 (N_2230,N_2154,N_2192);
nand U2231 (N_2231,N_2162,N_2131);
nor U2232 (N_2232,N_2196,N_2125);
and U2233 (N_2233,N_2175,N_2174);
and U2234 (N_2234,N_2101,N_2194);
nor U2235 (N_2235,N_2130,N_2121);
or U2236 (N_2236,N_2119,N_2164);
nor U2237 (N_2237,N_2172,N_2179);
nor U2238 (N_2238,N_2153,N_2166);
nor U2239 (N_2239,N_2124,N_2135);
or U2240 (N_2240,N_2129,N_2132);
nand U2241 (N_2241,N_2105,N_2152);
xnor U2242 (N_2242,N_2134,N_2126);
nand U2243 (N_2243,N_2137,N_2136);
nor U2244 (N_2244,N_2160,N_2115);
and U2245 (N_2245,N_2158,N_2148);
nand U2246 (N_2246,N_2186,N_2109);
or U2247 (N_2247,N_2108,N_2193);
nor U2248 (N_2248,N_2199,N_2168);
xnor U2249 (N_2249,N_2107,N_2151);
xnor U2250 (N_2250,N_2140,N_2126);
xnor U2251 (N_2251,N_2161,N_2128);
xor U2252 (N_2252,N_2193,N_2172);
nor U2253 (N_2253,N_2102,N_2133);
nand U2254 (N_2254,N_2121,N_2185);
and U2255 (N_2255,N_2162,N_2175);
nor U2256 (N_2256,N_2163,N_2143);
xnor U2257 (N_2257,N_2157,N_2177);
xor U2258 (N_2258,N_2134,N_2145);
or U2259 (N_2259,N_2129,N_2165);
xnor U2260 (N_2260,N_2145,N_2173);
nand U2261 (N_2261,N_2165,N_2142);
nor U2262 (N_2262,N_2184,N_2119);
xor U2263 (N_2263,N_2185,N_2122);
or U2264 (N_2264,N_2192,N_2132);
or U2265 (N_2265,N_2149,N_2125);
or U2266 (N_2266,N_2164,N_2191);
or U2267 (N_2267,N_2127,N_2139);
or U2268 (N_2268,N_2103,N_2199);
nor U2269 (N_2269,N_2151,N_2181);
xnor U2270 (N_2270,N_2185,N_2162);
or U2271 (N_2271,N_2123,N_2105);
or U2272 (N_2272,N_2111,N_2179);
nand U2273 (N_2273,N_2175,N_2166);
nand U2274 (N_2274,N_2122,N_2182);
or U2275 (N_2275,N_2199,N_2167);
and U2276 (N_2276,N_2176,N_2190);
nor U2277 (N_2277,N_2109,N_2140);
nand U2278 (N_2278,N_2134,N_2177);
xor U2279 (N_2279,N_2100,N_2102);
nor U2280 (N_2280,N_2123,N_2176);
nand U2281 (N_2281,N_2150,N_2138);
nor U2282 (N_2282,N_2164,N_2181);
nor U2283 (N_2283,N_2134,N_2122);
nand U2284 (N_2284,N_2162,N_2168);
nand U2285 (N_2285,N_2123,N_2153);
and U2286 (N_2286,N_2124,N_2134);
xnor U2287 (N_2287,N_2144,N_2128);
nor U2288 (N_2288,N_2188,N_2172);
nand U2289 (N_2289,N_2103,N_2154);
nand U2290 (N_2290,N_2163,N_2184);
nand U2291 (N_2291,N_2119,N_2166);
nand U2292 (N_2292,N_2153,N_2168);
xor U2293 (N_2293,N_2116,N_2110);
and U2294 (N_2294,N_2148,N_2101);
and U2295 (N_2295,N_2145,N_2157);
nand U2296 (N_2296,N_2144,N_2153);
nand U2297 (N_2297,N_2168,N_2190);
and U2298 (N_2298,N_2121,N_2119);
nor U2299 (N_2299,N_2131,N_2192);
nand U2300 (N_2300,N_2277,N_2273);
nand U2301 (N_2301,N_2234,N_2271);
and U2302 (N_2302,N_2263,N_2244);
xor U2303 (N_2303,N_2243,N_2269);
nand U2304 (N_2304,N_2268,N_2290);
nor U2305 (N_2305,N_2232,N_2236);
nand U2306 (N_2306,N_2251,N_2213);
or U2307 (N_2307,N_2227,N_2279);
xnor U2308 (N_2308,N_2250,N_2267);
and U2309 (N_2309,N_2201,N_2286);
nand U2310 (N_2310,N_2288,N_2247);
nor U2311 (N_2311,N_2298,N_2294);
nand U2312 (N_2312,N_2262,N_2221);
nand U2313 (N_2313,N_2278,N_2259);
or U2314 (N_2314,N_2235,N_2241);
nand U2315 (N_2315,N_2295,N_2257);
nor U2316 (N_2316,N_2210,N_2216);
xnor U2317 (N_2317,N_2228,N_2224);
and U2318 (N_2318,N_2214,N_2297);
xor U2319 (N_2319,N_2208,N_2287);
nor U2320 (N_2320,N_2264,N_2209);
nand U2321 (N_2321,N_2296,N_2248);
nor U2322 (N_2322,N_2299,N_2292);
xnor U2323 (N_2323,N_2217,N_2239);
or U2324 (N_2324,N_2289,N_2276);
or U2325 (N_2325,N_2212,N_2260);
xnor U2326 (N_2326,N_2200,N_2270);
and U2327 (N_2327,N_2242,N_2275);
or U2328 (N_2328,N_2205,N_2256);
xnor U2329 (N_2329,N_2253,N_2246);
or U2330 (N_2330,N_2202,N_2231);
and U2331 (N_2331,N_2258,N_2240);
nand U2332 (N_2332,N_2249,N_2274);
xor U2333 (N_2333,N_2283,N_2293);
nor U2334 (N_2334,N_2284,N_2206);
or U2335 (N_2335,N_2245,N_2266);
nor U2336 (N_2336,N_2238,N_2211);
xor U2337 (N_2337,N_2204,N_2203);
xor U2338 (N_2338,N_2282,N_2229);
or U2339 (N_2339,N_2223,N_2220);
nor U2340 (N_2340,N_2254,N_2215);
nor U2341 (N_2341,N_2230,N_2218);
nor U2342 (N_2342,N_2219,N_2207);
and U2343 (N_2343,N_2252,N_2225);
or U2344 (N_2344,N_2233,N_2285);
nand U2345 (N_2345,N_2255,N_2280);
nor U2346 (N_2346,N_2265,N_2226);
or U2347 (N_2347,N_2237,N_2222);
and U2348 (N_2348,N_2281,N_2272);
or U2349 (N_2349,N_2261,N_2291);
and U2350 (N_2350,N_2262,N_2206);
nor U2351 (N_2351,N_2289,N_2210);
and U2352 (N_2352,N_2202,N_2293);
or U2353 (N_2353,N_2292,N_2244);
nor U2354 (N_2354,N_2249,N_2210);
xor U2355 (N_2355,N_2283,N_2260);
or U2356 (N_2356,N_2240,N_2263);
or U2357 (N_2357,N_2296,N_2268);
nand U2358 (N_2358,N_2200,N_2224);
nor U2359 (N_2359,N_2233,N_2292);
nor U2360 (N_2360,N_2245,N_2232);
or U2361 (N_2361,N_2244,N_2256);
and U2362 (N_2362,N_2219,N_2279);
or U2363 (N_2363,N_2228,N_2214);
nand U2364 (N_2364,N_2201,N_2284);
nand U2365 (N_2365,N_2236,N_2214);
nand U2366 (N_2366,N_2270,N_2247);
nand U2367 (N_2367,N_2279,N_2235);
nor U2368 (N_2368,N_2282,N_2221);
nand U2369 (N_2369,N_2222,N_2296);
or U2370 (N_2370,N_2265,N_2200);
and U2371 (N_2371,N_2264,N_2226);
or U2372 (N_2372,N_2292,N_2257);
nor U2373 (N_2373,N_2217,N_2245);
nor U2374 (N_2374,N_2205,N_2268);
nand U2375 (N_2375,N_2236,N_2274);
and U2376 (N_2376,N_2294,N_2250);
or U2377 (N_2377,N_2273,N_2252);
nor U2378 (N_2378,N_2278,N_2202);
xor U2379 (N_2379,N_2223,N_2250);
or U2380 (N_2380,N_2229,N_2270);
nand U2381 (N_2381,N_2288,N_2255);
xnor U2382 (N_2382,N_2285,N_2240);
xnor U2383 (N_2383,N_2257,N_2279);
and U2384 (N_2384,N_2224,N_2265);
and U2385 (N_2385,N_2211,N_2255);
xor U2386 (N_2386,N_2233,N_2273);
or U2387 (N_2387,N_2272,N_2296);
or U2388 (N_2388,N_2255,N_2249);
nand U2389 (N_2389,N_2295,N_2277);
nor U2390 (N_2390,N_2269,N_2201);
and U2391 (N_2391,N_2239,N_2277);
nor U2392 (N_2392,N_2253,N_2222);
xor U2393 (N_2393,N_2298,N_2255);
xnor U2394 (N_2394,N_2264,N_2283);
or U2395 (N_2395,N_2251,N_2281);
and U2396 (N_2396,N_2244,N_2210);
nor U2397 (N_2397,N_2212,N_2290);
and U2398 (N_2398,N_2264,N_2299);
and U2399 (N_2399,N_2201,N_2257);
xor U2400 (N_2400,N_2394,N_2308);
and U2401 (N_2401,N_2338,N_2378);
and U2402 (N_2402,N_2384,N_2319);
or U2403 (N_2403,N_2322,N_2367);
xnor U2404 (N_2404,N_2302,N_2301);
xnor U2405 (N_2405,N_2383,N_2387);
and U2406 (N_2406,N_2329,N_2368);
nand U2407 (N_2407,N_2300,N_2390);
or U2408 (N_2408,N_2366,N_2375);
or U2409 (N_2409,N_2357,N_2381);
xor U2410 (N_2410,N_2376,N_2309);
xnor U2411 (N_2411,N_2356,N_2398);
nor U2412 (N_2412,N_2328,N_2347);
nor U2413 (N_2413,N_2336,N_2343);
xor U2414 (N_2414,N_2303,N_2314);
and U2415 (N_2415,N_2345,N_2323);
nand U2416 (N_2416,N_2310,N_2353);
and U2417 (N_2417,N_2316,N_2327);
xor U2418 (N_2418,N_2324,N_2351);
xnor U2419 (N_2419,N_2306,N_2313);
nand U2420 (N_2420,N_2382,N_2307);
nor U2421 (N_2421,N_2371,N_2385);
nor U2422 (N_2422,N_2388,N_2305);
or U2423 (N_2423,N_2393,N_2339);
nor U2424 (N_2424,N_2365,N_2349);
xor U2425 (N_2425,N_2379,N_2374);
nor U2426 (N_2426,N_2392,N_2331);
or U2427 (N_2427,N_2311,N_2330);
xnor U2428 (N_2428,N_2317,N_2362);
xnor U2429 (N_2429,N_2358,N_2363);
and U2430 (N_2430,N_2377,N_2373);
xor U2431 (N_2431,N_2335,N_2380);
nand U2432 (N_2432,N_2315,N_2372);
or U2433 (N_2433,N_2304,N_2364);
xnor U2434 (N_2434,N_2320,N_2348);
xnor U2435 (N_2435,N_2352,N_2321);
or U2436 (N_2436,N_2334,N_2396);
and U2437 (N_2437,N_2361,N_2397);
nand U2438 (N_2438,N_2350,N_2370);
xnor U2439 (N_2439,N_2399,N_2389);
nand U2440 (N_2440,N_2340,N_2346);
nor U2441 (N_2441,N_2342,N_2344);
nor U2442 (N_2442,N_2318,N_2360);
nor U2443 (N_2443,N_2325,N_2395);
or U2444 (N_2444,N_2355,N_2386);
and U2445 (N_2445,N_2333,N_2341);
or U2446 (N_2446,N_2391,N_2332);
and U2447 (N_2447,N_2326,N_2359);
nand U2448 (N_2448,N_2312,N_2337);
nor U2449 (N_2449,N_2354,N_2369);
xor U2450 (N_2450,N_2389,N_2364);
and U2451 (N_2451,N_2376,N_2343);
and U2452 (N_2452,N_2386,N_2357);
xnor U2453 (N_2453,N_2325,N_2373);
nor U2454 (N_2454,N_2339,N_2353);
or U2455 (N_2455,N_2370,N_2340);
or U2456 (N_2456,N_2308,N_2383);
nand U2457 (N_2457,N_2340,N_2325);
nor U2458 (N_2458,N_2356,N_2357);
and U2459 (N_2459,N_2341,N_2397);
and U2460 (N_2460,N_2386,N_2370);
xnor U2461 (N_2461,N_2362,N_2341);
and U2462 (N_2462,N_2352,N_2392);
xnor U2463 (N_2463,N_2318,N_2379);
xor U2464 (N_2464,N_2395,N_2300);
or U2465 (N_2465,N_2349,N_2387);
nor U2466 (N_2466,N_2393,N_2371);
nand U2467 (N_2467,N_2333,N_2383);
nor U2468 (N_2468,N_2315,N_2350);
nor U2469 (N_2469,N_2305,N_2358);
and U2470 (N_2470,N_2379,N_2322);
xnor U2471 (N_2471,N_2312,N_2389);
nor U2472 (N_2472,N_2384,N_2393);
or U2473 (N_2473,N_2343,N_2305);
nor U2474 (N_2474,N_2313,N_2354);
xnor U2475 (N_2475,N_2361,N_2335);
nand U2476 (N_2476,N_2306,N_2314);
nor U2477 (N_2477,N_2359,N_2381);
or U2478 (N_2478,N_2374,N_2321);
or U2479 (N_2479,N_2351,N_2366);
xor U2480 (N_2480,N_2348,N_2325);
and U2481 (N_2481,N_2338,N_2305);
and U2482 (N_2482,N_2340,N_2362);
nor U2483 (N_2483,N_2352,N_2373);
and U2484 (N_2484,N_2393,N_2351);
xor U2485 (N_2485,N_2376,N_2397);
xnor U2486 (N_2486,N_2345,N_2336);
or U2487 (N_2487,N_2382,N_2325);
xor U2488 (N_2488,N_2370,N_2355);
xor U2489 (N_2489,N_2363,N_2338);
or U2490 (N_2490,N_2319,N_2308);
nor U2491 (N_2491,N_2312,N_2379);
xnor U2492 (N_2492,N_2312,N_2310);
xor U2493 (N_2493,N_2312,N_2380);
xor U2494 (N_2494,N_2310,N_2335);
nor U2495 (N_2495,N_2334,N_2376);
nor U2496 (N_2496,N_2311,N_2383);
nand U2497 (N_2497,N_2345,N_2318);
and U2498 (N_2498,N_2382,N_2384);
nor U2499 (N_2499,N_2337,N_2345);
or U2500 (N_2500,N_2434,N_2421);
nor U2501 (N_2501,N_2482,N_2475);
and U2502 (N_2502,N_2493,N_2402);
nand U2503 (N_2503,N_2444,N_2450);
or U2504 (N_2504,N_2484,N_2423);
nor U2505 (N_2505,N_2454,N_2478);
and U2506 (N_2506,N_2472,N_2408);
xnor U2507 (N_2507,N_2433,N_2486);
nor U2508 (N_2508,N_2463,N_2452);
xor U2509 (N_2509,N_2449,N_2474);
xor U2510 (N_2510,N_2490,N_2424);
and U2511 (N_2511,N_2487,N_2414);
and U2512 (N_2512,N_2477,N_2473);
or U2513 (N_2513,N_2494,N_2426);
nor U2514 (N_2514,N_2411,N_2457);
nor U2515 (N_2515,N_2496,N_2455);
nand U2516 (N_2516,N_2442,N_2415);
or U2517 (N_2517,N_2435,N_2405);
nor U2518 (N_2518,N_2438,N_2495);
and U2519 (N_2519,N_2469,N_2497);
xnor U2520 (N_2520,N_2403,N_2400);
xnor U2521 (N_2521,N_2413,N_2499);
and U2522 (N_2522,N_2417,N_2464);
or U2523 (N_2523,N_2476,N_2489);
xor U2524 (N_2524,N_2458,N_2429);
xnor U2525 (N_2525,N_2447,N_2453);
xnor U2526 (N_2526,N_2462,N_2466);
nand U2527 (N_2527,N_2443,N_2491);
or U2528 (N_2528,N_2448,N_2460);
and U2529 (N_2529,N_2404,N_2427);
and U2530 (N_2530,N_2459,N_2465);
nor U2531 (N_2531,N_2430,N_2439);
or U2532 (N_2532,N_2445,N_2461);
or U2533 (N_2533,N_2428,N_2451);
and U2534 (N_2534,N_2468,N_2480);
and U2535 (N_2535,N_2446,N_2479);
nor U2536 (N_2536,N_2467,N_2492);
nand U2537 (N_2537,N_2456,N_2437);
nand U2538 (N_2538,N_2401,N_2485);
nor U2539 (N_2539,N_2431,N_2422);
or U2540 (N_2540,N_2488,N_2418);
nand U2541 (N_2541,N_2420,N_2498);
and U2542 (N_2542,N_2440,N_2409);
nor U2543 (N_2543,N_2412,N_2483);
nor U2544 (N_2544,N_2471,N_2419);
nor U2545 (N_2545,N_2441,N_2436);
xnor U2546 (N_2546,N_2432,N_2416);
and U2547 (N_2547,N_2481,N_2406);
nand U2548 (N_2548,N_2470,N_2410);
or U2549 (N_2549,N_2425,N_2407);
and U2550 (N_2550,N_2456,N_2488);
and U2551 (N_2551,N_2448,N_2430);
or U2552 (N_2552,N_2439,N_2434);
xnor U2553 (N_2553,N_2430,N_2432);
nor U2554 (N_2554,N_2448,N_2467);
nor U2555 (N_2555,N_2438,N_2421);
xnor U2556 (N_2556,N_2496,N_2414);
nand U2557 (N_2557,N_2415,N_2477);
or U2558 (N_2558,N_2477,N_2431);
nor U2559 (N_2559,N_2492,N_2432);
nand U2560 (N_2560,N_2440,N_2436);
or U2561 (N_2561,N_2431,N_2465);
nor U2562 (N_2562,N_2487,N_2437);
nand U2563 (N_2563,N_2474,N_2430);
nor U2564 (N_2564,N_2429,N_2414);
and U2565 (N_2565,N_2493,N_2405);
xor U2566 (N_2566,N_2418,N_2404);
nand U2567 (N_2567,N_2403,N_2471);
nand U2568 (N_2568,N_2484,N_2463);
nand U2569 (N_2569,N_2464,N_2492);
nand U2570 (N_2570,N_2410,N_2446);
and U2571 (N_2571,N_2414,N_2448);
nand U2572 (N_2572,N_2427,N_2454);
nand U2573 (N_2573,N_2417,N_2426);
xor U2574 (N_2574,N_2458,N_2488);
or U2575 (N_2575,N_2472,N_2458);
xor U2576 (N_2576,N_2459,N_2423);
and U2577 (N_2577,N_2404,N_2412);
nor U2578 (N_2578,N_2473,N_2415);
and U2579 (N_2579,N_2460,N_2464);
and U2580 (N_2580,N_2435,N_2447);
xnor U2581 (N_2581,N_2427,N_2403);
and U2582 (N_2582,N_2414,N_2470);
and U2583 (N_2583,N_2439,N_2422);
nor U2584 (N_2584,N_2452,N_2410);
nand U2585 (N_2585,N_2466,N_2479);
nor U2586 (N_2586,N_2452,N_2466);
nand U2587 (N_2587,N_2498,N_2421);
nand U2588 (N_2588,N_2484,N_2444);
nand U2589 (N_2589,N_2414,N_2476);
xnor U2590 (N_2590,N_2434,N_2435);
nor U2591 (N_2591,N_2467,N_2490);
nand U2592 (N_2592,N_2472,N_2497);
nor U2593 (N_2593,N_2489,N_2497);
nand U2594 (N_2594,N_2473,N_2484);
nand U2595 (N_2595,N_2407,N_2411);
nand U2596 (N_2596,N_2481,N_2444);
or U2597 (N_2597,N_2453,N_2468);
or U2598 (N_2598,N_2427,N_2449);
and U2599 (N_2599,N_2426,N_2463);
and U2600 (N_2600,N_2550,N_2541);
nor U2601 (N_2601,N_2503,N_2516);
and U2602 (N_2602,N_2543,N_2506);
nor U2603 (N_2603,N_2590,N_2599);
nand U2604 (N_2604,N_2597,N_2589);
and U2605 (N_2605,N_2560,N_2500);
nand U2606 (N_2606,N_2542,N_2548);
nand U2607 (N_2607,N_2524,N_2565);
nand U2608 (N_2608,N_2518,N_2585);
nor U2609 (N_2609,N_2593,N_2551);
or U2610 (N_2610,N_2569,N_2568);
xor U2611 (N_2611,N_2577,N_2526);
nand U2612 (N_2612,N_2538,N_2505);
nor U2613 (N_2613,N_2523,N_2509);
and U2614 (N_2614,N_2515,N_2508);
and U2615 (N_2615,N_2579,N_2535);
and U2616 (N_2616,N_2557,N_2582);
nor U2617 (N_2617,N_2576,N_2529);
nor U2618 (N_2618,N_2555,N_2536);
xor U2619 (N_2619,N_2513,N_2587);
xor U2620 (N_2620,N_2559,N_2507);
and U2621 (N_2621,N_2521,N_2595);
nand U2622 (N_2622,N_2522,N_2530);
and U2623 (N_2623,N_2511,N_2562);
nand U2624 (N_2624,N_2567,N_2502);
nor U2625 (N_2625,N_2574,N_2534);
or U2626 (N_2626,N_2592,N_2546);
or U2627 (N_2627,N_2591,N_2564);
nor U2628 (N_2628,N_2566,N_2561);
or U2629 (N_2629,N_2527,N_2533);
nor U2630 (N_2630,N_2544,N_2532);
and U2631 (N_2631,N_2572,N_2580);
nand U2632 (N_2632,N_2504,N_2552);
or U2633 (N_2633,N_2547,N_2588);
nand U2634 (N_2634,N_2510,N_2596);
and U2635 (N_2635,N_2531,N_2570);
and U2636 (N_2636,N_2571,N_2501);
xor U2637 (N_2637,N_2563,N_2553);
nor U2638 (N_2638,N_2583,N_2573);
xnor U2639 (N_2639,N_2556,N_2578);
nand U2640 (N_2640,N_2554,N_2537);
or U2641 (N_2641,N_2584,N_2581);
and U2642 (N_2642,N_2512,N_2520);
and U2643 (N_2643,N_2528,N_2525);
or U2644 (N_2644,N_2586,N_2598);
nand U2645 (N_2645,N_2558,N_2539);
nor U2646 (N_2646,N_2514,N_2575);
nor U2647 (N_2647,N_2545,N_2540);
nand U2648 (N_2648,N_2517,N_2594);
nand U2649 (N_2649,N_2519,N_2549);
nor U2650 (N_2650,N_2539,N_2544);
nor U2651 (N_2651,N_2573,N_2582);
nor U2652 (N_2652,N_2559,N_2566);
xor U2653 (N_2653,N_2549,N_2514);
xnor U2654 (N_2654,N_2542,N_2547);
nor U2655 (N_2655,N_2594,N_2565);
nand U2656 (N_2656,N_2562,N_2535);
xnor U2657 (N_2657,N_2583,N_2544);
and U2658 (N_2658,N_2592,N_2596);
xor U2659 (N_2659,N_2531,N_2509);
and U2660 (N_2660,N_2519,N_2576);
xor U2661 (N_2661,N_2536,N_2560);
nor U2662 (N_2662,N_2552,N_2558);
and U2663 (N_2663,N_2556,N_2545);
and U2664 (N_2664,N_2529,N_2509);
nor U2665 (N_2665,N_2578,N_2540);
nand U2666 (N_2666,N_2581,N_2566);
and U2667 (N_2667,N_2504,N_2558);
nor U2668 (N_2668,N_2575,N_2553);
or U2669 (N_2669,N_2571,N_2550);
and U2670 (N_2670,N_2563,N_2564);
nand U2671 (N_2671,N_2549,N_2510);
nor U2672 (N_2672,N_2584,N_2508);
nor U2673 (N_2673,N_2530,N_2580);
nand U2674 (N_2674,N_2544,N_2554);
nor U2675 (N_2675,N_2562,N_2583);
and U2676 (N_2676,N_2565,N_2539);
xnor U2677 (N_2677,N_2540,N_2566);
nand U2678 (N_2678,N_2544,N_2543);
nand U2679 (N_2679,N_2536,N_2578);
nand U2680 (N_2680,N_2549,N_2583);
and U2681 (N_2681,N_2567,N_2564);
nand U2682 (N_2682,N_2593,N_2584);
xnor U2683 (N_2683,N_2538,N_2582);
nand U2684 (N_2684,N_2586,N_2519);
nor U2685 (N_2685,N_2583,N_2548);
nand U2686 (N_2686,N_2521,N_2539);
nor U2687 (N_2687,N_2501,N_2547);
nor U2688 (N_2688,N_2587,N_2588);
or U2689 (N_2689,N_2526,N_2515);
or U2690 (N_2690,N_2532,N_2547);
xor U2691 (N_2691,N_2581,N_2576);
or U2692 (N_2692,N_2585,N_2553);
or U2693 (N_2693,N_2568,N_2596);
nor U2694 (N_2694,N_2522,N_2505);
nor U2695 (N_2695,N_2562,N_2542);
xor U2696 (N_2696,N_2583,N_2580);
and U2697 (N_2697,N_2589,N_2588);
xnor U2698 (N_2698,N_2590,N_2598);
nor U2699 (N_2699,N_2567,N_2500);
xor U2700 (N_2700,N_2617,N_2604);
or U2701 (N_2701,N_2673,N_2648);
xor U2702 (N_2702,N_2664,N_2678);
nor U2703 (N_2703,N_2644,N_2692);
nand U2704 (N_2704,N_2618,N_2683);
and U2705 (N_2705,N_2633,N_2666);
nor U2706 (N_2706,N_2600,N_2626);
nor U2707 (N_2707,N_2646,N_2651);
nor U2708 (N_2708,N_2643,N_2614);
or U2709 (N_2709,N_2625,N_2656);
and U2710 (N_2710,N_2647,N_2686);
or U2711 (N_2711,N_2663,N_2662);
nor U2712 (N_2712,N_2637,N_2695);
xnor U2713 (N_2713,N_2671,N_2681);
or U2714 (N_2714,N_2606,N_2658);
nand U2715 (N_2715,N_2690,N_2669);
and U2716 (N_2716,N_2632,N_2605);
and U2717 (N_2717,N_2650,N_2685);
and U2718 (N_2718,N_2602,N_2620);
nand U2719 (N_2719,N_2624,N_2608);
and U2720 (N_2720,N_2616,N_2612);
nand U2721 (N_2721,N_2688,N_2615);
and U2722 (N_2722,N_2672,N_2691);
xnor U2723 (N_2723,N_2634,N_2649);
nand U2724 (N_2724,N_2603,N_2670);
nand U2725 (N_2725,N_2653,N_2610);
xnor U2726 (N_2726,N_2641,N_2689);
and U2727 (N_2727,N_2657,N_2642);
xor U2728 (N_2728,N_2611,N_2694);
xnor U2729 (N_2729,N_2676,N_2682);
and U2730 (N_2730,N_2640,N_2645);
nor U2731 (N_2731,N_2696,N_2677);
xor U2732 (N_2732,N_2693,N_2667);
xor U2733 (N_2733,N_2655,N_2679);
nor U2734 (N_2734,N_2627,N_2631);
nand U2735 (N_2735,N_2684,N_2601);
xnor U2736 (N_2736,N_2607,N_2652);
xor U2737 (N_2737,N_2697,N_2639);
or U2738 (N_2738,N_2638,N_2630);
and U2739 (N_2739,N_2622,N_2636);
nor U2740 (N_2740,N_2680,N_2613);
and U2741 (N_2741,N_2699,N_2660);
or U2742 (N_2742,N_2675,N_2623);
nor U2743 (N_2743,N_2609,N_2635);
nor U2744 (N_2744,N_2621,N_2628);
xor U2745 (N_2745,N_2668,N_2661);
nor U2746 (N_2746,N_2619,N_2665);
and U2747 (N_2747,N_2654,N_2674);
nand U2748 (N_2748,N_2698,N_2629);
and U2749 (N_2749,N_2687,N_2659);
and U2750 (N_2750,N_2617,N_2602);
nand U2751 (N_2751,N_2650,N_2625);
nor U2752 (N_2752,N_2625,N_2626);
and U2753 (N_2753,N_2625,N_2639);
nand U2754 (N_2754,N_2659,N_2698);
nand U2755 (N_2755,N_2615,N_2679);
and U2756 (N_2756,N_2605,N_2666);
or U2757 (N_2757,N_2686,N_2687);
and U2758 (N_2758,N_2607,N_2669);
and U2759 (N_2759,N_2604,N_2641);
or U2760 (N_2760,N_2697,N_2684);
and U2761 (N_2761,N_2681,N_2664);
nor U2762 (N_2762,N_2608,N_2603);
nor U2763 (N_2763,N_2677,N_2614);
nand U2764 (N_2764,N_2633,N_2642);
or U2765 (N_2765,N_2680,N_2660);
or U2766 (N_2766,N_2640,N_2629);
xnor U2767 (N_2767,N_2625,N_2654);
or U2768 (N_2768,N_2676,N_2618);
nor U2769 (N_2769,N_2656,N_2665);
nand U2770 (N_2770,N_2609,N_2624);
or U2771 (N_2771,N_2628,N_2601);
and U2772 (N_2772,N_2626,N_2659);
nand U2773 (N_2773,N_2603,N_2644);
or U2774 (N_2774,N_2671,N_2697);
xnor U2775 (N_2775,N_2674,N_2645);
xnor U2776 (N_2776,N_2602,N_2647);
or U2777 (N_2777,N_2608,N_2655);
or U2778 (N_2778,N_2670,N_2620);
and U2779 (N_2779,N_2620,N_2682);
and U2780 (N_2780,N_2638,N_2698);
nor U2781 (N_2781,N_2693,N_2606);
and U2782 (N_2782,N_2644,N_2661);
and U2783 (N_2783,N_2640,N_2612);
nor U2784 (N_2784,N_2677,N_2682);
and U2785 (N_2785,N_2656,N_2676);
xnor U2786 (N_2786,N_2681,N_2685);
nor U2787 (N_2787,N_2624,N_2694);
xor U2788 (N_2788,N_2613,N_2693);
or U2789 (N_2789,N_2679,N_2656);
and U2790 (N_2790,N_2684,N_2696);
nor U2791 (N_2791,N_2604,N_2670);
and U2792 (N_2792,N_2698,N_2607);
and U2793 (N_2793,N_2625,N_2645);
and U2794 (N_2794,N_2619,N_2648);
nand U2795 (N_2795,N_2632,N_2602);
or U2796 (N_2796,N_2683,N_2616);
xnor U2797 (N_2797,N_2663,N_2618);
xnor U2798 (N_2798,N_2694,N_2632);
nand U2799 (N_2799,N_2627,N_2611);
nand U2800 (N_2800,N_2765,N_2731);
xor U2801 (N_2801,N_2777,N_2723);
nor U2802 (N_2802,N_2729,N_2781);
nor U2803 (N_2803,N_2745,N_2763);
nor U2804 (N_2804,N_2743,N_2741);
or U2805 (N_2805,N_2767,N_2785);
or U2806 (N_2806,N_2780,N_2733);
xor U2807 (N_2807,N_2758,N_2782);
nand U2808 (N_2808,N_2738,N_2751);
nor U2809 (N_2809,N_2728,N_2706);
or U2810 (N_2810,N_2714,N_2716);
or U2811 (N_2811,N_2725,N_2724);
or U2812 (N_2812,N_2702,N_2786);
nand U2813 (N_2813,N_2791,N_2754);
and U2814 (N_2814,N_2710,N_2713);
nand U2815 (N_2815,N_2736,N_2712);
xor U2816 (N_2816,N_2707,N_2726);
nand U2817 (N_2817,N_2737,N_2704);
nor U2818 (N_2818,N_2760,N_2730);
xor U2819 (N_2819,N_2766,N_2740);
nand U2820 (N_2820,N_2718,N_2739);
and U2821 (N_2821,N_2717,N_2701);
and U2822 (N_2822,N_2788,N_2794);
nand U2823 (N_2823,N_2773,N_2753);
xnor U2824 (N_2824,N_2746,N_2727);
nand U2825 (N_2825,N_2784,N_2711);
nor U2826 (N_2826,N_2769,N_2795);
and U2827 (N_2827,N_2742,N_2792);
or U2828 (N_2828,N_2756,N_2735);
or U2829 (N_2829,N_2700,N_2798);
nand U2830 (N_2830,N_2734,N_2719);
nor U2831 (N_2831,N_2774,N_2757);
and U2832 (N_2832,N_2797,N_2752);
and U2833 (N_2833,N_2761,N_2720);
xnor U2834 (N_2834,N_2747,N_2771);
or U2835 (N_2835,N_2759,N_2779);
nand U2836 (N_2836,N_2770,N_2787);
nand U2837 (N_2837,N_2764,N_2721);
or U2838 (N_2838,N_2775,N_2722);
nor U2839 (N_2839,N_2709,N_2744);
or U2840 (N_2840,N_2796,N_2715);
and U2841 (N_2841,N_2778,N_2708);
or U2842 (N_2842,N_2793,N_2768);
nor U2843 (N_2843,N_2799,N_2790);
nor U2844 (N_2844,N_2776,N_2789);
nand U2845 (N_2845,N_2748,N_2772);
and U2846 (N_2846,N_2749,N_2703);
nor U2847 (N_2847,N_2705,N_2750);
and U2848 (N_2848,N_2755,N_2732);
and U2849 (N_2849,N_2783,N_2762);
nor U2850 (N_2850,N_2776,N_2708);
xor U2851 (N_2851,N_2755,N_2748);
or U2852 (N_2852,N_2773,N_2724);
nor U2853 (N_2853,N_2707,N_2761);
nand U2854 (N_2854,N_2714,N_2701);
and U2855 (N_2855,N_2744,N_2794);
nor U2856 (N_2856,N_2743,N_2705);
xnor U2857 (N_2857,N_2761,N_2775);
or U2858 (N_2858,N_2785,N_2788);
nand U2859 (N_2859,N_2711,N_2727);
nor U2860 (N_2860,N_2771,N_2797);
xnor U2861 (N_2861,N_2783,N_2716);
or U2862 (N_2862,N_2738,N_2784);
xor U2863 (N_2863,N_2733,N_2720);
or U2864 (N_2864,N_2777,N_2700);
and U2865 (N_2865,N_2750,N_2793);
xor U2866 (N_2866,N_2799,N_2720);
and U2867 (N_2867,N_2748,N_2792);
and U2868 (N_2868,N_2723,N_2700);
nand U2869 (N_2869,N_2733,N_2701);
xor U2870 (N_2870,N_2722,N_2781);
and U2871 (N_2871,N_2782,N_2750);
or U2872 (N_2872,N_2733,N_2795);
nand U2873 (N_2873,N_2767,N_2771);
and U2874 (N_2874,N_2750,N_2727);
nand U2875 (N_2875,N_2774,N_2729);
or U2876 (N_2876,N_2760,N_2763);
and U2877 (N_2877,N_2709,N_2732);
or U2878 (N_2878,N_2792,N_2724);
nor U2879 (N_2879,N_2709,N_2752);
xnor U2880 (N_2880,N_2728,N_2766);
or U2881 (N_2881,N_2739,N_2719);
and U2882 (N_2882,N_2757,N_2796);
xor U2883 (N_2883,N_2710,N_2739);
nor U2884 (N_2884,N_2733,N_2773);
and U2885 (N_2885,N_2716,N_2790);
or U2886 (N_2886,N_2765,N_2791);
and U2887 (N_2887,N_2741,N_2794);
nand U2888 (N_2888,N_2718,N_2730);
or U2889 (N_2889,N_2721,N_2766);
or U2890 (N_2890,N_2739,N_2738);
nor U2891 (N_2891,N_2710,N_2730);
nor U2892 (N_2892,N_2778,N_2740);
and U2893 (N_2893,N_2764,N_2780);
xor U2894 (N_2894,N_2753,N_2719);
nand U2895 (N_2895,N_2765,N_2708);
nand U2896 (N_2896,N_2711,N_2730);
and U2897 (N_2897,N_2795,N_2784);
and U2898 (N_2898,N_2725,N_2721);
or U2899 (N_2899,N_2703,N_2702);
and U2900 (N_2900,N_2804,N_2864);
or U2901 (N_2901,N_2818,N_2837);
nand U2902 (N_2902,N_2831,N_2895);
nand U2903 (N_2903,N_2825,N_2898);
xnor U2904 (N_2904,N_2886,N_2806);
or U2905 (N_2905,N_2815,N_2809);
and U2906 (N_2906,N_2810,N_2826);
xor U2907 (N_2907,N_2820,N_2840);
or U2908 (N_2908,N_2827,N_2888);
or U2909 (N_2909,N_2821,N_2861);
xnor U2910 (N_2910,N_2883,N_2893);
nor U2911 (N_2911,N_2882,N_2805);
xor U2912 (N_2912,N_2867,N_2808);
nand U2913 (N_2913,N_2892,N_2817);
or U2914 (N_2914,N_2858,N_2862);
xnor U2915 (N_2915,N_2803,N_2833);
nand U2916 (N_2916,N_2830,N_2842);
nand U2917 (N_2917,N_2807,N_2816);
or U2918 (N_2918,N_2839,N_2850);
or U2919 (N_2919,N_2896,N_2868);
and U2920 (N_2920,N_2894,N_2851);
and U2921 (N_2921,N_2800,N_2845);
nor U2922 (N_2922,N_2853,N_2802);
xor U2923 (N_2923,N_2865,N_2801);
nor U2924 (N_2924,N_2866,N_2875);
and U2925 (N_2925,N_2854,N_2874);
or U2926 (N_2926,N_2855,N_2856);
xor U2927 (N_2927,N_2860,N_2828);
xnor U2928 (N_2928,N_2843,N_2869);
nand U2929 (N_2929,N_2849,N_2872);
or U2930 (N_2930,N_2891,N_2873);
or U2931 (N_2931,N_2844,N_2835);
xor U2932 (N_2932,N_2863,N_2811);
nand U2933 (N_2933,N_2829,N_2857);
and U2934 (N_2934,N_2887,N_2848);
and U2935 (N_2935,N_2824,N_2871);
nor U2936 (N_2936,N_2876,N_2823);
or U2937 (N_2937,N_2881,N_2899);
xor U2938 (N_2938,N_2832,N_2814);
or U2939 (N_2939,N_2889,N_2846);
xnor U2940 (N_2940,N_2879,N_2834);
xnor U2941 (N_2941,N_2838,N_2847);
or U2942 (N_2942,N_2877,N_2880);
and U2943 (N_2943,N_2852,N_2859);
nand U2944 (N_2944,N_2897,N_2812);
nand U2945 (N_2945,N_2870,N_2884);
or U2946 (N_2946,N_2819,N_2890);
or U2947 (N_2947,N_2836,N_2822);
or U2948 (N_2948,N_2841,N_2878);
xor U2949 (N_2949,N_2813,N_2885);
and U2950 (N_2950,N_2884,N_2878);
and U2951 (N_2951,N_2830,N_2876);
nor U2952 (N_2952,N_2841,N_2893);
or U2953 (N_2953,N_2849,N_2832);
or U2954 (N_2954,N_2893,N_2875);
or U2955 (N_2955,N_2876,N_2851);
nor U2956 (N_2956,N_2843,N_2833);
nor U2957 (N_2957,N_2897,N_2860);
nor U2958 (N_2958,N_2862,N_2853);
or U2959 (N_2959,N_2885,N_2883);
nor U2960 (N_2960,N_2861,N_2837);
xor U2961 (N_2961,N_2854,N_2882);
xor U2962 (N_2962,N_2836,N_2826);
xor U2963 (N_2963,N_2894,N_2820);
and U2964 (N_2964,N_2807,N_2845);
xnor U2965 (N_2965,N_2861,N_2849);
nand U2966 (N_2966,N_2890,N_2879);
xnor U2967 (N_2967,N_2855,N_2872);
nand U2968 (N_2968,N_2886,N_2838);
nand U2969 (N_2969,N_2864,N_2863);
nor U2970 (N_2970,N_2801,N_2848);
nor U2971 (N_2971,N_2805,N_2880);
and U2972 (N_2972,N_2826,N_2818);
or U2973 (N_2973,N_2805,N_2872);
nand U2974 (N_2974,N_2884,N_2844);
and U2975 (N_2975,N_2824,N_2810);
xor U2976 (N_2976,N_2878,N_2868);
or U2977 (N_2977,N_2864,N_2894);
and U2978 (N_2978,N_2889,N_2858);
or U2979 (N_2979,N_2876,N_2818);
and U2980 (N_2980,N_2805,N_2852);
nand U2981 (N_2981,N_2882,N_2878);
xnor U2982 (N_2982,N_2848,N_2874);
or U2983 (N_2983,N_2826,N_2835);
nand U2984 (N_2984,N_2857,N_2815);
and U2985 (N_2985,N_2861,N_2840);
and U2986 (N_2986,N_2806,N_2855);
and U2987 (N_2987,N_2875,N_2819);
or U2988 (N_2988,N_2863,N_2810);
nand U2989 (N_2989,N_2871,N_2831);
xnor U2990 (N_2990,N_2830,N_2834);
nand U2991 (N_2991,N_2884,N_2865);
nand U2992 (N_2992,N_2849,N_2851);
and U2993 (N_2993,N_2894,N_2811);
nand U2994 (N_2994,N_2856,N_2802);
and U2995 (N_2995,N_2861,N_2801);
nor U2996 (N_2996,N_2817,N_2836);
xnor U2997 (N_2997,N_2882,N_2881);
nand U2998 (N_2998,N_2867,N_2892);
nor U2999 (N_2999,N_2802,N_2820);
nand U3000 (N_3000,N_2962,N_2997);
nand U3001 (N_3001,N_2958,N_2981);
xnor U3002 (N_3002,N_2956,N_2938);
nand U3003 (N_3003,N_2924,N_2954);
and U3004 (N_3004,N_2952,N_2967);
or U3005 (N_3005,N_2931,N_2932);
nand U3006 (N_3006,N_2984,N_2994);
xor U3007 (N_3007,N_2953,N_2901);
nor U3008 (N_3008,N_2908,N_2946);
xnor U3009 (N_3009,N_2966,N_2930);
and U3010 (N_3010,N_2927,N_2988);
or U3011 (N_3011,N_2940,N_2982);
nor U3012 (N_3012,N_2973,N_2942);
or U3013 (N_3013,N_2985,N_2974);
or U3014 (N_3014,N_2909,N_2920);
xnor U3015 (N_3015,N_2928,N_2949);
and U3016 (N_3016,N_2947,N_2975);
nand U3017 (N_3017,N_2943,N_2944);
xnor U3018 (N_3018,N_2979,N_2995);
nor U3019 (N_3019,N_2916,N_2963);
or U3020 (N_3020,N_2987,N_2903);
xnor U3021 (N_3021,N_2929,N_2964);
xor U3022 (N_3022,N_2961,N_2976);
nand U3023 (N_3023,N_2977,N_2934);
nor U3024 (N_3024,N_2915,N_2965);
and U3025 (N_3025,N_2918,N_2970);
nand U3026 (N_3026,N_2939,N_2980);
or U3027 (N_3027,N_2926,N_2936);
nand U3028 (N_3028,N_2941,N_2907);
nand U3029 (N_3029,N_2935,N_2950);
and U3030 (N_3030,N_2951,N_2992);
xor U3031 (N_3031,N_2968,N_2986);
or U3032 (N_3032,N_2913,N_2996);
nand U3033 (N_3033,N_2914,N_2969);
or U3034 (N_3034,N_2937,N_2978);
nand U3035 (N_3035,N_2960,N_2906);
nand U3036 (N_3036,N_2990,N_2972);
xnor U3037 (N_3037,N_2919,N_2991);
nor U3038 (N_3038,N_2999,N_2945);
nand U3039 (N_3039,N_2910,N_2948);
nor U3040 (N_3040,N_2921,N_2971);
xnor U3041 (N_3041,N_2993,N_2998);
nand U3042 (N_3042,N_2989,N_2925);
or U3043 (N_3043,N_2905,N_2957);
nand U3044 (N_3044,N_2922,N_2917);
xnor U3045 (N_3045,N_2912,N_2983);
or U3046 (N_3046,N_2904,N_2933);
xnor U3047 (N_3047,N_2900,N_2959);
and U3048 (N_3048,N_2902,N_2923);
xor U3049 (N_3049,N_2955,N_2911);
and U3050 (N_3050,N_2986,N_2904);
xnor U3051 (N_3051,N_2960,N_2993);
and U3052 (N_3052,N_2982,N_2961);
nand U3053 (N_3053,N_2964,N_2916);
or U3054 (N_3054,N_2903,N_2991);
nand U3055 (N_3055,N_2984,N_2918);
or U3056 (N_3056,N_2900,N_2940);
nor U3057 (N_3057,N_2949,N_2988);
and U3058 (N_3058,N_2928,N_2923);
nand U3059 (N_3059,N_2903,N_2959);
nor U3060 (N_3060,N_2939,N_2941);
and U3061 (N_3061,N_2930,N_2982);
and U3062 (N_3062,N_2972,N_2929);
and U3063 (N_3063,N_2924,N_2971);
nand U3064 (N_3064,N_2984,N_2976);
xnor U3065 (N_3065,N_2909,N_2976);
nor U3066 (N_3066,N_2965,N_2989);
and U3067 (N_3067,N_2943,N_2999);
xor U3068 (N_3068,N_2999,N_2965);
or U3069 (N_3069,N_2941,N_2959);
nand U3070 (N_3070,N_2961,N_2924);
xor U3071 (N_3071,N_2992,N_2995);
or U3072 (N_3072,N_2977,N_2960);
and U3073 (N_3073,N_2972,N_2960);
xor U3074 (N_3074,N_2933,N_2986);
nand U3075 (N_3075,N_2986,N_2997);
nor U3076 (N_3076,N_2936,N_2951);
nor U3077 (N_3077,N_2966,N_2997);
or U3078 (N_3078,N_2910,N_2986);
nand U3079 (N_3079,N_2946,N_2944);
nor U3080 (N_3080,N_2940,N_2996);
nor U3081 (N_3081,N_2925,N_2995);
or U3082 (N_3082,N_2967,N_2978);
nand U3083 (N_3083,N_2916,N_2997);
nor U3084 (N_3084,N_2975,N_2973);
nand U3085 (N_3085,N_2949,N_2932);
nor U3086 (N_3086,N_2978,N_2976);
or U3087 (N_3087,N_2930,N_2943);
nand U3088 (N_3088,N_2969,N_2947);
xor U3089 (N_3089,N_2907,N_2929);
or U3090 (N_3090,N_2985,N_2987);
and U3091 (N_3091,N_2903,N_2915);
nor U3092 (N_3092,N_2977,N_2961);
nor U3093 (N_3093,N_2924,N_2986);
nand U3094 (N_3094,N_2977,N_2952);
nor U3095 (N_3095,N_2920,N_2930);
and U3096 (N_3096,N_2908,N_2966);
nor U3097 (N_3097,N_2972,N_2925);
or U3098 (N_3098,N_2949,N_2923);
nand U3099 (N_3099,N_2923,N_2985);
or U3100 (N_3100,N_3047,N_3027);
nor U3101 (N_3101,N_3060,N_3075);
xor U3102 (N_3102,N_3070,N_3088);
xor U3103 (N_3103,N_3004,N_3041);
nand U3104 (N_3104,N_3044,N_3040);
nor U3105 (N_3105,N_3032,N_3092);
xnor U3106 (N_3106,N_3081,N_3013);
and U3107 (N_3107,N_3058,N_3091);
nand U3108 (N_3108,N_3076,N_3093);
and U3109 (N_3109,N_3063,N_3006);
xnor U3110 (N_3110,N_3024,N_3048);
nor U3111 (N_3111,N_3071,N_3034);
nand U3112 (N_3112,N_3085,N_3011);
xor U3113 (N_3113,N_3018,N_3078);
or U3114 (N_3114,N_3003,N_3072);
or U3115 (N_3115,N_3080,N_3001);
or U3116 (N_3116,N_3045,N_3019);
and U3117 (N_3117,N_3065,N_3056);
and U3118 (N_3118,N_3010,N_3069);
nand U3119 (N_3119,N_3079,N_3016);
nand U3120 (N_3120,N_3014,N_3054);
nor U3121 (N_3121,N_3096,N_3005);
or U3122 (N_3122,N_3067,N_3084);
nor U3123 (N_3123,N_3025,N_3002);
or U3124 (N_3124,N_3055,N_3009);
or U3125 (N_3125,N_3083,N_3026);
and U3126 (N_3126,N_3017,N_3061);
nand U3127 (N_3127,N_3066,N_3073);
and U3128 (N_3128,N_3049,N_3098);
xnor U3129 (N_3129,N_3007,N_3052);
and U3130 (N_3130,N_3042,N_3012);
nor U3131 (N_3131,N_3029,N_3022);
or U3132 (N_3132,N_3035,N_3000);
nor U3133 (N_3133,N_3008,N_3090);
xnor U3134 (N_3134,N_3033,N_3059);
nor U3135 (N_3135,N_3051,N_3015);
xnor U3136 (N_3136,N_3062,N_3089);
nor U3137 (N_3137,N_3057,N_3031);
or U3138 (N_3138,N_3039,N_3097);
and U3139 (N_3139,N_3020,N_3082);
nor U3140 (N_3140,N_3021,N_3074);
nand U3141 (N_3141,N_3068,N_3095);
nand U3142 (N_3142,N_3037,N_3030);
xor U3143 (N_3143,N_3046,N_3086);
nor U3144 (N_3144,N_3064,N_3053);
or U3145 (N_3145,N_3023,N_3036);
xor U3146 (N_3146,N_3050,N_3043);
and U3147 (N_3147,N_3077,N_3038);
or U3148 (N_3148,N_3087,N_3099);
xor U3149 (N_3149,N_3094,N_3028);
xnor U3150 (N_3150,N_3082,N_3054);
nor U3151 (N_3151,N_3059,N_3040);
and U3152 (N_3152,N_3053,N_3019);
nor U3153 (N_3153,N_3069,N_3079);
or U3154 (N_3154,N_3061,N_3063);
or U3155 (N_3155,N_3052,N_3048);
and U3156 (N_3156,N_3098,N_3031);
nor U3157 (N_3157,N_3019,N_3005);
nor U3158 (N_3158,N_3092,N_3080);
and U3159 (N_3159,N_3093,N_3042);
nand U3160 (N_3160,N_3021,N_3016);
and U3161 (N_3161,N_3022,N_3056);
and U3162 (N_3162,N_3010,N_3027);
and U3163 (N_3163,N_3026,N_3064);
nor U3164 (N_3164,N_3042,N_3094);
nor U3165 (N_3165,N_3052,N_3030);
xor U3166 (N_3166,N_3017,N_3077);
nor U3167 (N_3167,N_3095,N_3008);
xnor U3168 (N_3168,N_3074,N_3022);
and U3169 (N_3169,N_3036,N_3038);
or U3170 (N_3170,N_3056,N_3058);
nand U3171 (N_3171,N_3059,N_3009);
xor U3172 (N_3172,N_3077,N_3014);
and U3173 (N_3173,N_3001,N_3002);
xor U3174 (N_3174,N_3035,N_3082);
or U3175 (N_3175,N_3060,N_3064);
and U3176 (N_3176,N_3038,N_3000);
xor U3177 (N_3177,N_3089,N_3064);
or U3178 (N_3178,N_3037,N_3057);
nand U3179 (N_3179,N_3043,N_3075);
xor U3180 (N_3180,N_3076,N_3061);
or U3181 (N_3181,N_3028,N_3079);
or U3182 (N_3182,N_3029,N_3021);
and U3183 (N_3183,N_3094,N_3083);
nand U3184 (N_3184,N_3092,N_3095);
or U3185 (N_3185,N_3083,N_3095);
or U3186 (N_3186,N_3049,N_3008);
and U3187 (N_3187,N_3097,N_3092);
or U3188 (N_3188,N_3076,N_3023);
and U3189 (N_3189,N_3036,N_3098);
nand U3190 (N_3190,N_3020,N_3033);
and U3191 (N_3191,N_3091,N_3037);
nor U3192 (N_3192,N_3033,N_3089);
xnor U3193 (N_3193,N_3055,N_3020);
nand U3194 (N_3194,N_3031,N_3012);
nand U3195 (N_3195,N_3037,N_3019);
nor U3196 (N_3196,N_3087,N_3091);
nor U3197 (N_3197,N_3032,N_3095);
xnor U3198 (N_3198,N_3005,N_3033);
xor U3199 (N_3199,N_3006,N_3053);
xnor U3200 (N_3200,N_3185,N_3175);
or U3201 (N_3201,N_3193,N_3125);
nor U3202 (N_3202,N_3171,N_3134);
and U3203 (N_3203,N_3168,N_3157);
nand U3204 (N_3204,N_3174,N_3187);
nor U3205 (N_3205,N_3121,N_3137);
or U3206 (N_3206,N_3128,N_3176);
nor U3207 (N_3207,N_3135,N_3144);
nor U3208 (N_3208,N_3199,N_3173);
xor U3209 (N_3209,N_3129,N_3120);
xor U3210 (N_3210,N_3126,N_3180);
or U3211 (N_3211,N_3118,N_3136);
or U3212 (N_3212,N_3159,N_3172);
nor U3213 (N_3213,N_3196,N_3177);
nand U3214 (N_3214,N_3104,N_3114);
or U3215 (N_3215,N_3167,N_3113);
xnor U3216 (N_3216,N_3111,N_3191);
nor U3217 (N_3217,N_3169,N_3183);
nand U3218 (N_3218,N_3101,N_3141);
nor U3219 (N_3219,N_3102,N_3153);
xor U3220 (N_3220,N_3146,N_3194);
nor U3221 (N_3221,N_3189,N_3116);
nand U3222 (N_3222,N_3163,N_3103);
nor U3223 (N_3223,N_3123,N_3149);
nand U3224 (N_3224,N_3127,N_3112);
nor U3225 (N_3225,N_3148,N_3162);
or U3226 (N_3226,N_3117,N_3186);
xor U3227 (N_3227,N_3122,N_3179);
xor U3228 (N_3228,N_3198,N_3119);
nand U3229 (N_3229,N_3166,N_3115);
nor U3230 (N_3230,N_3152,N_3161);
or U3231 (N_3231,N_3158,N_3156);
nand U3232 (N_3232,N_3107,N_3155);
and U3233 (N_3233,N_3145,N_3154);
nor U3234 (N_3234,N_3108,N_3150);
nand U3235 (N_3235,N_3109,N_3106);
nor U3236 (N_3236,N_3138,N_3100);
and U3237 (N_3237,N_3110,N_3140);
and U3238 (N_3238,N_3143,N_3188);
nor U3239 (N_3239,N_3124,N_3130);
xor U3240 (N_3240,N_3197,N_3178);
xnor U3241 (N_3241,N_3105,N_3195);
nor U3242 (N_3242,N_3131,N_3192);
nand U3243 (N_3243,N_3160,N_3165);
nor U3244 (N_3244,N_3151,N_3147);
nand U3245 (N_3245,N_3139,N_3170);
nand U3246 (N_3246,N_3142,N_3182);
nand U3247 (N_3247,N_3184,N_3190);
nor U3248 (N_3248,N_3133,N_3164);
nor U3249 (N_3249,N_3132,N_3181);
xor U3250 (N_3250,N_3179,N_3116);
nor U3251 (N_3251,N_3178,N_3174);
or U3252 (N_3252,N_3109,N_3146);
xor U3253 (N_3253,N_3148,N_3183);
nand U3254 (N_3254,N_3144,N_3119);
and U3255 (N_3255,N_3175,N_3100);
nand U3256 (N_3256,N_3116,N_3110);
xor U3257 (N_3257,N_3188,N_3141);
and U3258 (N_3258,N_3168,N_3186);
or U3259 (N_3259,N_3171,N_3141);
and U3260 (N_3260,N_3199,N_3132);
xnor U3261 (N_3261,N_3128,N_3195);
or U3262 (N_3262,N_3176,N_3124);
nand U3263 (N_3263,N_3141,N_3103);
xnor U3264 (N_3264,N_3168,N_3183);
and U3265 (N_3265,N_3138,N_3103);
nand U3266 (N_3266,N_3133,N_3182);
xor U3267 (N_3267,N_3101,N_3116);
xor U3268 (N_3268,N_3168,N_3176);
xor U3269 (N_3269,N_3147,N_3100);
xor U3270 (N_3270,N_3174,N_3145);
and U3271 (N_3271,N_3101,N_3140);
or U3272 (N_3272,N_3167,N_3140);
and U3273 (N_3273,N_3106,N_3198);
xnor U3274 (N_3274,N_3177,N_3161);
and U3275 (N_3275,N_3154,N_3156);
or U3276 (N_3276,N_3109,N_3137);
nand U3277 (N_3277,N_3140,N_3104);
or U3278 (N_3278,N_3156,N_3114);
xnor U3279 (N_3279,N_3126,N_3131);
nor U3280 (N_3280,N_3148,N_3126);
nand U3281 (N_3281,N_3174,N_3164);
nand U3282 (N_3282,N_3171,N_3126);
nand U3283 (N_3283,N_3177,N_3142);
nand U3284 (N_3284,N_3141,N_3115);
and U3285 (N_3285,N_3191,N_3112);
or U3286 (N_3286,N_3113,N_3174);
xor U3287 (N_3287,N_3131,N_3164);
and U3288 (N_3288,N_3174,N_3182);
and U3289 (N_3289,N_3158,N_3176);
nand U3290 (N_3290,N_3106,N_3149);
nand U3291 (N_3291,N_3153,N_3118);
and U3292 (N_3292,N_3135,N_3149);
nor U3293 (N_3293,N_3154,N_3199);
or U3294 (N_3294,N_3168,N_3143);
xor U3295 (N_3295,N_3115,N_3193);
or U3296 (N_3296,N_3106,N_3174);
and U3297 (N_3297,N_3127,N_3143);
and U3298 (N_3298,N_3113,N_3180);
nand U3299 (N_3299,N_3152,N_3101);
and U3300 (N_3300,N_3247,N_3263);
and U3301 (N_3301,N_3218,N_3257);
and U3302 (N_3302,N_3254,N_3238);
xor U3303 (N_3303,N_3214,N_3204);
nor U3304 (N_3304,N_3273,N_3241);
or U3305 (N_3305,N_3283,N_3271);
nor U3306 (N_3306,N_3223,N_3219);
nor U3307 (N_3307,N_3256,N_3230);
nand U3308 (N_3308,N_3226,N_3262);
nor U3309 (N_3309,N_3279,N_3258);
xnor U3310 (N_3310,N_3253,N_3291);
nand U3311 (N_3311,N_3286,N_3239);
nor U3312 (N_3312,N_3267,N_3295);
and U3313 (N_3313,N_3250,N_3270);
nand U3314 (N_3314,N_3206,N_3281);
and U3315 (N_3315,N_3287,N_3231);
or U3316 (N_3316,N_3248,N_3213);
nor U3317 (N_3317,N_3201,N_3289);
nor U3318 (N_3318,N_3245,N_3294);
and U3319 (N_3319,N_3210,N_3233);
or U3320 (N_3320,N_3275,N_3229);
nand U3321 (N_3321,N_3212,N_3269);
xor U3322 (N_3322,N_3278,N_3202);
nor U3323 (N_3323,N_3246,N_3298);
xnor U3324 (N_3324,N_3243,N_3222);
nand U3325 (N_3325,N_3293,N_3224);
xnor U3326 (N_3326,N_3288,N_3216);
nand U3327 (N_3327,N_3274,N_3217);
xnor U3328 (N_3328,N_3205,N_3252);
nor U3329 (N_3329,N_3236,N_3285);
nand U3330 (N_3330,N_3259,N_3215);
or U3331 (N_3331,N_3272,N_3284);
nand U3332 (N_3332,N_3297,N_3249);
and U3333 (N_3333,N_3266,N_3232);
or U3334 (N_3334,N_3235,N_3220);
xor U3335 (N_3335,N_3234,N_3208);
xnor U3336 (N_3336,N_3261,N_3207);
xor U3337 (N_3337,N_3240,N_3251);
nor U3338 (N_3338,N_3296,N_3264);
xor U3339 (N_3339,N_3228,N_3237);
or U3340 (N_3340,N_3225,N_3244);
xnor U3341 (N_3341,N_3277,N_3280);
nor U3342 (N_3342,N_3299,N_3200);
or U3343 (N_3343,N_3242,N_3260);
xnor U3344 (N_3344,N_3209,N_3265);
nand U3345 (N_3345,N_3227,N_3292);
nor U3346 (N_3346,N_3203,N_3268);
and U3347 (N_3347,N_3290,N_3282);
or U3348 (N_3348,N_3211,N_3221);
nand U3349 (N_3349,N_3276,N_3255);
and U3350 (N_3350,N_3236,N_3228);
and U3351 (N_3351,N_3229,N_3201);
nand U3352 (N_3352,N_3278,N_3213);
xnor U3353 (N_3353,N_3241,N_3213);
or U3354 (N_3354,N_3268,N_3221);
nor U3355 (N_3355,N_3268,N_3235);
nor U3356 (N_3356,N_3267,N_3217);
nor U3357 (N_3357,N_3297,N_3214);
and U3358 (N_3358,N_3204,N_3265);
and U3359 (N_3359,N_3213,N_3290);
xnor U3360 (N_3360,N_3233,N_3222);
nand U3361 (N_3361,N_3262,N_3280);
xnor U3362 (N_3362,N_3241,N_3282);
nor U3363 (N_3363,N_3224,N_3279);
nand U3364 (N_3364,N_3217,N_3210);
nand U3365 (N_3365,N_3217,N_3298);
or U3366 (N_3366,N_3207,N_3294);
xnor U3367 (N_3367,N_3224,N_3214);
and U3368 (N_3368,N_3204,N_3226);
xor U3369 (N_3369,N_3254,N_3261);
nand U3370 (N_3370,N_3256,N_3298);
or U3371 (N_3371,N_3215,N_3249);
xor U3372 (N_3372,N_3204,N_3224);
nor U3373 (N_3373,N_3262,N_3245);
nor U3374 (N_3374,N_3291,N_3241);
or U3375 (N_3375,N_3231,N_3259);
xor U3376 (N_3376,N_3285,N_3214);
or U3377 (N_3377,N_3240,N_3266);
nand U3378 (N_3378,N_3207,N_3292);
and U3379 (N_3379,N_3258,N_3251);
nand U3380 (N_3380,N_3251,N_3248);
nand U3381 (N_3381,N_3262,N_3274);
nor U3382 (N_3382,N_3243,N_3234);
nor U3383 (N_3383,N_3228,N_3205);
nand U3384 (N_3384,N_3201,N_3255);
nor U3385 (N_3385,N_3249,N_3208);
or U3386 (N_3386,N_3279,N_3298);
or U3387 (N_3387,N_3245,N_3297);
nor U3388 (N_3388,N_3258,N_3291);
and U3389 (N_3389,N_3227,N_3241);
xnor U3390 (N_3390,N_3225,N_3295);
nor U3391 (N_3391,N_3273,N_3201);
or U3392 (N_3392,N_3274,N_3200);
xor U3393 (N_3393,N_3282,N_3269);
or U3394 (N_3394,N_3221,N_3277);
nand U3395 (N_3395,N_3255,N_3272);
or U3396 (N_3396,N_3266,N_3219);
nand U3397 (N_3397,N_3250,N_3291);
or U3398 (N_3398,N_3216,N_3237);
xnor U3399 (N_3399,N_3290,N_3269);
nand U3400 (N_3400,N_3307,N_3370);
and U3401 (N_3401,N_3340,N_3315);
or U3402 (N_3402,N_3365,N_3376);
nand U3403 (N_3403,N_3361,N_3325);
or U3404 (N_3404,N_3367,N_3318);
xor U3405 (N_3405,N_3372,N_3396);
or U3406 (N_3406,N_3322,N_3369);
xor U3407 (N_3407,N_3314,N_3366);
or U3408 (N_3408,N_3323,N_3398);
xnor U3409 (N_3409,N_3304,N_3341);
nand U3410 (N_3410,N_3364,N_3309);
nor U3411 (N_3411,N_3379,N_3339);
nor U3412 (N_3412,N_3329,N_3332);
xnor U3413 (N_3413,N_3395,N_3333);
xnor U3414 (N_3414,N_3359,N_3338);
or U3415 (N_3415,N_3321,N_3399);
xor U3416 (N_3416,N_3382,N_3373);
or U3417 (N_3417,N_3397,N_3319);
or U3418 (N_3418,N_3383,N_3362);
nand U3419 (N_3419,N_3316,N_3393);
xnor U3420 (N_3420,N_3326,N_3378);
nor U3421 (N_3421,N_3375,N_3353);
nand U3422 (N_3422,N_3301,N_3380);
nand U3423 (N_3423,N_3337,N_3391);
and U3424 (N_3424,N_3368,N_3328);
xor U3425 (N_3425,N_3355,N_3346);
nand U3426 (N_3426,N_3331,N_3352);
nor U3427 (N_3427,N_3303,N_3312);
xor U3428 (N_3428,N_3343,N_3351);
nor U3429 (N_3429,N_3381,N_3363);
xnor U3430 (N_3430,N_3344,N_3308);
or U3431 (N_3431,N_3349,N_3358);
nor U3432 (N_3432,N_3345,N_3348);
and U3433 (N_3433,N_3377,N_3310);
and U3434 (N_3434,N_3330,N_3387);
nor U3435 (N_3435,N_3357,N_3335);
and U3436 (N_3436,N_3390,N_3354);
and U3437 (N_3437,N_3384,N_3374);
nand U3438 (N_3438,N_3305,N_3371);
xnor U3439 (N_3439,N_3360,N_3302);
or U3440 (N_3440,N_3306,N_3356);
and U3441 (N_3441,N_3385,N_3386);
xnor U3442 (N_3442,N_3342,N_3320);
or U3443 (N_3443,N_3347,N_3389);
and U3444 (N_3444,N_3336,N_3317);
nand U3445 (N_3445,N_3324,N_3300);
nand U3446 (N_3446,N_3311,N_3334);
nor U3447 (N_3447,N_3327,N_3350);
nand U3448 (N_3448,N_3392,N_3388);
nand U3449 (N_3449,N_3394,N_3313);
or U3450 (N_3450,N_3392,N_3359);
xor U3451 (N_3451,N_3353,N_3360);
xor U3452 (N_3452,N_3304,N_3340);
nor U3453 (N_3453,N_3375,N_3328);
and U3454 (N_3454,N_3365,N_3318);
xor U3455 (N_3455,N_3370,N_3387);
and U3456 (N_3456,N_3338,N_3370);
or U3457 (N_3457,N_3386,N_3360);
nor U3458 (N_3458,N_3357,N_3364);
nor U3459 (N_3459,N_3305,N_3397);
nand U3460 (N_3460,N_3381,N_3351);
nor U3461 (N_3461,N_3317,N_3301);
nor U3462 (N_3462,N_3332,N_3330);
and U3463 (N_3463,N_3383,N_3315);
nand U3464 (N_3464,N_3361,N_3309);
and U3465 (N_3465,N_3334,N_3364);
xnor U3466 (N_3466,N_3337,N_3371);
xnor U3467 (N_3467,N_3302,N_3383);
and U3468 (N_3468,N_3329,N_3353);
xor U3469 (N_3469,N_3360,N_3319);
nor U3470 (N_3470,N_3342,N_3328);
nor U3471 (N_3471,N_3301,N_3314);
and U3472 (N_3472,N_3367,N_3385);
nand U3473 (N_3473,N_3328,N_3301);
xor U3474 (N_3474,N_3368,N_3341);
or U3475 (N_3475,N_3324,N_3304);
nand U3476 (N_3476,N_3364,N_3388);
nand U3477 (N_3477,N_3399,N_3371);
nor U3478 (N_3478,N_3332,N_3346);
and U3479 (N_3479,N_3349,N_3398);
or U3480 (N_3480,N_3395,N_3352);
nand U3481 (N_3481,N_3345,N_3352);
nand U3482 (N_3482,N_3370,N_3337);
or U3483 (N_3483,N_3303,N_3397);
nand U3484 (N_3484,N_3376,N_3319);
nand U3485 (N_3485,N_3398,N_3319);
or U3486 (N_3486,N_3371,N_3379);
and U3487 (N_3487,N_3370,N_3363);
nand U3488 (N_3488,N_3383,N_3374);
nand U3489 (N_3489,N_3384,N_3395);
or U3490 (N_3490,N_3369,N_3386);
or U3491 (N_3491,N_3359,N_3331);
nand U3492 (N_3492,N_3352,N_3334);
nand U3493 (N_3493,N_3396,N_3338);
or U3494 (N_3494,N_3359,N_3379);
nor U3495 (N_3495,N_3374,N_3303);
xor U3496 (N_3496,N_3320,N_3302);
nor U3497 (N_3497,N_3351,N_3368);
nand U3498 (N_3498,N_3357,N_3391);
nand U3499 (N_3499,N_3340,N_3320);
or U3500 (N_3500,N_3484,N_3463);
and U3501 (N_3501,N_3481,N_3419);
nand U3502 (N_3502,N_3451,N_3425);
and U3503 (N_3503,N_3498,N_3466);
or U3504 (N_3504,N_3444,N_3421);
xnor U3505 (N_3505,N_3438,N_3439);
nor U3506 (N_3506,N_3448,N_3487);
nand U3507 (N_3507,N_3476,N_3437);
and U3508 (N_3508,N_3482,N_3488);
or U3509 (N_3509,N_3456,N_3489);
nor U3510 (N_3510,N_3415,N_3493);
nor U3511 (N_3511,N_3426,N_3467);
and U3512 (N_3512,N_3433,N_3441);
or U3513 (N_3513,N_3452,N_3409);
or U3514 (N_3514,N_3461,N_3442);
and U3515 (N_3515,N_3420,N_3462);
and U3516 (N_3516,N_3400,N_3492);
nand U3517 (N_3517,N_3403,N_3464);
and U3518 (N_3518,N_3423,N_3470);
nor U3519 (N_3519,N_3401,N_3480);
and U3520 (N_3520,N_3486,N_3471);
nor U3521 (N_3521,N_3496,N_3499);
nor U3522 (N_3522,N_3405,N_3474);
nand U3523 (N_3523,N_3413,N_3424);
xor U3524 (N_3524,N_3434,N_3477);
or U3525 (N_3525,N_3436,N_3495);
or U3526 (N_3526,N_3485,N_3478);
or U3527 (N_3527,N_3427,N_3490);
or U3528 (N_3528,N_3410,N_3475);
nor U3529 (N_3529,N_3491,N_3402);
nor U3530 (N_3530,N_3449,N_3472);
nor U3531 (N_3531,N_3411,N_3430);
nor U3532 (N_3532,N_3458,N_3422);
nand U3533 (N_3533,N_3408,N_3404);
or U3534 (N_3534,N_3497,N_3455);
xnor U3535 (N_3535,N_3406,N_3407);
xnor U3536 (N_3536,N_3445,N_3428);
and U3537 (N_3537,N_3460,N_3435);
xor U3538 (N_3538,N_3440,N_3473);
and U3539 (N_3539,N_3417,N_3465);
nand U3540 (N_3540,N_3446,N_3414);
nand U3541 (N_3541,N_3479,N_3447);
nor U3542 (N_3542,N_3469,N_3412);
and U3543 (N_3543,N_3418,N_3494);
xnor U3544 (N_3544,N_3429,N_3454);
nand U3545 (N_3545,N_3443,N_3453);
and U3546 (N_3546,N_3483,N_3431);
nand U3547 (N_3547,N_3450,N_3416);
and U3548 (N_3548,N_3432,N_3457);
nand U3549 (N_3549,N_3468,N_3459);
or U3550 (N_3550,N_3415,N_3419);
and U3551 (N_3551,N_3473,N_3496);
or U3552 (N_3552,N_3420,N_3447);
nand U3553 (N_3553,N_3430,N_3416);
and U3554 (N_3554,N_3487,N_3488);
and U3555 (N_3555,N_3451,N_3463);
xor U3556 (N_3556,N_3486,N_3401);
nand U3557 (N_3557,N_3415,N_3441);
nand U3558 (N_3558,N_3437,N_3483);
nand U3559 (N_3559,N_3449,N_3454);
and U3560 (N_3560,N_3486,N_3414);
and U3561 (N_3561,N_3482,N_3445);
nand U3562 (N_3562,N_3458,N_3460);
or U3563 (N_3563,N_3482,N_3401);
or U3564 (N_3564,N_3433,N_3458);
xnor U3565 (N_3565,N_3492,N_3450);
nor U3566 (N_3566,N_3409,N_3446);
and U3567 (N_3567,N_3472,N_3454);
or U3568 (N_3568,N_3421,N_3476);
and U3569 (N_3569,N_3471,N_3420);
or U3570 (N_3570,N_3445,N_3458);
and U3571 (N_3571,N_3468,N_3489);
or U3572 (N_3572,N_3429,N_3433);
or U3573 (N_3573,N_3492,N_3475);
and U3574 (N_3574,N_3490,N_3424);
or U3575 (N_3575,N_3440,N_3424);
nand U3576 (N_3576,N_3491,N_3431);
xor U3577 (N_3577,N_3453,N_3479);
or U3578 (N_3578,N_3409,N_3480);
nand U3579 (N_3579,N_3479,N_3441);
nor U3580 (N_3580,N_3419,N_3456);
nand U3581 (N_3581,N_3420,N_3494);
or U3582 (N_3582,N_3461,N_3469);
and U3583 (N_3583,N_3477,N_3430);
nor U3584 (N_3584,N_3476,N_3403);
or U3585 (N_3585,N_3429,N_3496);
nor U3586 (N_3586,N_3446,N_3413);
nand U3587 (N_3587,N_3493,N_3446);
nor U3588 (N_3588,N_3496,N_3408);
or U3589 (N_3589,N_3461,N_3488);
nor U3590 (N_3590,N_3438,N_3413);
and U3591 (N_3591,N_3481,N_3487);
nor U3592 (N_3592,N_3471,N_3460);
and U3593 (N_3593,N_3401,N_3468);
or U3594 (N_3594,N_3472,N_3405);
and U3595 (N_3595,N_3415,N_3431);
xnor U3596 (N_3596,N_3466,N_3438);
xnor U3597 (N_3597,N_3488,N_3420);
nor U3598 (N_3598,N_3459,N_3487);
and U3599 (N_3599,N_3411,N_3443);
nor U3600 (N_3600,N_3596,N_3558);
nor U3601 (N_3601,N_3525,N_3598);
nor U3602 (N_3602,N_3576,N_3562);
nand U3603 (N_3603,N_3566,N_3555);
nand U3604 (N_3604,N_3531,N_3585);
xor U3605 (N_3605,N_3586,N_3565);
xor U3606 (N_3606,N_3571,N_3503);
xor U3607 (N_3607,N_3504,N_3538);
or U3608 (N_3608,N_3501,N_3550);
and U3609 (N_3609,N_3595,N_3528);
xnor U3610 (N_3610,N_3588,N_3563);
and U3611 (N_3611,N_3579,N_3578);
xnor U3612 (N_3612,N_3582,N_3583);
or U3613 (N_3613,N_3553,N_3592);
xor U3614 (N_3614,N_3509,N_3544);
or U3615 (N_3615,N_3541,N_3518);
nand U3616 (N_3616,N_3536,N_3526);
or U3617 (N_3617,N_3546,N_3514);
xor U3618 (N_3618,N_3505,N_3527);
and U3619 (N_3619,N_3569,N_3534);
or U3620 (N_3620,N_3512,N_3519);
nand U3621 (N_3621,N_3502,N_3577);
and U3622 (N_3622,N_3572,N_3516);
xor U3623 (N_3623,N_3521,N_3549);
xor U3624 (N_3624,N_3581,N_3552);
or U3625 (N_3625,N_3575,N_3533);
and U3626 (N_3626,N_3537,N_3593);
or U3627 (N_3627,N_3591,N_3564);
and U3628 (N_3628,N_3517,N_3590);
nand U3629 (N_3629,N_3589,N_3530);
and U3630 (N_3630,N_3510,N_3507);
and U3631 (N_3631,N_3548,N_3597);
xor U3632 (N_3632,N_3570,N_3567);
nor U3633 (N_3633,N_3543,N_3554);
nand U3634 (N_3634,N_3511,N_3539);
xnor U3635 (N_3635,N_3557,N_3559);
and U3636 (N_3636,N_3535,N_3532);
nand U3637 (N_3637,N_3500,N_3513);
and U3638 (N_3638,N_3515,N_3580);
nand U3639 (N_3639,N_3542,N_3584);
nand U3640 (N_3640,N_3560,N_3573);
or U3641 (N_3641,N_3574,N_3587);
nor U3642 (N_3642,N_3545,N_3523);
xnor U3643 (N_3643,N_3599,N_3568);
and U3644 (N_3644,N_3508,N_3529);
nand U3645 (N_3645,N_3540,N_3522);
nand U3646 (N_3646,N_3561,N_3547);
nor U3647 (N_3647,N_3520,N_3556);
nor U3648 (N_3648,N_3506,N_3551);
xnor U3649 (N_3649,N_3594,N_3524);
or U3650 (N_3650,N_3591,N_3593);
nand U3651 (N_3651,N_3561,N_3546);
or U3652 (N_3652,N_3503,N_3504);
nor U3653 (N_3653,N_3558,N_3568);
and U3654 (N_3654,N_3544,N_3595);
and U3655 (N_3655,N_3532,N_3565);
nand U3656 (N_3656,N_3506,N_3552);
nand U3657 (N_3657,N_3565,N_3559);
or U3658 (N_3658,N_3558,N_3563);
or U3659 (N_3659,N_3516,N_3507);
and U3660 (N_3660,N_3595,N_3593);
and U3661 (N_3661,N_3536,N_3566);
xor U3662 (N_3662,N_3522,N_3587);
or U3663 (N_3663,N_3586,N_3551);
nand U3664 (N_3664,N_3560,N_3574);
nand U3665 (N_3665,N_3555,N_3592);
and U3666 (N_3666,N_3585,N_3599);
and U3667 (N_3667,N_3544,N_3505);
xor U3668 (N_3668,N_3532,N_3587);
and U3669 (N_3669,N_3562,N_3525);
nor U3670 (N_3670,N_3566,N_3598);
or U3671 (N_3671,N_3548,N_3593);
or U3672 (N_3672,N_3572,N_3560);
nand U3673 (N_3673,N_3545,N_3526);
nand U3674 (N_3674,N_3561,N_3584);
nand U3675 (N_3675,N_3515,N_3582);
and U3676 (N_3676,N_3562,N_3539);
xor U3677 (N_3677,N_3512,N_3598);
and U3678 (N_3678,N_3574,N_3514);
or U3679 (N_3679,N_3566,N_3510);
and U3680 (N_3680,N_3524,N_3558);
and U3681 (N_3681,N_3579,N_3519);
or U3682 (N_3682,N_3582,N_3558);
xnor U3683 (N_3683,N_3564,N_3578);
xor U3684 (N_3684,N_3547,N_3502);
nand U3685 (N_3685,N_3554,N_3544);
xnor U3686 (N_3686,N_3521,N_3591);
and U3687 (N_3687,N_3599,N_3519);
and U3688 (N_3688,N_3551,N_3524);
nor U3689 (N_3689,N_3565,N_3599);
xor U3690 (N_3690,N_3571,N_3540);
xor U3691 (N_3691,N_3531,N_3598);
nor U3692 (N_3692,N_3548,N_3591);
and U3693 (N_3693,N_3558,N_3538);
nor U3694 (N_3694,N_3579,N_3535);
xnor U3695 (N_3695,N_3505,N_3543);
and U3696 (N_3696,N_3500,N_3592);
nand U3697 (N_3697,N_3503,N_3566);
xor U3698 (N_3698,N_3563,N_3525);
nor U3699 (N_3699,N_3554,N_3588);
or U3700 (N_3700,N_3626,N_3650);
and U3701 (N_3701,N_3663,N_3619);
nor U3702 (N_3702,N_3644,N_3677);
nor U3703 (N_3703,N_3652,N_3634);
or U3704 (N_3704,N_3602,N_3675);
nor U3705 (N_3705,N_3670,N_3686);
and U3706 (N_3706,N_3654,N_3638);
xor U3707 (N_3707,N_3660,N_3695);
nand U3708 (N_3708,N_3694,N_3601);
or U3709 (N_3709,N_3631,N_3621);
nand U3710 (N_3710,N_3699,N_3646);
and U3711 (N_3711,N_3680,N_3698);
nor U3712 (N_3712,N_3679,N_3666);
nor U3713 (N_3713,N_3653,N_3665);
xnor U3714 (N_3714,N_3639,N_3618);
nor U3715 (N_3715,N_3625,N_3640);
and U3716 (N_3716,N_3692,N_3689);
xor U3717 (N_3717,N_3608,N_3629);
xor U3718 (N_3718,N_3648,N_3684);
nand U3719 (N_3719,N_3649,N_3678);
and U3720 (N_3720,N_3614,N_3656);
nand U3721 (N_3721,N_3668,N_3672);
xnor U3722 (N_3722,N_3633,N_3685);
xnor U3723 (N_3723,N_3661,N_3682);
and U3724 (N_3724,N_3647,N_3613);
nand U3725 (N_3725,N_3662,N_3683);
or U3726 (N_3726,N_3604,N_3645);
or U3727 (N_3727,N_3687,N_3671);
nand U3728 (N_3728,N_3655,N_3659);
and U3729 (N_3729,N_3632,N_3658);
or U3730 (N_3730,N_3615,N_3643);
or U3731 (N_3731,N_3669,N_3697);
or U3732 (N_3732,N_3630,N_3622);
or U3733 (N_3733,N_3620,N_3623);
xor U3734 (N_3734,N_3657,N_3603);
or U3735 (N_3735,N_3624,N_3693);
nand U3736 (N_3736,N_3600,N_3607);
nand U3737 (N_3737,N_3636,N_3606);
xnor U3738 (N_3738,N_3673,N_3651);
or U3739 (N_3739,N_3605,N_3690);
nand U3740 (N_3740,N_3691,N_3612);
or U3741 (N_3741,N_3609,N_3627);
xnor U3742 (N_3742,N_3635,N_3696);
and U3743 (N_3743,N_3676,N_3617);
nor U3744 (N_3744,N_3616,N_3641);
xnor U3745 (N_3745,N_3688,N_3611);
nand U3746 (N_3746,N_3637,N_3681);
and U3747 (N_3747,N_3674,N_3610);
and U3748 (N_3748,N_3642,N_3664);
or U3749 (N_3749,N_3667,N_3628);
nand U3750 (N_3750,N_3601,N_3642);
and U3751 (N_3751,N_3644,N_3655);
nand U3752 (N_3752,N_3674,N_3642);
and U3753 (N_3753,N_3699,N_3695);
nand U3754 (N_3754,N_3673,N_3637);
xor U3755 (N_3755,N_3661,N_3640);
and U3756 (N_3756,N_3658,N_3667);
nand U3757 (N_3757,N_3600,N_3613);
or U3758 (N_3758,N_3603,N_3604);
nor U3759 (N_3759,N_3657,N_3611);
xor U3760 (N_3760,N_3657,N_3623);
and U3761 (N_3761,N_3643,N_3606);
and U3762 (N_3762,N_3601,N_3635);
nand U3763 (N_3763,N_3666,N_3665);
or U3764 (N_3764,N_3688,N_3667);
nor U3765 (N_3765,N_3688,N_3699);
nor U3766 (N_3766,N_3653,N_3657);
nand U3767 (N_3767,N_3652,N_3654);
nor U3768 (N_3768,N_3638,N_3693);
nand U3769 (N_3769,N_3613,N_3652);
nand U3770 (N_3770,N_3608,N_3634);
nand U3771 (N_3771,N_3685,N_3686);
or U3772 (N_3772,N_3609,N_3636);
or U3773 (N_3773,N_3637,N_3674);
and U3774 (N_3774,N_3655,N_3611);
and U3775 (N_3775,N_3652,N_3678);
xor U3776 (N_3776,N_3636,N_3661);
nand U3777 (N_3777,N_3610,N_3695);
and U3778 (N_3778,N_3691,N_3654);
and U3779 (N_3779,N_3629,N_3604);
xor U3780 (N_3780,N_3690,N_3649);
nor U3781 (N_3781,N_3639,N_3692);
nand U3782 (N_3782,N_3676,N_3608);
xnor U3783 (N_3783,N_3611,N_3607);
xnor U3784 (N_3784,N_3671,N_3611);
nand U3785 (N_3785,N_3650,N_3616);
xor U3786 (N_3786,N_3658,N_3697);
or U3787 (N_3787,N_3665,N_3672);
nand U3788 (N_3788,N_3626,N_3634);
and U3789 (N_3789,N_3697,N_3663);
nor U3790 (N_3790,N_3662,N_3690);
or U3791 (N_3791,N_3625,N_3683);
and U3792 (N_3792,N_3671,N_3684);
and U3793 (N_3793,N_3691,N_3670);
nand U3794 (N_3794,N_3660,N_3624);
and U3795 (N_3795,N_3601,N_3627);
nor U3796 (N_3796,N_3674,N_3666);
and U3797 (N_3797,N_3679,N_3633);
or U3798 (N_3798,N_3630,N_3671);
or U3799 (N_3799,N_3606,N_3612);
nor U3800 (N_3800,N_3712,N_3720);
and U3801 (N_3801,N_3756,N_3713);
and U3802 (N_3802,N_3736,N_3705);
xor U3803 (N_3803,N_3767,N_3752);
nand U3804 (N_3804,N_3753,N_3750);
nor U3805 (N_3805,N_3790,N_3718);
xnor U3806 (N_3806,N_3735,N_3769);
or U3807 (N_3807,N_3768,N_3764);
nor U3808 (N_3808,N_3774,N_3717);
nor U3809 (N_3809,N_3723,N_3791);
and U3810 (N_3810,N_3737,N_3780);
nor U3811 (N_3811,N_3798,N_3708);
nand U3812 (N_3812,N_3711,N_3773);
xor U3813 (N_3813,N_3749,N_3793);
or U3814 (N_3814,N_3724,N_3761);
xnor U3815 (N_3815,N_3741,N_3746);
nor U3816 (N_3816,N_3770,N_3784);
nand U3817 (N_3817,N_3740,N_3799);
and U3818 (N_3818,N_3727,N_3794);
or U3819 (N_3819,N_3709,N_3760);
and U3820 (N_3820,N_3706,N_3754);
nor U3821 (N_3821,N_3771,N_3762);
xnor U3822 (N_3822,N_3797,N_3786);
or U3823 (N_3823,N_3703,N_3745);
and U3824 (N_3824,N_3795,N_3701);
xnor U3825 (N_3825,N_3731,N_3716);
and U3826 (N_3826,N_3747,N_3788);
nor U3827 (N_3827,N_3730,N_3772);
nor U3828 (N_3828,N_3765,N_3700);
and U3829 (N_3829,N_3783,N_3725);
or U3830 (N_3830,N_3751,N_3789);
nor U3831 (N_3831,N_3728,N_3710);
nor U3832 (N_3832,N_3758,N_3796);
nor U3833 (N_3833,N_3733,N_3782);
and U3834 (N_3834,N_3785,N_3787);
nand U3835 (N_3835,N_3702,N_3792);
nor U3836 (N_3836,N_3722,N_3757);
and U3837 (N_3837,N_3734,N_3779);
or U3838 (N_3838,N_3715,N_3742);
or U3839 (N_3839,N_3781,N_3704);
or U3840 (N_3840,N_3759,N_3766);
xnor U3841 (N_3841,N_3744,N_3719);
or U3842 (N_3842,N_3743,N_3775);
and U3843 (N_3843,N_3721,N_3755);
and U3844 (N_3844,N_3748,N_3726);
and U3845 (N_3845,N_3729,N_3778);
nand U3846 (N_3846,N_3776,N_3777);
nor U3847 (N_3847,N_3763,N_3732);
nor U3848 (N_3848,N_3739,N_3738);
xnor U3849 (N_3849,N_3714,N_3707);
xnor U3850 (N_3850,N_3770,N_3783);
xor U3851 (N_3851,N_3717,N_3779);
and U3852 (N_3852,N_3777,N_3766);
nor U3853 (N_3853,N_3760,N_3721);
or U3854 (N_3854,N_3738,N_3750);
or U3855 (N_3855,N_3720,N_3743);
nand U3856 (N_3856,N_3781,N_3709);
nand U3857 (N_3857,N_3706,N_3791);
and U3858 (N_3858,N_3706,N_3711);
nor U3859 (N_3859,N_3744,N_3738);
or U3860 (N_3860,N_3783,N_3784);
or U3861 (N_3861,N_3726,N_3777);
nor U3862 (N_3862,N_3734,N_3789);
or U3863 (N_3863,N_3789,N_3716);
xnor U3864 (N_3864,N_3727,N_3724);
or U3865 (N_3865,N_3749,N_3736);
or U3866 (N_3866,N_3774,N_3723);
or U3867 (N_3867,N_3775,N_3742);
nor U3868 (N_3868,N_3791,N_3732);
nand U3869 (N_3869,N_3726,N_3717);
xor U3870 (N_3870,N_3766,N_3770);
nand U3871 (N_3871,N_3774,N_3783);
and U3872 (N_3872,N_3769,N_3756);
xnor U3873 (N_3873,N_3738,N_3758);
nor U3874 (N_3874,N_3706,N_3776);
xor U3875 (N_3875,N_3750,N_3716);
nand U3876 (N_3876,N_3721,N_3708);
nor U3877 (N_3877,N_3719,N_3704);
nand U3878 (N_3878,N_3757,N_3735);
and U3879 (N_3879,N_3731,N_3740);
and U3880 (N_3880,N_3710,N_3787);
xor U3881 (N_3881,N_3728,N_3721);
and U3882 (N_3882,N_3703,N_3743);
nor U3883 (N_3883,N_3781,N_3777);
or U3884 (N_3884,N_3703,N_3796);
or U3885 (N_3885,N_3756,N_3737);
xnor U3886 (N_3886,N_3773,N_3754);
nor U3887 (N_3887,N_3728,N_3770);
nand U3888 (N_3888,N_3764,N_3758);
xnor U3889 (N_3889,N_3716,N_3708);
or U3890 (N_3890,N_3764,N_3766);
xor U3891 (N_3891,N_3782,N_3773);
nor U3892 (N_3892,N_3706,N_3725);
nor U3893 (N_3893,N_3772,N_3784);
nand U3894 (N_3894,N_3728,N_3716);
or U3895 (N_3895,N_3730,N_3793);
or U3896 (N_3896,N_3767,N_3777);
or U3897 (N_3897,N_3795,N_3778);
or U3898 (N_3898,N_3728,N_3705);
nor U3899 (N_3899,N_3799,N_3794);
nor U3900 (N_3900,N_3808,N_3867);
xor U3901 (N_3901,N_3885,N_3845);
and U3902 (N_3902,N_3864,N_3844);
nor U3903 (N_3903,N_3840,N_3828);
nand U3904 (N_3904,N_3850,N_3877);
nor U3905 (N_3905,N_3831,N_3841);
nor U3906 (N_3906,N_3849,N_3825);
nor U3907 (N_3907,N_3848,N_3815);
xnor U3908 (N_3908,N_3819,N_3878);
xor U3909 (N_3909,N_3807,N_3884);
or U3910 (N_3910,N_3860,N_3896);
and U3911 (N_3911,N_3846,N_3870);
nand U3912 (N_3912,N_3869,N_3824);
or U3913 (N_3913,N_3811,N_3855);
and U3914 (N_3914,N_3865,N_3895);
nand U3915 (N_3915,N_3843,N_3888);
and U3916 (N_3916,N_3879,N_3871);
or U3917 (N_3917,N_3829,N_3817);
and U3918 (N_3918,N_3803,N_3882);
or U3919 (N_3919,N_3886,N_3813);
xor U3920 (N_3920,N_3891,N_3894);
xnor U3921 (N_3921,N_3832,N_3881);
nand U3922 (N_3922,N_3821,N_3834);
and U3923 (N_3923,N_3826,N_3857);
and U3924 (N_3924,N_3875,N_3863);
and U3925 (N_3925,N_3837,N_3830);
or U3926 (N_3926,N_3839,N_3872);
nand U3927 (N_3927,N_3866,N_3823);
or U3928 (N_3928,N_3836,N_3810);
or U3929 (N_3929,N_3822,N_3801);
nand U3930 (N_3930,N_3809,N_3890);
or U3931 (N_3931,N_3851,N_3876);
xor U3932 (N_3932,N_3806,N_3838);
or U3933 (N_3933,N_3861,N_3892);
xnor U3934 (N_3934,N_3868,N_3816);
xor U3935 (N_3935,N_3842,N_3854);
nor U3936 (N_3936,N_3800,N_3812);
nand U3937 (N_3937,N_3880,N_3835);
or U3938 (N_3938,N_3862,N_3827);
nor U3939 (N_3939,N_3858,N_3833);
nand U3940 (N_3940,N_3873,N_3883);
nand U3941 (N_3941,N_3852,N_3804);
nand U3942 (N_3942,N_3874,N_3897);
or U3943 (N_3943,N_3893,N_3802);
and U3944 (N_3944,N_3847,N_3898);
or U3945 (N_3945,N_3889,N_3887);
or U3946 (N_3946,N_3820,N_3805);
nand U3947 (N_3947,N_3818,N_3856);
nor U3948 (N_3948,N_3814,N_3853);
or U3949 (N_3949,N_3859,N_3899);
or U3950 (N_3950,N_3818,N_3854);
xnor U3951 (N_3951,N_3879,N_3845);
xnor U3952 (N_3952,N_3837,N_3848);
nand U3953 (N_3953,N_3860,N_3865);
nor U3954 (N_3954,N_3886,N_3864);
or U3955 (N_3955,N_3890,N_3876);
and U3956 (N_3956,N_3877,N_3894);
xnor U3957 (N_3957,N_3838,N_3804);
nor U3958 (N_3958,N_3859,N_3864);
nor U3959 (N_3959,N_3810,N_3856);
nor U3960 (N_3960,N_3897,N_3801);
nand U3961 (N_3961,N_3806,N_3848);
and U3962 (N_3962,N_3815,N_3870);
and U3963 (N_3963,N_3877,N_3807);
nand U3964 (N_3964,N_3811,N_3833);
xnor U3965 (N_3965,N_3827,N_3897);
and U3966 (N_3966,N_3815,N_3898);
or U3967 (N_3967,N_3806,N_3829);
or U3968 (N_3968,N_3810,N_3806);
nand U3969 (N_3969,N_3896,N_3806);
xnor U3970 (N_3970,N_3874,N_3873);
and U3971 (N_3971,N_3825,N_3846);
xor U3972 (N_3972,N_3833,N_3824);
and U3973 (N_3973,N_3877,N_3832);
or U3974 (N_3974,N_3883,N_3891);
nand U3975 (N_3975,N_3877,N_3875);
xnor U3976 (N_3976,N_3890,N_3846);
nor U3977 (N_3977,N_3824,N_3806);
or U3978 (N_3978,N_3845,N_3855);
and U3979 (N_3979,N_3895,N_3820);
nor U3980 (N_3980,N_3812,N_3887);
nand U3981 (N_3981,N_3829,N_3885);
nor U3982 (N_3982,N_3873,N_3821);
nand U3983 (N_3983,N_3863,N_3830);
or U3984 (N_3984,N_3881,N_3887);
nand U3985 (N_3985,N_3835,N_3878);
nor U3986 (N_3986,N_3803,N_3832);
and U3987 (N_3987,N_3860,N_3862);
nor U3988 (N_3988,N_3827,N_3820);
xor U3989 (N_3989,N_3820,N_3898);
or U3990 (N_3990,N_3806,N_3846);
nor U3991 (N_3991,N_3815,N_3874);
nor U3992 (N_3992,N_3863,N_3867);
or U3993 (N_3993,N_3842,N_3875);
nand U3994 (N_3994,N_3801,N_3835);
nand U3995 (N_3995,N_3838,N_3811);
nor U3996 (N_3996,N_3890,N_3823);
nor U3997 (N_3997,N_3887,N_3826);
or U3998 (N_3998,N_3863,N_3872);
and U3999 (N_3999,N_3865,N_3836);
and U4000 (N_4000,N_3999,N_3985);
and U4001 (N_4001,N_3958,N_3981);
nor U4002 (N_4002,N_3984,N_3903);
and U4003 (N_4003,N_3991,N_3912);
nand U4004 (N_4004,N_3975,N_3972);
or U4005 (N_4005,N_3950,N_3964);
nand U4006 (N_4006,N_3966,N_3979);
and U4007 (N_4007,N_3987,N_3995);
nor U4008 (N_4008,N_3943,N_3938);
xnor U4009 (N_4009,N_3928,N_3986);
or U4010 (N_4010,N_3990,N_3937);
or U4011 (N_4011,N_3948,N_3947);
nand U4012 (N_4012,N_3942,N_3968);
nor U4013 (N_4013,N_3996,N_3926);
and U4014 (N_4014,N_3924,N_3982);
and U4015 (N_4015,N_3992,N_3967);
nand U4016 (N_4016,N_3901,N_3998);
nor U4017 (N_4017,N_3955,N_3956);
nand U4018 (N_4018,N_3946,N_3906);
and U4019 (N_4019,N_3909,N_3969);
nor U4020 (N_4020,N_3902,N_3963);
xnor U4021 (N_4021,N_3957,N_3951);
nand U4022 (N_4022,N_3934,N_3941);
or U4023 (N_4023,N_3915,N_3971);
and U4024 (N_4024,N_3904,N_3916);
and U4025 (N_4025,N_3918,N_3935);
nor U4026 (N_4026,N_3931,N_3932);
or U4027 (N_4027,N_3989,N_3921);
nor U4028 (N_4028,N_3940,N_3923);
or U4029 (N_4029,N_3959,N_3954);
or U4030 (N_4030,N_3939,N_3910);
and U4031 (N_4031,N_3927,N_3945);
and U4032 (N_4032,N_3922,N_3953);
nand U4033 (N_4033,N_3933,N_3930);
and U4034 (N_4034,N_3952,N_3978);
or U4035 (N_4035,N_3960,N_3907);
xnor U4036 (N_4036,N_3919,N_3980);
nor U4037 (N_4037,N_3900,N_3911);
nor U4038 (N_4038,N_3993,N_3983);
and U4039 (N_4039,N_3917,N_3929);
nor U4040 (N_4040,N_3974,N_3965);
or U4041 (N_4041,N_3976,N_3997);
xor U4042 (N_4042,N_3944,N_3977);
or U4043 (N_4043,N_3988,N_3949);
nand U4044 (N_4044,N_3961,N_3913);
nand U4045 (N_4045,N_3914,N_3920);
and U4046 (N_4046,N_3970,N_3908);
nand U4047 (N_4047,N_3905,N_3962);
nor U4048 (N_4048,N_3973,N_3925);
nor U4049 (N_4049,N_3994,N_3936);
and U4050 (N_4050,N_3971,N_3944);
xor U4051 (N_4051,N_3916,N_3932);
nor U4052 (N_4052,N_3955,N_3997);
or U4053 (N_4053,N_3998,N_3986);
or U4054 (N_4054,N_3954,N_3969);
xnor U4055 (N_4055,N_3923,N_3994);
xnor U4056 (N_4056,N_3944,N_3915);
or U4057 (N_4057,N_3996,N_3985);
nand U4058 (N_4058,N_3916,N_3966);
nand U4059 (N_4059,N_3918,N_3905);
nand U4060 (N_4060,N_3995,N_3922);
nor U4061 (N_4061,N_3925,N_3971);
or U4062 (N_4062,N_3909,N_3927);
nor U4063 (N_4063,N_3909,N_3976);
or U4064 (N_4064,N_3954,N_3961);
nand U4065 (N_4065,N_3916,N_3905);
or U4066 (N_4066,N_3981,N_3928);
and U4067 (N_4067,N_3978,N_3908);
xnor U4068 (N_4068,N_3969,N_3938);
xor U4069 (N_4069,N_3963,N_3906);
nor U4070 (N_4070,N_3915,N_3946);
or U4071 (N_4071,N_3952,N_3958);
xor U4072 (N_4072,N_3993,N_3959);
or U4073 (N_4073,N_3901,N_3915);
nor U4074 (N_4074,N_3989,N_3969);
and U4075 (N_4075,N_3913,N_3986);
nor U4076 (N_4076,N_3905,N_3990);
or U4077 (N_4077,N_3947,N_3906);
xnor U4078 (N_4078,N_3950,N_3915);
xor U4079 (N_4079,N_3926,N_3973);
xor U4080 (N_4080,N_3908,N_3925);
and U4081 (N_4081,N_3910,N_3937);
nor U4082 (N_4082,N_3990,N_3944);
nor U4083 (N_4083,N_3926,N_3933);
and U4084 (N_4084,N_3978,N_3925);
nand U4085 (N_4085,N_3958,N_3983);
and U4086 (N_4086,N_3915,N_3926);
xnor U4087 (N_4087,N_3904,N_3985);
nand U4088 (N_4088,N_3979,N_3938);
or U4089 (N_4089,N_3979,N_3916);
nand U4090 (N_4090,N_3945,N_3958);
or U4091 (N_4091,N_3970,N_3978);
nor U4092 (N_4092,N_3915,N_3931);
and U4093 (N_4093,N_3967,N_3926);
nor U4094 (N_4094,N_3952,N_3999);
nor U4095 (N_4095,N_3988,N_3908);
nand U4096 (N_4096,N_3929,N_3998);
and U4097 (N_4097,N_3931,N_3918);
nand U4098 (N_4098,N_3921,N_3965);
nor U4099 (N_4099,N_3950,N_3971);
or U4100 (N_4100,N_4049,N_4091);
and U4101 (N_4101,N_4047,N_4038);
nand U4102 (N_4102,N_4041,N_4045);
xnor U4103 (N_4103,N_4007,N_4065);
and U4104 (N_4104,N_4002,N_4016);
nor U4105 (N_4105,N_4009,N_4088);
and U4106 (N_4106,N_4015,N_4072);
xnor U4107 (N_4107,N_4095,N_4003);
nor U4108 (N_4108,N_4017,N_4010);
and U4109 (N_4109,N_4078,N_4066);
and U4110 (N_4110,N_4057,N_4068);
or U4111 (N_4111,N_4028,N_4004);
and U4112 (N_4112,N_4051,N_4096);
nand U4113 (N_4113,N_4055,N_4019);
nor U4114 (N_4114,N_4084,N_4060);
or U4115 (N_4115,N_4056,N_4021);
nor U4116 (N_4116,N_4062,N_4058);
nor U4117 (N_4117,N_4031,N_4027);
xor U4118 (N_4118,N_4013,N_4086);
nand U4119 (N_4119,N_4024,N_4073);
nor U4120 (N_4120,N_4067,N_4026);
nor U4121 (N_4121,N_4033,N_4040);
xor U4122 (N_4122,N_4050,N_4014);
xor U4123 (N_4123,N_4069,N_4097);
nor U4124 (N_4124,N_4048,N_4023);
xnor U4125 (N_4125,N_4099,N_4032);
nor U4126 (N_4126,N_4063,N_4018);
xor U4127 (N_4127,N_4092,N_4075);
or U4128 (N_4128,N_4089,N_4093);
xor U4129 (N_4129,N_4064,N_4074);
or U4130 (N_4130,N_4054,N_4034);
nor U4131 (N_4131,N_4044,N_4042);
nand U4132 (N_4132,N_4083,N_4029);
nor U4133 (N_4133,N_4071,N_4022);
or U4134 (N_4134,N_4081,N_4087);
nand U4135 (N_4135,N_4076,N_4053);
nand U4136 (N_4136,N_4020,N_4030);
nand U4137 (N_4137,N_4061,N_4039);
and U4138 (N_4138,N_4070,N_4052);
or U4139 (N_4139,N_4043,N_4059);
and U4140 (N_4140,N_4000,N_4006);
nor U4141 (N_4141,N_4011,N_4079);
xnor U4142 (N_4142,N_4077,N_4001);
nor U4143 (N_4143,N_4094,N_4005);
or U4144 (N_4144,N_4046,N_4008);
xor U4145 (N_4145,N_4025,N_4037);
or U4146 (N_4146,N_4098,N_4080);
or U4147 (N_4147,N_4085,N_4082);
xor U4148 (N_4148,N_4012,N_4036);
and U4149 (N_4149,N_4090,N_4035);
nor U4150 (N_4150,N_4062,N_4057);
nand U4151 (N_4151,N_4035,N_4040);
and U4152 (N_4152,N_4017,N_4070);
and U4153 (N_4153,N_4019,N_4015);
and U4154 (N_4154,N_4083,N_4047);
nand U4155 (N_4155,N_4074,N_4019);
nand U4156 (N_4156,N_4059,N_4034);
nor U4157 (N_4157,N_4064,N_4003);
or U4158 (N_4158,N_4055,N_4059);
nand U4159 (N_4159,N_4038,N_4082);
nand U4160 (N_4160,N_4046,N_4089);
and U4161 (N_4161,N_4068,N_4004);
nor U4162 (N_4162,N_4062,N_4068);
nor U4163 (N_4163,N_4026,N_4082);
xnor U4164 (N_4164,N_4078,N_4081);
and U4165 (N_4165,N_4093,N_4047);
or U4166 (N_4166,N_4098,N_4022);
nand U4167 (N_4167,N_4052,N_4048);
nand U4168 (N_4168,N_4017,N_4094);
or U4169 (N_4169,N_4096,N_4055);
xnor U4170 (N_4170,N_4034,N_4058);
xnor U4171 (N_4171,N_4061,N_4077);
or U4172 (N_4172,N_4040,N_4079);
xnor U4173 (N_4173,N_4083,N_4053);
and U4174 (N_4174,N_4028,N_4041);
and U4175 (N_4175,N_4078,N_4052);
nor U4176 (N_4176,N_4063,N_4007);
and U4177 (N_4177,N_4061,N_4017);
or U4178 (N_4178,N_4031,N_4038);
nand U4179 (N_4179,N_4073,N_4056);
nor U4180 (N_4180,N_4084,N_4009);
nand U4181 (N_4181,N_4010,N_4005);
nor U4182 (N_4182,N_4003,N_4007);
nor U4183 (N_4183,N_4004,N_4009);
and U4184 (N_4184,N_4098,N_4040);
or U4185 (N_4185,N_4053,N_4026);
xnor U4186 (N_4186,N_4008,N_4079);
or U4187 (N_4187,N_4056,N_4098);
xor U4188 (N_4188,N_4087,N_4069);
nor U4189 (N_4189,N_4007,N_4038);
nor U4190 (N_4190,N_4038,N_4093);
xnor U4191 (N_4191,N_4063,N_4032);
and U4192 (N_4192,N_4056,N_4057);
nor U4193 (N_4193,N_4097,N_4009);
or U4194 (N_4194,N_4056,N_4018);
xnor U4195 (N_4195,N_4039,N_4018);
nor U4196 (N_4196,N_4031,N_4021);
nor U4197 (N_4197,N_4034,N_4084);
nand U4198 (N_4198,N_4036,N_4033);
nand U4199 (N_4199,N_4035,N_4098);
and U4200 (N_4200,N_4193,N_4133);
xnor U4201 (N_4201,N_4113,N_4174);
xor U4202 (N_4202,N_4160,N_4170);
nor U4203 (N_4203,N_4126,N_4194);
or U4204 (N_4204,N_4123,N_4153);
or U4205 (N_4205,N_4192,N_4135);
or U4206 (N_4206,N_4129,N_4151);
xor U4207 (N_4207,N_4142,N_4122);
and U4208 (N_4208,N_4195,N_4163);
nand U4209 (N_4209,N_4152,N_4148);
or U4210 (N_4210,N_4141,N_4199);
nor U4211 (N_4211,N_4150,N_4182);
xnor U4212 (N_4212,N_4127,N_4100);
or U4213 (N_4213,N_4196,N_4118);
nand U4214 (N_4214,N_4146,N_4107);
xor U4215 (N_4215,N_4185,N_4155);
xor U4216 (N_4216,N_4168,N_4139);
nor U4217 (N_4217,N_4124,N_4131);
xor U4218 (N_4218,N_4156,N_4157);
xnor U4219 (N_4219,N_4119,N_4120);
and U4220 (N_4220,N_4191,N_4180);
or U4221 (N_4221,N_4109,N_4136);
and U4222 (N_4222,N_4110,N_4162);
and U4223 (N_4223,N_4128,N_4116);
and U4224 (N_4224,N_4172,N_4165);
nor U4225 (N_4225,N_4158,N_4145);
and U4226 (N_4226,N_4132,N_4198);
or U4227 (N_4227,N_4106,N_4167);
nor U4228 (N_4228,N_4114,N_4117);
or U4229 (N_4229,N_4112,N_4137);
xnor U4230 (N_4230,N_4104,N_4105);
xor U4231 (N_4231,N_4164,N_4177);
xnor U4232 (N_4232,N_4173,N_4103);
or U4233 (N_4233,N_4159,N_4115);
nor U4234 (N_4234,N_4149,N_4138);
nor U4235 (N_4235,N_4140,N_4161);
xor U4236 (N_4236,N_4183,N_4178);
or U4237 (N_4237,N_4175,N_4108);
nor U4238 (N_4238,N_4189,N_4101);
xor U4239 (N_4239,N_4184,N_4181);
xnor U4240 (N_4240,N_4187,N_4147);
and U4241 (N_4241,N_4179,N_4171);
or U4242 (N_4242,N_4121,N_4143);
or U4243 (N_4243,N_4102,N_4186);
nor U4244 (N_4244,N_4144,N_4197);
or U4245 (N_4245,N_4188,N_4130);
xor U4246 (N_4246,N_4190,N_4169);
or U4247 (N_4247,N_4176,N_4111);
nor U4248 (N_4248,N_4166,N_4125);
and U4249 (N_4249,N_4154,N_4134);
or U4250 (N_4250,N_4140,N_4145);
and U4251 (N_4251,N_4115,N_4157);
or U4252 (N_4252,N_4104,N_4193);
or U4253 (N_4253,N_4116,N_4166);
nand U4254 (N_4254,N_4147,N_4130);
and U4255 (N_4255,N_4128,N_4176);
nand U4256 (N_4256,N_4182,N_4151);
or U4257 (N_4257,N_4138,N_4129);
and U4258 (N_4258,N_4186,N_4191);
nor U4259 (N_4259,N_4130,N_4138);
xnor U4260 (N_4260,N_4123,N_4101);
and U4261 (N_4261,N_4197,N_4134);
xnor U4262 (N_4262,N_4116,N_4184);
and U4263 (N_4263,N_4196,N_4153);
xor U4264 (N_4264,N_4134,N_4114);
and U4265 (N_4265,N_4127,N_4114);
nand U4266 (N_4266,N_4108,N_4134);
or U4267 (N_4267,N_4191,N_4153);
or U4268 (N_4268,N_4152,N_4114);
and U4269 (N_4269,N_4185,N_4101);
nand U4270 (N_4270,N_4167,N_4132);
or U4271 (N_4271,N_4125,N_4160);
xor U4272 (N_4272,N_4142,N_4161);
nor U4273 (N_4273,N_4177,N_4116);
xor U4274 (N_4274,N_4198,N_4134);
xor U4275 (N_4275,N_4188,N_4118);
xnor U4276 (N_4276,N_4171,N_4187);
and U4277 (N_4277,N_4188,N_4195);
nand U4278 (N_4278,N_4142,N_4157);
nor U4279 (N_4279,N_4193,N_4126);
xnor U4280 (N_4280,N_4115,N_4119);
xor U4281 (N_4281,N_4125,N_4132);
xnor U4282 (N_4282,N_4128,N_4178);
nand U4283 (N_4283,N_4164,N_4102);
nand U4284 (N_4284,N_4148,N_4186);
or U4285 (N_4285,N_4151,N_4190);
or U4286 (N_4286,N_4142,N_4134);
xnor U4287 (N_4287,N_4172,N_4135);
xor U4288 (N_4288,N_4149,N_4191);
nand U4289 (N_4289,N_4156,N_4184);
nor U4290 (N_4290,N_4168,N_4122);
or U4291 (N_4291,N_4157,N_4170);
nor U4292 (N_4292,N_4123,N_4195);
xor U4293 (N_4293,N_4132,N_4106);
nand U4294 (N_4294,N_4175,N_4152);
nand U4295 (N_4295,N_4153,N_4131);
or U4296 (N_4296,N_4177,N_4167);
nor U4297 (N_4297,N_4147,N_4137);
and U4298 (N_4298,N_4144,N_4157);
xnor U4299 (N_4299,N_4107,N_4150);
nand U4300 (N_4300,N_4276,N_4215);
or U4301 (N_4301,N_4212,N_4245);
or U4302 (N_4302,N_4222,N_4299);
nor U4303 (N_4303,N_4219,N_4213);
xor U4304 (N_4304,N_4267,N_4252);
nor U4305 (N_4305,N_4255,N_4253);
or U4306 (N_4306,N_4209,N_4207);
nor U4307 (N_4307,N_4214,N_4229);
nand U4308 (N_4308,N_4247,N_4206);
and U4309 (N_4309,N_4208,N_4243);
nand U4310 (N_4310,N_4290,N_4224);
or U4311 (N_4311,N_4280,N_4272);
and U4312 (N_4312,N_4271,N_4204);
xnor U4313 (N_4313,N_4223,N_4251);
nor U4314 (N_4314,N_4234,N_4261);
nand U4315 (N_4315,N_4289,N_4286);
nor U4316 (N_4316,N_4244,N_4236);
nand U4317 (N_4317,N_4278,N_4266);
and U4318 (N_4318,N_4230,N_4295);
and U4319 (N_4319,N_4281,N_4233);
xnor U4320 (N_4320,N_4293,N_4220);
nand U4321 (N_4321,N_4227,N_4226);
or U4322 (N_4322,N_4202,N_4288);
and U4323 (N_4323,N_4274,N_4211);
and U4324 (N_4324,N_4218,N_4283);
xnor U4325 (N_4325,N_4260,N_4200);
nor U4326 (N_4326,N_4294,N_4250);
xor U4327 (N_4327,N_4254,N_4275);
nor U4328 (N_4328,N_4232,N_4259);
or U4329 (N_4329,N_4231,N_4264);
nand U4330 (N_4330,N_4285,N_4291);
nor U4331 (N_4331,N_4205,N_4269);
xnor U4332 (N_4332,N_4221,N_4297);
and U4333 (N_4333,N_4268,N_4228);
xnor U4334 (N_4334,N_4258,N_4265);
or U4335 (N_4335,N_4210,N_4298);
or U4336 (N_4336,N_4242,N_4287);
or U4337 (N_4337,N_4296,N_4235);
xor U4338 (N_4338,N_4292,N_4216);
or U4339 (N_4339,N_4239,N_4249);
nand U4340 (N_4340,N_4238,N_4263);
nand U4341 (N_4341,N_4246,N_4225);
nor U4342 (N_4342,N_4256,N_4241);
xnor U4343 (N_4343,N_4277,N_4201);
nand U4344 (N_4344,N_4240,N_4273);
nor U4345 (N_4345,N_4203,N_4257);
nand U4346 (N_4346,N_4237,N_4270);
and U4347 (N_4347,N_4262,N_4217);
nand U4348 (N_4348,N_4279,N_4282);
or U4349 (N_4349,N_4284,N_4248);
or U4350 (N_4350,N_4280,N_4279);
and U4351 (N_4351,N_4203,N_4207);
or U4352 (N_4352,N_4244,N_4270);
or U4353 (N_4353,N_4239,N_4242);
nor U4354 (N_4354,N_4251,N_4265);
xnor U4355 (N_4355,N_4293,N_4205);
xor U4356 (N_4356,N_4294,N_4295);
or U4357 (N_4357,N_4264,N_4278);
or U4358 (N_4358,N_4269,N_4246);
nor U4359 (N_4359,N_4262,N_4223);
nand U4360 (N_4360,N_4215,N_4251);
or U4361 (N_4361,N_4271,N_4225);
or U4362 (N_4362,N_4231,N_4269);
xor U4363 (N_4363,N_4291,N_4264);
and U4364 (N_4364,N_4253,N_4244);
and U4365 (N_4365,N_4244,N_4230);
xnor U4366 (N_4366,N_4288,N_4271);
nand U4367 (N_4367,N_4267,N_4264);
and U4368 (N_4368,N_4234,N_4246);
and U4369 (N_4369,N_4208,N_4214);
nand U4370 (N_4370,N_4209,N_4234);
xor U4371 (N_4371,N_4232,N_4290);
xnor U4372 (N_4372,N_4262,N_4214);
nand U4373 (N_4373,N_4215,N_4203);
or U4374 (N_4374,N_4295,N_4210);
xor U4375 (N_4375,N_4263,N_4225);
and U4376 (N_4376,N_4239,N_4216);
xor U4377 (N_4377,N_4283,N_4281);
and U4378 (N_4378,N_4204,N_4215);
xnor U4379 (N_4379,N_4252,N_4266);
and U4380 (N_4380,N_4201,N_4210);
nand U4381 (N_4381,N_4218,N_4238);
nor U4382 (N_4382,N_4247,N_4200);
and U4383 (N_4383,N_4200,N_4222);
and U4384 (N_4384,N_4256,N_4221);
and U4385 (N_4385,N_4242,N_4253);
and U4386 (N_4386,N_4205,N_4217);
nor U4387 (N_4387,N_4214,N_4225);
nor U4388 (N_4388,N_4225,N_4243);
or U4389 (N_4389,N_4282,N_4281);
xor U4390 (N_4390,N_4294,N_4272);
nor U4391 (N_4391,N_4253,N_4291);
nor U4392 (N_4392,N_4262,N_4202);
xnor U4393 (N_4393,N_4215,N_4202);
and U4394 (N_4394,N_4211,N_4231);
xor U4395 (N_4395,N_4233,N_4285);
and U4396 (N_4396,N_4294,N_4200);
nand U4397 (N_4397,N_4253,N_4216);
nand U4398 (N_4398,N_4208,N_4230);
and U4399 (N_4399,N_4221,N_4233);
nor U4400 (N_4400,N_4348,N_4392);
and U4401 (N_4401,N_4355,N_4395);
or U4402 (N_4402,N_4304,N_4353);
and U4403 (N_4403,N_4347,N_4331);
nor U4404 (N_4404,N_4374,N_4307);
nor U4405 (N_4405,N_4324,N_4337);
or U4406 (N_4406,N_4352,N_4356);
and U4407 (N_4407,N_4343,N_4351);
xor U4408 (N_4408,N_4373,N_4339);
xnor U4409 (N_4409,N_4384,N_4314);
nand U4410 (N_4410,N_4379,N_4359);
nor U4411 (N_4411,N_4377,N_4323);
nand U4412 (N_4412,N_4345,N_4391);
nor U4413 (N_4413,N_4309,N_4358);
and U4414 (N_4414,N_4388,N_4301);
and U4415 (N_4415,N_4378,N_4306);
or U4416 (N_4416,N_4372,N_4381);
or U4417 (N_4417,N_4399,N_4394);
xnor U4418 (N_4418,N_4310,N_4313);
nor U4419 (N_4419,N_4300,N_4375);
and U4420 (N_4420,N_4317,N_4383);
or U4421 (N_4421,N_4332,N_4369);
nand U4422 (N_4422,N_4311,N_4342);
and U4423 (N_4423,N_4334,N_4363);
or U4424 (N_4424,N_4329,N_4349);
xnor U4425 (N_4425,N_4326,N_4357);
or U4426 (N_4426,N_4341,N_4389);
or U4427 (N_4427,N_4344,N_4371);
nand U4428 (N_4428,N_4346,N_4328);
xor U4429 (N_4429,N_4318,N_4316);
nand U4430 (N_4430,N_4303,N_4396);
and U4431 (N_4431,N_4365,N_4302);
nor U4432 (N_4432,N_4319,N_4398);
or U4433 (N_4433,N_4362,N_4370);
nor U4434 (N_4434,N_4364,N_4335);
nor U4435 (N_4435,N_4336,N_4321);
nor U4436 (N_4436,N_4340,N_4308);
nor U4437 (N_4437,N_4322,N_4387);
nor U4438 (N_4438,N_4305,N_4390);
xor U4439 (N_4439,N_4315,N_4366);
nand U4440 (N_4440,N_4393,N_4380);
nor U4441 (N_4441,N_4338,N_4330);
xnor U4442 (N_4442,N_4385,N_4367);
and U4443 (N_4443,N_4320,N_4397);
xor U4444 (N_4444,N_4333,N_4360);
or U4445 (N_4445,N_4350,N_4361);
and U4446 (N_4446,N_4376,N_4312);
and U4447 (N_4447,N_4382,N_4327);
nand U4448 (N_4448,N_4368,N_4386);
or U4449 (N_4449,N_4325,N_4354);
or U4450 (N_4450,N_4347,N_4374);
nand U4451 (N_4451,N_4327,N_4323);
nor U4452 (N_4452,N_4368,N_4390);
nor U4453 (N_4453,N_4363,N_4322);
xor U4454 (N_4454,N_4305,N_4373);
or U4455 (N_4455,N_4336,N_4396);
nor U4456 (N_4456,N_4350,N_4371);
nand U4457 (N_4457,N_4370,N_4304);
nand U4458 (N_4458,N_4339,N_4367);
nand U4459 (N_4459,N_4352,N_4395);
nor U4460 (N_4460,N_4379,N_4319);
nand U4461 (N_4461,N_4374,N_4353);
or U4462 (N_4462,N_4364,N_4366);
or U4463 (N_4463,N_4388,N_4331);
xnor U4464 (N_4464,N_4381,N_4334);
or U4465 (N_4465,N_4392,N_4317);
nor U4466 (N_4466,N_4378,N_4395);
xnor U4467 (N_4467,N_4312,N_4399);
xnor U4468 (N_4468,N_4355,N_4351);
nor U4469 (N_4469,N_4304,N_4375);
nor U4470 (N_4470,N_4367,N_4389);
nor U4471 (N_4471,N_4396,N_4370);
nor U4472 (N_4472,N_4351,N_4323);
xor U4473 (N_4473,N_4376,N_4370);
xnor U4474 (N_4474,N_4348,N_4370);
nand U4475 (N_4475,N_4331,N_4307);
nand U4476 (N_4476,N_4373,N_4312);
nor U4477 (N_4477,N_4386,N_4397);
xnor U4478 (N_4478,N_4394,N_4370);
or U4479 (N_4479,N_4354,N_4337);
or U4480 (N_4480,N_4390,N_4328);
nand U4481 (N_4481,N_4354,N_4366);
nand U4482 (N_4482,N_4374,N_4375);
or U4483 (N_4483,N_4301,N_4331);
or U4484 (N_4484,N_4319,N_4321);
or U4485 (N_4485,N_4342,N_4303);
xor U4486 (N_4486,N_4364,N_4352);
xor U4487 (N_4487,N_4325,N_4379);
xor U4488 (N_4488,N_4370,N_4310);
xor U4489 (N_4489,N_4349,N_4308);
xnor U4490 (N_4490,N_4316,N_4367);
or U4491 (N_4491,N_4352,N_4399);
and U4492 (N_4492,N_4358,N_4302);
nor U4493 (N_4493,N_4312,N_4338);
and U4494 (N_4494,N_4334,N_4397);
nand U4495 (N_4495,N_4351,N_4365);
nand U4496 (N_4496,N_4349,N_4324);
nor U4497 (N_4497,N_4312,N_4365);
nor U4498 (N_4498,N_4391,N_4359);
xor U4499 (N_4499,N_4349,N_4348);
or U4500 (N_4500,N_4457,N_4487);
nor U4501 (N_4501,N_4497,N_4483);
xnor U4502 (N_4502,N_4458,N_4449);
nor U4503 (N_4503,N_4450,N_4433);
nor U4504 (N_4504,N_4400,N_4431);
or U4505 (N_4505,N_4437,N_4499);
xor U4506 (N_4506,N_4461,N_4448);
and U4507 (N_4507,N_4467,N_4492);
nor U4508 (N_4508,N_4496,N_4465);
or U4509 (N_4509,N_4444,N_4479);
nor U4510 (N_4510,N_4428,N_4459);
nor U4511 (N_4511,N_4481,N_4435);
xor U4512 (N_4512,N_4452,N_4469);
and U4513 (N_4513,N_4493,N_4468);
nand U4514 (N_4514,N_4427,N_4436);
or U4515 (N_4515,N_4418,N_4485);
xor U4516 (N_4516,N_4447,N_4422);
nand U4517 (N_4517,N_4421,N_4460);
xnor U4518 (N_4518,N_4474,N_4462);
and U4519 (N_4519,N_4408,N_4445);
xor U4520 (N_4520,N_4443,N_4470);
nor U4521 (N_4521,N_4410,N_4404);
or U4522 (N_4522,N_4464,N_4415);
nand U4523 (N_4523,N_4406,N_4432);
nor U4524 (N_4524,N_4453,N_4405);
and U4525 (N_4525,N_4407,N_4403);
nand U4526 (N_4526,N_4426,N_4429);
or U4527 (N_4527,N_4473,N_4489);
nand U4528 (N_4528,N_4401,N_4440);
and U4529 (N_4529,N_4476,N_4439);
or U4530 (N_4530,N_4425,N_4482);
nor U4531 (N_4531,N_4491,N_4419);
nor U4532 (N_4532,N_4451,N_4423);
nand U4533 (N_4533,N_4456,N_4455);
nor U4534 (N_4534,N_4494,N_4420);
nand U4535 (N_4535,N_4434,N_4402);
or U4536 (N_4536,N_4475,N_4477);
xor U4537 (N_4537,N_4417,N_4430);
and U4538 (N_4538,N_4441,N_4409);
and U4539 (N_4539,N_4478,N_4463);
or U4540 (N_4540,N_4471,N_4484);
or U4541 (N_4541,N_4416,N_4490);
and U4542 (N_4542,N_4438,N_4424);
nor U4543 (N_4543,N_4412,N_4480);
and U4544 (N_4544,N_4442,N_4498);
nand U4545 (N_4545,N_4454,N_4495);
and U4546 (N_4546,N_4413,N_4472);
and U4547 (N_4547,N_4414,N_4466);
xnor U4548 (N_4548,N_4488,N_4486);
or U4549 (N_4549,N_4411,N_4446);
and U4550 (N_4550,N_4418,N_4430);
or U4551 (N_4551,N_4432,N_4487);
xnor U4552 (N_4552,N_4401,N_4481);
xnor U4553 (N_4553,N_4444,N_4419);
nand U4554 (N_4554,N_4441,N_4427);
nand U4555 (N_4555,N_4408,N_4427);
nand U4556 (N_4556,N_4443,N_4491);
nor U4557 (N_4557,N_4456,N_4485);
xnor U4558 (N_4558,N_4467,N_4494);
xnor U4559 (N_4559,N_4493,N_4439);
or U4560 (N_4560,N_4413,N_4475);
and U4561 (N_4561,N_4486,N_4492);
or U4562 (N_4562,N_4472,N_4448);
xor U4563 (N_4563,N_4444,N_4469);
nand U4564 (N_4564,N_4436,N_4411);
xor U4565 (N_4565,N_4467,N_4487);
xnor U4566 (N_4566,N_4401,N_4418);
nand U4567 (N_4567,N_4408,N_4484);
xnor U4568 (N_4568,N_4499,N_4428);
nor U4569 (N_4569,N_4458,N_4429);
or U4570 (N_4570,N_4421,N_4401);
and U4571 (N_4571,N_4473,N_4478);
or U4572 (N_4572,N_4477,N_4420);
xor U4573 (N_4573,N_4455,N_4443);
or U4574 (N_4574,N_4430,N_4421);
nand U4575 (N_4575,N_4462,N_4469);
and U4576 (N_4576,N_4460,N_4481);
nand U4577 (N_4577,N_4482,N_4490);
and U4578 (N_4578,N_4457,N_4473);
nand U4579 (N_4579,N_4481,N_4461);
nand U4580 (N_4580,N_4493,N_4454);
xnor U4581 (N_4581,N_4486,N_4460);
nor U4582 (N_4582,N_4431,N_4420);
and U4583 (N_4583,N_4475,N_4448);
nand U4584 (N_4584,N_4472,N_4484);
nor U4585 (N_4585,N_4452,N_4440);
nand U4586 (N_4586,N_4473,N_4439);
nor U4587 (N_4587,N_4406,N_4485);
and U4588 (N_4588,N_4489,N_4458);
xnor U4589 (N_4589,N_4465,N_4485);
or U4590 (N_4590,N_4494,N_4405);
and U4591 (N_4591,N_4470,N_4447);
and U4592 (N_4592,N_4464,N_4496);
nor U4593 (N_4593,N_4470,N_4459);
nor U4594 (N_4594,N_4433,N_4454);
or U4595 (N_4595,N_4464,N_4495);
nand U4596 (N_4596,N_4439,N_4450);
nor U4597 (N_4597,N_4456,N_4425);
nand U4598 (N_4598,N_4489,N_4461);
and U4599 (N_4599,N_4444,N_4409);
or U4600 (N_4600,N_4577,N_4582);
or U4601 (N_4601,N_4553,N_4523);
or U4602 (N_4602,N_4566,N_4540);
nand U4603 (N_4603,N_4518,N_4544);
xnor U4604 (N_4604,N_4549,N_4501);
nand U4605 (N_4605,N_4531,N_4515);
nor U4606 (N_4606,N_4529,N_4586);
or U4607 (N_4607,N_4588,N_4516);
nor U4608 (N_4608,N_4576,N_4534);
xor U4609 (N_4609,N_4537,N_4507);
nand U4610 (N_4610,N_4597,N_4536);
or U4611 (N_4611,N_4567,N_4509);
and U4612 (N_4612,N_4522,N_4592);
xor U4613 (N_4613,N_4559,N_4506);
nor U4614 (N_4614,N_4551,N_4572);
or U4615 (N_4615,N_4532,N_4526);
and U4616 (N_4616,N_4517,N_4571);
or U4617 (N_4617,N_4505,N_4595);
or U4618 (N_4618,N_4574,N_4573);
nor U4619 (N_4619,N_4543,N_4520);
nand U4620 (N_4620,N_4599,N_4528);
nand U4621 (N_4621,N_4557,N_4555);
and U4622 (N_4622,N_4596,N_4589);
nor U4623 (N_4623,N_4569,N_4565);
nor U4624 (N_4624,N_4550,N_4538);
xor U4625 (N_4625,N_4547,N_4587);
or U4626 (N_4626,N_4580,N_4584);
nand U4627 (N_4627,N_4502,N_4560);
or U4628 (N_4628,N_4561,N_4521);
and U4629 (N_4629,N_4514,N_4500);
nand U4630 (N_4630,N_4510,N_4554);
nand U4631 (N_4631,N_4579,N_4591);
nand U4632 (N_4632,N_4558,N_4504);
nand U4633 (N_4633,N_4583,N_4548);
and U4634 (N_4634,N_4545,N_4585);
or U4635 (N_4635,N_4593,N_4535);
or U4636 (N_4636,N_4552,N_4542);
or U4637 (N_4637,N_4564,N_4524);
and U4638 (N_4638,N_4570,N_4563);
nor U4639 (N_4639,N_4581,N_4527);
or U4640 (N_4640,N_4590,N_4503);
and U4641 (N_4641,N_4512,N_4556);
xor U4642 (N_4642,N_4525,N_4513);
nor U4643 (N_4643,N_4562,N_4578);
nand U4644 (N_4644,N_4511,N_4539);
or U4645 (N_4645,N_4519,N_4568);
and U4646 (N_4646,N_4508,N_4533);
or U4647 (N_4647,N_4594,N_4541);
or U4648 (N_4648,N_4575,N_4598);
nand U4649 (N_4649,N_4546,N_4530);
or U4650 (N_4650,N_4535,N_4583);
or U4651 (N_4651,N_4577,N_4532);
or U4652 (N_4652,N_4569,N_4591);
nand U4653 (N_4653,N_4574,N_4598);
or U4654 (N_4654,N_4525,N_4504);
xnor U4655 (N_4655,N_4576,N_4569);
or U4656 (N_4656,N_4544,N_4521);
and U4657 (N_4657,N_4509,N_4591);
or U4658 (N_4658,N_4545,N_4587);
nand U4659 (N_4659,N_4594,N_4530);
nor U4660 (N_4660,N_4503,N_4572);
nor U4661 (N_4661,N_4537,N_4531);
nand U4662 (N_4662,N_4595,N_4537);
and U4663 (N_4663,N_4594,N_4538);
xor U4664 (N_4664,N_4532,N_4558);
xnor U4665 (N_4665,N_4513,N_4556);
and U4666 (N_4666,N_4589,N_4564);
or U4667 (N_4667,N_4558,N_4544);
nand U4668 (N_4668,N_4512,N_4528);
xor U4669 (N_4669,N_4593,N_4531);
xnor U4670 (N_4670,N_4536,N_4574);
or U4671 (N_4671,N_4513,N_4558);
nand U4672 (N_4672,N_4570,N_4551);
nand U4673 (N_4673,N_4512,N_4505);
or U4674 (N_4674,N_4561,N_4588);
nand U4675 (N_4675,N_4592,N_4505);
or U4676 (N_4676,N_4596,N_4515);
or U4677 (N_4677,N_4594,N_4535);
and U4678 (N_4678,N_4573,N_4520);
xor U4679 (N_4679,N_4572,N_4579);
xor U4680 (N_4680,N_4599,N_4508);
xor U4681 (N_4681,N_4536,N_4570);
and U4682 (N_4682,N_4523,N_4540);
or U4683 (N_4683,N_4525,N_4536);
nor U4684 (N_4684,N_4596,N_4521);
and U4685 (N_4685,N_4505,N_4502);
nand U4686 (N_4686,N_4557,N_4521);
nor U4687 (N_4687,N_4577,N_4501);
xnor U4688 (N_4688,N_4514,N_4558);
or U4689 (N_4689,N_4512,N_4561);
nor U4690 (N_4690,N_4552,N_4574);
nand U4691 (N_4691,N_4536,N_4530);
xor U4692 (N_4692,N_4585,N_4549);
xor U4693 (N_4693,N_4531,N_4500);
and U4694 (N_4694,N_4541,N_4573);
and U4695 (N_4695,N_4599,N_4541);
and U4696 (N_4696,N_4534,N_4556);
nand U4697 (N_4697,N_4514,N_4594);
xnor U4698 (N_4698,N_4579,N_4538);
nor U4699 (N_4699,N_4590,N_4512);
nor U4700 (N_4700,N_4668,N_4692);
xor U4701 (N_4701,N_4612,N_4679);
and U4702 (N_4702,N_4605,N_4611);
and U4703 (N_4703,N_4644,N_4663);
nor U4704 (N_4704,N_4628,N_4637);
xnor U4705 (N_4705,N_4673,N_4696);
nor U4706 (N_4706,N_4684,N_4689);
or U4707 (N_4707,N_4655,N_4608);
or U4708 (N_4708,N_4650,N_4687);
nor U4709 (N_4709,N_4653,N_4609);
nand U4710 (N_4710,N_4625,N_4613);
and U4711 (N_4711,N_4664,N_4680);
nor U4712 (N_4712,N_4630,N_4669);
xor U4713 (N_4713,N_4616,N_4620);
nand U4714 (N_4714,N_4659,N_4606);
and U4715 (N_4715,N_4670,N_4677);
nand U4716 (N_4716,N_4640,N_4683);
nor U4717 (N_4717,N_4686,N_4615);
or U4718 (N_4718,N_4666,N_4656);
or U4719 (N_4719,N_4646,N_4693);
and U4720 (N_4720,N_4685,N_4649);
xnor U4721 (N_4721,N_4642,N_4602);
xnor U4722 (N_4722,N_4672,N_4629);
and U4723 (N_4723,N_4651,N_4636);
or U4724 (N_4724,N_4676,N_4678);
or U4725 (N_4725,N_4658,N_4662);
xor U4726 (N_4726,N_4635,N_4652);
nor U4727 (N_4727,N_4614,N_4645);
nor U4728 (N_4728,N_4699,N_4648);
or U4729 (N_4729,N_4604,N_4607);
nand U4730 (N_4730,N_4691,N_4698);
xor U4731 (N_4731,N_4694,N_4633);
nor U4732 (N_4732,N_4674,N_4631);
and U4733 (N_4733,N_4621,N_4690);
or U4734 (N_4734,N_4682,N_4619);
xor U4735 (N_4735,N_4654,N_4665);
and U4736 (N_4736,N_4681,N_4618);
and U4737 (N_4737,N_4675,N_4695);
or U4738 (N_4738,N_4617,N_4661);
nand U4739 (N_4739,N_4688,N_4657);
or U4740 (N_4740,N_4603,N_4634);
nand U4741 (N_4741,N_4667,N_4639);
and U4742 (N_4742,N_4671,N_4601);
nand U4743 (N_4743,N_4632,N_4627);
xor U4744 (N_4744,N_4610,N_4647);
nor U4745 (N_4745,N_4641,N_4600);
nor U4746 (N_4746,N_4697,N_4660);
nand U4747 (N_4747,N_4638,N_4643);
xor U4748 (N_4748,N_4626,N_4623);
nand U4749 (N_4749,N_4624,N_4622);
nand U4750 (N_4750,N_4645,N_4610);
nand U4751 (N_4751,N_4634,N_4624);
or U4752 (N_4752,N_4606,N_4623);
xor U4753 (N_4753,N_4665,N_4692);
nand U4754 (N_4754,N_4615,N_4658);
nor U4755 (N_4755,N_4693,N_4696);
and U4756 (N_4756,N_4669,N_4631);
and U4757 (N_4757,N_4611,N_4601);
nand U4758 (N_4758,N_4680,N_4654);
and U4759 (N_4759,N_4643,N_4662);
nor U4760 (N_4760,N_4652,N_4639);
nor U4761 (N_4761,N_4655,N_4677);
nand U4762 (N_4762,N_4685,N_4661);
xor U4763 (N_4763,N_4644,N_4642);
or U4764 (N_4764,N_4677,N_4699);
nand U4765 (N_4765,N_4619,N_4666);
xnor U4766 (N_4766,N_4662,N_4683);
xnor U4767 (N_4767,N_4656,N_4672);
xor U4768 (N_4768,N_4626,N_4647);
or U4769 (N_4769,N_4600,N_4692);
nor U4770 (N_4770,N_4671,N_4677);
or U4771 (N_4771,N_4603,N_4678);
and U4772 (N_4772,N_4683,N_4613);
or U4773 (N_4773,N_4692,N_4655);
and U4774 (N_4774,N_4621,N_4652);
xnor U4775 (N_4775,N_4610,N_4621);
or U4776 (N_4776,N_4666,N_4669);
nand U4777 (N_4777,N_4601,N_4638);
nand U4778 (N_4778,N_4602,N_4692);
xnor U4779 (N_4779,N_4602,N_4629);
nand U4780 (N_4780,N_4622,N_4626);
nand U4781 (N_4781,N_4631,N_4670);
xor U4782 (N_4782,N_4604,N_4697);
nor U4783 (N_4783,N_4602,N_4684);
nor U4784 (N_4784,N_4603,N_4610);
xor U4785 (N_4785,N_4681,N_4640);
xnor U4786 (N_4786,N_4634,N_4630);
nand U4787 (N_4787,N_4654,N_4698);
xnor U4788 (N_4788,N_4666,N_4653);
or U4789 (N_4789,N_4602,N_4656);
nand U4790 (N_4790,N_4686,N_4650);
nand U4791 (N_4791,N_4644,N_4601);
and U4792 (N_4792,N_4660,N_4622);
nor U4793 (N_4793,N_4647,N_4616);
or U4794 (N_4794,N_4698,N_4674);
or U4795 (N_4795,N_4688,N_4668);
nand U4796 (N_4796,N_4604,N_4685);
nand U4797 (N_4797,N_4659,N_4665);
and U4798 (N_4798,N_4666,N_4686);
nor U4799 (N_4799,N_4688,N_4698);
nor U4800 (N_4800,N_4770,N_4736);
nor U4801 (N_4801,N_4784,N_4765);
nor U4802 (N_4802,N_4764,N_4734);
and U4803 (N_4803,N_4769,N_4741);
or U4804 (N_4804,N_4793,N_4711);
nand U4805 (N_4805,N_4754,N_4782);
nand U4806 (N_4806,N_4790,N_4788);
nand U4807 (N_4807,N_4757,N_4773);
or U4808 (N_4808,N_4705,N_4730);
or U4809 (N_4809,N_4727,N_4763);
nand U4810 (N_4810,N_4742,N_4771);
or U4811 (N_4811,N_4749,N_4707);
xor U4812 (N_4812,N_4724,N_4786);
xnor U4813 (N_4813,N_4712,N_4751);
or U4814 (N_4814,N_4789,N_4785);
xnor U4815 (N_4815,N_4746,N_4795);
and U4816 (N_4816,N_4783,N_4768);
xnor U4817 (N_4817,N_4796,N_4761);
xnor U4818 (N_4818,N_4728,N_4723);
nand U4819 (N_4819,N_4703,N_4718);
or U4820 (N_4820,N_4775,N_4731);
nor U4821 (N_4821,N_4762,N_4715);
nand U4822 (N_4822,N_4713,N_4708);
and U4823 (N_4823,N_4774,N_4791);
nor U4824 (N_4824,N_4755,N_4706);
nor U4825 (N_4825,N_4743,N_4759);
nand U4826 (N_4826,N_4722,N_4726);
nand U4827 (N_4827,N_4719,N_4778);
nand U4828 (N_4828,N_4752,N_4702);
or U4829 (N_4829,N_4758,N_4716);
nand U4830 (N_4830,N_4766,N_4777);
and U4831 (N_4831,N_4729,N_4704);
nor U4832 (N_4832,N_4709,N_4720);
or U4833 (N_4833,N_4772,N_4744);
nor U4834 (N_4834,N_4767,N_4794);
nand U4835 (N_4835,N_4747,N_4776);
xnor U4836 (N_4836,N_4700,N_4797);
and U4837 (N_4837,N_4753,N_4721);
nand U4838 (N_4838,N_4735,N_4725);
nor U4839 (N_4839,N_4739,N_4760);
nand U4840 (N_4840,N_4733,N_4714);
xor U4841 (N_4841,N_4737,N_4701);
xnor U4842 (N_4842,N_4799,N_4798);
nor U4843 (N_4843,N_4750,N_4738);
or U4844 (N_4844,N_4745,N_4781);
or U4845 (N_4845,N_4756,N_4748);
or U4846 (N_4846,N_4787,N_4732);
xor U4847 (N_4847,N_4717,N_4792);
xor U4848 (N_4848,N_4780,N_4710);
xnor U4849 (N_4849,N_4779,N_4740);
xnor U4850 (N_4850,N_4793,N_4745);
xnor U4851 (N_4851,N_4725,N_4701);
and U4852 (N_4852,N_4711,N_4753);
nand U4853 (N_4853,N_4793,N_4739);
or U4854 (N_4854,N_4789,N_4727);
nor U4855 (N_4855,N_4744,N_4735);
or U4856 (N_4856,N_4791,N_4726);
nor U4857 (N_4857,N_4795,N_4792);
nand U4858 (N_4858,N_4760,N_4727);
or U4859 (N_4859,N_4785,N_4712);
nand U4860 (N_4860,N_4763,N_4726);
xnor U4861 (N_4861,N_4779,N_4780);
or U4862 (N_4862,N_4792,N_4733);
or U4863 (N_4863,N_4767,N_4754);
nor U4864 (N_4864,N_4709,N_4794);
or U4865 (N_4865,N_4784,N_4719);
xor U4866 (N_4866,N_4724,N_4771);
nand U4867 (N_4867,N_4717,N_4756);
and U4868 (N_4868,N_4755,N_4748);
or U4869 (N_4869,N_4730,N_4741);
nand U4870 (N_4870,N_4792,N_4709);
xor U4871 (N_4871,N_4726,N_4728);
xnor U4872 (N_4872,N_4734,N_4770);
xor U4873 (N_4873,N_4754,N_4736);
or U4874 (N_4874,N_4790,N_4751);
nand U4875 (N_4875,N_4714,N_4771);
or U4876 (N_4876,N_4798,N_4749);
nand U4877 (N_4877,N_4721,N_4790);
nand U4878 (N_4878,N_4740,N_4755);
xor U4879 (N_4879,N_4712,N_4719);
nand U4880 (N_4880,N_4769,N_4795);
nand U4881 (N_4881,N_4725,N_4762);
or U4882 (N_4882,N_4710,N_4757);
xor U4883 (N_4883,N_4767,N_4790);
nand U4884 (N_4884,N_4767,N_4779);
or U4885 (N_4885,N_4786,N_4739);
xor U4886 (N_4886,N_4709,N_4711);
or U4887 (N_4887,N_4745,N_4769);
and U4888 (N_4888,N_4795,N_4741);
xnor U4889 (N_4889,N_4739,N_4737);
nand U4890 (N_4890,N_4790,N_4741);
xor U4891 (N_4891,N_4733,N_4703);
nor U4892 (N_4892,N_4727,N_4770);
nor U4893 (N_4893,N_4774,N_4789);
or U4894 (N_4894,N_4727,N_4783);
xnor U4895 (N_4895,N_4750,N_4704);
or U4896 (N_4896,N_4710,N_4784);
xnor U4897 (N_4897,N_4707,N_4730);
or U4898 (N_4898,N_4760,N_4746);
nand U4899 (N_4899,N_4703,N_4747);
nor U4900 (N_4900,N_4880,N_4810);
xnor U4901 (N_4901,N_4865,N_4848);
nor U4902 (N_4902,N_4889,N_4864);
nand U4903 (N_4903,N_4861,N_4844);
xor U4904 (N_4904,N_4804,N_4892);
and U4905 (N_4905,N_4821,N_4881);
xnor U4906 (N_4906,N_4859,N_4820);
or U4907 (N_4907,N_4825,N_4847);
nand U4908 (N_4908,N_4890,N_4818);
or U4909 (N_4909,N_4877,N_4826);
or U4910 (N_4910,N_4883,N_4805);
or U4911 (N_4911,N_4819,N_4824);
and U4912 (N_4912,N_4840,N_4868);
and U4913 (N_4913,N_4807,N_4841);
nor U4914 (N_4914,N_4802,N_4893);
nor U4915 (N_4915,N_4854,N_4834);
nand U4916 (N_4916,N_4855,N_4835);
or U4917 (N_4917,N_4858,N_4829);
and U4918 (N_4918,N_4851,N_4876);
or U4919 (N_4919,N_4846,N_4856);
and U4920 (N_4920,N_4857,N_4806);
and U4921 (N_4921,N_4872,N_4843);
nand U4922 (N_4922,N_4823,N_4811);
xor U4923 (N_4923,N_4871,N_4866);
and U4924 (N_4924,N_4800,N_4837);
and U4925 (N_4925,N_4845,N_4833);
nand U4926 (N_4926,N_4839,N_4886);
or U4927 (N_4927,N_4814,N_4875);
xor U4928 (N_4928,N_4853,N_4878);
xor U4929 (N_4929,N_4836,N_4812);
nor U4930 (N_4930,N_4838,N_4827);
or U4931 (N_4931,N_4816,N_4832);
xnor U4932 (N_4932,N_4879,N_4899);
nand U4933 (N_4933,N_4867,N_4831);
nor U4934 (N_4934,N_4813,N_4850);
nand U4935 (N_4935,N_4897,N_4849);
nor U4936 (N_4936,N_4896,N_4894);
and U4937 (N_4937,N_4809,N_4842);
xor U4938 (N_4938,N_4898,N_4885);
nor U4939 (N_4939,N_4887,N_4808);
xor U4940 (N_4940,N_4822,N_4895);
xor U4941 (N_4941,N_4852,N_4801);
and U4942 (N_4942,N_4882,N_4863);
and U4943 (N_4943,N_4862,N_4891);
and U4944 (N_4944,N_4888,N_4830);
or U4945 (N_4945,N_4869,N_4817);
nor U4946 (N_4946,N_4884,N_4873);
xor U4947 (N_4947,N_4803,N_4874);
xor U4948 (N_4948,N_4828,N_4870);
xnor U4949 (N_4949,N_4815,N_4860);
and U4950 (N_4950,N_4857,N_4882);
and U4951 (N_4951,N_4899,N_4811);
and U4952 (N_4952,N_4869,N_4816);
nor U4953 (N_4953,N_4840,N_4865);
nand U4954 (N_4954,N_4895,N_4834);
nand U4955 (N_4955,N_4884,N_4823);
and U4956 (N_4956,N_4844,N_4871);
nor U4957 (N_4957,N_4817,N_4872);
or U4958 (N_4958,N_4851,N_4829);
and U4959 (N_4959,N_4896,N_4832);
and U4960 (N_4960,N_4855,N_4828);
nand U4961 (N_4961,N_4843,N_4859);
nor U4962 (N_4962,N_4868,N_4869);
nor U4963 (N_4963,N_4869,N_4873);
nand U4964 (N_4964,N_4852,N_4873);
nand U4965 (N_4965,N_4873,N_4889);
and U4966 (N_4966,N_4828,N_4833);
xnor U4967 (N_4967,N_4855,N_4824);
or U4968 (N_4968,N_4836,N_4889);
and U4969 (N_4969,N_4896,N_4836);
nor U4970 (N_4970,N_4852,N_4851);
nor U4971 (N_4971,N_4883,N_4843);
nor U4972 (N_4972,N_4845,N_4819);
nand U4973 (N_4973,N_4814,N_4809);
and U4974 (N_4974,N_4833,N_4805);
and U4975 (N_4975,N_4826,N_4867);
nor U4976 (N_4976,N_4862,N_4858);
xor U4977 (N_4977,N_4841,N_4882);
xnor U4978 (N_4978,N_4824,N_4820);
and U4979 (N_4979,N_4881,N_4887);
or U4980 (N_4980,N_4857,N_4805);
or U4981 (N_4981,N_4867,N_4836);
nand U4982 (N_4982,N_4865,N_4825);
and U4983 (N_4983,N_4839,N_4867);
xnor U4984 (N_4984,N_4877,N_4847);
nor U4985 (N_4985,N_4881,N_4897);
nor U4986 (N_4986,N_4886,N_4880);
xnor U4987 (N_4987,N_4892,N_4829);
nor U4988 (N_4988,N_4859,N_4897);
and U4989 (N_4989,N_4858,N_4881);
nor U4990 (N_4990,N_4881,N_4832);
nor U4991 (N_4991,N_4834,N_4836);
and U4992 (N_4992,N_4848,N_4898);
xor U4993 (N_4993,N_4827,N_4816);
xnor U4994 (N_4994,N_4809,N_4847);
nand U4995 (N_4995,N_4885,N_4817);
xor U4996 (N_4996,N_4823,N_4831);
nor U4997 (N_4997,N_4881,N_4807);
and U4998 (N_4998,N_4883,N_4833);
or U4999 (N_4999,N_4844,N_4807);
nand U5000 (N_5000,N_4920,N_4990);
or U5001 (N_5001,N_4983,N_4937);
and U5002 (N_5002,N_4930,N_4948);
or U5003 (N_5003,N_4952,N_4975);
or U5004 (N_5004,N_4944,N_4905);
nor U5005 (N_5005,N_4909,N_4996);
xnor U5006 (N_5006,N_4982,N_4929);
xnor U5007 (N_5007,N_4907,N_4999);
nand U5008 (N_5008,N_4946,N_4991);
nand U5009 (N_5009,N_4973,N_4914);
and U5010 (N_5010,N_4970,N_4932);
xnor U5011 (N_5011,N_4960,N_4961);
nand U5012 (N_5012,N_4969,N_4945);
nand U5013 (N_5013,N_4979,N_4962);
or U5014 (N_5014,N_4994,N_4919);
nor U5015 (N_5015,N_4998,N_4916);
xor U5016 (N_5016,N_4935,N_4939);
or U5017 (N_5017,N_4908,N_4958);
and U5018 (N_5018,N_4957,N_4917);
nor U5019 (N_5019,N_4931,N_4906);
nand U5020 (N_5020,N_4995,N_4951);
xnor U5021 (N_5021,N_4940,N_4978);
nor U5022 (N_5022,N_4925,N_4943);
or U5023 (N_5023,N_4986,N_4976);
nand U5024 (N_5024,N_4984,N_4934);
nor U5025 (N_5025,N_4968,N_4959);
xnor U5026 (N_5026,N_4910,N_4923);
or U5027 (N_5027,N_4989,N_4933);
and U5028 (N_5028,N_4963,N_4936);
or U5029 (N_5029,N_4922,N_4942);
and U5030 (N_5030,N_4953,N_4950);
nor U5031 (N_5031,N_4904,N_4918);
and U5032 (N_5032,N_4955,N_4985);
nor U5033 (N_5033,N_4941,N_4902);
xnor U5034 (N_5034,N_4947,N_4993);
xnor U5035 (N_5035,N_4924,N_4965);
or U5036 (N_5036,N_4900,N_4981);
nand U5037 (N_5037,N_4987,N_4921);
and U5038 (N_5038,N_4980,N_4992);
or U5039 (N_5039,N_4926,N_4964);
nor U5040 (N_5040,N_4928,N_4901);
and U5041 (N_5041,N_4997,N_4949);
xnor U5042 (N_5042,N_4967,N_4938);
nor U5043 (N_5043,N_4977,N_4903);
or U5044 (N_5044,N_4915,N_4927);
xnor U5045 (N_5045,N_4971,N_4988);
xnor U5046 (N_5046,N_4954,N_4966);
and U5047 (N_5047,N_4974,N_4913);
nor U5048 (N_5048,N_4956,N_4911);
or U5049 (N_5049,N_4912,N_4972);
xor U5050 (N_5050,N_4994,N_4951);
or U5051 (N_5051,N_4936,N_4941);
and U5052 (N_5052,N_4918,N_4920);
nand U5053 (N_5053,N_4909,N_4968);
or U5054 (N_5054,N_4907,N_4943);
and U5055 (N_5055,N_4909,N_4956);
xor U5056 (N_5056,N_4975,N_4941);
or U5057 (N_5057,N_4909,N_4972);
and U5058 (N_5058,N_4944,N_4952);
nand U5059 (N_5059,N_4902,N_4947);
or U5060 (N_5060,N_4991,N_4967);
and U5061 (N_5061,N_4976,N_4972);
or U5062 (N_5062,N_4923,N_4981);
nand U5063 (N_5063,N_4995,N_4901);
nand U5064 (N_5064,N_4989,N_4932);
and U5065 (N_5065,N_4924,N_4930);
nor U5066 (N_5066,N_4992,N_4905);
nand U5067 (N_5067,N_4978,N_4997);
or U5068 (N_5068,N_4900,N_4906);
nand U5069 (N_5069,N_4960,N_4915);
xor U5070 (N_5070,N_4942,N_4999);
nand U5071 (N_5071,N_4995,N_4964);
nor U5072 (N_5072,N_4922,N_4974);
xnor U5073 (N_5073,N_4949,N_4977);
and U5074 (N_5074,N_4930,N_4955);
nand U5075 (N_5075,N_4989,N_4922);
or U5076 (N_5076,N_4946,N_4953);
xnor U5077 (N_5077,N_4961,N_4985);
nor U5078 (N_5078,N_4938,N_4968);
nor U5079 (N_5079,N_4979,N_4943);
or U5080 (N_5080,N_4949,N_4946);
nor U5081 (N_5081,N_4970,N_4964);
and U5082 (N_5082,N_4975,N_4998);
or U5083 (N_5083,N_4939,N_4902);
xor U5084 (N_5084,N_4964,N_4905);
and U5085 (N_5085,N_4950,N_4957);
nor U5086 (N_5086,N_4904,N_4909);
xnor U5087 (N_5087,N_4985,N_4982);
xnor U5088 (N_5088,N_4938,N_4972);
nand U5089 (N_5089,N_4974,N_4944);
nor U5090 (N_5090,N_4906,N_4903);
xnor U5091 (N_5091,N_4909,N_4969);
xor U5092 (N_5092,N_4938,N_4961);
or U5093 (N_5093,N_4997,N_4971);
nor U5094 (N_5094,N_4989,N_4963);
nand U5095 (N_5095,N_4979,N_4987);
xnor U5096 (N_5096,N_4900,N_4930);
and U5097 (N_5097,N_4911,N_4947);
and U5098 (N_5098,N_4997,N_4917);
nand U5099 (N_5099,N_4992,N_4935);
nand U5100 (N_5100,N_5075,N_5086);
nand U5101 (N_5101,N_5036,N_5082);
or U5102 (N_5102,N_5023,N_5094);
xnor U5103 (N_5103,N_5032,N_5038);
xnor U5104 (N_5104,N_5051,N_5029);
nand U5105 (N_5105,N_5045,N_5062);
xor U5106 (N_5106,N_5009,N_5002);
or U5107 (N_5107,N_5054,N_5074);
nand U5108 (N_5108,N_5056,N_5013);
and U5109 (N_5109,N_5070,N_5060);
nor U5110 (N_5110,N_5021,N_5090);
xnor U5111 (N_5111,N_5037,N_5025);
or U5112 (N_5112,N_5006,N_5096);
nor U5113 (N_5113,N_5011,N_5080);
or U5114 (N_5114,N_5088,N_5085);
or U5115 (N_5115,N_5053,N_5014);
or U5116 (N_5116,N_5039,N_5077);
and U5117 (N_5117,N_5018,N_5043);
or U5118 (N_5118,N_5015,N_5065);
xor U5119 (N_5119,N_5026,N_5098);
and U5120 (N_5120,N_5020,N_5034);
and U5121 (N_5121,N_5050,N_5059);
or U5122 (N_5122,N_5027,N_5007);
or U5123 (N_5123,N_5099,N_5000);
or U5124 (N_5124,N_5068,N_5005);
or U5125 (N_5125,N_5010,N_5008);
and U5126 (N_5126,N_5004,N_5024);
and U5127 (N_5127,N_5089,N_5061);
nor U5128 (N_5128,N_5063,N_5072);
or U5129 (N_5129,N_5041,N_5044);
or U5130 (N_5130,N_5092,N_5012);
xnor U5131 (N_5131,N_5001,N_5071);
nor U5132 (N_5132,N_5087,N_5067);
nand U5133 (N_5133,N_5022,N_5079);
nand U5134 (N_5134,N_5093,N_5033);
or U5135 (N_5135,N_5076,N_5083);
nor U5136 (N_5136,N_5081,N_5057);
nand U5137 (N_5137,N_5028,N_5048);
nor U5138 (N_5138,N_5049,N_5066);
or U5139 (N_5139,N_5052,N_5040);
xnor U5140 (N_5140,N_5003,N_5046);
xnor U5141 (N_5141,N_5035,N_5030);
nor U5142 (N_5142,N_5073,N_5091);
and U5143 (N_5143,N_5069,N_5095);
nor U5144 (N_5144,N_5058,N_5055);
nor U5145 (N_5145,N_5019,N_5042);
or U5146 (N_5146,N_5031,N_5016);
nor U5147 (N_5147,N_5047,N_5017);
nand U5148 (N_5148,N_5078,N_5064);
nand U5149 (N_5149,N_5097,N_5084);
and U5150 (N_5150,N_5074,N_5096);
nor U5151 (N_5151,N_5087,N_5090);
nand U5152 (N_5152,N_5087,N_5047);
nand U5153 (N_5153,N_5059,N_5093);
nor U5154 (N_5154,N_5048,N_5046);
or U5155 (N_5155,N_5091,N_5019);
nor U5156 (N_5156,N_5083,N_5041);
or U5157 (N_5157,N_5023,N_5073);
and U5158 (N_5158,N_5036,N_5098);
xor U5159 (N_5159,N_5053,N_5039);
nor U5160 (N_5160,N_5010,N_5056);
nand U5161 (N_5161,N_5024,N_5035);
and U5162 (N_5162,N_5054,N_5062);
and U5163 (N_5163,N_5082,N_5098);
and U5164 (N_5164,N_5021,N_5072);
nand U5165 (N_5165,N_5064,N_5095);
nand U5166 (N_5166,N_5059,N_5046);
or U5167 (N_5167,N_5051,N_5093);
and U5168 (N_5168,N_5055,N_5022);
nand U5169 (N_5169,N_5037,N_5069);
xor U5170 (N_5170,N_5018,N_5006);
nand U5171 (N_5171,N_5068,N_5027);
nand U5172 (N_5172,N_5090,N_5007);
nor U5173 (N_5173,N_5054,N_5070);
nand U5174 (N_5174,N_5043,N_5030);
and U5175 (N_5175,N_5096,N_5031);
nor U5176 (N_5176,N_5043,N_5088);
nand U5177 (N_5177,N_5072,N_5088);
and U5178 (N_5178,N_5033,N_5031);
nor U5179 (N_5179,N_5045,N_5055);
xor U5180 (N_5180,N_5005,N_5059);
xor U5181 (N_5181,N_5006,N_5069);
xnor U5182 (N_5182,N_5052,N_5060);
and U5183 (N_5183,N_5038,N_5034);
and U5184 (N_5184,N_5095,N_5097);
and U5185 (N_5185,N_5000,N_5089);
xnor U5186 (N_5186,N_5032,N_5071);
and U5187 (N_5187,N_5071,N_5003);
nand U5188 (N_5188,N_5060,N_5093);
xnor U5189 (N_5189,N_5070,N_5011);
or U5190 (N_5190,N_5003,N_5004);
nor U5191 (N_5191,N_5039,N_5057);
and U5192 (N_5192,N_5038,N_5097);
and U5193 (N_5193,N_5032,N_5066);
nor U5194 (N_5194,N_5014,N_5049);
xor U5195 (N_5195,N_5020,N_5098);
xor U5196 (N_5196,N_5043,N_5046);
or U5197 (N_5197,N_5063,N_5098);
xor U5198 (N_5198,N_5087,N_5063);
or U5199 (N_5199,N_5077,N_5021);
nor U5200 (N_5200,N_5160,N_5173);
nand U5201 (N_5201,N_5102,N_5165);
and U5202 (N_5202,N_5142,N_5198);
nor U5203 (N_5203,N_5185,N_5178);
and U5204 (N_5204,N_5134,N_5139);
nand U5205 (N_5205,N_5179,N_5155);
xor U5206 (N_5206,N_5146,N_5113);
nand U5207 (N_5207,N_5111,N_5177);
nand U5208 (N_5208,N_5121,N_5192);
nor U5209 (N_5209,N_5125,N_5123);
nand U5210 (N_5210,N_5144,N_5130);
nand U5211 (N_5211,N_5105,N_5137);
nand U5212 (N_5212,N_5110,N_5176);
nand U5213 (N_5213,N_5116,N_5157);
or U5214 (N_5214,N_5104,N_5145);
nor U5215 (N_5215,N_5147,N_5181);
or U5216 (N_5216,N_5184,N_5101);
xnor U5217 (N_5217,N_5191,N_5107);
nor U5218 (N_5218,N_5168,N_5100);
or U5219 (N_5219,N_5106,N_5141);
or U5220 (N_5220,N_5182,N_5136);
and U5221 (N_5221,N_5162,N_5149);
xnor U5222 (N_5222,N_5128,N_5131);
xnor U5223 (N_5223,N_5124,N_5156);
xor U5224 (N_5224,N_5186,N_5174);
or U5225 (N_5225,N_5195,N_5135);
xnor U5226 (N_5226,N_5154,N_5189);
and U5227 (N_5227,N_5127,N_5197);
xor U5228 (N_5228,N_5148,N_5140);
or U5229 (N_5229,N_5150,N_5159);
and U5230 (N_5230,N_5167,N_5193);
xnor U5231 (N_5231,N_5151,N_5108);
xor U5232 (N_5232,N_5172,N_5163);
and U5233 (N_5233,N_5129,N_5194);
nor U5234 (N_5234,N_5120,N_5199);
and U5235 (N_5235,N_5112,N_5164);
xnor U5236 (N_5236,N_5175,N_5169);
or U5237 (N_5237,N_5161,N_5166);
nand U5238 (N_5238,N_5152,N_5188);
or U5239 (N_5239,N_5114,N_5133);
nor U5240 (N_5240,N_5117,N_5103);
nor U5241 (N_5241,N_5187,N_5190);
or U5242 (N_5242,N_5126,N_5132);
and U5243 (N_5243,N_5143,N_5109);
nor U5244 (N_5244,N_5153,N_5180);
xnor U5245 (N_5245,N_5118,N_5158);
nor U5246 (N_5246,N_5119,N_5171);
nand U5247 (N_5247,N_5183,N_5115);
nor U5248 (N_5248,N_5196,N_5122);
or U5249 (N_5249,N_5170,N_5138);
nand U5250 (N_5250,N_5133,N_5167);
and U5251 (N_5251,N_5168,N_5194);
xnor U5252 (N_5252,N_5113,N_5197);
nand U5253 (N_5253,N_5191,N_5119);
nand U5254 (N_5254,N_5145,N_5171);
nor U5255 (N_5255,N_5198,N_5168);
or U5256 (N_5256,N_5195,N_5158);
nand U5257 (N_5257,N_5129,N_5164);
nand U5258 (N_5258,N_5162,N_5157);
xnor U5259 (N_5259,N_5184,N_5129);
and U5260 (N_5260,N_5107,N_5149);
and U5261 (N_5261,N_5199,N_5197);
nand U5262 (N_5262,N_5139,N_5151);
xor U5263 (N_5263,N_5140,N_5193);
nand U5264 (N_5264,N_5191,N_5126);
or U5265 (N_5265,N_5160,N_5120);
or U5266 (N_5266,N_5154,N_5176);
and U5267 (N_5267,N_5196,N_5193);
nor U5268 (N_5268,N_5166,N_5187);
or U5269 (N_5269,N_5146,N_5127);
or U5270 (N_5270,N_5124,N_5176);
xnor U5271 (N_5271,N_5135,N_5180);
and U5272 (N_5272,N_5105,N_5184);
nand U5273 (N_5273,N_5198,N_5116);
nor U5274 (N_5274,N_5185,N_5123);
xnor U5275 (N_5275,N_5106,N_5111);
xor U5276 (N_5276,N_5198,N_5149);
nor U5277 (N_5277,N_5119,N_5120);
and U5278 (N_5278,N_5197,N_5166);
and U5279 (N_5279,N_5164,N_5160);
nor U5280 (N_5280,N_5196,N_5101);
xor U5281 (N_5281,N_5159,N_5153);
or U5282 (N_5282,N_5130,N_5176);
xnor U5283 (N_5283,N_5122,N_5194);
nor U5284 (N_5284,N_5197,N_5107);
and U5285 (N_5285,N_5151,N_5181);
or U5286 (N_5286,N_5139,N_5175);
or U5287 (N_5287,N_5120,N_5150);
nand U5288 (N_5288,N_5198,N_5128);
nor U5289 (N_5289,N_5177,N_5113);
nor U5290 (N_5290,N_5191,N_5140);
xor U5291 (N_5291,N_5197,N_5156);
nor U5292 (N_5292,N_5103,N_5165);
xor U5293 (N_5293,N_5179,N_5180);
and U5294 (N_5294,N_5182,N_5124);
nand U5295 (N_5295,N_5135,N_5169);
or U5296 (N_5296,N_5117,N_5150);
nor U5297 (N_5297,N_5159,N_5110);
or U5298 (N_5298,N_5130,N_5113);
nand U5299 (N_5299,N_5172,N_5146);
nand U5300 (N_5300,N_5285,N_5234);
nand U5301 (N_5301,N_5240,N_5226);
and U5302 (N_5302,N_5213,N_5261);
xnor U5303 (N_5303,N_5265,N_5210);
xnor U5304 (N_5304,N_5294,N_5279);
nor U5305 (N_5305,N_5286,N_5263);
and U5306 (N_5306,N_5281,N_5217);
nor U5307 (N_5307,N_5298,N_5223);
and U5308 (N_5308,N_5266,N_5244);
or U5309 (N_5309,N_5274,N_5258);
or U5310 (N_5310,N_5260,N_5253);
or U5311 (N_5311,N_5252,N_5264);
nor U5312 (N_5312,N_5251,N_5299);
nand U5313 (N_5313,N_5228,N_5224);
and U5314 (N_5314,N_5229,N_5201);
xor U5315 (N_5315,N_5225,N_5259);
nor U5316 (N_5316,N_5297,N_5256);
and U5317 (N_5317,N_5248,N_5211);
and U5318 (N_5318,N_5236,N_5232);
xor U5319 (N_5319,N_5269,N_5241);
nor U5320 (N_5320,N_5222,N_5289);
xor U5321 (N_5321,N_5200,N_5245);
and U5322 (N_5322,N_5204,N_5278);
nor U5323 (N_5323,N_5207,N_5267);
xor U5324 (N_5324,N_5268,N_5250);
nor U5325 (N_5325,N_5288,N_5219);
or U5326 (N_5326,N_5276,N_5202);
and U5327 (N_5327,N_5221,N_5218);
nand U5328 (N_5328,N_5280,N_5214);
xnor U5329 (N_5329,N_5243,N_5249);
nor U5330 (N_5330,N_5292,N_5215);
or U5331 (N_5331,N_5233,N_5247);
or U5332 (N_5332,N_5295,N_5231);
and U5333 (N_5333,N_5239,N_5203);
or U5334 (N_5334,N_5205,N_5242);
and U5335 (N_5335,N_5212,N_5270);
xor U5336 (N_5336,N_5209,N_5277);
or U5337 (N_5337,N_5275,N_5220);
xor U5338 (N_5338,N_5230,N_5290);
or U5339 (N_5339,N_5262,N_5246);
xnor U5340 (N_5340,N_5238,N_5216);
nor U5341 (N_5341,N_5291,N_5293);
xor U5342 (N_5342,N_5227,N_5296);
xor U5343 (N_5343,N_5237,N_5282);
nor U5344 (N_5344,N_5254,N_5283);
and U5345 (N_5345,N_5255,N_5206);
or U5346 (N_5346,N_5235,N_5273);
xor U5347 (N_5347,N_5287,N_5257);
nor U5348 (N_5348,N_5284,N_5271);
nor U5349 (N_5349,N_5208,N_5272);
and U5350 (N_5350,N_5243,N_5209);
or U5351 (N_5351,N_5255,N_5213);
nor U5352 (N_5352,N_5200,N_5211);
or U5353 (N_5353,N_5234,N_5236);
and U5354 (N_5354,N_5204,N_5283);
or U5355 (N_5355,N_5267,N_5209);
or U5356 (N_5356,N_5222,N_5245);
xor U5357 (N_5357,N_5273,N_5277);
nand U5358 (N_5358,N_5266,N_5260);
or U5359 (N_5359,N_5247,N_5263);
xnor U5360 (N_5360,N_5204,N_5228);
xor U5361 (N_5361,N_5203,N_5281);
xnor U5362 (N_5362,N_5290,N_5284);
and U5363 (N_5363,N_5234,N_5215);
and U5364 (N_5364,N_5219,N_5233);
nor U5365 (N_5365,N_5222,N_5292);
and U5366 (N_5366,N_5258,N_5208);
nand U5367 (N_5367,N_5261,N_5217);
and U5368 (N_5368,N_5244,N_5291);
nor U5369 (N_5369,N_5293,N_5265);
and U5370 (N_5370,N_5219,N_5255);
xnor U5371 (N_5371,N_5238,N_5272);
or U5372 (N_5372,N_5282,N_5205);
nand U5373 (N_5373,N_5220,N_5277);
nand U5374 (N_5374,N_5224,N_5249);
xnor U5375 (N_5375,N_5273,N_5230);
or U5376 (N_5376,N_5268,N_5247);
or U5377 (N_5377,N_5239,N_5249);
nor U5378 (N_5378,N_5247,N_5291);
nor U5379 (N_5379,N_5280,N_5273);
nand U5380 (N_5380,N_5237,N_5235);
and U5381 (N_5381,N_5239,N_5228);
xor U5382 (N_5382,N_5219,N_5272);
nor U5383 (N_5383,N_5277,N_5230);
and U5384 (N_5384,N_5281,N_5257);
and U5385 (N_5385,N_5203,N_5209);
nand U5386 (N_5386,N_5289,N_5259);
or U5387 (N_5387,N_5249,N_5246);
and U5388 (N_5388,N_5217,N_5246);
xnor U5389 (N_5389,N_5203,N_5205);
and U5390 (N_5390,N_5243,N_5247);
and U5391 (N_5391,N_5247,N_5200);
and U5392 (N_5392,N_5277,N_5226);
nand U5393 (N_5393,N_5212,N_5242);
nand U5394 (N_5394,N_5252,N_5214);
nand U5395 (N_5395,N_5245,N_5292);
nor U5396 (N_5396,N_5202,N_5285);
nor U5397 (N_5397,N_5284,N_5235);
or U5398 (N_5398,N_5296,N_5226);
nor U5399 (N_5399,N_5286,N_5226);
nand U5400 (N_5400,N_5321,N_5306);
nor U5401 (N_5401,N_5319,N_5324);
nor U5402 (N_5402,N_5367,N_5300);
and U5403 (N_5403,N_5384,N_5332);
xor U5404 (N_5404,N_5337,N_5360);
nor U5405 (N_5405,N_5342,N_5318);
nand U5406 (N_5406,N_5343,N_5316);
or U5407 (N_5407,N_5315,N_5341);
nor U5408 (N_5408,N_5390,N_5383);
and U5409 (N_5409,N_5350,N_5377);
xor U5410 (N_5410,N_5355,N_5344);
and U5411 (N_5411,N_5331,N_5352);
and U5412 (N_5412,N_5326,N_5354);
nor U5413 (N_5413,N_5312,N_5361);
xor U5414 (N_5414,N_5363,N_5386);
nor U5415 (N_5415,N_5373,N_5393);
and U5416 (N_5416,N_5330,N_5339);
nor U5417 (N_5417,N_5357,N_5317);
nand U5418 (N_5418,N_5307,N_5385);
nor U5419 (N_5419,N_5309,N_5380);
nor U5420 (N_5420,N_5392,N_5314);
xnor U5421 (N_5421,N_5310,N_5388);
or U5422 (N_5422,N_5302,N_5334);
nand U5423 (N_5423,N_5372,N_5340);
xnor U5424 (N_5424,N_5327,N_5305);
xnor U5425 (N_5425,N_5378,N_5304);
and U5426 (N_5426,N_5325,N_5336);
nand U5427 (N_5427,N_5370,N_5351);
nor U5428 (N_5428,N_5313,N_5381);
nor U5429 (N_5429,N_5374,N_5328);
or U5430 (N_5430,N_5308,N_5396);
and U5431 (N_5431,N_5397,N_5391);
nand U5432 (N_5432,N_5329,N_5322);
nor U5433 (N_5433,N_5358,N_5366);
nand U5434 (N_5434,N_5356,N_5395);
xor U5435 (N_5435,N_5382,N_5398);
nand U5436 (N_5436,N_5368,N_5365);
nor U5437 (N_5437,N_5389,N_5353);
xor U5438 (N_5438,N_5362,N_5338);
nand U5439 (N_5439,N_5347,N_5349);
xnor U5440 (N_5440,N_5320,N_5359);
or U5441 (N_5441,N_5399,N_5379);
nor U5442 (N_5442,N_5345,N_5303);
xnor U5443 (N_5443,N_5301,N_5311);
or U5444 (N_5444,N_5371,N_5323);
or U5445 (N_5445,N_5394,N_5364);
or U5446 (N_5446,N_5348,N_5387);
or U5447 (N_5447,N_5346,N_5376);
nor U5448 (N_5448,N_5375,N_5333);
and U5449 (N_5449,N_5335,N_5369);
xor U5450 (N_5450,N_5320,N_5395);
or U5451 (N_5451,N_5386,N_5354);
or U5452 (N_5452,N_5357,N_5380);
and U5453 (N_5453,N_5348,N_5347);
or U5454 (N_5454,N_5342,N_5382);
nand U5455 (N_5455,N_5385,N_5367);
or U5456 (N_5456,N_5331,N_5361);
nor U5457 (N_5457,N_5339,N_5360);
nor U5458 (N_5458,N_5373,N_5300);
nand U5459 (N_5459,N_5380,N_5320);
nor U5460 (N_5460,N_5310,N_5300);
xor U5461 (N_5461,N_5311,N_5378);
nand U5462 (N_5462,N_5371,N_5306);
nor U5463 (N_5463,N_5353,N_5305);
and U5464 (N_5464,N_5394,N_5389);
or U5465 (N_5465,N_5329,N_5383);
nand U5466 (N_5466,N_5300,N_5366);
and U5467 (N_5467,N_5336,N_5323);
nor U5468 (N_5468,N_5330,N_5327);
and U5469 (N_5469,N_5351,N_5347);
nand U5470 (N_5470,N_5342,N_5344);
xor U5471 (N_5471,N_5383,N_5325);
nand U5472 (N_5472,N_5351,N_5312);
and U5473 (N_5473,N_5391,N_5390);
or U5474 (N_5474,N_5387,N_5367);
and U5475 (N_5475,N_5341,N_5396);
and U5476 (N_5476,N_5344,N_5359);
or U5477 (N_5477,N_5377,N_5371);
nor U5478 (N_5478,N_5396,N_5379);
nor U5479 (N_5479,N_5308,N_5324);
or U5480 (N_5480,N_5373,N_5347);
nand U5481 (N_5481,N_5350,N_5385);
nor U5482 (N_5482,N_5307,N_5384);
nor U5483 (N_5483,N_5365,N_5377);
or U5484 (N_5484,N_5354,N_5358);
or U5485 (N_5485,N_5395,N_5384);
nand U5486 (N_5486,N_5360,N_5364);
nor U5487 (N_5487,N_5351,N_5313);
or U5488 (N_5488,N_5360,N_5385);
xnor U5489 (N_5489,N_5381,N_5312);
nor U5490 (N_5490,N_5363,N_5335);
or U5491 (N_5491,N_5372,N_5355);
nor U5492 (N_5492,N_5392,N_5359);
and U5493 (N_5493,N_5352,N_5311);
xor U5494 (N_5494,N_5391,N_5389);
xor U5495 (N_5495,N_5399,N_5315);
nor U5496 (N_5496,N_5358,N_5367);
nand U5497 (N_5497,N_5340,N_5332);
or U5498 (N_5498,N_5361,N_5304);
nor U5499 (N_5499,N_5339,N_5300);
or U5500 (N_5500,N_5450,N_5452);
or U5501 (N_5501,N_5463,N_5462);
and U5502 (N_5502,N_5438,N_5408);
nor U5503 (N_5503,N_5440,N_5429);
nor U5504 (N_5504,N_5471,N_5489);
and U5505 (N_5505,N_5457,N_5401);
nand U5506 (N_5506,N_5494,N_5496);
xor U5507 (N_5507,N_5477,N_5424);
and U5508 (N_5508,N_5409,N_5407);
xor U5509 (N_5509,N_5479,N_5485);
xor U5510 (N_5510,N_5448,N_5447);
nand U5511 (N_5511,N_5483,N_5406);
nand U5512 (N_5512,N_5439,N_5473);
or U5513 (N_5513,N_5459,N_5419);
nand U5514 (N_5514,N_5418,N_5443);
xor U5515 (N_5515,N_5492,N_5461);
and U5516 (N_5516,N_5468,N_5414);
nand U5517 (N_5517,N_5458,N_5474);
nor U5518 (N_5518,N_5488,N_5495);
and U5519 (N_5519,N_5469,N_5432);
or U5520 (N_5520,N_5436,N_5491);
nor U5521 (N_5521,N_5405,N_5430);
or U5522 (N_5522,N_5472,N_5410);
xor U5523 (N_5523,N_5478,N_5434);
nor U5524 (N_5524,N_5465,N_5423);
and U5525 (N_5525,N_5415,N_5453);
and U5526 (N_5526,N_5411,N_5428);
nand U5527 (N_5527,N_5451,N_5446);
or U5528 (N_5528,N_5404,N_5420);
or U5529 (N_5529,N_5487,N_5466);
nor U5530 (N_5530,N_5490,N_5426);
nor U5531 (N_5531,N_5437,N_5422);
nor U5532 (N_5532,N_5425,N_5435);
and U5533 (N_5533,N_5416,N_5484);
xnor U5534 (N_5534,N_5412,N_5456);
nand U5535 (N_5535,N_5476,N_5431);
nand U5536 (N_5536,N_5493,N_5499);
nor U5537 (N_5537,N_5417,N_5486);
and U5538 (N_5538,N_5475,N_5470);
and U5539 (N_5539,N_5400,N_5449);
and U5540 (N_5540,N_5480,N_5421);
and U5541 (N_5541,N_5413,N_5464);
nand U5542 (N_5542,N_5445,N_5498);
nor U5543 (N_5543,N_5455,N_5403);
or U5544 (N_5544,N_5433,N_5444);
xor U5545 (N_5545,N_5481,N_5442);
or U5546 (N_5546,N_5497,N_5402);
and U5547 (N_5547,N_5460,N_5454);
nand U5548 (N_5548,N_5467,N_5482);
xor U5549 (N_5549,N_5441,N_5427);
nor U5550 (N_5550,N_5435,N_5420);
xnor U5551 (N_5551,N_5436,N_5472);
nor U5552 (N_5552,N_5449,N_5407);
xor U5553 (N_5553,N_5442,N_5446);
nor U5554 (N_5554,N_5414,N_5493);
or U5555 (N_5555,N_5400,N_5407);
nand U5556 (N_5556,N_5433,N_5496);
and U5557 (N_5557,N_5406,N_5468);
or U5558 (N_5558,N_5466,N_5402);
xnor U5559 (N_5559,N_5457,N_5492);
nand U5560 (N_5560,N_5413,N_5474);
nand U5561 (N_5561,N_5490,N_5477);
xor U5562 (N_5562,N_5435,N_5472);
nor U5563 (N_5563,N_5432,N_5438);
or U5564 (N_5564,N_5460,N_5455);
nand U5565 (N_5565,N_5438,N_5414);
or U5566 (N_5566,N_5404,N_5428);
or U5567 (N_5567,N_5418,N_5414);
xnor U5568 (N_5568,N_5493,N_5403);
xnor U5569 (N_5569,N_5447,N_5475);
nor U5570 (N_5570,N_5442,N_5478);
nor U5571 (N_5571,N_5406,N_5436);
nor U5572 (N_5572,N_5462,N_5433);
or U5573 (N_5573,N_5473,N_5478);
xnor U5574 (N_5574,N_5420,N_5412);
nand U5575 (N_5575,N_5478,N_5493);
and U5576 (N_5576,N_5403,N_5458);
xnor U5577 (N_5577,N_5450,N_5484);
or U5578 (N_5578,N_5469,N_5445);
xor U5579 (N_5579,N_5448,N_5481);
and U5580 (N_5580,N_5450,N_5466);
or U5581 (N_5581,N_5499,N_5434);
xor U5582 (N_5582,N_5445,N_5429);
xor U5583 (N_5583,N_5485,N_5421);
xnor U5584 (N_5584,N_5456,N_5453);
xor U5585 (N_5585,N_5421,N_5475);
xor U5586 (N_5586,N_5423,N_5490);
xnor U5587 (N_5587,N_5494,N_5483);
and U5588 (N_5588,N_5448,N_5406);
nor U5589 (N_5589,N_5415,N_5467);
nand U5590 (N_5590,N_5461,N_5464);
nand U5591 (N_5591,N_5409,N_5430);
and U5592 (N_5592,N_5455,N_5491);
xnor U5593 (N_5593,N_5460,N_5417);
or U5594 (N_5594,N_5422,N_5414);
xor U5595 (N_5595,N_5411,N_5433);
and U5596 (N_5596,N_5477,N_5407);
xnor U5597 (N_5597,N_5402,N_5448);
or U5598 (N_5598,N_5465,N_5400);
and U5599 (N_5599,N_5475,N_5451);
nor U5600 (N_5600,N_5578,N_5519);
and U5601 (N_5601,N_5543,N_5517);
xor U5602 (N_5602,N_5524,N_5564);
and U5603 (N_5603,N_5566,N_5588);
nand U5604 (N_5604,N_5551,N_5509);
or U5605 (N_5605,N_5529,N_5571);
nand U5606 (N_5606,N_5553,N_5514);
nand U5607 (N_5607,N_5504,N_5544);
or U5608 (N_5608,N_5542,N_5516);
or U5609 (N_5609,N_5550,N_5510);
xnor U5610 (N_5610,N_5523,N_5592);
xor U5611 (N_5611,N_5556,N_5573);
nand U5612 (N_5612,N_5557,N_5535);
and U5613 (N_5613,N_5552,N_5503);
and U5614 (N_5614,N_5549,N_5540);
nand U5615 (N_5615,N_5568,N_5539);
nand U5616 (N_5616,N_5545,N_5558);
nand U5617 (N_5617,N_5548,N_5528);
nand U5618 (N_5618,N_5563,N_5595);
xor U5619 (N_5619,N_5508,N_5541);
nand U5620 (N_5620,N_5527,N_5534);
xor U5621 (N_5621,N_5512,N_5507);
nand U5622 (N_5622,N_5582,N_5526);
nand U5623 (N_5623,N_5505,N_5532);
nand U5624 (N_5624,N_5577,N_5502);
xnor U5625 (N_5625,N_5565,N_5594);
or U5626 (N_5626,N_5580,N_5584);
xnor U5627 (N_5627,N_5533,N_5583);
and U5628 (N_5628,N_5547,N_5574);
nand U5629 (N_5629,N_5585,N_5500);
or U5630 (N_5630,N_5569,N_5591);
or U5631 (N_5631,N_5576,N_5593);
xnor U5632 (N_5632,N_5531,N_5598);
nand U5633 (N_5633,N_5596,N_5560);
nor U5634 (N_5634,N_5525,N_5562);
nand U5635 (N_5635,N_5575,N_5567);
and U5636 (N_5636,N_5572,N_5589);
xnor U5637 (N_5637,N_5513,N_5520);
xnor U5638 (N_5638,N_5506,N_5559);
xnor U5639 (N_5639,N_5521,N_5546);
xnor U5640 (N_5640,N_5522,N_5530);
xnor U5641 (N_5641,N_5586,N_5597);
or U5642 (N_5642,N_5536,N_5581);
and U5643 (N_5643,N_5587,N_5590);
and U5644 (N_5644,N_5555,N_5537);
and U5645 (N_5645,N_5599,N_5501);
nand U5646 (N_5646,N_5511,N_5518);
xor U5647 (N_5647,N_5515,N_5579);
and U5648 (N_5648,N_5561,N_5570);
nand U5649 (N_5649,N_5538,N_5554);
xnor U5650 (N_5650,N_5549,N_5575);
xnor U5651 (N_5651,N_5574,N_5592);
nor U5652 (N_5652,N_5502,N_5592);
or U5653 (N_5653,N_5571,N_5570);
or U5654 (N_5654,N_5555,N_5576);
and U5655 (N_5655,N_5588,N_5580);
and U5656 (N_5656,N_5574,N_5552);
nor U5657 (N_5657,N_5501,N_5548);
nand U5658 (N_5658,N_5549,N_5595);
nand U5659 (N_5659,N_5597,N_5510);
nor U5660 (N_5660,N_5588,N_5555);
nor U5661 (N_5661,N_5507,N_5531);
nand U5662 (N_5662,N_5559,N_5515);
nand U5663 (N_5663,N_5510,N_5505);
and U5664 (N_5664,N_5528,N_5573);
and U5665 (N_5665,N_5519,N_5561);
nor U5666 (N_5666,N_5535,N_5579);
nand U5667 (N_5667,N_5565,N_5529);
nor U5668 (N_5668,N_5543,N_5540);
nand U5669 (N_5669,N_5523,N_5565);
nand U5670 (N_5670,N_5534,N_5500);
and U5671 (N_5671,N_5559,N_5542);
or U5672 (N_5672,N_5582,N_5592);
and U5673 (N_5673,N_5599,N_5532);
xnor U5674 (N_5674,N_5595,N_5555);
or U5675 (N_5675,N_5524,N_5557);
or U5676 (N_5676,N_5527,N_5573);
nor U5677 (N_5677,N_5524,N_5508);
and U5678 (N_5678,N_5558,N_5564);
nand U5679 (N_5679,N_5515,N_5523);
and U5680 (N_5680,N_5592,N_5504);
and U5681 (N_5681,N_5510,N_5543);
nor U5682 (N_5682,N_5596,N_5579);
nand U5683 (N_5683,N_5537,N_5594);
or U5684 (N_5684,N_5592,N_5570);
or U5685 (N_5685,N_5588,N_5514);
nor U5686 (N_5686,N_5507,N_5569);
nand U5687 (N_5687,N_5528,N_5534);
and U5688 (N_5688,N_5592,N_5546);
nand U5689 (N_5689,N_5531,N_5502);
nand U5690 (N_5690,N_5545,N_5511);
nand U5691 (N_5691,N_5500,N_5565);
and U5692 (N_5692,N_5565,N_5585);
and U5693 (N_5693,N_5504,N_5510);
nand U5694 (N_5694,N_5597,N_5537);
nor U5695 (N_5695,N_5548,N_5596);
nand U5696 (N_5696,N_5509,N_5541);
nand U5697 (N_5697,N_5507,N_5508);
or U5698 (N_5698,N_5580,N_5545);
and U5699 (N_5699,N_5507,N_5589);
nand U5700 (N_5700,N_5696,N_5639);
or U5701 (N_5701,N_5681,N_5620);
nor U5702 (N_5702,N_5668,N_5631);
and U5703 (N_5703,N_5601,N_5646);
xnor U5704 (N_5704,N_5687,N_5651);
or U5705 (N_5705,N_5664,N_5606);
xnor U5706 (N_5706,N_5675,N_5649);
xnor U5707 (N_5707,N_5695,N_5641);
nor U5708 (N_5708,N_5636,N_5673);
nand U5709 (N_5709,N_5634,N_5627);
nand U5710 (N_5710,N_5655,N_5604);
nand U5711 (N_5711,N_5629,N_5633);
nand U5712 (N_5712,N_5632,N_5667);
or U5713 (N_5713,N_5659,N_5672);
nand U5714 (N_5714,N_5692,N_5623);
nor U5715 (N_5715,N_5698,N_5607);
nor U5716 (N_5716,N_5615,N_5626);
nand U5717 (N_5717,N_5657,N_5621);
or U5718 (N_5718,N_5622,N_5661);
nand U5719 (N_5719,N_5628,N_5686);
and U5720 (N_5720,N_5652,N_5603);
xnor U5721 (N_5721,N_5650,N_5699);
or U5722 (N_5722,N_5635,N_5637);
and U5723 (N_5723,N_5624,N_5653);
nor U5724 (N_5724,N_5612,N_5658);
or U5725 (N_5725,N_5645,N_5670);
and U5726 (N_5726,N_5647,N_5656);
nand U5727 (N_5727,N_5617,N_5618);
nand U5728 (N_5728,N_5642,N_5654);
nor U5729 (N_5729,N_5676,N_5697);
xor U5730 (N_5730,N_5669,N_5671);
xor U5731 (N_5731,N_5643,N_5663);
or U5732 (N_5732,N_5600,N_5605);
or U5733 (N_5733,N_5640,N_5613);
or U5734 (N_5734,N_5625,N_5666);
or U5735 (N_5735,N_5648,N_5660);
and U5736 (N_5736,N_5682,N_5679);
nor U5737 (N_5737,N_5614,N_5691);
or U5738 (N_5738,N_5674,N_5683);
and U5739 (N_5739,N_5685,N_5693);
and U5740 (N_5740,N_5689,N_5694);
nor U5741 (N_5741,N_5680,N_5638);
nor U5742 (N_5742,N_5690,N_5602);
and U5743 (N_5743,N_5610,N_5677);
xor U5744 (N_5744,N_5619,N_5678);
xor U5745 (N_5745,N_5630,N_5665);
and U5746 (N_5746,N_5616,N_5609);
or U5747 (N_5747,N_5611,N_5608);
or U5748 (N_5748,N_5644,N_5684);
nor U5749 (N_5749,N_5662,N_5688);
nor U5750 (N_5750,N_5604,N_5636);
or U5751 (N_5751,N_5665,N_5655);
nor U5752 (N_5752,N_5646,N_5620);
and U5753 (N_5753,N_5674,N_5686);
or U5754 (N_5754,N_5642,N_5682);
nand U5755 (N_5755,N_5638,N_5652);
nor U5756 (N_5756,N_5658,N_5676);
or U5757 (N_5757,N_5604,N_5630);
nand U5758 (N_5758,N_5646,N_5639);
and U5759 (N_5759,N_5687,N_5658);
nor U5760 (N_5760,N_5613,N_5662);
nor U5761 (N_5761,N_5682,N_5603);
xor U5762 (N_5762,N_5618,N_5616);
xor U5763 (N_5763,N_5688,N_5617);
and U5764 (N_5764,N_5638,N_5649);
xnor U5765 (N_5765,N_5618,N_5647);
nand U5766 (N_5766,N_5683,N_5628);
nand U5767 (N_5767,N_5632,N_5606);
and U5768 (N_5768,N_5624,N_5678);
nor U5769 (N_5769,N_5638,N_5665);
or U5770 (N_5770,N_5605,N_5612);
and U5771 (N_5771,N_5632,N_5611);
nand U5772 (N_5772,N_5604,N_5639);
and U5773 (N_5773,N_5696,N_5628);
nor U5774 (N_5774,N_5665,N_5667);
nand U5775 (N_5775,N_5651,N_5686);
nand U5776 (N_5776,N_5635,N_5663);
nor U5777 (N_5777,N_5658,N_5665);
and U5778 (N_5778,N_5644,N_5650);
or U5779 (N_5779,N_5656,N_5613);
xnor U5780 (N_5780,N_5614,N_5603);
nor U5781 (N_5781,N_5683,N_5692);
xnor U5782 (N_5782,N_5634,N_5661);
xor U5783 (N_5783,N_5678,N_5692);
or U5784 (N_5784,N_5656,N_5648);
xnor U5785 (N_5785,N_5654,N_5634);
and U5786 (N_5786,N_5695,N_5620);
nor U5787 (N_5787,N_5671,N_5652);
nor U5788 (N_5788,N_5689,N_5680);
or U5789 (N_5789,N_5616,N_5614);
or U5790 (N_5790,N_5624,N_5631);
or U5791 (N_5791,N_5603,N_5623);
nor U5792 (N_5792,N_5632,N_5686);
or U5793 (N_5793,N_5664,N_5669);
xor U5794 (N_5794,N_5693,N_5686);
and U5795 (N_5795,N_5618,N_5603);
nor U5796 (N_5796,N_5640,N_5689);
nand U5797 (N_5797,N_5686,N_5629);
nor U5798 (N_5798,N_5697,N_5623);
xor U5799 (N_5799,N_5635,N_5672);
xnor U5800 (N_5800,N_5701,N_5760);
or U5801 (N_5801,N_5783,N_5779);
nor U5802 (N_5802,N_5705,N_5726);
or U5803 (N_5803,N_5741,N_5796);
or U5804 (N_5804,N_5777,N_5743);
nor U5805 (N_5805,N_5757,N_5712);
nand U5806 (N_5806,N_5717,N_5758);
nor U5807 (N_5807,N_5713,N_5710);
and U5808 (N_5808,N_5723,N_5739);
nand U5809 (N_5809,N_5771,N_5750);
xor U5810 (N_5810,N_5788,N_5745);
nor U5811 (N_5811,N_5703,N_5774);
nand U5812 (N_5812,N_5744,N_5700);
and U5813 (N_5813,N_5704,N_5763);
and U5814 (N_5814,N_5715,N_5793);
nand U5815 (N_5815,N_5791,N_5714);
or U5816 (N_5816,N_5786,N_5748);
or U5817 (N_5817,N_5768,N_5759);
xnor U5818 (N_5818,N_5761,N_5719);
nand U5819 (N_5819,N_5747,N_5752);
nand U5820 (N_5820,N_5780,N_5749);
and U5821 (N_5821,N_5732,N_5733);
nor U5822 (N_5822,N_5770,N_5756);
xnor U5823 (N_5823,N_5728,N_5798);
and U5824 (N_5824,N_5792,N_5736);
and U5825 (N_5825,N_5727,N_5799);
or U5826 (N_5826,N_5716,N_5785);
or U5827 (N_5827,N_5797,N_5720);
xnor U5828 (N_5828,N_5735,N_5773);
xor U5829 (N_5829,N_5782,N_5762);
or U5830 (N_5830,N_5746,N_5787);
and U5831 (N_5831,N_5794,N_5775);
and U5832 (N_5832,N_5766,N_5795);
nor U5833 (N_5833,N_5781,N_5724);
and U5834 (N_5834,N_5769,N_5772);
nand U5835 (N_5835,N_5730,N_5731);
nand U5836 (N_5836,N_5742,N_5734);
nand U5837 (N_5837,N_5755,N_5776);
xor U5838 (N_5838,N_5711,N_5738);
and U5839 (N_5839,N_5754,N_5751);
or U5840 (N_5840,N_5764,N_5778);
and U5841 (N_5841,N_5753,N_5718);
xor U5842 (N_5842,N_5789,N_5725);
or U5843 (N_5843,N_5708,N_5790);
or U5844 (N_5844,N_5729,N_5767);
nor U5845 (N_5845,N_5706,N_5740);
xnor U5846 (N_5846,N_5784,N_5721);
nor U5847 (N_5847,N_5702,N_5737);
xor U5848 (N_5848,N_5709,N_5707);
nand U5849 (N_5849,N_5722,N_5765);
or U5850 (N_5850,N_5757,N_5761);
nor U5851 (N_5851,N_5709,N_5755);
nand U5852 (N_5852,N_5740,N_5702);
and U5853 (N_5853,N_5780,N_5741);
nor U5854 (N_5854,N_5739,N_5777);
nor U5855 (N_5855,N_5748,N_5700);
or U5856 (N_5856,N_5793,N_5778);
and U5857 (N_5857,N_5707,N_5765);
or U5858 (N_5858,N_5733,N_5768);
xnor U5859 (N_5859,N_5786,N_5771);
xnor U5860 (N_5860,N_5751,N_5735);
xnor U5861 (N_5861,N_5798,N_5708);
and U5862 (N_5862,N_5793,N_5761);
nand U5863 (N_5863,N_5760,N_5782);
nor U5864 (N_5864,N_5773,N_5712);
or U5865 (N_5865,N_5746,N_5754);
nor U5866 (N_5866,N_5799,N_5772);
and U5867 (N_5867,N_5732,N_5727);
xnor U5868 (N_5868,N_5725,N_5774);
nor U5869 (N_5869,N_5787,N_5728);
and U5870 (N_5870,N_5767,N_5736);
xnor U5871 (N_5871,N_5756,N_5743);
or U5872 (N_5872,N_5748,N_5706);
and U5873 (N_5873,N_5786,N_5700);
or U5874 (N_5874,N_5707,N_5778);
and U5875 (N_5875,N_5719,N_5713);
xnor U5876 (N_5876,N_5748,N_5790);
nor U5877 (N_5877,N_5743,N_5782);
nand U5878 (N_5878,N_5762,N_5734);
xnor U5879 (N_5879,N_5765,N_5780);
nor U5880 (N_5880,N_5739,N_5765);
or U5881 (N_5881,N_5789,N_5723);
nand U5882 (N_5882,N_5754,N_5722);
xnor U5883 (N_5883,N_5700,N_5752);
and U5884 (N_5884,N_5726,N_5761);
nand U5885 (N_5885,N_5777,N_5700);
or U5886 (N_5886,N_5755,N_5758);
xnor U5887 (N_5887,N_5767,N_5749);
and U5888 (N_5888,N_5796,N_5768);
or U5889 (N_5889,N_5791,N_5743);
or U5890 (N_5890,N_5730,N_5799);
or U5891 (N_5891,N_5700,N_5712);
or U5892 (N_5892,N_5705,N_5742);
and U5893 (N_5893,N_5705,N_5708);
nand U5894 (N_5894,N_5777,N_5797);
or U5895 (N_5895,N_5766,N_5732);
xor U5896 (N_5896,N_5734,N_5747);
nor U5897 (N_5897,N_5760,N_5785);
nor U5898 (N_5898,N_5716,N_5709);
xnor U5899 (N_5899,N_5744,N_5759);
or U5900 (N_5900,N_5862,N_5822);
nor U5901 (N_5901,N_5856,N_5877);
nor U5902 (N_5902,N_5832,N_5826);
and U5903 (N_5903,N_5853,N_5897);
nand U5904 (N_5904,N_5879,N_5852);
nor U5905 (N_5905,N_5867,N_5821);
or U5906 (N_5906,N_5813,N_5845);
nor U5907 (N_5907,N_5887,N_5869);
nand U5908 (N_5908,N_5824,N_5870);
nor U5909 (N_5909,N_5895,N_5894);
nor U5910 (N_5910,N_5866,N_5817);
xnor U5911 (N_5911,N_5806,N_5881);
xnor U5912 (N_5912,N_5854,N_5814);
xor U5913 (N_5913,N_5892,N_5863);
nand U5914 (N_5914,N_5888,N_5860);
xor U5915 (N_5915,N_5899,N_5811);
and U5916 (N_5916,N_5830,N_5868);
nand U5917 (N_5917,N_5840,N_5898);
or U5918 (N_5918,N_5818,N_5828);
and U5919 (N_5919,N_5873,N_5855);
and U5920 (N_5920,N_5893,N_5843);
nand U5921 (N_5921,N_5861,N_5802);
xnor U5922 (N_5922,N_5833,N_5882);
nand U5923 (N_5923,N_5835,N_5801);
or U5924 (N_5924,N_5889,N_5857);
and U5925 (N_5925,N_5871,N_5859);
and U5926 (N_5926,N_5875,N_5807);
and U5927 (N_5927,N_5849,N_5876);
or U5928 (N_5928,N_5883,N_5880);
nand U5929 (N_5929,N_5805,N_5841);
or U5930 (N_5930,N_5823,N_5884);
or U5931 (N_5931,N_5831,N_5896);
and U5932 (N_5932,N_5850,N_5839);
or U5933 (N_5933,N_5803,N_5827);
nor U5934 (N_5934,N_5872,N_5836);
or U5935 (N_5935,N_5858,N_5885);
nand U5936 (N_5936,N_5809,N_5838);
or U5937 (N_5937,N_5844,N_5819);
and U5938 (N_5938,N_5851,N_5846);
and U5939 (N_5939,N_5820,N_5878);
xnor U5940 (N_5940,N_5804,N_5829);
nand U5941 (N_5941,N_5816,N_5842);
nand U5942 (N_5942,N_5865,N_5886);
and U5943 (N_5943,N_5890,N_5808);
nand U5944 (N_5944,N_5834,N_5864);
and U5945 (N_5945,N_5812,N_5847);
or U5946 (N_5946,N_5874,N_5891);
nor U5947 (N_5947,N_5837,N_5825);
or U5948 (N_5948,N_5810,N_5800);
and U5949 (N_5949,N_5848,N_5815);
nand U5950 (N_5950,N_5887,N_5832);
and U5951 (N_5951,N_5814,N_5846);
and U5952 (N_5952,N_5863,N_5802);
xnor U5953 (N_5953,N_5859,N_5880);
nand U5954 (N_5954,N_5894,N_5808);
xnor U5955 (N_5955,N_5882,N_5857);
and U5956 (N_5956,N_5849,N_5869);
xor U5957 (N_5957,N_5892,N_5896);
nor U5958 (N_5958,N_5864,N_5800);
and U5959 (N_5959,N_5872,N_5862);
nor U5960 (N_5960,N_5871,N_5886);
or U5961 (N_5961,N_5891,N_5875);
and U5962 (N_5962,N_5888,N_5814);
xnor U5963 (N_5963,N_5844,N_5824);
nand U5964 (N_5964,N_5804,N_5856);
and U5965 (N_5965,N_5894,N_5854);
or U5966 (N_5966,N_5838,N_5821);
or U5967 (N_5967,N_5811,N_5873);
nand U5968 (N_5968,N_5886,N_5838);
or U5969 (N_5969,N_5883,N_5867);
xnor U5970 (N_5970,N_5876,N_5858);
or U5971 (N_5971,N_5869,N_5873);
xor U5972 (N_5972,N_5894,N_5897);
and U5973 (N_5973,N_5811,N_5895);
xor U5974 (N_5974,N_5846,N_5894);
or U5975 (N_5975,N_5865,N_5897);
and U5976 (N_5976,N_5811,N_5844);
nor U5977 (N_5977,N_5825,N_5850);
xor U5978 (N_5978,N_5897,N_5852);
xor U5979 (N_5979,N_5820,N_5893);
nor U5980 (N_5980,N_5852,N_5856);
nor U5981 (N_5981,N_5860,N_5865);
or U5982 (N_5982,N_5801,N_5865);
and U5983 (N_5983,N_5822,N_5845);
nor U5984 (N_5984,N_5801,N_5898);
and U5985 (N_5985,N_5887,N_5856);
xor U5986 (N_5986,N_5861,N_5871);
or U5987 (N_5987,N_5899,N_5879);
or U5988 (N_5988,N_5810,N_5835);
xnor U5989 (N_5989,N_5885,N_5888);
and U5990 (N_5990,N_5828,N_5832);
or U5991 (N_5991,N_5841,N_5851);
and U5992 (N_5992,N_5861,N_5848);
xnor U5993 (N_5993,N_5885,N_5813);
xnor U5994 (N_5994,N_5861,N_5867);
or U5995 (N_5995,N_5803,N_5825);
xor U5996 (N_5996,N_5811,N_5855);
or U5997 (N_5997,N_5803,N_5828);
xor U5998 (N_5998,N_5832,N_5823);
xnor U5999 (N_5999,N_5848,N_5855);
xnor U6000 (N_6000,N_5967,N_5905);
nand U6001 (N_6001,N_5986,N_5900);
xor U6002 (N_6002,N_5930,N_5981);
nand U6003 (N_6003,N_5964,N_5938);
or U6004 (N_6004,N_5979,N_5973);
xor U6005 (N_6005,N_5925,N_5966);
nand U6006 (N_6006,N_5984,N_5923);
nand U6007 (N_6007,N_5965,N_5951);
nor U6008 (N_6008,N_5968,N_5918);
or U6009 (N_6009,N_5928,N_5929);
and U6010 (N_6010,N_5901,N_5940);
or U6011 (N_6011,N_5956,N_5957);
xor U6012 (N_6012,N_5960,N_5955);
nand U6013 (N_6013,N_5907,N_5982);
nor U6014 (N_6014,N_5946,N_5961);
and U6015 (N_6015,N_5948,N_5992);
xnor U6016 (N_6016,N_5989,N_5920);
nand U6017 (N_6017,N_5902,N_5987);
nor U6018 (N_6018,N_5937,N_5936);
and U6019 (N_6019,N_5963,N_5993);
xor U6020 (N_6020,N_5995,N_5911);
or U6021 (N_6021,N_5926,N_5903);
nand U6022 (N_6022,N_5917,N_5978);
nor U6023 (N_6023,N_5962,N_5924);
xor U6024 (N_6024,N_5942,N_5908);
nand U6025 (N_6025,N_5935,N_5972);
and U6026 (N_6026,N_5976,N_5922);
or U6027 (N_6027,N_5934,N_5932);
nand U6028 (N_6028,N_5980,N_5970);
nand U6029 (N_6029,N_5941,N_5953);
xnor U6030 (N_6030,N_5931,N_5959);
nand U6031 (N_6031,N_5983,N_5991);
xnor U6032 (N_6032,N_5969,N_5996);
and U6033 (N_6033,N_5947,N_5921);
and U6034 (N_6034,N_5914,N_5927);
xnor U6035 (N_6035,N_5975,N_5919);
and U6036 (N_6036,N_5943,N_5913);
xor U6037 (N_6037,N_5971,N_5974);
xor U6038 (N_6038,N_5949,N_5988);
or U6039 (N_6039,N_5952,N_5939);
xnor U6040 (N_6040,N_5904,N_5916);
nand U6041 (N_6041,N_5997,N_5915);
or U6042 (N_6042,N_5954,N_5994);
xnor U6043 (N_6043,N_5909,N_5958);
nand U6044 (N_6044,N_5950,N_5944);
nand U6045 (N_6045,N_5945,N_5933);
nor U6046 (N_6046,N_5998,N_5985);
xor U6047 (N_6047,N_5999,N_5977);
nor U6048 (N_6048,N_5912,N_5910);
xor U6049 (N_6049,N_5906,N_5990);
nand U6050 (N_6050,N_5913,N_5980);
nor U6051 (N_6051,N_5903,N_5949);
or U6052 (N_6052,N_5955,N_5931);
nor U6053 (N_6053,N_5938,N_5985);
nor U6054 (N_6054,N_5911,N_5939);
nand U6055 (N_6055,N_5918,N_5946);
nand U6056 (N_6056,N_5920,N_5925);
and U6057 (N_6057,N_5902,N_5984);
and U6058 (N_6058,N_5974,N_5934);
and U6059 (N_6059,N_5990,N_5966);
or U6060 (N_6060,N_5990,N_5911);
or U6061 (N_6061,N_5988,N_5919);
xor U6062 (N_6062,N_5969,N_5979);
or U6063 (N_6063,N_5913,N_5967);
and U6064 (N_6064,N_5938,N_5927);
nand U6065 (N_6065,N_5961,N_5937);
nand U6066 (N_6066,N_5924,N_5997);
nor U6067 (N_6067,N_5933,N_5949);
or U6068 (N_6068,N_5904,N_5942);
xnor U6069 (N_6069,N_5912,N_5988);
nand U6070 (N_6070,N_5922,N_5903);
or U6071 (N_6071,N_5989,N_5906);
or U6072 (N_6072,N_5945,N_5954);
or U6073 (N_6073,N_5937,N_5981);
nor U6074 (N_6074,N_5948,N_5972);
xor U6075 (N_6075,N_5948,N_5919);
nor U6076 (N_6076,N_5999,N_5949);
xor U6077 (N_6077,N_5992,N_5933);
and U6078 (N_6078,N_5964,N_5972);
or U6079 (N_6079,N_5910,N_5939);
xor U6080 (N_6080,N_5909,N_5988);
nand U6081 (N_6081,N_5972,N_5971);
nor U6082 (N_6082,N_5907,N_5912);
nor U6083 (N_6083,N_5946,N_5947);
nand U6084 (N_6084,N_5920,N_5992);
or U6085 (N_6085,N_5935,N_5907);
nor U6086 (N_6086,N_5937,N_5972);
nor U6087 (N_6087,N_5922,N_5951);
nor U6088 (N_6088,N_5957,N_5996);
xor U6089 (N_6089,N_5970,N_5923);
nor U6090 (N_6090,N_5970,N_5917);
nor U6091 (N_6091,N_5918,N_5958);
xor U6092 (N_6092,N_5964,N_5980);
xor U6093 (N_6093,N_5950,N_5931);
nor U6094 (N_6094,N_5995,N_5953);
nand U6095 (N_6095,N_5940,N_5932);
or U6096 (N_6096,N_5955,N_5912);
and U6097 (N_6097,N_5970,N_5992);
nor U6098 (N_6098,N_5914,N_5932);
and U6099 (N_6099,N_5963,N_5942);
xnor U6100 (N_6100,N_6082,N_6004);
nand U6101 (N_6101,N_6075,N_6052);
nor U6102 (N_6102,N_6059,N_6044);
xnor U6103 (N_6103,N_6067,N_6024);
nor U6104 (N_6104,N_6023,N_6021);
and U6105 (N_6105,N_6042,N_6049);
nand U6106 (N_6106,N_6010,N_6097);
or U6107 (N_6107,N_6090,N_6095);
and U6108 (N_6108,N_6048,N_6071);
or U6109 (N_6109,N_6045,N_6093);
nor U6110 (N_6110,N_6047,N_6013);
or U6111 (N_6111,N_6036,N_6041);
nand U6112 (N_6112,N_6068,N_6035);
nand U6113 (N_6113,N_6043,N_6072);
nor U6114 (N_6114,N_6055,N_6098);
xnor U6115 (N_6115,N_6096,N_6064);
nand U6116 (N_6116,N_6066,N_6094);
nor U6117 (N_6117,N_6011,N_6025);
or U6118 (N_6118,N_6062,N_6017);
nand U6119 (N_6119,N_6050,N_6002);
and U6120 (N_6120,N_6091,N_6074);
and U6121 (N_6121,N_6056,N_6081);
xnor U6122 (N_6122,N_6026,N_6019);
xnor U6123 (N_6123,N_6018,N_6046);
nand U6124 (N_6124,N_6084,N_6009);
nor U6125 (N_6125,N_6032,N_6063);
nand U6126 (N_6126,N_6078,N_6007);
nand U6127 (N_6127,N_6080,N_6073);
or U6128 (N_6128,N_6092,N_6015);
and U6129 (N_6129,N_6037,N_6088);
nand U6130 (N_6130,N_6087,N_6057);
and U6131 (N_6131,N_6076,N_6030);
xor U6132 (N_6132,N_6038,N_6006);
nand U6133 (N_6133,N_6085,N_6039);
xor U6134 (N_6134,N_6089,N_6000);
xor U6135 (N_6135,N_6028,N_6001);
and U6136 (N_6136,N_6054,N_6060);
and U6137 (N_6137,N_6053,N_6070);
and U6138 (N_6138,N_6083,N_6022);
nor U6139 (N_6139,N_6029,N_6061);
nor U6140 (N_6140,N_6034,N_6027);
nand U6141 (N_6141,N_6040,N_6099);
xnor U6142 (N_6142,N_6086,N_6031);
nand U6143 (N_6143,N_6077,N_6003);
and U6144 (N_6144,N_6020,N_6079);
nor U6145 (N_6145,N_6065,N_6005);
or U6146 (N_6146,N_6058,N_6014);
nor U6147 (N_6147,N_6008,N_6016);
or U6148 (N_6148,N_6069,N_6033);
nand U6149 (N_6149,N_6051,N_6012);
xor U6150 (N_6150,N_6090,N_6061);
or U6151 (N_6151,N_6025,N_6032);
nor U6152 (N_6152,N_6049,N_6014);
and U6153 (N_6153,N_6070,N_6085);
xnor U6154 (N_6154,N_6017,N_6036);
and U6155 (N_6155,N_6033,N_6053);
and U6156 (N_6156,N_6043,N_6024);
or U6157 (N_6157,N_6091,N_6084);
nand U6158 (N_6158,N_6087,N_6072);
or U6159 (N_6159,N_6039,N_6054);
and U6160 (N_6160,N_6050,N_6018);
nor U6161 (N_6161,N_6066,N_6077);
nor U6162 (N_6162,N_6060,N_6069);
nor U6163 (N_6163,N_6078,N_6004);
nand U6164 (N_6164,N_6031,N_6033);
xor U6165 (N_6165,N_6058,N_6056);
xor U6166 (N_6166,N_6090,N_6060);
or U6167 (N_6167,N_6097,N_6005);
and U6168 (N_6168,N_6072,N_6076);
nand U6169 (N_6169,N_6035,N_6017);
and U6170 (N_6170,N_6013,N_6056);
nand U6171 (N_6171,N_6001,N_6088);
or U6172 (N_6172,N_6016,N_6094);
nand U6173 (N_6173,N_6085,N_6046);
xnor U6174 (N_6174,N_6088,N_6044);
or U6175 (N_6175,N_6033,N_6088);
nand U6176 (N_6176,N_6051,N_6070);
nor U6177 (N_6177,N_6074,N_6087);
nor U6178 (N_6178,N_6084,N_6008);
nand U6179 (N_6179,N_6025,N_6063);
and U6180 (N_6180,N_6083,N_6063);
or U6181 (N_6181,N_6059,N_6016);
or U6182 (N_6182,N_6014,N_6069);
nand U6183 (N_6183,N_6063,N_6034);
and U6184 (N_6184,N_6097,N_6080);
or U6185 (N_6185,N_6057,N_6036);
nand U6186 (N_6186,N_6039,N_6050);
and U6187 (N_6187,N_6035,N_6073);
and U6188 (N_6188,N_6042,N_6037);
or U6189 (N_6189,N_6025,N_6061);
or U6190 (N_6190,N_6027,N_6010);
nand U6191 (N_6191,N_6079,N_6076);
and U6192 (N_6192,N_6070,N_6017);
nand U6193 (N_6193,N_6097,N_6002);
or U6194 (N_6194,N_6072,N_6091);
or U6195 (N_6195,N_6090,N_6039);
nand U6196 (N_6196,N_6097,N_6066);
and U6197 (N_6197,N_6093,N_6000);
nand U6198 (N_6198,N_6075,N_6079);
xor U6199 (N_6199,N_6057,N_6076);
and U6200 (N_6200,N_6166,N_6194);
nor U6201 (N_6201,N_6107,N_6106);
nor U6202 (N_6202,N_6184,N_6191);
xnor U6203 (N_6203,N_6192,N_6160);
nor U6204 (N_6204,N_6111,N_6198);
nand U6205 (N_6205,N_6159,N_6153);
and U6206 (N_6206,N_6151,N_6158);
and U6207 (N_6207,N_6183,N_6149);
and U6208 (N_6208,N_6117,N_6131);
nand U6209 (N_6209,N_6142,N_6120);
nand U6210 (N_6210,N_6125,N_6197);
nand U6211 (N_6211,N_6177,N_6167);
or U6212 (N_6212,N_6190,N_6127);
xor U6213 (N_6213,N_6102,N_6123);
nor U6214 (N_6214,N_6163,N_6143);
and U6215 (N_6215,N_6148,N_6108);
nand U6216 (N_6216,N_6115,N_6196);
or U6217 (N_6217,N_6112,N_6155);
nor U6218 (N_6218,N_6134,N_6100);
or U6219 (N_6219,N_6119,N_6193);
or U6220 (N_6220,N_6162,N_6116);
and U6221 (N_6221,N_6145,N_6103);
and U6222 (N_6222,N_6129,N_6122);
and U6223 (N_6223,N_6124,N_6121);
xnor U6224 (N_6224,N_6136,N_6140);
xnor U6225 (N_6225,N_6173,N_6157);
or U6226 (N_6226,N_6175,N_6152);
nor U6227 (N_6227,N_6195,N_6133);
xnor U6228 (N_6228,N_6179,N_6135);
and U6229 (N_6229,N_6137,N_6174);
nor U6230 (N_6230,N_6154,N_6178);
xor U6231 (N_6231,N_6156,N_6130);
and U6232 (N_6232,N_6141,N_6199);
nand U6233 (N_6233,N_6144,N_6168);
nor U6234 (N_6234,N_6185,N_6109);
or U6235 (N_6235,N_6182,N_6176);
nand U6236 (N_6236,N_6164,N_6126);
and U6237 (N_6237,N_6114,N_6181);
or U6238 (N_6238,N_6161,N_6150);
nand U6239 (N_6239,N_6180,N_6147);
nand U6240 (N_6240,N_6132,N_6172);
nand U6241 (N_6241,N_6169,N_6104);
xor U6242 (N_6242,N_6101,N_6110);
and U6243 (N_6243,N_6128,N_6118);
or U6244 (N_6244,N_6113,N_6189);
xor U6245 (N_6245,N_6138,N_6105);
nor U6246 (N_6246,N_6139,N_6170);
xor U6247 (N_6247,N_6171,N_6187);
nor U6248 (N_6248,N_6146,N_6165);
nand U6249 (N_6249,N_6188,N_6186);
nand U6250 (N_6250,N_6121,N_6153);
and U6251 (N_6251,N_6178,N_6199);
nor U6252 (N_6252,N_6143,N_6149);
nand U6253 (N_6253,N_6199,N_6169);
or U6254 (N_6254,N_6116,N_6130);
xnor U6255 (N_6255,N_6130,N_6170);
or U6256 (N_6256,N_6187,N_6174);
and U6257 (N_6257,N_6102,N_6191);
nand U6258 (N_6258,N_6188,N_6129);
nor U6259 (N_6259,N_6159,N_6143);
xor U6260 (N_6260,N_6127,N_6186);
or U6261 (N_6261,N_6137,N_6136);
or U6262 (N_6262,N_6199,N_6174);
nand U6263 (N_6263,N_6191,N_6113);
nand U6264 (N_6264,N_6171,N_6190);
or U6265 (N_6265,N_6109,N_6144);
and U6266 (N_6266,N_6182,N_6165);
and U6267 (N_6267,N_6145,N_6189);
xnor U6268 (N_6268,N_6192,N_6190);
xor U6269 (N_6269,N_6137,N_6111);
xnor U6270 (N_6270,N_6109,N_6111);
nor U6271 (N_6271,N_6137,N_6187);
nand U6272 (N_6272,N_6166,N_6141);
or U6273 (N_6273,N_6166,N_6100);
or U6274 (N_6274,N_6142,N_6176);
nor U6275 (N_6275,N_6177,N_6117);
xor U6276 (N_6276,N_6185,N_6174);
nor U6277 (N_6277,N_6125,N_6123);
or U6278 (N_6278,N_6189,N_6183);
xor U6279 (N_6279,N_6178,N_6141);
and U6280 (N_6280,N_6134,N_6188);
nor U6281 (N_6281,N_6160,N_6115);
xnor U6282 (N_6282,N_6113,N_6115);
nor U6283 (N_6283,N_6153,N_6170);
or U6284 (N_6284,N_6142,N_6125);
nand U6285 (N_6285,N_6170,N_6109);
nor U6286 (N_6286,N_6117,N_6186);
or U6287 (N_6287,N_6123,N_6179);
or U6288 (N_6288,N_6135,N_6149);
nor U6289 (N_6289,N_6145,N_6181);
xor U6290 (N_6290,N_6160,N_6131);
and U6291 (N_6291,N_6198,N_6112);
xor U6292 (N_6292,N_6164,N_6109);
nor U6293 (N_6293,N_6127,N_6111);
and U6294 (N_6294,N_6182,N_6102);
xnor U6295 (N_6295,N_6187,N_6168);
xor U6296 (N_6296,N_6170,N_6103);
xnor U6297 (N_6297,N_6115,N_6154);
and U6298 (N_6298,N_6155,N_6116);
and U6299 (N_6299,N_6164,N_6151);
xnor U6300 (N_6300,N_6244,N_6250);
nor U6301 (N_6301,N_6226,N_6296);
or U6302 (N_6302,N_6234,N_6202);
or U6303 (N_6303,N_6222,N_6221);
nand U6304 (N_6304,N_6239,N_6203);
xnor U6305 (N_6305,N_6282,N_6256);
nor U6306 (N_6306,N_6268,N_6267);
nor U6307 (N_6307,N_6270,N_6261);
xor U6308 (N_6308,N_6232,N_6272);
nand U6309 (N_6309,N_6266,N_6257);
or U6310 (N_6310,N_6269,N_6292);
and U6311 (N_6311,N_6290,N_6213);
and U6312 (N_6312,N_6207,N_6249);
or U6313 (N_6313,N_6260,N_6209);
and U6314 (N_6314,N_6230,N_6218);
nand U6315 (N_6315,N_6289,N_6200);
nor U6316 (N_6316,N_6219,N_6220);
nor U6317 (N_6317,N_6287,N_6225);
nor U6318 (N_6318,N_6262,N_6237);
nand U6319 (N_6319,N_6280,N_6201);
xor U6320 (N_6320,N_6279,N_6274);
nand U6321 (N_6321,N_6214,N_6295);
nor U6322 (N_6322,N_6228,N_6286);
xor U6323 (N_6323,N_6277,N_6271);
xor U6324 (N_6324,N_6251,N_6255);
nand U6325 (N_6325,N_6281,N_6208);
or U6326 (N_6326,N_6224,N_6233);
nand U6327 (N_6327,N_6241,N_6273);
or U6328 (N_6328,N_6247,N_6297);
nor U6329 (N_6329,N_6253,N_6211);
nor U6330 (N_6330,N_6283,N_6293);
nor U6331 (N_6331,N_6254,N_6288);
and U6332 (N_6332,N_6284,N_6265);
or U6333 (N_6333,N_6276,N_6258);
or U6334 (N_6334,N_6291,N_6259);
xor U6335 (N_6335,N_6263,N_6227);
xnor U6336 (N_6336,N_6236,N_6246);
nand U6337 (N_6337,N_6240,N_6204);
and U6338 (N_6338,N_6205,N_6217);
xnor U6339 (N_6339,N_6248,N_6206);
and U6340 (N_6340,N_6285,N_6229);
nand U6341 (N_6341,N_6243,N_6216);
or U6342 (N_6342,N_6215,N_6235);
nand U6343 (N_6343,N_6210,N_6264);
nand U6344 (N_6344,N_6231,N_6245);
nand U6345 (N_6345,N_6212,N_6238);
nand U6346 (N_6346,N_6275,N_6223);
xor U6347 (N_6347,N_6278,N_6252);
xnor U6348 (N_6348,N_6294,N_6298);
xor U6349 (N_6349,N_6242,N_6299);
nor U6350 (N_6350,N_6229,N_6208);
or U6351 (N_6351,N_6224,N_6229);
nor U6352 (N_6352,N_6289,N_6245);
nand U6353 (N_6353,N_6207,N_6224);
or U6354 (N_6354,N_6248,N_6254);
nand U6355 (N_6355,N_6267,N_6218);
nand U6356 (N_6356,N_6226,N_6252);
nand U6357 (N_6357,N_6231,N_6235);
nor U6358 (N_6358,N_6207,N_6213);
or U6359 (N_6359,N_6211,N_6254);
and U6360 (N_6360,N_6297,N_6287);
xnor U6361 (N_6361,N_6287,N_6234);
xnor U6362 (N_6362,N_6255,N_6202);
or U6363 (N_6363,N_6242,N_6244);
or U6364 (N_6364,N_6233,N_6228);
nor U6365 (N_6365,N_6244,N_6218);
or U6366 (N_6366,N_6283,N_6233);
or U6367 (N_6367,N_6211,N_6281);
nand U6368 (N_6368,N_6247,N_6281);
nand U6369 (N_6369,N_6231,N_6256);
nand U6370 (N_6370,N_6205,N_6237);
and U6371 (N_6371,N_6206,N_6226);
nor U6372 (N_6372,N_6216,N_6286);
xor U6373 (N_6373,N_6245,N_6203);
xnor U6374 (N_6374,N_6297,N_6214);
and U6375 (N_6375,N_6259,N_6223);
or U6376 (N_6376,N_6287,N_6289);
or U6377 (N_6377,N_6216,N_6263);
xor U6378 (N_6378,N_6271,N_6293);
and U6379 (N_6379,N_6268,N_6273);
and U6380 (N_6380,N_6288,N_6207);
or U6381 (N_6381,N_6202,N_6262);
xnor U6382 (N_6382,N_6256,N_6273);
xnor U6383 (N_6383,N_6293,N_6230);
xor U6384 (N_6384,N_6237,N_6271);
or U6385 (N_6385,N_6203,N_6288);
nor U6386 (N_6386,N_6297,N_6299);
xor U6387 (N_6387,N_6261,N_6236);
and U6388 (N_6388,N_6277,N_6285);
nand U6389 (N_6389,N_6246,N_6255);
nand U6390 (N_6390,N_6227,N_6232);
nor U6391 (N_6391,N_6299,N_6255);
or U6392 (N_6392,N_6233,N_6270);
nand U6393 (N_6393,N_6297,N_6245);
nand U6394 (N_6394,N_6209,N_6221);
or U6395 (N_6395,N_6279,N_6241);
nor U6396 (N_6396,N_6214,N_6232);
nor U6397 (N_6397,N_6278,N_6266);
or U6398 (N_6398,N_6272,N_6299);
and U6399 (N_6399,N_6223,N_6217);
nand U6400 (N_6400,N_6361,N_6306);
and U6401 (N_6401,N_6367,N_6326);
or U6402 (N_6402,N_6382,N_6358);
nand U6403 (N_6403,N_6374,N_6381);
nor U6404 (N_6404,N_6320,N_6334);
xor U6405 (N_6405,N_6378,N_6304);
and U6406 (N_6406,N_6388,N_6341);
xor U6407 (N_6407,N_6318,N_6302);
xnor U6408 (N_6408,N_6389,N_6323);
or U6409 (N_6409,N_6317,N_6357);
or U6410 (N_6410,N_6309,N_6359);
nor U6411 (N_6411,N_6360,N_6344);
or U6412 (N_6412,N_6371,N_6363);
and U6413 (N_6413,N_6351,N_6368);
and U6414 (N_6414,N_6312,N_6394);
and U6415 (N_6415,N_6379,N_6325);
nor U6416 (N_6416,N_6376,N_6375);
nand U6417 (N_6417,N_6397,N_6337);
nand U6418 (N_6418,N_6340,N_6315);
nor U6419 (N_6419,N_6398,N_6321);
or U6420 (N_6420,N_6353,N_6333);
xnor U6421 (N_6421,N_6310,N_6342);
and U6422 (N_6422,N_6339,N_6327);
or U6423 (N_6423,N_6355,N_6332);
or U6424 (N_6424,N_6328,N_6364);
or U6425 (N_6425,N_6380,N_6301);
and U6426 (N_6426,N_6319,N_6343);
and U6427 (N_6427,N_6350,N_6347);
xor U6428 (N_6428,N_6393,N_6322);
nor U6429 (N_6429,N_6356,N_6392);
and U6430 (N_6430,N_6324,N_6335);
and U6431 (N_6431,N_6399,N_6354);
and U6432 (N_6432,N_6345,N_6372);
or U6433 (N_6433,N_6305,N_6331);
xnor U6434 (N_6434,N_6300,N_6395);
nand U6435 (N_6435,N_6330,N_6391);
nand U6436 (N_6436,N_6313,N_6370);
and U6437 (N_6437,N_6303,N_6385);
and U6438 (N_6438,N_6386,N_6308);
nand U6439 (N_6439,N_6366,N_6349);
or U6440 (N_6440,N_6346,N_6311);
nor U6441 (N_6441,N_6314,N_6338);
nand U6442 (N_6442,N_6390,N_6336);
nor U6443 (N_6443,N_6383,N_6348);
xor U6444 (N_6444,N_6377,N_6384);
or U6445 (N_6445,N_6352,N_6387);
xnor U6446 (N_6446,N_6316,N_6365);
nor U6447 (N_6447,N_6369,N_6373);
or U6448 (N_6448,N_6307,N_6396);
nor U6449 (N_6449,N_6329,N_6362);
nor U6450 (N_6450,N_6338,N_6343);
nor U6451 (N_6451,N_6355,N_6365);
or U6452 (N_6452,N_6355,N_6379);
xnor U6453 (N_6453,N_6378,N_6356);
nand U6454 (N_6454,N_6303,N_6333);
or U6455 (N_6455,N_6366,N_6308);
nor U6456 (N_6456,N_6340,N_6338);
nand U6457 (N_6457,N_6375,N_6304);
or U6458 (N_6458,N_6359,N_6361);
nand U6459 (N_6459,N_6302,N_6390);
nor U6460 (N_6460,N_6372,N_6366);
and U6461 (N_6461,N_6398,N_6389);
or U6462 (N_6462,N_6363,N_6349);
and U6463 (N_6463,N_6363,N_6396);
nand U6464 (N_6464,N_6320,N_6301);
and U6465 (N_6465,N_6336,N_6327);
or U6466 (N_6466,N_6347,N_6310);
or U6467 (N_6467,N_6358,N_6370);
xor U6468 (N_6468,N_6308,N_6348);
and U6469 (N_6469,N_6376,N_6379);
or U6470 (N_6470,N_6318,N_6352);
xnor U6471 (N_6471,N_6312,N_6326);
nor U6472 (N_6472,N_6317,N_6362);
xnor U6473 (N_6473,N_6329,N_6348);
or U6474 (N_6474,N_6351,N_6347);
nor U6475 (N_6475,N_6366,N_6376);
or U6476 (N_6476,N_6399,N_6306);
xor U6477 (N_6477,N_6365,N_6374);
nand U6478 (N_6478,N_6316,N_6303);
xnor U6479 (N_6479,N_6309,N_6352);
xnor U6480 (N_6480,N_6318,N_6322);
and U6481 (N_6481,N_6374,N_6303);
nor U6482 (N_6482,N_6363,N_6348);
nor U6483 (N_6483,N_6315,N_6349);
or U6484 (N_6484,N_6334,N_6328);
xnor U6485 (N_6485,N_6360,N_6395);
or U6486 (N_6486,N_6375,N_6380);
nand U6487 (N_6487,N_6393,N_6380);
or U6488 (N_6488,N_6335,N_6380);
and U6489 (N_6489,N_6398,N_6349);
nand U6490 (N_6490,N_6319,N_6346);
xor U6491 (N_6491,N_6399,N_6352);
and U6492 (N_6492,N_6330,N_6323);
and U6493 (N_6493,N_6360,N_6333);
nand U6494 (N_6494,N_6375,N_6361);
nor U6495 (N_6495,N_6308,N_6350);
and U6496 (N_6496,N_6362,N_6315);
xnor U6497 (N_6497,N_6315,N_6319);
nand U6498 (N_6498,N_6348,N_6307);
nor U6499 (N_6499,N_6365,N_6363);
nand U6500 (N_6500,N_6444,N_6400);
or U6501 (N_6501,N_6467,N_6484);
nor U6502 (N_6502,N_6402,N_6499);
xor U6503 (N_6503,N_6434,N_6431);
and U6504 (N_6504,N_6414,N_6410);
and U6505 (N_6505,N_6416,N_6439);
nand U6506 (N_6506,N_6405,N_6436);
and U6507 (N_6507,N_6475,N_6492);
or U6508 (N_6508,N_6403,N_6426);
nor U6509 (N_6509,N_6415,N_6401);
and U6510 (N_6510,N_6461,N_6470);
nor U6511 (N_6511,N_6407,N_6428);
or U6512 (N_6512,N_6411,N_6447);
and U6513 (N_6513,N_6430,N_6455);
nor U6514 (N_6514,N_6423,N_6483);
xor U6515 (N_6515,N_6429,N_6469);
xnor U6516 (N_6516,N_6438,N_6462);
xor U6517 (N_6517,N_6420,N_6445);
nand U6518 (N_6518,N_6456,N_6487);
xnor U6519 (N_6519,N_6422,N_6424);
nor U6520 (N_6520,N_6408,N_6457);
and U6521 (N_6521,N_6441,N_6409);
and U6522 (N_6522,N_6448,N_6480);
or U6523 (N_6523,N_6450,N_6471);
nand U6524 (N_6524,N_6419,N_6442);
nor U6525 (N_6525,N_6498,N_6493);
and U6526 (N_6526,N_6474,N_6421);
nand U6527 (N_6527,N_6459,N_6496);
or U6528 (N_6528,N_6473,N_6440);
nand U6529 (N_6529,N_6481,N_6465);
nor U6530 (N_6530,N_6449,N_6463);
xor U6531 (N_6531,N_6482,N_6466);
nor U6532 (N_6532,N_6472,N_6451);
xor U6533 (N_6533,N_6413,N_6406);
nor U6534 (N_6534,N_6418,N_6490);
nand U6535 (N_6535,N_6489,N_6458);
or U6536 (N_6536,N_6468,N_6477);
nand U6537 (N_6537,N_6497,N_6460);
or U6538 (N_6538,N_6404,N_6488);
and U6539 (N_6539,N_6412,N_6478);
nand U6540 (N_6540,N_6464,N_6425);
nand U6541 (N_6541,N_6433,N_6479);
or U6542 (N_6542,N_6446,N_6437);
or U6543 (N_6543,N_6452,N_6432);
nor U6544 (N_6544,N_6491,N_6417);
xnor U6545 (N_6545,N_6443,N_6495);
nor U6546 (N_6546,N_6476,N_6454);
nor U6547 (N_6547,N_6485,N_6427);
or U6548 (N_6548,N_6435,N_6453);
and U6549 (N_6549,N_6494,N_6486);
nor U6550 (N_6550,N_6472,N_6476);
nor U6551 (N_6551,N_6473,N_6454);
xnor U6552 (N_6552,N_6448,N_6409);
and U6553 (N_6553,N_6431,N_6495);
xor U6554 (N_6554,N_6462,N_6422);
and U6555 (N_6555,N_6484,N_6473);
xnor U6556 (N_6556,N_6497,N_6462);
xor U6557 (N_6557,N_6463,N_6405);
nor U6558 (N_6558,N_6420,N_6455);
and U6559 (N_6559,N_6429,N_6440);
and U6560 (N_6560,N_6496,N_6482);
nor U6561 (N_6561,N_6481,N_6428);
and U6562 (N_6562,N_6424,N_6406);
nand U6563 (N_6563,N_6443,N_6409);
xnor U6564 (N_6564,N_6472,N_6470);
nor U6565 (N_6565,N_6494,N_6460);
or U6566 (N_6566,N_6499,N_6488);
and U6567 (N_6567,N_6496,N_6450);
nand U6568 (N_6568,N_6449,N_6418);
nor U6569 (N_6569,N_6403,N_6479);
xnor U6570 (N_6570,N_6432,N_6415);
xnor U6571 (N_6571,N_6464,N_6438);
nand U6572 (N_6572,N_6476,N_6409);
and U6573 (N_6573,N_6495,N_6453);
nor U6574 (N_6574,N_6401,N_6409);
and U6575 (N_6575,N_6477,N_6420);
and U6576 (N_6576,N_6470,N_6440);
nand U6577 (N_6577,N_6464,N_6441);
xnor U6578 (N_6578,N_6476,N_6482);
and U6579 (N_6579,N_6456,N_6449);
nand U6580 (N_6580,N_6429,N_6459);
xnor U6581 (N_6581,N_6415,N_6408);
or U6582 (N_6582,N_6414,N_6490);
or U6583 (N_6583,N_6498,N_6419);
or U6584 (N_6584,N_6489,N_6465);
xor U6585 (N_6585,N_6469,N_6427);
nor U6586 (N_6586,N_6479,N_6494);
xor U6587 (N_6587,N_6441,N_6472);
or U6588 (N_6588,N_6466,N_6456);
or U6589 (N_6589,N_6402,N_6439);
or U6590 (N_6590,N_6465,N_6412);
nor U6591 (N_6591,N_6404,N_6412);
or U6592 (N_6592,N_6443,N_6469);
or U6593 (N_6593,N_6461,N_6400);
xnor U6594 (N_6594,N_6492,N_6482);
or U6595 (N_6595,N_6434,N_6455);
xnor U6596 (N_6596,N_6418,N_6436);
or U6597 (N_6597,N_6474,N_6457);
xor U6598 (N_6598,N_6473,N_6478);
nor U6599 (N_6599,N_6481,N_6403);
xor U6600 (N_6600,N_6566,N_6533);
or U6601 (N_6601,N_6589,N_6541);
and U6602 (N_6602,N_6515,N_6588);
and U6603 (N_6603,N_6507,N_6580);
nor U6604 (N_6604,N_6511,N_6538);
and U6605 (N_6605,N_6597,N_6586);
nor U6606 (N_6606,N_6524,N_6577);
and U6607 (N_6607,N_6548,N_6528);
xnor U6608 (N_6608,N_6519,N_6549);
xor U6609 (N_6609,N_6501,N_6517);
nor U6610 (N_6610,N_6504,N_6520);
or U6611 (N_6611,N_6530,N_6522);
nor U6612 (N_6612,N_6521,N_6572);
nor U6613 (N_6613,N_6540,N_6553);
or U6614 (N_6614,N_6557,N_6559);
xor U6615 (N_6615,N_6596,N_6569);
and U6616 (N_6616,N_6510,N_6527);
xnor U6617 (N_6617,N_6568,N_6509);
nor U6618 (N_6618,N_6532,N_6582);
nor U6619 (N_6619,N_6581,N_6594);
xnor U6620 (N_6620,N_6561,N_6575);
xnor U6621 (N_6621,N_6556,N_6560);
and U6622 (N_6622,N_6535,N_6514);
and U6623 (N_6623,N_6508,N_6570);
and U6624 (N_6624,N_6547,N_6593);
nor U6625 (N_6625,N_6573,N_6564);
nand U6626 (N_6626,N_6546,N_6591);
or U6627 (N_6627,N_6526,N_6552);
or U6628 (N_6628,N_6525,N_6562);
nand U6629 (N_6629,N_6579,N_6523);
or U6630 (N_6630,N_6583,N_6574);
nor U6631 (N_6631,N_6536,N_6554);
nand U6632 (N_6632,N_6503,N_6543);
or U6633 (N_6633,N_6513,N_6584);
nor U6634 (N_6634,N_6500,N_6578);
nor U6635 (N_6635,N_6565,N_6590);
or U6636 (N_6636,N_6537,N_6576);
nand U6637 (N_6637,N_6558,N_6516);
nand U6638 (N_6638,N_6505,N_6567);
nand U6639 (N_6639,N_6544,N_6502);
xor U6640 (N_6640,N_6595,N_6539);
xnor U6641 (N_6641,N_6563,N_6518);
or U6642 (N_6642,N_6599,N_6571);
or U6643 (N_6643,N_6587,N_6592);
nor U6644 (N_6644,N_6529,N_6534);
or U6645 (N_6645,N_6555,N_6542);
and U6646 (N_6646,N_6551,N_6585);
xor U6647 (N_6647,N_6598,N_6531);
or U6648 (N_6648,N_6545,N_6512);
or U6649 (N_6649,N_6550,N_6506);
xor U6650 (N_6650,N_6520,N_6547);
nand U6651 (N_6651,N_6556,N_6512);
or U6652 (N_6652,N_6567,N_6516);
or U6653 (N_6653,N_6549,N_6556);
nand U6654 (N_6654,N_6535,N_6576);
xor U6655 (N_6655,N_6583,N_6564);
or U6656 (N_6656,N_6599,N_6590);
nand U6657 (N_6657,N_6554,N_6516);
nand U6658 (N_6658,N_6530,N_6575);
nor U6659 (N_6659,N_6526,N_6591);
or U6660 (N_6660,N_6526,N_6522);
and U6661 (N_6661,N_6585,N_6552);
and U6662 (N_6662,N_6557,N_6522);
xnor U6663 (N_6663,N_6521,N_6591);
xor U6664 (N_6664,N_6582,N_6508);
or U6665 (N_6665,N_6560,N_6585);
nor U6666 (N_6666,N_6563,N_6545);
and U6667 (N_6667,N_6516,N_6528);
nor U6668 (N_6668,N_6536,N_6568);
and U6669 (N_6669,N_6587,N_6509);
xor U6670 (N_6670,N_6523,N_6515);
xor U6671 (N_6671,N_6592,N_6510);
and U6672 (N_6672,N_6519,N_6567);
or U6673 (N_6673,N_6510,N_6562);
xor U6674 (N_6674,N_6526,N_6530);
and U6675 (N_6675,N_6509,N_6577);
or U6676 (N_6676,N_6526,N_6534);
or U6677 (N_6677,N_6509,N_6542);
nand U6678 (N_6678,N_6556,N_6528);
xor U6679 (N_6679,N_6555,N_6526);
or U6680 (N_6680,N_6572,N_6541);
nor U6681 (N_6681,N_6571,N_6583);
and U6682 (N_6682,N_6593,N_6595);
nand U6683 (N_6683,N_6587,N_6521);
nand U6684 (N_6684,N_6537,N_6512);
nand U6685 (N_6685,N_6531,N_6539);
xnor U6686 (N_6686,N_6529,N_6506);
xnor U6687 (N_6687,N_6501,N_6561);
nor U6688 (N_6688,N_6591,N_6547);
nor U6689 (N_6689,N_6560,N_6525);
nor U6690 (N_6690,N_6511,N_6541);
xor U6691 (N_6691,N_6526,N_6543);
or U6692 (N_6692,N_6577,N_6523);
or U6693 (N_6693,N_6563,N_6503);
nand U6694 (N_6694,N_6536,N_6544);
or U6695 (N_6695,N_6522,N_6561);
and U6696 (N_6696,N_6535,N_6555);
xor U6697 (N_6697,N_6598,N_6543);
or U6698 (N_6698,N_6595,N_6587);
nor U6699 (N_6699,N_6541,N_6530);
xor U6700 (N_6700,N_6670,N_6682);
and U6701 (N_6701,N_6684,N_6605);
xnor U6702 (N_6702,N_6678,N_6661);
xor U6703 (N_6703,N_6602,N_6627);
nand U6704 (N_6704,N_6623,N_6610);
xnor U6705 (N_6705,N_6679,N_6674);
xor U6706 (N_6706,N_6696,N_6657);
nor U6707 (N_6707,N_6638,N_6631);
nand U6708 (N_6708,N_6690,N_6676);
nand U6709 (N_6709,N_6667,N_6653);
nor U6710 (N_6710,N_6629,N_6683);
nand U6711 (N_6711,N_6611,N_6642);
xnor U6712 (N_6712,N_6680,N_6644);
nand U6713 (N_6713,N_6665,N_6616);
or U6714 (N_6714,N_6688,N_6632);
and U6715 (N_6715,N_6660,N_6613);
nor U6716 (N_6716,N_6615,N_6621);
and U6717 (N_6717,N_6601,N_6675);
nand U6718 (N_6718,N_6636,N_6640);
nor U6719 (N_6719,N_6687,N_6612);
xnor U6720 (N_6720,N_6689,N_6607);
nor U6721 (N_6721,N_6697,N_6659);
nor U6722 (N_6722,N_6645,N_6622);
nand U6723 (N_6723,N_6698,N_6648);
nand U6724 (N_6724,N_6641,N_6604);
nor U6725 (N_6725,N_6647,N_6656);
nand U6726 (N_6726,N_6658,N_6649);
nor U6727 (N_6727,N_6633,N_6608);
and U6728 (N_6728,N_6692,N_6695);
or U6729 (N_6729,N_6668,N_6618);
xnor U6730 (N_6730,N_6691,N_6639);
nand U6731 (N_6731,N_6663,N_6606);
nor U6732 (N_6732,N_6625,N_6630);
or U6733 (N_6733,N_6664,N_6651);
or U6734 (N_6734,N_6617,N_6672);
and U6735 (N_6735,N_6673,N_6634);
nand U6736 (N_6736,N_6646,N_6609);
xor U6737 (N_6737,N_6677,N_6603);
and U6738 (N_6738,N_6614,N_6619);
nor U6739 (N_6739,N_6662,N_6624);
xor U6740 (N_6740,N_6600,N_6693);
nand U6741 (N_6741,N_6643,N_6635);
nor U6742 (N_6742,N_6654,N_6620);
nand U6743 (N_6743,N_6669,N_6655);
nand U6744 (N_6744,N_6681,N_6699);
and U6745 (N_6745,N_6628,N_6685);
and U6746 (N_6746,N_6626,N_6650);
or U6747 (N_6747,N_6637,N_6694);
nand U6748 (N_6748,N_6671,N_6652);
or U6749 (N_6749,N_6666,N_6686);
nor U6750 (N_6750,N_6655,N_6647);
or U6751 (N_6751,N_6658,N_6690);
or U6752 (N_6752,N_6622,N_6665);
nand U6753 (N_6753,N_6636,N_6643);
xnor U6754 (N_6754,N_6634,N_6647);
and U6755 (N_6755,N_6658,N_6622);
xor U6756 (N_6756,N_6691,N_6622);
xnor U6757 (N_6757,N_6619,N_6632);
nor U6758 (N_6758,N_6650,N_6632);
and U6759 (N_6759,N_6659,N_6687);
nor U6760 (N_6760,N_6691,N_6609);
xor U6761 (N_6761,N_6651,N_6615);
nor U6762 (N_6762,N_6628,N_6657);
nand U6763 (N_6763,N_6641,N_6670);
xnor U6764 (N_6764,N_6658,N_6667);
and U6765 (N_6765,N_6648,N_6642);
xor U6766 (N_6766,N_6655,N_6608);
or U6767 (N_6767,N_6654,N_6657);
nand U6768 (N_6768,N_6613,N_6669);
xor U6769 (N_6769,N_6651,N_6635);
and U6770 (N_6770,N_6627,N_6682);
nor U6771 (N_6771,N_6603,N_6665);
nor U6772 (N_6772,N_6648,N_6604);
nand U6773 (N_6773,N_6600,N_6624);
xnor U6774 (N_6774,N_6697,N_6653);
nor U6775 (N_6775,N_6638,N_6673);
and U6776 (N_6776,N_6626,N_6682);
and U6777 (N_6777,N_6606,N_6647);
or U6778 (N_6778,N_6661,N_6675);
and U6779 (N_6779,N_6682,N_6631);
xor U6780 (N_6780,N_6628,N_6647);
or U6781 (N_6781,N_6690,N_6611);
nand U6782 (N_6782,N_6635,N_6628);
xnor U6783 (N_6783,N_6652,N_6615);
xnor U6784 (N_6784,N_6659,N_6635);
or U6785 (N_6785,N_6614,N_6629);
nand U6786 (N_6786,N_6680,N_6630);
nor U6787 (N_6787,N_6617,N_6690);
nor U6788 (N_6788,N_6602,N_6616);
and U6789 (N_6789,N_6644,N_6635);
nor U6790 (N_6790,N_6610,N_6680);
or U6791 (N_6791,N_6658,N_6665);
or U6792 (N_6792,N_6672,N_6656);
nor U6793 (N_6793,N_6623,N_6605);
xnor U6794 (N_6794,N_6648,N_6635);
nor U6795 (N_6795,N_6616,N_6624);
nand U6796 (N_6796,N_6672,N_6601);
nand U6797 (N_6797,N_6640,N_6693);
nand U6798 (N_6798,N_6674,N_6664);
nor U6799 (N_6799,N_6605,N_6662);
xor U6800 (N_6800,N_6752,N_6702);
nand U6801 (N_6801,N_6734,N_6706);
and U6802 (N_6802,N_6709,N_6733);
xor U6803 (N_6803,N_6744,N_6764);
or U6804 (N_6804,N_6714,N_6725);
xnor U6805 (N_6805,N_6776,N_6793);
nor U6806 (N_6806,N_6739,N_6710);
and U6807 (N_6807,N_6729,N_6700);
xor U6808 (N_6808,N_6773,N_6770);
nand U6809 (N_6809,N_6727,N_6790);
nor U6810 (N_6810,N_6799,N_6741);
or U6811 (N_6811,N_6759,N_6757);
or U6812 (N_6812,N_6748,N_6747);
or U6813 (N_6813,N_6753,N_6781);
xnor U6814 (N_6814,N_6762,N_6792);
nor U6815 (N_6815,N_6769,N_6794);
and U6816 (N_6816,N_6778,N_6713);
nand U6817 (N_6817,N_6705,N_6701);
xnor U6818 (N_6818,N_6775,N_6761);
xor U6819 (N_6819,N_6708,N_6771);
nor U6820 (N_6820,N_6740,N_6784);
nand U6821 (N_6821,N_6749,N_6787);
xnor U6822 (N_6822,N_6715,N_6758);
nand U6823 (N_6823,N_6719,N_6712);
or U6824 (N_6824,N_6766,N_6751);
or U6825 (N_6825,N_6724,N_6798);
nand U6826 (N_6826,N_6703,N_6716);
nor U6827 (N_6827,N_6726,N_6723);
and U6828 (N_6828,N_6782,N_6738);
xor U6829 (N_6829,N_6718,N_6704);
nand U6830 (N_6830,N_6786,N_6767);
or U6831 (N_6831,N_6750,N_6772);
and U6832 (N_6832,N_6721,N_6765);
xnor U6833 (N_6833,N_6783,N_6797);
or U6834 (N_6834,N_6763,N_6754);
or U6835 (N_6835,N_6737,N_6785);
or U6836 (N_6836,N_6774,N_6796);
and U6837 (N_6837,N_6731,N_6756);
nand U6838 (N_6838,N_6745,N_6728);
or U6839 (N_6839,N_6746,N_6722);
nand U6840 (N_6840,N_6755,N_6791);
nand U6841 (N_6841,N_6743,N_6788);
or U6842 (N_6842,N_6779,N_6780);
xnor U6843 (N_6843,N_6789,N_6742);
xor U6844 (N_6844,N_6795,N_6777);
or U6845 (N_6845,N_6717,N_6707);
xor U6846 (N_6846,N_6732,N_6720);
and U6847 (N_6847,N_6730,N_6760);
and U6848 (N_6848,N_6768,N_6735);
and U6849 (N_6849,N_6711,N_6736);
and U6850 (N_6850,N_6743,N_6784);
or U6851 (N_6851,N_6760,N_6762);
or U6852 (N_6852,N_6740,N_6717);
and U6853 (N_6853,N_6786,N_6737);
xor U6854 (N_6854,N_6748,N_6709);
xnor U6855 (N_6855,N_6740,N_6788);
nor U6856 (N_6856,N_6756,N_6728);
and U6857 (N_6857,N_6776,N_6758);
nor U6858 (N_6858,N_6725,N_6796);
nor U6859 (N_6859,N_6799,N_6735);
or U6860 (N_6860,N_6752,N_6797);
xor U6861 (N_6861,N_6707,N_6702);
and U6862 (N_6862,N_6778,N_6770);
and U6863 (N_6863,N_6751,N_6709);
nor U6864 (N_6864,N_6725,N_6726);
nand U6865 (N_6865,N_6719,N_6786);
and U6866 (N_6866,N_6724,N_6793);
and U6867 (N_6867,N_6775,N_6760);
nand U6868 (N_6868,N_6797,N_6758);
xor U6869 (N_6869,N_6713,N_6757);
nor U6870 (N_6870,N_6737,N_6744);
nand U6871 (N_6871,N_6715,N_6735);
xor U6872 (N_6872,N_6744,N_6771);
xor U6873 (N_6873,N_6767,N_6773);
xor U6874 (N_6874,N_6782,N_6702);
nand U6875 (N_6875,N_6753,N_6700);
nand U6876 (N_6876,N_6705,N_6768);
or U6877 (N_6877,N_6717,N_6748);
nand U6878 (N_6878,N_6784,N_6734);
and U6879 (N_6879,N_6731,N_6759);
and U6880 (N_6880,N_6724,N_6776);
nor U6881 (N_6881,N_6717,N_6771);
nand U6882 (N_6882,N_6752,N_6709);
or U6883 (N_6883,N_6710,N_6793);
xnor U6884 (N_6884,N_6798,N_6753);
xnor U6885 (N_6885,N_6701,N_6752);
and U6886 (N_6886,N_6718,N_6703);
nand U6887 (N_6887,N_6721,N_6730);
xor U6888 (N_6888,N_6756,N_6763);
nor U6889 (N_6889,N_6741,N_6714);
and U6890 (N_6890,N_6768,N_6763);
xor U6891 (N_6891,N_6704,N_6791);
xnor U6892 (N_6892,N_6721,N_6799);
nor U6893 (N_6893,N_6720,N_6753);
and U6894 (N_6894,N_6760,N_6791);
nand U6895 (N_6895,N_6781,N_6744);
nand U6896 (N_6896,N_6793,N_6758);
and U6897 (N_6897,N_6731,N_6739);
xor U6898 (N_6898,N_6748,N_6787);
nand U6899 (N_6899,N_6728,N_6744);
xnor U6900 (N_6900,N_6882,N_6825);
nor U6901 (N_6901,N_6865,N_6859);
nor U6902 (N_6902,N_6888,N_6873);
and U6903 (N_6903,N_6813,N_6847);
and U6904 (N_6904,N_6869,N_6836);
nor U6905 (N_6905,N_6887,N_6858);
and U6906 (N_6906,N_6817,N_6895);
nor U6907 (N_6907,N_6831,N_6848);
or U6908 (N_6908,N_6893,N_6840);
nand U6909 (N_6909,N_6855,N_6883);
nor U6910 (N_6910,N_6896,N_6846);
or U6911 (N_6911,N_6853,N_6800);
and U6912 (N_6912,N_6886,N_6878);
xnor U6913 (N_6913,N_6829,N_6837);
and U6914 (N_6914,N_6826,N_6872);
and U6915 (N_6915,N_6897,N_6870);
nor U6916 (N_6916,N_6818,N_6835);
xnor U6917 (N_6917,N_6832,N_6806);
nor U6918 (N_6918,N_6820,N_6851);
nand U6919 (N_6919,N_6821,N_6889);
nor U6920 (N_6920,N_6849,N_6845);
xnor U6921 (N_6921,N_6808,N_6894);
and U6922 (N_6922,N_6875,N_6876);
nor U6923 (N_6923,N_6854,N_6802);
nor U6924 (N_6924,N_6824,N_6884);
nand U6925 (N_6925,N_6871,N_6843);
nor U6926 (N_6926,N_6804,N_6899);
or U6927 (N_6927,N_6850,N_6857);
nor U6928 (N_6928,N_6863,N_6856);
nand U6929 (N_6929,N_6892,N_6877);
nor U6930 (N_6930,N_6842,N_6866);
xnor U6931 (N_6931,N_6867,N_6880);
or U6932 (N_6932,N_6874,N_6828);
nand U6933 (N_6933,N_6803,N_6898);
nor U6934 (N_6934,N_6861,N_6812);
xnor U6935 (N_6935,N_6868,N_6823);
or U6936 (N_6936,N_6811,N_6816);
nor U6937 (N_6937,N_6890,N_6815);
or U6938 (N_6938,N_6805,N_6822);
nor U6939 (N_6939,N_6834,N_6885);
nand U6940 (N_6940,N_6814,N_6827);
nor U6941 (N_6941,N_6819,N_6864);
or U6942 (N_6942,N_6833,N_6809);
nand U6943 (N_6943,N_6879,N_6862);
and U6944 (N_6944,N_6801,N_6838);
and U6945 (N_6945,N_6810,N_6830);
or U6946 (N_6946,N_6881,N_6839);
nand U6947 (N_6947,N_6841,N_6807);
xor U6948 (N_6948,N_6860,N_6852);
xor U6949 (N_6949,N_6844,N_6891);
xor U6950 (N_6950,N_6844,N_6899);
xnor U6951 (N_6951,N_6809,N_6843);
xnor U6952 (N_6952,N_6802,N_6840);
or U6953 (N_6953,N_6864,N_6811);
nand U6954 (N_6954,N_6833,N_6899);
nor U6955 (N_6955,N_6819,N_6888);
nand U6956 (N_6956,N_6820,N_6838);
nor U6957 (N_6957,N_6868,N_6852);
nand U6958 (N_6958,N_6846,N_6801);
xor U6959 (N_6959,N_6856,N_6882);
or U6960 (N_6960,N_6827,N_6887);
and U6961 (N_6961,N_6840,N_6825);
and U6962 (N_6962,N_6874,N_6801);
or U6963 (N_6963,N_6847,N_6860);
or U6964 (N_6964,N_6813,N_6868);
and U6965 (N_6965,N_6833,N_6854);
or U6966 (N_6966,N_6828,N_6838);
or U6967 (N_6967,N_6818,N_6851);
xnor U6968 (N_6968,N_6859,N_6823);
nor U6969 (N_6969,N_6854,N_6807);
nand U6970 (N_6970,N_6890,N_6878);
nor U6971 (N_6971,N_6872,N_6882);
nor U6972 (N_6972,N_6816,N_6888);
xor U6973 (N_6973,N_6840,N_6879);
nand U6974 (N_6974,N_6875,N_6894);
or U6975 (N_6975,N_6894,N_6822);
xnor U6976 (N_6976,N_6879,N_6852);
xor U6977 (N_6977,N_6827,N_6885);
nor U6978 (N_6978,N_6802,N_6887);
xnor U6979 (N_6979,N_6828,N_6860);
nor U6980 (N_6980,N_6823,N_6827);
nor U6981 (N_6981,N_6814,N_6810);
xor U6982 (N_6982,N_6870,N_6859);
nand U6983 (N_6983,N_6868,N_6863);
nor U6984 (N_6984,N_6895,N_6859);
or U6985 (N_6985,N_6876,N_6879);
and U6986 (N_6986,N_6837,N_6800);
nand U6987 (N_6987,N_6865,N_6878);
nand U6988 (N_6988,N_6845,N_6833);
xnor U6989 (N_6989,N_6833,N_6861);
nand U6990 (N_6990,N_6884,N_6845);
and U6991 (N_6991,N_6814,N_6854);
and U6992 (N_6992,N_6890,N_6898);
and U6993 (N_6993,N_6848,N_6866);
and U6994 (N_6994,N_6877,N_6880);
xnor U6995 (N_6995,N_6893,N_6855);
or U6996 (N_6996,N_6833,N_6810);
and U6997 (N_6997,N_6830,N_6836);
nand U6998 (N_6998,N_6837,N_6893);
nand U6999 (N_6999,N_6887,N_6816);
and U7000 (N_7000,N_6948,N_6918);
xor U7001 (N_7001,N_6906,N_6966);
nand U7002 (N_7002,N_6996,N_6951);
nor U7003 (N_7003,N_6922,N_6911);
and U7004 (N_7004,N_6968,N_6999);
nand U7005 (N_7005,N_6984,N_6923);
and U7006 (N_7006,N_6965,N_6942);
nand U7007 (N_7007,N_6915,N_6931);
nor U7008 (N_7008,N_6946,N_6961);
nand U7009 (N_7009,N_6977,N_6995);
nor U7010 (N_7010,N_6905,N_6909);
nand U7011 (N_7011,N_6932,N_6903);
or U7012 (N_7012,N_6901,N_6970);
nor U7013 (N_7013,N_6907,N_6939);
or U7014 (N_7014,N_6992,N_6954);
nand U7015 (N_7015,N_6971,N_6952);
xor U7016 (N_7016,N_6941,N_6917);
nor U7017 (N_7017,N_6927,N_6964);
or U7018 (N_7018,N_6930,N_6900);
nor U7019 (N_7019,N_6997,N_6963);
and U7020 (N_7020,N_6934,N_6985);
and U7021 (N_7021,N_6945,N_6913);
and U7022 (N_7022,N_6944,N_6975);
xnor U7023 (N_7023,N_6955,N_6983);
xor U7024 (N_7024,N_6926,N_6912);
nand U7025 (N_7025,N_6978,N_6914);
xor U7026 (N_7026,N_6981,N_6976);
or U7027 (N_7027,N_6950,N_6993);
nand U7028 (N_7028,N_6902,N_6933);
and U7029 (N_7029,N_6979,N_6937);
and U7030 (N_7030,N_6910,N_6947);
and U7031 (N_7031,N_6959,N_6972);
or U7032 (N_7032,N_6908,N_6960);
xor U7033 (N_7033,N_6991,N_6943);
xnor U7034 (N_7034,N_6998,N_6990);
or U7035 (N_7035,N_6980,N_6994);
and U7036 (N_7036,N_6920,N_6928);
or U7037 (N_7037,N_6956,N_6940);
nand U7038 (N_7038,N_6936,N_6957);
nand U7039 (N_7039,N_6987,N_6982);
or U7040 (N_7040,N_6958,N_6919);
nand U7041 (N_7041,N_6953,N_6949);
xor U7042 (N_7042,N_6973,N_6967);
nand U7043 (N_7043,N_6929,N_6989);
nor U7044 (N_7044,N_6938,N_6988);
xor U7045 (N_7045,N_6925,N_6904);
xor U7046 (N_7046,N_6935,N_6924);
nand U7047 (N_7047,N_6916,N_6974);
xnor U7048 (N_7048,N_6969,N_6986);
nand U7049 (N_7049,N_6921,N_6962);
or U7050 (N_7050,N_6953,N_6923);
or U7051 (N_7051,N_6986,N_6963);
nor U7052 (N_7052,N_6909,N_6954);
nand U7053 (N_7053,N_6920,N_6900);
xor U7054 (N_7054,N_6981,N_6937);
xnor U7055 (N_7055,N_6968,N_6949);
and U7056 (N_7056,N_6988,N_6918);
or U7057 (N_7057,N_6993,N_6918);
xnor U7058 (N_7058,N_6928,N_6921);
nor U7059 (N_7059,N_6929,N_6962);
xor U7060 (N_7060,N_6977,N_6933);
or U7061 (N_7061,N_6964,N_6947);
nand U7062 (N_7062,N_6902,N_6995);
and U7063 (N_7063,N_6973,N_6995);
or U7064 (N_7064,N_6972,N_6966);
xnor U7065 (N_7065,N_6949,N_6912);
nor U7066 (N_7066,N_6925,N_6973);
and U7067 (N_7067,N_6955,N_6920);
or U7068 (N_7068,N_6955,N_6959);
nor U7069 (N_7069,N_6903,N_6943);
and U7070 (N_7070,N_6993,N_6983);
nor U7071 (N_7071,N_6987,N_6976);
nor U7072 (N_7072,N_6902,N_6958);
and U7073 (N_7073,N_6929,N_6969);
nor U7074 (N_7074,N_6986,N_6910);
nand U7075 (N_7075,N_6926,N_6958);
nor U7076 (N_7076,N_6948,N_6967);
or U7077 (N_7077,N_6973,N_6988);
nand U7078 (N_7078,N_6928,N_6919);
nand U7079 (N_7079,N_6916,N_6969);
and U7080 (N_7080,N_6986,N_6993);
or U7081 (N_7081,N_6942,N_6991);
nand U7082 (N_7082,N_6910,N_6962);
and U7083 (N_7083,N_6988,N_6913);
xor U7084 (N_7084,N_6925,N_6931);
nor U7085 (N_7085,N_6945,N_6979);
or U7086 (N_7086,N_6909,N_6918);
nand U7087 (N_7087,N_6978,N_6962);
or U7088 (N_7088,N_6971,N_6996);
nand U7089 (N_7089,N_6952,N_6931);
nand U7090 (N_7090,N_6926,N_6989);
nor U7091 (N_7091,N_6901,N_6904);
and U7092 (N_7092,N_6945,N_6924);
or U7093 (N_7093,N_6923,N_6937);
xor U7094 (N_7094,N_6917,N_6903);
xor U7095 (N_7095,N_6971,N_6947);
and U7096 (N_7096,N_6992,N_6986);
and U7097 (N_7097,N_6945,N_6948);
xor U7098 (N_7098,N_6926,N_6943);
xor U7099 (N_7099,N_6999,N_6933);
and U7100 (N_7100,N_7024,N_7088);
xnor U7101 (N_7101,N_7004,N_7021);
and U7102 (N_7102,N_7066,N_7002);
nor U7103 (N_7103,N_7038,N_7069);
nand U7104 (N_7104,N_7093,N_7036);
or U7105 (N_7105,N_7040,N_7037);
or U7106 (N_7106,N_7051,N_7027);
xor U7107 (N_7107,N_7011,N_7048);
nand U7108 (N_7108,N_7063,N_7000);
or U7109 (N_7109,N_7030,N_7031);
or U7110 (N_7110,N_7080,N_7059);
xnor U7111 (N_7111,N_7095,N_7001);
and U7112 (N_7112,N_7009,N_7057);
nor U7113 (N_7113,N_7028,N_7097);
nor U7114 (N_7114,N_7065,N_7098);
xnor U7115 (N_7115,N_7055,N_7035);
xor U7116 (N_7116,N_7073,N_7013);
xnor U7117 (N_7117,N_7014,N_7070);
or U7118 (N_7118,N_7020,N_7015);
and U7119 (N_7119,N_7075,N_7086);
and U7120 (N_7120,N_7019,N_7079);
and U7121 (N_7121,N_7096,N_7050);
and U7122 (N_7122,N_7044,N_7023);
nand U7123 (N_7123,N_7033,N_7082);
or U7124 (N_7124,N_7029,N_7076);
and U7125 (N_7125,N_7090,N_7071);
or U7126 (N_7126,N_7092,N_7064);
nor U7127 (N_7127,N_7049,N_7005);
or U7128 (N_7128,N_7026,N_7085);
nor U7129 (N_7129,N_7043,N_7018);
nand U7130 (N_7130,N_7062,N_7025);
nor U7131 (N_7131,N_7006,N_7058);
and U7132 (N_7132,N_7067,N_7012);
or U7133 (N_7133,N_7017,N_7010);
and U7134 (N_7134,N_7099,N_7056);
xor U7135 (N_7135,N_7084,N_7078);
and U7136 (N_7136,N_7061,N_7087);
xnor U7137 (N_7137,N_7047,N_7089);
nor U7138 (N_7138,N_7003,N_7016);
or U7139 (N_7139,N_7039,N_7053);
xnor U7140 (N_7140,N_7041,N_7054);
xnor U7141 (N_7141,N_7022,N_7046);
or U7142 (N_7142,N_7032,N_7074);
nor U7143 (N_7143,N_7072,N_7007);
nand U7144 (N_7144,N_7045,N_7068);
xnor U7145 (N_7145,N_7081,N_7077);
xor U7146 (N_7146,N_7008,N_7034);
nand U7147 (N_7147,N_7042,N_7083);
nor U7148 (N_7148,N_7091,N_7052);
nand U7149 (N_7149,N_7060,N_7094);
nand U7150 (N_7150,N_7050,N_7032);
nor U7151 (N_7151,N_7056,N_7087);
nand U7152 (N_7152,N_7051,N_7015);
nor U7153 (N_7153,N_7014,N_7055);
and U7154 (N_7154,N_7080,N_7043);
nand U7155 (N_7155,N_7047,N_7074);
or U7156 (N_7156,N_7021,N_7091);
xnor U7157 (N_7157,N_7010,N_7041);
nor U7158 (N_7158,N_7031,N_7088);
and U7159 (N_7159,N_7021,N_7026);
xnor U7160 (N_7160,N_7025,N_7009);
xnor U7161 (N_7161,N_7011,N_7056);
and U7162 (N_7162,N_7049,N_7029);
nor U7163 (N_7163,N_7084,N_7016);
xnor U7164 (N_7164,N_7035,N_7049);
nor U7165 (N_7165,N_7056,N_7020);
nand U7166 (N_7166,N_7064,N_7042);
and U7167 (N_7167,N_7001,N_7026);
and U7168 (N_7168,N_7013,N_7030);
nand U7169 (N_7169,N_7094,N_7070);
nand U7170 (N_7170,N_7057,N_7008);
nand U7171 (N_7171,N_7082,N_7044);
and U7172 (N_7172,N_7079,N_7008);
and U7173 (N_7173,N_7069,N_7070);
xor U7174 (N_7174,N_7053,N_7032);
and U7175 (N_7175,N_7029,N_7024);
nand U7176 (N_7176,N_7020,N_7067);
or U7177 (N_7177,N_7094,N_7059);
xnor U7178 (N_7178,N_7059,N_7016);
xor U7179 (N_7179,N_7009,N_7035);
xnor U7180 (N_7180,N_7078,N_7079);
and U7181 (N_7181,N_7052,N_7026);
nor U7182 (N_7182,N_7087,N_7004);
nor U7183 (N_7183,N_7046,N_7062);
nor U7184 (N_7184,N_7013,N_7055);
and U7185 (N_7185,N_7086,N_7053);
or U7186 (N_7186,N_7069,N_7063);
xor U7187 (N_7187,N_7003,N_7066);
nand U7188 (N_7188,N_7069,N_7059);
or U7189 (N_7189,N_7017,N_7078);
xnor U7190 (N_7190,N_7010,N_7089);
nand U7191 (N_7191,N_7096,N_7000);
nand U7192 (N_7192,N_7079,N_7014);
or U7193 (N_7193,N_7082,N_7084);
and U7194 (N_7194,N_7099,N_7088);
xnor U7195 (N_7195,N_7007,N_7039);
nand U7196 (N_7196,N_7042,N_7072);
nand U7197 (N_7197,N_7065,N_7016);
or U7198 (N_7198,N_7095,N_7049);
xnor U7199 (N_7199,N_7054,N_7024);
xnor U7200 (N_7200,N_7164,N_7191);
nand U7201 (N_7201,N_7107,N_7112);
nand U7202 (N_7202,N_7132,N_7116);
nor U7203 (N_7203,N_7162,N_7196);
nand U7204 (N_7204,N_7165,N_7111);
nor U7205 (N_7205,N_7175,N_7156);
or U7206 (N_7206,N_7144,N_7188);
xnor U7207 (N_7207,N_7115,N_7177);
and U7208 (N_7208,N_7185,N_7142);
nand U7209 (N_7209,N_7182,N_7148);
xnor U7210 (N_7210,N_7110,N_7180);
or U7211 (N_7211,N_7150,N_7181);
nand U7212 (N_7212,N_7163,N_7127);
and U7213 (N_7213,N_7179,N_7199);
nor U7214 (N_7214,N_7168,N_7171);
xnor U7215 (N_7215,N_7125,N_7197);
nor U7216 (N_7216,N_7120,N_7134);
and U7217 (N_7217,N_7178,N_7103);
and U7218 (N_7218,N_7131,N_7173);
and U7219 (N_7219,N_7130,N_7135);
nand U7220 (N_7220,N_7198,N_7190);
or U7221 (N_7221,N_7184,N_7146);
and U7222 (N_7222,N_7119,N_7193);
nor U7223 (N_7223,N_7101,N_7151);
xnor U7224 (N_7224,N_7137,N_7114);
nand U7225 (N_7225,N_7195,N_7154);
and U7226 (N_7226,N_7166,N_7157);
or U7227 (N_7227,N_7170,N_7159);
nor U7228 (N_7228,N_7122,N_7128);
nand U7229 (N_7229,N_7187,N_7139);
or U7230 (N_7230,N_7105,N_7186);
nor U7231 (N_7231,N_7192,N_7136);
and U7232 (N_7232,N_7117,N_7169);
or U7233 (N_7233,N_7124,N_7147);
xor U7234 (N_7234,N_7183,N_7160);
nor U7235 (N_7235,N_7152,N_7167);
and U7236 (N_7236,N_7153,N_7189);
xnor U7237 (N_7237,N_7109,N_7126);
nand U7238 (N_7238,N_7158,N_7138);
nand U7239 (N_7239,N_7143,N_7133);
or U7240 (N_7240,N_7123,N_7118);
nor U7241 (N_7241,N_7113,N_7140);
xnor U7242 (N_7242,N_7106,N_7141);
xnor U7243 (N_7243,N_7149,N_7194);
nand U7244 (N_7244,N_7161,N_7174);
nand U7245 (N_7245,N_7155,N_7100);
nor U7246 (N_7246,N_7102,N_7129);
xor U7247 (N_7247,N_7172,N_7121);
and U7248 (N_7248,N_7145,N_7176);
nand U7249 (N_7249,N_7104,N_7108);
or U7250 (N_7250,N_7133,N_7165);
nand U7251 (N_7251,N_7193,N_7160);
nand U7252 (N_7252,N_7106,N_7168);
and U7253 (N_7253,N_7104,N_7178);
or U7254 (N_7254,N_7175,N_7168);
xnor U7255 (N_7255,N_7179,N_7116);
xnor U7256 (N_7256,N_7197,N_7136);
xnor U7257 (N_7257,N_7196,N_7147);
nor U7258 (N_7258,N_7132,N_7152);
or U7259 (N_7259,N_7136,N_7154);
xor U7260 (N_7260,N_7127,N_7110);
or U7261 (N_7261,N_7138,N_7129);
or U7262 (N_7262,N_7167,N_7111);
and U7263 (N_7263,N_7135,N_7120);
xnor U7264 (N_7264,N_7189,N_7175);
nand U7265 (N_7265,N_7140,N_7115);
xnor U7266 (N_7266,N_7130,N_7165);
or U7267 (N_7267,N_7178,N_7100);
nor U7268 (N_7268,N_7169,N_7123);
nor U7269 (N_7269,N_7183,N_7163);
nor U7270 (N_7270,N_7117,N_7183);
nand U7271 (N_7271,N_7121,N_7164);
xnor U7272 (N_7272,N_7180,N_7123);
or U7273 (N_7273,N_7132,N_7154);
nand U7274 (N_7274,N_7162,N_7165);
and U7275 (N_7275,N_7105,N_7120);
and U7276 (N_7276,N_7175,N_7181);
nand U7277 (N_7277,N_7180,N_7109);
nand U7278 (N_7278,N_7165,N_7112);
or U7279 (N_7279,N_7181,N_7122);
xnor U7280 (N_7280,N_7126,N_7180);
nor U7281 (N_7281,N_7147,N_7134);
or U7282 (N_7282,N_7184,N_7165);
xor U7283 (N_7283,N_7191,N_7113);
nand U7284 (N_7284,N_7105,N_7115);
xnor U7285 (N_7285,N_7172,N_7153);
or U7286 (N_7286,N_7191,N_7166);
or U7287 (N_7287,N_7102,N_7164);
nand U7288 (N_7288,N_7123,N_7167);
xor U7289 (N_7289,N_7199,N_7130);
or U7290 (N_7290,N_7160,N_7108);
and U7291 (N_7291,N_7182,N_7117);
xnor U7292 (N_7292,N_7110,N_7186);
nor U7293 (N_7293,N_7193,N_7106);
and U7294 (N_7294,N_7150,N_7125);
or U7295 (N_7295,N_7117,N_7115);
nor U7296 (N_7296,N_7144,N_7158);
and U7297 (N_7297,N_7149,N_7197);
nor U7298 (N_7298,N_7134,N_7143);
nand U7299 (N_7299,N_7172,N_7160);
nor U7300 (N_7300,N_7225,N_7228);
nand U7301 (N_7301,N_7258,N_7221);
nor U7302 (N_7302,N_7240,N_7286);
and U7303 (N_7303,N_7274,N_7268);
xor U7304 (N_7304,N_7233,N_7296);
and U7305 (N_7305,N_7244,N_7235);
nand U7306 (N_7306,N_7298,N_7205);
or U7307 (N_7307,N_7250,N_7276);
and U7308 (N_7308,N_7226,N_7246);
or U7309 (N_7309,N_7253,N_7210);
nor U7310 (N_7310,N_7299,N_7272);
and U7311 (N_7311,N_7290,N_7242);
or U7312 (N_7312,N_7212,N_7245);
nor U7313 (N_7313,N_7247,N_7281);
or U7314 (N_7314,N_7280,N_7275);
and U7315 (N_7315,N_7236,N_7294);
xor U7316 (N_7316,N_7237,N_7252);
nor U7317 (N_7317,N_7289,N_7265);
and U7318 (N_7318,N_7208,N_7215);
nand U7319 (N_7319,N_7264,N_7230);
xnor U7320 (N_7320,N_7219,N_7254);
or U7321 (N_7321,N_7256,N_7224);
xnor U7322 (N_7322,N_7223,N_7232);
or U7323 (N_7323,N_7277,N_7295);
nand U7324 (N_7324,N_7216,N_7266);
xnor U7325 (N_7325,N_7217,N_7202);
and U7326 (N_7326,N_7218,N_7220);
nand U7327 (N_7327,N_7201,N_7292);
xor U7328 (N_7328,N_7227,N_7278);
or U7329 (N_7329,N_7273,N_7270);
xor U7330 (N_7330,N_7238,N_7287);
nand U7331 (N_7331,N_7271,N_7269);
xnor U7332 (N_7332,N_7255,N_7257);
nand U7333 (N_7333,N_7262,N_7248);
or U7334 (N_7334,N_7204,N_7207);
xor U7335 (N_7335,N_7234,N_7261);
and U7336 (N_7336,N_7241,N_7251);
and U7337 (N_7337,N_7263,N_7283);
nand U7338 (N_7338,N_7213,N_7267);
or U7339 (N_7339,N_7239,N_7211);
and U7340 (N_7340,N_7209,N_7243);
nor U7341 (N_7341,N_7259,N_7229);
and U7342 (N_7342,N_7288,N_7293);
xor U7343 (N_7343,N_7200,N_7291);
xor U7344 (N_7344,N_7285,N_7206);
and U7345 (N_7345,N_7260,N_7231);
xor U7346 (N_7346,N_7284,N_7214);
or U7347 (N_7347,N_7249,N_7222);
nor U7348 (N_7348,N_7203,N_7297);
xor U7349 (N_7349,N_7279,N_7282);
xor U7350 (N_7350,N_7278,N_7252);
nand U7351 (N_7351,N_7223,N_7282);
nand U7352 (N_7352,N_7253,N_7235);
xnor U7353 (N_7353,N_7274,N_7278);
xor U7354 (N_7354,N_7203,N_7249);
and U7355 (N_7355,N_7237,N_7227);
nor U7356 (N_7356,N_7240,N_7271);
and U7357 (N_7357,N_7204,N_7278);
or U7358 (N_7358,N_7212,N_7264);
or U7359 (N_7359,N_7224,N_7266);
or U7360 (N_7360,N_7212,N_7202);
xnor U7361 (N_7361,N_7231,N_7290);
nand U7362 (N_7362,N_7227,N_7215);
nand U7363 (N_7363,N_7210,N_7265);
nand U7364 (N_7364,N_7267,N_7287);
xnor U7365 (N_7365,N_7261,N_7298);
nand U7366 (N_7366,N_7273,N_7288);
xnor U7367 (N_7367,N_7271,N_7268);
or U7368 (N_7368,N_7208,N_7283);
and U7369 (N_7369,N_7200,N_7208);
or U7370 (N_7370,N_7236,N_7218);
xnor U7371 (N_7371,N_7293,N_7247);
nor U7372 (N_7372,N_7250,N_7275);
nand U7373 (N_7373,N_7206,N_7202);
and U7374 (N_7374,N_7246,N_7294);
xor U7375 (N_7375,N_7238,N_7227);
nand U7376 (N_7376,N_7268,N_7266);
xor U7377 (N_7377,N_7248,N_7250);
nor U7378 (N_7378,N_7211,N_7260);
or U7379 (N_7379,N_7286,N_7245);
and U7380 (N_7380,N_7272,N_7226);
or U7381 (N_7381,N_7221,N_7247);
and U7382 (N_7382,N_7256,N_7230);
and U7383 (N_7383,N_7235,N_7275);
and U7384 (N_7384,N_7202,N_7262);
xor U7385 (N_7385,N_7229,N_7293);
or U7386 (N_7386,N_7207,N_7212);
nand U7387 (N_7387,N_7236,N_7215);
xor U7388 (N_7388,N_7285,N_7262);
xor U7389 (N_7389,N_7251,N_7220);
nor U7390 (N_7390,N_7286,N_7257);
nor U7391 (N_7391,N_7230,N_7285);
and U7392 (N_7392,N_7297,N_7241);
or U7393 (N_7393,N_7261,N_7278);
nor U7394 (N_7394,N_7225,N_7204);
and U7395 (N_7395,N_7261,N_7240);
nor U7396 (N_7396,N_7280,N_7223);
nor U7397 (N_7397,N_7216,N_7290);
nand U7398 (N_7398,N_7299,N_7297);
and U7399 (N_7399,N_7206,N_7247);
and U7400 (N_7400,N_7307,N_7360);
xnor U7401 (N_7401,N_7345,N_7326);
nand U7402 (N_7402,N_7392,N_7339);
nor U7403 (N_7403,N_7321,N_7368);
xor U7404 (N_7404,N_7300,N_7361);
xnor U7405 (N_7405,N_7377,N_7315);
nor U7406 (N_7406,N_7370,N_7344);
nor U7407 (N_7407,N_7365,N_7375);
or U7408 (N_7408,N_7371,N_7362);
xnor U7409 (N_7409,N_7373,N_7357);
nor U7410 (N_7410,N_7309,N_7396);
nand U7411 (N_7411,N_7343,N_7305);
or U7412 (N_7412,N_7332,N_7322);
nor U7413 (N_7413,N_7383,N_7324);
or U7414 (N_7414,N_7387,N_7359);
nand U7415 (N_7415,N_7313,N_7395);
or U7416 (N_7416,N_7301,N_7353);
or U7417 (N_7417,N_7323,N_7331);
nor U7418 (N_7418,N_7317,N_7372);
xnor U7419 (N_7419,N_7329,N_7378);
and U7420 (N_7420,N_7342,N_7341);
and U7421 (N_7421,N_7367,N_7363);
or U7422 (N_7422,N_7391,N_7312);
xnor U7423 (N_7423,N_7390,N_7310);
or U7424 (N_7424,N_7389,N_7308);
nor U7425 (N_7425,N_7354,N_7348);
and U7426 (N_7426,N_7398,N_7350);
nand U7427 (N_7427,N_7349,N_7318);
nand U7428 (N_7428,N_7330,N_7358);
nand U7429 (N_7429,N_7397,N_7338);
nor U7430 (N_7430,N_7304,N_7320);
or U7431 (N_7431,N_7352,N_7382);
and U7432 (N_7432,N_7316,N_7385);
and U7433 (N_7433,N_7302,N_7347);
nand U7434 (N_7434,N_7346,N_7388);
nor U7435 (N_7435,N_7381,N_7340);
xnor U7436 (N_7436,N_7374,N_7335);
nand U7437 (N_7437,N_7356,N_7334);
nor U7438 (N_7438,N_7337,N_7314);
xnor U7439 (N_7439,N_7366,N_7393);
and U7440 (N_7440,N_7333,N_7336);
and U7441 (N_7441,N_7364,N_7306);
nand U7442 (N_7442,N_7376,N_7369);
and U7443 (N_7443,N_7384,N_7327);
nor U7444 (N_7444,N_7355,N_7303);
nand U7445 (N_7445,N_7319,N_7380);
and U7446 (N_7446,N_7328,N_7379);
and U7447 (N_7447,N_7386,N_7351);
nor U7448 (N_7448,N_7394,N_7311);
and U7449 (N_7449,N_7399,N_7325);
nand U7450 (N_7450,N_7380,N_7361);
xnor U7451 (N_7451,N_7395,N_7322);
nor U7452 (N_7452,N_7310,N_7328);
nor U7453 (N_7453,N_7388,N_7315);
xor U7454 (N_7454,N_7327,N_7385);
nor U7455 (N_7455,N_7367,N_7332);
nand U7456 (N_7456,N_7307,N_7389);
nand U7457 (N_7457,N_7306,N_7390);
and U7458 (N_7458,N_7365,N_7340);
or U7459 (N_7459,N_7313,N_7383);
nand U7460 (N_7460,N_7319,N_7339);
nand U7461 (N_7461,N_7327,N_7316);
or U7462 (N_7462,N_7361,N_7335);
nor U7463 (N_7463,N_7310,N_7363);
and U7464 (N_7464,N_7398,N_7319);
xnor U7465 (N_7465,N_7329,N_7332);
nor U7466 (N_7466,N_7313,N_7341);
xor U7467 (N_7467,N_7343,N_7356);
xor U7468 (N_7468,N_7391,N_7314);
xnor U7469 (N_7469,N_7309,N_7379);
nor U7470 (N_7470,N_7353,N_7313);
nand U7471 (N_7471,N_7346,N_7309);
nand U7472 (N_7472,N_7325,N_7329);
or U7473 (N_7473,N_7398,N_7363);
and U7474 (N_7474,N_7347,N_7306);
nand U7475 (N_7475,N_7303,N_7370);
and U7476 (N_7476,N_7372,N_7388);
or U7477 (N_7477,N_7306,N_7360);
nor U7478 (N_7478,N_7335,N_7360);
nand U7479 (N_7479,N_7370,N_7395);
and U7480 (N_7480,N_7377,N_7347);
nor U7481 (N_7481,N_7359,N_7377);
nand U7482 (N_7482,N_7392,N_7341);
xor U7483 (N_7483,N_7324,N_7360);
nor U7484 (N_7484,N_7320,N_7354);
nand U7485 (N_7485,N_7354,N_7385);
and U7486 (N_7486,N_7305,N_7364);
and U7487 (N_7487,N_7372,N_7381);
and U7488 (N_7488,N_7350,N_7335);
nand U7489 (N_7489,N_7331,N_7310);
or U7490 (N_7490,N_7327,N_7309);
xnor U7491 (N_7491,N_7358,N_7367);
and U7492 (N_7492,N_7387,N_7395);
nor U7493 (N_7493,N_7393,N_7371);
nand U7494 (N_7494,N_7346,N_7318);
xor U7495 (N_7495,N_7394,N_7378);
xor U7496 (N_7496,N_7365,N_7355);
xor U7497 (N_7497,N_7368,N_7323);
and U7498 (N_7498,N_7348,N_7305);
nor U7499 (N_7499,N_7355,N_7302);
xnor U7500 (N_7500,N_7426,N_7423);
nor U7501 (N_7501,N_7497,N_7404);
nand U7502 (N_7502,N_7412,N_7452);
xnor U7503 (N_7503,N_7473,N_7499);
or U7504 (N_7504,N_7446,N_7488);
and U7505 (N_7505,N_7450,N_7493);
and U7506 (N_7506,N_7443,N_7433);
xor U7507 (N_7507,N_7476,N_7491);
xor U7508 (N_7508,N_7448,N_7409);
nand U7509 (N_7509,N_7477,N_7422);
and U7510 (N_7510,N_7451,N_7429);
or U7511 (N_7511,N_7484,N_7425);
or U7512 (N_7512,N_7413,N_7419);
or U7513 (N_7513,N_7495,N_7457);
nand U7514 (N_7514,N_7449,N_7427);
or U7515 (N_7515,N_7424,N_7456);
and U7516 (N_7516,N_7406,N_7474);
nand U7517 (N_7517,N_7432,N_7434);
xnor U7518 (N_7518,N_7469,N_7479);
or U7519 (N_7519,N_7421,N_7441);
nand U7520 (N_7520,N_7407,N_7482);
nor U7521 (N_7521,N_7417,N_7444);
nand U7522 (N_7522,N_7408,N_7416);
xor U7523 (N_7523,N_7405,N_7496);
nand U7524 (N_7524,N_7445,N_7400);
xnor U7525 (N_7525,N_7455,N_7437);
nor U7526 (N_7526,N_7464,N_7489);
nor U7527 (N_7527,N_7498,N_7439);
and U7528 (N_7528,N_7483,N_7466);
and U7529 (N_7529,N_7420,N_7442);
nand U7530 (N_7530,N_7430,N_7460);
xnor U7531 (N_7531,N_7461,N_7494);
or U7532 (N_7532,N_7453,N_7480);
nand U7533 (N_7533,N_7478,N_7435);
or U7534 (N_7534,N_7475,N_7462);
nand U7535 (N_7535,N_7463,N_7485);
and U7536 (N_7536,N_7440,N_7428);
nand U7537 (N_7537,N_7447,N_7410);
or U7538 (N_7538,N_7438,N_7431);
xor U7539 (N_7539,N_7490,N_7487);
xnor U7540 (N_7540,N_7471,N_7486);
nand U7541 (N_7541,N_7470,N_7411);
and U7542 (N_7542,N_7402,N_7414);
xnor U7543 (N_7543,N_7468,N_7401);
or U7544 (N_7544,N_7418,N_7465);
xor U7545 (N_7545,N_7472,N_7403);
xor U7546 (N_7546,N_7459,N_7454);
nor U7547 (N_7547,N_7436,N_7458);
or U7548 (N_7548,N_7467,N_7415);
or U7549 (N_7549,N_7492,N_7481);
xnor U7550 (N_7550,N_7433,N_7494);
and U7551 (N_7551,N_7403,N_7449);
and U7552 (N_7552,N_7488,N_7482);
xor U7553 (N_7553,N_7417,N_7451);
nand U7554 (N_7554,N_7464,N_7415);
xnor U7555 (N_7555,N_7482,N_7486);
xnor U7556 (N_7556,N_7441,N_7498);
or U7557 (N_7557,N_7426,N_7489);
nor U7558 (N_7558,N_7448,N_7461);
nor U7559 (N_7559,N_7440,N_7474);
or U7560 (N_7560,N_7409,N_7444);
nand U7561 (N_7561,N_7434,N_7461);
or U7562 (N_7562,N_7407,N_7408);
xor U7563 (N_7563,N_7415,N_7461);
nand U7564 (N_7564,N_7476,N_7457);
xor U7565 (N_7565,N_7407,N_7499);
or U7566 (N_7566,N_7436,N_7425);
or U7567 (N_7567,N_7480,N_7415);
and U7568 (N_7568,N_7451,N_7498);
and U7569 (N_7569,N_7478,N_7457);
nor U7570 (N_7570,N_7428,N_7493);
and U7571 (N_7571,N_7471,N_7407);
nand U7572 (N_7572,N_7488,N_7439);
and U7573 (N_7573,N_7404,N_7472);
xnor U7574 (N_7574,N_7404,N_7405);
nand U7575 (N_7575,N_7411,N_7478);
and U7576 (N_7576,N_7465,N_7471);
or U7577 (N_7577,N_7406,N_7424);
nor U7578 (N_7578,N_7409,N_7445);
xnor U7579 (N_7579,N_7433,N_7402);
xor U7580 (N_7580,N_7429,N_7490);
or U7581 (N_7581,N_7496,N_7452);
xnor U7582 (N_7582,N_7436,N_7487);
or U7583 (N_7583,N_7455,N_7465);
nor U7584 (N_7584,N_7493,N_7488);
and U7585 (N_7585,N_7450,N_7444);
xnor U7586 (N_7586,N_7418,N_7488);
nand U7587 (N_7587,N_7410,N_7473);
nor U7588 (N_7588,N_7441,N_7474);
or U7589 (N_7589,N_7437,N_7444);
or U7590 (N_7590,N_7466,N_7423);
or U7591 (N_7591,N_7419,N_7455);
nor U7592 (N_7592,N_7407,N_7415);
xnor U7593 (N_7593,N_7422,N_7498);
nand U7594 (N_7594,N_7472,N_7401);
xnor U7595 (N_7595,N_7448,N_7490);
and U7596 (N_7596,N_7406,N_7481);
or U7597 (N_7597,N_7457,N_7440);
or U7598 (N_7598,N_7404,N_7403);
nand U7599 (N_7599,N_7419,N_7449);
and U7600 (N_7600,N_7577,N_7538);
nand U7601 (N_7601,N_7522,N_7558);
nand U7602 (N_7602,N_7588,N_7505);
nor U7603 (N_7603,N_7515,N_7587);
nand U7604 (N_7604,N_7532,N_7525);
and U7605 (N_7605,N_7573,N_7542);
xnor U7606 (N_7606,N_7581,N_7585);
or U7607 (N_7607,N_7544,N_7531);
or U7608 (N_7608,N_7530,N_7503);
xor U7609 (N_7609,N_7528,N_7584);
or U7610 (N_7610,N_7574,N_7561);
nand U7611 (N_7611,N_7580,N_7509);
nor U7612 (N_7612,N_7545,N_7570);
xor U7613 (N_7613,N_7511,N_7567);
nor U7614 (N_7614,N_7516,N_7506);
nand U7615 (N_7615,N_7521,N_7526);
xor U7616 (N_7616,N_7576,N_7514);
or U7617 (N_7617,N_7512,N_7510);
xor U7618 (N_7618,N_7508,N_7583);
nand U7619 (N_7619,N_7593,N_7575);
or U7620 (N_7620,N_7547,N_7537);
nor U7621 (N_7621,N_7571,N_7565);
xnor U7622 (N_7622,N_7549,N_7523);
nand U7623 (N_7623,N_7572,N_7535);
nor U7624 (N_7624,N_7527,N_7539);
nor U7625 (N_7625,N_7598,N_7533);
nor U7626 (N_7626,N_7550,N_7502);
nand U7627 (N_7627,N_7568,N_7529);
or U7628 (N_7628,N_7562,N_7520);
nand U7629 (N_7629,N_7579,N_7595);
nand U7630 (N_7630,N_7540,N_7524);
nand U7631 (N_7631,N_7507,N_7501);
or U7632 (N_7632,N_7541,N_7504);
nor U7633 (N_7633,N_7556,N_7548);
or U7634 (N_7634,N_7590,N_7599);
or U7635 (N_7635,N_7543,N_7563);
nor U7636 (N_7636,N_7534,N_7569);
xor U7637 (N_7637,N_7582,N_7519);
or U7638 (N_7638,N_7554,N_7536);
and U7639 (N_7639,N_7546,N_7551);
or U7640 (N_7640,N_7564,N_7555);
nand U7641 (N_7641,N_7578,N_7592);
xnor U7642 (N_7642,N_7557,N_7596);
xnor U7643 (N_7643,N_7566,N_7597);
or U7644 (N_7644,N_7517,N_7591);
and U7645 (N_7645,N_7559,N_7586);
nand U7646 (N_7646,N_7513,N_7552);
xnor U7647 (N_7647,N_7589,N_7553);
xor U7648 (N_7648,N_7500,N_7518);
xnor U7649 (N_7649,N_7594,N_7560);
nor U7650 (N_7650,N_7524,N_7575);
or U7651 (N_7651,N_7564,N_7593);
or U7652 (N_7652,N_7507,N_7519);
or U7653 (N_7653,N_7553,N_7531);
nand U7654 (N_7654,N_7562,N_7566);
and U7655 (N_7655,N_7579,N_7596);
xnor U7656 (N_7656,N_7567,N_7539);
nand U7657 (N_7657,N_7507,N_7511);
or U7658 (N_7658,N_7561,N_7545);
and U7659 (N_7659,N_7544,N_7525);
nand U7660 (N_7660,N_7569,N_7503);
xnor U7661 (N_7661,N_7533,N_7555);
nor U7662 (N_7662,N_7593,N_7518);
nand U7663 (N_7663,N_7521,N_7506);
nand U7664 (N_7664,N_7560,N_7540);
nor U7665 (N_7665,N_7508,N_7566);
nand U7666 (N_7666,N_7589,N_7555);
xnor U7667 (N_7667,N_7576,N_7596);
or U7668 (N_7668,N_7580,N_7583);
or U7669 (N_7669,N_7536,N_7595);
or U7670 (N_7670,N_7595,N_7522);
nand U7671 (N_7671,N_7568,N_7521);
nor U7672 (N_7672,N_7523,N_7599);
and U7673 (N_7673,N_7553,N_7528);
and U7674 (N_7674,N_7529,N_7507);
xor U7675 (N_7675,N_7508,N_7530);
xor U7676 (N_7676,N_7535,N_7503);
nand U7677 (N_7677,N_7527,N_7515);
or U7678 (N_7678,N_7588,N_7514);
or U7679 (N_7679,N_7563,N_7565);
nand U7680 (N_7680,N_7509,N_7528);
nor U7681 (N_7681,N_7557,N_7567);
or U7682 (N_7682,N_7515,N_7505);
xor U7683 (N_7683,N_7534,N_7550);
xor U7684 (N_7684,N_7599,N_7511);
nand U7685 (N_7685,N_7573,N_7538);
or U7686 (N_7686,N_7553,N_7504);
or U7687 (N_7687,N_7529,N_7582);
and U7688 (N_7688,N_7565,N_7596);
and U7689 (N_7689,N_7595,N_7590);
or U7690 (N_7690,N_7599,N_7538);
nand U7691 (N_7691,N_7563,N_7510);
or U7692 (N_7692,N_7589,N_7566);
xor U7693 (N_7693,N_7554,N_7567);
xor U7694 (N_7694,N_7568,N_7570);
and U7695 (N_7695,N_7542,N_7563);
and U7696 (N_7696,N_7530,N_7544);
xnor U7697 (N_7697,N_7594,N_7548);
nand U7698 (N_7698,N_7559,N_7585);
nand U7699 (N_7699,N_7552,N_7598);
nor U7700 (N_7700,N_7668,N_7697);
and U7701 (N_7701,N_7671,N_7673);
and U7702 (N_7702,N_7694,N_7674);
and U7703 (N_7703,N_7601,N_7698);
nor U7704 (N_7704,N_7679,N_7634);
nor U7705 (N_7705,N_7630,N_7629);
nor U7706 (N_7706,N_7619,N_7669);
nand U7707 (N_7707,N_7696,N_7639);
xor U7708 (N_7708,N_7614,N_7618);
and U7709 (N_7709,N_7627,N_7677);
and U7710 (N_7710,N_7699,N_7670);
xor U7711 (N_7711,N_7605,N_7653);
nor U7712 (N_7712,N_7644,N_7603);
and U7713 (N_7713,N_7636,N_7678);
nand U7714 (N_7714,N_7632,N_7611);
xor U7715 (N_7715,N_7622,N_7667);
xnor U7716 (N_7716,N_7662,N_7672);
or U7717 (N_7717,N_7665,N_7610);
nor U7718 (N_7718,N_7675,N_7650);
xnor U7719 (N_7719,N_7695,N_7623);
or U7720 (N_7720,N_7654,N_7663);
and U7721 (N_7721,N_7621,N_7666);
xor U7722 (N_7722,N_7642,N_7692);
or U7723 (N_7723,N_7649,N_7658);
nor U7724 (N_7724,N_7628,N_7635);
xnor U7725 (N_7725,N_7615,N_7617);
or U7726 (N_7726,N_7633,N_7689);
nor U7727 (N_7727,N_7626,N_7625);
and U7728 (N_7728,N_7606,N_7657);
nor U7729 (N_7729,N_7690,N_7655);
and U7730 (N_7730,N_7609,N_7648);
nand U7731 (N_7731,N_7691,N_7664);
nor U7732 (N_7732,N_7647,N_7612);
nor U7733 (N_7733,N_7660,N_7602);
nand U7734 (N_7734,N_7680,N_7687);
nand U7735 (N_7735,N_7682,N_7604);
and U7736 (N_7736,N_7651,N_7641);
nand U7737 (N_7737,N_7683,N_7616);
or U7738 (N_7738,N_7688,N_7640);
and U7739 (N_7739,N_7620,N_7637);
nand U7740 (N_7740,N_7652,N_7638);
and U7741 (N_7741,N_7643,N_7646);
xnor U7742 (N_7742,N_7600,N_7661);
nand U7743 (N_7743,N_7685,N_7624);
and U7744 (N_7744,N_7608,N_7686);
or U7745 (N_7745,N_7607,N_7656);
nor U7746 (N_7746,N_7693,N_7659);
and U7747 (N_7747,N_7676,N_7681);
nor U7748 (N_7748,N_7613,N_7684);
or U7749 (N_7749,N_7631,N_7645);
and U7750 (N_7750,N_7645,N_7686);
and U7751 (N_7751,N_7617,N_7638);
nand U7752 (N_7752,N_7699,N_7678);
nor U7753 (N_7753,N_7622,N_7675);
nand U7754 (N_7754,N_7650,N_7632);
or U7755 (N_7755,N_7629,N_7625);
and U7756 (N_7756,N_7638,N_7697);
or U7757 (N_7757,N_7611,N_7637);
xnor U7758 (N_7758,N_7688,N_7658);
xnor U7759 (N_7759,N_7652,N_7621);
xnor U7760 (N_7760,N_7654,N_7670);
nor U7761 (N_7761,N_7624,N_7619);
nand U7762 (N_7762,N_7604,N_7679);
nand U7763 (N_7763,N_7671,N_7634);
nor U7764 (N_7764,N_7619,N_7616);
xnor U7765 (N_7765,N_7679,N_7633);
nand U7766 (N_7766,N_7678,N_7618);
or U7767 (N_7767,N_7625,N_7609);
and U7768 (N_7768,N_7619,N_7652);
or U7769 (N_7769,N_7672,N_7613);
and U7770 (N_7770,N_7608,N_7603);
nand U7771 (N_7771,N_7646,N_7693);
and U7772 (N_7772,N_7671,N_7612);
xnor U7773 (N_7773,N_7625,N_7631);
nand U7774 (N_7774,N_7679,N_7632);
xor U7775 (N_7775,N_7658,N_7615);
xor U7776 (N_7776,N_7663,N_7616);
and U7777 (N_7777,N_7614,N_7696);
xor U7778 (N_7778,N_7653,N_7640);
nor U7779 (N_7779,N_7645,N_7638);
nand U7780 (N_7780,N_7699,N_7608);
nor U7781 (N_7781,N_7649,N_7669);
nand U7782 (N_7782,N_7670,N_7624);
nand U7783 (N_7783,N_7665,N_7609);
and U7784 (N_7784,N_7601,N_7691);
or U7785 (N_7785,N_7663,N_7674);
or U7786 (N_7786,N_7602,N_7622);
and U7787 (N_7787,N_7636,N_7657);
and U7788 (N_7788,N_7652,N_7651);
xor U7789 (N_7789,N_7631,N_7604);
nor U7790 (N_7790,N_7678,N_7670);
and U7791 (N_7791,N_7636,N_7614);
or U7792 (N_7792,N_7678,N_7648);
or U7793 (N_7793,N_7627,N_7657);
xor U7794 (N_7794,N_7643,N_7661);
or U7795 (N_7795,N_7693,N_7668);
xnor U7796 (N_7796,N_7637,N_7685);
nor U7797 (N_7797,N_7617,N_7655);
xor U7798 (N_7798,N_7683,N_7693);
and U7799 (N_7799,N_7622,N_7677);
or U7800 (N_7800,N_7744,N_7795);
nand U7801 (N_7801,N_7760,N_7747);
nand U7802 (N_7802,N_7749,N_7781);
nor U7803 (N_7803,N_7707,N_7796);
xnor U7804 (N_7804,N_7730,N_7769);
or U7805 (N_7805,N_7761,N_7743);
and U7806 (N_7806,N_7784,N_7780);
and U7807 (N_7807,N_7778,N_7798);
nor U7808 (N_7808,N_7797,N_7788);
nor U7809 (N_7809,N_7782,N_7776);
nand U7810 (N_7810,N_7792,N_7767);
xor U7811 (N_7811,N_7751,N_7721);
nor U7812 (N_7812,N_7771,N_7736);
nor U7813 (N_7813,N_7762,N_7772);
nor U7814 (N_7814,N_7729,N_7703);
or U7815 (N_7815,N_7706,N_7724);
or U7816 (N_7816,N_7716,N_7741);
and U7817 (N_7817,N_7779,N_7726);
or U7818 (N_7818,N_7756,N_7754);
and U7819 (N_7819,N_7758,N_7725);
nand U7820 (N_7820,N_7700,N_7712);
xor U7821 (N_7821,N_7764,N_7787);
xor U7822 (N_7822,N_7714,N_7799);
xor U7823 (N_7823,N_7757,N_7765);
or U7824 (N_7824,N_7777,N_7702);
nor U7825 (N_7825,N_7735,N_7775);
xnor U7826 (N_7826,N_7718,N_7755);
and U7827 (N_7827,N_7705,N_7745);
nor U7828 (N_7828,N_7783,N_7750);
or U7829 (N_7829,N_7773,N_7733);
and U7830 (N_7830,N_7752,N_7793);
and U7831 (N_7831,N_7731,N_7728);
xor U7832 (N_7832,N_7709,N_7786);
nor U7833 (N_7833,N_7791,N_7734);
nor U7834 (N_7834,N_7766,N_7710);
nor U7835 (N_7835,N_7722,N_7720);
xnor U7836 (N_7836,N_7704,N_7790);
and U7837 (N_7837,N_7732,N_7713);
or U7838 (N_7838,N_7746,N_7715);
or U7839 (N_7839,N_7759,N_7774);
xnor U7840 (N_7840,N_7708,N_7768);
xnor U7841 (N_7841,N_7723,N_7742);
and U7842 (N_7842,N_7794,N_7740);
nor U7843 (N_7843,N_7711,N_7785);
and U7844 (N_7844,N_7770,N_7727);
xnor U7845 (N_7845,N_7763,N_7737);
and U7846 (N_7846,N_7748,N_7719);
and U7847 (N_7847,N_7738,N_7739);
and U7848 (N_7848,N_7701,N_7789);
nor U7849 (N_7849,N_7753,N_7717);
and U7850 (N_7850,N_7771,N_7776);
nor U7851 (N_7851,N_7778,N_7702);
nor U7852 (N_7852,N_7753,N_7739);
nor U7853 (N_7853,N_7774,N_7792);
nor U7854 (N_7854,N_7704,N_7726);
xnor U7855 (N_7855,N_7737,N_7754);
and U7856 (N_7856,N_7741,N_7704);
nand U7857 (N_7857,N_7701,N_7745);
or U7858 (N_7858,N_7700,N_7755);
and U7859 (N_7859,N_7720,N_7768);
nand U7860 (N_7860,N_7723,N_7765);
and U7861 (N_7861,N_7778,N_7786);
nand U7862 (N_7862,N_7737,N_7797);
and U7863 (N_7863,N_7708,N_7795);
xnor U7864 (N_7864,N_7743,N_7768);
xor U7865 (N_7865,N_7755,N_7759);
nand U7866 (N_7866,N_7749,N_7728);
nand U7867 (N_7867,N_7752,N_7765);
xnor U7868 (N_7868,N_7750,N_7706);
nand U7869 (N_7869,N_7773,N_7758);
nor U7870 (N_7870,N_7732,N_7765);
nand U7871 (N_7871,N_7700,N_7715);
or U7872 (N_7872,N_7709,N_7735);
nand U7873 (N_7873,N_7792,N_7715);
xor U7874 (N_7874,N_7775,N_7784);
nand U7875 (N_7875,N_7778,N_7715);
nor U7876 (N_7876,N_7764,N_7710);
and U7877 (N_7877,N_7752,N_7741);
and U7878 (N_7878,N_7765,N_7753);
nor U7879 (N_7879,N_7732,N_7797);
nor U7880 (N_7880,N_7756,N_7791);
nand U7881 (N_7881,N_7739,N_7771);
and U7882 (N_7882,N_7754,N_7753);
nor U7883 (N_7883,N_7772,N_7737);
nor U7884 (N_7884,N_7737,N_7758);
nand U7885 (N_7885,N_7781,N_7710);
xnor U7886 (N_7886,N_7761,N_7746);
and U7887 (N_7887,N_7794,N_7732);
and U7888 (N_7888,N_7792,N_7799);
nand U7889 (N_7889,N_7756,N_7708);
and U7890 (N_7890,N_7722,N_7735);
nor U7891 (N_7891,N_7794,N_7739);
and U7892 (N_7892,N_7746,N_7723);
and U7893 (N_7893,N_7787,N_7720);
or U7894 (N_7894,N_7766,N_7760);
nand U7895 (N_7895,N_7784,N_7759);
nand U7896 (N_7896,N_7753,N_7774);
nor U7897 (N_7897,N_7762,N_7763);
and U7898 (N_7898,N_7757,N_7725);
and U7899 (N_7899,N_7749,N_7780);
and U7900 (N_7900,N_7825,N_7823);
nand U7901 (N_7901,N_7859,N_7897);
or U7902 (N_7902,N_7841,N_7803);
xnor U7903 (N_7903,N_7895,N_7888);
or U7904 (N_7904,N_7804,N_7892);
or U7905 (N_7905,N_7840,N_7843);
or U7906 (N_7906,N_7828,N_7879);
nor U7907 (N_7907,N_7839,N_7865);
nand U7908 (N_7908,N_7827,N_7864);
nor U7909 (N_7909,N_7874,N_7883);
and U7910 (N_7910,N_7800,N_7819);
nor U7911 (N_7911,N_7834,N_7830);
nand U7912 (N_7912,N_7814,N_7816);
or U7913 (N_7913,N_7811,N_7854);
nor U7914 (N_7914,N_7880,N_7875);
or U7915 (N_7915,N_7867,N_7899);
xnor U7916 (N_7916,N_7858,N_7881);
or U7917 (N_7917,N_7852,N_7870);
nor U7918 (N_7918,N_7862,N_7866);
nor U7919 (N_7919,N_7860,N_7877);
or U7920 (N_7920,N_7894,N_7876);
or U7921 (N_7921,N_7855,N_7846);
xor U7922 (N_7922,N_7857,N_7863);
xor U7923 (N_7923,N_7878,N_7849);
nor U7924 (N_7924,N_7842,N_7810);
nand U7925 (N_7925,N_7808,N_7838);
nand U7926 (N_7926,N_7801,N_7833);
nor U7927 (N_7927,N_7821,N_7882);
xnor U7928 (N_7928,N_7805,N_7807);
nor U7929 (N_7929,N_7837,N_7832);
and U7930 (N_7930,N_7891,N_7847);
or U7931 (N_7931,N_7826,N_7884);
or U7932 (N_7932,N_7872,N_7822);
nand U7933 (N_7933,N_7848,N_7851);
and U7934 (N_7934,N_7886,N_7890);
and U7935 (N_7935,N_7861,N_7824);
nor U7936 (N_7936,N_7802,N_7817);
or U7937 (N_7937,N_7829,N_7845);
xnor U7938 (N_7938,N_7856,N_7812);
nand U7939 (N_7939,N_7836,N_7835);
or U7940 (N_7940,N_7844,N_7871);
nand U7941 (N_7941,N_7806,N_7873);
or U7942 (N_7942,N_7869,N_7896);
nor U7943 (N_7943,N_7898,N_7809);
nand U7944 (N_7944,N_7850,N_7831);
nor U7945 (N_7945,N_7818,N_7820);
or U7946 (N_7946,N_7889,N_7815);
and U7947 (N_7947,N_7893,N_7885);
nand U7948 (N_7948,N_7868,N_7853);
nand U7949 (N_7949,N_7887,N_7813);
and U7950 (N_7950,N_7845,N_7813);
nand U7951 (N_7951,N_7864,N_7808);
nor U7952 (N_7952,N_7808,N_7832);
xnor U7953 (N_7953,N_7823,N_7871);
or U7954 (N_7954,N_7806,N_7854);
nand U7955 (N_7955,N_7886,N_7862);
nand U7956 (N_7956,N_7841,N_7810);
nor U7957 (N_7957,N_7802,N_7846);
and U7958 (N_7958,N_7856,N_7875);
xor U7959 (N_7959,N_7825,N_7833);
nand U7960 (N_7960,N_7871,N_7836);
and U7961 (N_7961,N_7896,N_7899);
and U7962 (N_7962,N_7891,N_7848);
nand U7963 (N_7963,N_7831,N_7848);
nor U7964 (N_7964,N_7882,N_7827);
nand U7965 (N_7965,N_7854,N_7896);
or U7966 (N_7966,N_7878,N_7863);
or U7967 (N_7967,N_7810,N_7825);
nor U7968 (N_7968,N_7826,N_7856);
and U7969 (N_7969,N_7870,N_7840);
or U7970 (N_7970,N_7887,N_7804);
or U7971 (N_7971,N_7806,N_7869);
nor U7972 (N_7972,N_7889,N_7850);
or U7973 (N_7973,N_7883,N_7822);
or U7974 (N_7974,N_7857,N_7822);
nand U7975 (N_7975,N_7887,N_7806);
or U7976 (N_7976,N_7827,N_7840);
and U7977 (N_7977,N_7831,N_7809);
nor U7978 (N_7978,N_7858,N_7893);
and U7979 (N_7979,N_7800,N_7869);
xnor U7980 (N_7980,N_7864,N_7837);
nor U7981 (N_7981,N_7826,N_7807);
nand U7982 (N_7982,N_7891,N_7845);
and U7983 (N_7983,N_7844,N_7869);
xor U7984 (N_7984,N_7864,N_7826);
and U7985 (N_7985,N_7885,N_7873);
and U7986 (N_7986,N_7810,N_7830);
xnor U7987 (N_7987,N_7858,N_7859);
xor U7988 (N_7988,N_7885,N_7879);
nand U7989 (N_7989,N_7895,N_7885);
or U7990 (N_7990,N_7809,N_7872);
or U7991 (N_7991,N_7847,N_7835);
or U7992 (N_7992,N_7804,N_7811);
nand U7993 (N_7993,N_7816,N_7882);
xor U7994 (N_7994,N_7804,N_7806);
or U7995 (N_7995,N_7882,N_7838);
xnor U7996 (N_7996,N_7818,N_7839);
nand U7997 (N_7997,N_7847,N_7833);
xor U7998 (N_7998,N_7813,N_7885);
nand U7999 (N_7999,N_7841,N_7856);
or U8000 (N_8000,N_7939,N_7995);
nand U8001 (N_8001,N_7961,N_7986);
xor U8002 (N_8002,N_7931,N_7982);
or U8003 (N_8003,N_7936,N_7908);
xnor U8004 (N_8004,N_7934,N_7944);
or U8005 (N_8005,N_7994,N_7941);
nor U8006 (N_8006,N_7918,N_7924);
nor U8007 (N_8007,N_7921,N_7946);
nor U8008 (N_8008,N_7912,N_7923);
xnor U8009 (N_8009,N_7922,N_7905);
or U8010 (N_8010,N_7926,N_7963);
nor U8011 (N_8011,N_7950,N_7917);
and U8012 (N_8012,N_7956,N_7910);
xor U8013 (N_8013,N_7919,N_7988);
or U8014 (N_8014,N_7999,N_7985);
nor U8015 (N_8015,N_7993,N_7984);
nor U8016 (N_8016,N_7914,N_7955);
nor U8017 (N_8017,N_7940,N_7962);
nand U8018 (N_8018,N_7929,N_7951);
or U8019 (N_8019,N_7987,N_7983);
xor U8020 (N_8020,N_7978,N_7900);
or U8021 (N_8021,N_7954,N_7952);
nand U8022 (N_8022,N_7968,N_7997);
or U8023 (N_8023,N_7901,N_7949);
and U8024 (N_8024,N_7937,N_7948);
nand U8025 (N_8025,N_7915,N_7998);
nand U8026 (N_8026,N_7960,N_7958);
or U8027 (N_8027,N_7916,N_7903);
or U8028 (N_8028,N_7907,N_7964);
and U8029 (N_8029,N_7974,N_7935);
and U8030 (N_8030,N_7959,N_7925);
xor U8031 (N_8031,N_7980,N_7973);
xnor U8032 (N_8032,N_7938,N_7957);
xor U8033 (N_8033,N_7975,N_7911);
and U8034 (N_8034,N_7990,N_7913);
nand U8035 (N_8035,N_7966,N_7945);
nand U8036 (N_8036,N_7920,N_7930);
and U8037 (N_8037,N_7976,N_7989);
and U8038 (N_8038,N_7992,N_7933);
nor U8039 (N_8039,N_7902,N_7981);
xor U8040 (N_8040,N_7977,N_7970);
nor U8041 (N_8041,N_7969,N_7928);
and U8042 (N_8042,N_7904,N_7932);
and U8043 (N_8043,N_7927,N_7909);
nand U8044 (N_8044,N_7947,N_7967);
nand U8045 (N_8045,N_7943,N_7953);
or U8046 (N_8046,N_7972,N_7942);
nor U8047 (N_8047,N_7906,N_7965);
and U8048 (N_8048,N_7996,N_7971);
and U8049 (N_8049,N_7979,N_7991);
and U8050 (N_8050,N_7918,N_7916);
or U8051 (N_8051,N_7977,N_7936);
nand U8052 (N_8052,N_7984,N_7929);
nor U8053 (N_8053,N_7950,N_7901);
xor U8054 (N_8054,N_7996,N_7915);
xor U8055 (N_8055,N_7996,N_7978);
xnor U8056 (N_8056,N_7975,N_7974);
and U8057 (N_8057,N_7951,N_7950);
and U8058 (N_8058,N_7934,N_7930);
nor U8059 (N_8059,N_7985,N_7963);
xnor U8060 (N_8060,N_7930,N_7972);
and U8061 (N_8061,N_7926,N_7984);
and U8062 (N_8062,N_7950,N_7911);
or U8063 (N_8063,N_7991,N_7920);
nand U8064 (N_8064,N_7928,N_7962);
and U8065 (N_8065,N_7998,N_7975);
and U8066 (N_8066,N_7936,N_7998);
or U8067 (N_8067,N_7994,N_7900);
nor U8068 (N_8068,N_7944,N_7905);
and U8069 (N_8069,N_7929,N_7977);
nand U8070 (N_8070,N_7990,N_7994);
xor U8071 (N_8071,N_7907,N_7911);
nor U8072 (N_8072,N_7916,N_7957);
nor U8073 (N_8073,N_7962,N_7970);
and U8074 (N_8074,N_7937,N_7999);
or U8075 (N_8075,N_7962,N_7984);
nand U8076 (N_8076,N_7956,N_7938);
nor U8077 (N_8077,N_7973,N_7965);
xnor U8078 (N_8078,N_7939,N_7953);
nand U8079 (N_8079,N_7982,N_7940);
and U8080 (N_8080,N_7999,N_7911);
or U8081 (N_8081,N_7916,N_7901);
nor U8082 (N_8082,N_7981,N_7988);
nand U8083 (N_8083,N_7961,N_7917);
xor U8084 (N_8084,N_7900,N_7984);
nor U8085 (N_8085,N_7904,N_7963);
and U8086 (N_8086,N_7929,N_7914);
xnor U8087 (N_8087,N_7961,N_7938);
or U8088 (N_8088,N_7979,N_7977);
nand U8089 (N_8089,N_7935,N_7992);
and U8090 (N_8090,N_7991,N_7964);
or U8091 (N_8091,N_7924,N_7964);
or U8092 (N_8092,N_7969,N_7933);
nand U8093 (N_8093,N_7977,N_7973);
nor U8094 (N_8094,N_7906,N_7998);
or U8095 (N_8095,N_7947,N_7916);
nand U8096 (N_8096,N_7926,N_7981);
or U8097 (N_8097,N_7955,N_7990);
nor U8098 (N_8098,N_7911,N_7961);
or U8099 (N_8099,N_7975,N_7934);
nor U8100 (N_8100,N_8018,N_8041);
xnor U8101 (N_8101,N_8033,N_8068);
xnor U8102 (N_8102,N_8061,N_8059);
nor U8103 (N_8103,N_8014,N_8080);
and U8104 (N_8104,N_8028,N_8010);
nor U8105 (N_8105,N_8044,N_8015);
xnor U8106 (N_8106,N_8000,N_8004);
or U8107 (N_8107,N_8078,N_8070);
nand U8108 (N_8108,N_8052,N_8020);
or U8109 (N_8109,N_8003,N_8009);
or U8110 (N_8110,N_8057,N_8049);
xor U8111 (N_8111,N_8096,N_8082);
or U8112 (N_8112,N_8094,N_8038);
nor U8113 (N_8113,N_8050,N_8087);
and U8114 (N_8114,N_8021,N_8005);
and U8115 (N_8115,N_8090,N_8019);
nor U8116 (N_8116,N_8086,N_8079);
nor U8117 (N_8117,N_8013,N_8055);
or U8118 (N_8118,N_8073,N_8025);
xor U8119 (N_8119,N_8043,N_8074);
or U8120 (N_8120,N_8022,N_8062);
nand U8121 (N_8121,N_8042,N_8060);
nand U8122 (N_8122,N_8046,N_8032);
xor U8123 (N_8123,N_8035,N_8002);
or U8124 (N_8124,N_8037,N_8095);
xnor U8125 (N_8125,N_8051,N_8047);
or U8126 (N_8126,N_8006,N_8081);
and U8127 (N_8127,N_8001,N_8026);
xor U8128 (N_8128,N_8024,N_8012);
nor U8129 (N_8129,N_8039,N_8099);
and U8130 (N_8130,N_8008,N_8084);
and U8131 (N_8131,N_8034,N_8011);
or U8132 (N_8132,N_8027,N_8097);
nand U8133 (N_8133,N_8031,N_8029);
and U8134 (N_8134,N_8017,N_8076);
xor U8135 (N_8135,N_8093,N_8098);
xnor U8136 (N_8136,N_8075,N_8036);
nor U8137 (N_8137,N_8056,N_8072);
xnor U8138 (N_8138,N_8091,N_8092);
xor U8139 (N_8139,N_8089,N_8048);
xor U8140 (N_8140,N_8045,N_8064);
nand U8141 (N_8141,N_8088,N_8083);
nand U8142 (N_8142,N_8067,N_8058);
nor U8143 (N_8143,N_8069,N_8077);
and U8144 (N_8144,N_8085,N_8063);
nand U8145 (N_8145,N_8071,N_8007);
and U8146 (N_8146,N_8065,N_8054);
or U8147 (N_8147,N_8030,N_8023);
nor U8148 (N_8148,N_8016,N_8066);
nor U8149 (N_8149,N_8040,N_8053);
nor U8150 (N_8150,N_8082,N_8004);
xnor U8151 (N_8151,N_8065,N_8094);
xor U8152 (N_8152,N_8033,N_8019);
and U8153 (N_8153,N_8073,N_8068);
or U8154 (N_8154,N_8041,N_8074);
or U8155 (N_8155,N_8012,N_8076);
xnor U8156 (N_8156,N_8004,N_8019);
nor U8157 (N_8157,N_8098,N_8087);
and U8158 (N_8158,N_8098,N_8022);
xor U8159 (N_8159,N_8067,N_8044);
or U8160 (N_8160,N_8011,N_8075);
nor U8161 (N_8161,N_8055,N_8096);
nand U8162 (N_8162,N_8041,N_8082);
and U8163 (N_8163,N_8057,N_8043);
or U8164 (N_8164,N_8066,N_8028);
and U8165 (N_8165,N_8071,N_8081);
and U8166 (N_8166,N_8080,N_8023);
or U8167 (N_8167,N_8024,N_8058);
or U8168 (N_8168,N_8012,N_8053);
or U8169 (N_8169,N_8028,N_8078);
nor U8170 (N_8170,N_8023,N_8076);
xor U8171 (N_8171,N_8091,N_8082);
nor U8172 (N_8172,N_8044,N_8080);
and U8173 (N_8173,N_8086,N_8005);
nand U8174 (N_8174,N_8062,N_8078);
nor U8175 (N_8175,N_8046,N_8050);
and U8176 (N_8176,N_8093,N_8074);
and U8177 (N_8177,N_8085,N_8087);
nand U8178 (N_8178,N_8002,N_8003);
and U8179 (N_8179,N_8030,N_8077);
and U8180 (N_8180,N_8086,N_8060);
xor U8181 (N_8181,N_8012,N_8092);
nor U8182 (N_8182,N_8052,N_8010);
nor U8183 (N_8183,N_8087,N_8047);
xor U8184 (N_8184,N_8067,N_8034);
nor U8185 (N_8185,N_8020,N_8017);
nand U8186 (N_8186,N_8090,N_8068);
or U8187 (N_8187,N_8069,N_8042);
nor U8188 (N_8188,N_8045,N_8086);
xnor U8189 (N_8189,N_8091,N_8037);
nand U8190 (N_8190,N_8000,N_8044);
nor U8191 (N_8191,N_8063,N_8081);
nor U8192 (N_8192,N_8071,N_8067);
nor U8193 (N_8193,N_8010,N_8012);
nand U8194 (N_8194,N_8069,N_8093);
nor U8195 (N_8195,N_8015,N_8033);
and U8196 (N_8196,N_8060,N_8046);
nor U8197 (N_8197,N_8092,N_8014);
or U8198 (N_8198,N_8094,N_8003);
nand U8199 (N_8199,N_8027,N_8035);
or U8200 (N_8200,N_8177,N_8102);
nand U8201 (N_8201,N_8198,N_8152);
nand U8202 (N_8202,N_8133,N_8164);
xor U8203 (N_8203,N_8139,N_8100);
nand U8204 (N_8204,N_8147,N_8157);
nand U8205 (N_8205,N_8193,N_8131);
and U8206 (N_8206,N_8109,N_8156);
and U8207 (N_8207,N_8163,N_8170);
nor U8208 (N_8208,N_8107,N_8155);
or U8209 (N_8209,N_8117,N_8140);
nand U8210 (N_8210,N_8116,N_8118);
and U8211 (N_8211,N_8122,N_8101);
nor U8212 (N_8212,N_8148,N_8180);
and U8213 (N_8213,N_8144,N_8153);
or U8214 (N_8214,N_8127,N_8136);
nor U8215 (N_8215,N_8128,N_8108);
or U8216 (N_8216,N_8125,N_8197);
or U8217 (N_8217,N_8151,N_8146);
nand U8218 (N_8218,N_8134,N_8114);
or U8219 (N_8219,N_8112,N_8103);
xnor U8220 (N_8220,N_8124,N_8135);
or U8221 (N_8221,N_8104,N_8175);
nor U8222 (N_8222,N_8169,N_8154);
or U8223 (N_8223,N_8161,N_8115);
nor U8224 (N_8224,N_8191,N_8126);
or U8225 (N_8225,N_8187,N_8188);
nand U8226 (N_8226,N_8159,N_8137);
nor U8227 (N_8227,N_8168,N_8184);
and U8228 (N_8228,N_8179,N_8183);
xor U8229 (N_8229,N_8194,N_8120);
or U8230 (N_8230,N_8165,N_8113);
nor U8231 (N_8231,N_8119,N_8174);
and U8232 (N_8232,N_8171,N_8199);
nor U8233 (N_8233,N_8158,N_8178);
xor U8234 (N_8234,N_8138,N_8142);
nor U8235 (N_8235,N_8149,N_8173);
nand U8236 (N_8236,N_8176,N_8162);
nand U8237 (N_8237,N_8166,N_8132);
and U8238 (N_8238,N_8182,N_8141);
and U8239 (N_8239,N_8111,N_8105);
and U8240 (N_8240,N_8130,N_8121);
or U8241 (N_8241,N_8150,N_8110);
and U8242 (N_8242,N_8129,N_8145);
nand U8243 (N_8243,N_8190,N_8172);
or U8244 (N_8244,N_8181,N_8196);
and U8245 (N_8245,N_8143,N_8167);
and U8246 (N_8246,N_8186,N_8160);
xor U8247 (N_8247,N_8123,N_8195);
or U8248 (N_8248,N_8189,N_8192);
nor U8249 (N_8249,N_8185,N_8106);
nand U8250 (N_8250,N_8106,N_8131);
or U8251 (N_8251,N_8139,N_8127);
nand U8252 (N_8252,N_8163,N_8144);
xnor U8253 (N_8253,N_8144,N_8147);
or U8254 (N_8254,N_8189,N_8167);
or U8255 (N_8255,N_8126,N_8177);
or U8256 (N_8256,N_8198,N_8196);
xnor U8257 (N_8257,N_8109,N_8193);
xnor U8258 (N_8258,N_8159,N_8135);
or U8259 (N_8259,N_8171,N_8155);
or U8260 (N_8260,N_8193,N_8151);
or U8261 (N_8261,N_8145,N_8168);
nand U8262 (N_8262,N_8170,N_8162);
nor U8263 (N_8263,N_8186,N_8131);
xnor U8264 (N_8264,N_8144,N_8121);
xor U8265 (N_8265,N_8116,N_8125);
xnor U8266 (N_8266,N_8142,N_8103);
and U8267 (N_8267,N_8121,N_8170);
nor U8268 (N_8268,N_8190,N_8145);
or U8269 (N_8269,N_8106,N_8181);
nor U8270 (N_8270,N_8152,N_8172);
and U8271 (N_8271,N_8134,N_8188);
or U8272 (N_8272,N_8147,N_8128);
and U8273 (N_8273,N_8192,N_8126);
and U8274 (N_8274,N_8155,N_8189);
xor U8275 (N_8275,N_8133,N_8193);
nor U8276 (N_8276,N_8114,N_8115);
or U8277 (N_8277,N_8157,N_8107);
xnor U8278 (N_8278,N_8132,N_8157);
and U8279 (N_8279,N_8123,N_8156);
and U8280 (N_8280,N_8152,N_8139);
and U8281 (N_8281,N_8179,N_8187);
nor U8282 (N_8282,N_8111,N_8126);
or U8283 (N_8283,N_8177,N_8108);
nand U8284 (N_8284,N_8161,N_8167);
nand U8285 (N_8285,N_8161,N_8104);
and U8286 (N_8286,N_8128,N_8126);
nor U8287 (N_8287,N_8143,N_8123);
xnor U8288 (N_8288,N_8191,N_8141);
or U8289 (N_8289,N_8117,N_8112);
nand U8290 (N_8290,N_8109,N_8119);
xor U8291 (N_8291,N_8182,N_8194);
xor U8292 (N_8292,N_8173,N_8137);
nand U8293 (N_8293,N_8129,N_8189);
or U8294 (N_8294,N_8106,N_8116);
or U8295 (N_8295,N_8156,N_8178);
nand U8296 (N_8296,N_8187,N_8107);
and U8297 (N_8297,N_8146,N_8161);
xnor U8298 (N_8298,N_8106,N_8136);
and U8299 (N_8299,N_8173,N_8157);
nor U8300 (N_8300,N_8209,N_8289);
nor U8301 (N_8301,N_8284,N_8269);
and U8302 (N_8302,N_8275,N_8239);
nor U8303 (N_8303,N_8254,N_8272);
nand U8304 (N_8304,N_8235,N_8286);
or U8305 (N_8305,N_8212,N_8291);
or U8306 (N_8306,N_8297,N_8264);
and U8307 (N_8307,N_8270,N_8253);
and U8308 (N_8308,N_8206,N_8279);
xor U8309 (N_8309,N_8220,N_8203);
and U8310 (N_8310,N_8233,N_8245);
nor U8311 (N_8311,N_8295,N_8277);
nor U8312 (N_8312,N_8221,N_8256);
nor U8313 (N_8313,N_8283,N_8280);
and U8314 (N_8314,N_8200,N_8262);
nor U8315 (N_8315,N_8230,N_8225);
xnor U8316 (N_8316,N_8274,N_8266);
and U8317 (N_8317,N_8278,N_8271);
and U8318 (N_8318,N_8282,N_8268);
or U8319 (N_8319,N_8213,N_8241);
and U8320 (N_8320,N_8219,N_8251);
nand U8321 (N_8321,N_8255,N_8208);
nand U8322 (N_8322,N_8248,N_8226);
or U8323 (N_8323,N_8201,N_8257);
and U8324 (N_8324,N_8234,N_8218);
nor U8325 (N_8325,N_8246,N_8242);
xnor U8326 (N_8326,N_8252,N_8227);
or U8327 (N_8327,N_8236,N_8231);
or U8328 (N_8328,N_8215,N_8267);
nor U8329 (N_8329,N_8228,N_8294);
nand U8330 (N_8330,N_8240,N_8216);
nand U8331 (N_8331,N_8232,N_8276);
nand U8332 (N_8332,N_8288,N_8204);
or U8333 (N_8333,N_8237,N_8290);
nor U8334 (N_8334,N_8210,N_8287);
or U8335 (N_8335,N_8258,N_8285);
or U8336 (N_8336,N_8224,N_8273);
and U8337 (N_8337,N_8229,N_8299);
nand U8338 (N_8338,N_8261,N_8244);
nand U8339 (N_8339,N_8247,N_8238);
and U8340 (N_8340,N_8292,N_8202);
xnor U8341 (N_8341,N_8296,N_8205);
xnor U8342 (N_8342,N_8249,N_8250);
nor U8343 (N_8343,N_8223,N_8263);
nor U8344 (N_8344,N_8265,N_8293);
nor U8345 (N_8345,N_8211,N_8281);
and U8346 (N_8346,N_8207,N_8217);
and U8347 (N_8347,N_8243,N_8298);
or U8348 (N_8348,N_8214,N_8260);
xnor U8349 (N_8349,N_8259,N_8222);
nand U8350 (N_8350,N_8209,N_8288);
xnor U8351 (N_8351,N_8270,N_8211);
and U8352 (N_8352,N_8263,N_8225);
nor U8353 (N_8353,N_8242,N_8214);
or U8354 (N_8354,N_8270,N_8291);
and U8355 (N_8355,N_8242,N_8280);
nand U8356 (N_8356,N_8274,N_8298);
nor U8357 (N_8357,N_8241,N_8275);
and U8358 (N_8358,N_8287,N_8298);
and U8359 (N_8359,N_8238,N_8232);
nand U8360 (N_8360,N_8271,N_8217);
nor U8361 (N_8361,N_8291,N_8211);
nand U8362 (N_8362,N_8266,N_8217);
and U8363 (N_8363,N_8272,N_8209);
or U8364 (N_8364,N_8298,N_8252);
xor U8365 (N_8365,N_8214,N_8280);
nor U8366 (N_8366,N_8258,N_8204);
or U8367 (N_8367,N_8299,N_8211);
and U8368 (N_8368,N_8250,N_8213);
and U8369 (N_8369,N_8202,N_8221);
and U8370 (N_8370,N_8298,N_8203);
or U8371 (N_8371,N_8244,N_8201);
xnor U8372 (N_8372,N_8231,N_8247);
and U8373 (N_8373,N_8258,N_8226);
or U8374 (N_8374,N_8233,N_8228);
and U8375 (N_8375,N_8274,N_8280);
xor U8376 (N_8376,N_8291,N_8214);
nand U8377 (N_8377,N_8211,N_8236);
nand U8378 (N_8378,N_8261,N_8232);
or U8379 (N_8379,N_8206,N_8291);
and U8380 (N_8380,N_8268,N_8239);
nor U8381 (N_8381,N_8212,N_8237);
and U8382 (N_8382,N_8227,N_8262);
nand U8383 (N_8383,N_8230,N_8297);
or U8384 (N_8384,N_8218,N_8285);
or U8385 (N_8385,N_8232,N_8297);
nor U8386 (N_8386,N_8226,N_8275);
nor U8387 (N_8387,N_8226,N_8252);
xor U8388 (N_8388,N_8248,N_8220);
nor U8389 (N_8389,N_8296,N_8273);
xnor U8390 (N_8390,N_8286,N_8269);
and U8391 (N_8391,N_8271,N_8211);
and U8392 (N_8392,N_8264,N_8298);
or U8393 (N_8393,N_8263,N_8275);
xor U8394 (N_8394,N_8252,N_8273);
or U8395 (N_8395,N_8204,N_8240);
and U8396 (N_8396,N_8286,N_8255);
nand U8397 (N_8397,N_8250,N_8245);
xnor U8398 (N_8398,N_8299,N_8236);
xnor U8399 (N_8399,N_8266,N_8218);
and U8400 (N_8400,N_8379,N_8354);
or U8401 (N_8401,N_8306,N_8334);
xor U8402 (N_8402,N_8330,N_8392);
xnor U8403 (N_8403,N_8322,N_8359);
and U8404 (N_8404,N_8372,N_8373);
and U8405 (N_8405,N_8376,N_8309);
nand U8406 (N_8406,N_8367,N_8333);
xor U8407 (N_8407,N_8363,N_8349);
nor U8408 (N_8408,N_8331,N_8353);
or U8409 (N_8409,N_8320,N_8312);
or U8410 (N_8410,N_8303,N_8381);
and U8411 (N_8411,N_8326,N_8339);
or U8412 (N_8412,N_8399,N_8397);
nand U8413 (N_8413,N_8348,N_8338);
and U8414 (N_8414,N_8398,N_8346);
nor U8415 (N_8415,N_8323,N_8384);
and U8416 (N_8416,N_8393,N_8318);
nand U8417 (N_8417,N_8394,N_8345);
or U8418 (N_8418,N_8355,N_8328);
nand U8419 (N_8419,N_8307,N_8341);
nor U8420 (N_8420,N_8327,N_8332);
nor U8421 (N_8421,N_8357,N_8377);
and U8422 (N_8422,N_8383,N_8308);
nor U8423 (N_8423,N_8311,N_8321);
or U8424 (N_8424,N_8370,N_8368);
xor U8425 (N_8425,N_8387,N_8364);
or U8426 (N_8426,N_8386,N_8380);
nor U8427 (N_8427,N_8324,N_8350);
nor U8428 (N_8428,N_8371,N_8391);
or U8429 (N_8429,N_8329,N_8302);
or U8430 (N_8430,N_8314,N_8390);
nand U8431 (N_8431,N_8356,N_8382);
or U8432 (N_8432,N_8336,N_8347);
or U8433 (N_8433,N_8378,N_8343);
and U8434 (N_8434,N_8315,N_8365);
xnor U8435 (N_8435,N_8310,N_8388);
nor U8436 (N_8436,N_8301,N_8340);
nand U8437 (N_8437,N_8352,N_8389);
nand U8438 (N_8438,N_8316,N_8317);
or U8439 (N_8439,N_8342,N_8358);
and U8440 (N_8440,N_8351,N_8385);
nor U8441 (N_8441,N_8361,N_8369);
xnor U8442 (N_8442,N_8396,N_8300);
nand U8443 (N_8443,N_8362,N_8374);
or U8444 (N_8444,N_8325,N_8344);
nor U8445 (N_8445,N_8313,N_8305);
nand U8446 (N_8446,N_8395,N_8319);
or U8447 (N_8447,N_8304,N_8360);
xor U8448 (N_8448,N_8337,N_8375);
or U8449 (N_8449,N_8366,N_8335);
or U8450 (N_8450,N_8347,N_8325);
or U8451 (N_8451,N_8303,N_8341);
xor U8452 (N_8452,N_8306,N_8319);
nor U8453 (N_8453,N_8383,N_8342);
xnor U8454 (N_8454,N_8378,N_8369);
and U8455 (N_8455,N_8313,N_8341);
xor U8456 (N_8456,N_8330,N_8340);
nor U8457 (N_8457,N_8312,N_8347);
and U8458 (N_8458,N_8311,N_8397);
and U8459 (N_8459,N_8380,N_8332);
nand U8460 (N_8460,N_8350,N_8312);
nor U8461 (N_8461,N_8352,N_8314);
xnor U8462 (N_8462,N_8399,N_8335);
nand U8463 (N_8463,N_8312,N_8331);
nand U8464 (N_8464,N_8356,N_8319);
and U8465 (N_8465,N_8320,N_8332);
nand U8466 (N_8466,N_8349,N_8371);
or U8467 (N_8467,N_8312,N_8303);
and U8468 (N_8468,N_8361,N_8346);
xnor U8469 (N_8469,N_8311,N_8335);
xor U8470 (N_8470,N_8349,N_8394);
xnor U8471 (N_8471,N_8334,N_8391);
nor U8472 (N_8472,N_8383,N_8320);
nand U8473 (N_8473,N_8318,N_8376);
nand U8474 (N_8474,N_8386,N_8330);
or U8475 (N_8475,N_8347,N_8373);
nand U8476 (N_8476,N_8378,N_8316);
nor U8477 (N_8477,N_8343,N_8360);
and U8478 (N_8478,N_8336,N_8399);
nand U8479 (N_8479,N_8319,N_8349);
or U8480 (N_8480,N_8356,N_8395);
or U8481 (N_8481,N_8328,N_8378);
xor U8482 (N_8482,N_8344,N_8316);
and U8483 (N_8483,N_8381,N_8370);
nor U8484 (N_8484,N_8323,N_8388);
or U8485 (N_8485,N_8316,N_8350);
xor U8486 (N_8486,N_8343,N_8359);
nand U8487 (N_8487,N_8377,N_8304);
or U8488 (N_8488,N_8308,N_8365);
nand U8489 (N_8489,N_8358,N_8373);
xnor U8490 (N_8490,N_8390,N_8331);
nor U8491 (N_8491,N_8381,N_8397);
nor U8492 (N_8492,N_8304,N_8320);
nor U8493 (N_8493,N_8337,N_8358);
and U8494 (N_8494,N_8324,N_8304);
xor U8495 (N_8495,N_8319,N_8379);
nor U8496 (N_8496,N_8351,N_8300);
or U8497 (N_8497,N_8325,N_8367);
nor U8498 (N_8498,N_8328,N_8344);
or U8499 (N_8499,N_8369,N_8362);
or U8500 (N_8500,N_8443,N_8419);
and U8501 (N_8501,N_8477,N_8431);
nand U8502 (N_8502,N_8469,N_8488);
nand U8503 (N_8503,N_8448,N_8491);
or U8504 (N_8504,N_8406,N_8497);
and U8505 (N_8505,N_8430,N_8420);
nand U8506 (N_8506,N_8499,N_8471);
xor U8507 (N_8507,N_8427,N_8466);
and U8508 (N_8508,N_8454,N_8439);
and U8509 (N_8509,N_8445,N_8459);
and U8510 (N_8510,N_8412,N_8464);
or U8511 (N_8511,N_8403,N_8410);
or U8512 (N_8512,N_8467,N_8409);
nor U8513 (N_8513,N_8493,N_8438);
nor U8514 (N_8514,N_8475,N_8463);
nor U8515 (N_8515,N_8444,N_8436);
nor U8516 (N_8516,N_8429,N_8424);
and U8517 (N_8517,N_8452,N_8423);
nor U8518 (N_8518,N_8442,N_8451);
or U8519 (N_8519,N_8405,N_8449);
or U8520 (N_8520,N_8489,N_8411);
nand U8521 (N_8521,N_8418,N_8421);
nor U8522 (N_8522,N_8441,N_8458);
or U8523 (N_8523,N_8447,N_8422);
and U8524 (N_8524,N_8428,N_8415);
or U8525 (N_8525,N_8446,N_8496);
nand U8526 (N_8526,N_8416,N_8432);
xnor U8527 (N_8527,N_8479,N_8465);
xnor U8528 (N_8528,N_8478,N_8484);
and U8529 (N_8529,N_8482,N_8435);
nand U8530 (N_8530,N_8461,N_8470);
nor U8531 (N_8531,N_8460,N_8473);
nand U8532 (N_8532,N_8485,N_8414);
and U8533 (N_8533,N_8453,N_8404);
and U8534 (N_8534,N_8455,N_8456);
nand U8535 (N_8535,N_8407,N_8425);
and U8536 (N_8536,N_8437,N_8495);
nand U8537 (N_8537,N_8490,N_8400);
nor U8538 (N_8538,N_8462,N_8413);
or U8539 (N_8539,N_8498,N_8408);
nor U8540 (N_8540,N_8401,N_8417);
and U8541 (N_8541,N_8486,N_8492);
nor U8542 (N_8542,N_8450,N_8480);
nand U8543 (N_8543,N_8457,N_8468);
or U8544 (N_8544,N_8481,N_8487);
or U8545 (N_8545,N_8426,N_8483);
nand U8546 (N_8546,N_8474,N_8433);
xnor U8547 (N_8547,N_8472,N_8434);
xnor U8548 (N_8548,N_8402,N_8476);
nand U8549 (N_8549,N_8440,N_8494);
xnor U8550 (N_8550,N_8488,N_8425);
and U8551 (N_8551,N_8434,N_8493);
xor U8552 (N_8552,N_8423,N_8415);
nand U8553 (N_8553,N_8407,N_8463);
nor U8554 (N_8554,N_8414,N_8467);
xor U8555 (N_8555,N_8431,N_8440);
and U8556 (N_8556,N_8491,N_8484);
or U8557 (N_8557,N_8446,N_8486);
xor U8558 (N_8558,N_8434,N_8459);
or U8559 (N_8559,N_8498,N_8402);
nor U8560 (N_8560,N_8489,N_8456);
and U8561 (N_8561,N_8451,N_8496);
nor U8562 (N_8562,N_8453,N_8440);
and U8563 (N_8563,N_8475,N_8495);
xor U8564 (N_8564,N_8466,N_8489);
nor U8565 (N_8565,N_8427,N_8499);
and U8566 (N_8566,N_8412,N_8456);
xnor U8567 (N_8567,N_8419,N_8471);
nand U8568 (N_8568,N_8481,N_8436);
and U8569 (N_8569,N_8461,N_8433);
xor U8570 (N_8570,N_8466,N_8434);
and U8571 (N_8571,N_8435,N_8450);
and U8572 (N_8572,N_8455,N_8408);
and U8573 (N_8573,N_8470,N_8486);
or U8574 (N_8574,N_8408,N_8477);
or U8575 (N_8575,N_8445,N_8419);
nor U8576 (N_8576,N_8419,N_8456);
or U8577 (N_8577,N_8458,N_8437);
or U8578 (N_8578,N_8453,N_8402);
or U8579 (N_8579,N_8498,N_8467);
nor U8580 (N_8580,N_8475,N_8490);
and U8581 (N_8581,N_8478,N_8447);
xnor U8582 (N_8582,N_8411,N_8407);
xnor U8583 (N_8583,N_8405,N_8450);
or U8584 (N_8584,N_8403,N_8472);
and U8585 (N_8585,N_8433,N_8479);
xnor U8586 (N_8586,N_8404,N_8437);
and U8587 (N_8587,N_8475,N_8427);
nand U8588 (N_8588,N_8401,N_8419);
and U8589 (N_8589,N_8405,N_8409);
nor U8590 (N_8590,N_8443,N_8499);
xnor U8591 (N_8591,N_8413,N_8466);
xnor U8592 (N_8592,N_8494,N_8400);
xor U8593 (N_8593,N_8464,N_8445);
and U8594 (N_8594,N_8449,N_8451);
nor U8595 (N_8595,N_8493,N_8483);
or U8596 (N_8596,N_8425,N_8458);
xnor U8597 (N_8597,N_8417,N_8444);
nand U8598 (N_8598,N_8448,N_8442);
xnor U8599 (N_8599,N_8430,N_8444);
xnor U8600 (N_8600,N_8536,N_8585);
or U8601 (N_8601,N_8553,N_8587);
or U8602 (N_8602,N_8582,N_8505);
xor U8603 (N_8603,N_8573,N_8520);
or U8604 (N_8604,N_8535,N_8533);
xnor U8605 (N_8605,N_8547,N_8576);
nor U8606 (N_8606,N_8597,N_8593);
or U8607 (N_8607,N_8529,N_8530);
nor U8608 (N_8608,N_8524,N_8516);
and U8609 (N_8609,N_8564,N_8534);
and U8610 (N_8610,N_8518,N_8548);
xnor U8611 (N_8611,N_8571,N_8592);
or U8612 (N_8612,N_8565,N_8567);
xor U8613 (N_8613,N_8577,N_8523);
or U8614 (N_8614,N_8583,N_8508);
xnor U8615 (N_8615,N_8570,N_8588);
nand U8616 (N_8616,N_8537,N_8580);
nor U8617 (N_8617,N_8541,N_8558);
xor U8618 (N_8618,N_8584,N_8557);
or U8619 (N_8619,N_8568,N_8543);
or U8620 (N_8620,N_8532,N_8554);
and U8621 (N_8621,N_8539,N_8544);
nor U8622 (N_8622,N_8515,N_8578);
nand U8623 (N_8623,N_8531,N_8510);
xnor U8624 (N_8624,N_8589,N_8598);
nand U8625 (N_8625,N_8575,N_8512);
and U8626 (N_8626,N_8560,N_8513);
nor U8627 (N_8627,N_8522,N_8507);
or U8628 (N_8628,N_8549,N_8519);
nand U8629 (N_8629,N_8506,N_8555);
xnor U8630 (N_8630,N_8546,N_8562);
and U8631 (N_8631,N_8503,N_8552);
nand U8632 (N_8632,N_8590,N_8509);
or U8633 (N_8633,N_8591,N_8569);
or U8634 (N_8634,N_8502,N_8517);
and U8635 (N_8635,N_8563,N_8594);
nor U8636 (N_8636,N_8538,N_8525);
nor U8637 (N_8637,N_8551,N_8511);
xor U8638 (N_8638,N_8542,N_8527);
or U8639 (N_8639,N_8521,N_8572);
nor U8640 (N_8640,N_8514,N_8545);
and U8641 (N_8641,N_8579,N_8528);
nand U8642 (N_8642,N_8599,N_8500);
or U8643 (N_8643,N_8540,N_8595);
nor U8644 (N_8644,N_8526,N_8559);
xor U8645 (N_8645,N_8550,N_8586);
or U8646 (N_8646,N_8501,N_8504);
nor U8647 (N_8647,N_8596,N_8574);
nand U8648 (N_8648,N_8581,N_8556);
nor U8649 (N_8649,N_8566,N_8561);
or U8650 (N_8650,N_8536,N_8563);
xor U8651 (N_8651,N_8529,N_8560);
nor U8652 (N_8652,N_8531,N_8591);
nand U8653 (N_8653,N_8574,N_8550);
nor U8654 (N_8654,N_8581,N_8567);
and U8655 (N_8655,N_8515,N_8517);
and U8656 (N_8656,N_8520,N_8538);
nand U8657 (N_8657,N_8597,N_8572);
and U8658 (N_8658,N_8505,N_8529);
and U8659 (N_8659,N_8548,N_8569);
xnor U8660 (N_8660,N_8586,N_8516);
nand U8661 (N_8661,N_8568,N_8512);
or U8662 (N_8662,N_8543,N_8596);
and U8663 (N_8663,N_8513,N_8561);
xnor U8664 (N_8664,N_8583,N_8527);
and U8665 (N_8665,N_8507,N_8526);
xnor U8666 (N_8666,N_8530,N_8565);
or U8667 (N_8667,N_8518,N_8574);
xnor U8668 (N_8668,N_8570,N_8530);
and U8669 (N_8669,N_8521,N_8541);
nor U8670 (N_8670,N_8522,N_8545);
and U8671 (N_8671,N_8528,N_8545);
or U8672 (N_8672,N_8563,N_8590);
nor U8673 (N_8673,N_8598,N_8511);
xnor U8674 (N_8674,N_8516,N_8573);
nor U8675 (N_8675,N_8588,N_8563);
xnor U8676 (N_8676,N_8579,N_8554);
nand U8677 (N_8677,N_8567,N_8525);
nor U8678 (N_8678,N_8596,N_8591);
or U8679 (N_8679,N_8581,N_8548);
and U8680 (N_8680,N_8520,N_8563);
nor U8681 (N_8681,N_8567,N_8548);
nor U8682 (N_8682,N_8552,N_8581);
and U8683 (N_8683,N_8502,N_8539);
and U8684 (N_8684,N_8538,N_8539);
or U8685 (N_8685,N_8575,N_8522);
and U8686 (N_8686,N_8596,N_8517);
nand U8687 (N_8687,N_8594,N_8547);
or U8688 (N_8688,N_8595,N_8509);
or U8689 (N_8689,N_8570,N_8594);
or U8690 (N_8690,N_8577,N_8567);
nand U8691 (N_8691,N_8575,N_8561);
or U8692 (N_8692,N_8501,N_8589);
and U8693 (N_8693,N_8570,N_8546);
and U8694 (N_8694,N_8537,N_8573);
and U8695 (N_8695,N_8505,N_8579);
nor U8696 (N_8696,N_8536,N_8566);
nor U8697 (N_8697,N_8511,N_8590);
or U8698 (N_8698,N_8566,N_8509);
or U8699 (N_8699,N_8529,N_8534);
nor U8700 (N_8700,N_8672,N_8619);
nor U8701 (N_8701,N_8694,N_8628);
nor U8702 (N_8702,N_8604,N_8644);
xor U8703 (N_8703,N_8654,N_8651);
nand U8704 (N_8704,N_8617,N_8647);
nand U8705 (N_8705,N_8699,N_8693);
nor U8706 (N_8706,N_8675,N_8678);
nor U8707 (N_8707,N_8603,N_8660);
or U8708 (N_8708,N_8600,N_8618);
or U8709 (N_8709,N_8645,N_8670);
xnor U8710 (N_8710,N_8643,N_8697);
nor U8711 (N_8711,N_8659,N_8632);
xor U8712 (N_8712,N_8641,N_8629);
or U8713 (N_8713,N_8634,N_8689);
and U8714 (N_8714,N_8614,N_8625);
and U8715 (N_8715,N_8658,N_8686);
nand U8716 (N_8716,N_8695,N_8633);
or U8717 (N_8717,N_8650,N_8674);
nor U8718 (N_8718,N_8676,N_8683);
nor U8719 (N_8719,N_8649,N_8665);
and U8720 (N_8720,N_8606,N_8640);
and U8721 (N_8721,N_8685,N_8622);
xnor U8722 (N_8722,N_8691,N_8682);
and U8723 (N_8723,N_8624,N_8601);
nand U8724 (N_8724,N_8637,N_8671);
and U8725 (N_8725,N_8679,N_8636);
and U8726 (N_8726,N_8620,N_8609);
nand U8727 (N_8727,N_8661,N_8669);
xor U8728 (N_8728,N_8653,N_8698);
nor U8729 (N_8729,N_8687,N_8616);
nand U8730 (N_8730,N_8613,N_8673);
nand U8731 (N_8731,N_8615,N_8608);
nor U8732 (N_8732,N_8692,N_8623);
and U8733 (N_8733,N_8655,N_8602);
and U8734 (N_8734,N_8662,N_8656);
and U8735 (N_8735,N_8681,N_8667);
nor U8736 (N_8736,N_8652,N_8680);
nand U8737 (N_8737,N_8638,N_8648);
or U8738 (N_8738,N_8611,N_8612);
or U8739 (N_8739,N_8664,N_8677);
nor U8740 (N_8740,N_8688,N_8646);
nor U8741 (N_8741,N_8639,N_8657);
nor U8742 (N_8742,N_8684,N_8696);
nand U8743 (N_8743,N_8663,N_8626);
and U8744 (N_8744,N_8627,N_8607);
or U8745 (N_8745,N_8690,N_8631);
xor U8746 (N_8746,N_8621,N_8668);
or U8747 (N_8747,N_8666,N_8610);
xnor U8748 (N_8748,N_8642,N_8635);
and U8749 (N_8749,N_8605,N_8630);
and U8750 (N_8750,N_8651,N_8673);
nor U8751 (N_8751,N_8634,N_8696);
nor U8752 (N_8752,N_8651,N_8694);
xor U8753 (N_8753,N_8634,N_8632);
nand U8754 (N_8754,N_8688,N_8627);
or U8755 (N_8755,N_8609,N_8647);
and U8756 (N_8756,N_8607,N_8699);
nor U8757 (N_8757,N_8667,N_8614);
or U8758 (N_8758,N_8653,N_8666);
and U8759 (N_8759,N_8635,N_8649);
nand U8760 (N_8760,N_8601,N_8689);
or U8761 (N_8761,N_8697,N_8607);
nand U8762 (N_8762,N_8693,N_8634);
and U8763 (N_8763,N_8643,N_8650);
xor U8764 (N_8764,N_8608,N_8686);
nand U8765 (N_8765,N_8680,N_8666);
or U8766 (N_8766,N_8621,N_8611);
or U8767 (N_8767,N_8660,N_8651);
xor U8768 (N_8768,N_8634,N_8681);
xor U8769 (N_8769,N_8682,N_8657);
or U8770 (N_8770,N_8618,N_8655);
nand U8771 (N_8771,N_8653,N_8640);
nand U8772 (N_8772,N_8666,N_8641);
or U8773 (N_8773,N_8610,N_8662);
and U8774 (N_8774,N_8697,N_8678);
xnor U8775 (N_8775,N_8667,N_8689);
nand U8776 (N_8776,N_8607,N_8655);
nand U8777 (N_8777,N_8620,N_8678);
nand U8778 (N_8778,N_8602,N_8657);
or U8779 (N_8779,N_8697,N_8621);
nor U8780 (N_8780,N_8676,N_8688);
nor U8781 (N_8781,N_8627,N_8601);
and U8782 (N_8782,N_8633,N_8654);
nor U8783 (N_8783,N_8685,N_8606);
nor U8784 (N_8784,N_8674,N_8602);
nor U8785 (N_8785,N_8688,N_8612);
and U8786 (N_8786,N_8646,N_8680);
nand U8787 (N_8787,N_8633,N_8661);
nand U8788 (N_8788,N_8631,N_8653);
and U8789 (N_8789,N_8678,N_8640);
nor U8790 (N_8790,N_8639,N_8663);
and U8791 (N_8791,N_8661,N_8684);
nand U8792 (N_8792,N_8695,N_8674);
or U8793 (N_8793,N_8682,N_8606);
or U8794 (N_8794,N_8661,N_8608);
nor U8795 (N_8795,N_8676,N_8669);
or U8796 (N_8796,N_8625,N_8673);
nand U8797 (N_8797,N_8680,N_8617);
xor U8798 (N_8798,N_8602,N_8656);
nor U8799 (N_8799,N_8663,N_8675);
or U8800 (N_8800,N_8789,N_8745);
or U8801 (N_8801,N_8711,N_8758);
and U8802 (N_8802,N_8722,N_8768);
nor U8803 (N_8803,N_8739,N_8772);
xor U8804 (N_8804,N_8788,N_8792);
and U8805 (N_8805,N_8767,N_8703);
or U8806 (N_8806,N_8754,N_8763);
nor U8807 (N_8807,N_8764,N_8798);
xor U8808 (N_8808,N_8736,N_8738);
nand U8809 (N_8809,N_8720,N_8734);
nor U8810 (N_8810,N_8756,N_8706);
nor U8811 (N_8811,N_8721,N_8718);
and U8812 (N_8812,N_8760,N_8775);
xnor U8813 (N_8813,N_8723,N_8704);
nand U8814 (N_8814,N_8705,N_8707);
nor U8815 (N_8815,N_8786,N_8782);
nor U8816 (N_8816,N_8799,N_8759);
and U8817 (N_8817,N_8735,N_8748);
and U8818 (N_8818,N_8794,N_8791);
nor U8819 (N_8819,N_8765,N_8777);
or U8820 (N_8820,N_8742,N_8787);
nand U8821 (N_8821,N_8769,N_8749);
or U8822 (N_8822,N_8713,N_8773);
or U8823 (N_8823,N_8709,N_8761);
nor U8824 (N_8824,N_8728,N_8732);
or U8825 (N_8825,N_8755,N_8702);
xor U8826 (N_8826,N_8757,N_8778);
or U8827 (N_8827,N_8744,N_8710);
or U8828 (N_8828,N_8746,N_8724);
xnor U8829 (N_8829,N_8795,N_8725);
nor U8830 (N_8830,N_8700,N_8740);
or U8831 (N_8831,N_8715,N_8784);
xor U8832 (N_8832,N_8774,N_8779);
xor U8833 (N_8833,N_8733,N_8750);
or U8834 (N_8834,N_8727,N_8770);
nor U8835 (N_8835,N_8726,N_8701);
nand U8836 (N_8836,N_8796,N_8708);
xor U8837 (N_8837,N_8762,N_8785);
xor U8838 (N_8838,N_8719,N_8716);
xor U8839 (N_8839,N_8766,N_8712);
and U8840 (N_8840,N_8753,N_8714);
nor U8841 (N_8841,N_8781,N_8717);
nor U8842 (N_8842,N_8793,N_8730);
xnor U8843 (N_8843,N_8776,N_8783);
nor U8844 (N_8844,N_8752,N_8729);
or U8845 (N_8845,N_8737,N_8790);
nor U8846 (N_8846,N_8743,N_8741);
or U8847 (N_8847,N_8780,N_8747);
or U8848 (N_8848,N_8731,N_8751);
nand U8849 (N_8849,N_8797,N_8771);
nand U8850 (N_8850,N_8772,N_8780);
xor U8851 (N_8851,N_8748,N_8747);
nand U8852 (N_8852,N_8786,N_8727);
xnor U8853 (N_8853,N_8748,N_8764);
or U8854 (N_8854,N_8724,N_8716);
and U8855 (N_8855,N_8759,N_8710);
xor U8856 (N_8856,N_8751,N_8763);
nor U8857 (N_8857,N_8727,N_8780);
xnor U8858 (N_8858,N_8773,N_8737);
and U8859 (N_8859,N_8768,N_8774);
nor U8860 (N_8860,N_8795,N_8757);
xor U8861 (N_8861,N_8793,N_8716);
nor U8862 (N_8862,N_8726,N_8750);
nor U8863 (N_8863,N_8795,N_8750);
xor U8864 (N_8864,N_8765,N_8720);
nand U8865 (N_8865,N_8739,N_8712);
xnor U8866 (N_8866,N_8757,N_8721);
and U8867 (N_8867,N_8775,N_8732);
or U8868 (N_8868,N_8705,N_8768);
xor U8869 (N_8869,N_8776,N_8761);
nor U8870 (N_8870,N_8742,N_8728);
or U8871 (N_8871,N_8729,N_8767);
and U8872 (N_8872,N_8745,N_8727);
nor U8873 (N_8873,N_8794,N_8726);
or U8874 (N_8874,N_8734,N_8724);
and U8875 (N_8875,N_8779,N_8777);
and U8876 (N_8876,N_8702,N_8756);
nor U8877 (N_8877,N_8776,N_8765);
nand U8878 (N_8878,N_8741,N_8769);
nand U8879 (N_8879,N_8798,N_8793);
or U8880 (N_8880,N_8752,N_8707);
xnor U8881 (N_8881,N_8771,N_8776);
xor U8882 (N_8882,N_8771,N_8785);
nor U8883 (N_8883,N_8742,N_8775);
xor U8884 (N_8884,N_8757,N_8708);
or U8885 (N_8885,N_8738,N_8715);
nand U8886 (N_8886,N_8779,N_8771);
and U8887 (N_8887,N_8734,N_8745);
or U8888 (N_8888,N_8774,N_8782);
nor U8889 (N_8889,N_8719,N_8786);
nor U8890 (N_8890,N_8721,N_8720);
nand U8891 (N_8891,N_8704,N_8769);
and U8892 (N_8892,N_8743,N_8725);
and U8893 (N_8893,N_8710,N_8706);
or U8894 (N_8894,N_8748,N_8716);
nand U8895 (N_8895,N_8758,N_8704);
xor U8896 (N_8896,N_8791,N_8708);
or U8897 (N_8897,N_8710,N_8727);
xor U8898 (N_8898,N_8709,N_8731);
and U8899 (N_8899,N_8775,N_8771);
nor U8900 (N_8900,N_8806,N_8847);
or U8901 (N_8901,N_8800,N_8879);
or U8902 (N_8902,N_8880,N_8858);
xor U8903 (N_8903,N_8885,N_8822);
nor U8904 (N_8904,N_8894,N_8860);
and U8905 (N_8905,N_8876,N_8813);
nor U8906 (N_8906,N_8842,N_8841);
and U8907 (N_8907,N_8898,N_8854);
and U8908 (N_8908,N_8846,N_8896);
and U8909 (N_8909,N_8891,N_8801);
xnor U8910 (N_8910,N_8888,N_8838);
nor U8911 (N_8911,N_8877,N_8866);
nor U8912 (N_8912,N_8844,N_8850);
or U8913 (N_8913,N_8829,N_8881);
and U8914 (N_8914,N_8849,N_8859);
and U8915 (N_8915,N_8889,N_8864);
xor U8916 (N_8916,N_8819,N_8886);
or U8917 (N_8917,N_8878,N_8816);
nor U8918 (N_8918,N_8834,N_8865);
nor U8919 (N_8919,N_8855,N_8828);
and U8920 (N_8920,N_8852,N_8871);
and U8921 (N_8921,N_8812,N_8874);
or U8922 (N_8922,N_8868,N_8804);
or U8923 (N_8923,N_8805,N_8815);
nor U8924 (N_8924,N_8811,N_8820);
xnor U8925 (N_8925,N_8861,N_8848);
nor U8926 (N_8926,N_8863,N_8883);
and U8927 (N_8927,N_8824,N_8867);
or U8928 (N_8928,N_8839,N_8899);
nand U8929 (N_8929,N_8807,N_8826);
nor U8930 (N_8930,N_8856,N_8818);
nand U8931 (N_8931,N_8872,N_8830);
or U8932 (N_8932,N_8897,N_8895);
or U8933 (N_8933,N_8809,N_8832);
nand U8934 (N_8934,N_8831,N_8851);
and U8935 (N_8935,N_8823,N_8827);
xor U8936 (N_8936,N_8873,N_8833);
nand U8937 (N_8937,N_8810,N_8887);
nand U8938 (N_8938,N_8884,N_8843);
and U8939 (N_8939,N_8836,N_8837);
nor U8940 (N_8940,N_8853,N_8808);
xor U8941 (N_8941,N_8835,N_8893);
xnor U8942 (N_8942,N_8862,N_8817);
and U8943 (N_8943,N_8840,N_8845);
and U8944 (N_8944,N_8857,N_8869);
nand U8945 (N_8945,N_8892,N_8882);
nor U8946 (N_8946,N_8803,N_8875);
nor U8947 (N_8947,N_8814,N_8890);
nand U8948 (N_8948,N_8825,N_8802);
and U8949 (N_8949,N_8870,N_8821);
nand U8950 (N_8950,N_8856,N_8855);
or U8951 (N_8951,N_8843,N_8891);
nor U8952 (N_8952,N_8899,N_8835);
xnor U8953 (N_8953,N_8855,N_8811);
nand U8954 (N_8954,N_8850,N_8895);
nor U8955 (N_8955,N_8837,N_8822);
xor U8956 (N_8956,N_8825,N_8866);
or U8957 (N_8957,N_8898,N_8803);
nand U8958 (N_8958,N_8822,N_8832);
xnor U8959 (N_8959,N_8883,N_8838);
xnor U8960 (N_8960,N_8803,N_8830);
and U8961 (N_8961,N_8821,N_8882);
nand U8962 (N_8962,N_8808,N_8880);
or U8963 (N_8963,N_8819,N_8854);
and U8964 (N_8964,N_8823,N_8893);
and U8965 (N_8965,N_8839,N_8819);
nor U8966 (N_8966,N_8841,N_8827);
nor U8967 (N_8967,N_8893,N_8870);
and U8968 (N_8968,N_8851,N_8894);
or U8969 (N_8969,N_8826,N_8859);
xnor U8970 (N_8970,N_8870,N_8833);
and U8971 (N_8971,N_8878,N_8825);
or U8972 (N_8972,N_8867,N_8842);
nand U8973 (N_8973,N_8862,N_8890);
and U8974 (N_8974,N_8816,N_8835);
xor U8975 (N_8975,N_8892,N_8845);
nor U8976 (N_8976,N_8868,N_8824);
xor U8977 (N_8977,N_8846,N_8898);
and U8978 (N_8978,N_8870,N_8881);
xor U8979 (N_8979,N_8831,N_8806);
or U8980 (N_8980,N_8821,N_8867);
nand U8981 (N_8981,N_8813,N_8870);
nand U8982 (N_8982,N_8820,N_8803);
or U8983 (N_8983,N_8880,N_8847);
nor U8984 (N_8984,N_8860,N_8826);
xor U8985 (N_8985,N_8830,N_8801);
nand U8986 (N_8986,N_8858,N_8866);
nand U8987 (N_8987,N_8833,N_8882);
or U8988 (N_8988,N_8875,N_8847);
nor U8989 (N_8989,N_8822,N_8896);
nand U8990 (N_8990,N_8864,N_8845);
and U8991 (N_8991,N_8857,N_8899);
and U8992 (N_8992,N_8805,N_8854);
nand U8993 (N_8993,N_8812,N_8884);
or U8994 (N_8994,N_8879,N_8807);
or U8995 (N_8995,N_8867,N_8859);
nor U8996 (N_8996,N_8876,N_8812);
or U8997 (N_8997,N_8831,N_8821);
or U8998 (N_8998,N_8885,N_8855);
nand U8999 (N_8999,N_8811,N_8835);
nor U9000 (N_9000,N_8935,N_8982);
xor U9001 (N_9001,N_8956,N_8963);
nor U9002 (N_9002,N_8954,N_8937);
nor U9003 (N_9003,N_8911,N_8941);
nand U9004 (N_9004,N_8989,N_8928);
or U9005 (N_9005,N_8903,N_8991);
xnor U9006 (N_9006,N_8957,N_8907);
and U9007 (N_9007,N_8917,N_8925);
or U9008 (N_9008,N_8908,N_8923);
or U9009 (N_9009,N_8944,N_8951);
and U9010 (N_9010,N_8999,N_8993);
xnor U9011 (N_9011,N_8942,N_8924);
or U9012 (N_9012,N_8926,N_8998);
or U9013 (N_9013,N_8965,N_8930);
nor U9014 (N_9014,N_8940,N_8969);
xnor U9015 (N_9015,N_8945,N_8988);
nor U9016 (N_9016,N_8984,N_8946);
nand U9017 (N_9017,N_8948,N_8915);
xor U9018 (N_9018,N_8986,N_8977);
xnor U9019 (N_9019,N_8916,N_8976);
nand U9020 (N_9020,N_8905,N_8978);
nand U9021 (N_9021,N_8901,N_8960);
or U9022 (N_9022,N_8961,N_8932);
and U9023 (N_9023,N_8934,N_8918);
nand U9024 (N_9024,N_8971,N_8962);
xnor U9025 (N_9025,N_8992,N_8938);
and U9026 (N_9026,N_8975,N_8952);
or U9027 (N_9027,N_8912,N_8981);
and U9028 (N_9028,N_8931,N_8933);
and U9029 (N_9029,N_8990,N_8955);
or U9030 (N_9030,N_8922,N_8979);
and U9031 (N_9031,N_8966,N_8939);
xnor U9032 (N_9032,N_8913,N_8983);
and U9033 (N_9033,N_8921,N_8972);
nand U9034 (N_9034,N_8964,N_8953);
or U9035 (N_9035,N_8994,N_8949);
or U9036 (N_9036,N_8995,N_8919);
or U9037 (N_9037,N_8950,N_8959);
or U9038 (N_9038,N_8947,N_8904);
and U9039 (N_9039,N_8996,N_8958);
and U9040 (N_9040,N_8920,N_8985);
or U9041 (N_9041,N_8906,N_8980);
nor U9042 (N_9042,N_8968,N_8910);
nand U9043 (N_9043,N_8967,N_8943);
and U9044 (N_9044,N_8909,N_8974);
nand U9045 (N_9045,N_8987,N_8902);
xnor U9046 (N_9046,N_8927,N_8929);
or U9047 (N_9047,N_8900,N_8914);
nor U9048 (N_9048,N_8936,N_8970);
nor U9049 (N_9049,N_8973,N_8997);
and U9050 (N_9050,N_8908,N_8924);
nand U9051 (N_9051,N_8989,N_8932);
and U9052 (N_9052,N_8977,N_8975);
and U9053 (N_9053,N_8941,N_8962);
and U9054 (N_9054,N_8966,N_8974);
and U9055 (N_9055,N_8955,N_8945);
nor U9056 (N_9056,N_8953,N_8997);
xnor U9057 (N_9057,N_8966,N_8999);
nand U9058 (N_9058,N_8993,N_8981);
nand U9059 (N_9059,N_8981,N_8982);
nand U9060 (N_9060,N_8961,N_8942);
and U9061 (N_9061,N_8961,N_8982);
nand U9062 (N_9062,N_8939,N_8962);
nand U9063 (N_9063,N_8969,N_8900);
xor U9064 (N_9064,N_8904,N_8966);
nor U9065 (N_9065,N_8931,N_8963);
xnor U9066 (N_9066,N_8932,N_8931);
xor U9067 (N_9067,N_8919,N_8951);
nor U9068 (N_9068,N_8986,N_8947);
xnor U9069 (N_9069,N_8924,N_8904);
and U9070 (N_9070,N_8970,N_8966);
nor U9071 (N_9071,N_8948,N_8990);
or U9072 (N_9072,N_8916,N_8986);
and U9073 (N_9073,N_8989,N_8906);
or U9074 (N_9074,N_8966,N_8996);
nor U9075 (N_9075,N_8970,N_8997);
xnor U9076 (N_9076,N_8972,N_8958);
nor U9077 (N_9077,N_8991,N_8984);
xnor U9078 (N_9078,N_8948,N_8937);
nand U9079 (N_9079,N_8979,N_8912);
nor U9080 (N_9080,N_8942,N_8932);
nand U9081 (N_9081,N_8988,N_8989);
or U9082 (N_9082,N_8906,N_8962);
xnor U9083 (N_9083,N_8968,N_8928);
and U9084 (N_9084,N_8971,N_8969);
and U9085 (N_9085,N_8910,N_8941);
nand U9086 (N_9086,N_8975,N_8915);
xnor U9087 (N_9087,N_8922,N_8907);
xnor U9088 (N_9088,N_8994,N_8903);
xor U9089 (N_9089,N_8939,N_8992);
and U9090 (N_9090,N_8955,N_8922);
xor U9091 (N_9091,N_8934,N_8971);
nor U9092 (N_9092,N_8988,N_8973);
xor U9093 (N_9093,N_8935,N_8908);
nor U9094 (N_9094,N_8978,N_8943);
or U9095 (N_9095,N_8976,N_8993);
nor U9096 (N_9096,N_8956,N_8968);
nand U9097 (N_9097,N_8959,N_8923);
nor U9098 (N_9098,N_8901,N_8967);
and U9099 (N_9099,N_8993,N_8987);
nor U9100 (N_9100,N_9066,N_9029);
xor U9101 (N_9101,N_9032,N_9056);
nand U9102 (N_9102,N_9092,N_9033);
nand U9103 (N_9103,N_9099,N_9084);
or U9104 (N_9104,N_9011,N_9000);
nor U9105 (N_9105,N_9040,N_9002);
and U9106 (N_9106,N_9052,N_9037);
and U9107 (N_9107,N_9085,N_9076);
nand U9108 (N_9108,N_9096,N_9058);
and U9109 (N_9109,N_9068,N_9048);
or U9110 (N_9110,N_9057,N_9006);
nand U9111 (N_9111,N_9051,N_9072);
nor U9112 (N_9112,N_9042,N_9007);
or U9113 (N_9113,N_9045,N_9049);
nand U9114 (N_9114,N_9064,N_9091);
nor U9115 (N_9115,N_9044,N_9025);
or U9116 (N_9116,N_9038,N_9019);
or U9117 (N_9117,N_9009,N_9089);
nand U9118 (N_9118,N_9024,N_9003);
and U9119 (N_9119,N_9078,N_9086);
xor U9120 (N_9120,N_9021,N_9039);
nor U9121 (N_9121,N_9030,N_9081);
nand U9122 (N_9122,N_9035,N_9055);
xor U9123 (N_9123,N_9015,N_9034);
nand U9124 (N_9124,N_9073,N_9074);
nand U9125 (N_9125,N_9079,N_9001);
nand U9126 (N_9126,N_9046,N_9062);
and U9127 (N_9127,N_9077,N_9054);
nor U9128 (N_9128,N_9083,N_9065);
and U9129 (N_9129,N_9080,N_9090);
xnor U9130 (N_9130,N_9036,N_9008);
or U9131 (N_9131,N_9004,N_9012);
and U9132 (N_9132,N_9071,N_9047);
or U9133 (N_9133,N_9050,N_9005);
xnor U9134 (N_9134,N_9060,N_9059);
nor U9135 (N_9135,N_9026,N_9067);
or U9136 (N_9136,N_9016,N_9022);
nand U9137 (N_9137,N_9069,N_9010);
nor U9138 (N_9138,N_9095,N_9087);
or U9139 (N_9139,N_9020,N_9094);
nand U9140 (N_9140,N_9031,N_9043);
xor U9141 (N_9141,N_9070,N_9014);
xor U9142 (N_9142,N_9063,N_9053);
nand U9143 (N_9143,N_9088,N_9027);
and U9144 (N_9144,N_9023,N_9098);
nand U9145 (N_9145,N_9082,N_9013);
nor U9146 (N_9146,N_9093,N_9028);
or U9147 (N_9147,N_9017,N_9097);
and U9148 (N_9148,N_9018,N_9075);
nand U9149 (N_9149,N_9041,N_9061);
nand U9150 (N_9150,N_9092,N_9007);
and U9151 (N_9151,N_9091,N_9066);
or U9152 (N_9152,N_9013,N_9056);
or U9153 (N_9153,N_9032,N_9089);
nor U9154 (N_9154,N_9021,N_9030);
or U9155 (N_9155,N_9022,N_9058);
xnor U9156 (N_9156,N_9082,N_9025);
and U9157 (N_9157,N_9013,N_9022);
xnor U9158 (N_9158,N_9072,N_9021);
nand U9159 (N_9159,N_9088,N_9018);
or U9160 (N_9160,N_9098,N_9003);
and U9161 (N_9161,N_9058,N_9079);
or U9162 (N_9162,N_9027,N_9096);
or U9163 (N_9163,N_9082,N_9026);
or U9164 (N_9164,N_9088,N_9037);
and U9165 (N_9165,N_9018,N_9028);
nand U9166 (N_9166,N_9085,N_9042);
xor U9167 (N_9167,N_9038,N_9043);
or U9168 (N_9168,N_9099,N_9087);
or U9169 (N_9169,N_9076,N_9053);
nand U9170 (N_9170,N_9093,N_9078);
nor U9171 (N_9171,N_9095,N_9073);
and U9172 (N_9172,N_9053,N_9002);
or U9173 (N_9173,N_9083,N_9078);
nor U9174 (N_9174,N_9030,N_9090);
or U9175 (N_9175,N_9043,N_9089);
and U9176 (N_9176,N_9098,N_9041);
or U9177 (N_9177,N_9040,N_9029);
nand U9178 (N_9178,N_9058,N_9004);
nor U9179 (N_9179,N_9067,N_9062);
nand U9180 (N_9180,N_9002,N_9057);
nand U9181 (N_9181,N_9073,N_9008);
xnor U9182 (N_9182,N_9037,N_9057);
xnor U9183 (N_9183,N_9096,N_9045);
nor U9184 (N_9184,N_9021,N_9087);
nor U9185 (N_9185,N_9093,N_9018);
or U9186 (N_9186,N_9044,N_9007);
xor U9187 (N_9187,N_9059,N_9039);
and U9188 (N_9188,N_9052,N_9007);
nor U9189 (N_9189,N_9030,N_9077);
nor U9190 (N_9190,N_9019,N_9013);
nand U9191 (N_9191,N_9051,N_9059);
and U9192 (N_9192,N_9014,N_9028);
and U9193 (N_9193,N_9068,N_9089);
or U9194 (N_9194,N_9026,N_9088);
xor U9195 (N_9195,N_9026,N_9095);
or U9196 (N_9196,N_9040,N_9071);
or U9197 (N_9197,N_9039,N_9072);
xnor U9198 (N_9198,N_9086,N_9051);
xor U9199 (N_9199,N_9098,N_9020);
nand U9200 (N_9200,N_9182,N_9151);
or U9201 (N_9201,N_9159,N_9127);
and U9202 (N_9202,N_9187,N_9105);
nand U9203 (N_9203,N_9146,N_9108);
nor U9204 (N_9204,N_9168,N_9130);
nand U9205 (N_9205,N_9158,N_9157);
and U9206 (N_9206,N_9116,N_9142);
xor U9207 (N_9207,N_9125,N_9144);
xnor U9208 (N_9208,N_9135,N_9185);
and U9209 (N_9209,N_9112,N_9141);
nor U9210 (N_9210,N_9198,N_9106);
nand U9211 (N_9211,N_9174,N_9179);
or U9212 (N_9212,N_9194,N_9124);
or U9213 (N_9213,N_9152,N_9166);
nor U9214 (N_9214,N_9181,N_9196);
xnor U9215 (N_9215,N_9119,N_9155);
or U9216 (N_9216,N_9126,N_9128);
nand U9217 (N_9217,N_9115,N_9122);
and U9218 (N_9218,N_9114,N_9117);
nand U9219 (N_9219,N_9191,N_9193);
and U9220 (N_9220,N_9180,N_9154);
and U9221 (N_9221,N_9192,N_9165);
and U9222 (N_9222,N_9173,N_9118);
xor U9223 (N_9223,N_9149,N_9175);
nor U9224 (N_9224,N_9199,N_9123);
nand U9225 (N_9225,N_9186,N_9147);
nand U9226 (N_9226,N_9183,N_9101);
or U9227 (N_9227,N_9163,N_9120);
xnor U9228 (N_9228,N_9190,N_9121);
xor U9229 (N_9229,N_9104,N_9138);
xor U9230 (N_9230,N_9164,N_9100);
nor U9231 (N_9231,N_9134,N_9169);
nand U9232 (N_9232,N_9103,N_9167);
and U9233 (N_9233,N_9189,N_9113);
or U9234 (N_9234,N_9129,N_9156);
nand U9235 (N_9235,N_9195,N_9188);
xnor U9236 (N_9236,N_9133,N_9150);
or U9237 (N_9237,N_9148,N_9153);
nor U9238 (N_9238,N_9140,N_9111);
and U9239 (N_9239,N_9160,N_9136);
xor U9240 (N_9240,N_9145,N_9177);
and U9241 (N_9241,N_9176,N_9161);
nor U9242 (N_9242,N_9171,N_9139);
nand U9243 (N_9243,N_9143,N_9109);
nand U9244 (N_9244,N_9110,N_9131);
xnor U9245 (N_9245,N_9170,N_9162);
or U9246 (N_9246,N_9184,N_9132);
nand U9247 (N_9247,N_9137,N_9178);
and U9248 (N_9248,N_9107,N_9172);
and U9249 (N_9249,N_9102,N_9197);
xor U9250 (N_9250,N_9159,N_9129);
and U9251 (N_9251,N_9116,N_9185);
xnor U9252 (N_9252,N_9191,N_9141);
nor U9253 (N_9253,N_9151,N_9113);
nor U9254 (N_9254,N_9106,N_9150);
nand U9255 (N_9255,N_9115,N_9104);
or U9256 (N_9256,N_9168,N_9166);
or U9257 (N_9257,N_9112,N_9184);
and U9258 (N_9258,N_9125,N_9192);
nand U9259 (N_9259,N_9196,N_9101);
and U9260 (N_9260,N_9172,N_9193);
or U9261 (N_9261,N_9122,N_9119);
or U9262 (N_9262,N_9183,N_9113);
and U9263 (N_9263,N_9188,N_9131);
and U9264 (N_9264,N_9105,N_9175);
nand U9265 (N_9265,N_9167,N_9141);
nor U9266 (N_9266,N_9169,N_9127);
nor U9267 (N_9267,N_9140,N_9182);
or U9268 (N_9268,N_9105,N_9149);
nand U9269 (N_9269,N_9143,N_9142);
nand U9270 (N_9270,N_9117,N_9147);
nand U9271 (N_9271,N_9196,N_9111);
xnor U9272 (N_9272,N_9139,N_9137);
and U9273 (N_9273,N_9135,N_9158);
xnor U9274 (N_9274,N_9130,N_9132);
or U9275 (N_9275,N_9105,N_9182);
nand U9276 (N_9276,N_9171,N_9156);
and U9277 (N_9277,N_9183,N_9111);
xnor U9278 (N_9278,N_9118,N_9190);
nand U9279 (N_9279,N_9163,N_9197);
nand U9280 (N_9280,N_9107,N_9195);
nand U9281 (N_9281,N_9131,N_9145);
or U9282 (N_9282,N_9139,N_9125);
xor U9283 (N_9283,N_9177,N_9193);
nor U9284 (N_9284,N_9105,N_9120);
or U9285 (N_9285,N_9199,N_9120);
nor U9286 (N_9286,N_9135,N_9114);
or U9287 (N_9287,N_9124,N_9115);
xnor U9288 (N_9288,N_9174,N_9148);
nor U9289 (N_9289,N_9139,N_9195);
xnor U9290 (N_9290,N_9190,N_9138);
nor U9291 (N_9291,N_9190,N_9142);
nor U9292 (N_9292,N_9125,N_9162);
nand U9293 (N_9293,N_9155,N_9121);
and U9294 (N_9294,N_9145,N_9159);
nand U9295 (N_9295,N_9179,N_9125);
or U9296 (N_9296,N_9171,N_9148);
nand U9297 (N_9297,N_9198,N_9151);
and U9298 (N_9298,N_9178,N_9175);
or U9299 (N_9299,N_9170,N_9110);
nor U9300 (N_9300,N_9219,N_9292);
xor U9301 (N_9301,N_9223,N_9285);
nand U9302 (N_9302,N_9245,N_9224);
xor U9303 (N_9303,N_9288,N_9216);
or U9304 (N_9304,N_9242,N_9297);
nand U9305 (N_9305,N_9240,N_9262);
xor U9306 (N_9306,N_9210,N_9284);
xnor U9307 (N_9307,N_9296,N_9215);
or U9308 (N_9308,N_9264,N_9295);
nand U9309 (N_9309,N_9269,N_9253);
and U9310 (N_9310,N_9291,N_9230);
nor U9311 (N_9311,N_9212,N_9254);
xor U9312 (N_9312,N_9247,N_9246);
xnor U9313 (N_9313,N_9244,N_9208);
nor U9314 (N_9314,N_9290,N_9252);
or U9315 (N_9315,N_9275,N_9221);
nor U9316 (N_9316,N_9237,N_9255);
nor U9317 (N_9317,N_9299,N_9203);
nand U9318 (N_9318,N_9217,N_9226);
nor U9319 (N_9319,N_9206,N_9232);
and U9320 (N_9320,N_9241,N_9248);
nor U9321 (N_9321,N_9233,N_9222);
nor U9322 (N_9322,N_9276,N_9213);
or U9323 (N_9323,N_9205,N_9286);
xnor U9324 (N_9324,N_9257,N_9228);
and U9325 (N_9325,N_9293,N_9298);
xor U9326 (N_9326,N_9214,N_9229);
nor U9327 (N_9327,N_9268,N_9218);
xor U9328 (N_9328,N_9243,N_9207);
xor U9329 (N_9329,N_9270,N_9271);
or U9330 (N_9330,N_9235,N_9267);
or U9331 (N_9331,N_9220,N_9266);
xnor U9332 (N_9332,N_9258,N_9260);
xnor U9333 (N_9333,N_9227,N_9225);
and U9334 (N_9334,N_9277,N_9287);
nand U9335 (N_9335,N_9294,N_9280);
nor U9336 (N_9336,N_9289,N_9200);
xnor U9337 (N_9337,N_9234,N_9281);
and U9338 (N_9338,N_9272,N_9256);
xor U9339 (N_9339,N_9202,N_9259);
nor U9340 (N_9340,N_9249,N_9211);
xor U9341 (N_9341,N_9251,N_9209);
nand U9342 (N_9342,N_9250,N_9283);
xor U9343 (N_9343,N_9273,N_9265);
xnor U9344 (N_9344,N_9238,N_9278);
and U9345 (N_9345,N_9279,N_9261);
nand U9346 (N_9346,N_9263,N_9274);
nor U9347 (N_9347,N_9236,N_9204);
nand U9348 (N_9348,N_9282,N_9231);
xnor U9349 (N_9349,N_9239,N_9201);
nand U9350 (N_9350,N_9232,N_9224);
nand U9351 (N_9351,N_9210,N_9270);
and U9352 (N_9352,N_9202,N_9279);
xnor U9353 (N_9353,N_9295,N_9268);
xnor U9354 (N_9354,N_9284,N_9235);
nand U9355 (N_9355,N_9215,N_9207);
or U9356 (N_9356,N_9220,N_9274);
and U9357 (N_9357,N_9219,N_9284);
nor U9358 (N_9358,N_9264,N_9235);
and U9359 (N_9359,N_9213,N_9255);
nand U9360 (N_9360,N_9216,N_9207);
nor U9361 (N_9361,N_9247,N_9271);
or U9362 (N_9362,N_9243,N_9234);
and U9363 (N_9363,N_9216,N_9225);
nand U9364 (N_9364,N_9282,N_9221);
nor U9365 (N_9365,N_9296,N_9295);
or U9366 (N_9366,N_9281,N_9254);
nand U9367 (N_9367,N_9267,N_9250);
and U9368 (N_9368,N_9240,N_9244);
or U9369 (N_9369,N_9234,N_9236);
or U9370 (N_9370,N_9276,N_9284);
or U9371 (N_9371,N_9238,N_9232);
nand U9372 (N_9372,N_9260,N_9285);
or U9373 (N_9373,N_9263,N_9214);
xnor U9374 (N_9374,N_9224,N_9273);
xnor U9375 (N_9375,N_9246,N_9280);
nor U9376 (N_9376,N_9251,N_9200);
nand U9377 (N_9377,N_9261,N_9201);
or U9378 (N_9378,N_9224,N_9283);
and U9379 (N_9379,N_9292,N_9232);
nor U9380 (N_9380,N_9218,N_9293);
nor U9381 (N_9381,N_9228,N_9243);
nor U9382 (N_9382,N_9290,N_9248);
nor U9383 (N_9383,N_9265,N_9248);
nand U9384 (N_9384,N_9290,N_9233);
nor U9385 (N_9385,N_9240,N_9206);
nand U9386 (N_9386,N_9253,N_9264);
and U9387 (N_9387,N_9284,N_9273);
nand U9388 (N_9388,N_9277,N_9208);
and U9389 (N_9389,N_9277,N_9221);
nand U9390 (N_9390,N_9296,N_9272);
xor U9391 (N_9391,N_9234,N_9245);
or U9392 (N_9392,N_9243,N_9299);
and U9393 (N_9393,N_9248,N_9282);
nor U9394 (N_9394,N_9247,N_9261);
xor U9395 (N_9395,N_9261,N_9204);
and U9396 (N_9396,N_9211,N_9298);
and U9397 (N_9397,N_9244,N_9292);
and U9398 (N_9398,N_9251,N_9208);
and U9399 (N_9399,N_9255,N_9287);
nor U9400 (N_9400,N_9399,N_9381);
or U9401 (N_9401,N_9324,N_9375);
xor U9402 (N_9402,N_9367,N_9387);
nand U9403 (N_9403,N_9357,N_9341);
nor U9404 (N_9404,N_9388,N_9345);
nand U9405 (N_9405,N_9316,N_9333);
and U9406 (N_9406,N_9360,N_9302);
or U9407 (N_9407,N_9348,N_9398);
nand U9408 (N_9408,N_9350,N_9376);
nand U9409 (N_9409,N_9374,N_9311);
or U9410 (N_9410,N_9339,N_9300);
nand U9411 (N_9411,N_9319,N_9330);
nand U9412 (N_9412,N_9327,N_9310);
and U9413 (N_9413,N_9328,N_9305);
and U9414 (N_9414,N_9307,N_9340);
xnor U9415 (N_9415,N_9347,N_9373);
or U9416 (N_9416,N_9346,N_9335);
nor U9417 (N_9417,N_9336,N_9383);
nor U9418 (N_9418,N_9308,N_9384);
or U9419 (N_9419,N_9358,N_9363);
and U9420 (N_9420,N_9366,N_9362);
or U9421 (N_9421,N_9304,N_9355);
nor U9422 (N_9422,N_9317,N_9309);
nor U9423 (N_9423,N_9395,N_9326);
or U9424 (N_9424,N_9378,N_9323);
and U9425 (N_9425,N_9322,N_9334);
nand U9426 (N_9426,N_9392,N_9318);
or U9427 (N_9427,N_9342,N_9331);
nand U9428 (N_9428,N_9329,N_9337);
and U9429 (N_9429,N_9306,N_9321);
nand U9430 (N_9430,N_9314,N_9354);
or U9431 (N_9431,N_9382,N_9385);
and U9432 (N_9432,N_9315,N_9389);
and U9433 (N_9433,N_9394,N_9386);
and U9434 (N_9434,N_9359,N_9365);
and U9435 (N_9435,N_9301,N_9332);
or U9436 (N_9436,N_9344,N_9396);
or U9437 (N_9437,N_9351,N_9370);
xnor U9438 (N_9438,N_9361,N_9390);
and U9439 (N_9439,N_9380,N_9312);
and U9440 (N_9440,N_9325,N_9353);
xnor U9441 (N_9441,N_9303,N_9356);
nor U9442 (N_9442,N_9352,N_9369);
xor U9443 (N_9443,N_9371,N_9320);
and U9444 (N_9444,N_9397,N_9349);
or U9445 (N_9445,N_9364,N_9368);
nand U9446 (N_9446,N_9377,N_9379);
and U9447 (N_9447,N_9313,N_9393);
and U9448 (N_9448,N_9391,N_9338);
xor U9449 (N_9449,N_9343,N_9372);
nor U9450 (N_9450,N_9332,N_9368);
and U9451 (N_9451,N_9303,N_9308);
nor U9452 (N_9452,N_9384,N_9366);
nand U9453 (N_9453,N_9320,N_9344);
or U9454 (N_9454,N_9364,N_9366);
and U9455 (N_9455,N_9338,N_9315);
and U9456 (N_9456,N_9394,N_9349);
and U9457 (N_9457,N_9380,N_9321);
nor U9458 (N_9458,N_9370,N_9319);
nand U9459 (N_9459,N_9376,N_9306);
nand U9460 (N_9460,N_9361,N_9322);
xor U9461 (N_9461,N_9364,N_9378);
nor U9462 (N_9462,N_9364,N_9396);
nor U9463 (N_9463,N_9332,N_9309);
and U9464 (N_9464,N_9378,N_9309);
nand U9465 (N_9465,N_9356,N_9354);
xor U9466 (N_9466,N_9396,N_9320);
or U9467 (N_9467,N_9367,N_9391);
nor U9468 (N_9468,N_9354,N_9381);
and U9469 (N_9469,N_9364,N_9388);
and U9470 (N_9470,N_9367,N_9302);
xnor U9471 (N_9471,N_9353,N_9378);
nand U9472 (N_9472,N_9325,N_9373);
or U9473 (N_9473,N_9322,N_9328);
and U9474 (N_9474,N_9320,N_9399);
xor U9475 (N_9475,N_9358,N_9365);
or U9476 (N_9476,N_9306,N_9302);
or U9477 (N_9477,N_9357,N_9353);
nand U9478 (N_9478,N_9315,N_9316);
or U9479 (N_9479,N_9387,N_9383);
or U9480 (N_9480,N_9353,N_9324);
or U9481 (N_9481,N_9367,N_9312);
xor U9482 (N_9482,N_9397,N_9307);
nor U9483 (N_9483,N_9345,N_9302);
nand U9484 (N_9484,N_9312,N_9359);
and U9485 (N_9485,N_9340,N_9342);
or U9486 (N_9486,N_9371,N_9344);
nor U9487 (N_9487,N_9335,N_9304);
nor U9488 (N_9488,N_9361,N_9340);
or U9489 (N_9489,N_9392,N_9397);
xor U9490 (N_9490,N_9344,N_9383);
nand U9491 (N_9491,N_9355,N_9332);
xor U9492 (N_9492,N_9389,N_9381);
xor U9493 (N_9493,N_9328,N_9390);
or U9494 (N_9494,N_9383,N_9397);
and U9495 (N_9495,N_9320,N_9380);
or U9496 (N_9496,N_9342,N_9321);
nand U9497 (N_9497,N_9348,N_9395);
or U9498 (N_9498,N_9303,N_9394);
or U9499 (N_9499,N_9340,N_9360);
nand U9500 (N_9500,N_9464,N_9434);
nor U9501 (N_9501,N_9496,N_9435);
nor U9502 (N_9502,N_9462,N_9487);
and U9503 (N_9503,N_9445,N_9480);
and U9504 (N_9504,N_9473,N_9484);
or U9505 (N_9505,N_9499,N_9483);
xnor U9506 (N_9506,N_9429,N_9472);
and U9507 (N_9507,N_9466,N_9460);
and U9508 (N_9508,N_9448,N_9433);
or U9509 (N_9509,N_9467,N_9410);
nor U9510 (N_9510,N_9489,N_9456);
nor U9511 (N_9511,N_9405,N_9481);
and U9512 (N_9512,N_9401,N_9490);
nand U9513 (N_9513,N_9418,N_9424);
or U9514 (N_9514,N_9408,N_9474);
or U9515 (N_9515,N_9469,N_9409);
or U9516 (N_9516,N_9427,N_9411);
xnor U9517 (N_9517,N_9493,N_9485);
or U9518 (N_9518,N_9439,N_9479);
or U9519 (N_9519,N_9419,N_9422);
xor U9520 (N_9520,N_9415,N_9498);
xnor U9521 (N_9521,N_9416,N_9444);
nand U9522 (N_9522,N_9482,N_9406);
and U9523 (N_9523,N_9438,N_9426);
nand U9524 (N_9524,N_9453,N_9468);
and U9525 (N_9525,N_9454,N_9457);
nor U9526 (N_9526,N_9459,N_9425);
nor U9527 (N_9527,N_9431,N_9470);
nor U9528 (N_9528,N_9437,N_9428);
nor U9529 (N_9529,N_9495,N_9465);
or U9530 (N_9530,N_9423,N_9458);
xor U9531 (N_9531,N_9492,N_9420);
nor U9532 (N_9532,N_9436,N_9451);
or U9533 (N_9533,N_9461,N_9449);
or U9534 (N_9534,N_9494,N_9446);
nor U9535 (N_9535,N_9476,N_9413);
or U9536 (N_9536,N_9402,N_9452);
xor U9537 (N_9537,N_9442,N_9497);
and U9538 (N_9538,N_9430,N_9440);
nand U9539 (N_9539,N_9404,N_9412);
nor U9540 (N_9540,N_9421,N_9403);
xnor U9541 (N_9541,N_9475,N_9407);
or U9542 (N_9542,N_9443,N_9432);
nor U9543 (N_9543,N_9414,N_9478);
and U9544 (N_9544,N_9486,N_9417);
and U9545 (N_9545,N_9471,N_9463);
nand U9546 (N_9546,N_9488,N_9441);
and U9547 (N_9547,N_9400,N_9491);
nor U9548 (N_9548,N_9477,N_9450);
nor U9549 (N_9549,N_9455,N_9447);
xor U9550 (N_9550,N_9495,N_9489);
nor U9551 (N_9551,N_9494,N_9480);
and U9552 (N_9552,N_9491,N_9466);
and U9553 (N_9553,N_9403,N_9430);
nand U9554 (N_9554,N_9492,N_9440);
and U9555 (N_9555,N_9470,N_9402);
nand U9556 (N_9556,N_9439,N_9408);
nor U9557 (N_9557,N_9433,N_9409);
nand U9558 (N_9558,N_9436,N_9443);
xnor U9559 (N_9559,N_9475,N_9491);
xnor U9560 (N_9560,N_9470,N_9406);
and U9561 (N_9561,N_9461,N_9447);
nor U9562 (N_9562,N_9406,N_9401);
and U9563 (N_9563,N_9497,N_9472);
nor U9564 (N_9564,N_9480,N_9406);
nor U9565 (N_9565,N_9491,N_9438);
xnor U9566 (N_9566,N_9479,N_9472);
xnor U9567 (N_9567,N_9493,N_9440);
nand U9568 (N_9568,N_9463,N_9421);
or U9569 (N_9569,N_9488,N_9422);
or U9570 (N_9570,N_9465,N_9490);
xnor U9571 (N_9571,N_9457,N_9470);
or U9572 (N_9572,N_9403,N_9481);
xor U9573 (N_9573,N_9452,N_9492);
and U9574 (N_9574,N_9482,N_9441);
nor U9575 (N_9575,N_9474,N_9455);
nand U9576 (N_9576,N_9402,N_9489);
xor U9577 (N_9577,N_9488,N_9457);
nand U9578 (N_9578,N_9441,N_9439);
or U9579 (N_9579,N_9411,N_9414);
nor U9580 (N_9580,N_9430,N_9454);
nor U9581 (N_9581,N_9434,N_9444);
or U9582 (N_9582,N_9488,N_9456);
and U9583 (N_9583,N_9425,N_9421);
nor U9584 (N_9584,N_9432,N_9495);
and U9585 (N_9585,N_9484,N_9476);
nand U9586 (N_9586,N_9475,N_9422);
nor U9587 (N_9587,N_9455,N_9427);
xor U9588 (N_9588,N_9475,N_9440);
or U9589 (N_9589,N_9446,N_9436);
xor U9590 (N_9590,N_9488,N_9499);
and U9591 (N_9591,N_9408,N_9475);
xnor U9592 (N_9592,N_9439,N_9472);
nand U9593 (N_9593,N_9499,N_9455);
xnor U9594 (N_9594,N_9424,N_9413);
or U9595 (N_9595,N_9442,N_9498);
nand U9596 (N_9596,N_9497,N_9432);
nor U9597 (N_9597,N_9424,N_9486);
nor U9598 (N_9598,N_9475,N_9458);
or U9599 (N_9599,N_9456,N_9468);
nor U9600 (N_9600,N_9507,N_9564);
and U9601 (N_9601,N_9569,N_9591);
nor U9602 (N_9602,N_9585,N_9543);
xor U9603 (N_9603,N_9504,N_9511);
xnor U9604 (N_9604,N_9520,N_9548);
nor U9605 (N_9605,N_9537,N_9573);
and U9606 (N_9606,N_9522,N_9553);
and U9607 (N_9607,N_9536,N_9549);
nand U9608 (N_9608,N_9597,N_9596);
nor U9609 (N_9609,N_9550,N_9515);
nor U9610 (N_9610,N_9586,N_9584);
xor U9611 (N_9611,N_9524,N_9580);
nand U9612 (N_9612,N_9525,N_9516);
xor U9613 (N_9613,N_9535,N_9575);
nor U9614 (N_9614,N_9576,N_9574);
nand U9615 (N_9615,N_9558,N_9508);
nor U9616 (N_9616,N_9503,N_9519);
or U9617 (N_9617,N_9577,N_9599);
nand U9618 (N_9618,N_9560,N_9512);
nand U9619 (N_9619,N_9563,N_9583);
nand U9620 (N_9620,N_9565,N_9534);
nor U9621 (N_9621,N_9559,N_9547);
nand U9622 (N_9622,N_9555,N_9598);
or U9623 (N_9623,N_9566,N_9518);
xor U9624 (N_9624,N_9546,N_9513);
nor U9625 (N_9625,N_9538,N_9593);
and U9626 (N_9626,N_9567,N_9579);
xnor U9627 (N_9627,N_9590,N_9587);
or U9628 (N_9628,N_9545,N_9544);
xor U9629 (N_9629,N_9556,N_9562);
or U9630 (N_9630,N_9500,N_9514);
or U9631 (N_9631,N_9527,N_9592);
or U9632 (N_9632,N_9557,N_9541);
and U9633 (N_9633,N_9581,N_9501);
or U9634 (N_9634,N_9505,N_9540);
xor U9635 (N_9635,N_9570,N_9539);
nor U9636 (N_9636,N_9530,N_9517);
nand U9637 (N_9637,N_9572,N_9506);
nand U9638 (N_9638,N_9552,N_9509);
or U9639 (N_9639,N_9551,N_9528);
nor U9640 (N_9640,N_9568,N_9529);
and U9641 (N_9641,N_9521,N_9561);
xnor U9642 (N_9642,N_9582,N_9533);
nand U9643 (N_9643,N_9526,N_9571);
and U9644 (N_9644,N_9510,N_9532);
or U9645 (N_9645,N_9588,N_9531);
and U9646 (N_9646,N_9523,N_9595);
nand U9647 (N_9647,N_9594,N_9578);
nor U9648 (N_9648,N_9542,N_9554);
nand U9649 (N_9649,N_9502,N_9589);
and U9650 (N_9650,N_9546,N_9582);
nor U9651 (N_9651,N_9565,N_9560);
xnor U9652 (N_9652,N_9595,N_9528);
and U9653 (N_9653,N_9516,N_9511);
or U9654 (N_9654,N_9543,N_9507);
nor U9655 (N_9655,N_9584,N_9599);
and U9656 (N_9656,N_9594,N_9513);
or U9657 (N_9657,N_9565,N_9595);
or U9658 (N_9658,N_9506,N_9584);
and U9659 (N_9659,N_9561,N_9553);
nor U9660 (N_9660,N_9578,N_9548);
nor U9661 (N_9661,N_9510,N_9540);
and U9662 (N_9662,N_9570,N_9525);
nor U9663 (N_9663,N_9575,N_9543);
and U9664 (N_9664,N_9525,N_9562);
and U9665 (N_9665,N_9577,N_9562);
nand U9666 (N_9666,N_9590,N_9556);
nand U9667 (N_9667,N_9592,N_9543);
and U9668 (N_9668,N_9593,N_9568);
nand U9669 (N_9669,N_9515,N_9531);
and U9670 (N_9670,N_9570,N_9551);
or U9671 (N_9671,N_9549,N_9539);
xor U9672 (N_9672,N_9505,N_9567);
nor U9673 (N_9673,N_9573,N_9550);
nor U9674 (N_9674,N_9572,N_9511);
and U9675 (N_9675,N_9595,N_9502);
and U9676 (N_9676,N_9524,N_9570);
nand U9677 (N_9677,N_9509,N_9573);
nand U9678 (N_9678,N_9552,N_9519);
nand U9679 (N_9679,N_9513,N_9598);
nor U9680 (N_9680,N_9558,N_9560);
and U9681 (N_9681,N_9506,N_9538);
nand U9682 (N_9682,N_9570,N_9594);
nor U9683 (N_9683,N_9586,N_9514);
or U9684 (N_9684,N_9518,N_9543);
and U9685 (N_9685,N_9549,N_9550);
or U9686 (N_9686,N_9580,N_9560);
xnor U9687 (N_9687,N_9550,N_9576);
xor U9688 (N_9688,N_9500,N_9517);
and U9689 (N_9689,N_9522,N_9579);
or U9690 (N_9690,N_9571,N_9524);
xor U9691 (N_9691,N_9518,N_9588);
nand U9692 (N_9692,N_9564,N_9505);
xnor U9693 (N_9693,N_9599,N_9518);
nor U9694 (N_9694,N_9566,N_9579);
xnor U9695 (N_9695,N_9559,N_9523);
or U9696 (N_9696,N_9515,N_9537);
nor U9697 (N_9697,N_9504,N_9514);
and U9698 (N_9698,N_9508,N_9584);
and U9699 (N_9699,N_9551,N_9512);
xor U9700 (N_9700,N_9671,N_9614);
xnor U9701 (N_9701,N_9692,N_9690);
xor U9702 (N_9702,N_9681,N_9605);
or U9703 (N_9703,N_9637,N_9627);
nor U9704 (N_9704,N_9630,N_9642);
nor U9705 (N_9705,N_9641,N_9615);
and U9706 (N_9706,N_9662,N_9611);
or U9707 (N_9707,N_9658,N_9680);
nor U9708 (N_9708,N_9607,N_9617);
and U9709 (N_9709,N_9693,N_9687);
or U9710 (N_9710,N_9640,N_9646);
xor U9711 (N_9711,N_9663,N_9612);
or U9712 (N_9712,N_9679,N_9665);
nor U9713 (N_9713,N_9653,N_9623);
nor U9714 (N_9714,N_9686,N_9684);
nand U9715 (N_9715,N_9699,N_9600);
xor U9716 (N_9716,N_9661,N_9628);
and U9717 (N_9717,N_9669,N_9606);
xnor U9718 (N_9718,N_9626,N_9618);
and U9719 (N_9719,N_9644,N_9685);
and U9720 (N_9720,N_9609,N_9672);
nor U9721 (N_9721,N_9650,N_9622);
xor U9722 (N_9722,N_9682,N_9655);
or U9723 (N_9723,N_9602,N_9643);
or U9724 (N_9724,N_9647,N_9619);
nand U9725 (N_9725,N_9675,N_9698);
or U9726 (N_9726,N_9657,N_9688);
and U9727 (N_9727,N_9670,N_9610);
nor U9728 (N_9728,N_9616,N_9678);
nor U9729 (N_9729,N_9632,N_9697);
nor U9730 (N_9730,N_9659,N_9621);
and U9731 (N_9731,N_9634,N_9638);
xnor U9732 (N_9732,N_9668,N_9654);
and U9733 (N_9733,N_9673,N_9656);
and U9734 (N_9734,N_9601,N_9677);
xnor U9735 (N_9735,N_9645,N_9691);
nand U9736 (N_9736,N_9674,N_9695);
nor U9737 (N_9737,N_9625,N_9636);
xnor U9738 (N_9738,N_9676,N_9604);
or U9739 (N_9739,N_9629,N_9649);
nand U9740 (N_9740,N_9631,N_9624);
nor U9741 (N_9741,N_9694,N_9652);
and U9742 (N_9742,N_9664,N_9689);
or U9743 (N_9743,N_9696,N_9666);
and U9744 (N_9744,N_9648,N_9660);
nand U9745 (N_9745,N_9608,N_9603);
nand U9746 (N_9746,N_9639,N_9635);
nor U9747 (N_9747,N_9683,N_9620);
or U9748 (N_9748,N_9667,N_9651);
xor U9749 (N_9749,N_9613,N_9633);
nand U9750 (N_9750,N_9647,N_9630);
nand U9751 (N_9751,N_9612,N_9679);
nand U9752 (N_9752,N_9693,N_9625);
nand U9753 (N_9753,N_9666,N_9687);
nand U9754 (N_9754,N_9630,N_9668);
nor U9755 (N_9755,N_9603,N_9657);
and U9756 (N_9756,N_9679,N_9671);
nor U9757 (N_9757,N_9616,N_9672);
and U9758 (N_9758,N_9664,N_9641);
xnor U9759 (N_9759,N_9694,N_9640);
nor U9760 (N_9760,N_9664,N_9692);
xnor U9761 (N_9761,N_9699,N_9668);
or U9762 (N_9762,N_9609,N_9608);
or U9763 (N_9763,N_9668,N_9611);
nor U9764 (N_9764,N_9668,N_9603);
or U9765 (N_9765,N_9609,N_9654);
and U9766 (N_9766,N_9623,N_9673);
nor U9767 (N_9767,N_9617,N_9689);
and U9768 (N_9768,N_9650,N_9606);
and U9769 (N_9769,N_9688,N_9679);
nand U9770 (N_9770,N_9602,N_9699);
and U9771 (N_9771,N_9610,N_9604);
xor U9772 (N_9772,N_9665,N_9675);
and U9773 (N_9773,N_9621,N_9641);
nand U9774 (N_9774,N_9611,N_9600);
and U9775 (N_9775,N_9668,N_9661);
nand U9776 (N_9776,N_9627,N_9697);
nor U9777 (N_9777,N_9604,N_9645);
xor U9778 (N_9778,N_9613,N_9625);
nor U9779 (N_9779,N_9623,N_9677);
and U9780 (N_9780,N_9606,N_9647);
nor U9781 (N_9781,N_9634,N_9658);
and U9782 (N_9782,N_9673,N_9618);
xnor U9783 (N_9783,N_9623,N_9680);
xor U9784 (N_9784,N_9646,N_9634);
nand U9785 (N_9785,N_9646,N_9661);
nor U9786 (N_9786,N_9658,N_9603);
and U9787 (N_9787,N_9686,N_9673);
xnor U9788 (N_9788,N_9698,N_9693);
nor U9789 (N_9789,N_9628,N_9620);
nor U9790 (N_9790,N_9639,N_9610);
xnor U9791 (N_9791,N_9683,N_9640);
nand U9792 (N_9792,N_9678,N_9674);
and U9793 (N_9793,N_9643,N_9677);
nand U9794 (N_9794,N_9617,N_9610);
or U9795 (N_9795,N_9623,N_9652);
nor U9796 (N_9796,N_9668,N_9656);
nor U9797 (N_9797,N_9608,N_9671);
and U9798 (N_9798,N_9685,N_9613);
xnor U9799 (N_9799,N_9606,N_9662);
nor U9800 (N_9800,N_9723,N_9728);
and U9801 (N_9801,N_9737,N_9739);
or U9802 (N_9802,N_9744,N_9720);
nand U9803 (N_9803,N_9719,N_9769);
or U9804 (N_9804,N_9708,N_9735);
and U9805 (N_9805,N_9792,N_9774);
xnor U9806 (N_9806,N_9732,N_9799);
nand U9807 (N_9807,N_9784,N_9795);
or U9808 (N_9808,N_9789,N_9788);
and U9809 (N_9809,N_9781,N_9714);
nor U9810 (N_9810,N_9700,N_9747);
xnor U9811 (N_9811,N_9791,N_9751);
xnor U9812 (N_9812,N_9725,N_9777);
nand U9813 (N_9813,N_9772,N_9797);
or U9814 (N_9814,N_9766,N_9734);
nor U9815 (N_9815,N_9753,N_9717);
nor U9816 (N_9816,N_9738,N_9706);
xnor U9817 (N_9817,N_9743,N_9780);
or U9818 (N_9818,N_9710,N_9783);
nand U9819 (N_9819,N_9745,N_9730);
and U9820 (N_9820,N_9713,N_9740);
or U9821 (N_9821,N_9731,N_9757);
nand U9822 (N_9822,N_9704,N_9798);
nand U9823 (N_9823,N_9760,N_9768);
or U9824 (N_9824,N_9773,N_9707);
or U9825 (N_9825,N_9721,N_9701);
and U9826 (N_9826,N_9787,N_9771);
nor U9827 (N_9827,N_9748,N_9715);
nor U9828 (N_9828,N_9709,N_9750);
and U9829 (N_9829,N_9765,N_9742);
nand U9830 (N_9830,N_9767,N_9786);
and U9831 (N_9831,N_9729,N_9736);
and U9832 (N_9832,N_9741,N_9727);
or U9833 (N_9833,N_9762,N_9770);
and U9834 (N_9834,N_9782,N_9726);
or U9835 (N_9835,N_9761,N_9716);
and U9836 (N_9836,N_9794,N_9796);
and U9837 (N_9837,N_9722,N_9712);
xor U9838 (N_9838,N_9755,N_9711);
nor U9839 (N_9839,N_9705,N_9793);
nor U9840 (N_9840,N_9703,N_9749);
and U9841 (N_9841,N_9775,N_9759);
or U9842 (N_9842,N_9763,N_9754);
or U9843 (N_9843,N_9724,N_9756);
xor U9844 (N_9844,N_9746,N_9752);
or U9845 (N_9845,N_9779,N_9764);
nor U9846 (N_9846,N_9718,N_9776);
xor U9847 (N_9847,N_9733,N_9778);
and U9848 (N_9848,N_9758,N_9702);
or U9849 (N_9849,N_9785,N_9790);
nand U9850 (N_9850,N_9717,N_9758);
nand U9851 (N_9851,N_9747,N_9714);
xor U9852 (N_9852,N_9708,N_9788);
nor U9853 (N_9853,N_9712,N_9784);
nor U9854 (N_9854,N_9785,N_9771);
or U9855 (N_9855,N_9739,N_9747);
nand U9856 (N_9856,N_9792,N_9713);
nor U9857 (N_9857,N_9721,N_9708);
nor U9858 (N_9858,N_9788,N_9711);
and U9859 (N_9859,N_9720,N_9726);
nand U9860 (N_9860,N_9775,N_9739);
nor U9861 (N_9861,N_9738,N_9746);
nand U9862 (N_9862,N_9798,N_9708);
xnor U9863 (N_9863,N_9788,N_9724);
and U9864 (N_9864,N_9706,N_9731);
and U9865 (N_9865,N_9755,N_9749);
or U9866 (N_9866,N_9713,N_9782);
xor U9867 (N_9867,N_9712,N_9727);
xnor U9868 (N_9868,N_9755,N_9701);
nand U9869 (N_9869,N_9702,N_9796);
nor U9870 (N_9870,N_9785,N_9759);
and U9871 (N_9871,N_9713,N_9711);
and U9872 (N_9872,N_9798,N_9792);
nand U9873 (N_9873,N_9713,N_9724);
nand U9874 (N_9874,N_9758,N_9798);
xnor U9875 (N_9875,N_9770,N_9790);
and U9876 (N_9876,N_9707,N_9746);
nand U9877 (N_9877,N_9718,N_9799);
or U9878 (N_9878,N_9703,N_9788);
and U9879 (N_9879,N_9759,N_9702);
nor U9880 (N_9880,N_9745,N_9736);
or U9881 (N_9881,N_9729,N_9793);
nor U9882 (N_9882,N_9726,N_9730);
xnor U9883 (N_9883,N_9705,N_9704);
xnor U9884 (N_9884,N_9760,N_9769);
nand U9885 (N_9885,N_9763,N_9701);
xnor U9886 (N_9886,N_9791,N_9734);
nand U9887 (N_9887,N_9721,N_9775);
nor U9888 (N_9888,N_9746,N_9782);
or U9889 (N_9889,N_9757,N_9730);
xor U9890 (N_9890,N_9765,N_9747);
xor U9891 (N_9891,N_9742,N_9760);
or U9892 (N_9892,N_9794,N_9746);
and U9893 (N_9893,N_9781,N_9754);
nor U9894 (N_9894,N_9798,N_9701);
nor U9895 (N_9895,N_9704,N_9777);
nand U9896 (N_9896,N_9747,N_9781);
or U9897 (N_9897,N_9782,N_9739);
or U9898 (N_9898,N_9735,N_9780);
nor U9899 (N_9899,N_9759,N_9798);
or U9900 (N_9900,N_9885,N_9807);
nand U9901 (N_9901,N_9882,N_9878);
and U9902 (N_9902,N_9896,N_9826);
nand U9903 (N_9903,N_9804,N_9894);
xnor U9904 (N_9904,N_9845,N_9856);
or U9905 (N_9905,N_9805,N_9869);
nand U9906 (N_9906,N_9834,N_9867);
and U9907 (N_9907,N_9886,N_9838);
or U9908 (N_9908,N_9846,N_9880);
xor U9909 (N_9909,N_9831,N_9810);
or U9910 (N_9910,N_9897,N_9876);
nand U9911 (N_9911,N_9841,N_9888);
nand U9912 (N_9912,N_9854,N_9812);
xnor U9913 (N_9913,N_9803,N_9870);
xor U9914 (N_9914,N_9828,N_9836);
and U9915 (N_9915,N_9879,N_9801);
xnor U9916 (N_9916,N_9815,N_9862);
and U9917 (N_9917,N_9835,N_9844);
nor U9918 (N_9918,N_9814,N_9825);
nor U9919 (N_9919,N_9802,N_9823);
nand U9920 (N_9920,N_9827,N_9893);
xnor U9921 (N_9921,N_9857,N_9850);
xnor U9922 (N_9922,N_9853,N_9830);
and U9923 (N_9923,N_9819,N_9800);
or U9924 (N_9924,N_9892,N_9861);
nand U9925 (N_9925,N_9891,N_9871);
nor U9926 (N_9926,N_9817,N_9872);
and U9927 (N_9927,N_9887,N_9890);
xnor U9928 (N_9928,N_9848,N_9818);
and U9929 (N_9929,N_9813,N_9806);
nor U9930 (N_9930,N_9883,N_9829);
nand U9931 (N_9931,N_9881,N_9809);
and U9932 (N_9932,N_9852,N_9858);
nand U9933 (N_9933,N_9884,N_9816);
nor U9934 (N_9934,N_9849,N_9855);
nand U9935 (N_9935,N_9889,N_9866);
nor U9936 (N_9936,N_9820,N_9842);
nor U9937 (N_9937,N_9899,N_9877);
nor U9938 (N_9938,N_9847,N_9808);
nor U9939 (N_9939,N_9865,N_9833);
nand U9940 (N_9940,N_9860,N_9840);
xor U9941 (N_9941,N_9864,N_9859);
nand U9942 (N_9942,N_9824,N_9839);
nor U9943 (N_9943,N_9821,N_9822);
nor U9944 (N_9944,N_9874,N_9832);
or U9945 (N_9945,N_9843,N_9837);
nor U9946 (N_9946,N_9811,N_9851);
or U9947 (N_9947,N_9863,N_9898);
nor U9948 (N_9948,N_9895,N_9873);
or U9949 (N_9949,N_9868,N_9875);
xor U9950 (N_9950,N_9894,N_9896);
nand U9951 (N_9951,N_9872,N_9889);
or U9952 (N_9952,N_9898,N_9807);
nand U9953 (N_9953,N_9833,N_9816);
nor U9954 (N_9954,N_9899,N_9832);
or U9955 (N_9955,N_9858,N_9895);
and U9956 (N_9956,N_9854,N_9851);
nand U9957 (N_9957,N_9804,N_9887);
nor U9958 (N_9958,N_9868,N_9891);
xnor U9959 (N_9959,N_9844,N_9852);
xnor U9960 (N_9960,N_9843,N_9802);
or U9961 (N_9961,N_9808,N_9812);
xor U9962 (N_9962,N_9835,N_9884);
nand U9963 (N_9963,N_9847,N_9835);
or U9964 (N_9964,N_9874,N_9802);
xor U9965 (N_9965,N_9883,N_9875);
and U9966 (N_9966,N_9894,N_9898);
or U9967 (N_9967,N_9816,N_9870);
and U9968 (N_9968,N_9886,N_9873);
xnor U9969 (N_9969,N_9875,N_9835);
nor U9970 (N_9970,N_9869,N_9816);
xor U9971 (N_9971,N_9800,N_9895);
or U9972 (N_9972,N_9861,N_9837);
xnor U9973 (N_9973,N_9895,N_9874);
nand U9974 (N_9974,N_9801,N_9834);
or U9975 (N_9975,N_9899,N_9894);
and U9976 (N_9976,N_9895,N_9870);
xnor U9977 (N_9977,N_9813,N_9866);
xor U9978 (N_9978,N_9898,N_9819);
or U9979 (N_9979,N_9850,N_9821);
xnor U9980 (N_9980,N_9800,N_9890);
nand U9981 (N_9981,N_9883,N_9861);
xor U9982 (N_9982,N_9851,N_9883);
nand U9983 (N_9983,N_9833,N_9873);
nor U9984 (N_9984,N_9819,N_9828);
nor U9985 (N_9985,N_9807,N_9856);
and U9986 (N_9986,N_9849,N_9891);
and U9987 (N_9987,N_9861,N_9813);
or U9988 (N_9988,N_9858,N_9812);
xnor U9989 (N_9989,N_9867,N_9890);
nand U9990 (N_9990,N_9806,N_9851);
nor U9991 (N_9991,N_9872,N_9873);
or U9992 (N_9992,N_9813,N_9857);
nand U9993 (N_9993,N_9886,N_9868);
and U9994 (N_9994,N_9884,N_9829);
nand U9995 (N_9995,N_9890,N_9883);
nand U9996 (N_9996,N_9818,N_9849);
and U9997 (N_9997,N_9886,N_9877);
or U9998 (N_9998,N_9872,N_9869);
nor U9999 (N_9999,N_9807,N_9897);
or UO_0 (O_0,N_9966,N_9963);
nor UO_1 (O_1,N_9943,N_9985);
nor UO_2 (O_2,N_9925,N_9979);
nand UO_3 (O_3,N_9915,N_9956);
nor UO_4 (O_4,N_9965,N_9914);
and UO_5 (O_5,N_9903,N_9992);
and UO_6 (O_6,N_9958,N_9909);
nor UO_7 (O_7,N_9996,N_9972);
nand UO_8 (O_8,N_9905,N_9951);
nand UO_9 (O_9,N_9994,N_9975);
nand UO_10 (O_10,N_9962,N_9938);
or UO_11 (O_11,N_9982,N_9954);
nor UO_12 (O_12,N_9976,N_9947);
nand UO_13 (O_13,N_9997,N_9939);
xnor UO_14 (O_14,N_9998,N_9901);
xnor UO_15 (O_15,N_9912,N_9987);
or UO_16 (O_16,N_9959,N_9904);
or UO_17 (O_17,N_9967,N_9908);
and UO_18 (O_18,N_9932,N_9906);
and UO_19 (O_19,N_9961,N_9928);
and UO_20 (O_20,N_9920,N_9968);
nor UO_21 (O_21,N_9940,N_9984);
nor UO_22 (O_22,N_9964,N_9937);
or UO_23 (O_23,N_9907,N_9945);
xnor UO_24 (O_24,N_9921,N_9977);
xor UO_25 (O_25,N_9980,N_9936);
xor UO_26 (O_26,N_9924,N_9929);
xor UO_27 (O_27,N_9923,N_9931);
nand UO_28 (O_28,N_9970,N_9910);
nor UO_29 (O_29,N_9974,N_9917);
and UO_30 (O_30,N_9969,N_9973);
nand UO_31 (O_31,N_9955,N_9990);
xor UO_32 (O_32,N_9991,N_9950);
and UO_33 (O_33,N_9900,N_9957);
nand UO_34 (O_34,N_9978,N_9918);
or UO_35 (O_35,N_9948,N_9935);
or UO_36 (O_36,N_9988,N_9926);
and UO_37 (O_37,N_9952,N_9919);
nand UO_38 (O_38,N_9981,N_9989);
or UO_39 (O_39,N_9953,N_9911);
nand UO_40 (O_40,N_9902,N_9960);
nor UO_41 (O_41,N_9983,N_9971);
xnor UO_42 (O_42,N_9933,N_9913);
xnor UO_43 (O_43,N_9946,N_9941);
nor UO_44 (O_44,N_9999,N_9922);
and UO_45 (O_45,N_9993,N_9942);
xnor UO_46 (O_46,N_9944,N_9934);
nor UO_47 (O_47,N_9995,N_9949);
nor UO_48 (O_48,N_9930,N_9916);
nor UO_49 (O_49,N_9927,N_9986);
xor UO_50 (O_50,N_9917,N_9945);
nand UO_51 (O_51,N_9958,N_9904);
or UO_52 (O_52,N_9910,N_9916);
and UO_53 (O_53,N_9939,N_9995);
and UO_54 (O_54,N_9962,N_9908);
xnor UO_55 (O_55,N_9964,N_9910);
nor UO_56 (O_56,N_9975,N_9936);
nand UO_57 (O_57,N_9917,N_9967);
nand UO_58 (O_58,N_9965,N_9962);
xnor UO_59 (O_59,N_9929,N_9981);
and UO_60 (O_60,N_9911,N_9938);
nand UO_61 (O_61,N_9916,N_9992);
or UO_62 (O_62,N_9907,N_9980);
nor UO_63 (O_63,N_9933,N_9972);
or UO_64 (O_64,N_9968,N_9992);
nand UO_65 (O_65,N_9942,N_9964);
or UO_66 (O_66,N_9920,N_9917);
xnor UO_67 (O_67,N_9998,N_9959);
or UO_68 (O_68,N_9956,N_9985);
xnor UO_69 (O_69,N_9911,N_9906);
or UO_70 (O_70,N_9909,N_9906);
nor UO_71 (O_71,N_9962,N_9985);
xor UO_72 (O_72,N_9955,N_9925);
nand UO_73 (O_73,N_9920,N_9907);
and UO_74 (O_74,N_9940,N_9927);
or UO_75 (O_75,N_9925,N_9938);
or UO_76 (O_76,N_9990,N_9923);
or UO_77 (O_77,N_9904,N_9927);
nand UO_78 (O_78,N_9946,N_9970);
or UO_79 (O_79,N_9987,N_9909);
or UO_80 (O_80,N_9961,N_9951);
and UO_81 (O_81,N_9959,N_9961);
nand UO_82 (O_82,N_9995,N_9967);
xor UO_83 (O_83,N_9950,N_9970);
or UO_84 (O_84,N_9924,N_9922);
nand UO_85 (O_85,N_9992,N_9915);
and UO_86 (O_86,N_9958,N_9963);
or UO_87 (O_87,N_9914,N_9987);
nand UO_88 (O_88,N_9957,N_9985);
nor UO_89 (O_89,N_9918,N_9939);
and UO_90 (O_90,N_9949,N_9920);
nor UO_91 (O_91,N_9948,N_9932);
and UO_92 (O_92,N_9996,N_9955);
nor UO_93 (O_93,N_9980,N_9900);
and UO_94 (O_94,N_9989,N_9900);
nor UO_95 (O_95,N_9952,N_9949);
nand UO_96 (O_96,N_9981,N_9935);
or UO_97 (O_97,N_9924,N_9975);
nand UO_98 (O_98,N_9910,N_9942);
or UO_99 (O_99,N_9930,N_9998);
nor UO_100 (O_100,N_9932,N_9983);
and UO_101 (O_101,N_9900,N_9942);
nor UO_102 (O_102,N_9995,N_9990);
or UO_103 (O_103,N_9987,N_9904);
and UO_104 (O_104,N_9934,N_9993);
nand UO_105 (O_105,N_9901,N_9958);
or UO_106 (O_106,N_9960,N_9982);
nand UO_107 (O_107,N_9935,N_9901);
nand UO_108 (O_108,N_9945,N_9948);
and UO_109 (O_109,N_9948,N_9983);
and UO_110 (O_110,N_9981,N_9994);
or UO_111 (O_111,N_9953,N_9932);
nor UO_112 (O_112,N_9920,N_9940);
xnor UO_113 (O_113,N_9941,N_9957);
nand UO_114 (O_114,N_9922,N_9955);
or UO_115 (O_115,N_9929,N_9977);
nand UO_116 (O_116,N_9932,N_9980);
xor UO_117 (O_117,N_9951,N_9911);
or UO_118 (O_118,N_9950,N_9943);
nand UO_119 (O_119,N_9904,N_9928);
and UO_120 (O_120,N_9954,N_9987);
xnor UO_121 (O_121,N_9983,N_9928);
nand UO_122 (O_122,N_9933,N_9947);
xnor UO_123 (O_123,N_9924,N_9912);
and UO_124 (O_124,N_9945,N_9994);
xnor UO_125 (O_125,N_9984,N_9990);
nand UO_126 (O_126,N_9923,N_9997);
and UO_127 (O_127,N_9967,N_9949);
nor UO_128 (O_128,N_9932,N_9993);
nor UO_129 (O_129,N_9951,N_9901);
and UO_130 (O_130,N_9931,N_9961);
and UO_131 (O_131,N_9974,N_9922);
nor UO_132 (O_132,N_9957,N_9925);
or UO_133 (O_133,N_9921,N_9963);
xnor UO_134 (O_134,N_9954,N_9943);
nor UO_135 (O_135,N_9949,N_9923);
or UO_136 (O_136,N_9943,N_9923);
nand UO_137 (O_137,N_9983,N_9939);
or UO_138 (O_138,N_9973,N_9939);
and UO_139 (O_139,N_9995,N_9938);
nand UO_140 (O_140,N_9990,N_9910);
and UO_141 (O_141,N_9928,N_9907);
or UO_142 (O_142,N_9906,N_9976);
nand UO_143 (O_143,N_9993,N_9939);
nor UO_144 (O_144,N_9971,N_9915);
nor UO_145 (O_145,N_9981,N_9946);
nor UO_146 (O_146,N_9941,N_9966);
nor UO_147 (O_147,N_9924,N_9963);
xnor UO_148 (O_148,N_9926,N_9936);
nor UO_149 (O_149,N_9916,N_9909);
nand UO_150 (O_150,N_9983,N_9974);
nor UO_151 (O_151,N_9926,N_9992);
and UO_152 (O_152,N_9948,N_9950);
nor UO_153 (O_153,N_9993,N_9994);
or UO_154 (O_154,N_9931,N_9972);
or UO_155 (O_155,N_9906,N_9929);
and UO_156 (O_156,N_9908,N_9910);
or UO_157 (O_157,N_9969,N_9971);
xor UO_158 (O_158,N_9979,N_9999);
nand UO_159 (O_159,N_9963,N_9936);
xor UO_160 (O_160,N_9973,N_9909);
nand UO_161 (O_161,N_9996,N_9936);
nand UO_162 (O_162,N_9928,N_9941);
xnor UO_163 (O_163,N_9918,N_9913);
xnor UO_164 (O_164,N_9982,N_9924);
and UO_165 (O_165,N_9959,N_9997);
and UO_166 (O_166,N_9995,N_9923);
nand UO_167 (O_167,N_9959,N_9941);
and UO_168 (O_168,N_9931,N_9940);
nand UO_169 (O_169,N_9973,N_9953);
or UO_170 (O_170,N_9992,N_9952);
or UO_171 (O_171,N_9939,N_9977);
or UO_172 (O_172,N_9953,N_9942);
and UO_173 (O_173,N_9992,N_9921);
nor UO_174 (O_174,N_9958,N_9965);
or UO_175 (O_175,N_9972,N_9915);
or UO_176 (O_176,N_9927,N_9929);
xor UO_177 (O_177,N_9966,N_9971);
xor UO_178 (O_178,N_9934,N_9926);
or UO_179 (O_179,N_9932,N_9910);
and UO_180 (O_180,N_9919,N_9926);
xnor UO_181 (O_181,N_9927,N_9965);
and UO_182 (O_182,N_9975,N_9968);
nor UO_183 (O_183,N_9924,N_9923);
nor UO_184 (O_184,N_9967,N_9968);
and UO_185 (O_185,N_9993,N_9906);
or UO_186 (O_186,N_9991,N_9937);
or UO_187 (O_187,N_9932,N_9974);
and UO_188 (O_188,N_9902,N_9972);
xor UO_189 (O_189,N_9963,N_9904);
and UO_190 (O_190,N_9981,N_9913);
and UO_191 (O_191,N_9914,N_9955);
nand UO_192 (O_192,N_9943,N_9920);
nand UO_193 (O_193,N_9943,N_9933);
nand UO_194 (O_194,N_9908,N_9949);
nor UO_195 (O_195,N_9905,N_9919);
nor UO_196 (O_196,N_9969,N_9988);
and UO_197 (O_197,N_9925,N_9978);
or UO_198 (O_198,N_9984,N_9915);
xor UO_199 (O_199,N_9963,N_9948);
or UO_200 (O_200,N_9961,N_9974);
nor UO_201 (O_201,N_9972,N_9927);
or UO_202 (O_202,N_9937,N_9936);
nor UO_203 (O_203,N_9944,N_9915);
nand UO_204 (O_204,N_9947,N_9931);
and UO_205 (O_205,N_9969,N_9917);
nor UO_206 (O_206,N_9907,N_9918);
nand UO_207 (O_207,N_9925,N_9960);
nand UO_208 (O_208,N_9936,N_9925);
nand UO_209 (O_209,N_9941,N_9944);
nor UO_210 (O_210,N_9929,N_9948);
and UO_211 (O_211,N_9918,N_9914);
nor UO_212 (O_212,N_9944,N_9996);
or UO_213 (O_213,N_9974,N_9946);
xor UO_214 (O_214,N_9925,N_9941);
xnor UO_215 (O_215,N_9977,N_9954);
nor UO_216 (O_216,N_9977,N_9957);
nor UO_217 (O_217,N_9918,N_9916);
nand UO_218 (O_218,N_9992,N_9964);
and UO_219 (O_219,N_9939,N_9967);
and UO_220 (O_220,N_9908,N_9917);
or UO_221 (O_221,N_9914,N_9945);
or UO_222 (O_222,N_9931,N_9945);
nor UO_223 (O_223,N_9934,N_9953);
xnor UO_224 (O_224,N_9965,N_9959);
nor UO_225 (O_225,N_9976,N_9958);
or UO_226 (O_226,N_9955,N_9942);
or UO_227 (O_227,N_9927,N_9984);
nand UO_228 (O_228,N_9941,N_9909);
xnor UO_229 (O_229,N_9984,N_9965);
nand UO_230 (O_230,N_9975,N_9937);
xnor UO_231 (O_231,N_9912,N_9977);
or UO_232 (O_232,N_9950,N_9931);
xnor UO_233 (O_233,N_9912,N_9983);
nand UO_234 (O_234,N_9912,N_9958);
nor UO_235 (O_235,N_9920,N_9948);
or UO_236 (O_236,N_9906,N_9962);
nor UO_237 (O_237,N_9944,N_9946);
xor UO_238 (O_238,N_9946,N_9999);
or UO_239 (O_239,N_9954,N_9946);
or UO_240 (O_240,N_9994,N_9964);
nor UO_241 (O_241,N_9919,N_9906);
nor UO_242 (O_242,N_9910,N_9971);
or UO_243 (O_243,N_9929,N_9943);
and UO_244 (O_244,N_9947,N_9904);
or UO_245 (O_245,N_9946,N_9900);
nor UO_246 (O_246,N_9978,N_9951);
nand UO_247 (O_247,N_9902,N_9971);
or UO_248 (O_248,N_9954,N_9930);
or UO_249 (O_249,N_9976,N_9987);
or UO_250 (O_250,N_9996,N_9900);
and UO_251 (O_251,N_9932,N_9925);
or UO_252 (O_252,N_9997,N_9932);
xor UO_253 (O_253,N_9980,N_9953);
xor UO_254 (O_254,N_9931,N_9968);
xnor UO_255 (O_255,N_9936,N_9956);
nor UO_256 (O_256,N_9933,N_9961);
and UO_257 (O_257,N_9908,N_9957);
nand UO_258 (O_258,N_9998,N_9991);
xor UO_259 (O_259,N_9963,N_9915);
nand UO_260 (O_260,N_9983,N_9991);
and UO_261 (O_261,N_9978,N_9953);
and UO_262 (O_262,N_9995,N_9919);
nor UO_263 (O_263,N_9965,N_9936);
nand UO_264 (O_264,N_9993,N_9997);
and UO_265 (O_265,N_9990,N_9911);
or UO_266 (O_266,N_9937,N_9902);
and UO_267 (O_267,N_9908,N_9921);
xnor UO_268 (O_268,N_9953,N_9941);
and UO_269 (O_269,N_9911,N_9999);
nor UO_270 (O_270,N_9919,N_9966);
or UO_271 (O_271,N_9929,N_9990);
and UO_272 (O_272,N_9951,N_9908);
xnor UO_273 (O_273,N_9986,N_9912);
nor UO_274 (O_274,N_9907,N_9978);
nor UO_275 (O_275,N_9939,N_9921);
xnor UO_276 (O_276,N_9919,N_9908);
xnor UO_277 (O_277,N_9910,N_9980);
nand UO_278 (O_278,N_9920,N_9981);
and UO_279 (O_279,N_9900,N_9969);
nor UO_280 (O_280,N_9929,N_9946);
nor UO_281 (O_281,N_9944,N_9980);
nor UO_282 (O_282,N_9913,N_9998);
nand UO_283 (O_283,N_9919,N_9911);
and UO_284 (O_284,N_9987,N_9930);
or UO_285 (O_285,N_9939,N_9940);
nand UO_286 (O_286,N_9978,N_9945);
nor UO_287 (O_287,N_9930,N_9984);
and UO_288 (O_288,N_9996,N_9925);
nor UO_289 (O_289,N_9957,N_9915);
nand UO_290 (O_290,N_9933,N_9942);
xnor UO_291 (O_291,N_9921,N_9925);
or UO_292 (O_292,N_9924,N_9961);
and UO_293 (O_293,N_9947,N_9991);
and UO_294 (O_294,N_9911,N_9943);
xnor UO_295 (O_295,N_9916,N_9960);
nand UO_296 (O_296,N_9901,N_9968);
nor UO_297 (O_297,N_9959,N_9908);
nand UO_298 (O_298,N_9971,N_9922);
xor UO_299 (O_299,N_9989,N_9905);
and UO_300 (O_300,N_9926,N_9980);
xnor UO_301 (O_301,N_9907,N_9933);
nor UO_302 (O_302,N_9910,N_9904);
or UO_303 (O_303,N_9980,N_9940);
nor UO_304 (O_304,N_9911,N_9967);
xnor UO_305 (O_305,N_9901,N_9911);
nand UO_306 (O_306,N_9995,N_9932);
and UO_307 (O_307,N_9903,N_9957);
xor UO_308 (O_308,N_9933,N_9901);
or UO_309 (O_309,N_9931,N_9951);
nor UO_310 (O_310,N_9927,N_9938);
or UO_311 (O_311,N_9943,N_9915);
and UO_312 (O_312,N_9990,N_9979);
and UO_313 (O_313,N_9984,N_9988);
or UO_314 (O_314,N_9991,N_9946);
nand UO_315 (O_315,N_9951,N_9932);
or UO_316 (O_316,N_9913,N_9983);
or UO_317 (O_317,N_9970,N_9976);
and UO_318 (O_318,N_9928,N_9934);
nor UO_319 (O_319,N_9905,N_9975);
and UO_320 (O_320,N_9991,N_9935);
xor UO_321 (O_321,N_9925,N_9974);
xor UO_322 (O_322,N_9996,N_9984);
nor UO_323 (O_323,N_9960,N_9966);
and UO_324 (O_324,N_9969,N_9993);
nor UO_325 (O_325,N_9976,N_9942);
xor UO_326 (O_326,N_9974,N_9935);
xnor UO_327 (O_327,N_9964,N_9954);
and UO_328 (O_328,N_9973,N_9934);
nand UO_329 (O_329,N_9935,N_9961);
xor UO_330 (O_330,N_9905,N_9928);
nand UO_331 (O_331,N_9959,N_9953);
or UO_332 (O_332,N_9915,N_9931);
and UO_333 (O_333,N_9959,N_9986);
and UO_334 (O_334,N_9960,N_9977);
or UO_335 (O_335,N_9989,N_9923);
or UO_336 (O_336,N_9967,N_9952);
or UO_337 (O_337,N_9907,N_9923);
nor UO_338 (O_338,N_9941,N_9936);
nand UO_339 (O_339,N_9924,N_9936);
or UO_340 (O_340,N_9961,N_9968);
xor UO_341 (O_341,N_9914,N_9966);
and UO_342 (O_342,N_9969,N_9987);
xor UO_343 (O_343,N_9906,N_9912);
nor UO_344 (O_344,N_9964,N_9924);
xnor UO_345 (O_345,N_9934,N_9940);
xor UO_346 (O_346,N_9930,N_9973);
nor UO_347 (O_347,N_9925,N_9926);
nand UO_348 (O_348,N_9987,N_9947);
nor UO_349 (O_349,N_9926,N_9945);
nand UO_350 (O_350,N_9919,N_9992);
nand UO_351 (O_351,N_9983,N_9988);
or UO_352 (O_352,N_9969,N_9963);
nor UO_353 (O_353,N_9963,N_9906);
nand UO_354 (O_354,N_9973,N_9985);
or UO_355 (O_355,N_9985,N_9986);
or UO_356 (O_356,N_9986,N_9928);
xnor UO_357 (O_357,N_9906,N_9941);
and UO_358 (O_358,N_9933,N_9996);
nor UO_359 (O_359,N_9991,N_9913);
nor UO_360 (O_360,N_9944,N_9924);
nand UO_361 (O_361,N_9985,N_9983);
or UO_362 (O_362,N_9986,N_9968);
nand UO_363 (O_363,N_9976,N_9901);
xor UO_364 (O_364,N_9925,N_9937);
nand UO_365 (O_365,N_9993,N_9933);
nand UO_366 (O_366,N_9936,N_9950);
and UO_367 (O_367,N_9998,N_9995);
nor UO_368 (O_368,N_9990,N_9953);
nor UO_369 (O_369,N_9958,N_9966);
nor UO_370 (O_370,N_9994,N_9935);
and UO_371 (O_371,N_9924,N_9960);
or UO_372 (O_372,N_9964,N_9965);
nor UO_373 (O_373,N_9951,N_9960);
nor UO_374 (O_374,N_9933,N_9992);
nor UO_375 (O_375,N_9922,N_9985);
and UO_376 (O_376,N_9933,N_9988);
and UO_377 (O_377,N_9910,N_9967);
or UO_378 (O_378,N_9967,N_9919);
xnor UO_379 (O_379,N_9944,N_9995);
or UO_380 (O_380,N_9945,N_9959);
nand UO_381 (O_381,N_9912,N_9901);
or UO_382 (O_382,N_9923,N_9940);
nand UO_383 (O_383,N_9927,N_9909);
nand UO_384 (O_384,N_9939,N_9910);
nor UO_385 (O_385,N_9968,N_9981);
nand UO_386 (O_386,N_9926,N_9907);
xnor UO_387 (O_387,N_9954,N_9921);
xor UO_388 (O_388,N_9998,N_9943);
nor UO_389 (O_389,N_9995,N_9904);
xor UO_390 (O_390,N_9995,N_9952);
nor UO_391 (O_391,N_9953,N_9943);
nand UO_392 (O_392,N_9956,N_9970);
nand UO_393 (O_393,N_9908,N_9974);
or UO_394 (O_394,N_9906,N_9961);
or UO_395 (O_395,N_9953,N_9931);
nor UO_396 (O_396,N_9951,N_9965);
nor UO_397 (O_397,N_9956,N_9928);
xnor UO_398 (O_398,N_9915,N_9904);
nand UO_399 (O_399,N_9963,N_9998);
and UO_400 (O_400,N_9943,N_9977);
xor UO_401 (O_401,N_9979,N_9969);
nand UO_402 (O_402,N_9962,N_9959);
or UO_403 (O_403,N_9937,N_9966);
xor UO_404 (O_404,N_9951,N_9985);
or UO_405 (O_405,N_9970,N_9915);
and UO_406 (O_406,N_9914,N_9959);
nand UO_407 (O_407,N_9945,N_9927);
xor UO_408 (O_408,N_9996,N_9992);
nand UO_409 (O_409,N_9948,N_9930);
xnor UO_410 (O_410,N_9958,N_9936);
or UO_411 (O_411,N_9944,N_9966);
and UO_412 (O_412,N_9922,N_9960);
and UO_413 (O_413,N_9982,N_9928);
nand UO_414 (O_414,N_9904,N_9994);
and UO_415 (O_415,N_9998,N_9979);
nor UO_416 (O_416,N_9973,N_9984);
or UO_417 (O_417,N_9950,N_9905);
or UO_418 (O_418,N_9926,N_9962);
xnor UO_419 (O_419,N_9997,N_9969);
xor UO_420 (O_420,N_9997,N_9912);
xor UO_421 (O_421,N_9920,N_9929);
xor UO_422 (O_422,N_9903,N_9927);
and UO_423 (O_423,N_9949,N_9968);
xnor UO_424 (O_424,N_9991,N_9933);
nand UO_425 (O_425,N_9975,N_9934);
nor UO_426 (O_426,N_9992,N_9907);
nor UO_427 (O_427,N_9978,N_9931);
and UO_428 (O_428,N_9964,N_9915);
nor UO_429 (O_429,N_9917,N_9994);
xnor UO_430 (O_430,N_9929,N_9914);
and UO_431 (O_431,N_9924,N_9930);
and UO_432 (O_432,N_9921,N_9931);
xnor UO_433 (O_433,N_9937,N_9944);
nand UO_434 (O_434,N_9903,N_9919);
and UO_435 (O_435,N_9949,N_9941);
and UO_436 (O_436,N_9973,N_9938);
nand UO_437 (O_437,N_9936,N_9907);
nand UO_438 (O_438,N_9903,N_9951);
or UO_439 (O_439,N_9988,N_9932);
xnor UO_440 (O_440,N_9954,N_9910);
and UO_441 (O_441,N_9916,N_9998);
nor UO_442 (O_442,N_9997,N_9952);
nand UO_443 (O_443,N_9974,N_9960);
xor UO_444 (O_444,N_9979,N_9924);
xor UO_445 (O_445,N_9940,N_9905);
nand UO_446 (O_446,N_9971,N_9937);
nand UO_447 (O_447,N_9978,N_9961);
nor UO_448 (O_448,N_9913,N_9904);
and UO_449 (O_449,N_9901,N_9904);
nor UO_450 (O_450,N_9926,N_9991);
or UO_451 (O_451,N_9901,N_9910);
and UO_452 (O_452,N_9935,N_9949);
nand UO_453 (O_453,N_9950,N_9995);
and UO_454 (O_454,N_9927,N_9912);
nand UO_455 (O_455,N_9998,N_9950);
or UO_456 (O_456,N_9983,N_9973);
nor UO_457 (O_457,N_9999,N_9945);
and UO_458 (O_458,N_9991,N_9993);
and UO_459 (O_459,N_9924,N_9965);
nor UO_460 (O_460,N_9957,N_9949);
nor UO_461 (O_461,N_9908,N_9964);
nand UO_462 (O_462,N_9944,N_9909);
and UO_463 (O_463,N_9952,N_9936);
xor UO_464 (O_464,N_9967,N_9973);
or UO_465 (O_465,N_9969,N_9952);
and UO_466 (O_466,N_9904,N_9983);
nor UO_467 (O_467,N_9934,N_9999);
or UO_468 (O_468,N_9945,N_9980);
and UO_469 (O_469,N_9914,N_9915);
or UO_470 (O_470,N_9984,N_9923);
and UO_471 (O_471,N_9951,N_9976);
nand UO_472 (O_472,N_9971,N_9914);
xor UO_473 (O_473,N_9939,N_9917);
or UO_474 (O_474,N_9961,N_9985);
nand UO_475 (O_475,N_9958,N_9970);
and UO_476 (O_476,N_9922,N_9940);
and UO_477 (O_477,N_9930,N_9952);
nor UO_478 (O_478,N_9945,N_9942);
nand UO_479 (O_479,N_9995,N_9907);
xor UO_480 (O_480,N_9918,N_9934);
xor UO_481 (O_481,N_9964,N_9926);
nand UO_482 (O_482,N_9969,N_9926);
nor UO_483 (O_483,N_9988,N_9900);
nor UO_484 (O_484,N_9919,N_9933);
or UO_485 (O_485,N_9900,N_9972);
or UO_486 (O_486,N_9907,N_9902);
nor UO_487 (O_487,N_9971,N_9944);
and UO_488 (O_488,N_9999,N_9905);
xnor UO_489 (O_489,N_9909,N_9954);
nor UO_490 (O_490,N_9993,N_9920);
xor UO_491 (O_491,N_9914,N_9981);
nor UO_492 (O_492,N_9950,N_9992);
or UO_493 (O_493,N_9912,N_9936);
or UO_494 (O_494,N_9971,N_9901);
and UO_495 (O_495,N_9918,N_9923);
nor UO_496 (O_496,N_9957,N_9982);
nor UO_497 (O_497,N_9904,N_9979);
and UO_498 (O_498,N_9924,N_9916);
or UO_499 (O_499,N_9978,N_9976);
and UO_500 (O_500,N_9935,N_9989);
and UO_501 (O_501,N_9993,N_9974);
nor UO_502 (O_502,N_9924,N_9977);
xor UO_503 (O_503,N_9988,N_9936);
nand UO_504 (O_504,N_9921,N_9972);
nand UO_505 (O_505,N_9987,N_9925);
xnor UO_506 (O_506,N_9902,N_9923);
or UO_507 (O_507,N_9980,N_9977);
or UO_508 (O_508,N_9941,N_9992);
nand UO_509 (O_509,N_9930,N_9911);
nor UO_510 (O_510,N_9922,N_9958);
nand UO_511 (O_511,N_9908,N_9946);
xnor UO_512 (O_512,N_9962,N_9990);
or UO_513 (O_513,N_9987,N_9988);
nand UO_514 (O_514,N_9997,N_9918);
and UO_515 (O_515,N_9994,N_9983);
and UO_516 (O_516,N_9925,N_9970);
nand UO_517 (O_517,N_9989,N_9920);
and UO_518 (O_518,N_9977,N_9940);
xnor UO_519 (O_519,N_9927,N_9953);
nand UO_520 (O_520,N_9990,N_9970);
xor UO_521 (O_521,N_9988,N_9915);
or UO_522 (O_522,N_9980,N_9924);
and UO_523 (O_523,N_9923,N_9926);
nor UO_524 (O_524,N_9961,N_9922);
or UO_525 (O_525,N_9989,N_9931);
nand UO_526 (O_526,N_9902,N_9984);
nand UO_527 (O_527,N_9923,N_9964);
and UO_528 (O_528,N_9928,N_9968);
xor UO_529 (O_529,N_9993,N_9938);
nand UO_530 (O_530,N_9913,N_9992);
or UO_531 (O_531,N_9936,N_9946);
or UO_532 (O_532,N_9936,N_9944);
nand UO_533 (O_533,N_9930,N_9901);
and UO_534 (O_534,N_9964,N_9932);
xnor UO_535 (O_535,N_9912,N_9943);
or UO_536 (O_536,N_9968,N_9964);
nand UO_537 (O_537,N_9966,N_9992);
and UO_538 (O_538,N_9928,N_9950);
nor UO_539 (O_539,N_9952,N_9941);
and UO_540 (O_540,N_9968,N_9970);
or UO_541 (O_541,N_9901,N_9994);
xor UO_542 (O_542,N_9987,N_9927);
xor UO_543 (O_543,N_9949,N_9915);
nor UO_544 (O_544,N_9953,N_9933);
or UO_545 (O_545,N_9913,N_9962);
nor UO_546 (O_546,N_9923,N_9978);
or UO_547 (O_547,N_9965,N_9969);
xnor UO_548 (O_548,N_9980,N_9985);
and UO_549 (O_549,N_9917,N_9933);
or UO_550 (O_550,N_9925,N_9975);
nand UO_551 (O_551,N_9919,N_9976);
or UO_552 (O_552,N_9934,N_9931);
nor UO_553 (O_553,N_9922,N_9901);
xnor UO_554 (O_554,N_9978,N_9929);
nand UO_555 (O_555,N_9961,N_9921);
xnor UO_556 (O_556,N_9996,N_9969);
or UO_557 (O_557,N_9930,N_9963);
nor UO_558 (O_558,N_9969,N_9923);
nand UO_559 (O_559,N_9910,N_9965);
nand UO_560 (O_560,N_9991,N_9905);
nor UO_561 (O_561,N_9986,N_9974);
nand UO_562 (O_562,N_9983,N_9930);
nand UO_563 (O_563,N_9944,N_9904);
xor UO_564 (O_564,N_9909,N_9924);
and UO_565 (O_565,N_9961,N_9992);
nor UO_566 (O_566,N_9955,N_9950);
nand UO_567 (O_567,N_9929,N_9974);
nand UO_568 (O_568,N_9929,N_9910);
and UO_569 (O_569,N_9939,N_9905);
nor UO_570 (O_570,N_9918,N_9973);
and UO_571 (O_571,N_9960,N_9904);
and UO_572 (O_572,N_9975,N_9992);
xnor UO_573 (O_573,N_9982,N_9909);
or UO_574 (O_574,N_9936,N_9991);
and UO_575 (O_575,N_9950,N_9994);
nand UO_576 (O_576,N_9916,N_9997);
or UO_577 (O_577,N_9986,N_9981);
nand UO_578 (O_578,N_9914,N_9901);
or UO_579 (O_579,N_9933,N_9998);
xor UO_580 (O_580,N_9997,N_9973);
or UO_581 (O_581,N_9930,N_9957);
and UO_582 (O_582,N_9908,N_9983);
and UO_583 (O_583,N_9998,N_9974);
nor UO_584 (O_584,N_9972,N_9971);
or UO_585 (O_585,N_9947,N_9906);
or UO_586 (O_586,N_9914,N_9932);
and UO_587 (O_587,N_9965,N_9932);
nand UO_588 (O_588,N_9941,N_9942);
and UO_589 (O_589,N_9935,N_9916);
nor UO_590 (O_590,N_9953,N_9923);
and UO_591 (O_591,N_9934,N_9958);
and UO_592 (O_592,N_9931,N_9962);
nand UO_593 (O_593,N_9969,N_9922);
nand UO_594 (O_594,N_9918,N_9984);
nor UO_595 (O_595,N_9976,N_9975);
xor UO_596 (O_596,N_9945,N_9955);
xnor UO_597 (O_597,N_9961,N_9918);
nor UO_598 (O_598,N_9987,N_9931);
nand UO_599 (O_599,N_9944,N_9962);
nand UO_600 (O_600,N_9938,N_9916);
nor UO_601 (O_601,N_9958,N_9972);
nor UO_602 (O_602,N_9923,N_9983);
or UO_603 (O_603,N_9999,N_9963);
nor UO_604 (O_604,N_9932,N_9923);
and UO_605 (O_605,N_9907,N_9954);
or UO_606 (O_606,N_9927,N_9931);
nor UO_607 (O_607,N_9948,N_9958);
nor UO_608 (O_608,N_9914,N_9902);
nor UO_609 (O_609,N_9916,N_9996);
or UO_610 (O_610,N_9911,N_9983);
xnor UO_611 (O_611,N_9991,N_9954);
nor UO_612 (O_612,N_9947,N_9919);
and UO_613 (O_613,N_9979,N_9917);
and UO_614 (O_614,N_9954,N_9970);
and UO_615 (O_615,N_9983,N_9918);
or UO_616 (O_616,N_9924,N_9949);
and UO_617 (O_617,N_9977,N_9947);
and UO_618 (O_618,N_9965,N_9941);
nand UO_619 (O_619,N_9957,N_9963);
or UO_620 (O_620,N_9946,N_9935);
and UO_621 (O_621,N_9991,N_9930);
nand UO_622 (O_622,N_9990,N_9915);
nand UO_623 (O_623,N_9933,N_9900);
and UO_624 (O_624,N_9959,N_9972);
nand UO_625 (O_625,N_9965,N_9975);
xor UO_626 (O_626,N_9939,N_9946);
and UO_627 (O_627,N_9920,N_9970);
or UO_628 (O_628,N_9923,N_9937);
xor UO_629 (O_629,N_9950,N_9907);
nor UO_630 (O_630,N_9983,N_9986);
and UO_631 (O_631,N_9952,N_9905);
and UO_632 (O_632,N_9991,N_9996);
and UO_633 (O_633,N_9941,N_9969);
nor UO_634 (O_634,N_9972,N_9924);
and UO_635 (O_635,N_9995,N_9958);
nor UO_636 (O_636,N_9975,N_9951);
xor UO_637 (O_637,N_9959,N_9970);
nand UO_638 (O_638,N_9996,N_9980);
xor UO_639 (O_639,N_9928,N_9972);
or UO_640 (O_640,N_9963,N_9900);
nor UO_641 (O_641,N_9948,N_9986);
or UO_642 (O_642,N_9961,N_9997);
xnor UO_643 (O_643,N_9900,N_9956);
and UO_644 (O_644,N_9957,N_9989);
nand UO_645 (O_645,N_9948,N_9936);
nor UO_646 (O_646,N_9942,N_9988);
xnor UO_647 (O_647,N_9997,N_9953);
nand UO_648 (O_648,N_9993,N_9915);
nand UO_649 (O_649,N_9955,N_9995);
or UO_650 (O_650,N_9976,N_9912);
xor UO_651 (O_651,N_9922,N_9972);
nor UO_652 (O_652,N_9918,N_9966);
nor UO_653 (O_653,N_9912,N_9940);
nand UO_654 (O_654,N_9959,N_9943);
nand UO_655 (O_655,N_9967,N_9927);
or UO_656 (O_656,N_9900,N_9986);
and UO_657 (O_657,N_9999,N_9948);
or UO_658 (O_658,N_9924,N_9956);
xor UO_659 (O_659,N_9979,N_9972);
nand UO_660 (O_660,N_9985,N_9900);
xnor UO_661 (O_661,N_9987,N_9982);
and UO_662 (O_662,N_9971,N_9928);
or UO_663 (O_663,N_9924,N_9902);
nor UO_664 (O_664,N_9907,N_9942);
nor UO_665 (O_665,N_9923,N_9914);
or UO_666 (O_666,N_9921,N_9951);
xor UO_667 (O_667,N_9994,N_9990);
xor UO_668 (O_668,N_9996,N_9956);
or UO_669 (O_669,N_9993,N_9964);
and UO_670 (O_670,N_9929,N_9938);
or UO_671 (O_671,N_9949,N_9910);
xnor UO_672 (O_672,N_9944,N_9908);
nor UO_673 (O_673,N_9985,N_9989);
xor UO_674 (O_674,N_9956,N_9950);
nand UO_675 (O_675,N_9911,N_9925);
nor UO_676 (O_676,N_9988,N_9977);
or UO_677 (O_677,N_9965,N_9997);
and UO_678 (O_678,N_9970,N_9981);
nor UO_679 (O_679,N_9973,N_9901);
nor UO_680 (O_680,N_9986,N_9969);
nand UO_681 (O_681,N_9997,N_9944);
nor UO_682 (O_682,N_9971,N_9979);
or UO_683 (O_683,N_9948,N_9917);
xnor UO_684 (O_684,N_9995,N_9969);
nor UO_685 (O_685,N_9977,N_9970);
or UO_686 (O_686,N_9989,N_9999);
nor UO_687 (O_687,N_9980,N_9990);
and UO_688 (O_688,N_9914,N_9924);
nor UO_689 (O_689,N_9966,N_9916);
or UO_690 (O_690,N_9981,N_9923);
and UO_691 (O_691,N_9918,N_9932);
xor UO_692 (O_692,N_9906,N_9916);
nor UO_693 (O_693,N_9927,N_9914);
nand UO_694 (O_694,N_9900,N_9953);
or UO_695 (O_695,N_9972,N_9946);
nor UO_696 (O_696,N_9950,N_9983);
nor UO_697 (O_697,N_9926,N_9954);
or UO_698 (O_698,N_9953,N_9916);
and UO_699 (O_699,N_9925,N_9945);
and UO_700 (O_700,N_9942,N_9934);
nor UO_701 (O_701,N_9965,N_9920);
or UO_702 (O_702,N_9960,N_9979);
or UO_703 (O_703,N_9991,N_9953);
nand UO_704 (O_704,N_9965,N_9938);
or UO_705 (O_705,N_9928,N_9996);
nand UO_706 (O_706,N_9926,N_9965);
or UO_707 (O_707,N_9907,N_9913);
nand UO_708 (O_708,N_9934,N_9981);
nand UO_709 (O_709,N_9945,N_9972);
nor UO_710 (O_710,N_9946,N_9984);
xnor UO_711 (O_711,N_9910,N_9972);
xnor UO_712 (O_712,N_9999,N_9933);
nand UO_713 (O_713,N_9932,N_9900);
and UO_714 (O_714,N_9987,N_9903);
or UO_715 (O_715,N_9922,N_9991);
or UO_716 (O_716,N_9910,N_9900);
nor UO_717 (O_717,N_9989,N_9971);
nand UO_718 (O_718,N_9989,N_9995);
nor UO_719 (O_719,N_9997,N_9975);
and UO_720 (O_720,N_9901,N_9902);
or UO_721 (O_721,N_9919,N_9941);
xor UO_722 (O_722,N_9918,N_9922);
nor UO_723 (O_723,N_9916,N_9970);
and UO_724 (O_724,N_9912,N_9925);
or UO_725 (O_725,N_9967,N_9931);
xor UO_726 (O_726,N_9916,N_9945);
xor UO_727 (O_727,N_9947,N_9922);
or UO_728 (O_728,N_9988,N_9954);
nand UO_729 (O_729,N_9921,N_9962);
or UO_730 (O_730,N_9999,N_9993);
and UO_731 (O_731,N_9974,N_9931);
or UO_732 (O_732,N_9938,N_9913);
or UO_733 (O_733,N_9955,N_9940);
and UO_734 (O_734,N_9938,N_9907);
and UO_735 (O_735,N_9941,N_9971);
and UO_736 (O_736,N_9955,N_9932);
or UO_737 (O_737,N_9904,N_9925);
and UO_738 (O_738,N_9973,N_9927);
or UO_739 (O_739,N_9975,N_9927);
nor UO_740 (O_740,N_9970,N_9914);
or UO_741 (O_741,N_9979,N_9993);
xnor UO_742 (O_742,N_9948,N_9944);
and UO_743 (O_743,N_9986,N_9918);
or UO_744 (O_744,N_9934,N_9903);
and UO_745 (O_745,N_9998,N_9926);
xnor UO_746 (O_746,N_9909,N_9966);
xnor UO_747 (O_747,N_9928,N_9909);
nand UO_748 (O_748,N_9938,N_9919);
xnor UO_749 (O_749,N_9986,N_9990);
or UO_750 (O_750,N_9992,N_9949);
xor UO_751 (O_751,N_9984,N_9995);
or UO_752 (O_752,N_9916,N_9942);
and UO_753 (O_753,N_9915,N_9954);
or UO_754 (O_754,N_9946,N_9980);
xnor UO_755 (O_755,N_9953,N_9994);
nand UO_756 (O_756,N_9942,N_9996);
nor UO_757 (O_757,N_9934,N_9920);
or UO_758 (O_758,N_9907,N_9937);
or UO_759 (O_759,N_9950,N_9903);
nor UO_760 (O_760,N_9926,N_9947);
and UO_761 (O_761,N_9937,N_9951);
nor UO_762 (O_762,N_9957,N_9928);
xnor UO_763 (O_763,N_9923,N_9973);
nor UO_764 (O_764,N_9999,N_9940);
xnor UO_765 (O_765,N_9920,N_9904);
nand UO_766 (O_766,N_9993,N_9918);
or UO_767 (O_767,N_9991,N_9929);
xor UO_768 (O_768,N_9927,N_9968);
and UO_769 (O_769,N_9980,N_9938);
or UO_770 (O_770,N_9958,N_9969);
or UO_771 (O_771,N_9986,N_9926);
nor UO_772 (O_772,N_9945,N_9947);
nor UO_773 (O_773,N_9910,N_9999);
nand UO_774 (O_774,N_9998,N_9972);
or UO_775 (O_775,N_9956,N_9992);
xnor UO_776 (O_776,N_9988,N_9989);
xor UO_777 (O_777,N_9982,N_9959);
xor UO_778 (O_778,N_9936,N_9961);
or UO_779 (O_779,N_9918,N_9980);
nor UO_780 (O_780,N_9914,N_9906);
nor UO_781 (O_781,N_9903,N_9971);
and UO_782 (O_782,N_9917,N_9998);
xnor UO_783 (O_783,N_9914,N_9986);
xor UO_784 (O_784,N_9912,N_9962);
nand UO_785 (O_785,N_9938,N_9923);
nor UO_786 (O_786,N_9916,N_9900);
nand UO_787 (O_787,N_9908,N_9997);
or UO_788 (O_788,N_9987,N_9998);
nor UO_789 (O_789,N_9972,N_9935);
nor UO_790 (O_790,N_9906,N_9934);
or UO_791 (O_791,N_9922,N_9949);
or UO_792 (O_792,N_9909,N_9908);
xor UO_793 (O_793,N_9982,N_9913);
or UO_794 (O_794,N_9968,N_9978);
xnor UO_795 (O_795,N_9915,N_9932);
xnor UO_796 (O_796,N_9990,N_9926);
nor UO_797 (O_797,N_9963,N_9996);
and UO_798 (O_798,N_9991,N_9927);
and UO_799 (O_799,N_9951,N_9981);
xor UO_800 (O_800,N_9953,N_9905);
or UO_801 (O_801,N_9913,N_9944);
xnor UO_802 (O_802,N_9960,N_9943);
xnor UO_803 (O_803,N_9916,N_9926);
xnor UO_804 (O_804,N_9919,N_9961);
and UO_805 (O_805,N_9931,N_9963);
xor UO_806 (O_806,N_9922,N_9934);
nor UO_807 (O_807,N_9911,N_9949);
xor UO_808 (O_808,N_9947,N_9988);
and UO_809 (O_809,N_9961,N_9925);
nand UO_810 (O_810,N_9924,N_9953);
and UO_811 (O_811,N_9909,N_9930);
or UO_812 (O_812,N_9912,N_9949);
and UO_813 (O_813,N_9987,N_9919);
or UO_814 (O_814,N_9977,N_9914);
xor UO_815 (O_815,N_9958,N_9918);
and UO_816 (O_816,N_9989,N_9903);
nand UO_817 (O_817,N_9987,N_9906);
or UO_818 (O_818,N_9953,N_9946);
xor UO_819 (O_819,N_9904,N_9975);
and UO_820 (O_820,N_9965,N_9928);
or UO_821 (O_821,N_9985,N_9959);
nor UO_822 (O_822,N_9955,N_9912);
and UO_823 (O_823,N_9943,N_9913);
or UO_824 (O_824,N_9994,N_9948);
or UO_825 (O_825,N_9997,N_9951);
and UO_826 (O_826,N_9997,N_9999);
and UO_827 (O_827,N_9901,N_9934);
nand UO_828 (O_828,N_9965,N_9963);
or UO_829 (O_829,N_9912,N_9957);
nor UO_830 (O_830,N_9964,N_9998);
or UO_831 (O_831,N_9929,N_9987);
or UO_832 (O_832,N_9967,N_9901);
or UO_833 (O_833,N_9943,N_9952);
or UO_834 (O_834,N_9925,N_9963);
or UO_835 (O_835,N_9935,N_9962);
nor UO_836 (O_836,N_9960,N_9996);
or UO_837 (O_837,N_9914,N_9990);
xnor UO_838 (O_838,N_9937,N_9933);
and UO_839 (O_839,N_9927,N_9932);
and UO_840 (O_840,N_9903,N_9973);
or UO_841 (O_841,N_9986,N_9930);
nand UO_842 (O_842,N_9971,N_9936);
xnor UO_843 (O_843,N_9921,N_9967);
or UO_844 (O_844,N_9907,N_9986);
or UO_845 (O_845,N_9946,N_9904);
nand UO_846 (O_846,N_9953,N_9926);
xor UO_847 (O_847,N_9970,N_9996);
or UO_848 (O_848,N_9996,N_9924);
nor UO_849 (O_849,N_9923,N_9996);
and UO_850 (O_850,N_9933,N_9923);
xor UO_851 (O_851,N_9917,N_9903);
xnor UO_852 (O_852,N_9910,N_9920);
or UO_853 (O_853,N_9908,N_9939);
nor UO_854 (O_854,N_9987,N_9934);
nor UO_855 (O_855,N_9981,N_9976);
xor UO_856 (O_856,N_9901,N_9919);
and UO_857 (O_857,N_9923,N_9929);
or UO_858 (O_858,N_9975,N_9974);
nor UO_859 (O_859,N_9940,N_9909);
or UO_860 (O_860,N_9965,N_9911);
nor UO_861 (O_861,N_9999,N_9985);
xor UO_862 (O_862,N_9992,N_9973);
xor UO_863 (O_863,N_9982,N_9996);
nor UO_864 (O_864,N_9995,N_9991);
nor UO_865 (O_865,N_9907,N_9941);
or UO_866 (O_866,N_9997,N_9936);
or UO_867 (O_867,N_9991,N_9963);
xor UO_868 (O_868,N_9999,N_9953);
nand UO_869 (O_869,N_9917,N_9996);
or UO_870 (O_870,N_9943,N_9956);
or UO_871 (O_871,N_9977,N_9997);
and UO_872 (O_872,N_9919,N_9978);
and UO_873 (O_873,N_9919,N_9962);
xnor UO_874 (O_874,N_9943,N_9989);
nor UO_875 (O_875,N_9912,N_9974);
or UO_876 (O_876,N_9976,N_9907);
nand UO_877 (O_877,N_9994,N_9949);
or UO_878 (O_878,N_9970,N_9942);
and UO_879 (O_879,N_9986,N_9964);
xor UO_880 (O_880,N_9932,N_9961);
nand UO_881 (O_881,N_9964,N_9990);
or UO_882 (O_882,N_9949,N_9991);
xor UO_883 (O_883,N_9923,N_9999);
or UO_884 (O_884,N_9945,N_9924);
nand UO_885 (O_885,N_9956,N_9910);
nor UO_886 (O_886,N_9915,N_9935);
nand UO_887 (O_887,N_9964,N_9985);
nand UO_888 (O_888,N_9908,N_9969);
and UO_889 (O_889,N_9952,N_9927);
and UO_890 (O_890,N_9996,N_9908);
nand UO_891 (O_891,N_9939,N_9959);
nor UO_892 (O_892,N_9934,N_9983);
xnor UO_893 (O_893,N_9954,N_9937);
nor UO_894 (O_894,N_9934,N_9924);
and UO_895 (O_895,N_9917,N_9992);
nand UO_896 (O_896,N_9921,N_9990);
or UO_897 (O_897,N_9960,N_9936);
nand UO_898 (O_898,N_9934,N_9969);
or UO_899 (O_899,N_9915,N_9933);
and UO_900 (O_900,N_9907,N_9981);
xor UO_901 (O_901,N_9962,N_9948);
nand UO_902 (O_902,N_9945,N_9909);
or UO_903 (O_903,N_9950,N_9916);
nand UO_904 (O_904,N_9931,N_9905);
and UO_905 (O_905,N_9974,N_9997);
nand UO_906 (O_906,N_9923,N_9961);
and UO_907 (O_907,N_9919,N_9972);
nor UO_908 (O_908,N_9962,N_9951);
and UO_909 (O_909,N_9966,N_9962);
nor UO_910 (O_910,N_9969,N_9909);
xor UO_911 (O_911,N_9991,N_9976);
nor UO_912 (O_912,N_9998,N_9942);
and UO_913 (O_913,N_9941,N_9916);
and UO_914 (O_914,N_9924,N_9984);
nor UO_915 (O_915,N_9975,N_9914);
or UO_916 (O_916,N_9910,N_9937);
nand UO_917 (O_917,N_9912,N_9930);
and UO_918 (O_918,N_9917,N_9916);
nor UO_919 (O_919,N_9947,N_9944);
nor UO_920 (O_920,N_9940,N_9957);
or UO_921 (O_921,N_9939,N_9986);
nor UO_922 (O_922,N_9917,N_9982);
or UO_923 (O_923,N_9955,N_9982);
and UO_924 (O_924,N_9918,N_9915);
nand UO_925 (O_925,N_9997,N_9947);
xor UO_926 (O_926,N_9948,N_9975);
and UO_927 (O_927,N_9913,N_9985);
xor UO_928 (O_928,N_9969,N_9992);
nand UO_929 (O_929,N_9979,N_9922);
nor UO_930 (O_930,N_9949,N_9996);
and UO_931 (O_931,N_9900,N_9978);
or UO_932 (O_932,N_9938,N_9926);
or UO_933 (O_933,N_9932,N_9971);
nor UO_934 (O_934,N_9909,N_9991);
or UO_935 (O_935,N_9906,N_9980);
or UO_936 (O_936,N_9995,N_9983);
or UO_937 (O_937,N_9917,N_9928);
xnor UO_938 (O_938,N_9905,N_9973);
and UO_939 (O_939,N_9938,N_9976);
and UO_940 (O_940,N_9985,N_9939);
or UO_941 (O_941,N_9908,N_9972);
nand UO_942 (O_942,N_9923,N_9972);
xnor UO_943 (O_943,N_9913,N_9995);
or UO_944 (O_944,N_9932,N_9998);
and UO_945 (O_945,N_9940,N_9956);
or UO_946 (O_946,N_9917,N_9988);
nor UO_947 (O_947,N_9991,N_9902);
or UO_948 (O_948,N_9959,N_9917);
or UO_949 (O_949,N_9998,N_9948);
and UO_950 (O_950,N_9907,N_9947);
nor UO_951 (O_951,N_9999,N_9971);
and UO_952 (O_952,N_9963,N_9981);
and UO_953 (O_953,N_9978,N_9924);
or UO_954 (O_954,N_9908,N_9993);
nand UO_955 (O_955,N_9913,N_9970);
xor UO_956 (O_956,N_9991,N_9999);
xor UO_957 (O_957,N_9918,N_9953);
or UO_958 (O_958,N_9924,N_9985);
nor UO_959 (O_959,N_9949,N_9947);
nor UO_960 (O_960,N_9973,N_9991);
nor UO_961 (O_961,N_9921,N_9927);
xnor UO_962 (O_962,N_9915,N_9937);
nand UO_963 (O_963,N_9902,N_9989);
xnor UO_964 (O_964,N_9982,N_9923);
and UO_965 (O_965,N_9901,N_9992);
and UO_966 (O_966,N_9974,N_9977);
nor UO_967 (O_967,N_9954,N_9975);
and UO_968 (O_968,N_9980,N_9997);
nand UO_969 (O_969,N_9966,N_9900);
or UO_970 (O_970,N_9910,N_9977);
nor UO_971 (O_971,N_9945,N_9935);
nor UO_972 (O_972,N_9933,N_9948);
xnor UO_973 (O_973,N_9956,N_9916);
and UO_974 (O_974,N_9982,N_9916);
or UO_975 (O_975,N_9990,N_9999);
nand UO_976 (O_976,N_9982,N_9905);
xnor UO_977 (O_977,N_9910,N_9918);
xnor UO_978 (O_978,N_9958,N_9979);
and UO_979 (O_979,N_9936,N_9922);
or UO_980 (O_980,N_9934,N_9950);
xor UO_981 (O_981,N_9989,N_9955);
nand UO_982 (O_982,N_9924,N_9900);
or UO_983 (O_983,N_9937,N_9981);
xnor UO_984 (O_984,N_9974,N_9965);
nor UO_985 (O_985,N_9970,N_9971);
xor UO_986 (O_986,N_9909,N_9948);
and UO_987 (O_987,N_9941,N_9976);
or UO_988 (O_988,N_9938,N_9997);
or UO_989 (O_989,N_9946,N_9977);
nor UO_990 (O_990,N_9999,N_9977);
xnor UO_991 (O_991,N_9928,N_9970);
and UO_992 (O_992,N_9931,N_9949);
nor UO_993 (O_993,N_9976,N_9982);
nor UO_994 (O_994,N_9902,N_9959);
and UO_995 (O_995,N_9925,N_9959);
and UO_996 (O_996,N_9909,N_9905);
or UO_997 (O_997,N_9948,N_9919);
xnor UO_998 (O_998,N_9928,N_9995);
nor UO_999 (O_999,N_9981,N_9924);
or UO_1000 (O_1000,N_9910,N_9997);
nand UO_1001 (O_1001,N_9933,N_9949);
nor UO_1002 (O_1002,N_9985,N_9982);
xor UO_1003 (O_1003,N_9991,N_9984);
or UO_1004 (O_1004,N_9906,N_9978);
nor UO_1005 (O_1005,N_9939,N_9954);
xnor UO_1006 (O_1006,N_9904,N_9948);
nand UO_1007 (O_1007,N_9900,N_9906);
nor UO_1008 (O_1008,N_9995,N_9968);
nor UO_1009 (O_1009,N_9968,N_9979);
nor UO_1010 (O_1010,N_9959,N_9923);
nor UO_1011 (O_1011,N_9951,N_9900);
and UO_1012 (O_1012,N_9918,N_9940);
or UO_1013 (O_1013,N_9993,N_9944);
and UO_1014 (O_1014,N_9947,N_9921);
xnor UO_1015 (O_1015,N_9967,N_9986);
nor UO_1016 (O_1016,N_9926,N_9970);
nor UO_1017 (O_1017,N_9962,N_9977);
xnor UO_1018 (O_1018,N_9981,N_9992);
xnor UO_1019 (O_1019,N_9917,N_9940);
nor UO_1020 (O_1020,N_9994,N_9984);
or UO_1021 (O_1021,N_9999,N_9965);
xnor UO_1022 (O_1022,N_9948,N_9913);
nor UO_1023 (O_1023,N_9961,N_9969);
or UO_1024 (O_1024,N_9907,N_9934);
xnor UO_1025 (O_1025,N_9943,N_9935);
or UO_1026 (O_1026,N_9982,N_9946);
or UO_1027 (O_1027,N_9974,N_9989);
nand UO_1028 (O_1028,N_9925,N_9913);
xor UO_1029 (O_1029,N_9977,N_9927);
xor UO_1030 (O_1030,N_9945,N_9953);
and UO_1031 (O_1031,N_9977,N_9911);
nor UO_1032 (O_1032,N_9999,N_9982);
nor UO_1033 (O_1033,N_9992,N_9985);
or UO_1034 (O_1034,N_9976,N_9964);
and UO_1035 (O_1035,N_9939,N_9907);
or UO_1036 (O_1036,N_9901,N_9918);
nand UO_1037 (O_1037,N_9929,N_9937);
nand UO_1038 (O_1038,N_9947,N_9957);
xor UO_1039 (O_1039,N_9989,N_9934);
or UO_1040 (O_1040,N_9950,N_9953);
or UO_1041 (O_1041,N_9960,N_9952);
nand UO_1042 (O_1042,N_9929,N_9916);
or UO_1043 (O_1043,N_9929,N_9922);
nor UO_1044 (O_1044,N_9970,N_9999);
and UO_1045 (O_1045,N_9928,N_9999);
xor UO_1046 (O_1046,N_9987,N_9901);
xnor UO_1047 (O_1047,N_9906,N_9988);
nor UO_1048 (O_1048,N_9962,N_9987);
nor UO_1049 (O_1049,N_9988,N_9927);
xnor UO_1050 (O_1050,N_9959,N_9915);
and UO_1051 (O_1051,N_9940,N_9988);
and UO_1052 (O_1052,N_9945,N_9975);
nand UO_1053 (O_1053,N_9909,N_9918);
nor UO_1054 (O_1054,N_9975,N_9929);
or UO_1055 (O_1055,N_9997,N_9914);
and UO_1056 (O_1056,N_9905,N_9943);
nand UO_1057 (O_1057,N_9955,N_9904);
nor UO_1058 (O_1058,N_9967,N_9998);
and UO_1059 (O_1059,N_9909,N_9996);
nand UO_1060 (O_1060,N_9926,N_9971);
and UO_1061 (O_1061,N_9950,N_9938);
nor UO_1062 (O_1062,N_9939,N_9976);
and UO_1063 (O_1063,N_9998,N_9951);
nand UO_1064 (O_1064,N_9920,N_9975);
xor UO_1065 (O_1065,N_9934,N_9976);
nor UO_1066 (O_1066,N_9968,N_9902);
nand UO_1067 (O_1067,N_9923,N_9942);
nand UO_1068 (O_1068,N_9915,N_9910);
and UO_1069 (O_1069,N_9940,N_9981);
nand UO_1070 (O_1070,N_9921,N_9928);
nand UO_1071 (O_1071,N_9926,N_9976);
and UO_1072 (O_1072,N_9929,N_9933);
xnor UO_1073 (O_1073,N_9926,N_9920);
nand UO_1074 (O_1074,N_9990,N_9938);
nand UO_1075 (O_1075,N_9953,N_9979);
xnor UO_1076 (O_1076,N_9974,N_9904);
or UO_1077 (O_1077,N_9944,N_9950);
nor UO_1078 (O_1078,N_9938,N_9971);
nor UO_1079 (O_1079,N_9962,N_9904);
nand UO_1080 (O_1080,N_9924,N_9931);
xor UO_1081 (O_1081,N_9901,N_9907);
xor UO_1082 (O_1082,N_9908,N_9990);
xnor UO_1083 (O_1083,N_9951,N_9910);
xnor UO_1084 (O_1084,N_9952,N_9916);
xor UO_1085 (O_1085,N_9993,N_9922);
and UO_1086 (O_1086,N_9952,N_9978);
nor UO_1087 (O_1087,N_9986,N_9934);
xnor UO_1088 (O_1088,N_9983,N_9976);
or UO_1089 (O_1089,N_9945,N_9988);
or UO_1090 (O_1090,N_9929,N_9921);
nand UO_1091 (O_1091,N_9908,N_9920);
nand UO_1092 (O_1092,N_9918,N_9970);
and UO_1093 (O_1093,N_9963,N_9902);
or UO_1094 (O_1094,N_9940,N_9936);
xnor UO_1095 (O_1095,N_9966,N_9928);
and UO_1096 (O_1096,N_9935,N_9926);
nand UO_1097 (O_1097,N_9961,N_9911);
xor UO_1098 (O_1098,N_9975,N_9931);
and UO_1099 (O_1099,N_9916,N_9915);
or UO_1100 (O_1100,N_9973,N_9989);
xnor UO_1101 (O_1101,N_9904,N_9933);
xnor UO_1102 (O_1102,N_9912,N_9959);
and UO_1103 (O_1103,N_9960,N_9990);
and UO_1104 (O_1104,N_9993,N_9909);
nand UO_1105 (O_1105,N_9956,N_9966);
nand UO_1106 (O_1106,N_9973,N_9955);
nand UO_1107 (O_1107,N_9968,N_9953);
nor UO_1108 (O_1108,N_9980,N_9922);
nand UO_1109 (O_1109,N_9922,N_9944);
nand UO_1110 (O_1110,N_9901,N_9959);
nand UO_1111 (O_1111,N_9962,N_9997);
or UO_1112 (O_1112,N_9976,N_9954);
nor UO_1113 (O_1113,N_9916,N_9976);
or UO_1114 (O_1114,N_9933,N_9951);
nand UO_1115 (O_1115,N_9968,N_9973);
xor UO_1116 (O_1116,N_9951,N_9983);
nand UO_1117 (O_1117,N_9949,N_9998);
nor UO_1118 (O_1118,N_9945,N_9964);
xor UO_1119 (O_1119,N_9989,N_9978);
and UO_1120 (O_1120,N_9980,N_9971);
and UO_1121 (O_1121,N_9980,N_9911);
and UO_1122 (O_1122,N_9982,N_9903);
nand UO_1123 (O_1123,N_9943,N_9909);
xor UO_1124 (O_1124,N_9987,N_9942);
or UO_1125 (O_1125,N_9938,N_9904);
and UO_1126 (O_1126,N_9974,N_9934);
and UO_1127 (O_1127,N_9912,N_9939);
nand UO_1128 (O_1128,N_9939,N_9923);
nand UO_1129 (O_1129,N_9933,N_9952);
nand UO_1130 (O_1130,N_9954,N_9986);
or UO_1131 (O_1131,N_9929,N_9980);
and UO_1132 (O_1132,N_9957,N_9946);
nand UO_1133 (O_1133,N_9960,N_9930);
nand UO_1134 (O_1134,N_9923,N_9956);
nand UO_1135 (O_1135,N_9999,N_9947);
xor UO_1136 (O_1136,N_9934,N_9911);
or UO_1137 (O_1137,N_9906,N_9983);
xnor UO_1138 (O_1138,N_9988,N_9913);
xor UO_1139 (O_1139,N_9905,N_9932);
and UO_1140 (O_1140,N_9942,N_9989);
and UO_1141 (O_1141,N_9918,N_9900);
and UO_1142 (O_1142,N_9950,N_9904);
nor UO_1143 (O_1143,N_9940,N_9983);
or UO_1144 (O_1144,N_9959,N_9995);
xnor UO_1145 (O_1145,N_9935,N_9956);
nand UO_1146 (O_1146,N_9990,N_9945);
nand UO_1147 (O_1147,N_9926,N_9983);
nand UO_1148 (O_1148,N_9977,N_9919);
or UO_1149 (O_1149,N_9993,N_9992);
and UO_1150 (O_1150,N_9953,N_9983);
and UO_1151 (O_1151,N_9942,N_9902);
or UO_1152 (O_1152,N_9913,N_9957);
xnor UO_1153 (O_1153,N_9933,N_9980);
nand UO_1154 (O_1154,N_9901,N_9927);
and UO_1155 (O_1155,N_9944,N_9991);
and UO_1156 (O_1156,N_9938,N_9918);
nand UO_1157 (O_1157,N_9936,N_9972);
nand UO_1158 (O_1158,N_9911,N_9947);
nand UO_1159 (O_1159,N_9970,N_9944);
or UO_1160 (O_1160,N_9961,N_9946);
xor UO_1161 (O_1161,N_9978,N_9988);
nor UO_1162 (O_1162,N_9981,N_9959);
nand UO_1163 (O_1163,N_9968,N_9909);
xor UO_1164 (O_1164,N_9975,N_9907);
xor UO_1165 (O_1165,N_9983,N_9962);
or UO_1166 (O_1166,N_9917,N_9987);
and UO_1167 (O_1167,N_9988,N_9938);
or UO_1168 (O_1168,N_9952,N_9993);
nor UO_1169 (O_1169,N_9906,N_9968);
xor UO_1170 (O_1170,N_9999,N_9967);
or UO_1171 (O_1171,N_9982,N_9918);
and UO_1172 (O_1172,N_9933,N_9971);
xor UO_1173 (O_1173,N_9909,N_9981);
and UO_1174 (O_1174,N_9907,N_9946);
and UO_1175 (O_1175,N_9919,N_9980);
xnor UO_1176 (O_1176,N_9916,N_9907);
nor UO_1177 (O_1177,N_9926,N_9978);
and UO_1178 (O_1178,N_9952,N_9935);
and UO_1179 (O_1179,N_9990,N_9956);
and UO_1180 (O_1180,N_9979,N_9977);
xnor UO_1181 (O_1181,N_9999,N_9914);
xor UO_1182 (O_1182,N_9933,N_9935);
xnor UO_1183 (O_1183,N_9925,N_9903);
xnor UO_1184 (O_1184,N_9989,N_9939);
and UO_1185 (O_1185,N_9950,N_9963);
nor UO_1186 (O_1186,N_9967,N_9978);
xnor UO_1187 (O_1187,N_9900,N_9991);
or UO_1188 (O_1188,N_9901,N_9916);
and UO_1189 (O_1189,N_9963,N_9976);
nand UO_1190 (O_1190,N_9981,N_9947);
xnor UO_1191 (O_1191,N_9984,N_9974);
xor UO_1192 (O_1192,N_9955,N_9970);
and UO_1193 (O_1193,N_9911,N_9996);
xor UO_1194 (O_1194,N_9947,N_9950);
and UO_1195 (O_1195,N_9982,N_9988);
or UO_1196 (O_1196,N_9919,N_9955);
xnor UO_1197 (O_1197,N_9900,N_9954);
and UO_1198 (O_1198,N_9967,N_9980);
nor UO_1199 (O_1199,N_9904,N_9977);
nor UO_1200 (O_1200,N_9926,N_9984);
xnor UO_1201 (O_1201,N_9988,N_9923);
nor UO_1202 (O_1202,N_9950,N_9933);
or UO_1203 (O_1203,N_9963,N_9943);
and UO_1204 (O_1204,N_9997,N_9990);
nand UO_1205 (O_1205,N_9940,N_9929);
nand UO_1206 (O_1206,N_9924,N_9919);
or UO_1207 (O_1207,N_9946,N_9947);
nand UO_1208 (O_1208,N_9982,N_9949);
xor UO_1209 (O_1209,N_9942,N_9924);
xnor UO_1210 (O_1210,N_9962,N_9988);
nand UO_1211 (O_1211,N_9966,N_9998);
and UO_1212 (O_1212,N_9948,N_9988);
or UO_1213 (O_1213,N_9987,N_9921);
or UO_1214 (O_1214,N_9979,N_9906);
nand UO_1215 (O_1215,N_9964,N_9929);
nand UO_1216 (O_1216,N_9948,N_9961);
and UO_1217 (O_1217,N_9998,N_9909);
nand UO_1218 (O_1218,N_9924,N_9973);
xor UO_1219 (O_1219,N_9919,N_9918);
xor UO_1220 (O_1220,N_9933,N_9966);
nand UO_1221 (O_1221,N_9972,N_9973);
nor UO_1222 (O_1222,N_9943,N_9988);
nand UO_1223 (O_1223,N_9948,N_9960);
nand UO_1224 (O_1224,N_9971,N_9998);
or UO_1225 (O_1225,N_9943,N_9986);
nand UO_1226 (O_1226,N_9950,N_9917);
or UO_1227 (O_1227,N_9911,N_9900);
nand UO_1228 (O_1228,N_9918,N_9946);
nand UO_1229 (O_1229,N_9920,N_9925);
or UO_1230 (O_1230,N_9961,N_9966);
nor UO_1231 (O_1231,N_9914,N_9912);
nand UO_1232 (O_1232,N_9938,N_9920);
xnor UO_1233 (O_1233,N_9947,N_9914);
and UO_1234 (O_1234,N_9928,N_9998);
and UO_1235 (O_1235,N_9968,N_9993);
xnor UO_1236 (O_1236,N_9969,N_9936);
xnor UO_1237 (O_1237,N_9982,N_9950);
nor UO_1238 (O_1238,N_9951,N_9964);
nor UO_1239 (O_1239,N_9976,N_9995);
nand UO_1240 (O_1240,N_9999,N_9949);
nor UO_1241 (O_1241,N_9948,N_9967);
and UO_1242 (O_1242,N_9964,N_9970);
nor UO_1243 (O_1243,N_9934,N_9935);
or UO_1244 (O_1244,N_9980,N_9954);
nand UO_1245 (O_1245,N_9939,N_9968);
nand UO_1246 (O_1246,N_9956,N_9998);
xnor UO_1247 (O_1247,N_9922,N_9975);
or UO_1248 (O_1248,N_9991,N_9934);
nand UO_1249 (O_1249,N_9984,N_9911);
or UO_1250 (O_1250,N_9934,N_9933);
nor UO_1251 (O_1251,N_9963,N_9952);
xnor UO_1252 (O_1252,N_9910,N_9953);
nand UO_1253 (O_1253,N_9903,N_9978);
nor UO_1254 (O_1254,N_9925,N_9908);
nor UO_1255 (O_1255,N_9901,N_9920);
nor UO_1256 (O_1256,N_9975,N_9985);
xnor UO_1257 (O_1257,N_9940,N_9996);
xor UO_1258 (O_1258,N_9942,N_9972);
nor UO_1259 (O_1259,N_9966,N_9952);
and UO_1260 (O_1260,N_9967,N_9912);
or UO_1261 (O_1261,N_9938,N_9910);
nand UO_1262 (O_1262,N_9948,N_9966);
or UO_1263 (O_1263,N_9945,N_9946);
nor UO_1264 (O_1264,N_9993,N_9958);
and UO_1265 (O_1265,N_9905,N_9972);
or UO_1266 (O_1266,N_9982,N_9962);
and UO_1267 (O_1267,N_9911,N_9908);
and UO_1268 (O_1268,N_9956,N_9903);
xnor UO_1269 (O_1269,N_9982,N_9980);
nor UO_1270 (O_1270,N_9988,N_9974);
or UO_1271 (O_1271,N_9935,N_9902);
nor UO_1272 (O_1272,N_9928,N_9927);
xor UO_1273 (O_1273,N_9900,N_9931);
or UO_1274 (O_1274,N_9931,N_9981);
or UO_1275 (O_1275,N_9992,N_9971);
or UO_1276 (O_1276,N_9979,N_9959);
nand UO_1277 (O_1277,N_9986,N_9976);
and UO_1278 (O_1278,N_9926,N_9966);
nand UO_1279 (O_1279,N_9989,N_9993);
and UO_1280 (O_1280,N_9966,N_9955);
nor UO_1281 (O_1281,N_9920,N_9915);
xnor UO_1282 (O_1282,N_9942,N_9994);
or UO_1283 (O_1283,N_9930,N_9935);
or UO_1284 (O_1284,N_9934,N_9909);
and UO_1285 (O_1285,N_9989,N_9921);
and UO_1286 (O_1286,N_9920,N_9950);
xor UO_1287 (O_1287,N_9946,N_9950);
nand UO_1288 (O_1288,N_9997,N_9915);
xnor UO_1289 (O_1289,N_9900,N_9960);
nand UO_1290 (O_1290,N_9990,N_9949);
and UO_1291 (O_1291,N_9971,N_9921);
and UO_1292 (O_1292,N_9930,N_9958);
nand UO_1293 (O_1293,N_9973,N_9906);
or UO_1294 (O_1294,N_9923,N_9993);
and UO_1295 (O_1295,N_9990,N_9903);
xor UO_1296 (O_1296,N_9902,N_9964);
xor UO_1297 (O_1297,N_9999,N_9941);
and UO_1298 (O_1298,N_9932,N_9996);
xor UO_1299 (O_1299,N_9912,N_9934);
nor UO_1300 (O_1300,N_9990,N_9954);
and UO_1301 (O_1301,N_9989,N_9926);
or UO_1302 (O_1302,N_9946,N_9985);
xor UO_1303 (O_1303,N_9951,N_9988);
or UO_1304 (O_1304,N_9976,N_9925);
or UO_1305 (O_1305,N_9978,N_9991);
nand UO_1306 (O_1306,N_9911,N_9928);
and UO_1307 (O_1307,N_9998,N_9927);
xor UO_1308 (O_1308,N_9912,N_9963);
nand UO_1309 (O_1309,N_9939,N_9937);
nand UO_1310 (O_1310,N_9930,N_9975);
or UO_1311 (O_1311,N_9942,N_9950);
or UO_1312 (O_1312,N_9997,N_9904);
and UO_1313 (O_1313,N_9968,N_9903);
nor UO_1314 (O_1314,N_9997,N_9922);
xnor UO_1315 (O_1315,N_9976,N_9945);
and UO_1316 (O_1316,N_9957,N_9958);
nor UO_1317 (O_1317,N_9976,N_9953);
or UO_1318 (O_1318,N_9946,N_9905);
nand UO_1319 (O_1319,N_9992,N_9958);
nor UO_1320 (O_1320,N_9907,N_9927);
nor UO_1321 (O_1321,N_9956,N_9974);
and UO_1322 (O_1322,N_9913,N_9967);
and UO_1323 (O_1323,N_9910,N_9958);
nand UO_1324 (O_1324,N_9970,N_9967);
nand UO_1325 (O_1325,N_9950,N_9958);
or UO_1326 (O_1326,N_9971,N_9909);
nand UO_1327 (O_1327,N_9928,N_9955);
xnor UO_1328 (O_1328,N_9910,N_9944);
xor UO_1329 (O_1329,N_9902,N_9977);
or UO_1330 (O_1330,N_9941,N_9920);
nor UO_1331 (O_1331,N_9987,N_9946);
and UO_1332 (O_1332,N_9906,N_9936);
or UO_1333 (O_1333,N_9944,N_9902);
and UO_1334 (O_1334,N_9957,N_9936);
nand UO_1335 (O_1335,N_9960,N_9958);
nor UO_1336 (O_1336,N_9919,N_9907);
nand UO_1337 (O_1337,N_9904,N_9937);
xnor UO_1338 (O_1338,N_9954,N_9994);
xnor UO_1339 (O_1339,N_9929,N_9942);
and UO_1340 (O_1340,N_9957,N_9983);
nand UO_1341 (O_1341,N_9907,N_9914);
nor UO_1342 (O_1342,N_9923,N_9979);
nand UO_1343 (O_1343,N_9962,N_9980);
or UO_1344 (O_1344,N_9916,N_9937);
nor UO_1345 (O_1345,N_9929,N_9904);
nor UO_1346 (O_1346,N_9973,N_9995);
xnor UO_1347 (O_1347,N_9916,N_9904);
nand UO_1348 (O_1348,N_9983,N_9937);
xor UO_1349 (O_1349,N_9935,N_9910);
nor UO_1350 (O_1350,N_9960,N_9947);
xnor UO_1351 (O_1351,N_9932,N_9976);
nand UO_1352 (O_1352,N_9911,N_9923);
nor UO_1353 (O_1353,N_9969,N_9943);
xnor UO_1354 (O_1354,N_9972,N_9947);
xor UO_1355 (O_1355,N_9936,N_9977);
and UO_1356 (O_1356,N_9912,N_9920);
nor UO_1357 (O_1357,N_9969,N_9950);
xor UO_1358 (O_1358,N_9951,N_9977);
xor UO_1359 (O_1359,N_9944,N_9912);
nor UO_1360 (O_1360,N_9921,N_9960);
nand UO_1361 (O_1361,N_9924,N_9918);
or UO_1362 (O_1362,N_9914,N_9958);
and UO_1363 (O_1363,N_9908,N_9932);
nand UO_1364 (O_1364,N_9928,N_9969);
nor UO_1365 (O_1365,N_9926,N_9930);
or UO_1366 (O_1366,N_9963,N_9929);
xnor UO_1367 (O_1367,N_9907,N_9971);
and UO_1368 (O_1368,N_9942,N_9919);
xor UO_1369 (O_1369,N_9936,N_9992);
nor UO_1370 (O_1370,N_9982,N_9927);
xor UO_1371 (O_1371,N_9917,N_9946);
xnor UO_1372 (O_1372,N_9941,N_9905);
and UO_1373 (O_1373,N_9923,N_9915);
or UO_1374 (O_1374,N_9921,N_9953);
nor UO_1375 (O_1375,N_9976,N_9985);
or UO_1376 (O_1376,N_9933,N_9921);
xor UO_1377 (O_1377,N_9911,N_9998);
or UO_1378 (O_1378,N_9934,N_9957);
and UO_1379 (O_1379,N_9911,N_9976);
and UO_1380 (O_1380,N_9964,N_9913);
nor UO_1381 (O_1381,N_9923,N_9921);
nor UO_1382 (O_1382,N_9939,N_9962);
and UO_1383 (O_1383,N_9967,N_9926);
or UO_1384 (O_1384,N_9917,N_9977);
nor UO_1385 (O_1385,N_9914,N_9994);
or UO_1386 (O_1386,N_9930,N_9969);
or UO_1387 (O_1387,N_9973,N_9980);
nor UO_1388 (O_1388,N_9975,N_9953);
or UO_1389 (O_1389,N_9906,N_9902);
nor UO_1390 (O_1390,N_9944,N_9985);
nor UO_1391 (O_1391,N_9951,N_9953);
and UO_1392 (O_1392,N_9939,N_9969);
or UO_1393 (O_1393,N_9930,N_9932);
nand UO_1394 (O_1394,N_9946,N_9983);
nor UO_1395 (O_1395,N_9936,N_9979);
nand UO_1396 (O_1396,N_9902,N_9917);
or UO_1397 (O_1397,N_9906,N_9999);
nand UO_1398 (O_1398,N_9967,N_9922);
nand UO_1399 (O_1399,N_9914,N_9995);
and UO_1400 (O_1400,N_9946,N_9934);
nor UO_1401 (O_1401,N_9949,N_9914);
nand UO_1402 (O_1402,N_9951,N_9986);
nand UO_1403 (O_1403,N_9937,N_9924);
xnor UO_1404 (O_1404,N_9975,N_9966);
and UO_1405 (O_1405,N_9923,N_9941);
and UO_1406 (O_1406,N_9985,N_9929);
xor UO_1407 (O_1407,N_9978,N_9913);
or UO_1408 (O_1408,N_9962,N_9914);
xor UO_1409 (O_1409,N_9974,N_9944);
nor UO_1410 (O_1410,N_9955,N_9994);
and UO_1411 (O_1411,N_9961,N_9980);
nor UO_1412 (O_1412,N_9919,N_9956);
nand UO_1413 (O_1413,N_9920,N_9999);
or UO_1414 (O_1414,N_9951,N_9957);
nor UO_1415 (O_1415,N_9956,N_9933);
nor UO_1416 (O_1416,N_9991,N_9928);
and UO_1417 (O_1417,N_9926,N_9918);
xor UO_1418 (O_1418,N_9952,N_9970);
nand UO_1419 (O_1419,N_9938,N_9969);
or UO_1420 (O_1420,N_9994,N_9997);
nand UO_1421 (O_1421,N_9962,N_9918);
xnor UO_1422 (O_1422,N_9990,N_9987);
nand UO_1423 (O_1423,N_9901,N_9960);
and UO_1424 (O_1424,N_9973,N_9959);
xnor UO_1425 (O_1425,N_9974,N_9990);
or UO_1426 (O_1426,N_9923,N_9903);
and UO_1427 (O_1427,N_9904,N_9989);
nor UO_1428 (O_1428,N_9976,N_9917);
nor UO_1429 (O_1429,N_9939,N_9930);
nor UO_1430 (O_1430,N_9959,N_9947);
or UO_1431 (O_1431,N_9955,N_9960);
or UO_1432 (O_1432,N_9908,N_9918);
and UO_1433 (O_1433,N_9909,N_9915);
xor UO_1434 (O_1434,N_9977,N_9916);
or UO_1435 (O_1435,N_9913,N_9934);
nor UO_1436 (O_1436,N_9905,N_9920);
xor UO_1437 (O_1437,N_9926,N_9960);
nand UO_1438 (O_1438,N_9962,N_9933);
xor UO_1439 (O_1439,N_9925,N_9968);
xnor UO_1440 (O_1440,N_9911,N_9978);
and UO_1441 (O_1441,N_9942,N_9931);
nor UO_1442 (O_1442,N_9906,N_9982);
and UO_1443 (O_1443,N_9921,N_9994);
xor UO_1444 (O_1444,N_9911,N_9971);
or UO_1445 (O_1445,N_9957,N_9970);
or UO_1446 (O_1446,N_9964,N_9927);
nor UO_1447 (O_1447,N_9935,N_9987);
xor UO_1448 (O_1448,N_9968,N_9916);
nor UO_1449 (O_1449,N_9938,N_9940);
or UO_1450 (O_1450,N_9983,N_9959);
xnor UO_1451 (O_1451,N_9990,N_9934);
and UO_1452 (O_1452,N_9997,N_9934);
nand UO_1453 (O_1453,N_9949,N_9970);
and UO_1454 (O_1454,N_9906,N_9937);
and UO_1455 (O_1455,N_9965,N_9944);
nand UO_1456 (O_1456,N_9979,N_9962);
nor UO_1457 (O_1457,N_9958,N_9906);
nand UO_1458 (O_1458,N_9972,N_9966);
and UO_1459 (O_1459,N_9921,N_9980);
xnor UO_1460 (O_1460,N_9917,N_9991);
and UO_1461 (O_1461,N_9960,N_9910);
nand UO_1462 (O_1462,N_9938,N_9921);
nand UO_1463 (O_1463,N_9901,N_9955);
nor UO_1464 (O_1464,N_9991,N_9960);
nor UO_1465 (O_1465,N_9963,N_9933);
xor UO_1466 (O_1466,N_9941,N_9975);
xnor UO_1467 (O_1467,N_9905,N_9987);
nor UO_1468 (O_1468,N_9949,N_9986);
nor UO_1469 (O_1469,N_9907,N_9949);
xor UO_1470 (O_1470,N_9940,N_9924);
xor UO_1471 (O_1471,N_9949,N_9997);
nand UO_1472 (O_1472,N_9936,N_9916);
or UO_1473 (O_1473,N_9918,N_9975);
and UO_1474 (O_1474,N_9907,N_9952);
nor UO_1475 (O_1475,N_9944,N_9914);
xnor UO_1476 (O_1476,N_9922,N_9935);
and UO_1477 (O_1477,N_9904,N_9952);
xor UO_1478 (O_1478,N_9965,N_9903);
xor UO_1479 (O_1479,N_9977,N_9964);
nor UO_1480 (O_1480,N_9955,N_9961);
nor UO_1481 (O_1481,N_9930,N_9943);
and UO_1482 (O_1482,N_9976,N_9950);
nand UO_1483 (O_1483,N_9959,N_9956);
xnor UO_1484 (O_1484,N_9968,N_9972);
nand UO_1485 (O_1485,N_9930,N_9981);
and UO_1486 (O_1486,N_9973,N_9982);
or UO_1487 (O_1487,N_9987,N_9939);
xnor UO_1488 (O_1488,N_9997,N_9988);
xnor UO_1489 (O_1489,N_9906,N_9928);
nand UO_1490 (O_1490,N_9957,N_9923);
nor UO_1491 (O_1491,N_9991,N_9958);
nand UO_1492 (O_1492,N_9985,N_9965);
nor UO_1493 (O_1493,N_9962,N_9946);
or UO_1494 (O_1494,N_9979,N_9984);
nand UO_1495 (O_1495,N_9980,N_9902);
nand UO_1496 (O_1496,N_9902,N_9995);
nand UO_1497 (O_1497,N_9952,N_9923);
nand UO_1498 (O_1498,N_9943,N_9995);
xnor UO_1499 (O_1499,N_9935,N_9959);
endmodule