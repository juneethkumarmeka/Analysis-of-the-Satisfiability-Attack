module basic_1000_10000_1500_2_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5003,N_5004,N_5005,N_5009,N_5011,N_5012,N_5015,N_5016,N_5017,N_5018,N_5021,N_5025,N_5026,N_5027,N_5028,N_5030,N_5031,N_5033,N_5034,N_5037,N_5038,N_5040,N_5043,N_5046,N_5047,N_5048,N_5051,N_5054,N_5056,N_5057,N_5060,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5074,N_5076,N_5077,N_5078,N_5081,N_5083,N_5084,N_5085,N_5086,N_5093,N_5094,N_5096,N_5097,N_5098,N_5100,N_5102,N_5107,N_5109,N_5110,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5120,N_5121,N_5122,N_5123,N_5126,N_5127,N_5128,N_5130,N_5132,N_5134,N_5137,N_5138,N_5142,N_5143,N_5145,N_5146,N_5147,N_5148,N_5149,N_5151,N_5153,N_5154,N_5156,N_5160,N_5161,N_5163,N_5164,N_5165,N_5168,N_5169,N_5170,N_5172,N_5173,N_5178,N_5179,N_5180,N_5181,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5192,N_5194,N_5195,N_5197,N_5198,N_5199,N_5201,N_5202,N_5209,N_5210,N_5211,N_5213,N_5217,N_5218,N_5221,N_5222,N_5223,N_5226,N_5227,N_5230,N_5231,N_5233,N_5234,N_5236,N_5240,N_5241,N_5243,N_5244,N_5248,N_5249,N_5251,N_5252,N_5253,N_5256,N_5257,N_5259,N_5260,N_5264,N_5265,N_5266,N_5268,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5278,N_5280,N_5281,N_5284,N_5286,N_5288,N_5290,N_5292,N_5293,N_5295,N_5296,N_5297,N_5299,N_5300,N_5303,N_5304,N_5307,N_5308,N_5309,N_5310,N_5312,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5323,N_5324,N_5326,N_5327,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5338,N_5339,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5361,N_5363,N_5365,N_5366,N_5367,N_5370,N_5371,N_5372,N_5375,N_5376,N_5378,N_5379,N_5383,N_5384,N_5385,N_5386,N_5388,N_5390,N_5391,N_5393,N_5395,N_5396,N_5397,N_5399,N_5400,N_5403,N_5404,N_5405,N_5406,N_5412,N_5413,N_5414,N_5415,N_5418,N_5419,N_5421,N_5422,N_5424,N_5427,N_5428,N_5430,N_5431,N_5432,N_5433,N_5434,N_5437,N_5440,N_5441,N_5443,N_5446,N_5447,N_5449,N_5450,N_5451,N_5452,N_5454,N_5457,N_5458,N_5459,N_5460,N_5461,N_5463,N_5464,N_5465,N_5466,N_5468,N_5469,N_5470,N_5473,N_5474,N_5475,N_5477,N_5483,N_5485,N_5486,N_5487,N_5489,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5502,N_5503,N_5504,N_5507,N_5508,N_5509,N_5511,N_5512,N_5515,N_5516,N_5519,N_5520,N_5521,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5533,N_5534,N_5538,N_5539,N_5544,N_5545,N_5546,N_5548,N_5549,N_5553,N_5557,N_5558,N_5560,N_5561,N_5564,N_5565,N_5566,N_5568,N_5569,N_5570,N_5572,N_5574,N_5575,N_5577,N_5579,N_5583,N_5584,N_5586,N_5587,N_5591,N_5594,N_5597,N_5598,N_5599,N_5600,N_5601,N_5603,N_5604,N_5605,N_5608,N_5609,N_5611,N_5612,N_5613,N_5614,N_5621,N_5622,N_5625,N_5627,N_5628,N_5629,N_5630,N_5633,N_5636,N_5639,N_5640,N_5641,N_5642,N_5644,N_5645,N_5649,N_5651,N_5652,N_5653,N_5654,N_5655,N_5660,N_5662,N_5664,N_5665,N_5666,N_5668,N_5669,N_5670,N_5671,N_5672,N_5674,N_5675,N_5676,N_5678,N_5680,N_5683,N_5684,N_5685,N_5686,N_5688,N_5690,N_5693,N_5694,N_5696,N_5697,N_5698,N_5700,N_5704,N_5705,N_5706,N_5708,N_5712,N_5713,N_5714,N_5716,N_5717,N_5718,N_5719,N_5721,N_5722,N_5724,N_5726,N_5727,N_5730,N_5732,N_5735,N_5736,N_5737,N_5739,N_5740,N_5741,N_5742,N_5745,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5755,N_5756,N_5757,N_5759,N_5760,N_5761,N_5765,N_5766,N_5767,N_5772,N_5773,N_5774,N_5775,N_5777,N_5779,N_5780,N_5782,N_5786,N_5787,N_5788,N_5790,N_5793,N_5796,N_5798,N_5799,N_5807,N_5812,N_5813,N_5815,N_5818,N_5820,N_5821,N_5822,N_5825,N_5828,N_5829,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5840,N_5841,N_5842,N_5843,N_5844,N_5846,N_5848,N_5851,N_5853,N_5854,N_5856,N_5857,N_5858,N_5861,N_5864,N_5865,N_5866,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5883,N_5884,N_5886,N_5887,N_5890,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5900,N_5902,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5920,N_5921,N_5922,N_5926,N_5927,N_5929,N_5933,N_5937,N_5938,N_5939,N_5940,N_5942,N_5943,N_5944,N_5946,N_5947,N_5948,N_5949,N_5950,N_5955,N_5956,N_5957,N_5961,N_5963,N_5964,N_5966,N_5967,N_5969,N_5970,N_5972,N_5973,N_5975,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5990,N_5991,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_6000,N_6003,N_6004,N_6008,N_6010,N_6011,N_6012,N_6015,N_6016,N_6017,N_6018,N_6020,N_6022,N_6029,N_6030,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6042,N_6043,N_6044,N_6045,N_6046,N_6048,N_6049,N_6050,N_6051,N_6054,N_6056,N_6057,N_6060,N_6062,N_6063,N_6066,N_6068,N_6069,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6081,N_6082,N_6086,N_6088,N_6090,N_6095,N_6096,N_6097,N_6099,N_6103,N_6105,N_6106,N_6108,N_6109,N_6115,N_6116,N_6117,N_6120,N_6122,N_6124,N_6125,N_6127,N_6128,N_6129,N_6135,N_6138,N_6139,N_6140,N_6141,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6151,N_6152,N_6153,N_6155,N_6160,N_6161,N_6162,N_6163,N_6164,N_6166,N_6167,N_6168,N_6169,N_6170,N_6173,N_6174,N_6175,N_6176,N_6177,N_6179,N_6180,N_6182,N_6185,N_6187,N_6190,N_6191,N_6194,N_6195,N_6197,N_6198,N_6200,N_6204,N_6206,N_6211,N_6212,N_6213,N_6216,N_6218,N_6219,N_6221,N_6223,N_6225,N_6226,N_6230,N_6231,N_6233,N_6234,N_6236,N_6237,N_6238,N_6241,N_6242,N_6243,N_6244,N_6246,N_6247,N_6248,N_6249,N_6251,N_6253,N_6254,N_6255,N_6256,N_6257,N_6261,N_6263,N_6266,N_6267,N_6268,N_6270,N_6272,N_6273,N_6275,N_6276,N_6278,N_6280,N_6281,N_6282,N_6283,N_6284,N_6287,N_6289,N_6292,N_6293,N_6294,N_6295,N_6296,N_6298,N_6299,N_6300,N_6301,N_6303,N_6304,N_6305,N_6306,N_6308,N_6309,N_6311,N_6312,N_6314,N_6315,N_6316,N_6321,N_6322,N_6324,N_6328,N_6330,N_6331,N_6332,N_6333,N_6334,N_6337,N_6339,N_6341,N_6344,N_6345,N_6346,N_6349,N_6350,N_6352,N_6353,N_6354,N_6355,N_6358,N_6359,N_6361,N_6364,N_6365,N_6366,N_6367,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6376,N_6378,N_6384,N_6385,N_6388,N_6389,N_6394,N_6395,N_6397,N_6400,N_6401,N_6402,N_6404,N_6405,N_6406,N_6407,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6418,N_6420,N_6422,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6432,N_6434,N_6437,N_6438,N_6443,N_6448,N_6451,N_6454,N_6456,N_6457,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6472,N_6473,N_6475,N_6482,N_6483,N_6484,N_6486,N_6487,N_6488,N_6490,N_6492,N_6493,N_6494,N_6495,N_6496,N_6498,N_6500,N_6502,N_6505,N_6506,N_6512,N_6515,N_6517,N_6519,N_6520,N_6521,N_6523,N_6524,N_6526,N_6531,N_6532,N_6535,N_6537,N_6538,N_6540,N_6542,N_6543,N_6548,N_6551,N_6555,N_6557,N_6558,N_6559,N_6560,N_6565,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6579,N_6580,N_6581,N_6583,N_6584,N_6587,N_6588,N_6591,N_6592,N_6593,N_6594,N_6595,N_6597,N_6598,N_6600,N_6601,N_6604,N_6606,N_6608,N_6612,N_6613,N_6620,N_6621,N_6622,N_6625,N_6627,N_6631,N_6632,N_6633,N_6635,N_6636,N_6637,N_6641,N_6644,N_6645,N_6646,N_6647,N_6648,N_6651,N_6652,N_6653,N_6658,N_6659,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6674,N_6675,N_6676,N_6680,N_6681,N_6683,N_6685,N_6686,N_6687,N_6689,N_6690,N_6692,N_6693,N_6694,N_6696,N_6697,N_6698,N_6699,N_6700,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6710,N_6713,N_6714,N_6716,N_6717,N_6720,N_6721,N_6722,N_6723,N_6725,N_6727,N_6728,N_6729,N_6730,N_6733,N_6734,N_6735,N_6737,N_6738,N_6743,N_6745,N_6748,N_6750,N_6751,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6760,N_6761,N_6762,N_6763,N_6765,N_6768,N_6770,N_6772,N_6774,N_6775,N_6779,N_6782,N_6785,N_6786,N_6787,N_6789,N_6791,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6808,N_6809,N_6812,N_6813,N_6816,N_6817,N_6822,N_6824,N_6825,N_6826,N_6827,N_6829,N_6830,N_6832,N_6834,N_6835,N_6836,N_6842,N_6845,N_6848,N_6849,N_6851,N_6852,N_6854,N_6857,N_6858,N_6859,N_6861,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6871,N_6873,N_6874,N_6876,N_6877,N_6878,N_6879,N_6880,N_6882,N_6883,N_6884,N_6885,N_6886,N_6888,N_6889,N_6892,N_6894,N_6896,N_6898,N_6899,N_6900,N_6902,N_6905,N_6907,N_6908,N_6909,N_6912,N_6913,N_6914,N_6915,N_6919,N_6920,N_6922,N_6925,N_6927,N_6928,N_6930,N_6936,N_6937,N_6938,N_6940,N_6942,N_6944,N_6946,N_6947,N_6949,N_6951,N_6953,N_6956,N_6957,N_6958,N_6961,N_6962,N_6963,N_6965,N_6966,N_6967,N_6969,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6980,N_6981,N_6983,N_6984,N_6985,N_6987,N_6988,N_6989,N_6993,N_6994,N_6996,N_6998,N_6999,N_7000,N_7001,N_7002,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7021,N_7023,N_7024,N_7027,N_7028,N_7029,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7039,N_7040,N_7044,N_7045,N_7047,N_7052,N_7053,N_7056,N_7057,N_7058,N_7059,N_7060,N_7062,N_7063,N_7065,N_7067,N_7070,N_7072,N_7076,N_7081,N_7084,N_7087,N_7092,N_7093,N_7095,N_7096,N_7097,N_7099,N_7100,N_7101,N_7103,N_7104,N_7105,N_7108,N_7109,N_7111,N_7114,N_7117,N_7118,N_7119,N_7120,N_7123,N_7126,N_7127,N_7128,N_7130,N_7131,N_7133,N_7134,N_7135,N_7137,N_7140,N_7141,N_7143,N_7147,N_7149,N_7151,N_7152,N_7154,N_7155,N_7157,N_7158,N_7159,N_7160,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7173,N_7174,N_7175,N_7177,N_7178,N_7181,N_7182,N_7183,N_7184,N_7187,N_7188,N_7191,N_7192,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7211,N_7212,N_7214,N_7215,N_7216,N_7218,N_7219,N_7220,N_7223,N_7225,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7245,N_7246,N_7248,N_7251,N_7252,N_7253,N_7256,N_7257,N_7258,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7268,N_7269,N_7271,N_7273,N_7280,N_7282,N_7284,N_7286,N_7288,N_7290,N_7292,N_7293,N_7295,N_7296,N_7297,N_7298,N_7301,N_7303,N_7304,N_7305,N_7306,N_7311,N_7312,N_7313,N_7314,N_7316,N_7321,N_7324,N_7325,N_7326,N_7327,N_7329,N_7331,N_7334,N_7335,N_7338,N_7340,N_7343,N_7344,N_7346,N_7347,N_7350,N_7353,N_7354,N_7355,N_7356,N_7357,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7377,N_7378,N_7380,N_7381,N_7382,N_7383,N_7387,N_7388,N_7391,N_7393,N_7394,N_7395,N_7396,N_7398,N_7399,N_7400,N_7403,N_7404,N_7408,N_7410,N_7411,N_7412,N_7413,N_7414,N_7416,N_7417,N_7418,N_7420,N_7421,N_7423,N_7425,N_7426,N_7427,N_7430,N_7431,N_7433,N_7434,N_7435,N_7437,N_7438,N_7439,N_7441,N_7442,N_7443,N_7444,N_7445,N_7447,N_7448,N_7452,N_7453,N_7454,N_7456,N_7457,N_7458,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7469,N_7470,N_7472,N_7474,N_7476,N_7478,N_7481,N_7482,N_7483,N_7485,N_7486,N_7487,N_7488,N_7492,N_7496,N_7497,N_7500,N_7501,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7513,N_7514,N_7515,N_7516,N_7517,N_7519,N_7521,N_7522,N_7523,N_7526,N_7527,N_7530,N_7531,N_7532,N_7534,N_7538,N_7539,N_7540,N_7543,N_7544,N_7545,N_7547,N_7548,N_7550,N_7551,N_7554,N_7555,N_7556,N_7557,N_7567,N_7568,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7580,N_7581,N_7582,N_7584,N_7585,N_7586,N_7590,N_7591,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7602,N_7604,N_7605,N_7606,N_7607,N_7608,N_7610,N_7612,N_7614,N_7615,N_7616,N_7618,N_7621,N_7623,N_7624,N_7625,N_7627,N_7628,N_7633,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7645,N_7647,N_7648,N_7650,N_7653,N_7658,N_7661,N_7664,N_7665,N_7667,N_7668,N_7669,N_7673,N_7674,N_7675,N_7677,N_7678,N_7679,N_7680,N_7683,N_7684,N_7685,N_7686,N_7688,N_7689,N_7690,N_7691,N_7693,N_7696,N_7698,N_7704,N_7705,N_7707,N_7709,N_7711,N_7712,N_7716,N_7717,N_7719,N_7726,N_7728,N_7729,N_7730,N_7731,N_7732,N_7734,N_7736,N_7738,N_7744,N_7745,N_7748,N_7749,N_7753,N_7755,N_7756,N_7758,N_7759,N_7763,N_7764,N_7766,N_7769,N_7771,N_7772,N_7773,N_7776,N_7777,N_7778,N_7781,N_7782,N_7783,N_7784,N_7786,N_7787,N_7788,N_7789,N_7791,N_7792,N_7793,N_7795,N_7800,N_7802,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7811,N_7812,N_7813,N_7814,N_7815,N_7817,N_7818,N_7819,N_7820,N_7830,N_7831,N_7832,N_7834,N_7836,N_7837,N_7839,N_7840,N_7842,N_7843,N_7844,N_7845,N_7847,N_7848,N_7850,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7864,N_7865,N_7867,N_7868,N_7869,N_7870,N_7872,N_7874,N_7876,N_7877,N_7880,N_7881,N_7882,N_7884,N_7888,N_7890,N_7893,N_7894,N_7895,N_7896,N_7898,N_7901,N_7903,N_7904,N_7905,N_7906,N_7907,N_7910,N_7912,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7924,N_7925,N_7926,N_7929,N_7933,N_7934,N_7936,N_7937,N_7938,N_7939,N_7943,N_7944,N_7945,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7956,N_7957,N_7960,N_7961,N_7962,N_7964,N_7965,N_7969,N_7970,N_7972,N_7973,N_7974,N_7976,N_7977,N_7978,N_7980,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7992,N_7993,N_7994,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8004,N_8005,N_8010,N_8014,N_8015,N_8017,N_8018,N_8019,N_8021,N_8022,N_8023,N_8024,N_8032,N_8033,N_8035,N_8037,N_8038,N_8039,N_8041,N_8043,N_8049,N_8051,N_8061,N_8062,N_8064,N_8065,N_8066,N_8067,N_8071,N_8072,N_8076,N_8078,N_8079,N_8081,N_8082,N_8083,N_8085,N_8086,N_8088,N_8090,N_8092,N_8093,N_8098,N_8101,N_8103,N_8107,N_8108,N_8109,N_8112,N_8113,N_8114,N_8115,N_8116,N_8118,N_8119,N_8120,N_8124,N_8126,N_8127,N_8128,N_8130,N_8131,N_8132,N_8133,N_8135,N_8136,N_8138,N_8141,N_8142,N_8143,N_8144,N_8145,N_8147,N_8148,N_8149,N_8150,N_8152,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8170,N_8171,N_8172,N_8173,N_8177,N_8178,N_8179,N_8181,N_8184,N_8186,N_8187,N_8188,N_8189,N_8190,N_8193,N_8194,N_8195,N_8197,N_8199,N_8200,N_8201,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8213,N_8214,N_8215,N_8223,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8238,N_8241,N_8242,N_8243,N_8245,N_8246,N_8247,N_8249,N_8252,N_8253,N_8257,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8276,N_8278,N_8280,N_8281,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8294,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8307,N_8308,N_8309,N_8311,N_8313,N_8315,N_8316,N_8317,N_8318,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8336,N_8338,N_8339,N_8342,N_8343,N_8344,N_8345,N_8351,N_8352,N_8353,N_8355,N_8357,N_8358,N_8359,N_8360,N_8370,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8380,N_8381,N_8383,N_8385,N_8387,N_8388,N_8389,N_8390,N_8391,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8401,N_8402,N_8403,N_8405,N_8406,N_8407,N_8410,N_8411,N_8413,N_8414,N_8415,N_8416,N_8418,N_8420,N_8421,N_8423,N_8424,N_8425,N_8428,N_8429,N_8431,N_8433,N_8435,N_8437,N_8439,N_8440,N_8442,N_8443,N_8444,N_8448,N_8449,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8458,N_8459,N_8462,N_8463,N_8464,N_8466,N_8467,N_8468,N_8469,N_8470,N_8472,N_8473,N_8474,N_8476,N_8477,N_8479,N_8480,N_8481,N_8482,N_8484,N_8485,N_8486,N_8487,N_8488,N_8490,N_8491,N_8492,N_8493,N_8495,N_8496,N_8497,N_8498,N_8499,N_8503,N_8504,N_8505,N_8508,N_8511,N_8515,N_8517,N_8518,N_8522,N_8524,N_8526,N_8529,N_8531,N_8532,N_8533,N_8534,N_8535,N_8539,N_8541,N_8542,N_8544,N_8545,N_8547,N_8549,N_8550,N_8552,N_8554,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8568,N_8569,N_8570,N_8571,N_8573,N_8574,N_8575,N_8576,N_8577,N_8579,N_8580,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8593,N_8594,N_8596,N_8597,N_8598,N_8600,N_8602,N_8603,N_8605,N_8606,N_8609,N_8610,N_8612,N_8613,N_8614,N_8615,N_8616,N_8618,N_8620,N_8621,N_8622,N_8623,N_8624,N_8626,N_8627,N_8628,N_8629,N_8632,N_8634,N_8636,N_8640,N_8641,N_8643,N_8644,N_8649,N_8650,N_8653,N_8656,N_8657,N_8660,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8672,N_8673,N_8674,N_8675,N_8677,N_8679,N_8680,N_8683,N_8684,N_8686,N_8687,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8697,N_8700,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8716,N_8719,N_8720,N_8721,N_8723,N_8724,N_8729,N_8732,N_8733,N_8734,N_8735,N_8736,N_8738,N_8739,N_8741,N_8743,N_8744,N_8745,N_8746,N_8748,N_8750,N_8751,N_8752,N_8753,N_8756,N_8759,N_8760,N_8762,N_8763,N_8765,N_8766,N_8768,N_8772,N_8775,N_8777,N_8778,N_8779,N_8780,N_8783,N_8786,N_8787,N_8791,N_8793,N_8794,N_8796,N_8800,N_8802,N_8805,N_8806,N_8807,N_8808,N_8810,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8820,N_8821,N_8824,N_8825,N_8826,N_8828,N_8830,N_8831,N_8832,N_8833,N_8834,N_8837,N_8838,N_8840,N_8842,N_8843,N_8844,N_8845,N_8846,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8858,N_8863,N_8864,N_8865,N_8871,N_8872,N_8875,N_8876,N_8877,N_8878,N_8880,N_8881,N_8882,N_8883,N_8886,N_8888,N_8891,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8902,N_8903,N_8909,N_8910,N_8911,N_8912,N_8914,N_8915,N_8917,N_8918,N_8920,N_8923,N_8924,N_8925,N_8926,N_8927,N_8929,N_8931,N_8933,N_8934,N_8935,N_8937,N_8938,N_8939,N_8943,N_8945,N_8946,N_8949,N_8951,N_8952,N_8953,N_8955,N_8957,N_8958,N_8960,N_8961,N_8962,N_8964,N_8965,N_8966,N_8968,N_8969,N_8970,N_8972,N_8974,N_8975,N_8976,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8992,N_8993,N_8995,N_8997,N_9002,N_9004,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9013,N_9014,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9023,N_9024,N_9025,N_9028,N_9029,N_9032,N_9033,N_9034,N_9035,N_9037,N_9038,N_9039,N_9040,N_9041,N_9043,N_9044,N_9046,N_9053,N_9054,N_9055,N_9058,N_9062,N_9063,N_9065,N_9067,N_9069,N_9073,N_9075,N_9076,N_9077,N_9078,N_9080,N_9081,N_9082,N_9083,N_9090,N_9092,N_9093,N_9094,N_9100,N_9101,N_9102,N_9103,N_9104,N_9106,N_9108,N_9110,N_9112,N_9115,N_9116,N_9117,N_9118,N_9121,N_9123,N_9124,N_9126,N_9127,N_9132,N_9133,N_9137,N_9138,N_9139,N_9140,N_9142,N_9143,N_9144,N_9145,N_9147,N_9149,N_9150,N_9153,N_9154,N_9155,N_9156,N_9157,N_9161,N_9162,N_9163,N_9164,N_9165,N_9167,N_9170,N_9173,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9185,N_9189,N_9190,N_9191,N_9193,N_9195,N_9198,N_9199,N_9200,N_9202,N_9204,N_9205,N_9207,N_9208,N_9209,N_9211,N_9213,N_9214,N_9216,N_9217,N_9218,N_9220,N_9222,N_9223,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9237,N_9239,N_9240,N_9241,N_9242,N_9245,N_9247,N_9250,N_9251,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9260,N_9264,N_9265,N_9266,N_9268,N_9269,N_9272,N_9273,N_9275,N_9276,N_9277,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9287,N_9288,N_9289,N_9290,N_9294,N_9296,N_9297,N_9298,N_9299,N_9302,N_9305,N_9306,N_9307,N_9308,N_9309,N_9311,N_9312,N_9318,N_9319,N_9321,N_9324,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9335,N_9337,N_9339,N_9342,N_9344,N_9345,N_9348,N_9350,N_9351,N_9352,N_9353,N_9354,N_9357,N_9358,N_9362,N_9363,N_9365,N_9368,N_9369,N_9371,N_9375,N_9377,N_9380,N_9383,N_9386,N_9387,N_9390,N_9392,N_9393,N_9394,N_9395,N_9396,N_9398,N_9399,N_9400,N_9402,N_9403,N_9404,N_9405,N_9407,N_9408,N_9410,N_9412,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9430,N_9432,N_9433,N_9434,N_9435,N_9437,N_9438,N_9440,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9449,N_9452,N_9454,N_9456,N_9457,N_9462,N_9463,N_9464,N_9465,N_9467,N_9468,N_9469,N_9472,N_9473,N_9474,N_9475,N_9478,N_9480,N_9481,N_9482,N_9483,N_9484,N_9486,N_9488,N_9489,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9507,N_9509,N_9511,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9523,N_9524,N_9526,N_9527,N_9530,N_9532,N_9533,N_9534,N_9537,N_9539,N_9541,N_9543,N_9546,N_9547,N_9553,N_9554,N_9555,N_9557,N_9560,N_9561,N_9563,N_9564,N_9565,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9580,N_9581,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9590,N_9591,N_9592,N_9594,N_9595,N_9598,N_9599,N_9600,N_9601,N_9604,N_9605,N_9607,N_9609,N_9612,N_9613,N_9614,N_9616,N_9618,N_9619,N_9620,N_9622,N_9624,N_9626,N_9627,N_9629,N_9630,N_9631,N_9635,N_9636,N_9638,N_9639,N_9641,N_9642,N_9643,N_9646,N_9650,N_9651,N_9654,N_9655,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9667,N_9670,N_9671,N_9672,N_9673,N_9675,N_9676,N_9679,N_9680,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9690,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9701,N_9702,N_9703,N_9705,N_9706,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9716,N_9717,N_9719,N_9720,N_9721,N_9723,N_9724,N_9726,N_9729,N_9730,N_9732,N_9734,N_9738,N_9739,N_9742,N_9744,N_9747,N_9748,N_9749,N_9753,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9764,N_9765,N_9766,N_9768,N_9769,N_9770,N_9771,N_9772,N_9774,N_9775,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9788,N_9792,N_9797,N_9801,N_9804,N_9807,N_9808,N_9809,N_9811,N_9812,N_9813,N_9815,N_9817,N_9818,N_9819,N_9821,N_9822,N_9827,N_9828,N_9829,N_9830,N_9832,N_9833,N_9837,N_9839,N_9840,N_9841,N_9843,N_9844,N_9847,N_9850,N_9852,N_9854,N_9856,N_9858,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9878,N_9880,N_9885,N_9887,N_9888,N_9889,N_9890,N_9892,N_9893,N_9894,N_9895,N_9898,N_9899,N_9900,N_9901,N_9902,N_9904,N_9907,N_9908,N_9910,N_9913,N_9916,N_9917,N_9918,N_9919,N_9921,N_9922,N_9923,N_9925,N_9926,N_9927,N_9928,N_9930,N_9932,N_9936,N_9938,N_9939,N_9940,N_9941,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9950,N_9952,N_9954,N_9956,N_9957,N_9963,N_9964,N_9968,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9977,N_9979,N_9980,N_9981,N_9984,N_9985,N_9988,N_9989,N_9990,N_9991,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_329,In_612);
nor U1 (N_1,In_143,In_847);
and U2 (N_2,In_253,In_732);
nand U3 (N_3,In_121,In_830);
and U4 (N_4,In_359,In_488);
nand U5 (N_5,In_13,In_567);
nor U6 (N_6,In_614,In_366);
nand U7 (N_7,In_991,In_970);
nand U8 (N_8,In_996,In_517);
xnor U9 (N_9,In_499,In_151);
nand U10 (N_10,In_465,In_459);
xnor U11 (N_11,In_32,In_495);
and U12 (N_12,In_355,In_518);
nor U13 (N_13,In_96,In_295);
or U14 (N_14,In_158,In_907);
and U15 (N_15,In_906,In_916);
and U16 (N_16,In_255,In_525);
or U17 (N_17,In_988,In_282);
or U18 (N_18,In_850,In_183);
nor U19 (N_19,In_526,In_56);
or U20 (N_20,In_442,In_912);
nor U21 (N_21,In_723,In_217);
and U22 (N_22,In_305,In_694);
xor U23 (N_23,In_936,In_507);
and U24 (N_24,In_64,In_709);
or U25 (N_25,In_628,In_589);
nor U26 (N_26,In_479,In_212);
and U27 (N_27,In_289,In_62);
nor U28 (N_28,In_86,In_326);
or U29 (N_29,In_123,In_740);
and U30 (N_30,In_215,In_801);
or U31 (N_31,In_481,In_873);
xor U32 (N_32,In_30,In_239);
nand U33 (N_33,In_568,In_776);
and U34 (N_34,In_361,In_337);
and U35 (N_35,In_486,In_680);
and U36 (N_36,In_487,In_927);
and U37 (N_37,In_642,In_266);
nand U38 (N_38,In_303,In_720);
nor U39 (N_39,In_10,In_50);
or U40 (N_40,In_840,In_675);
nand U41 (N_41,In_6,In_169);
and U42 (N_42,In_549,In_245);
xor U43 (N_43,In_216,In_322);
xor U44 (N_44,In_339,In_226);
xor U45 (N_45,In_102,In_108);
xnor U46 (N_46,In_650,In_800);
and U47 (N_47,In_336,In_707);
nand U48 (N_48,In_914,In_460);
and U49 (N_49,In_613,In_942);
nand U50 (N_50,In_957,In_979);
nor U51 (N_51,In_144,In_718);
nand U52 (N_52,In_861,In_691);
xor U53 (N_53,In_235,In_824);
or U54 (N_54,In_423,In_997);
nor U55 (N_55,In_351,In_389);
nor U56 (N_56,In_51,In_752);
or U57 (N_57,In_975,In_416);
or U58 (N_58,In_424,In_999);
xnor U59 (N_59,In_941,In_888);
and U60 (N_60,In_120,In_894);
and U61 (N_61,In_616,In_982);
and U62 (N_62,In_828,In_94);
nor U63 (N_63,In_803,In_107);
and U64 (N_64,In_441,In_280);
and U65 (N_65,In_952,In_190);
nor U66 (N_66,In_431,In_191);
nand U67 (N_67,In_265,In_584);
xor U68 (N_68,In_33,In_736);
and U69 (N_69,In_655,In_474);
nor U70 (N_70,In_370,In_529);
nand U71 (N_71,In_576,In_367);
xor U72 (N_72,In_247,In_885);
and U73 (N_73,In_382,In_268);
nand U74 (N_74,In_793,In_218);
nor U75 (N_75,In_357,In_348);
and U76 (N_76,In_381,In_500);
nand U77 (N_77,In_449,In_210);
and U78 (N_78,In_597,In_135);
nand U79 (N_79,In_19,In_409);
or U80 (N_80,In_739,In_106);
or U81 (N_81,In_882,In_260);
nand U82 (N_82,In_994,In_175);
nor U83 (N_83,In_114,In_512);
and U84 (N_84,In_977,In_903);
nor U85 (N_85,In_3,In_635);
xnor U86 (N_86,In_588,In_703);
xnor U87 (N_87,In_947,In_973);
and U88 (N_88,In_890,In_541);
nand U89 (N_89,In_412,In_674);
nor U90 (N_90,In_789,In_77);
nand U91 (N_91,In_437,In_570);
nand U92 (N_92,In_178,In_782);
nand U93 (N_93,In_700,In_572);
nand U94 (N_94,In_751,In_147);
nor U95 (N_95,In_42,In_76);
nand U96 (N_96,In_365,In_234);
nand U97 (N_97,In_791,In_261);
nand U98 (N_98,In_574,In_632);
nor U99 (N_99,In_626,In_594);
nand U100 (N_100,In_187,In_176);
and U101 (N_101,In_11,In_902);
nor U102 (N_102,In_561,In_75);
or U103 (N_103,In_236,In_754);
or U104 (N_104,In_884,In_786);
and U105 (N_105,In_331,In_358);
xnor U106 (N_106,In_644,In_457);
xnor U107 (N_107,In_761,In_814);
or U108 (N_108,In_730,In_137);
nor U109 (N_109,In_298,In_271);
nor U110 (N_110,In_922,In_772);
and U111 (N_111,In_250,In_596);
nor U112 (N_112,In_595,In_609);
and U113 (N_113,In_748,In_44);
nand U114 (N_114,In_390,In_400);
nand U115 (N_115,In_648,In_124);
and U116 (N_116,In_695,In_787);
nand U117 (N_117,In_606,In_946);
and U118 (N_118,In_540,In_634);
nand U119 (N_119,In_484,In_909);
nand U120 (N_120,In_434,In_910);
and U121 (N_121,In_471,In_12);
xnor U122 (N_122,In_100,In_607);
xnor U123 (N_123,In_164,In_931);
or U124 (N_124,In_535,In_360);
or U125 (N_125,In_981,In_649);
or U126 (N_126,In_189,In_654);
xor U127 (N_127,In_84,In_556);
xnor U128 (N_128,In_463,In_119);
and U129 (N_129,In_569,In_113);
nor U130 (N_130,In_395,In_625);
and U131 (N_131,In_797,In_118);
nand U132 (N_132,In_321,In_264);
and U133 (N_133,In_392,In_188);
or U134 (N_134,In_200,In_41);
nor U135 (N_135,In_919,In_69);
or U136 (N_136,In_901,In_523);
nand U137 (N_137,In_29,In_619);
and U138 (N_138,In_808,In_283);
nand U139 (N_139,In_811,In_429);
nand U140 (N_140,In_213,In_258);
xnor U141 (N_141,In_203,In_746);
or U142 (N_142,In_766,In_439);
xnor U143 (N_143,In_843,In_263);
nor U144 (N_144,In_886,In_599);
or U145 (N_145,In_445,In_324);
nor U146 (N_146,In_496,In_276);
nor U147 (N_147,In_172,In_640);
and U148 (N_148,In_727,In_246);
and U149 (N_149,In_834,In_984);
and U150 (N_150,In_611,In_109);
nor U151 (N_151,In_696,In_658);
and U152 (N_152,In_469,In_9);
or U153 (N_153,In_224,In_45);
nor U154 (N_154,In_364,In_586);
or U155 (N_155,In_697,In_4);
and U156 (N_156,In_908,In_548);
and U157 (N_157,In_878,In_664);
nand U158 (N_158,In_472,In_554);
nand U159 (N_159,In_145,In_539);
nand U160 (N_160,In_320,In_156);
nor U161 (N_161,In_799,In_140);
and U162 (N_162,In_598,In_284);
or U163 (N_163,In_874,In_287);
or U164 (N_164,In_252,In_842);
xor U165 (N_165,In_784,In_755);
and U166 (N_166,In_604,In_790);
nor U167 (N_167,In_775,In_180);
nor U168 (N_168,In_404,In_31);
xor U169 (N_169,In_722,In_573);
nor U170 (N_170,In_506,In_24);
nor U171 (N_171,In_756,In_951);
nor U172 (N_172,In_273,In_557);
or U173 (N_173,In_621,In_98);
or U174 (N_174,In_617,In_478);
nand U175 (N_175,In_115,In_49);
and U176 (N_176,In_848,In_600);
and U177 (N_177,In_489,In_763);
and U178 (N_178,In_1,In_37);
nor U179 (N_179,In_698,In_403);
nand U180 (N_180,In_527,In_862);
and U181 (N_181,In_867,In_352);
and U182 (N_182,In_921,In_998);
xnor U183 (N_183,In_724,In_181);
xor U184 (N_184,In_876,In_464);
nor U185 (N_185,In_513,In_945);
and U186 (N_186,In_950,In_670);
nor U187 (N_187,In_221,In_836);
nor U188 (N_188,In_310,In_306);
xnor U189 (N_189,In_79,In_232);
xor U190 (N_190,In_854,In_555);
and U191 (N_191,In_290,In_993);
nand U192 (N_192,In_543,In_810);
or U193 (N_193,In_323,In_293);
and U194 (N_194,In_207,In_451);
nor U195 (N_195,In_230,In_821);
and U196 (N_196,In_238,In_858);
or U197 (N_197,In_411,In_671);
or U198 (N_198,In_802,In_421);
or U199 (N_199,In_159,In_913);
nor U200 (N_200,In_661,In_22);
nand U201 (N_201,In_519,In_682);
nor U202 (N_202,In_122,In_815);
xnor U203 (N_203,In_627,In_297);
nor U204 (N_204,In_546,In_376);
nand U205 (N_205,In_482,In_769);
and U206 (N_206,In_925,In_373);
nor U207 (N_207,In_141,In_978);
nand U208 (N_208,In_804,In_388);
nand U209 (N_209,In_228,In_335);
nor U210 (N_210,In_167,In_537);
nand U211 (N_211,In_476,In_277);
nand U212 (N_212,In_562,In_798);
and U213 (N_213,In_443,In_980);
nor U214 (N_214,In_807,In_729);
nor U215 (N_215,In_87,In_129);
and U216 (N_216,In_413,In_39);
nor U217 (N_217,In_949,In_139);
nor U218 (N_218,In_14,In_349);
nand U219 (N_219,In_163,In_468);
and U220 (N_220,In_737,In_173);
nor U221 (N_221,In_338,In_54);
nor U222 (N_222,In_844,In_20);
or U223 (N_223,In_354,In_623);
or U224 (N_224,In_929,In_580);
nand U225 (N_225,In_877,In_485);
or U226 (N_226,In_656,In_48);
or U227 (N_227,In_397,In_958);
nand U228 (N_228,In_446,In_863);
nand U229 (N_229,In_651,In_544);
nand U230 (N_230,In_719,In_288);
nand U231 (N_231,In_347,In_933);
nand U232 (N_232,In_711,In_565);
and U233 (N_233,In_833,In_470);
xor U234 (N_234,In_768,In_944);
nor U235 (N_235,In_932,In_383);
or U236 (N_236,In_508,In_155);
nand U237 (N_237,In_179,In_918);
nand U238 (N_238,In_672,In_208);
nor U239 (N_239,In_521,In_192);
nand U240 (N_240,In_101,In_857);
nor U241 (N_241,In_0,In_795);
nor U242 (N_242,In_524,In_771);
nor U243 (N_243,In_67,In_204);
nor U244 (N_244,In_510,In_504);
or U245 (N_245,In_964,In_201);
nand U246 (N_246,In_160,In_294);
or U247 (N_247,In_972,In_679);
and U248 (N_248,In_317,In_829);
nand U249 (N_249,In_65,In_928);
xor U250 (N_250,In_622,In_715);
nor U251 (N_251,In_615,In_18);
nor U252 (N_252,In_516,In_40);
nor U253 (N_253,In_47,In_839);
nor U254 (N_254,In_827,In_742);
and U255 (N_255,In_292,In_301);
nand U256 (N_256,In_864,In_350);
nand U257 (N_257,In_385,In_330);
nor U258 (N_258,In_831,In_35);
nor U259 (N_259,In_564,In_865);
and U260 (N_260,In_805,In_796);
nand U261 (N_261,In_681,In_125);
nor U262 (N_262,In_285,In_809);
nor U263 (N_263,In_315,In_665);
or U264 (N_264,In_103,In_243);
nor U265 (N_265,In_327,In_71);
and U266 (N_266,In_353,In_643);
or U267 (N_267,In_825,In_386);
nand U268 (N_268,In_375,In_820);
nand U269 (N_269,In_450,In_153);
xnor U270 (N_270,In_780,In_503);
or U271 (N_271,In_837,In_165);
and U272 (N_272,In_15,In_242);
xnor U273 (N_273,In_610,In_197);
and U274 (N_274,In_377,In_438);
and U275 (N_275,In_304,In_309);
nand U276 (N_276,In_579,In_897);
and U277 (N_277,In_152,In_566);
and U278 (N_278,In_774,In_689);
and U279 (N_279,In_325,In_923);
or U280 (N_280,In_195,In_444);
nand U281 (N_281,In_209,In_162);
nor U282 (N_282,In_88,In_686);
and U283 (N_283,In_231,In_2);
and U284 (N_284,In_659,In_186);
nand U285 (N_285,In_78,In_251);
xnor U286 (N_286,In_146,In_91);
nor U287 (N_287,In_134,In_462);
xnor U288 (N_288,In_668,In_533);
or U289 (N_289,In_747,In_105);
or U290 (N_290,In_177,In_117);
or U291 (N_291,In_552,In_227);
and U292 (N_292,In_286,In_369);
nor U293 (N_293,In_708,In_531);
nor U294 (N_294,In_97,In_168);
nand U295 (N_295,In_157,In_80);
and U296 (N_296,In_859,In_577);
or U297 (N_297,In_362,In_955);
nor U298 (N_298,In_743,In_571);
nand U299 (N_299,In_498,In_866);
nand U300 (N_300,In_111,In_713);
and U301 (N_301,In_428,In_259);
nor U302 (N_302,In_647,In_989);
nor U303 (N_303,In_716,In_812);
nor U304 (N_304,In_136,In_959);
nor U305 (N_305,In_705,In_311);
and U306 (N_306,In_248,In_639);
and U307 (N_307,In_773,In_57);
and U308 (N_308,In_641,In_783);
nor U309 (N_309,In_398,In_161);
or U310 (N_310,In_710,In_371);
and U311 (N_311,In_911,In_717);
and U312 (N_312,In_467,In_396);
nor U313 (N_313,In_781,In_174);
nand U314 (N_314,In_454,In_995);
nor U315 (N_315,In_683,In_560);
nand U316 (N_316,In_917,In_419);
or U317 (N_317,In_726,In_883);
nor U318 (N_318,In_992,In_819);
xnor U319 (N_319,In_150,In_592);
nor U320 (N_320,In_760,In_983);
nand U321 (N_321,In_70,In_406);
or U322 (N_322,In_532,In_662);
xnor U323 (N_323,In_758,In_466);
xnor U324 (N_324,In_823,In_127);
and U325 (N_325,In_838,In_701);
nand U326 (N_326,In_334,In_193);
or U327 (N_327,In_891,In_966);
nor U328 (N_328,In_856,In_687);
and U329 (N_329,In_530,In_104);
or U330 (N_330,In_765,In_593);
nand U331 (N_331,In_704,In_855);
nor U332 (N_332,In_868,In_956);
nand U333 (N_333,In_852,In_667);
nor U334 (N_334,In_948,In_433);
nor U335 (N_335,In_887,In_110);
nor U336 (N_336,In_849,In_59);
and U337 (N_337,In_28,In_341);
or U338 (N_338,In_990,In_985);
nor U339 (N_339,In_368,In_7);
or U340 (N_340,In_393,In_402);
nand U341 (N_341,In_378,In_72);
or U342 (N_342,In_583,In_26);
nor U343 (N_343,In_99,In_624);
or U344 (N_344,In_262,In_477);
nand U345 (N_345,In_900,In_267);
and U346 (N_346,In_328,In_545);
and U347 (N_347,In_300,In_971);
and U348 (N_348,In_291,In_953);
or U349 (N_349,In_733,In_74);
nand U350 (N_350,In_631,In_963);
or U351 (N_351,In_407,In_777);
nor U352 (N_352,In_678,In_590);
xnor U353 (N_353,In_603,In_551);
and U354 (N_354,In_116,In_757);
and U355 (N_355,In_205,In_128);
and U356 (N_356,In_170,In_826);
or U357 (N_357,In_85,In_645);
nor U358 (N_358,In_881,In_36);
and U359 (N_359,In_987,In_148);
and U360 (N_360,In_835,In_166);
nor U361 (N_361,In_53,In_677);
nor U362 (N_362,In_938,In_490);
xor U363 (N_363,In_346,In_870);
or U364 (N_364,In_872,In_646);
nor U365 (N_365,In_278,In_734);
xnor U366 (N_366,In_892,In_374);
nor U367 (N_367,In_394,In_296);
or U368 (N_368,In_27,In_425);
nor U369 (N_369,In_199,In_976);
xor U370 (N_370,In_92,In_550);
nor U371 (N_371,In_587,In_281);
nand U372 (N_372,In_220,In_249);
or U373 (N_373,In_794,In_17);
and U374 (N_374,In_61,In_256);
and U375 (N_375,In_274,In_456);
nor U376 (N_376,In_95,In_422);
nor U377 (N_377,In_860,In_816);
xor U378 (N_378,In_73,In_663);
nand U379 (N_379,In_738,In_960);
nand U380 (N_380,In_458,In_935);
nor U381 (N_381,In_307,In_43);
and U382 (N_382,In_275,In_214);
xnor U383 (N_383,In_898,In_171);
nor U384 (N_384,In_806,In_319);
nand U385 (N_385,In_961,In_915);
nor U386 (N_386,In_491,In_967);
and U387 (N_387,In_501,In_502);
or U388 (N_388,In_954,In_379);
nor U389 (N_389,In_83,In_629);
and U390 (N_390,In_986,In_16);
and U391 (N_391,In_563,In_131);
or U392 (N_392,In_82,In_391);
and U393 (N_393,In_405,In_68);
nor U394 (N_394,In_493,In_684);
nand U395 (N_395,In_21,In_871);
nand U396 (N_396,In_924,In_879);
nand U397 (N_397,In_414,In_542);
nand U398 (N_398,In_528,In_721);
nor U399 (N_399,In_608,In_475);
nand U400 (N_400,In_93,In_618);
or U401 (N_401,In_962,In_822);
and U402 (N_402,In_706,In_461);
nand U403 (N_403,In_142,In_930);
and U404 (N_404,In_699,In_669);
and U405 (N_405,In_257,In_575);
nand U406 (N_406,In_853,In_714);
or U407 (N_407,In_889,In_591);
or U408 (N_408,In_483,In_427);
nor U409 (N_409,In_452,In_448);
nand U410 (N_410,In_581,In_895);
nand U411 (N_411,In_332,In_869);
or U412 (N_412,In_968,In_340);
and U413 (N_413,In_430,In_55);
nand U414 (N_414,In_426,In_60);
and U415 (N_415,In_342,In_818);
nand U416 (N_416,In_25,In_473);
and U417 (N_417,In_940,In_211);
nand U418 (N_418,In_130,In_813);
and U419 (N_419,In_841,In_279);
nor U420 (N_420,In_372,In_553);
nand U421 (N_421,In_497,In_676);
or U422 (N_422,In_558,In_194);
nor U423 (N_423,In_511,In_435);
nor U424 (N_424,In_749,In_845);
or U425 (N_425,In_712,In_89);
or U426 (N_426,In_90,In_410);
nand U427 (N_427,In_202,In_578);
xnor U428 (N_428,In_728,In_934);
or U429 (N_429,In_222,In_81);
xor U430 (N_430,In_240,In_363);
nor U431 (N_431,In_313,In_345);
and U432 (N_432,In_318,In_380);
nor U433 (N_433,In_943,In_744);
nor U434 (N_434,In_184,In_126);
or U435 (N_435,In_229,In_219);
nand U436 (N_436,In_893,In_492);
nand U437 (N_437,In_602,In_133);
and U438 (N_438,In_965,In_225);
and U439 (N_439,In_690,In_384);
and U440 (N_440,In_316,In_272);
and U441 (N_441,In_241,In_447);
nand U442 (N_442,In_5,In_52);
xnor U443 (N_443,In_817,In_440);
nor U444 (N_444,In_38,In_905);
and U445 (N_445,In_436,In_630);
or U446 (N_446,In_269,In_725);
or U447 (N_447,In_233,In_939);
nand U448 (N_448,In_23,In_750);
xor U449 (N_449,In_198,In_731);
nand U450 (N_450,In_753,In_223);
and U451 (N_451,In_899,In_633);
nand U452 (N_452,In_969,In_112);
or U453 (N_453,In_455,In_759);
and U454 (N_454,In_254,In_926);
or U455 (N_455,In_741,In_333);
and U456 (N_456,In_453,In_536);
and U457 (N_457,In_244,In_653);
and U458 (N_458,In_312,In_778);
xor U459 (N_459,In_299,In_693);
xor U460 (N_460,In_601,In_415);
or U461 (N_461,In_764,In_343);
xor U462 (N_462,In_779,In_237);
xnor U463 (N_463,In_308,In_58);
and U464 (N_464,In_417,In_387);
nor U465 (N_465,In_638,In_660);
nor U466 (N_466,In_46,In_66);
or U467 (N_467,In_185,In_685);
nand U468 (N_468,In_636,In_420);
nand U469 (N_469,In_132,In_605);
nand U470 (N_470,In_585,In_832);
or U471 (N_471,In_770,In_792);
nor U472 (N_472,In_620,In_182);
nand U473 (N_473,In_480,In_344);
nor U474 (N_474,In_846,In_408);
xnor U475 (N_475,In_514,In_937);
or U476 (N_476,In_206,In_196);
nand U477 (N_477,In_559,In_538);
and U478 (N_478,In_34,In_904);
nor U479 (N_479,In_356,In_399);
nor U480 (N_480,In_637,In_767);
and U481 (N_481,In_547,In_745);
or U482 (N_482,In_880,In_652);
nand U483 (N_483,In_154,In_505);
nand U484 (N_484,In_735,In_788);
nand U485 (N_485,In_401,In_138);
or U486 (N_486,In_520,In_896);
nand U487 (N_487,In_494,In_534);
and U488 (N_488,In_875,In_149);
nor U489 (N_489,In_688,In_762);
or U490 (N_490,In_702,In_785);
or U491 (N_491,In_851,In_302);
or U492 (N_492,In_666,In_673);
nand U493 (N_493,In_270,In_63);
nand U494 (N_494,In_8,In_515);
and U495 (N_495,In_974,In_582);
nor U496 (N_496,In_692,In_920);
nor U497 (N_497,In_314,In_432);
and U498 (N_498,In_522,In_509);
and U499 (N_499,In_657,In_418);
and U500 (N_500,In_54,In_872);
nand U501 (N_501,In_426,In_64);
or U502 (N_502,In_573,In_884);
and U503 (N_503,In_907,In_430);
or U504 (N_504,In_192,In_749);
nor U505 (N_505,In_520,In_959);
nor U506 (N_506,In_495,In_868);
nor U507 (N_507,In_101,In_273);
nand U508 (N_508,In_87,In_655);
xor U509 (N_509,In_358,In_115);
xnor U510 (N_510,In_966,In_960);
and U511 (N_511,In_272,In_485);
nor U512 (N_512,In_421,In_31);
or U513 (N_513,In_927,In_435);
or U514 (N_514,In_117,In_775);
nand U515 (N_515,In_274,In_442);
nor U516 (N_516,In_748,In_28);
and U517 (N_517,In_586,In_73);
nand U518 (N_518,In_931,In_568);
and U519 (N_519,In_517,In_303);
nand U520 (N_520,In_896,In_562);
nand U521 (N_521,In_134,In_547);
and U522 (N_522,In_182,In_40);
nor U523 (N_523,In_491,In_161);
and U524 (N_524,In_257,In_964);
and U525 (N_525,In_903,In_839);
and U526 (N_526,In_946,In_37);
nor U527 (N_527,In_221,In_304);
and U528 (N_528,In_608,In_556);
nor U529 (N_529,In_71,In_646);
xnor U530 (N_530,In_912,In_460);
nor U531 (N_531,In_99,In_745);
nor U532 (N_532,In_314,In_900);
or U533 (N_533,In_370,In_353);
nor U534 (N_534,In_343,In_592);
and U535 (N_535,In_67,In_472);
nand U536 (N_536,In_740,In_861);
nor U537 (N_537,In_642,In_290);
and U538 (N_538,In_47,In_561);
or U539 (N_539,In_824,In_869);
or U540 (N_540,In_660,In_466);
nand U541 (N_541,In_375,In_646);
nand U542 (N_542,In_134,In_722);
or U543 (N_543,In_895,In_727);
nor U544 (N_544,In_129,In_501);
nor U545 (N_545,In_987,In_396);
nor U546 (N_546,In_601,In_845);
or U547 (N_547,In_47,In_761);
and U548 (N_548,In_859,In_107);
xnor U549 (N_549,In_210,In_762);
nand U550 (N_550,In_994,In_525);
or U551 (N_551,In_12,In_783);
nand U552 (N_552,In_699,In_962);
or U553 (N_553,In_244,In_66);
xor U554 (N_554,In_687,In_497);
xor U555 (N_555,In_718,In_940);
xnor U556 (N_556,In_529,In_466);
xnor U557 (N_557,In_378,In_277);
xnor U558 (N_558,In_870,In_650);
nand U559 (N_559,In_71,In_3);
nor U560 (N_560,In_838,In_51);
nand U561 (N_561,In_659,In_261);
nand U562 (N_562,In_875,In_813);
nand U563 (N_563,In_878,In_83);
and U564 (N_564,In_313,In_632);
nor U565 (N_565,In_575,In_209);
nand U566 (N_566,In_571,In_394);
and U567 (N_567,In_117,In_803);
xnor U568 (N_568,In_294,In_915);
or U569 (N_569,In_216,In_60);
nor U570 (N_570,In_660,In_589);
nor U571 (N_571,In_564,In_516);
and U572 (N_572,In_817,In_595);
nand U573 (N_573,In_107,In_564);
nand U574 (N_574,In_210,In_328);
nand U575 (N_575,In_582,In_827);
nor U576 (N_576,In_462,In_964);
nor U577 (N_577,In_257,In_578);
nor U578 (N_578,In_761,In_260);
or U579 (N_579,In_169,In_262);
xnor U580 (N_580,In_31,In_635);
nand U581 (N_581,In_918,In_556);
or U582 (N_582,In_292,In_812);
and U583 (N_583,In_43,In_508);
nand U584 (N_584,In_20,In_735);
and U585 (N_585,In_247,In_45);
and U586 (N_586,In_238,In_453);
nor U587 (N_587,In_42,In_166);
nand U588 (N_588,In_650,In_109);
nor U589 (N_589,In_954,In_279);
nand U590 (N_590,In_627,In_802);
and U591 (N_591,In_866,In_961);
nand U592 (N_592,In_535,In_656);
nand U593 (N_593,In_372,In_810);
and U594 (N_594,In_308,In_411);
and U595 (N_595,In_345,In_508);
nand U596 (N_596,In_801,In_615);
or U597 (N_597,In_396,In_744);
xnor U598 (N_598,In_538,In_391);
nand U599 (N_599,In_322,In_908);
and U600 (N_600,In_390,In_510);
xor U601 (N_601,In_65,In_809);
nand U602 (N_602,In_17,In_401);
nor U603 (N_603,In_588,In_39);
and U604 (N_604,In_845,In_485);
and U605 (N_605,In_138,In_738);
nor U606 (N_606,In_150,In_914);
and U607 (N_607,In_964,In_783);
nor U608 (N_608,In_69,In_650);
nand U609 (N_609,In_916,In_646);
and U610 (N_610,In_884,In_843);
or U611 (N_611,In_100,In_600);
and U612 (N_612,In_46,In_922);
nor U613 (N_613,In_384,In_968);
or U614 (N_614,In_871,In_908);
nand U615 (N_615,In_282,In_346);
nand U616 (N_616,In_383,In_177);
nor U617 (N_617,In_842,In_774);
or U618 (N_618,In_929,In_139);
and U619 (N_619,In_880,In_446);
and U620 (N_620,In_817,In_463);
nand U621 (N_621,In_601,In_170);
or U622 (N_622,In_587,In_58);
or U623 (N_623,In_349,In_875);
nand U624 (N_624,In_913,In_430);
xnor U625 (N_625,In_184,In_658);
and U626 (N_626,In_899,In_197);
and U627 (N_627,In_992,In_627);
nor U628 (N_628,In_883,In_925);
nand U629 (N_629,In_718,In_126);
nor U630 (N_630,In_123,In_684);
nor U631 (N_631,In_457,In_584);
nand U632 (N_632,In_132,In_876);
and U633 (N_633,In_675,In_627);
nand U634 (N_634,In_811,In_253);
and U635 (N_635,In_232,In_435);
or U636 (N_636,In_537,In_87);
or U637 (N_637,In_827,In_918);
xnor U638 (N_638,In_524,In_38);
xnor U639 (N_639,In_610,In_130);
or U640 (N_640,In_700,In_921);
or U641 (N_641,In_511,In_256);
nand U642 (N_642,In_486,In_455);
and U643 (N_643,In_868,In_648);
and U644 (N_644,In_981,In_570);
nand U645 (N_645,In_357,In_897);
nand U646 (N_646,In_48,In_822);
nand U647 (N_647,In_185,In_81);
and U648 (N_648,In_739,In_139);
or U649 (N_649,In_385,In_678);
or U650 (N_650,In_565,In_52);
nand U651 (N_651,In_298,In_175);
and U652 (N_652,In_963,In_946);
nand U653 (N_653,In_619,In_115);
nand U654 (N_654,In_816,In_859);
or U655 (N_655,In_227,In_300);
or U656 (N_656,In_110,In_502);
nor U657 (N_657,In_303,In_549);
xor U658 (N_658,In_952,In_850);
xnor U659 (N_659,In_529,In_206);
nor U660 (N_660,In_387,In_227);
or U661 (N_661,In_397,In_14);
xnor U662 (N_662,In_562,In_50);
nand U663 (N_663,In_303,In_130);
or U664 (N_664,In_219,In_153);
nand U665 (N_665,In_611,In_370);
nor U666 (N_666,In_707,In_396);
nand U667 (N_667,In_214,In_659);
nor U668 (N_668,In_827,In_911);
nand U669 (N_669,In_227,In_184);
xor U670 (N_670,In_119,In_780);
or U671 (N_671,In_908,In_808);
and U672 (N_672,In_102,In_37);
nand U673 (N_673,In_631,In_265);
nor U674 (N_674,In_417,In_50);
nand U675 (N_675,In_651,In_102);
and U676 (N_676,In_567,In_29);
nand U677 (N_677,In_653,In_881);
and U678 (N_678,In_295,In_120);
nor U679 (N_679,In_936,In_87);
nand U680 (N_680,In_991,In_439);
or U681 (N_681,In_899,In_685);
and U682 (N_682,In_144,In_536);
and U683 (N_683,In_534,In_597);
and U684 (N_684,In_181,In_816);
xnor U685 (N_685,In_459,In_959);
nor U686 (N_686,In_785,In_705);
or U687 (N_687,In_461,In_382);
and U688 (N_688,In_923,In_967);
or U689 (N_689,In_366,In_812);
or U690 (N_690,In_869,In_973);
nand U691 (N_691,In_492,In_930);
nor U692 (N_692,In_755,In_283);
or U693 (N_693,In_611,In_221);
nand U694 (N_694,In_476,In_289);
or U695 (N_695,In_355,In_430);
nand U696 (N_696,In_719,In_492);
and U697 (N_697,In_974,In_753);
and U698 (N_698,In_220,In_298);
or U699 (N_699,In_919,In_700);
nor U700 (N_700,In_549,In_15);
and U701 (N_701,In_949,In_980);
or U702 (N_702,In_954,In_341);
or U703 (N_703,In_923,In_634);
nand U704 (N_704,In_781,In_974);
and U705 (N_705,In_827,In_986);
or U706 (N_706,In_509,In_153);
or U707 (N_707,In_19,In_390);
and U708 (N_708,In_340,In_150);
xnor U709 (N_709,In_788,In_855);
xnor U710 (N_710,In_53,In_444);
nand U711 (N_711,In_646,In_532);
nand U712 (N_712,In_311,In_557);
or U713 (N_713,In_318,In_72);
and U714 (N_714,In_564,In_800);
nand U715 (N_715,In_617,In_846);
nand U716 (N_716,In_897,In_111);
and U717 (N_717,In_225,In_294);
nor U718 (N_718,In_562,In_641);
or U719 (N_719,In_62,In_196);
or U720 (N_720,In_366,In_590);
or U721 (N_721,In_703,In_321);
or U722 (N_722,In_674,In_424);
xnor U723 (N_723,In_466,In_649);
nand U724 (N_724,In_522,In_550);
nor U725 (N_725,In_380,In_889);
nand U726 (N_726,In_838,In_137);
nor U727 (N_727,In_232,In_898);
nand U728 (N_728,In_317,In_847);
nor U729 (N_729,In_962,In_112);
or U730 (N_730,In_841,In_958);
or U731 (N_731,In_668,In_459);
xor U732 (N_732,In_259,In_710);
nor U733 (N_733,In_453,In_50);
and U734 (N_734,In_971,In_99);
nand U735 (N_735,In_459,In_160);
and U736 (N_736,In_690,In_849);
or U737 (N_737,In_819,In_837);
nor U738 (N_738,In_828,In_492);
xnor U739 (N_739,In_849,In_400);
nor U740 (N_740,In_508,In_10);
nor U741 (N_741,In_445,In_858);
nor U742 (N_742,In_292,In_593);
and U743 (N_743,In_719,In_143);
and U744 (N_744,In_485,In_943);
and U745 (N_745,In_167,In_114);
and U746 (N_746,In_670,In_970);
and U747 (N_747,In_702,In_682);
nand U748 (N_748,In_447,In_450);
nand U749 (N_749,In_241,In_501);
or U750 (N_750,In_364,In_481);
xor U751 (N_751,In_112,In_708);
nor U752 (N_752,In_549,In_725);
or U753 (N_753,In_660,In_20);
and U754 (N_754,In_368,In_40);
nor U755 (N_755,In_115,In_77);
nand U756 (N_756,In_632,In_595);
xnor U757 (N_757,In_696,In_21);
and U758 (N_758,In_135,In_397);
and U759 (N_759,In_173,In_859);
nand U760 (N_760,In_867,In_199);
xnor U761 (N_761,In_484,In_469);
nor U762 (N_762,In_439,In_965);
and U763 (N_763,In_478,In_125);
nor U764 (N_764,In_695,In_206);
or U765 (N_765,In_218,In_99);
nor U766 (N_766,In_752,In_605);
nor U767 (N_767,In_779,In_432);
xor U768 (N_768,In_242,In_7);
or U769 (N_769,In_379,In_42);
and U770 (N_770,In_537,In_245);
xor U771 (N_771,In_412,In_829);
xor U772 (N_772,In_216,In_176);
nor U773 (N_773,In_556,In_569);
nor U774 (N_774,In_397,In_902);
nor U775 (N_775,In_989,In_66);
xnor U776 (N_776,In_940,In_510);
nor U777 (N_777,In_238,In_246);
xor U778 (N_778,In_204,In_791);
or U779 (N_779,In_28,In_884);
nor U780 (N_780,In_523,In_940);
nand U781 (N_781,In_605,In_758);
or U782 (N_782,In_518,In_541);
nor U783 (N_783,In_258,In_688);
or U784 (N_784,In_590,In_242);
nand U785 (N_785,In_491,In_655);
nand U786 (N_786,In_524,In_84);
nor U787 (N_787,In_2,In_604);
nand U788 (N_788,In_235,In_984);
or U789 (N_789,In_433,In_887);
and U790 (N_790,In_962,In_188);
nand U791 (N_791,In_233,In_865);
nand U792 (N_792,In_300,In_419);
nor U793 (N_793,In_602,In_618);
or U794 (N_794,In_259,In_618);
and U795 (N_795,In_396,In_218);
nand U796 (N_796,In_752,In_912);
nor U797 (N_797,In_564,In_600);
and U798 (N_798,In_854,In_916);
or U799 (N_799,In_708,In_681);
or U800 (N_800,In_651,In_668);
or U801 (N_801,In_635,In_402);
nor U802 (N_802,In_267,In_439);
nand U803 (N_803,In_918,In_30);
and U804 (N_804,In_900,In_325);
nand U805 (N_805,In_801,In_646);
or U806 (N_806,In_24,In_941);
nand U807 (N_807,In_446,In_799);
nor U808 (N_808,In_154,In_731);
and U809 (N_809,In_598,In_39);
or U810 (N_810,In_220,In_251);
and U811 (N_811,In_190,In_776);
nor U812 (N_812,In_54,In_110);
nor U813 (N_813,In_260,In_785);
or U814 (N_814,In_854,In_627);
nand U815 (N_815,In_825,In_755);
nor U816 (N_816,In_534,In_900);
nand U817 (N_817,In_555,In_775);
nor U818 (N_818,In_266,In_111);
or U819 (N_819,In_49,In_858);
or U820 (N_820,In_475,In_547);
xor U821 (N_821,In_410,In_436);
xnor U822 (N_822,In_29,In_404);
and U823 (N_823,In_297,In_255);
and U824 (N_824,In_81,In_588);
and U825 (N_825,In_273,In_587);
nor U826 (N_826,In_245,In_785);
nand U827 (N_827,In_794,In_304);
nor U828 (N_828,In_394,In_961);
nor U829 (N_829,In_247,In_929);
nor U830 (N_830,In_265,In_965);
xnor U831 (N_831,In_144,In_148);
nand U832 (N_832,In_490,In_103);
xor U833 (N_833,In_302,In_379);
and U834 (N_834,In_604,In_504);
and U835 (N_835,In_577,In_151);
and U836 (N_836,In_290,In_663);
and U837 (N_837,In_934,In_843);
nand U838 (N_838,In_580,In_566);
nand U839 (N_839,In_697,In_744);
nor U840 (N_840,In_607,In_741);
nand U841 (N_841,In_472,In_34);
and U842 (N_842,In_189,In_321);
or U843 (N_843,In_316,In_754);
nor U844 (N_844,In_405,In_548);
nand U845 (N_845,In_364,In_218);
nor U846 (N_846,In_473,In_674);
xor U847 (N_847,In_34,In_293);
nor U848 (N_848,In_663,In_106);
nand U849 (N_849,In_730,In_122);
nand U850 (N_850,In_629,In_231);
nor U851 (N_851,In_244,In_993);
nand U852 (N_852,In_881,In_991);
or U853 (N_853,In_189,In_257);
and U854 (N_854,In_47,In_802);
nand U855 (N_855,In_266,In_976);
and U856 (N_856,In_288,In_431);
and U857 (N_857,In_371,In_864);
and U858 (N_858,In_250,In_753);
nand U859 (N_859,In_821,In_890);
xor U860 (N_860,In_566,In_284);
and U861 (N_861,In_973,In_388);
and U862 (N_862,In_389,In_87);
nor U863 (N_863,In_916,In_695);
or U864 (N_864,In_582,In_382);
nand U865 (N_865,In_613,In_276);
xnor U866 (N_866,In_532,In_716);
nor U867 (N_867,In_760,In_208);
nand U868 (N_868,In_573,In_74);
nand U869 (N_869,In_466,In_129);
and U870 (N_870,In_971,In_116);
and U871 (N_871,In_443,In_762);
nor U872 (N_872,In_127,In_252);
or U873 (N_873,In_414,In_230);
and U874 (N_874,In_770,In_315);
and U875 (N_875,In_357,In_170);
nor U876 (N_876,In_244,In_723);
and U877 (N_877,In_509,In_35);
nand U878 (N_878,In_556,In_756);
and U879 (N_879,In_303,In_283);
nor U880 (N_880,In_117,In_311);
nand U881 (N_881,In_798,In_359);
xor U882 (N_882,In_547,In_215);
and U883 (N_883,In_530,In_793);
and U884 (N_884,In_689,In_375);
nor U885 (N_885,In_942,In_35);
nand U886 (N_886,In_64,In_319);
nand U887 (N_887,In_498,In_549);
and U888 (N_888,In_23,In_295);
or U889 (N_889,In_569,In_633);
nand U890 (N_890,In_380,In_312);
nor U891 (N_891,In_925,In_46);
and U892 (N_892,In_407,In_843);
and U893 (N_893,In_302,In_958);
nand U894 (N_894,In_268,In_996);
nor U895 (N_895,In_382,In_251);
or U896 (N_896,In_842,In_481);
nor U897 (N_897,In_221,In_114);
nand U898 (N_898,In_374,In_544);
and U899 (N_899,In_246,In_83);
nor U900 (N_900,In_884,In_2);
and U901 (N_901,In_771,In_142);
or U902 (N_902,In_109,In_119);
and U903 (N_903,In_664,In_952);
and U904 (N_904,In_551,In_226);
nand U905 (N_905,In_855,In_196);
nand U906 (N_906,In_744,In_54);
nor U907 (N_907,In_833,In_183);
and U908 (N_908,In_303,In_97);
xnor U909 (N_909,In_977,In_36);
and U910 (N_910,In_138,In_729);
or U911 (N_911,In_451,In_221);
nor U912 (N_912,In_617,In_833);
and U913 (N_913,In_410,In_809);
or U914 (N_914,In_462,In_223);
or U915 (N_915,In_637,In_610);
nor U916 (N_916,In_852,In_166);
nand U917 (N_917,In_456,In_234);
nand U918 (N_918,In_995,In_315);
and U919 (N_919,In_81,In_116);
nor U920 (N_920,In_67,In_222);
and U921 (N_921,In_713,In_812);
and U922 (N_922,In_977,In_217);
nor U923 (N_923,In_552,In_170);
nand U924 (N_924,In_821,In_463);
and U925 (N_925,In_366,In_376);
nand U926 (N_926,In_931,In_692);
nor U927 (N_927,In_805,In_365);
and U928 (N_928,In_265,In_94);
xnor U929 (N_929,In_599,In_210);
and U930 (N_930,In_526,In_92);
and U931 (N_931,In_326,In_341);
nand U932 (N_932,In_788,In_679);
nand U933 (N_933,In_566,In_234);
or U934 (N_934,In_250,In_384);
xor U935 (N_935,In_973,In_520);
and U936 (N_936,In_462,In_556);
and U937 (N_937,In_19,In_599);
and U938 (N_938,In_534,In_519);
and U939 (N_939,In_364,In_181);
xor U940 (N_940,In_427,In_165);
nor U941 (N_941,In_867,In_264);
nand U942 (N_942,In_867,In_786);
or U943 (N_943,In_213,In_902);
nand U944 (N_944,In_147,In_371);
and U945 (N_945,In_127,In_701);
nor U946 (N_946,In_881,In_310);
and U947 (N_947,In_645,In_592);
or U948 (N_948,In_317,In_351);
nand U949 (N_949,In_423,In_129);
nor U950 (N_950,In_517,In_399);
nor U951 (N_951,In_874,In_69);
xnor U952 (N_952,In_496,In_957);
nand U953 (N_953,In_46,In_147);
nand U954 (N_954,In_550,In_326);
nand U955 (N_955,In_268,In_612);
or U956 (N_956,In_938,In_886);
nand U957 (N_957,In_371,In_616);
nand U958 (N_958,In_308,In_262);
and U959 (N_959,In_215,In_240);
nor U960 (N_960,In_288,In_593);
nor U961 (N_961,In_346,In_731);
and U962 (N_962,In_929,In_353);
or U963 (N_963,In_443,In_449);
nand U964 (N_964,In_461,In_588);
nand U965 (N_965,In_342,In_493);
or U966 (N_966,In_532,In_6);
nand U967 (N_967,In_400,In_163);
nand U968 (N_968,In_185,In_256);
nand U969 (N_969,In_554,In_359);
or U970 (N_970,In_586,In_222);
nand U971 (N_971,In_154,In_468);
nand U972 (N_972,In_36,In_757);
and U973 (N_973,In_645,In_256);
nand U974 (N_974,In_889,In_460);
nand U975 (N_975,In_547,In_609);
nor U976 (N_976,In_743,In_972);
xor U977 (N_977,In_903,In_214);
or U978 (N_978,In_312,In_3);
or U979 (N_979,In_433,In_728);
and U980 (N_980,In_802,In_302);
or U981 (N_981,In_795,In_781);
nand U982 (N_982,In_963,In_244);
or U983 (N_983,In_256,In_501);
or U984 (N_984,In_428,In_314);
xnor U985 (N_985,In_224,In_947);
nor U986 (N_986,In_429,In_722);
nor U987 (N_987,In_504,In_974);
or U988 (N_988,In_939,In_924);
and U989 (N_989,In_351,In_157);
nor U990 (N_990,In_747,In_985);
nand U991 (N_991,In_181,In_970);
and U992 (N_992,In_257,In_564);
nand U993 (N_993,In_929,In_349);
nor U994 (N_994,In_602,In_984);
nor U995 (N_995,In_124,In_283);
nand U996 (N_996,In_745,In_567);
and U997 (N_997,In_704,In_452);
and U998 (N_998,In_329,In_189);
nand U999 (N_999,In_755,In_675);
or U1000 (N_1000,In_629,In_987);
or U1001 (N_1001,In_917,In_160);
or U1002 (N_1002,In_625,In_278);
and U1003 (N_1003,In_331,In_555);
or U1004 (N_1004,In_326,In_971);
and U1005 (N_1005,In_456,In_915);
nand U1006 (N_1006,In_328,In_97);
and U1007 (N_1007,In_726,In_870);
nor U1008 (N_1008,In_852,In_937);
and U1009 (N_1009,In_326,In_945);
and U1010 (N_1010,In_825,In_374);
xnor U1011 (N_1011,In_673,In_465);
and U1012 (N_1012,In_6,In_632);
nor U1013 (N_1013,In_877,In_495);
and U1014 (N_1014,In_308,In_565);
or U1015 (N_1015,In_801,In_439);
and U1016 (N_1016,In_175,In_360);
nor U1017 (N_1017,In_707,In_187);
or U1018 (N_1018,In_746,In_294);
or U1019 (N_1019,In_590,In_21);
nor U1020 (N_1020,In_687,In_546);
and U1021 (N_1021,In_155,In_509);
nand U1022 (N_1022,In_99,In_228);
xor U1023 (N_1023,In_637,In_770);
nor U1024 (N_1024,In_732,In_846);
and U1025 (N_1025,In_557,In_855);
or U1026 (N_1026,In_658,In_822);
nand U1027 (N_1027,In_966,In_679);
xnor U1028 (N_1028,In_472,In_923);
nor U1029 (N_1029,In_520,In_256);
or U1030 (N_1030,In_192,In_404);
and U1031 (N_1031,In_913,In_928);
nand U1032 (N_1032,In_265,In_328);
nor U1033 (N_1033,In_325,In_743);
and U1034 (N_1034,In_59,In_610);
or U1035 (N_1035,In_176,In_589);
or U1036 (N_1036,In_695,In_775);
nand U1037 (N_1037,In_243,In_67);
and U1038 (N_1038,In_383,In_158);
nor U1039 (N_1039,In_664,In_194);
or U1040 (N_1040,In_208,In_786);
nand U1041 (N_1041,In_851,In_655);
nor U1042 (N_1042,In_487,In_860);
and U1043 (N_1043,In_359,In_95);
or U1044 (N_1044,In_626,In_834);
nor U1045 (N_1045,In_41,In_661);
nand U1046 (N_1046,In_388,In_734);
nor U1047 (N_1047,In_801,In_544);
nand U1048 (N_1048,In_580,In_573);
nand U1049 (N_1049,In_148,In_898);
nand U1050 (N_1050,In_129,In_93);
nand U1051 (N_1051,In_628,In_950);
and U1052 (N_1052,In_966,In_827);
or U1053 (N_1053,In_859,In_247);
nor U1054 (N_1054,In_732,In_858);
nor U1055 (N_1055,In_732,In_132);
and U1056 (N_1056,In_290,In_763);
nand U1057 (N_1057,In_504,In_773);
and U1058 (N_1058,In_255,In_258);
and U1059 (N_1059,In_926,In_744);
or U1060 (N_1060,In_884,In_581);
nor U1061 (N_1061,In_542,In_434);
nand U1062 (N_1062,In_416,In_485);
or U1063 (N_1063,In_904,In_184);
and U1064 (N_1064,In_46,In_109);
nand U1065 (N_1065,In_432,In_202);
xor U1066 (N_1066,In_277,In_859);
nor U1067 (N_1067,In_476,In_927);
xor U1068 (N_1068,In_28,In_875);
nor U1069 (N_1069,In_885,In_96);
or U1070 (N_1070,In_804,In_943);
xnor U1071 (N_1071,In_764,In_123);
nor U1072 (N_1072,In_102,In_65);
or U1073 (N_1073,In_645,In_410);
or U1074 (N_1074,In_683,In_399);
and U1075 (N_1075,In_530,In_943);
and U1076 (N_1076,In_286,In_529);
and U1077 (N_1077,In_422,In_625);
xor U1078 (N_1078,In_0,In_693);
or U1079 (N_1079,In_619,In_934);
nand U1080 (N_1080,In_701,In_158);
or U1081 (N_1081,In_866,In_596);
nand U1082 (N_1082,In_135,In_618);
nand U1083 (N_1083,In_196,In_654);
or U1084 (N_1084,In_828,In_772);
nor U1085 (N_1085,In_994,In_530);
and U1086 (N_1086,In_808,In_122);
nor U1087 (N_1087,In_4,In_790);
or U1088 (N_1088,In_463,In_249);
or U1089 (N_1089,In_723,In_616);
and U1090 (N_1090,In_649,In_390);
nand U1091 (N_1091,In_17,In_71);
nor U1092 (N_1092,In_820,In_543);
xnor U1093 (N_1093,In_872,In_184);
nor U1094 (N_1094,In_629,In_227);
nand U1095 (N_1095,In_205,In_424);
or U1096 (N_1096,In_397,In_405);
nand U1097 (N_1097,In_673,In_939);
nor U1098 (N_1098,In_340,In_254);
and U1099 (N_1099,In_687,In_678);
nor U1100 (N_1100,In_114,In_430);
and U1101 (N_1101,In_764,In_247);
nor U1102 (N_1102,In_554,In_571);
and U1103 (N_1103,In_983,In_994);
and U1104 (N_1104,In_371,In_647);
and U1105 (N_1105,In_26,In_742);
nor U1106 (N_1106,In_649,In_274);
nand U1107 (N_1107,In_351,In_874);
nand U1108 (N_1108,In_834,In_541);
nor U1109 (N_1109,In_300,In_794);
nand U1110 (N_1110,In_961,In_384);
nor U1111 (N_1111,In_984,In_93);
nor U1112 (N_1112,In_814,In_980);
nand U1113 (N_1113,In_767,In_2);
nand U1114 (N_1114,In_478,In_869);
nor U1115 (N_1115,In_911,In_471);
nor U1116 (N_1116,In_744,In_871);
nand U1117 (N_1117,In_306,In_568);
nor U1118 (N_1118,In_718,In_725);
nand U1119 (N_1119,In_423,In_930);
or U1120 (N_1120,In_293,In_764);
or U1121 (N_1121,In_775,In_506);
xor U1122 (N_1122,In_879,In_914);
nand U1123 (N_1123,In_473,In_882);
and U1124 (N_1124,In_926,In_937);
and U1125 (N_1125,In_198,In_300);
nor U1126 (N_1126,In_352,In_818);
nor U1127 (N_1127,In_829,In_998);
and U1128 (N_1128,In_591,In_911);
xor U1129 (N_1129,In_731,In_873);
and U1130 (N_1130,In_567,In_124);
or U1131 (N_1131,In_344,In_646);
nor U1132 (N_1132,In_911,In_224);
or U1133 (N_1133,In_205,In_150);
nor U1134 (N_1134,In_1,In_377);
or U1135 (N_1135,In_918,In_791);
and U1136 (N_1136,In_508,In_89);
nand U1137 (N_1137,In_536,In_830);
and U1138 (N_1138,In_866,In_485);
xnor U1139 (N_1139,In_192,In_442);
nor U1140 (N_1140,In_536,In_869);
or U1141 (N_1141,In_956,In_223);
and U1142 (N_1142,In_68,In_485);
or U1143 (N_1143,In_160,In_773);
nor U1144 (N_1144,In_230,In_998);
nor U1145 (N_1145,In_109,In_107);
nor U1146 (N_1146,In_499,In_445);
nor U1147 (N_1147,In_738,In_250);
and U1148 (N_1148,In_600,In_131);
nand U1149 (N_1149,In_220,In_441);
and U1150 (N_1150,In_961,In_545);
nor U1151 (N_1151,In_781,In_21);
or U1152 (N_1152,In_118,In_28);
or U1153 (N_1153,In_672,In_921);
and U1154 (N_1154,In_263,In_265);
nor U1155 (N_1155,In_303,In_325);
and U1156 (N_1156,In_473,In_332);
nand U1157 (N_1157,In_209,In_215);
xor U1158 (N_1158,In_134,In_830);
and U1159 (N_1159,In_526,In_187);
and U1160 (N_1160,In_557,In_762);
or U1161 (N_1161,In_205,In_802);
nand U1162 (N_1162,In_502,In_789);
or U1163 (N_1163,In_775,In_600);
nor U1164 (N_1164,In_211,In_630);
or U1165 (N_1165,In_587,In_2);
nand U1166 (N_1166,In_210,In_849);
and U1167 (N_1167,In_241,In_526);
nor U1168 (N_1168,In_851,In_456);
nor U1169 (N_1169,In_810,In_442);
and U1170 (N_1170,In_337,In_522);
and U1171 (N_1171,In_892,In_718);
nor U1172 (N_1172,In_612,In_97);
nand U1173 (N_1173,In_279,In_742);
nand U1174 (N_1174,In_469,In_612);
or U1175 (N_1175,In_628,In_679);
and U1176 (N_1176,In_121,In_845);
and U1177 (N_1177,In_415,In_577);
and U1178 (N_1178,In_155,In_150);
nand U1179 (N_1179,In_180,In_98);
nor U1180 (N_1180,In_233,In_354);
and U1181 (N_1181,In_636,In_3);
and U1182 (N_1182,In_799,In_457);
or U1183 (N_1183,In_447,In_271);
nor U1184 (N_1184,In_263,In_668);
or U1185 (N_1185,In_72,In_260);
and U1186 (N_1186,In_635,In_772);
and U1187 (N_1187,In_442,In_6);
and U1188 (N_1188,In_786,In_77);
xor U1189 (N_1189,In_400,In_21);
xnor U1190 (N_1190,In_12,In_518);
and U1191 (N_1191,In_395,In_412);
and U1192 (N_1192,In_658,In_355);
and U1193 (N_1193,In_964,In_815);
or U1194 (N_1194,In_489,In_36);
xor U1195 (N_1195,In_262,In_137);
nand U1196 (N_1196,In_113,In_871);
nand U1197 (N_1197,In_88,In_395);
nor U1198 (N_1198,In_469,In_30);
xnor U1199 (N_1199,In_607,In_991);
and U1200 (N_1200,In_634,In_555);
nand U1201 (N_1201,In_390,In_314);
nor U1202 (N_1202,In_180,In_901);
or U1203 (N_1203,In_780,In_647);
nor U1204 (N_1204,In_235,In_544);
nor U1205 (N_1205,In_807,In_382);
and U1206 (N_1206,In_788,In_406);
and U1207 (N_1207,In_599,In_95);
nand U1208 (N_1208,In_597,In_114);
nor U1209 (N_1209,In_937,In_556);
nor U1210 (N_1210,In_69,In_46);
nand U1211 (N_1211,In_631,In_61);
xor U1212 (N_1212,In_276,In_390);
or U1213 (N_1213,In_487,In_347);
nor U1214 (N_1214,In_539,In_93);
or U1215 (N_1215,In_363,In_523);
and U1216 (N_1216,In_428,In_874);
or U1217 (N_1217,In_603,In_370);
nand U1218 (N_1218,In_645,In_778);
or U1219 (N_1219,In_613,In_121);
nor U1220 (N_1220,In_44,In_95);
nor U1221 (N_1221,In_844,In_545);
or U1222 (N_1222,In_769,In_721);
or U1223 (N_1223,In_388,In_391);
and U1224 (N_1224,In_299,In_623);
and U1225 (N_1225,In_585,In_964);
nor U1226 (N_1226,In_222,In_628);
nor U1227 (N_1227,In_301,In_369);
nor U1228 (N_1228,In_606,In_300);
or U1229 (N_1229,In_431,In_316);
and U1230 (N_1230,In_346,In_8);
or U1231 (N_1231,In_805,In_942);
nand U1232 (N_1232,In_878,In_972);
xnor U1233 (N_1233,In_802,In_408);
and U1234 (N_1234,In_529,In_534);
nor U1235 (N_1235,In_493,In_932);
nor U1236 (N_1236,In_293,In_268);
or U1237 (N_1237,In_111,In_590);
and U1238 (N_1238,In_811,In_132);
nand U1239 (N_1239,In_465,In_26);
and U1240 (N_1240,In_57,In_911);
and U1241 (N_1241,In_943,In_679);
nor U1242 (N_1242,In_164,In_700);
or U1243 (N_1243,In_887,In_507);
nand U1244 (N_1244,In_75,In_835);
nand U1245 (N_1245,In_559,In_989);
nor U1246 (N_1246,In_188,In_271);
and U1247 (N_1247,In_624,In_851);
xnor U1248 (N_1248,In_716,In_216);
or U1249 (N_1249,In_593,In_228);
nor U1250 (N_1250,In_437,In_408);
or U1251 (N_1251,In_856,In_780);
or U1252 (N_1252,In_934,In_572);
and U1253 (N_1253,In_498,In_832);
nor U1254 (N_1254,In_678,In_979);
nand U1255 (N_1255,In_297,In_151);
and U1256 (N_1256,In_634,In_486);
or U1257 (N_1257,In_323,In_952);
nor U1258 (N_1258,In_766,In_275);
nand U1259 (N_1259,In_342,In_433);
nor U1260 (N_1260,In_618,In_227);
or U1261 (N_1261,In_960,In_632);
or U1262 (N_1262,In_410,In_885);
or U1263 (N_1263,In_166,In_821);
xnor U1264 (N_1264,In_596,In_788);
or U1265 (N_1265,In_290,In_75);
and U1266 (N_1266,In_655,In_81);
or U1267 (N_1267,In_968,In_811);
or U1268 (N_1268,In_522,In_961);
nor U1269 (N_1269,In_462,In_555);
or U1270 (N_1270,In_658,In_40);
nor U1271 (N_1271,In_146,In_610);
nor U1272 (N_1272,In_249,In_884);
nor U1273 (N_1273,In_151,In_723);
nand U1274 (N_1274,In_32,In_578);
nor U1275 (N_1275,In_239,In_382);
nand U1276 (N_1276,In_413,In_443);
or U1277 (N_1277,In_712,In_938);
nand U1278 (N_1278,In_961,In_462);
xnor U1279 (N_1279,In_946,In_919);
nor U1280 (N_1280,In_684,In_310);
and U1281 (N_1281,In_870,In_842);
xnor U1282 (N_1282,In_189,In_752);
nand U1283 (N_1283,In_52,In_700);
nor U1284 (N_1284,In_167,In_53);
and U1285 (N_1285,In_763,In_757);
nor U1286 (N_1286,In_710,In_573);
nor U1287 (N_1287,In_264,In_467);
and U1288 (N_1288,In_133,In_546);
or U1289 (N_1289,In_437,In_276);
nor U1290 (N_1290,In_96,In_90);
nand U1291 (N_1291,In_856,In_644);
or U1292 (N_1292,In_885,In_182);
or U1293 (N_1293,In_631,In_579);
xnor U1294 (N_1294,In_868,In_949);
nor U1295 (N_1295,In_158,In_905);
or U1296 (N_1296,In_980,In_617);
nand U1297 (N_1297,In_404,In_57);
nor U1298 (N_1298,In_416,In_728);
nand U1299 (N_1299,In_425,In_342);
and U1300 (N_1300,In_197,In_602);
nor U1301 (N_1301,In_926,In_880);
and U1302 (N_1302,In_113,In_555);
and U1303 (N_1303,In_25,In_187);
nand U1304 (N_1304,In_699,In_743);
nand U1305 (N_1305,In_584,In_717);
nor U1306 (N_1306,In_85,In_679);
or U1307 (N_1307,In_495,In_693);
or U1308 (N_1308,In_806,In_99);
nor U1309 (N_1309,In_556,In_444);
and U1310 (N_1310,In_668,In_113);
and U1311 (N_1311,In_684,In_978);
or U1312 (N_1312,In_61,In_779);
nand U1313 (N_1313,In_967,In_537);
nand U1314 (N_1314,In_4,In_288);
or U1315 (N_1315,In_824,In_648);
nand U1316 (N_1316,In_862,In_444);
and U1317 (N_1317,In_717,In_659);
or U1318 (N_1318,In_623,In_220);
nor U1319 (N_1319,In_591,In_705);
nor U1320 (N_1320,In_206,In_936);
nor U1321 (N_1321,In_776,In_368);
nor U1322 (N_1322,In_325,In_370);
or U1323 (N_1323,In_234,In_398);
nor U1324 (N_1324,In_144,In_580);
and U1325 (N_1325,In_232,In_923);
and U1326 (N_1326,In_935,In_288);
and U1327 (N_1327,In_798,In_178);
and U1328 (N_1328,In_149,In_776);
and U1329 (N_1329,In_392,In_4);
or U1330 (N_1330,In_484,In_848);
and U1331 (N_1331,In_936,In_589);
or U1332 (N_1332,In_442,In_660);
nor U1333 (N_1333,In_770,In_607);
nand U1334 (N_1334,In_174,In_399);
and U1335 (N_1335,In_550,In_968);
nand U1336 (N_1336,In_888,In_158);
nand U1337 (N_1337,In_474,In_45);
nor U1338 (N_1338,In_294,In_942);
nor U1339 (N_1339,In_303,In_54);
nor U1340 (N_1340,In_194,In_44);
or U1341 (N_1341,In_995,In_604);
nand U1342 (N_1342,In_783,In_751);
and U1343 (N_1343,In_584,In_193);
xor U1344 (N_1344,In_911,In_209);
or U1345 (N_1345,In_837,In_895);
and U1346 (N_1346,In_656,In_231);
and U1347 (N_1347,In_139,In_547);
or U1348 (N_1348,In_537,In_907);
nor U1349 (N_1349,In_858,In_930);
nand U1350 (N_1350,In_70,In_29);
nand U1351 (N_1351,In_503,In_981);
or U1352 (N_1352,In_680,In_344);
and U1353 (N_1353,In_269,In_359);
or U1354 (N_1354,In_568,In_911);
or U1355 (N_1355,In_32,In_874);
xor U1356 (N_1356,In_811,In_374);
or U1357 (N_1357,In_613,In_815);
and U1358 (N_1358,In_370,In_155);
nor U1359 (N_1359,In_845,In_554);
nand U1360 (N_1360,In_474,In_592);
or U1361 (N_1361,In_793,In_994);
nor U1362 (N_1362,In_3,In_321);
nand U1363 (N_1363,In_843,In_251);
or U1364 (N_1364,In_153,In_794);
nand U1365 (N_1365,In_87,In_985);
nor U1366 (N_1366,In_778,In_926);
or U1367 (N_1367,In_815,In_599);
or U1368 (N_1368,In_508,In_662);
nor U1369 (N_1369,In_467,In_207);
and U1370 (N_1370,In_292,In_474);
nor U1371 (N_1371,In_454,In_955);
and U1372 (N_1372,In_923,In_961);
nor U1373 (N_1373,In_978,In_641);
nor U1374 (N_1374,In_662,In_650);
and U1375 (N_1375,In_375,In_973);
nand U1376 (N_1376,In_355,In_855);
or U1377 (N_1377,In_624,In_706);
and U1378 (N_1378,In_958,In_827);
nor U1379 (N_1379,In_375,In_781);
or U1380 (N_1380,In_996,In_122);
nand U1381 (N_1381,In_630,In_243);
nand U1382 (N_1382,In_241,In_398);
nor U1383 (N_1383,In_114,In_49);
nand U1384 (N_1384,In_829,In_265);
or U1385 (N_1385,In_535,In_686);
nor U1386 (N_1386,In_888,In_622);
and U1387 (N_1387,In_140,In_950);
nor U1388 (N_1388,In_507,In_582);
nor U1389 (N_1389,In_112,In_992);
nand U1390 (N_1390,In_250,In_284);
nor U1391 (N_1391,In_378,In_679);
nand U1392 (N_1392,In_352,In_929);
or U1393 (N_1393,In_281,In_838);
and U1394 (N_1394,In_664,In_391);
xnor U1395 (N_1395,In_670,In_150);
nor U1396 (N_1396,In_701,In_754);
and U1397 (N_1397,In_755,In_911);
nor U1398 (N_1398,In_622,In_725);
nor U1399 (N_1399,In_611,In_182);
nor U1400 (N_1400,In_123,In_767);
nand U1401 (N_1401,In_909,In_364);
nand U1402 (N_1402,In_185,In_80);
nand U1403 (N_1403,In_55,In_275);
nor U1404 (N_1404,In_363,In_289);
nor U1405 (N_1405,In_733,In_10);
or U1406 (N_1406,In_998,In_930);
nand U1407 (N_1407,In_576,In_699);
nor U1408 (N_1408,In_488,In_973);
nor U1409 (N_1409,In_734,In_633);
nand U1410 (N_1410,In_610,In_474);
nor U1411 (N_1411,In_788,In_200);
nand U1412 (N_1412,In_42,In_210);
nor U1413 (N_1413,In_606,In_320);
nor U1414 (N_1414,In_554,In_734);
nand U1415 (N_1415,In_793,In_813);
nor U1416 (N_1416,In_401,In_880);
nor U1417 (N_1417,In_494,In_936);
or U1418 (N_1418,In_936,In_145);
or U1419 (N_1419,In_850,In_710);
and U1420 (N_1420,In_751,In_582);
nand U1421 (N_1421,In_980,In_193);
or U1422 (N_1422,In_967,In_616);
and U1423 (N_1423,In_344,In_837);
nor U1424 (N_1424,In_500,In_575);
xor U1425 (N_1425,In_858,In_149);
or U1426 (N_1426,In_236,In_577);
nor U1427 (N_1427,In_525,In_999);
and U1428 (N_1428,In_20,In_292);
xor U1429 (N_1429,In_174,In_305);
xor U1430 (N_1430,In_720,In_410);
nand U1431 (N_1431,In_856,In_638);
and U1432 (N_1432,In_937,In_77);
or U1433 (N_1433,In_290,In_14);
nand U1434 (N_1434,In_842,In_610);
nor U1435 (N_1435,In_439,In_21);
nor U1436 (N_1436,In_870,In_579);
nand U1437 (N_1437,In_776,In_967);
or U1438 (N_1438,In_867,In_540);
nand U1439 (N_1439,In_166,In_295);
nand U1440 (N_1440,In_957,In_161);
and U1441 (N_1441,In_340,In_667);
and U1442 (N_1442,In_16,In_258);
and U1443 (N_1443,In_273,In_768);
and U1444 (N_1444,In_21,In_240);
or U1445 (N_1445,In_274,In_26);
nor U1446 (N_1446,In_805,In_121);
nand U1447 (N_1447,In_653,In_586);
and U1448 (N_1448,In_183,In_615);
nand U1449 (N_1449,In_60,In_773);
and U1450 (N_1450,In_175,In_613);
nand U1451 (N_1451,In_31,In_710);
or U1452 (N_1452,In_368,In_103);
nor U1453 (N_1453,In_952,In_12);
nor U1454 (N_1454,In_96,In_487);
nand U1455 (N_1455,In_156,In_189);
nor U1456 (N_1456,In_302,In_886);
xor U1457 (N_1457,In_366,In_636);
nand U1458 (N_1458,In_588,In_100);
nand U1459 (N_1459,In_697,In_101);
or U1460 (N_1460,In_489,In_228);
nand U1461 (N_1461,In_127,In_521);
and U1462 (N_1462,In_809,In_563);
and U1463 (N_1463,In_64,In_831);
xnor U1464 (N_1464,In_273,In_832);
and U1465 (N_1465,In_725,In_648);
xnor U1466 (N_1466,In_830,In_5);
or U1467 (N_1467,In_50,In_616);
and U1468 (N_1468,In_202,In_836);
and U1469 (N_1469,In_195,In_604);
or U1470 (N_1470,In_253,In_710);
nor U1471 (N_1471,In_872,In_837);
nand U1472 (N_1472,In_748,In_841);
or U1473 (N_1473,In_229,In_617);
or U1474 (N_1474,In_886,In_346);
nor U1475 (N_1475,In_878,In_46);
nor U1476 (N_1476,In_398,In_257);
nand U1477 (N_1477,In_199,In_685);
nor U1478 (N_1478,In_831,In_526);
nor U1479 (N_1479,In_27,In_11);
nor U1480 (N_1480,In_402,In_680);
nand U1481 (N_1481,In_97,In_961);
and U1482 (N_1482,In_735,In_247);
xor U1483 (N_1483,In_48,In_385);
or U1484 (N_1484,In_222,In_220);
nor U1485 (N_1485,In_130,In_852);
or U1486 (N_1486,In_946,In_424);
nand U1487 (N_1487,In_951,In_36);
or U1488 (N_1488,In_93,In_583);
or U1489 (N_1489,In_587,In_576);
nor U1490 (N_1490,In_733,In_154);
nand U1491 (N_1491,In_38,In_224);
nor U1492 (N_1492,In_201,In_828);
nor U1493 (N_1493,In_592,In_448);
nand U1494 (N_1494,In_992,In_488);
or U1495 (N_1495,In_979,In_764);
nor U1496 (N_1496,In_669,In_477);
and U1497 (N_1497,In_578,In_483);
or U1498 (N_1498,In_493,In_440);
and U1499 (N_1499,In_461,In_393);
or U1500 (N_1500,In_968,In_567);
nor U1501 (N_1501,In_726,In_49);
and U1502 (N_1502,In_270,In_390);
and U1503 (N_1503,In_176,In_235);
nor U1504 (N_1504,In_809,In_617);
nand U1505 (N_1505,In_44,In_877);
nand U1506 (N_1506,In_181,In_10);
and U1507 (N_1507,In_214,In_426);
nor U1508 (N_1508,In_831,In_349);
nand U1509 (N_1509,In_574,In_18);
nor U1510 (N_1510,In_225,In_666);
xnor U1511 (N_1511,In_560,In_390);
nand U1512 (N_1512,In_340,In_769);
nor U1513 (N_1513,In_652,In_537);
and U1514 (N_1514,In_674,In_777);
xnor U1515 (N_1515,In_743,In_354);
nand U1516 (N_1516,In_245,In_885);
or U1517 (N_1517,In_723,In_671);
nor U1518 (N_1518,In_160,In_25);
nand U1519 (N_1519,In_783,In_927);
xor U1520 (N_1520,In_455,In_270);
nand U1521 (N_1521,In_793,In_491);
nand U1522 (N_1522,In_795,In_793);
and U1523 (N_1523,In_120,In_144);
nand U1524 (N_1524,In_154,In_437);
or U1525 (N_1525,In_812,In_800);
and U1526 (N_1526,In_547,In_410);
and U1527 (N_1527,In_3,In_305);
nor U1528 (N_1528,In_461,In_12);
or U1529 (N_1529,In_176,In_365);
nor U1530 (N_1530,In_586,In_338);
and U1531 (N_1531,In_243,In_628);
and U1532 (N_1532,In_957,In_463);
and U1533 (N_1533,In_13,In_430);
or U1534 (N_1534,In_428,In_929);
or U1535 (N_1535,In_280,In_846);
or U1536 (N_1536,In_850,In_475);
nand U1537 (N_1537,In_726,In_880);
or U1538 (N_1538,In_864,In_259);
or U1539 (N_1539,In_778,In_984);
or U1540 (N_1540,In_144,In_472);
nor U1541 (N_1541,In_291,In_902);
or U1542 (N_1542,In_437,In_492);
nand U1543 (N_1543,In_31,In_332);
or U1544 (N_1544,In_185,In_564);
or U1545 (N_1545,In_656,In_277);
and U1546 (N_1546,In_690,In_928);
nand U1547 (N_1547,In_508,In_551);
and U1548 (N_1548,In_98,In_498);
nor U1549 (N_1549,In_644,In_161);
or U1550 (N_1550,In_441,In_972);
xnor U1551 (N_1551,In_818,In_411);
nor U1552 (N_1552,In_349,In_404);
xnor U1553 (N_1553,In_752,In_627);
nor U1554 (N_1554,In_550,In_454);
and U1555 (N_1555,In_724,In_613);
or U1556 (N_1556,In_601,In_286);
or U1557 (N_1557,In_981,In_770);
xor U1558 (N_1558,In_706,In_951);
nor U1559 (N_1559,In_190,In_250);
nand U1560 (N_1560,In_235,In_831);
or U1561 (N_1561,In_625,In_74);
and U1562 (N_1562,In_726,In_209);
nor U1563 (N_1563,In_796,In_292);
nand U1564 (N_1564,In_486,In_176);
nand U1565 (N_1565,In_676,In_553);
or U1566 (N_1566,In_102,In_781);
and U1567 (N_1567,In_676,In_750);
nor U1568 (N_1568,In_508,In_154);
and U1569 (N_1569,In_86,In_843);
xor U1570 (N_1570,In_158,In_739);
xor U1571 (N_1571,In_969,In_671);
nand U1572 (N_1572,In_603,In_342);
or U1573 (N_1573,In_557,In_196);
nand U1574 (N_1574,In_84,In_750);
or U1575 (N_1575,In_302,In_185);
and U1576 (N_1576,In_728,In_521);
nand U1577 (N_1577,In_318,In_76);
nand U1578 (N_1578,In_814,In_380);
nor U1579 (N_1579,In_916,In_204);
xnor U1580 (N_1580,In_225,In_742);
nand U1581 (N_1581,In_956,In_491);
or U1582 (N_1582,In_333,In_415);
or U1583 (N_1583,In_266,In_909);
or U1584 (N_1584,In_618,In_94);
nand U1585 (N_1585,In_203,In_640);
and U1586 (N_1586,In_861,In_372);
nand U1587 (N_1587,In_861,In_608);
nor U1588 (N_1588,In_205,In_762);
or U1589 (N_1589,In_895,In_122);
and U1590 (N_1590,In_608,In_311);
nor U1591 (N_1591,In_386,In_634);
xor U1592 (N_1592,In_417,In_960);
and U1593 (N_1593,In_785,In_721);
nand U1594 (N_1594,In_51,In_617);
or U1595 (N_1595,In_24,In_272);
nand U1596 (N_1596,In_713,In_483);
and U1597 (N_1597,In_415,In_863);
nand U1598 (N_1598,In_13,In_135);
nor U1599 (N_1599,In_748,In_20);
and U1600 (N_1600,In_749,In_318);
or U1601 (N_1601,In_725,In_768);
and U1602 (N_1602,In_206,In_89);
nand U1603 (N_1603,In_348,In_724);
and U1604 (N_1604,In_713,In_947);
or U1605 (N_1605,In_230,In_397);
nand U1606 (N_1606,In_989,In_6);
and U1607 (N_1607,In_782,In_805);
and U1608 (N_1608,In_543,In_665);
nand U1609 (N_1609,In_163,In_691);
nor U1610 (N_1610,In_626,In_58);
or U1611 (N_1611,In_669,In_384);
and U1612 (N_1612,In_455,In_979);
or U1613 (N_1613,In_124,In_73);
xor U1614 (N_1614,In_665,In_961);
nor U1615 (N_1615,In_980,In_124);
or U1616 (N_1616,In_594,In_407);
and U1617 (N_1617,In_927,In_131);
or U1618 (N_1618,In_82,In_128);
nand U1619 (N_1619,In_859,In_203);
nand U1620 (N_1620,In_291,In_920);
and U1621 (N_1621,In_945,In_36);
or U1622 (N_1622,In_882,In_422);
and U1623 (N_1623,In_577,In_283);
or U1624 (N_1624,In_513,In_146);
xnor U1625 (N_1625,In_478,In_324);
nand U1626 (N_1626,In_869,In_822);
nand U1627 (N_1627,In_468,In_270);
or U1628 (N_1628,In_51,In_847);
nor U1629 (N_1629,In_363,In_973);
xor U1630 (N_1630,In_605,In_713);
or U1631 (N_1631,In_872,In_685);
nor U1632 (N_1632,In_352,In_869);
and U1633 (N_1633,In_385,In_961);
or U1634 (N_1634,In_200,In_452);
or U1635 (N_1635,In_532,In_943);
or U1636 (N_1636,In_24,In_110);
nand U1637 (N_1637,In_463,In_179);
or U1638 (N_1638,In_326,In_393);
nor U1639 (N_1639,In_222,In_446);
or U1640 (N_1640,In_253,In_547);
and U1641 (N_1641,In_834,In_437);
nor U1642 (N_1642,In_888,In_966);
or U1643 (N_1643,In_440,In_888);
or U1644 (N_1644,In_837,In_876);
nand U1645 (N_1645,In_525,In_197);
xnor U1646 (N_1646,In_0,In_816);
or U1647 (N_1647,In_989,In_444);
and U1648 (N_1648,In_783,In_800);
nor U1649 (N_1649,In_600,In_901);
and U1650 (N_1650,In_979,In_48);
nand U1651 (N_1651,In_546,In_782);
nand U1652 (N_1652,In_238,In_5);
nor U1653 (N_1653,In_295,In_805);
nor U1654 (N_1654,In_293,In_888);
nor U1655 (N_1655,In_475,In_698);
nand U1656 (N_1656,In_51,In_996);
nor U1657 (N_1657,In_751,In_875);
nor U1658 (N_1658,In_131,In_823);
nor U1659 (N_1659,In_504,In_458);
nand U1660 (N_1660,In_2,In_574);
nand U1661 (N_1661,In_681,In_733);
xor U1662 (N_1662,In_931,In_675);
and U1663 (N_1663,In_403,In_91);
or U1664 (N_1664,In_927,In_967);
or U1665 (N_1665,In_180,In_92);
and U1666 (N_1666,In_963,In_866);
and U1667 (N_1667,In_116,In_695);
nor U1668 (N_1668,In_519,In_10);
and U1669 (N_1669,In_976,In_947);
xor U1670 (N_1670,In_919,In_755);
xnor U1671 (N_1671,In_73,In_917);
xnor U1672 (N_1672,In_774,In_617);
nor U1673 (N_1673,In_819,In_506);
xor U1674 (N_1674,In_264,In_496);
xor U1675 (N_1675,In_441,In_722);
nand U1676 (N_1676,In_736,In_315);
or U1677 (N_1677,In_595,In_390);
xor U1678 (N_1678,In_469,In_107);
nor U1679 (N_1679,In_125,In_972);
nor U1680 (N_1680,In_463,In_223);
xnor U1681 (N_1681,In_499,In_76);
and U1682 (N_1682,In_123,In_392);
or U1683 (N_1683,In_533,In_342);
nand U1684 (N_1684,In_137,In_418);
nor U1685 (N_1685,In_256,In_794);
and U1686 (N_1686,In_842,In_486);
xor U1687 (N_1687,In_43,In_391);
nand U1688 (N_1688,In_421,In_209);
or U1689 (N_1689,In_852,In_271);
xor U1690 (N_1690,In_853,In_477);
and U1691 (N_1691,In_863,In_508);
nor U1692 (N_1692,In_634,In_252);
or U1693 (N_1693,In_896,In_122);
nor U1694 (N_1694,In_136,In_761);
nor U1695 (N_1695,In_217,In_280);
nor U1696 (N_1696,In_332,In_990);
and U1697 (N_1697,In_416,In_96);
or U1698 (N_1698,In_690,In_817);
and U1699 (N_1699,In_167,In_778);
nand U1700 (N_1700,In_304,In_926);
xnor U1701 (N_1701,In_809,In_346);
nor U1702 (N_1702,In_696,In_96);
nor U1703 (N_1703,In_131,In_726);
nand U1704 (N_1704,In_340,In_772);
nor U1705 (N_1705,In_390,In_263);
nand U1706 (N_1706,In_545,In_217);
nand U1707 (N_1707,In_797,In_530);
xor U1708 (N_1708,In_474,In_629);
and U1709 (N_1709,In_212,In_298);
xor U1710 (N_1710,In_783,In_288);
nor U1711 (N_1711,In_516,In_401);
nand U1712 (N_1712,In_82,In_810);
nor U1713 (N_1713,In_38,In_491);
or U1714 (N_1714,In_449,In_53);
or U1715 (N_1715,In_833,In_469);
nor U1716 (N_1716,In_111,In_559);
and U1717 (N_1717,In_380,In_633);
and U1718 (N_1718,In_723,In_265);
and U1719 (N_1719,In_403,In_511);
nor U1720 (N_1720,In_0,In_344);
nor U1721 (N_1721,In_174,In_555);
or U1722 (N_1722,In_147,In_772);
nor U1723 (N_1723,In_819,In_946);
xor U1724 (N_1724,In_763,In_808);
and U1725 (N_1725,In_95,In_41);
nor U1726 (N_1726,In_991,In_497);
nand U1727 (N_1727,In_864,In_345);
nand U1728 (N_1728,In_839,In_764);
xor U1729 (N_1729,In_863,In_520);
xnor U1730 (N_1730,In_724,In_786);
nand U1731 (N_1731,In_323,In_367);
or U1732 (N_1732,In_349,In_81);
xor U1733 (N_1733,In_847,In_503);
or U1734 (N_1734,In_815,In_630);
or U1735 (N_1735,In_372,In_358);
nor U1736 (N_1736,In_94,In_705);
or U1737 (N_1737,In_683,In_255);
nor U1738 (N_1738,In_779,In_26);
nor U1739 (N_1739,In_685,In_319);
and U1740 (N_1740,In_879,In_645);
xnor U1741 (N_1741,In_679,In_152);
nor U1742 (N_1742,In_245,In_421);
or U1743 (N_1743,In_262,In_807);
or U1744 (N_1744,In_182,In_177);
nand U1745 (N_1745,In_354,In_15);
or U1746 (N_1746,In_792,In_204);
and U1747 (N_1747,In_871,In_742);
or U1748 (N_1748,In_828,In_816);
xor U1749 (N_1749,In_548,In_640);
and U1750 (N_1750,In_742,In_765);
and U1751 (N_1751,In_889,In_765);
or U1752 (N_1752,In_993,In_746);
nor U1753 (N_1753,In_361,In_446);
nor U1754 (N_1754,In_555,In_70);
or U1755 (N_1755,In_877,In_7);
nand U1756 (N_1756,In_86,In_338);
nor U1757 (N_1757,In_64,In_259);
and U1758 (N_1758,In_525,In_285);
and U1759 (N_1759,In_4,In_672);
or U1760 (N_1760,In_777,In_781);
nand U1761 (N_1761,In_741,In_316);
or U1762 (N_1762,In_493,In_172);
nor U1763 (N_1763,In_601,In_776);
nor U1764 (N_1764,In_420,In_15);
and U1765 (N_1765,In_44,In_401);
or U1766 (N_1766,In_28,In_712);
nor U1767 (N_1767,In_147,In_388);
and U1768 (N_1768,In_348,In_84);
or U1769 (N_1769,In_237,In_408);
or U1770 (N_1770,In_640,In_753);
or U1771 (N_1771,In_723,In_103);
nor U1772 (N_1772,In_635,In_132);
or U1773 (N_1773,In_959,In_598);
and U1774 (N_1774,In_96,In_934);
or U1775 (N_1775,In_158,In_52);
and U1776 (N_1776,In_929,In_381);
nand U1777 (N_1777,In_35,In_529);
nor U1778 (N_1778,In_777,In_92);
and U1779 (N_1779,In_682,In_442);
nand U1780 (N_1780,In_7,In_180);
or U1781 (N_1781,In_754,In_906);
nor U1782 (N_1782,In_381,In_305);
nand U1783 (N_1783,In_836,In_106);
xor U1784 (N_1784,In_434,In_802);
nand U1785 (N_1785,In_426,In_770);
or U1786 (N_1786,In_2,In_744);
nand U1787 (N_1787,In_663,In_985);
or U1788 (N_1788,In_372,In_814);
nor U1789 (N_1789,In_90,In_614);
or U1790 (N_1790,In_738,In_796);
nand U1791 (N_1791,In_10,In_642);
nand U1792 (N_1792,In_976,In_471);
or U1793 (N_1793,In_36,In_849);
or U1794 (N_1794,In_582,In_730);
and U1795 (N_1795,In_731,In_147);
nand U1796 (N_1796,In_270,In_172);
and U1797 (N_1797,In_825,In_753);
or U1798 (N_1798,In_988,In_484);
xor U1799 (N_1799,In_860,In_395);
and U1800 (N_1800,In_715,In_518);
nor U1801 (N_1801,In_437,In_935);
nor U1802 (N_1802,In_488,In_974);
nor U1803 (N_1803,In_163,In_19);
and U1804 (N_1804,In_224,In_575);
nor U1805 (N_1805,In_422,In_21);
nor U1806 (N_1806,In_177,In_545);
nand U1807 (N_1807,In_968,In_944);
xnor U1808 (N_1808,In_661,In_618);
xor U1809 (N_1809,In_193,In_302);
nor U1810 (N_1810,In_96,In_957);
or U1811 (N_1811,In_116,In_47);
nand U1812 (N_1812,In_270,In_340);
and U1813 (N_1813,In_837,In_623);
nand U1814 (N_1814,In_853,In_285);
and U1815 (N_1815,In_651,In_211);
nand U1816 (N_1816,In_839,In_465);
xnor U1817 (N_1817,In_445,In_16);
and U1818 (N_1818,In_812,In_394);
or U1819 (N_1819,In_722,In_494);
and U1820 (N_1820,In_484,In_935);
or U1821 (N_1821,In_802,In_797);
and U1822 (N_1822,In_719,In_586);
nor U1823 (N_1823,In_522,In_86);
nor U1824 (N_1824,In_841,In_128);
and U1825 (N_1825,In_894,In_272);
or U1826 (N_1826,In_778,In_26);
and U1827 (N_1827,In_648,In_688);
or U1828 (N_1828,In_377,In_698);
nor U1829 (N_1829,In_982,In_834);
nand U1830 (N_1830,In_982,In_411);
nor U1831 (N_1831,In_446,In_289);
nand U1832 (N_1832,In_847,In_249);
nand U1833 (N_1833,In_965,In_887);
nor U1834 (N_1834,In_324,In_147);
nand U1835 (N_1835,In_42,In_419);
or U1836 (N_1836,In_509,In_798);
nor U1837 (N_1837,In_645,In_12);
xor U1838 (N_1838,In_539,In_801);
and U1839 (N_1839,In_140,In_139);
and U1840 (N_1840,In_537,In_320);
nand U1841 (N_1841,In_998,In_23);
nand U1842 (N_1842,In_155,In_448);
and U1843 (N_1843,In_547,In_367);
or U1844 (N_1844,In_340,In_156);
and U1845 (N_1845,In_912,In_642);
nand U1846 (N_1846,In_49,In_71);
nand U1847 (N_1847,In_371,In_288);
and U1848 (N_1848,In_746,In_634);
nand U1849 (N_1849,In_482,In_574);
nand U1850 (N_1850,In_315,In_392);
nor U1851 (N_1851,In_935,In_169);
nand U1852 (N_1852,In_49,In_93);
nand U1853 (N_1853,In_708,In_166);
or U1854 (N_1854,In_978,In_777);
or U1855 (N_1855,In_266,In_655);
or U1856 (N_1856,In_627,In_654);
xor U1857 (N_1857,In_499,In_546);
nand U1858 (N_1858,In_602,In_737);
or U1859 (N_1859,In_494,In_896);
or U1860 (N_1860,In_176,In_450);
xnor U1861 (N_1861,In_65,In_555);
xor U1862 (N_1862,In_874,In_446);
and U1863 (N_1863,In_773,In_457);
nor U1864 (N_1864,In_931,In_547);
or U1865 (N_1865,In_26,In_986);
and U1866 (N_1866,In_45,In_633);
nand U1867 (N_1867,In_715,In_684);
and U1868 (N_1868,In_79,In_319);
and U1869 (N_1869,In_368,In_974);
and U1870 (N_1870,In_604,In_322);
nand U1871 (N_1871,In_677,In_867);
xnor U1872 (N_1872,In_134,In_872);
or U1873 (N_1873,In_865,In_608);
nand U1874 (N_1874,In_489,In_113);
or U1875 (N_1875,In_489,In_4);
and U1876 (N_1876,In_301,In_822);
xnor U1877 (N_1877,In_540,In_489);
xnor U1878 (N_1878,In_318,In_649);
or U1879 (N_1879,In_34,In_46);
and U1880 (N_1880,In_138,In_497);
and U1881 (N_1881,In_979,In_660);
or U1882 (N_1882,In_228,In_151);
and U1883 (N_1883,In_230,In_442);
or U1884 (N_1884,In_395,In_431);
nand U1885 (N_1885,In_984,In_485);
and U1886 (N_1886,In_145,In_883);
nand U1887 (N_1887,In_925,In_99);
and U1888 (N_1888,In_120,In_852);
nand U1889 (N_1889,In_154,In_120);
nand U1890 (N_1890,In_689,In_964);
nand U1891 (N_1891,In_110,In_722);
xor U1892 (N_1892,In_130,In_12);
and U1893 (N_1893,In_120,In_959);
and U1894 (N_1894,In_138,In_919);
xnor U1895 (N_1895,In_107,In_227);
xor U1896 (N_1896,In_694,In_503);
and U1897 (N_1897,In_684,In_730);
nor U1898 (N_1898,In_296,In_961);
nor U1899 (N_1899,In_310,In_112);
nor U1900 (N_1900,In_777,In_328);
and U1901 (N_1901,In_849,In_738);
nor U1902 (N_1902,In_329,In_397);
or U1903 (N_1903,In_387,In_94);
or U1904 (N_1904,In_746,In_275);
nand U1905 (N_1905,In_310,In_892);
and U1906 (N_1906,In_38,In_84);
nor U1907 (N_1907,In_531,In_757);
nor U1908 (N_1908,In_376,In_681);
nand U1909 (N_1909,In_127,In_119);
nor U1910 (N_1910,In_118,In_923);
xor U1911 (N_1911,In_381,In_578);
and U1912 (N_1912,In_748,In_984);
nor U1913 (N_1913,In_638,In_603);
xnor U1914 (N_1914,In_23,In_950);
or U1915 (N_1915,In_348,In_806);
nor U1916 (N_1916,In_258,In_201);
nor U1917 (N_1917,In_401,In_136);
nand U1918 (N_1918,In_610,In_258);
xnor U1919 (N_1919,In_990,In_571);
xnor U1920 (N_1920,In_855,In_858);
nor U1921 (N_1921,In_992,In_371);
or U1922 (N_1922,In_787,In_821);
xnor U1923 (N_1923,In_186,In_417);
or U1924 (N_1924,In_237,In_965);
and U1925 (N_1925,In_658,In_982);
and U1926 (N_1926,In_378,In_521);
nor U1927 (N_1927,In_772,In_49);
nand U1928 (N_1928,In_684,In_263);
nand U1929 (N_1929,In_73,In_234);
nor U1930 (N_1930,In_998,In_700);
xor U1931 (N_1931,In_135,In_170);
or U1932 (N_1932,In_828,In_734);
and U1933 (N_1933,In_878,In_407);
and U1934 (N_1934,In_308,In_549);
and U1935 (N_1935,In_273,In_975);
nand U1936 (N_1936,In_880,In_452);
and U1937 (N_1937,In_229,In_34);
and U1938 (N_1938,In_305,In_580);
nand U1939 (N_1939,In_0,In_870);
and U1940 (N_1940,In_921,In_690);
nor U1941 (N_1941,In_523,In_275);
nor U1942 (N_1942,In_536,In_893);
and U1943 (N_1943,In_511,In_125);
nor U1944 (N_1944,In_334,In_757);
nor U1945 (N_1945,In_511,In_231);
nand U1946 (N_1946,In_773,In_16);
or U1947 (N_1947,In_379,In_618);
nor U1948 (N_1948,In_831,In_538);
and U1949 (N_1949,In_306,In_421);
nor U1950 (N_1950,In_985,In_226);
and U1951 (N_1951,In_59,In_708);
or U1952 (N_1952,In_872,In_419);
or U1953 (N_1953,In_63,In_85);
or U1954 (N_1954,In_462,In_784);
and U1955 (N_1955,In_999,In_360);
xor U1956 (N_1956,In_320,In_810);
nand U1957 (N_1957,In_660,In_740);
or U1958 (N_1958,In_393,In_444);
xor U1959 (N_1959,In_343,In_204);
or U1960 (N_1960,In_718,In_979);
xnor U1961 (N_1961,In_906,In_772);
or U1962 (N_1962,In_510,In_86);
and U1963 (N_1963,In_835,In_602);
nor U1964 (N_1964,In_403,In_130);
and U1965 (N_1965,In_155,In_514);
nor U1966 (N_1966,In_715,In_270);
nor U1967 (N_1967,In_651,In_976);
nor U1968 (N_1968,In_772,In_508);
nand U1969 (N_1969,In_359,In_620);
nor U1970 (N_1970,In_833,In_896);
nor U1971 (N_1971,In_928,In_851);
nand U1972 (N_1972,In_340,In_114);
and U1973 (N_1973,In_117,In_337);
or U1974 (N_1974,In_206,In_468);
or U1975 (N_1975,In_355,In_547);
nor U1976 (N_1976,In_110,In_881);
or U1977 (N_1977,In_551,In_930);
or U1978 (N_1978,In_686,In_857);
nand U1979 (N_1979,In_117,In_746);
and U1980 (N_1980,In_200,In_357);
or U1981 (N_1981,In_537,In_845);
and U1982 (N_1982,In_258,In_620);
nor U1983 (N_1983,In_275,In_911);
nand U1984 (N_1984,In_307,In_893);
or U1985 (N_1985,In_258,In_653);
or U1986 (N_1986,In_181,In_191);
nand U1987 (N_1987,In_297,In_230);
nand U1988 (N_1988,In_698,In_323);
nor U1989 (N_1989,In_224,In_51);
nand U1990 (N_1990,In_455,In_606);
nor U1991 (N_1991,In_456,In_860);
or U1992 (N_1992,In_862,In_71);
xor U1993 (N_1993,In_53,In_259);
and U1994 (N_1994,In_725,In_596);
and U1995 (N_1995,In_657,In_70);
or U1996 (N_1996,In_860,In_626);
and U1997 (N_1997,In_97,In_321);
nand U1998 (N_1998,In_691,In_83);
nor U1999 (N_1999,In_629,In_613);
nand U2000 (N_2000,In_824,In_310);
nand U2001 (N_2001,In_533,In_983);
nand U2002 (N_2002,In_782,In_281);
nor U2003 (N_2003,In_786,In_172);
and U2004 (N_2004,In_898,In_679);
and U2005 (N_2005,In_137,In_971);
and U2006 (N_2006,In_960,In_806);
and U2007 (N_2007,In_757,In_545);
and U2008 (N_2008,In_25,In_743);
and U2009 (N_2009,In_926,In_890);
nand U2010 (N_2010,In_894,In_167);
nor U2011 (N_2011,In_493,In_577);
and U2012 (N_2012,In_621,In_568);
nand U2013 (N_2013,In_52,In_218);
nor U2014 (N_2014,In_89,In_399);
and U2015 (N_2015,In_594,In_108);
nand U2016 (N_2016,In_545,In_252);
or U2017 (N_2017,In_866,In_408);
nand U2018 (N_2018,In_11,In_819);
or U2019 (N_2019,In_348,In_708);
nor U2020 (N_2020,In_488,In_241);
or U2021 (N_2021,In_564,In_164);
and U2022 (N_2022,In_128,In_715);
nand U2023 (N_2023,In_187,In_949);
nor U2024 (N_2024,In_976,In_411);
or U2025 (N_2025,In_50,In_171);
nor U2026 (N_2026,In_783,In_481);
nor U2027 (N_2027,In_509,In_388);
and U2028 (N_2028,In_32,In_392);
nand U2029 (N_2029,In_109,In_843);
or U2030 (N_2030,In_425,In_761);
or U2031 (N_2031,In_97,In_693);
and U2032 (N_2032,In_583,In_896);
or U2033 (N_2033,In_640,In_273);
xor U2034 (N_2034,In_488,In_855);
nand U2035 (N_2035,In_206,In_569);
nand U2036 (N_2036,In_773,In_573);
and U2037 (N_2037,In_363,In_352);
nand U2038 (N_2038,In_326,In_773);
nand U2039 (N_2039,In_52,In_119);
nand U2040 (N_2040,In_146,In_333);
or U2041 (N_2041,In_345,In_913);
nand U2042 (N_2042,In_684,In_917);
or U2043 (N_2043,In_91,In_579);
nand U2044 (N_2044,In_700,In_951);
or U2045 (N_2045,In_417,In_642);
nand U2046 (N_2046,In_117,In_634);
nor U2047 (N_2047,In_424,In_763);
or U2048 (N_2048,In_936,In_760);
nand U2049 (N_2049,In_61,In_367);
and U2050 (N_2050,In_473,In_292);
or U2051 (N_2051,In_778,In_454);
nand U2052 (N_2052,In_304,In_101);
xor U2053 (N_2053,In_652,In_744);
nand U2054 (N_2054,In_263,In_319);
nand U2055 (N_2055,In_132,In_890);
nor U2056 (N_2056,In_915,In_110);
nand U2057 (N_2057,In_766,In_313);
and U2058 (N_2058,In_804,In_636);
and U2059 (N_2059,In_558,In_313);
and U2060 (N_2060,In_695,In_484);
or U2061 (N_2061,In_727,In_69);
xnor U2062 (N_2062,In_135,In_888);
nand U2063 (N_2063,In_853,In_247);
nor U2064 (N_2064,In_435,In_199);
nand U2065 (N_2065,In_777,In_972);
xnor U2066 (N_2066,In_407,In_890);
nand U2067 (N_2067,In_555,In_980);
or U2068 (N_2068,In_678,In_366);
and U2069 (N_2069,In_70,In_389);
and U2070 (N_2070,In_786,In_665);
and U2071 (N_2071,In_242,In_303);
nor U2072 (N_2072,In_729,In_702);
nand U2073 (N_2073,In_662,In_83);
nor U2074 (N_2074,In_476,In_261);
or U2075 (N_2075,In_739,In_805);
nand U2076 (N_2076,In_317,In_146);
nand U2077 (N_2077,In_381,In_952);
or U2078 (N_2078,In_914,In_168);
and U2079 (N_2079,In_322,In_855);
or U2080 (N_2080,In_835,In_538);
nand U2081 (N_2081,In_465,In_27);
nor U2082 (N_2082,In_623,In_902);
nand U2083 (N_2083,In_443,In_683);
nand U2084 (N_2084,In_797,In_426);
nand U2085 (N_2085,In_143,In_514);
xor U2086 (N_2086,In_313,In_670);
nand U2087 (N_2087,In_618,In_620);
xor U2088 (N_2088,In_976,In_824);
nand U2089 (N_2089,In_266,In_155);
nor U2090 (N_2090,In_226,In_35);
nor U2091 (N_2091,In_945,In_332);
nand U2092 (N_2092,In_413,In_51);
nand U2093 (N_2093,In_63,In_632);
and U2094 (N_2094,In_568,In_81);
and U2095 (N_2095,In_218,In_511);
nor U2096 (N_2096,In_805,In_815);
or U2097 (N_2097,In_823,In_612);
and U2098 (N_2098,In_769,In_798);
or U2099 (N_2099,In_836,In_105);
nand U2100 (N_2100,In_276,In_462);
or U2101 (N_2101,In_208,In_840);
and U2102 (N_2102,In_559,In_299);
or U2103 (N_2103,In_495,In_370);
or U2104 (N_2104,In_741,In_25);
nor U2105 (N_2105,In_726,In_467);
nor U2106 (N_2106,In_31,In_779);
and U2107 (N_2107,In_177,In_818);
and U2108 (N_2108,In_116,In_7);
nand U2109 (N_2109,In_370,In_313);
nand U2110 (N_2110,In_900,In_862);
and U2111 (N_2111,In_181,In_11);
and U2112 (N_2112,In_275,In_69);
nand U2113 (N_2113,In_990,In_349);
nor U2114 (N_2114,In_122,In_616);
or U2115 (N_2115,In_571,In_832);
nand U2116 (N_2116,In_205,In_815);
nand U2117 (N_2117,In_348,In_211);
nand U2118 (N_2118,In_764,In_626);
or U2119 (N_2119,In_390,In_770);
and U2120 (N_2120,In_700,In_941);
or U2121 (N_2121,In_790,In_7);
nor U2122 (N_2122,In_45,In_811);
and U2123 (N_2123,In_148,In_127);
or U2124 (N_2124,In_7,In_277);
or U2125 (N_2125,In_680,In_427);
xor U2126 (N_2126,In_507,In_915);
xnor U2127 (N_2127,In_167,In_250);
or U2128 (N_2128,In_576,In_718);
nor U2129 (N_2129,In_154,In_940);
nor U2130 (N_2130,In_68,In_239);
and U2131 (N_2131,In_628,In_552);
nand U2132 (N_2132,In_573,In_859);
and U2133 (N_2133,In_501,In_554);
nor U2134 (N_2134,In_984,In_396);
nand U2135 (N_2135,In_534,In_357);
or U2136 (N_2136,In_280,In_328);
and U2137 (N_2137,In_651,In_222);
nand U2138 (N_2138,In_902,In_3);
or U2139 (N_2139,In_913,In_24);
or U2140 (N_2140,In_142,In_966);
nand U2141 (N_2141,In_310,In_990);
and U2142 (N_2142,In_815,In_467);
nand U2143 (N_2143,In_218,In_468);
nand U2144 (N_2144,In_74,In_492);
nor U2145 (N_2145,In_629,In_102);
or U2146 (N_2146,In_655,In_953);
xor U2147 (N_2147,In_85,In_410);
and U2148 (N_2148,In_434,In_780);
nand U2149 (N_2149,In_190,In_514);
or U2150 (N_2150,In_442,In_408);
and U2151 (N_2151,In_399,In_453);
and U2152 (N_2152,In_208,In_328);
and U2153 (N_2153,In_126,In_324);
and U2154 (N_2154,In_247,In_740);
and U2155 (N_2155,In_653,In_240);
or U2156 (N_2156,In_614,In_935);
or U2157 (N_2157,In_382,In_822);
or U2158 (N_2158,In_841,In_727);
nand U2159 (N_2159,In_528,In_467);
or U2160 (N_2160,In_934,In_540);
nor U2161 (N_2161,In_743,In_376);
nor U2162 (N_2162,In_44,In_302);
nor U2163 (N_2163,In_66,In_24);
and U2164 (N_2164,In_41,In_938);
nor U2165 (N_2165,In_15,In_946);
xnor U2166 (N_2166,In_580,In_470);
and U2167 (N_2167,In_164,In_173);
nor U2168 (N_2168,In_160,In_106);
and U2169 (N_2169,In_594,In_267);
nor U2170 (N_2170,In_965,In_714);
nor U2171 (N_2171,In_970,In_278);
nand U2172 (N_2172,In_354,In_6);
and U2173 (N_2173,In_546,In_443);
nand U2174 (N_2174,In_387,In_773);
and U2175 (N_2175,In_220,In_627);
nor U2176 (N_2176,In_463,In_80);
nor U2177 (N_2177,In_285,In_721);
or U2178 (N_2178,In_838,In_945);
nor U2179 (N_2179,In_272,In_794);
or U2180 (N_2180,In_268,In_701);
or U2181 (N_2181,In_821,In_205);
or U2182 (N_2182,In_0,In_496);
and U2183 (N_2183,In_611,In_650);
or U2184 (N_2184,In_745,In_501);
and U2185 (N_2185,In_221,In_438);
nand U2186 (N_2186,In_242,In_698);
nand U2187 (N_2187,In_172,In_168);
and U2188 (N_2188,In_521,In_180);
or U2189 (N_2189,In_368,In_327);
or U2190 (N_2190,In_545,In_421);
nor U2191 (N_2191,In_709,In_551);
nor U2192 (N_2192,In_97,In_731);
xnor U2193 (N_2193,In_870,In_241);
xnor U2194 (N_2194,In_161,In_672);
nand U2195 (N_2195,In_389,In_695);
nand U2196 (N_2196,In_418,In_54);
xnor U2197 (N_2197,In_179,In_781);
nand U2198 (N_2198,In_957,In_200);
xnor U2199 (N_2199,In_512,In_189);
and U2200 (N_2200,In_679,In_56);
nor U2201 (N_2201,In_164,In_952);
xnor U2202 (N_2202,In_491,In_847);
and U2203 (N_2203,In_835,In_276);
nor U2204 (N_2204,In_122,In_328);
or U2205 (N_2205,In_658,In_899);
nor U2206 (N_2206,In_346,In_853);
nand U2207 (N_2207,In_412,In_694);
and U2208 (N_2208,In_653,In_458);
nand U2209 (N_2209,In_95,In_630);
and U2210 (N_2210,In_974,In_270);
and U2211 (N_2211,In_824,In_563);
nand U2212 (N_2212,In_986,In_437);
or U2213 (N_2213,In_872,In_103);
nor U2214 (N_2214,In_374,In_785);
nand U2215 (N_2215,In_388,In_796);
or U2216 (N_2216,In_56,In_559);
xnor U2217 (N_2217,In_320,In_197);
xnor U2218 (N_2218,In_262,In_881);
nand U2219 (N_2219,In_156,In_462);
xnor U2220 (N_2220,In_198,In_273);
and U2221 (N_2221,In_905,In_335);
or U2222 (N_2222,In_563,In_137);
and U2223 (N_2223,In_473,In_554);
or U2224 (N_2224,In_588,In_411);
and U2225 (N_2225,In_62,In_98);
nand U2226 (N_2226,In_960,In_16);
and U2227 (N_2227,In_282,In_795);
or U2228 (N_2228,In_100,In_318);
nor U2229 (N_2229,In_52,In_999);
or U2230 (N_2230,In_768,In_303);
or U2231 (N_2231,In_423,In_43);
and U2232 (N_2232,In_334,In_989);
nand U2233 (N_2233,In_867,In_607);
nand U2234 (N_2234,In_698,In_600);
nand U2235 (N_2235,In_622,In_93);
or U2236 (N_2236,In_382,In_80);
and U2237 (N_2237,In_744,In_489);
or U2238 (N_2238,In_293,In_620);
nor U2239 (N_2239,In_866,In_29);
and U2240 (N_2240,In_195,In_406);
nor U2241 (N_2241,In_206,In_533);
or U2242 (N_2242,In_394,In_581);
or U2243 (N_2243,In_979,In_828);
nand U2244 (N_2244,In_744,In_793);
or U2245 (N_2245,In_617,In_201);
nand U2246 (N_2246,In_918,In_51);
nor U2247 (N_2247,In_757,In_68);
and U2248 (N_2248,In_323,In_236);
nand U2249 (N_2249,In_633,In_144);
nor U2250 (N_2250,In_230,In_514);
nor U2251 (N_2251,In_982,In_939);
or U2252 (N_2252,In_320,In_171);
and U2253 (N_2253,In_970,In_708);
or U2254 (N_2254,In_407,In_211);
nor U2255 (N_2255,In_950,In_426);
and U2256 (N_2256,In_970,In_718);
nor U2257 (N_2257,In_808,In_259);
xnor U2258 (N_2258,In_103,In_207);
nor U2259 (N_2259,In_487,In_729);
or U2260 (N_2260,In_918,In_44);
or U2261 (N_2261,In_160,In_687);
or U2262 (N_2262,In_928,In_108);
nor U2263 (N_2263,In_569,In_786);
nor U2264 (N_2264,In_392,In_695);
and U2265 (N_2265,In_577,In_529);
or U2266 (N_2266,In_519,In_120);
nand U2267 (N_2267,In_254,In_893);
or U2268 (N_2268,In_858,In_844);
nor U2269 (N_2269,In_490,In_285);
xnor U2270 (N_2270,In_848,In_308);
nand U2271 (N_2271,In_19,In_872);
or U2272 (N_2272,In_646,In_488);
nand U2273 (N_2273,In_448,In_437);
xnor U2274 (N_2274,In_666,In_921);
nand U2275 (N_2275,In_303,In_424);
and U2276 (N_2276,In_11,In_949);
and U2277 (N_2277,In_923,In_192);
or U2278 (N_2278,In_518,In_449);
and U2279 (N_2279,In_509,In_934);
xor U2280 (N_2280,In_776,In_816);
nand U2281 (N_2281,In_134,In_342);
or U2282 (N_2282,In_837,In_83);
or U2283 (N_2283,In_778,In_721);
or U2284 (N_2284,In_177,In_949);
or U2285 (N_2285,In_264,In_760);
nand U2286 (N_2286,In_364,In_227);
or U2287 (N_2287,In_821,In_648);
nand U2288 (N_2288,In_323,In_268);
nor U2289 (N_2289,In_130,In_498);
nor U2290 (N_2290,In_726,In_901);
and U2291 (N_2291,In_245,In_300);
or U2292 (N_2292,In_103,In_574);
and U2293 (N_2293,In_283,In_368);
and U2294 (N_2294,In_831,In_457);
and U2295 (N_2295,In_175,In_407);
xor U2296 (N_2296,In_62,In_288);
nand U2297 (N_2297,In_297,In_618);
nand U2298 (N_2298,In_683,In_743);
and U2299 (N_2299,In_369,In_155);
nor U2300 (N_2300,In_518,In_54);
or U2301 (N_2301,In_175,In_242);
nor U2302 (N_2302,In_689,In_116);
nand U2303 (N_2303,In_591,In_239);
and U2304 (N_2304,In_476,In_145);
or U2305 (N_2305,In_791,In_157);
nand U2306 (N_2306,In_448,In_60);
or U2307 (N_2307,In_80,In_766);
nor U2308 (N_2308,In_343,In_475);
or U2309 (N_2309,In_51,In_621);
and U2310 (N_2310,In_559,In_783);
nor U2311 (N_2311,In_631,In_771);
or U2312 (N_2312,In_634,In_547);
and U2313 (N_2313,In_30,In_206);
nor U2314 (N_2314,In_942,In_0);
nand U2315 (N_2315,In_354,In_359);
xnor U2316 (N_2316,In_60,In_315);
xnor U2317 (N_2317,In_265,In_499);
nor U2318 (N_2318,In_850,In_834);
and U2319 (N_2319,In_699,In_36);
and U2320 (N_2320,In_798,In_862);
xor U2321 (N_2321,In_130,In_142);
and U2322 (N_2322,In_584,In_867);
or U2323 (N_2323,In_730,In_619);
and U2324 (N_2324,In_271,In_82);
and U2325 (N_2325,In_274,In_570);
and U2326 (N_2326,In_72,In_245);
nand U2327 (N_2327,In_298,In_166);
and U2328 (N_2328,In_549,In_538);
nor U2329 (N_2329,In_854,In_270);
nand U2330 (N_2330,In_484,In_976);
nor U2331 (N_2331,In_675,In_554);
and U2332 (N_2332,In_96,In_269);
nor U2333 (N_2333,In_872,In_711);
xnor U2334 (N_2334,In_726,In_165);
nand U2335 (N_2335,In_50,In_665);
or U2336 (N_2336,In_904,In_622);
and U2337 (N_2337,In_14,In_3);
xnor U2338 (N_2338,In_941,In_431);
nand U2339 (N_2339,In_30,In_755);
nand U2340 (N_2340,In_102,In_324);
or U2341 (N_2341,In_418,In_218);
and U2342 (N_2342,In_929,In_995);
and U2343 (N_2343,In_557,In_23);
and U2344 (N_2344,In_371,In_407);
and U2345 (N_2345,In_233,In_86);
nand U2346 (N_2346,In_782,In_104);
and U2347 (N_2347,In_687,In_701);
nor U2348 (N_2348,In_745,In_538);
nor U2349 (N_2349,In_563,In_981);
nand U2350 (N_2350,In_921,In_580);
nor U2351 (N_2351,In_327,In_446);
or U2352 (N_2352,In_392,In_906);
or U2353 (N_2353,In_998,In_471);
or U2354 (N_2354,In_852,In_207);
nand U2355 (N_2355,In_718,In_409);
or U2356 (N_2356,In_969,In_541);
xnor U2357 (N_2357,In_931,In_560);
nand U2358 (N_2358,In_493,In_970);
xnor U2359 (N_2359,In_803,In_493);
or U2360 (N_2360,In_841,In_425);
nor U2361 (N_2361,In_341,In_346);
or U2362 (N_2362,In_136,In_121);
nand U2363 (N_2363,In_217,In_855);
nor U2364 (N_2364,In_508,In_511);
nor U2365 (N_2365,In_207,In_393);
or U2366 (N_2366,In_828,In_6);
nand U2367 (N_2367,In_415,In_106);
nor U2368 (N_2368,In_681,In_80);
nand U2369 (N_2369,In_793,In_266);
nor U2370 (N_2370,In_847,In_596);
and U2371 (N_2371,In_245,In_89);
or U2372 (N_2372,In_196,In_525);
and U2373 (N_2373,In_459,In_515);
or U2374 (N_2374,In_547,In_273);
nor U2375 (N_2375,In_436,In_298);
and U2376 (N_2376,In_930,In_714);
or U2377 (N_2377,In_6,In_48);
or U2378 (N_2378,In_281,In_658);
nor U2379 (N_2379,In_137,In_184);
or U2380 (N_2380,In_907,In_531);
xnor U2381 (N_2381,In_467,In_650);
nand U2382 (N_2382,In_269,In_674);
or U2383 (N_2383,In_983,In_786);
or U2384 (N_2384,In_105,In_786);
xor U2385 (N_2385,In_232,In_521);
nand U2386 (N_2386,In_243,In_136);
nor U2387 (N_2387,In_686,In_723);
or U2388 (N_2388,In_814,In_257);
nor U2389 (N_2389,In_212,In_148);
nor U2390 (N_2390,In_441,In_926);
or U2391 (N_2391,In_538,In_251);
and U2392 (N_2392,In_792,In_667);
or U2393 (N_2393,In_542,In_644);
nor U2394 (N_2394,In_338,In_0);
and U2395 (N_2395,In_974,In_273);
and U2396 (N_2396,In_926,In_521);
or U2397 (N_2397,In_860,In_506);
xor U2398 (N_2398,In_340,In_888);
nand U2399 (N_2399,In_42,In_175);
nand U2400 (N_2400,In_405,In_235);
or U2401 (N_2401,In_786,In_186);
or U2402 (N_2402,In_819,In_728);
or U2403 (N_2403,In_682,In_566);
xnor U2404 (N_2404,In_279,In_656);
nand U2405 (N_2405,In_242,In_187);
nand U2406 (N_2406,In_9,In_247);
nand U2407 (N_2407,In_905,In_540);
or U2408 (N_2408,In_269,In_309);
or U2409 (N_2409,In_592,In_476);
xnor U2410 (N_2410,In_290,In_830);
nand U2411 (N_2411,In_313,In_199);
nor U2412 (N_2412,In_785,In_32);
nand U2413 (N_2413,In_729,In_641);
nand U2414 (N_2414,In_821,In_492);
nor U2415 (N_2415,In_816,In_41);
nor U2416 (N_2416,In_50,In_60);
or U2417 (N_2417,In_93,In_713);
or U2418 (N_2418,In_844,In_467);
nand U2419 (N_2419,In_355,In_489);
and U2420 (N_2420,In_565,In_617);
nand U2421 (N_2421,In_677,In_766);
and U2422 (N_2422,In_279,In_77);
nand U2423 (N_2423,In_340,In_596);
nand U2424 (N_2424,In_704,In_845);
nand U2425 (N_2425,In_116,In_600);
nor U2426 (N_2426,In_204,In_374);
nor U2427 (N_2427,In_341,In_442);
nor U2428 (N_2428,In_775,In_891);
xnor U2429 (N_2429,In_114,In_698);
xnor U2430 (N_2430,In_115,In_800);
nor U2431 (N_2431,In_895,In_292);
nand U2432 (N_2432,In_716,In_101);
nor U2433 (N_2433,In_603,In_372);
nand U2434 (N_2434,In_261,In_206);
nor U2435 (N_2435,In_967,In_451);
or U2436 (N_2436,In_881,In_861);
or U2437 (N_2437,In_823,In_659);
and U2438 (N_2438,In_596,In_758);
nand U2439 (N_2439,In_869,In_980);
or U2440 (N_2440,In_560,In_346);
nand U2441 (N_2441,In_560,In_286);
or U2442 (N_2442,In_914,In_141);
nor U2443 (N_2443,In_159,In_985);
nand U2444 (N_2444,In_650,In_276);
or U2445 (N_2445,In_858,In_154);
nor U2446 (N_2446,In_796,In_810);
or U2447 (N_2447,In_694,In_189);
and U2448 (N_2448,In_193,In_452);
nor U2449 (N_2449,In_941,In_949);
or U2450 (N_2450,In_531,In_453);
and U2451 (N_2451,In_305,In_507);
nor U2452 (N_2452,In_364,In_780);
nor U2453 (N_2453,In_490,In_456);
nor U2454 (N_2454,In_825,In_54);
nand U2455 (N_2455,In_979,In_798);
and U2456 (N_2456,In_709,In_455);
or U2457 (N_2457,In_954,In_532);
and U2458 (N_2458,In_940,In_392);
nand U2459 (N_2459,In_416,In_831);
and U2460 (N_2460,In_85,In_901);
xor U2461 (N_2461,In_478,In_917);
or U2462 (N_2462,In_811,In_637);
nand U2463 (N_2463,In_363,In_71);
and U2464 (N_2464,In_103,In_655);
and U2465 (N_2465,In_934,In_753);
nand U2466 (N_2466,In_862,In_601);
xnor U2467 (N_2467,In_650,In_832);
xnor U2468 (N_2468,In_199,In_615);
or U2469 (N_2469,In_628,In_112);
xor U2470 (N_2470,In_164,In_813);
and U2471 (N_2471,In_889,In_797);
nand U2472 (N_2472,In_733,In_908);
nand U2473 (N_2473,In_182,In_496);
or U2474 (N_2474,In_724,In_260);
or U2475 (N_2475,In_164,In_510);
nand U2476 (N_2476,In_717,In_50);
xor U2477 (N_2477,In_349,In_421);
or U2478 (N_2478,In_45,In_611);
nor U2479 (N_2479,In_293,In_657);
and U2480 (N_2480,In_452,In_690);
and U2481 (N_2481,In_733,In_868);
and U2482 (N_2482,In_211,In_769);
nand U2483 (N_2483,In_926,In_931);
or U2484 (N_2484,In_326,In_745);
and U2485 (N_2485,In_667,In_725);
nor U2486 (N_2486,In_582,In_318);
or U2487 (N_2487,In_35,In_818);
and U2488 (N_2488,In_116,In_95);
and U2489 (N_2489,In_693,In_488);
or U2490 (N_2490,In_378,In_961);
or U2491 (N_2491,In_395,In_632);
nand U2492 (N_2492,In_948,In_175);
and U2493 (N_2493,In_150,In_675);
or U2494 (N_2494,In_704,In_796);
and U2495 (N_2495,In_533,In_329);
nand U2496 (N_2496,In_370,In_532);
nor U2497 (N_2497,In_764,In_604);
or U2498 (N_2498,In_822,In_30);
and U2499 (N_2499,In_54,In_463);
or U2500 (N_2500,In_414,In_952);
nor U2501 (N_2501,In_363,In_816);
or U2502 (N_2502,In_687,In_142);
nand U2503 (N_2503,In_236,In_945);
nor U2504 (N_2504,In_553,In_122);
or U2505 (N_2505,In_669,In_975);
xnor U2506 (N_2506,In_617,In_438);
or U2507 (N_2507,In_289,In_249);
and U2508 (N_2508,In_796,In_611);
and U2509 (N_2509,In_688,In_192);
and U2510 (N_2510,In_41,In_267);
nand U2511 (N_2511,In_391,In_643);
xnor U2512 (N_2512,In_860,In_697);
nand U2513 (N_2513,In_142,In_772);
and U2514 (N_2514,In_678,In_914);
nor U2515 (N_2515,In_357,In_207);
and U2516 (N_2516,In_69,In_460);
nor U2517 (N_2517,In_289,In_14);
nand U2518 (N_2518,In_853,In_17);
xnor U2519 (N_2519,In_386,In_694);
nand U2520 (N_2520,In_469,In_78);
nor U2521 (N_2521,In_615,In_45);
nand U2522 (N_2522,In_545,In_679);
and U2523 (N_2523,In_300,In_573);
or U2524 (N_2524,In_687,In_562);
or U2525 (N_2525,In_283,In_220);
nor U2526 (N_2526,In_291,In_68);
or U2527 (N_2527,In_770,In_465);
nand U2528 (N_2528,In_226,In_466);
and U2529 (N_2529,In_125,In_389);
or U2530 (N_2530,In_819,In_637);
nor U2531 (N_2531,In_748,In_575);
nor U2532 (N_2532,In_677,In_558);
nor U2533 (N_2533,In_769,In_322);
nand U2534 (N_2534,In_304,In_6);
xnor U2535 (N_2535,In_547,In_265);
nor U2536 (N_2536,In_898,In_781);
nand U2537 (N_2537,In_368,In_570);
nor U2538 (N_2538,In_952,In_940);
nor U2539 (N_2539,In_193,In_171);
and U2540 (N_2540,In_594,In_959);
xor U2541 (N_2541,In_420,In_959);
nor U2542 (N_2542,In_592,In_678);
nor U2543 (N_2543,In_724,In_717);
and U2544 (N_2544,In_411,In_287);
or U2545 (N_2545,In_502,In_214);
or U2546 (N_2546,In_484,In_630);
xor U2547 (N_2547,In_505,In_625);
and U2548 (N_2548,In_526,In_435);
and U2549 (N_2549,In_786,In_428);
nor U2550 (N_2550,In_618,In_938);
nand U2551 (N_2551,In_686,In_399);
and U2552 (N_2552,In_539,In_183);
xor U2553 (N_2553,In_786,In_319);
xor U2554 (N_2554,In_120,In_1);
and U2555 (N_2555,In_936,In_392);
nor U2556 (N_2556,In_660,In_196);
nand U2557 (N_2557,In_609,In_765);
nor U2558 (N_2558,In_323,In_465);
or U2559 (N_2559,In_643,In_718);
nand U2560 (N_2560,In_445,In_151);
and U2561 (N_2561,In_824,In_848);
or U2562 (N_2562,In_787,In_476);
and U2563 (N_2563,In_92,In_718);
and U2564 (N_2564,In_919,In_959);
and U2565 (N_2565,In_311,In_550);
nor U2566 (N_2566,In_484,In_194);
nand U2567 (N_2567,In_801,In_941);
or U2568 (N_2568,In_415,In_456);
and U2569 (N_2569,In_178,In_393);
nand U2570 (N_2570,In_854,In_27);
nand U2571 (N_2571,In_4,In_694);
xnor U2572 (N_2572,In_408,In_510);
and U2573 (N_2573,In_299,In_913);
nand U2574 (N_2574,In_246,In_755);
and U2575 (N_2575,In_938,In_451);
and U2576 (N_2576,In_698,In_472);
nor U2577 (N_2577,In_883,In_775);
nand U2578 (N_2578,In_857,In_486);
or U2579 (N_2579,In_649,In_456);
or U2580 (N_2580,In_410,In_905);
nor U2581 (N_2581,In_496,In_332);
or U2582 (N_2582,In_483,In_171);
or U2583 (N_2583,In_654,In_591);
or U2584 (N_2584,In_470,In_880);
nor U2585 (N_2585,In_850,In_198);
or U2586 (N_2586,In_198,In_939);
and U2587 (N_2587,In_95,In_104);
or U2588 (N_2588,In_560,In_820);
nor U2589 (N_2589,In_923,In_44);
or U2590 (N_2590,In_428,In_421);
or U2591 (N_2591,In_7,In_596);
or U2592 (N_2592,In_566,In_175);
nand U2593 (N_2593,In_146,In_651);
or U2594 (N_2594,In_801,In_382);
nand U2595 (N_2595,In_968,In_92);
nand U2596 (N_2596,In_532,In_219);
nand U2597 (N_2597,In_253,In_336);
or U2598 (N_2598,In_647,In_431);
nor U2599 (N_2599,In_44,In_269);
and U2600 (N_2600,In_249,In_70);
nand U2601 (N_2601,In_979,In_457);
xor U2602 (N_2602,In_950,In_37);
and U2603 (N_2603,In_769,In_178);
xor U2604 (N_2604,In_53,In_774);
nand U2605 (N_2605,In_758,In_650);
and U2606 (N_2606,In_923,In_672);
xor U2607 (N_2607,In_488,In_475);
nor U2608 (N_2608,In_428,In_361);
and U2609 (N_2609,In_293,In_806);
or U2610 (N_2610,In_525,In_724);
and U2611 (N_2611,In_991,In_127);
nor U2612 (N_2612,In_122,In_971);
nand U2613 (N_2613,In_462,In_976);
xor U2614 (N_2614,In_646,In_798);
or U2615 (N_2615,In_524,In_311);
and U2616 (N_2616,In_576,In_939);
xor U2617 (N_2617,In_390,In_983);
nand U2618 (N_2618,In_315,In_74);
nor U2619 (N_2619,In_222,In_889);
and U2620 (N_2620,In_84,In_976);
or U2621 (N_2621,In_419,In_517);
or U2622 (N_2622,In_56,In_902);
or U2623 (N_2623,In_575,In_751);
or U2624 (N_2624,In_58,In_528);
nor U2625 (N_2625,In_389,In_357);
nand U2626 (N_2626,In_674,In_734);
nor U2627 (N_2627,In_557,In_784);
nand U2628 (N_2628,In_416,In_393);
and U2629 (N_2629,In_225,In_100);
nor U2630 (N_2630,In_245,In_624);
xnor U2631 (N_2631,In_453,In_190);
and U2632 (N_2632,In_899,In_571);
and U2633 (N_2633,In_808,In_709);
and U2634 (N_2634,In_741,In_808);
nand U2635 (N_2635,In_485,In_630);
xor U2636 (N_2636,In_162,In_781);
and U2637 (N_2637,In_452,In_196);
nor U2638 (N_2638,In_853,In_817);
nand U2639 (N_2639,In_368,In_671);
and U2640 (N_2640,In_311,In_939);
or U2641 (N_2641,In_271,In_923);
or U2642 (N_2642,In_538,In_31);
and U2643 (N_2643,In_954,In_544);
or U2644 (N_2644,In_612,In_407);
nor U2645 (N_2645,In_545,In_459);
or U2646 (N_2646,In_146,In_857);
or U2647 (N_2647,In_138,In_392);
and U2648 (N_2648,In_502,In_396);
or U2649 (N_2649,In_472,In_558);
or U2650 (N_2650,In_827,In_639);
and U2651 (N_2651,In_270,In_889);
nand U2652 (N_2652,In_915,In_843);
or U2653 (N_2653,In_579,In_304);
or U2654 (N_2654,In_216,In_847);
nand U2655 (N_2655,In_933,In_117);
nand U2656 (N_2656,In_822,In_837);
or U2657 (N_2657,In_358,In_576);
and U2658 (N_2658,In_781,In_746);
or U2659 (N_2659,In_811,In_246);
nand U2660 (N_2660,In_470,In_256);
and U2661 (N_2661,In_764,In_271);
or U2662 (N_2662,In_383,In_437);
xor U2663 (N_2663,In_29,In_957);
nand U2664 (N_2664,In_722,In_818);
or U2665 (N_2665,In_756,In_899);
or U2666 (N_2666,In_563,In_292);
nand U2667 (N_2667,In_922,In_272);
or U2668 (N_2668,In_552,In_143);
and U2669 (N_2669,In_45,In_833);
xor U2670 (N_2670,In_598,In_554);
or U2671 (N_2671,In_983,In_632);
and U2672 (N_2672,In_44,In_47);
nor U2673 (N_2673,In_378,In_751);
or U2674 (N_2674,In_26,In_851);
and U2675 (N_2675,In_546,In_914);
nand U2676 (N_2676,In_499,In_117);
nand U2677 (N_2677,In_656,In_411);
or U2678 (N_2678,In_249,In_541);
or U2679 (N_2679,In_947,In_233);
and U2680 (N_2680,In_805,In_880);
or U2681 (N_2681,In_584,In_233);
or U2682 (N_2682,In_229,In_31);
and U2683 (N_2683,In_381,In_274);
and U2684 (N_2684,In_817,In_858);
nor U2685 (N_2685,In_491,In_138);
xnor U2686 (N_2686,In_611,In_315);
nor U2687 (N_2687,In_994,In_59);
nor U2688 (N_2688,In_880,In_658);
and U2689 (N_2689,In_767,In_326);
nand U2690 (N_2690,In_346,In_933);
xnor U2691 (N_2691,In_581,In_782);
or U2692 (N_2692,In_212,In_541);
or U2693 (N_2693,In_838,In_518);
nor U2694 (N_2694,In_726,In_775);
nand U2695 (N_2695,In_25,In_873);
and U2696 (N_2696,In_102,In_311);
nor U2697 (N_2697,In_415,In_514);
and U2698 (N_2698,In_277,In_226);
nand U2699 (N_2699,In_806,In_233);
or U2700 (N_2700,In_970,In_233);
or U2701 (N_2701,In_336,In_650);
xnor U2702 (N_2702,In_210,In_819);
nor U2703 (N_2703,In_670,In_58);
and U2704 (N_2704,In_398,In_488);
or U2705 (N_2705,In_704,In_393);
or U2706 (N_2706,In_322,In_469);
nand U2707 (N_2707,In_362,In_296);
nand U2708 (N_2708,In_388,In_278);
nand U2709 (N_2709,In_311,In_154);
or U2710 (N_2710,In_164,In_590);
nand U2711 (N_2711,In_345,In_723);
nand U2712 (N_2712,In_306,In_960);
nor U2713 (N_2713,In_876,In_573);
nor U2714 (N_2714,In_300,In_885);
or U2715 (N_2715,In_200,In_725);
nand U2716 (N_2716,In_838,In_678);
or U2717 (N_2717,In_596,In_946);
or U2718 (N_2718,In_333,In_461);
and U2719 (N_2719,In_910,In_927);
and U2720 (N_2720,In_501,In_278);
nand U2721 (N_2721,In_868,In_689);
xnor U2722 (N_2722,In_433,In_317);
and U2723 (N_2723,In_756,In_969);
or U2724 (N_2724,In_403,In_887);
or U2725 (N_2725,In_981,In_970);
and U2726 (N_2726,In_961,In_607);
nand U2727 (N_2727,In_618,In_977);
nor U2728 (N_2728,In_537,In_186);
or U2729 (N_2729,In_950,In_210);
nand U2730 (N_2730,In_295,In_614);
nand U2731 (N_2731,In_274,In_4);
nor U2732 (N_2732,In_246,In_209);
nand U2733 (N_2733,In_819,In_853);
and U2734 (N_2734,In_582,In_941);
or U2735 (N_2735,In_571,In_369);
or U2736 (N_2736,In_350,In_231);
nor U2737 (N_2737,In_365,In_693);
nand U2738 (N_2738,In_396,In_873);
and U2739 (N_2739,In_555,In_199);
or U2740 (N_2740,In_133,In_882);
nand U2741 (N_2741,In_460,In_621);
nand U2742 (N_2742,In_161,In_38);
and U2743 (N_2743,In_306,In_379);
nor U2744 (N_2744,In_18,In_111);
and U2745 (N_2745,In_516,In_463);
xnor U2746 (N_2746,In_538,In_701);
or U2747 (N_2747,In_18,In_359);
xnor U2748 (N_2748,In_569,In_293);
or U2749 (N_2749,In_526,In_44);
nand U2750 (N_2750,In_984,In_90);
nor U2751 (N_2751,In_553,In_13);
nor U2752 (N_2752,In_603,In_373);
and U2753 (N_2753,In_942,In_105);
nand U2754 (N_2754,In_520,In_677);
nand U2755 (N_2755,In_525,In_5);
nand U2756 (N_2756,In_16,In_364);
nor U2757 (N_2757,In_612,In_862);
and U2758 (N_2758,In_892,In_10);
nand U2759 (N_2759,In_937,In_975);
or U2760 (N_2760,In_447,In_445);
xor U2761 (N_2761,In_669,In_621);
nand U2762 (N_2762,In_66,In_165);
and U2763 (N_2763,In_418,In_708);
nor U2764 (N_2764,In_738,In_84);
or U2765 (N_2765,In_608,In_893);
or U2766 (N_2766,In_64,In_462);
and U2767 (N_2767,In_183,In_352);
nand U2768 (N_2768,In_567,In_580);
nand U2769 (N_2769,In_140,In_754);
or U2770 (N_2770,In_858,In_318);
nand U2771 (N_2771,In_677,In_179);
and U2772 (N_2772,In_998,In_928);
and U2773 (N_2773,In_620,In_999);
or U2774 (N_2774,In_264,In_354);
and U2775 (N_2775,In_215,In_350);
and U2776 (N_2776,In_874,In_889);
or U2777 (N_2777,In_348,In_525);
or U2778 (N_2778,In_313,In_324);
xor U2779 (N_2779,In_173,In_16);
or U2780 (N_2780,In_865,In_973);
nand U2781 (N_2781,In_409,In_542);
xor U2782 (N_2782,In_29,In_69);
nor U2783 (N_2783,In_168,In_51);
nand U2784 (N_2784,In_369,In_938);
and U2785 (N_2785,In_504,In_286);
nor U2786 (N_2786,In_992,In_624);
nand U2787 (N_2787,In_475,In_1);
nor U2788 (N_2788,In_926,In_924);
and U2789 (N_2789,In_744,In_172);
and U2790 (N_2790,In_600,In_188);
or U2791 (N_2791,In_241,In_833);
nor U2792 (N_2792,In_317,In_194);
and U2793 (N_2793,In_518,In_816);
xnor U2794 (N_2794,In_59,In_24);
nor U2795 (N_2795,In_727,In_73);
xnor U2796 (N_2796,In_964,In_756);
nor U2797 (N_2797,In_221,In_868);
nor U2798 (N_2798,In_218,In_254);
or U2799 (N_2799,In_4,In_458);
nand U2800 (N_2800,In_175,In_308);
and U2801 (N_2801,In_43,In_516);
and U2802 (N_2802,In_442,In_784);
and U2803 (N_2803,In_642,In_190);
xnor U2804 (N_2804,In_612,In_828);
or U2805 (N_2805,In_386,In_933);
and U2806 (N_2806,In_412,In_545);
nand U2807 (N_2807,In_842,In_773);
nand U2808 (N_2808,In_484,In_911);
xor U2809 (N_2809,In_69,In_955);
nand U2810 (N_2810,In_989,In_296);
or U2811 (N_2811,In_942,In_334);
xnor U2812 (N_2812,In_255,In_325);
and U2813 (N_2813,In_395,In_516);
nor U2814 (N_2814,In_982,In_739);
and U2815 (N_2815,In_124,In_444);
and U2816 (N_2816,In_733,In_96);
xnor U2817 (N_2817,In_691,In_299);
nor U2818 (N_2818,In_455,In_473);
xor U2819 (N_2819,In_739,In_477);
nor U2820 (N_2820,In_599,In_608);
and U2821 (N_2821,In_882,In_153);
nor U2822 (N_2822,In_986,In_107);
xor U2823 (N_2823,In_858,In_841);
or U2824 (N_2824,In_475,In_227);
nand U2825 (N_2825,In_700,In_12);
and U2826 (N_2826,In_230,In_517);
or U2827 (N_2827,In_551,In_386);
nand U2828 (N_2828,In_652,In_428);
nor U2829 (N_2829,In_297,In_609);
nor U2830 (N_2830,In_25,In_220);
or U2831 (N_2831,In_544,In_57);
xnor U2832 (N_2832,In_43,In_847);
xor U2833 (N_2833,In_896,In_761);
nor U2834 (N_2834,In_342,In_143);
nand U2835 (N_2835,In_164,In_143);
nor U2836 (N_2836,In_936,In_768);
nand U2837 (N_2837,In_413,In_741);
and U2838 (N_2838,In_857,In_765);
and U2839 (N_2839,In_786,In_124);
or U2840 (N_2840,In_110,In_384);
and U2841 (N_2841,In_323,In_44);
nor U2842 (N_2842,In_974,In_1);
nand U2843 (N_2843,In_630,In_850);
and U2844 (N_2844,In_943,In_589);
nor U2845 (N_2845,In_412,In_821);
and U2846 (N_2846,In_928,In_657);
nor U2847 (N_2847,In_96,In_506);
and U2848 (N_2848,In_420,In_831);
or U2849 (N_2849,In_676,In_271);
and U2850 (N_2850,In_37,In_206);
nor U2851 (N_2851,In_630,In_564);
or U2852 (N_2852,In_956,In_382);
xor U2853 (N_2853,In_646,In_288);
nor U2854 (N_2854,In_797,In_217);
nor U2855 (N_2855,In_405,In_316);
nor U2856 (N_2856,In_441,In_36);
or U2857 (N_2857,In_767,In_876);
and U2858 (N_2858,In_28,In_263);
or U2859 (N_2859,In_158,In_861);
and U2860 (N_2860,In_53,In_601);
nand U2861 (N_2861,In_348,In_297);
nor U2862 (N_2862,In_665,In_422);
xnor U2863 (N_2863,In_492,In_549);
nand U2864 (N_2864,In_583,In_684);
or U2865 (N_2865,In_189,In_335);
and U2866 (N_2866,In_16,In_487);
and U2867 (N_2867,In_185,In_424);
nor U2868 (N_2868,In_108,In_109);
nor U2869 (N_2869,In_271,In_588);
or U2870 (N_2870,In_23,In_816);
and U2871 (N_2871,In_3,In_916);
nor U2872 (N_2872,In_131,In_639);
or U2873 (N_2873,In_430,In_699);
nor U2874 (N_2874,In_962,In_548);
or U2875 (N_2875,In_844,In_776);
or U2876 (N_2876,In_78,In_720);
xor U2877 (N_2877,In_57,In_88);
nand U2878 (N_2878,In_264,In_960);
or U2879 (N_2879,In_418,In_299);
nor U2880 (N_2880,In_475,In_130);
nor U2881 (N_2881,In_284,In_632);
nand U2882 (N_2882,In_635,In_896);
and U2883 (N_2883,In_674,In_162);
and U2884 (N_2884,In_354,In_571);
nand U2885 (N_2885,In_8,In_578);
and U2886 (N_2886,In_860,In_96);
nand U2887 (N_2887,In_847,In_587);
and U2888 (N_2888,In_660,In_931);
nand U2889 (N_2889,In_539,In_695);
nor U2890 (N_2890,In_244,In_575);
and U2891 (N_2891,In_223,In_750);
and U2892 (N_2892,In_188,In_702);
and U2893 (N_2893,In_812,In_186);
and U2894 (N_2894,In_408,In_595);
nand U2895 (N_2895,In_149,In_707);
nand U2896 (N_2896,In_667,In_336);
or U2897 (N_2897,In_117,In_915);
or U2898 (N_2898,In_329,In_509);
xor U2899 (N_2899,In_407,In_596);
or U2900 (N_2900,In_139,In_180);
nor U2901 (N_2901,In_23,In_869);
or U2902 (N_2902,In_892,In_728);
nand U2903 (N_2903,In_352,In_180);
nand U2904 (N_2904,In_271,In_484);
nand U2905 (N_2905,In_251,In_82);
and U2906 (N_2906,In_849,In_313);
and U2907 (N_2907,In_432,In_213);
nor U2908 (N_2908,In_379,In_762);
or U2909 (N_2909,In_692,In_376);
nor U2910 (N_2910,In_805,In_146);
nor U2911 (N_2911,In_27,In_906);
nor U2912 (N_2912,In_124,In_909);
nor U2913 (N_2913,In_62,In_821);
and U2914 (N_2914,In_706,In_687);
nand U2915 (N_2915,In_767,In_904);
nor U2916 (N_2916,In_419,In_639);
nand U2917 (N_2917,In_753,In_279);
and U2918 (N_2918,In_894,In_636);
and U2919 (N_2919,In_346,In_125);
or U2920 (N_2920,In_982,In_508);
or U2921 (N_2921,In_869,In_139);
and U2922 (N_2922,In_777,In_880);
nor U2923 (N_2923,In_170,In_727);
nor U2924 (N_2924,In_467,In_833);
nor U2925 (N_2925,In_100,In_738);
nand U2926 (N_2926,In_269,In_130);
nor U2927 (N_2927,In_709,In_331);
or U2928 (N_2928,In_813,In_201);
or U2929 (N_2929,In_88,In_646);
or U2930 (N_2930,In_361,In_603);
and U2931 (N_2931,In_966,In_213);
nand U2932 (N_2932,In_32,In_811);
or U2933 (N_2933,In_566,In_807);
nor U2934 (N_2934,In_652,In_930);
xor U2935 (N_2935,In_618,In_676);
xnor U2936 (N_2936,In_329,In_651);
and U2937 (N_2937,In_490,In_734);
and U2938 (N_2938,In_654,In_499);
nand U2939 (N_2939,In_980,In_155);
and U2940 (N_2940,In_811,In_292);
nand U2941 (N_2941,In_4,In_968);
nor U2942 (N_2942,In_740,In_898);
xor U2943 (N_2943,In_696,In_856);
or U2944 (N_2944,In_879,In_793);
and U2945 (N_2945,In_64,In_116);
nor U2946 (N_2946,In_161,In_253);
and U2947 (N_2947,In_437,In_580);
nand U2948 (N_2948,In_576,In_907);
nand U2949 (N_2949,In_513,In_784);
or U2950 (N_2950,In_649,In_720);
or U2951 (N_2951,In_841,In_679);
or U2952 (N_2952,In_447,In_327);
and U2953 (N_2953,In_63,In_644);
nor U2954 (N_2954,In_336,In_171);
and U2955 (N_2955,In_994,In_781);
and U2956 (N_2956,In_626,In_598);
nand U2957 (N_2957,In_117,In_72);
xor U2958 (N_2958,In_578,In_171);
nand U2959 (N_2959,In_897,In_310);
nand U2960 (N_2960,In_175,In_835);
and U2961 (N_2961,In_687,In_855);
and U2962 (N_2962,In_755,In_983);
or U2963 (N_2963,In_730,In_941);
and U2964 (N_2964,In_30,In_299);
nand U2965 (N_2965,In_132,In_548);
nand U2966 (N_2966,In_856,In_978);
nand U2967 (N_2967,In_611,In_393);
nand U2968 (N_2968,In_232,In_811);
and U2969 (N_2969,In_481,In_549);
nand U2970 (N_2970,In_897,In_131);
or U2971 (N_2971,In_752,In_989);
nand U2972 (N_2972,In_797,In_737);
nor U2973 (N_2973,In_410,In_810);
or U2974 (N_2974,In_517,In_475);
or U2975 (N_2975,In_810,In_747);
nor U2976 (N_2976,In_55,In_946);
nand U2977 (N_2977,In_215,In_603);
or U2978 (N_2978,In_690,In_836);
xor U2979 (N_2979,In_136,In_240);
nor U2980 (N_2980,In_927,In_577);
or U2981 (N_2981,In_20,In_333);
nand U2982 (N_2982,In_503,In_863);
or U2983 (N_2983,In_5,In_593);
nand U2984 (N_2984,In_577,In_308);
and U2985 (N_2985,In_278,In_144);
or U2986 (N_2986,In_558,In_88);
nor U2987 (N_2987,In_543,In_139);
or U2988 (N_2988,In_765,In_540);
and U2989 (N_2989,In_923,In_553);
nor U2990 (N_2990,In_595,In_844);
or U2991 (N_2991,In_233,In_668);
nand U2992 (N_2992,In_851,In_652);
xnor U2993 (N_2993,In_83,In_275);
xnor U2994 (N_2994,In_212,In_82);
or U2995 (N_2995,In_242,In_199);
and U2996 (N_2996,In_397,In_315);
nor U2997 (N_2997,In_316,In_988);
and U2998 (N_2998,In_480,In_288);
nand U2999 (N_2999,In_265,In_99);
or U3000 (N_3000,In_819,In_940);
nand U3001 (N_3001,In_995,In_675);
xnor U3002 (N_3002,In_600,In_352);
or U3003 (N_3003,In_195,In_592);
or U3004 (N_3004,In_365,In_338);
nor U3005 (N_3005,In_343,In_938);
and U3006 (N_3006,In_859,In_846);
nand U3007 (N_3007,In_428,In_213);
or U3008 (N_3008,In_380,In_29);
nand U3009 (N_3009,In_633,In_767);
nor U3010 (N_3010,In_206,In_125);
and U3011 (N_3011,In_620,In_554);
or U3012 (N_3012,In_331,In_986);
nor U3013 (N_3013,In_764,In_236);
nor U3014 (N_3014,In_7,In_20);
and U3015 (N_3015,In_230,In_117);
or U3016 (N_3016,In_114,In_539);
and U3017 (N_3017,In_188,In_296);
nand U3018 (N_3018,In_875,In_697);
nand U3019 (N_3019,In_886,In_33);
nand U3020 (N_3020,In_405,In_731);
or U3021 (N_3021,In_779,In_42);
and U3022 (N_3022,In_835,In_785);
and U3023 (N_3023,In_489,In_741);
or U3024 (N_3024,In_572,In_96);
nand U3025 (N_3025,In_685,In_531);
nor U3026 (N_3026,In_410,In_882);
nor U3027 (N_3027,In_616,In_770);
and U3028 (N_3028,In_328,In_724);
nor U3029 (N_3029,In_622,In_596);
and U3030 (N_3030,In_179,In_586);
nor U3031 (N_3031,In_129,In_645);
and U3032 (N_3032,In_305,In_767);
or U3033 (N_3033,In_987,In_607);
nor U3034 (N_3034,In_546,In_363);
xnor U3035 (N_3035,In_42,In_34);
or U3036 (N_3036,In_513,In_659);
nand U3037 (N_3037,In_554,In_574);
or U3038 (N_3038,In_303,In_129);
nor U3039 (N_3039,In_532,In_214);
or U3040 (N_3040,In_270,In_415);
nor U3041 (N_3041,In_185,In_54);
nand U3042 (N_3042,In_558,In_98);
nor U3043 (N_3043,In_790,In_451);
and U3044 (N_3044,In_358,In_94);
nor U3045 (N_3045,In_674,In_158);
nor U3046 (N_3046,In_17,In_801);
nor U3047 (N_3047,In_582,In_702);
and U3048 (N_3048,In_623,In_501);
nor U3049 (N_3049,In_207,In_784);
nor U3050 (N_3050,In_198,In_957);
nor U3051 (N_3051,In_60,In_596);
nor U3052 (N_3052,In_585,In_121);
xor U3053 (N_3053,In_221,In_945);
or U3054 (N_3054,In_564,In_72);
and U3055 (N_3055,In_755,In_750);
and U3056 (N_3056,In_45,In_951);
or U3057 (N_3057,In_449,In_586);
nand U3058 (N_3058,In_29,In_840);
and U3059 (N_3059,In_551,In_577);
nor U3060 (N_3060,In_219,In_620);
and U3061 (N_3061,In_872,In_76);
nor U3062 (N_3062,In_311,In_234);
xnor U3063 (N_3063,In_803,In_637);
and U3064 (N_3064,In_366,In_213);
nand U3065 (N_3065,In_458,In_906);
nor U3066 (N_3066,In_676,In_484);
and U3067 (N_3067,In_25,In_544);
nor U3068 (N_3068,In_169,In_391);
or U3069 (N_3069,In_975,In_467);
nor U3070 (N_3070,In_681,In_320);
or U3071 (N_3071,In_327,In_15);
and U3072 (N_3072,In_190,In_486);
nand U3073 (N_3073,In_241,In_155);
and U3074 (N_3074,In_791,In_659);
and U3075 (N_3075,In_547,In_875);
nand U3076 (N_3076,In_245,In_728);
and U3077 (N_3077,In_574,In_248);
and U3078 (N_3078,In_664,In_626);
nand U3079 (N_3079,In_923,In_71);
nor U3080 (N_3080,In_870,In_125);
nor U3081 (N_3081,In_165,In_348);
xnor U3082 (N_3082,In_649,In_890);
nor U3083 (N_3083,In_342,In_93);
or U3084 (N_3084,In_550,In_82);
nor U3085 (N_3085,In_732,In_635);
nor U3086 (N_3086,In_564,In_569);
nor U3087 (N_3087,In_576,In_872);
nand U3088 (N_3088,In_236,In_253);
nand U3089 (N_3089,In_939,In_448);
and U3090 (N_3090,In_238,In_450);
or U3091 (N_3091,In_553,In_695);
nor U3092 (N_3092,In_702,In_742);
xnor U3093 (N_3093,In_308,In_497);
nand U3094 (N_3094,In_972,In_31);
and U3095 (N_3095,In_180,In_284);
or U3096 (N_3096,In_983,In_565);
nor U3097 (N_3097,In_750,In_358);
and U3098 (N_3098,In_899,In_366);
nand U3099 (N_3099,In_783,In_761);
nor U3100 (N_3100,In_928,In_575);
and U3101 (N_3101,In_718,In_55);
xor U3102 (N_3102,In_230,In_778);
and U3103 (N_3103,In_116,In_361);
xnor U3104 (N_3104,In_816,In_941);
nand U3105 (N_3105,In_889,In_279);
or U3106 (N_3106,In_72,In_178);
nor U3107 (N_3107,In_760,In_405);
nand U3108 (N_3108,In_555,In_793);
and U3109 (N_3109,In_49,In_749);
nand U3110 (N_3110,In_711,In_981);
nand U3111 (N_3111,In_282,In_92);
nor U3112 (N_3112,In_321,In_682);
and U3113 (N_3113,In_537,In_854);
and U3114 (N_3114,In_888,In_45);
and U3115 (N_3115,In_138,In_685);
nor U3116 (N_3116,In_524,In_529);
nor U3117 (N_3117,In_165,In_80);
nor U3118 (N_3118,In_299,In_812);
nor U3119 (N_3119,In_388,In_874);
nor U3120 (N_3120,In_733,In_696);
and U3121 (N_3121,In_108,In_453);
nor U3122 (N_3122,In_482,In_114);
or U3123 (N_3123,In_672,In_301);
nand U3124 (N_3124,In_395,In_803);
nor U3125 (N_3125,In_655,In_660);
or U3126 (N_3126,In_296,In_191);
nand U3127 (N_3127,In_453,In_308);
nor U3128 (N_3128,In_111,In_859);
and U3129 (N_3129,In_453,In_901);
nand U3130 (N_3130,In_723,In_941);
nand U3131 (N_3131,In_566,In_616);
nand U3132 (N_3132,In_223,In_736);
nor U3133 (N_3133,In_774,In_714);
nor U3134 (N_3134,In_18,In_879);
xnor U3135 (N_3135,In_960,In_190);
nor U3136 (N_3136,In_933,In_902);
and U3137 (N_3137,In_836,In_189);
or U3138 (N_3138,In_254,In_870);
xnor U3139 (N_3139,In_462,In_996);
nand U3140 (N_3140,In_767,In_814);
nand U3141 (N_3141,In_625,In_466);
xor U3142 (N_3142,In_264,In_216);
xnor U3143 (N_3143,In_374,In_337);
nand U3144 (N_3144,In_146,In_684);
and U3145 (N_3145,In_876,In_127);
or U3146 (N_3146,In_532,In_986);
nor U3147 (N_3147,In_256,In_124);
nand U3148 (N_3148,In_327,In_912);
nor U3149 (N_3149,In_790,In_126);
and U3150 (N_3150,In_696,In_32);
and U3151 (N_3151,In_187,In_600);
nor U3152 (N_3152,In_720,In_416);
and U3153 (N_3153,In_302,In_167);
or U3154 (N_3154,In_433,In_950);
nand U3155 (N_3155,In_446,In_6);
nand U3156 (N_3156,In_706,In_877);
nor U3157 (N_3157,In_457,In_162);
or U3158 (N_3158,In_889,In_41);
or U3159 (N_3159,In_155,In_429);
and U3160 (N_3160,In_52,In_698);
nand U3161 (N_3161,In_382,In_937);
and U3162 (N_3162,In_830,In_368);
and U3163 (N_3163,In_758,In_659);
nand U3164 (N_3164,In_849,In_95);
nor U3165 (N_3165,In_245,In_807);
nor U3166 (N_3166,In_704,In_156);
nand U3167 (N_3167,In_719,In_449);
nor U3168 (N_3168,In_116,In_93);
nor U3169 (N_3169,In_157,In_836);
and U3170 (N_3170,In_6,In_62);
and U3171 (N_3171,In_801,In_427);
nor U3172 (N_3172,In_801,In_993);
or U3173 (N_3173,In_902,In_675);
nor U3174 (N_3174,In_398,In_15);
nand U3175 (N_3175,In_764,In_957);
nand U3176 (N_3176,In_452,In_173);
nor U3177 (N_3177,In_972,In_404);
or U3178 (N_3178,In_767,In_610);
or U3179 (N_3179,In_152,In_408);
nor U3180 (N_3180,In_727,In_819);
and U3181 (N_3181,In_865,In_444);
nor U3182 (N_3182,In_977,In_663);
nand U3183 (N_3183,In_960,In_298);
and U3184 (N_3184,In_453,In_668);
xor U3185 (N_3185,In_357,In_974);
and U3186 (N_3186,In_186,In_808);
or U3187 (N_3187,In_166,In_220);
and U3188 (N_3188,In_424,In_34);
and U3189 (N_3189,In_730,In_665);
xor U3190 (N_3190,In_921,In_918);
xor U3191 (N_3191,In_491,In_366);
nor U3192 (N_3192,In_644,In_385);
xnor U3193 (N_3193,In_55,In_961);
or U3194 (N_3194,In_112,In_552);
nand U3195 (N_3195,In_39,In_959);
or U3196 (N_3196,In_950,In_185);
and U3197 (N_3197,In_906,In_572);
nor U3198 (N_3198,In_930,In_854);
or U3199 (N_3199,In_252,In_636);
and U3200 (N_3200,In_303,In_544);
and U3201 (N_3201,In_623,In_848);
and U3202 (N_3202,In_72,In_756);
nor U3203 (N_3203,In_84,In_511);
xnor U3204 (N_3204,In_233,In_30);
or U3205 (N_3205,In_787,In_874);
nand U3206 (N_3206,In_744,In_192);
and U3207 (N_3207,In_497,In_883);
nand U3208 (N_3208,In_357,In_973);
nand U3209 (N_3209,In_695,In_450);
nand U3210 (N_3210,In_777,In_758);
and U3211 (N_3211,In_895,In_891);
xnor U3212 (N_3212,In_90,In_780);
or U3213 (N_3213,In_400,In_176);
or U3214 (N_3214,In_733,In_880);
and U3215 (N_3215,In_266,In_806);
nor U3216 (N_3216,In_913,In_212);
nor U3217 (N_3217,In_611,In_396);
xnor U3218 (N_3218,In_320,In_994);
and U3219 (N_3219,In_849,In_977);
xnor U3220 (N_3220,In_237,In_110);
nand U3221 (N_3221,In_928,In_856);
or U3222 (N_3222,In_38,In_482);
and U3223 (N_3223,In_890,In_436);
nand U3224 (N_3224,In_682,In_550);
nor U3225 (N_3225,In_536,In_782);
and U3226 (N_3226,In_560,In_225);
nor U3227 (N_3227,In_837,In_538);
nand U3228 (N_3228,In_909,In_668);
nand U3229 (N_3229,In_416,In_381);
and U3230 (N_3230,In_342,In_538);
nor U3231 (N_3231,In_609,In_472);
nor U3232 (N_3232,In_924,In_369);
or U3233 (N_3233,In_595,In_953);
nor U3234 (N_3234,In_980,In_907);
or U3235 (N_3235,In_826,In_448);
nor U3236 (N_3236,In_576,In_163);
or U3237 (N_3237,In_68,In_72);
xor U3238 (N_3238,In_190,In_261);
nand U3239 (N_3239,In_886,In_711);
nor U3240 (N_3240,In_389,In_782);
or U3241 (N_3241,In_960,In_622);
xnor U3242 (N_3242,In_272,In_172);
or U3243 (N_3243,In_550,In_656);
or U3244 (N_3244,In_577,In_475);
nor U3245 (N_3245,In_409,In_853);
nor U3246 (N_3246,In_757,In_533);
or U3247 (N_3247,In_315,In_429);
nor U3248 (N_3248,In_69,In_515);
nor U3249 (N_3249,In_803,In_780);
and U3250 (N_3250,In_307,In_767);
or U3251 (N_3251,In_457,In_45);
xnor U3252 (N_3252,In_165,In_353);
nand U3253 (N_3253,In_111,In_849);
nand U3254 (N_3254,In_55,In_53);
or U3255 (N_3255,In_18,In_513);
or U3256 (N_3256,In_977,In_458);
nand U3257 (N_3257,In_617,In_612);
nand U3258 (N_3258,In_354,In_996);
or U3259 (N_3259,In_295,In_790);
nand U3260 (N_3260,In_513,In_479);
and U3261 (N_3261,In_660,In_104);
xor U3262 (N_3262,In_169,In_420);
or U3263 (N_3263,In_812,In_604);
and U3264 (N_3264,In_622,In_327);
or U3265 (N_3265,In_333,In_25);
or U3266 (N_3266,In_570,In_762);
or U3267 (N_3267,In_784,In_102);
nand U3268 (N_3268,In_916,In_933);
nand U3269 (N_3269,In_114,In_479);
and U3270 (N_3270,In_313,In_522);
and U3271 (N_3271,In_673,In_210);
xnor U3272 (N_3272,In_412,In_189);
nor U3273 (N_3273,In_332,In_805);
nor U3274 (N_3274,In_25,In_742);
nand U3275 (N_3275,In_282,In_166);
or U3276 (N_3276,In_835,In_102);
nand U3277 (N_3277,In_887,In_831);
and U3278 (N_3278,In_834,In_309);
nor U3279 (N_3279,In_458,In_814);
or U3280 (N_3280,In_820,In_781);
or U3281 (N_3281,In_535,In_21);
nor U3282 (N_3282,In_119,In_47);
nand U3283 (N_3283,In_520,In_647);
nand U3284 (N_3284,In_195,In_559);
and U3285 (N_3285,In_936,In_186);
nor U3286 (N_3286,In_981,In_369);
nor U3287 (N_3287,In_239,In_38);
nor U3288 (N_3288,In_158,In_832);
and U3289 (N_3289,In_825,In_254);
and U3290 (N_3290,In_351,In_976);
or U3291 (N_3291,In_777,In_87);
nor U3292 (N_3292,In_426,In_559);
or U3293 (N_3293,In_234,In_463);
and U3294 (N_3294,In_591,In_532);
or U3295 (N_3295,In_615,In_323);
nand U3296 (N_3296,In_947,In_916);
and U3297 (N_3297,In_193,In_624);
and U3298 (N_3298,In_184,In_128);
nor U3299 (N_3299,In_472,In_373);
nor U3300 (N_3300,In_466,In_236);
or U3301 (N_3301,In_692,In_30);
nand U3302 (N_3302,In_786,In_170);
or U3303 (N_3303,In_544,In_389);
nand U3304 (N_3304,In_433,In_389);
or U3305 (N_3305,In_826,In_486);
nor U3306 (N_3306,In_362,In_548);
and U3307 (N_3307,In_837,In_894);
or U3308 (N_3308,In_360,In_898);
or U3309 (N_3309,In_507,In_344);
xor U3310 (N_3310,In_536,In_562);
and U3311 (N_3311,In_282,In_338);
nor U3312 (N_3312,In_427,In_192);
xor U3313 (N_3313,In_871,In_159);
or U3314 (N_3314,In_685,In_28);
xor U3315 (N_3315,In_466,In_14);
nand U3316 (N_3316,In_147,In_912);
nor U3317 (N_3317,In_488,In_478);
or U3318 (N_3318,In_544,In_779);
or U3319 (N_3319,In_623,In_649);
nand U3320 (N_3320,In_492,In_539);
nand U3321 (N_3321,In_583,In_140);
or U3322 (N_3322,In_706,In_302);
and U3323 (N_3323,In_213,In_164);
nand U3324 (N_3324,In_402,In_79);
nand U3325 (N_3325,In_740,In_949);
nand U3326 (N_3326,In_511,In_853);
and U3327 (N_3327,In_762,In_331);
and U3328 (N_3328,In_713,In_266);
nor U3329 (N_3329,In_517,In_938);
xnor U3330 (N_3330,In_534,In_683);
nand U3331 (N_3331,In_65,In_515);
nand U3332 (N_3332,In_182,In_3);
and U3333 (N_3333,In_82,In_364);
and U3334 (N_3334,In_788,In_30);
nor U3335 (N_3335,In_811,In_342);
or U3336 (N_3336,In_457,In_402);
or U3337 (N_3337,In_100,In_572);
or U3338 (N_3338,In_953,In_494);
nor U3339 (N_3339,In_605,In_397);
and U3340 (N_3340,In_63,In_987);
nor U3341 (N_3341,In_846,In_395);
and U3342 (N_3342,In_552,In_762);
nor U3343 (N_3343,In_928,In_696);
nand U3344 (N_3344,In_78,In_428);
nand U3345 (N_3345,In_672,In_606);
or U3346 (N_3346,In_623,In_821);
or U3347 (N_3347,In_796,In_740);
nor U3348 (N_3348,In_342,In_951);
nor U3349 (N_3349,In_630,In_737);
and U3350 (N_3350,In_623,In_982);
nor U3351 (N_3351,In_248,In_486);
and U3352 (N_3352,In_374,In_668);
and U3353 (N_3353,In_58,In_574);
nand U3354 (N_3354,In_855,In_652);
xnor U3355 (N_3355,In_514,In_291);
nand U3356 (N_3356,In_763,In_67);
nor U3357 (N_3357,In_972,In_576);
nand U3358 (N_3358,In_416,In_419);
nand U3359 (N_3359,In_1,In_452);
nor U3360 (N_3360,In_216,In_732);
or U3361 (N_3361,In_762,In_180);
nor U3362 (N_3362,In_565,In_750);
and U3363 (N_3363,In_659,In_603);
nand U3364 (N_3364,In_382,In_361);
nor U3365 (N_3365,In_560,In_649);
nand U3366 (N_3366,In_483,In_383);
nand U3367 (N_3367,In_6,In_816);
nand U3368 (N_3368,In_798,In_714);
or U3369 (N_3369,In_233,In_296);
nor U3370 (N_3370,In_524,In_359);
xnor U3371 (N_3371,In_819,In_547);
or U3372 (N_3372,In_860,In_445);
nand U3373 (N_3373,In_263,In_218);
nand U3374 (N_3374,In_681,In_789);
or U3375 (N_3375,In_529,In_353);
or U3376 (N_3376,In_547,In_426);
nand U3377 (N_3377,In_366,In_347);
nand U3378 (N_3378,In_799,In_170);
nand U3379 (N_3379,In_633,In_200);
nor U3380 (N_3380,In_633,In_46);
nand U3381 (N_3381,In_857,In_541);
and U3382 (N_3382,In_779,In_725);
and U3383 (N_3383,In_766,In_973);
nor U3384 (N_3384,In_710,In_986);
and U3385 (N_3385,In_958,In_944);
or U3386 (N_3386,In_670,In_209);
xor U3387 (N_3387,In_449,In_402);
and U3388 (N_3388,In_443,In_223);
and U3389 (N_3389,In_511,In_364);
or U3390 (N_3390,In_928,In_702);
or U3391 (N_3391,In_983,In_996);
nand U3392 (N_3392,In_74,In_566);
nor U3393 (N_3393,In_61,In_892);
nand U3394 (N_3394,In_612,In_939);
nand U3395 (N_3395,In_218,In_930);
or U3396 (N_3396,In_815,In_235);
and U3397 (N_3397,In_255,In_397);
or U3398 (N_3398,In_106,In_456);
or U3399 (N_3399,In_911,In_851);
nor U3400 (N_3400,In_881,In_674);
nor U3401 (N_3401,In_712,In_690);
and U3402 (N_3402,In_98,In_119);
or U3403 (N_3403,In_234,In_356);
xnor U3404 (N_3404,In_41,In_162);
or U3405 (N_3405,In_787,In_178);
or U3406 (N_3406,In_344,In_461);
nand U3407 (N_3407,In_286,In_429);
or U3408 (N_3408,In_696,In_542);
nor U3409 (N_3409,In_107,In_610);
and U3410 (N_3410,In_605,In_620);
and U3411 (N_3411,In_450,In_91);
xor U3412 (N_3412,In_437,In_29);
nor U3413 (N_3413,In_180,In_718);
or U3414 (N_3414,In_266,In_396);
or U3415 (N_3415,In_411,In_377);
and U3416 (N_3416,In_90,In_845);
or U3417 (N_3417,In_908,In_348);
or U3418 (N_3418,In_958,In_501);
xnor U3419 (N_3419,In_592,In_465);
or U3420 (N_3420,In_304,In_41);
and U3421 (N_3421,In_426,In_81);
nand U3422 (N_3422,In_669,In_63);
nand U3423 (N_3423,In_81,In_117);
xnor U3424 (N_3424,In_84,In_213);
and U3425 (N_3425,In_231,In_173);
nor U3426 (N_3426,In_156,In_260);
or U3427 (N_3427,In_688,In_418);
and U3428 (N_3428,In_942,In_344);
nor U3429 (N_3429,In_530,In_830);
nand U3430 (N_3430,In_810,In_315);
and U3431 (N_3431,In_150,In_134);
nand U3432 (N_3432,In_733,In_826);
nand U3433 (N_3433,In_973,In_75);
and U3434 (N_3434,In_719,In_297);
nand U3435 (N_3435,In_367,In_815);
nor U3436 (N_3436,In_101,In_881);
nand U3437 (N_3437,In_98,In_819);
nor U3438 (N_3438,In_481,In_924);
nand U3439 (N_3439,In_218,In_16);
nor U3440 (N_3440,In_930,In_398);
nand U3441 (N_3441,In_673,In_115);
nor U3442 (N_3442,In_869,In_615);
nand U3443 (N_3443,In_262,In_978);
nor U3444 (N_3444,In_725,In_160);
nand U3445 (N_3445,In_3,In_628);
nor U3446 (N_3446,In_868,In_377);
and U3447 (N_3447,In_698,In_501);
nand U3448 (N_3448,In_595,In_755);
nor U3449 (N_3449,In_755,In_174);
or U3450 (N_3450,In_541,In_677);
nor U3451 (N_3451,In_2,In_373);
nand U3452 (N_3452,In_407,In_188);
or U3453 (N_3453,In_922,In_641);
nor U3454 (N_3454,In_448,In_843);
nand U3455 (N_3455,In_915,In_781);
xor U3456 (N_3456,In_568,In_838);
nand U3457 (N_3457,In_1,In_272);
nor U3458 (N_3458,In_433,In_290);
nor U3459 (N_3459,In_659,In_698);
nor U3460 (N_3460,In_771,In_962);
or U3461 (N_3461,In_211,In_344);
nor U3462 (N_3462,In_324,In_931);
nor U3463 (N_3463,In_510,In_869);
or U3464 (N_3464,In_855,In_543);
nor U3465 (N_3465,In_27,In_505);
nor U3466 (N_3466,In_393,In_590);
and U3467 (N_3467,In_856,In_445);
xnor U3468 (N_3468,In_730,In_229);
nor U3469 (N_3469,In_130,In_435);
xnor U3470 (N_3470,In_779,In_529);
nor U3471 (N_3471,In_262,In_836);
or U3472 (N_3472,In_767,In_201);
nor U3473 (N_3473,In_992,In_787);
and U3474 (N_3474,In_386,In_604);
or U3475 (N_3475,In_224,In_972);
nand U3476 (N_3476,In_533,In_231);
nor U3477 (N_3477,In_400,In_997);
nand U3478 (N_3478,In_280,In_305);
and U3479 (N_3479,In_656,In_865);
or U3480 (N_3480,In_926,In_7);
and U3481 (N_3481,In_475,In_452);
or U3482 (N_3482,In_396,In_954);
xnor U3483 (N_3483,In_278,In_6);
nor U3484 (N_3484,In_153,In_556);
or U3485 (N_3485,In_753,In_983);
nor U3486 (N_3486,In_978,In_839);
nor U3487 (N_3487,In_881,In_596);
xnor U3488 (N_3488,In_145,In_357);
or U3489 (N_3489,In_961,In_194);
and U3490 (N_3490,In_40,In_508);
or U3491 (N_3491,In_635,In_202);
nand U3492 (N_3492,In_225,In_439);
nand U3493 (N_3493,In_907,In_888);
and U3494 (N_3494,In_703,In_285);
nand U3495 (N_3495,In_121,In_919);
xnor U3496 (N_3496,In_917,In_873);
nor U3497 (N_3497,In_816,In_221);
and U3498 (N_3498,In_668,In_107);
or U3499 (N_3499,In_241,In_76);
nand U3500 (N_3500,In_277,In_129);
nand U3501 (N_3501,In_714,In_787);
and U3502 (N_3502,In_77,In_304);
or U3503 (N_3503,In_45,In_952);
nand U3504 (N_3504,In_140,In_125);
or U3505 (N_3505,In_398,In_849);
or U3506 (N_3506,In_33,In_54);
nor U3507 (N_3507,In_905,In_509);
or U3508 (N_3508,In_936,In_703);
nor U3509 (N_3509,In_955,In_75);
or U3510 (N_3510,In_310,In_770);
and U3511 (N_3511,In_340,In_509);
nor U3512 (N_3512,In_474,In_601);
xor U3513 (N_3513,In_700,In_638);
nand U3514 (N_3514,In_944,In_72);
xor U3515 (N_3515,In_81,In_897);
and U3516 (N_3516,In_978,In_257);
or U3517 (N_3517,In_520,In_114);
and U3518 (N_3518,In_6,In_630);
and U3519 (N_3519,In_491,In_486);
or U3520 (N_3520,In_516,In_826);
nand U3521 (N_3521,In_80,In_853);
nor U3522 (N_3522,In_628,In_732);
xor U3523 (N_3523,In_491,In_867);
nor U3524 (N_3524,In_762,In_295);
or U3525 (N_3525,In_900,In_577);
nor U3526 (N_3526,In_455,In_415);
nand U3527 (N_3527,In_902,In_840);
nor U3528 (N_3528,In_769,In_916);
and U3529 (N_3529,In_615,In_897);
nand U3530 (N_3530,In_223,In_56);
xor U3531 (N_3531,In_624,In_355);
or U3532 (N_3532,In_703,In_229);
and U3533 (N_3533,In_601,In_784);
nor U3534 (N_3534,In_245,In_738);
nand U3535 (N_3535,In_801,In_642);
xnor U3536 (N_3536,In_411,In_541);
or U3537 (N_3537,In_762,In_406);
nand U3538 (N_3538,In_86,In_41);
and U3539 (N_3539,In_929,In_31);
nor U3540 (N_3540,In_806,In_648);
nand U3541 (N_3541,In_222,In_96);
or U3542 (N_3542,In_541,In_772);
nand U3543 (N_3543,In_426,In_336);
nor U3544 (N_3544,In_721,In_786);
nand U3545 (N_3545,In_314,In_90);
or U3546 (N_3546,In_922,In_129);
or U3547 (N_3547,In_655,In_808);
or U3548 (N_3548,In_793,In_504);
nand U3549 (N_3549,In_93,In_3);
and U3550 (N_3550,In_370,In_6);
xnor U3551 (N_3551,In_304,In_685);
and U3552 (N_3552,In_136,In_675);
or U3553 (N_3553,In_956,In_695);
nand U3554 (N_3554,In_155,In_61);
nor U3555 (N_3555,In_529,In_719);
nand U3556 (N_3556,In_666,In_640);
nand U3557 (N_3557,In_488,In_917);
or U3558 (N_3558,In_356,In_35);
nand U3559 (N_3559,In_620,In_410);
nor U3560 (N_3560,In_452,In_100);
xor U3561 (N_3561,In_285,In_394);
and U3562 (N_3562,In_617,In_887);
and U3563 (N_3563,In_147,In_854);
nand U3564 (N_3564,In_864,In_550);
and U3565 (N_3565,In_493,In_233);
or U3566 (N_3566,In_976,In_995);
nor U3567 (N_3567,In_738,In_143);
or U3568 (N_3568,In_39,In_342);
nor U3569 (N_3569,In_325,In_645);
nor U3570 (N_3570,In_494,In_38);
nand U3571 (N_3571,In_421,In_905);
or U3572 (N_3572,In_402,In_451);
nand U3573 (N_3573,In_945,In_917);
and U3574 (N_3574,In_977,In_707);
xnor U3575 (N_3575,In_272,In_455);
and U3576 (N_3576,In_382,In_722);
nor U3577 (N_3577,In_926,In_876);
nand U3578 (N_3578,In_107,In_503);
nor U3579 (N_3579,In_91,In_393);
and U3580 (N_3580,In_610,In_742);
or U3581 (N_3581,In_640,In_15);
and U3582 (N_3582,In_59,In_69);
or U3583 (N_3583,In_36,In_600);
or U3584 (N_3584,In_868,In_42);
or U3585 (N_3585,In_476,In_733);
or U3586 (N_3586,In_903,In_612);
nor U3587 (N_3587,In_912,In_981);
and U3588 (N_3588,In_416,In_270);
or U3589 (N_3589,In_997,In_429);
nand U3590 (N_3590,In_60,In_745);
nand U3591 (N_3591,In_923,In_89);
and U3592 (N_3592,In_728,In_853);
and U3593 (N_3593,In_598,In_630);
nor U3594 (N_3594,In_990,In_140);
or U3595 (N_3595,In_561,In_669);
nand U3596 (N_3596,In_609,In_425);
xnor U3597 (N_3597,In_862,In_723);
or U3598 (N_3598,In_241,In_596);
or U3599 (N_3599,In_340,In_609);
and U3600 (N_3600,In_445,In_52);
nand U3601 (N_3601,In_824,In_93);
nor U3602 (N_3602,In_213,In_167);
or U3603 (N_3603,In_987,In_93);
or U3604 (N_3604,In_246,In_828);
nand U3605 (N_3605,In_761,In_816);
and U3606 (N_3606,In_868,In_989);
nand U3607 (N_3607,In_506,In_806);
nand U3608 (N_3608,In_477,In_189);
nor U3609 (N_3609,In_339,In_568);
nand U3610 (N_3610,In_843,In_812);
nand U3611 (N_3611,In_120,In_461);
and U3612 (N_3612,In_454,In_290);
nand U3613 (N_3613,In_827,In_650);
nand U3614 (N_3614,In_365,In_341);
nand U3615 (N_3615,In_935,In_641);
nor U3616 (N_3616,In_677,In_777);
or U3617 (N_3617,In_408,In_714);
nor U3618 (N_3618,In_745,In_931);
nor U3619 (N_3619,In_496,In_158);
nor U3620 (N_3620,In_310,In_89);
nand U3621 (N_3621,In_896,In_983);
nand U3622 (N_3622,In_972,In_445);
nor U3623 (N_3623,In_716,In_26);
nor U3624 (N_3624,In_923,In_364);
nand U3625 (N_3625,In_854,In_321);
or U3626 (N_3626,In_188,In_680);
or U3627 (N_3627,In_783,In_22);
and U3628 (N_3628,In_990,In_152);
nand U3629 (N_3629,In_539,In_667);
nor U3630 (N_3630,In_967,In_263);
nor U3631 (N_3631,In_417,In_258);
xnor U3632 (N_3632,In_171,In_21);
and U3633 (N_3633,In_144,In_977);
and U3634 (N_3634,In_564,In_488);
nand U3635 (N_3635,In_752,In_201);
nand U3636 (N_3636,In_497,In_744);
and U3637 (N_3637,In_586,In_226);
and U3638 (N_3638,In_172,In_312);
nand U3639 (N_3639,In_393,In_866);
nand U3640 (N_3640,In_626,In_45);
nand U3641 (N_3641,In_58,In_911);
or U3642 (N_3642,In_748,In_15);
nor U3643 (N_3643,In_491,In_18);
nor U3644 (N_3644,In_366,In_946);
or U3645 (N_3645,In_964,In_836);
and U3646 (N_3646,In_681,In_61);
nor U3647 (N_3647,In_270,In_615);
nor U3648 (N_3648,In_4,In_934);
and U3649 (N_3649,In_412,In_234);
nor U3650 (N_3650,In_802,In_999);
or U3651 (N_3651,In_569,In_419);
xor U3652 (N_3652,In_300,In_387);
and U3653 (N_3653,In_477,In_254);
nor U3654 (N_3654,In_276,In_777);
or U3655 (N_3655,In_441,In_583);
nand U3656 (N_3656,In_81,In_617);
nor U3657 (N_3657,In_310,In_360);
and U3658 (N_3658,In_498,In_454);
or U3659 (N_3659,In_863,In_641);
nand U3660 (N_3660,In_301,In_29);
xor U3661 (N_3661,In_392,In_799);
and U3662 (N_3662,In_508,In_470);
and U3663 (N_3663,In_231,In_209);
nand U3664 (N_3664,In_203,In_798);
xor U3665 (N_3665,In_560,In_599);
or U3666 (N_3666,In_553,In_995);
or U3667 (N_3667,In_892,In_413);
nor U3668 (N_3668,In_580,In_254);
nor U3669 (N_3669,In_145,In_71);
nor U3670 (N_3670,In_347,In_452);
and U3671 (N_3671,In_618,In_483);
and U3672 (N_3672,In_921,In_354);
and U3673 (N_3673,In_993,In_52);
nor U3674 (N_3674,In_520,In_550);
nor U3675 (N_3675,In_229,In_131);
or U3676 (N_3676,In_395,In_875);
nand U3677 (N_3677,In_867,In_140);
xnor U3678 (N_3678,In_788,In_903);
and U3679 (N_3679,In_288,In_475);
or U3680 (N_3680,In_722,In_710);
nor U3681 (N_3681,In_218,In_791);
nand U3682 (N_3682,In_175,In_261);
xor U3683 (N_3683,In_263,In_105);
and U3684 (N_3684,In_394,In_237);
or U3685 (N_3685,In_526,In_568);
or U3686 (N_3686,In_690,In_922);
and U3687 (N_3687,In_637,In_941);
nor U3688 (N_3688,In_444,In_442);
nand U3689 (N_3689,In_470,In_888);
xor U3690 (N_3690,In_241,In_842);
nand U3691 (N_3691,In_724,In_430);
and U3692 (N_3692,In_472,In_926);
and U3693 (N_3693,In_7,In_958);
xor U3694 (N_3694,In_910,In_973);
nor U3695 (N_3695,In_153,In_297);
nand U3696 (N_3696,In_759,In_999);
and U3697 (N_3697,In_918,In_79);
nor U3698 (N_3698,In_891,In_767);
nand U3699 (N_3699,In_372,In_775);
or U3700 (N_3700,In_41,In_37);
nand U3701 (N_3701,In_777,In_653);
and U3702 (N_3702,In_212,In_51);
or U3703 (N_3703,In_818,In_519);
nor U3704 (N_3704,In_593,In_614);
and U3705 (N_3705,In_155,In_653);
nand U3706 (N_3706,In_675,In_619);
and U3707 (N_3707,In_747,In_175);
or U3708 (N_3708,In_990,In_126);
xor U3709 (N_3709,In_560,In_258);
nand U3710 (N_3710,In_822,In_256);
nand U3711 (N_3711,In_312,In_303);
nand U3712 (N_3712,In_503,In_47);
nand U3713 (N_3713,In_143,In_102);
xnor U3714 (N_3714,In_399,In_753);
nand U3715 (N_3715,In_593,In_599);
or U3716 (N_3716,In_542,In_52);
xor U3717 (N_3717,In_129,In_209);
and U3718 (N_3718,In_349,In_533);
and U3719 (N_3719,In_611,In_876);
nand U3720 (N_3720,In_522,In_638);
nor U3721 (N_3721,In_86,In_963);
and U3722 (N_3722,In_841,In_752);
and U3723 (N_3723,In_328,In_978);
xor U3724 (N_3724,In_632,In_454);
and U3725 (N_3725,In_513,In_385);
and U3726 (N_3726,In_454,In_48);
nor U3727 (N_3727,In_962,In_783);
nand U3728 (N_3728,In_286,In_594);
xnor U3729 (N_3729,In_865,In_679);
nor U3730 (N_3730,In_570,In_219);
nor U3731 (N_3731,In_664,In_116);
and U3732 (N_3732,In_132,In_315);
xnor U3733 (N_3733,In_984,In_101);
or U3734 (N_3734,In_949,In_192);
nand U3735 (N_3735,In_126,In_921);
or U3736 (N_3736,In_929,In_512);
and U3737 (N_3737,In_623,In_551);
or U3738 (N_3738,In_632,In_262);
and U3739 (N_3739,In_149,In_183);
and U3740 (N_3740,In_274,In_811);
nor U3741 (N_3741,In_734,In_437);
nor U3742 (N_3742,In_815,In_545);
nand U3743 (N_3743,In_903,In_268);
or U3744 (N_3744,In_139,In_796);
nor U3745 (N_3745,In_412,In_44);
nor U3746 (N_3746,In_380,In_259);
nor U3747 (N_3747,In_602,In_942);
nor U3748 (N_3748,In_512,In_973);
or U3749 (N_3749,In_955,In_411);
or U3750 (N_3750,In_196,In_843);
or U3751 (N_3751,In_82,In_78);
and U3752 (N_3752,In_307,In_694);
nor U3753 (N_3753,In_921,In_906);
xnor U3754 (N_3754,In_704,In_512);
and U3755 (N_3755,In_449,In_95);
and U3756 (N_3756,In_822,In_922);
and U3757 (N_3757,In_806,In_249);
nor U3758 (N_3758,In_110,In_431);
nand U3759 (N_3759,In_522,In_384);
xor U3760 (N_3760,In_590,In_909);
nor U3761 (N_3761,In_258,In_93);
or U3762 (N_3762,In_632,In_275);
or U3763 (N_3763,In_41,In_563);
nor U3764 (N_3764,In_392,In_29);
nor U3765 (N_3765,In_409,In_476);
or U3766 (N_3766,In_311,In_527);
nand U3767 (N_3767,In_904,In_4);
and U3768 (N_3768,In_395,In_965);
or U3769 (N_3769,In_499,In_854);
or U3770 (N_3770,In_576,In_74);
and U3771 (N_3771,In_185,In_970);
or U3772 (N_3772,In_268,In_797);
nor U3773 (N_3773,In_84,In_220);
nor U3774 (N_3774,In_259,In_437);
or U3775 (N_3775,In_980,In_182);
xor U3776 (N_3776,In_869,In_317);
and U3777 (N_3777,In_234,In_200);
or U3778 (N_3778,In_399,In_344);
or U3779 (N_3779,In_226,In_105);
nor U3780 (N_3780,In_79,In_595);
and U3781 (N_3781,In_912,In_45);
xnor U3782 (N_3782,In_227,In_442);
xnor U3783 (N_3783,In_852,In_496);
or U3784 (N_3784,In_729,In_48);
nor U3785 (N_3785,In_81,In_563);
nor U3786 (N_3786,In_521,In_387);
and U3787 (N_3787,In_214,In_553);
nor U3788 (N_3788,In_767,In_720);
and U3789 (N_3789,In_32,In_432);
nand U3790 (N_3790,In_11,In_256);
or U3791 (N_3791,In_465,In_620);
or U3792 (N_3792,In_525,In_734);
nand U3793 (N_3793,In_132,In_446);
or U3794 (N_3794,In_6,In_34);
nand U3795 (N_3795,In_76,In_973);
nand U3796 (N_3796,In_459,In_260);
nand U3797 (N_3797,In_608,In_788);
nor U3798 (N_3798,In_379,In_407);
nand U3799 (N_3799,In_896,In_594);
nand U3800 (N_3800,In_695,In_596);
nor U3801 (N_3801,In_683,In_7);
or U3802 (N_3802,In_353,In_702);
or U3803 (N_3803,In_227,In_457);
xnor U3804 (N_3804,In_723,In_180);
nand U3805 (N_3805,In_842,In_859);
or U3806 (N_3806,In_415,In_554);
nor U3807 (N_3807,In_622,In_310);
nand U3808 (N_3808,In_982,In_793);
nand U3809 (N_3809,In_573,In_482);
nor U3810 (N_3810,In_215,In_5);
nor U3811 (N_3811,In_865,In_328);
nor U3812 (N_3812,In_859,In_897);
nor U3813 (N_3813,In_228,In_863);
nor U3814 (N_3814,In_507,In_508);
nor U3815 (N_3815,In_181,In_323);
nor U3816 (N_3816,In_70,In_646);
and U3817 (N_3817,In_184,In_167);
nand U3818 (N_3818,In_704,In_492);
and U3819 (N_3819,In_768,In_625);
or U3820 (N_3820,In_546,In_862);
nor U3821 (N_3821,In_353,In_798);
nand U3822 (N_3822,In_783,In_179);
nor U3823 (N_3823,In_330,In_544);
nand U3824 (N_3824,In_35,In_954);
nand U3825 (N_3825,In_643,In_246);
nand U3826 (N_3826,In_942,In_437);
nor U3827 (N_3827,In_735,In_361);
or U3828 (N_3828,In_447,In_580);
and U3829 (N_3829,In_105,In_640);
xor U3830 (N_3830,In_508,In_361);
nand U3831 (N_3831,In_445,In_916);
xnor U3832 (N_3832,In_696,In_305);
or U3833 (N_3833,In_675,In_180);
and U3834 (N_3834,In_828,In_466);
nor U3835 (N_3835,In_120,In_262);
nor U3836 (N_3836,In_657,In_648);
or U3837 (N_3837,In_352,In_666);
or U3838 (N_3838,In_188,In_512);
and U3839 (N_3839,In_769,In_162);
or U3840 (N_3840,In_477,In_263);
nand U3841 (N_3841,In_109,In_285);
nand U3842 (N_3842,In_660,In_731);
nand U3843 (N_3843,In_821,In_484);
nor U3844 (N_3844,In_272,In_979);
nand U3845 (N_3845,In_292,In_764);
or U3846 (N_3846,In_991,In_222);
nor U3847 (N_3847,In_1,In_312);
and U3848 (N_3848,In_625,In_365);
nand U3849 (N_3849,In_784,In_54);
or U3850 (N_3850,In_423,In_422);
or U3851 (N_3851,In_958,In_579);
or U3852 (N_3852,In_290,In_746);
nor U3853 (N_3853,In_505,In_880);
or U3854 (N_3854,In_928,In_935);
and U3855 (N_3855,In_600,In_259);
xnor U3856 (N_3856,In_840,In_240);
nor U3857 (N_3857,In_677,In_998);
nand U3858 (N_3858,In_557,In_300);
and U3859 (N_3859,In_749,In_623);
nor U3860 (N_3860,In_128,In_597);
nor U3861 (N_3861,In_770,In_859);
and U3862 (N_3862,In_858,In_378);
nand U3863 (N_3863,In_446,In_31);
nor U3864 (N_3864,In_464,In_188);
or U3865 (N_3865,In_841,In_289);
nand U3866 (N_3866,In_510,In_747);
xnor U3867 (N_3867,In_764,In_19);
and U3868 (N_3868,In_666,In_249);
xnor U3869 (N_3869,In_176,In_411);
or U3870 (N_3870,In_304,In_563);
nor U3871 (N_3871,In_922,In_947);
or U3872 (N_3872,In_659,In_9);
and U3873 (N_3873,In_600,In_299);
or U3874 (N_3874,In_891,In_555);
or U3875 (N_3875,In_87,In_114);
nor U3876 (N_3876,In_302,In_113);
and U3877 (N_3877,In_795,In_710);
and U3878 (N_3878,In_608,In_942);
and U3879 (N_3879,In_873,In_958);
nor U3880 (N_3880,In_247,In_39);
nand U3881 (N_3881,In_34,In_755);
nand U3882 (N_3882,In_228,In_573);
and U3883 (N_3883,In_798,In_311);
nand U3884 (N_3884,In_346,In_802);
and U3885 (N_3885,In_838,In_43);
nor U3886 (N_3886,In_530,In_5);
nor U3887 (N_3887,In_422,In_383);
or U3888 (N_3888,In_411,In_909);
nor U3889 (N_3889,In_626,In_965);
nand U3890 (N_3890,In_380,In_547);
and U3891 (N_3891,In_103,In_333);
nand U3892 (N_3892,In_957,In_788);
nor U3893 (N_3893,In_190,In_535);
nand U3894 (N_3894,In_614,In_318);
and U3895 (N_3895,In_476,In_935);
and U3896 (N_3896,In_546,In_296);
xor U3897 (N_3897,In_479,In_473);
and U3898 (N_3898,In_831,In_133);
and U3899 (N_3899,In_182,In_320);
nor U3900 (N_3900,In_280,In_298);
nor U3901 (N_3901,In_101,In_368);
and U3902 (N_3902,In_870,In_978);
nor U3903 (N_3903,In_523,In_499);
xor U3904 (N_3904,In_531,In_984);
xnor U3905 (N_3905,In_456,In_119);
or U3906 (N_3906,In_155,In_314);
nand U3907 (N_3907,In_973,In_260);
nand U3908 (N_3908,In_677,In_808);
nor U3909 (N_3909,In_694,In_326);
nand U3910 (N_3910,In_354,In_316);
or U3911 (N_3911,In_169,In_537);
nand U3912 (N_3912,In_696,In_702);
nand U3913 (N_3913,In_300,In_714);
nand U3914 (N_3914,In_204,In_808);
and U3915 (N_3915,In_126,In_707);
or U3916 (N_3916,In_371,In_207);
nor U3917 (N_3917,In_738,In_981);
xnor U3918 (N_3918,In_163,In_855);
nor U3919 (N_3919,In_486,In_513);
nor U3920 (N_3920,In_676,In_74);
nor U3921 (N_3921,In_409,In_440);
nand U3922 (N_3922,In_493,In_21);
or U3923 (N_3923,In_316,In_438);
nor U3924 (N_3924,In_783,In_57);
and U3925 (N_3925,In_821,In_182);
and U3926 (N_3926,In_44,In_180);
or U3927 (N_3927,In_729,In_136);
nand U3928 (N_3928,In_634,In_998);
or U3929 (N_3929,In_811,In_338);
or U3930 (N_3930,In_673,In_311);
nand U3931 (N_3931,In_328,In_910);
or U3932 (N_3932,In_411,In_878);
or U3933 (N_3933,In_423,In_411);
nand U3934 (N_3934,In_140,In_551);
xor U3935 (N_3935,In_645,In_351);
nor U3936 (N_3936,In_710,In_260);
nand U3937 (N_3937,In_762,In_291);
and U3938 (N_3938,In_820,In_599);
or U3939 (N_3939,In_588,In_894);
nor U3940 (N_3940,In_375,In_762);
or U3941 (N_3941,In_959,In_461);
nor U3942 (N_3942,In_139,In_886);
nor U3943 (N_3943,In_679,In_651);
nand U3944 (N_3944,In_288,In_287);
xor U3945 (N_3945,In_322,In_426);
or U3946 (N_3946,In_917,In_61);
and U3947 (N_3947,In_700,In_99);
and U3948 (N_3948,In_713,In_432);
nor U3949 (N_3949,In_542,In_643);
nand U3950 (N_3950,In_910,In_813);
and U3951 (N_3951,In_773,In_298);
nor U3952 (N_3952,In_23,In_10);
and U3953 (N_3953,In_650,In_216);
or U3954 (N_3954,In_200,In_777);
or U3955 (N_3955,In_240,In_607);
nand U3956 (N_3956,In_230,In_275);
or U3957 (N_3957,In_967,In_814);
or U3958 (N_3958,In_924,In_0);
nor U3959 (N_3959,In_690,In_289);
and U3960 (N_3960,In_223,In_31);
and U3961 (N_3961,In_777,In_635);
or U3962 (N_3962,In_215,In_909);
and U3963 (N_3963,In_55,In_100);
xnor U3964 (N_3964,In_457,In_261);
or U3965 (N_3965,In_566,In_929);
or U3966 (N_3966,In_802,In_458);
and U3967 (N_3967,In_708,In_140);
nor U3968 (N_3968,In_680,In_162);
nand U3969 (N_3969,In_418,In_417);
xor U3970 (N_3970,In_804,In_148);
nand U3971 (N_3971,In_435,In_21);
and U3972 (N_3972,In_565,In_809);
nor U3973 (N_3973,In_760,In_256);
xor U3974 (N_3974,In_199,In_996);
xnor U3975 (N_3975,In_603,In_654);
nor U3976 (N_3976,In_545,In_647);
xor U3977 (N_3977,In_849,In_10);
nand U3978 (N_3978,In_15,In_183);
nor U3979 (N_3979,In_143,In_223);
or U3980 (N_3980,In_43,In_116);
xor U3981 (N_3981,In_243,In_314);
and U3982 (N_3982,In_837,In_394);
and U3983 (N_3983,In_142,In_636);
and U3984 (N_3984,In_212,In_389);
or U3985 (N_3985,In_342,In_770);
or U3986 (N_3986,In_522,In_899);
and U3987 (N_3987,In_804,In_711);
xnor U3988 (N_3988,In_456,In_722);
nor U3989 (N_3989,In_425,In_66);
nor U3990 (N_3990,In_327,In_504);
nor U3991 (N_3991,In_409,In_493);
nand U3992 (N_3992,In_21,In_268);
nor U3993 (N_3993,In_895,In_488);
or U3994 (N_3994,In_920,In_443);
nor U3995 (N_3995,In_487,In_728);
nand U3996 (N_3996,In_229,In_886);
or U3997 (N_3997,In_749,In_114);
or U3998 (N_3998,In_345,In_777);
nand U3999 (N_3999,In_544,In_759);
and U4000 (N_4000,In_397,In_985);
nand U4001 (N_4001,In_226,In_124);
nand U4002 (N_4002,In_58,In_643);
xor U4003 (N_4003,In_975,In_423);
or U4004 (N_4004,In_746,In_45);
or U4005 (N_4005,In_366,In_187);
nor U4006 (N_4006,In_560,In_808);
xnor U4007 (N_4007,In_617,In_297);
nor U4008 (N_4008,In_513,In_451);
or U4009 (N_4009,In_286,In_995);
nor U4010 (N_4010,In_949,In_188);
and U4011 (N_4011,In_660,In_3);
nand U4012 (N_4012,In_873,In_125);
or U4013 (N_4013,In_758,In_594);
nor U4014 (N_4014,In_945,In_323);
and U4015 (N_4015,In_458,In_571);
or U4016 (N_4016,In_427,In_809);
xnor U4017 (N_4017,In_235,In_155);
or U4018 (N_4018,In_784,In_496);
xor U4019 (N_4019,In_350,In_910);
or U4020 (N_4020,In_409,In_719);
and U4021 (N_4021,In_909,In_318);
xnor U4022 (N_4022,In_539,In_883);
nand U4023 (N_4023,In_394,In_754);
nor U4024 (N_4024,In_277,In_921);
or U4025 (N_4025,In_278,In_235);
and U4026 (N_4026,In_443,In_635);
and U4027 (N_4027,In_276,In_656);
or U4028 (N_4028,In_995,In_115);
and U4029 (N_4029,In_950,In_253);
or U4030 (N_4030,In_13,In_659);
nor U4031 (N_4031,In_224,In_76);
and U4032 (N_4032,In_670,In_105);
and U4033 (N_4033,In_488,In_735);
and U4034 (N_4034,In_574,In_339);
nand U4035 (N_4035,In_559,In_565);
nand U4036 (N_4036,In_114,In_573);
nand U4037 (N_4037,In_970,In_455);
nand U4038 (N_4038,In_206,In_106);
and U4039 (N_4039,In_122,In_95);
nand U4040 (N_4040,In_299,In_809);
nor U4041 (N_4041,In_768,In_617);
nand U4042 (N_4042,In_307,In_732);
nand U4043 (N_4043,In_990,In_857);
and U4044 (N_4044,In_182,In_114);
nand U4045 (N_4045,In_534,In_992);
nand U4046 (N_4046,In_983,In_716);
or U4047 (N_4047,In_164,In_74);
xnor U4048 (N_4048,In_576,In_811);
nand U4049 (N_4049,In_416,In_875);
nor U4050 (N_4050,In_0,In_897);
nand U4051 (N_4051,In_662,In_29);
nor U4052 (N_4052,In_902,In_704);
or U4053 (N_4053,In_389,In_358);
and U4054 (N_4054,In_616,In_492);
nand U4055 (N_4055,In_46,In_638);
and U4056 (N_4056,In_900,In_895);
xor U4057 (N_4057,In_776,In_665);
xnor U4058 (N_4058,In_567,In_550);
or U4059 (N_4059,In_683,In_236);
nand U4060 (N_4060,In_427,In_562);
xnor U4061 (N_4061,In_737,In_903);
and U4062 (N_4062,In_524,In_755);
nand U4063 (N_4063,In_628,In_871);
nor U4064 (N_4064,In_439,In_708);
or U4065 (N_4065,In_658,In_776);
or U4066 (N_4066,In_823,In_225);
nor U4067 (N_4067,In_57,In_167);
or U4068 (N_4068,In_970,In_154);
and U4069 (N_4069,In_655,In_777);
or U4070 (N_4070,In_814,In_897);
nor U4071 (N_4071,In_526,In_616);
and U4072 (N_4072,In_465,In_548);
nand U4073 (N_4073,In_144,In_888);
nand U4074 (N_4074,In_453,In_79);
and U4075 (N_4075,In_385,In_578);
and U4076 (N_4076,In_78,In_182);
nor U4077 (N_4077,In_620,In_56);
xnor U4078 (N_4078,In_184,In_615);
nor U4079 (N_4079,In_343,In_904);
nor U4080 (N_4080,In_794,In_773);
and U4081 (N_4081,In_44,In_240);
nand U4082 (N_4082,In_359,In_205);
xor U4083 (N_4083,In_722,In_491);
nand U4084 (N_4084,In_103,In_364);
and U4085 (N_4085,In_25,In_323);
nor U4086 (N_4086,In_484,In_753);
nor U4087 (N_4087,In_749,In_152);
nor U4088 (N_4088,In_436,In_546);
or U4089 (N_4089,In_597,In_885);
and U4090 (N_4090,In_85,In_225);
nand U4091 (N_4091,In_246,In_569);
and U4092 (N_4092,In_289,In_268);
or U4093 (N_4093,In_9,In_342);
and U4094 (N_4094,In_993,In_503);
and U4095 (N_4095,In_535,In_975);
xor U4096 (N_4096,In_694,In_77);
and U4097 (N_4097,In_872,In_501);
xnor U4098 (N_4098,In_511,In_917);
and U4099 (N_4099,In_851,In_526);
or U4100 (N_4100,In_388,In_255);
and U4101 (N_4101,In_562,In_432);
or U4102 (N_4102,In_48,In_493);
nand U4103 (N_4103,In_56,In_780);
and U4104 (N_4104,In_199,In_291);
or U4105 (N_4105,In_635,In_71);
xor U4106 (N_4106,In_856,In_353);
nor U4107 (N_4107,In_452,In_160);
nor U4108 (N_4108,In_808,In_245);
or U4109 (N_4109,In_71,In_810);
nand U4110 (N_4110,In_725,In_984);
nor U4111 (N_4111,In_81,In_423);
nand U4112 (N_4112,In_71,In_130);
and U4113 (N_4113,In_154,In_757);
or U4114 (N_4114,In_819,In_994);
and U4115 (N_4115,In_377,In_244);
nand U4116 (N_4116,In_331,In_483);
nand U4117 (N_4117,In_845,In_301);
nor U4118 (N_4118,In_700,In_141);
nor U4119 (N_4119,In_824,In_484);
nand U4120 (N_4120,In_327,In_261);
and U4121 (N_4121,In_227,In_889);
and U4122 (N_4122,In_183,In_24);
and U4123 (N_4123,In_52,In_972);
nor U4124 (N_4124,In_770,In_687);
nor U4125 (N_4125,In_689,In_104);
and U4126 (N_4126,In_945,In_730);
or U4127 (N_4127,In_87,In_305);
or U4128 (N_4128,In_887,In_862);
nand U4129 (N_4129,In_663,In_385);
nor U4130 (N_4130,In_580,In_402);
nor U4131 (N_4131,In_266,In_446);
nand U4132 (N_4132,In_759,In_200);
nand U4133 (N_4133,In_265,In_896);
nor U4134 (N_4134,In_579,In_36);
nor U4135 (N_4135,In_781,In_567);
nand U4136 (N_4136,In_185,In_234);
and U4137 (N_4137,In_674,In_140);
nand U4138 (N_4138,In_150,In_532);
nand U4139 (N_4139,In_466,In_368);
or U4140 (N_4140,In_804,In_695);
nand U4141 (N_4141,In_944,In_809);
xnor U4142 (N_4142,In_513,In_572);
nor U4143 (N_4143,In_36,In_919);
nor U4144 (N_4144,In_842,In_825);
xnor U4145 (N_4145,In_925,In_671);
nor U4146 (N_4146,In_143,In_86);
nand U4147 (N_4147,In_3,In_803);
or U4148 (N_4148,In_780,In_763);
and U4149 (N_4149,In_658,In_830);
nor U4150 (N_4150,In_4,In_939);
nor U4151 (N_4151,In_776,In_288);
and U4152 (N_4152,In_24,In_387);
nor U4153 (N_4153,In_307,In_439);
nor U4154 (N_4154,In_459,In_502);
and U4155 (N_4155,In_966,In_356);
nand U4156 (N_4156,In_153,In_836);
or U4157 (N_4157,In_908,In_440);
nand U4158 (N_4158,In_544,In_177);
nand U4159 (N_4159,In_202,In_329);
nand U4160 (N_4160,In_892,In_944);
nand U4161 (N_4161,In_433,In_421);
and U4162 (N_4162,In_668,In_180);
nand U4163 (N_4163,In_26,In_141);
nand U4164 (N_4164,In_802,In_72);
nor U4165 (N_4165,In_913,In_433);
nor U4166 (N_4166,In_375,In_478);
and U4167 (N_4167,In_279,In_231);
and U4168 (N_4168,In_757,In_555);
xnor U4169 (N_4169,In_741,In_605);
nor U4170 (N_4170,In_146,In_609);
xor U4171 (N_4171,In_363,In_198);
nand U4172 (N_4172,In_979,In_176);
and U4173 (N_4173,In_868,In_307);
nand U4174 (N_4174,In_464,In_155);
or U4175 (N_4175,In_516,In_841);
nor U4176 (N_4176,In_313,In_541);
and U4177 (N_4177,In_153,In_602);
nor U4178 (N_4178,In_524,In_863);
xnor U4179 (N_4179,In_293,In_447);
nor U4180 (N_4180,In_722,In_817);
or U4181 (N_4181,In_464,In_856);
xor U4182 (N_4182,In_105,In_78);
or U4183 (N_4183,In_492,In_546);
nand U4184 (N_4184,In_332,In_162);
xnor U4185 (N_4185,In_578,In_346);
nand U4186 (N_4186,In_47,In_397);
nand U4187 (N_4187,In_644,In_19);
xor U4188 (N_4188,In_239,In_601);
nand U4189 (N_4189,In_594,In_800);
nand U4190 (N_4190,In_672,In_412);
nor U4191 (N_4191,In_189,In_672);
nand U4192 (N_4192,In_596,In_774);
or U4193 (N_4193,In_266,In_604);
xnor U4194 (N_4194,In_485,In_506);
or U4195 (N_4195,In_570,In_478);
and U4196 (N_4196,In_379,In_726);
xnor U4197 (N_4197,In_132,In_776);
and U4198 (N_4198,In_204,In_880);
nor U4199 (N_4199,In_849,In_324);
and U4200 (N_4200,In_126,In_860);
xor U4201 (N_4201,In_803,In_423);
and U4202 (N_4202,In_251,In_509);
nor U4203 (N_4203,In_244,In_262);
and U4204 (N_4204,In_94,In_81);
nand U4205 (N_4205,In_820,In_245);
nor U4206 (N_4206,In_631,In_268);
or U4207 (N_4207,In_154,In_998);
nand U4208 (N_4208,In_905,In_642);
nor U4209 (N_4209,In_297,In_858);
nand U4210 (N_4210,In_359,In_683);
nor U4211 (N_4211,In_445,In_309);
xor U4212 (N_4212,In_119,In_203);
nand U4213 (N_4213,In_912,In_265);
or U4214 (N_4214,In_345,In_419);
nor U4215 (N_4215,In_322,In_755);
or U4216 (N_4216,In_182,In_629);
or U4217 (N_4217,In_481,In_878);
nand U4218 (N_4218,In_15,In_795);
nand U4219 (N_4219,In_851,In_929);
nor U4220 (N_4220,In_301,In_461);
nor U4221 (N_4221,In_685,In_228);
xnor U4222 (N_4222,In_29,In_398);
nor U4223 (N_4223,In_266,In_776);
nand U4224 (N_4224,In_871,In_718);
xor U4225 (N_4225,In_448,In_690);
or U4226 (N_4226,In_620,In_781);
nor U4227 (N_4227,In_106,In_960);
and U4228 (N_4228,In_125,In_761);
xor U4229 (N_4229,In_739,In_648);
and U4230 (N_4230,In_927,In_696);
and U4231 (N_4231,In_940,In_582);
or U4232 (N_4232,In_496,In_656);
or U4233 (N_4233,In_543,In_105);
nor U4234 (N_4234,In_668,In_389);
nor U4235 (N_4235,In_114,In_139);
nand U4236 (N_4236,In_314,In_120);
xor U4237 (N_4237,In_953,In_459);
nand U4238 (N_4238,In_314,In_106);
nand U4239 (N_4239,In_221,In_677);
and U4240 (N_4240,In_925,In_802);
nor U4241 (N_4241,In_264,In_558);
nor U4242 (N_4242,In_484,In_423);
or U4243 (N_4243,In_116,In_809);
nand U4244 (N_4244,In_183,In_372);
nor U4245 (N_4245,In_910,In_647);
or U4246 (N_4246,In_737,In_241);
nor U4247 (N_4247,In_866,In_388);
nor U4248 (N_4248,In_46,In_308);
and U4249 (N_4249,In_656,In_676);
xor U4250 (N_4250,In_804,In_485);
nor U4251 (N_4251,In_622,In_95);
or U4252 (N_4252,In_560,In_534);
and U4253 (N_4253,In_494,In_371);
and U4254 (N_4254,In_32,In_234);
xnor U4255 (N_4255,In_217,In_906);
nor U4256 (N_4256,In_638,In_781);
and U4257 (N_4257,In_152,In_645);
nor U4258 (N_4258,In_310,In_417);
nand U4259 (N_4259,In_940,In_904);
and U4260 (N_4260,In_62,In_733);
and U4261 (N_4261,In_48,In_550);
or U4262 (N_4262,In_215,In_395);
and U4263 (N_4263,In_381,In_968);
and U4264 (N_4264,In_874,In_146);
nand U4265 (N_4265,In_921,In_655);
nor U4266 (N_4266,In_701,In_8);
nand U4267 (N_4267,In_686,In_349);
and U4268 (N_4268,In_303,In_409);
xnor U4269 (N_4269,In_360,In_776);
or U4270 (N_4270,In_6,In_206);
nand U4271 (N_4271,In_61,In_967);
or U4272 (N_4272,In_492,In_462);
or U4273 (N_4273,In_249,In_990);
and U4274 (N_4274,In_857,In_700);
nand U4275 (N_4275,In_241,In_418);
or U4276 (N_4276,In_779,In_927);
nand U4277 (N_4277,In_199,In_744);
nor U4278 (N_4278,In_75,In_294);
nor U4279 (N_4279,In_967,In_421);
and U4280 (N_4280,In_659,In_554);
or U4281 (N_4281,In_572,In_585);
xnor U4282 (N_4282,In_797,In_913);
nor U4283 (N_4283,In_33,In_561);
xnor U4284 (N_4284,In_681,In_264);
and U4285 (N_4285,In_534,In_392);
nor U4286 (N_4286,In_267,In_921);
or U4287 (N_4287,In_648,In_9);
and U4288 (N_4288,In_73,In_671);
or U4289 (N_4289,In_706,In_389);
nand U4290 (N_4290,In_674,In_22);
nor U4291 (N_4291,In_20,In_3);
nand U4292 (N_4292,In_373,In_549);
nor U4293 (N_4293,In_179,In_934);
and U4294 (N_4294,In_123,In_931);
xor U4295 (N_4295,In_27,In_640);
or U4296 (N_4296,In_85,In_268);
and U4297 (N_4297,In_637,In_20);
nand U4298 (N_4298,In_511,In_309);
and U4299 (N_4299,In_658,In_481);
or U4300 (N_4300,In_252,In_405);
xor U4301 (N_4301,In_857,In_273);
nand U4302 (N_4302,In_394,In_71);
or U4303 (N_4303,In_585,In_909);
and U4304 (N_4304,In_815,In_685);
nand U4305 (N_4305,In_669,In_68);
or U4306 (N_4306,In_174,In_41);
or U4307 (N_4307,In_535,In_549);
nor U4308 (N_4308,In_921,In_218);
nand U4309 (N_4309,In_606,In_577);
or U4310 (N_4310,In_168,In_813);
nor U4311 (N_4311,In_447,In_768);
xor U4312 (N_4312,In_85,In_125);
and U4313 (N_4313,In_373,In_729);
nor U4314 (N_4314,In_804,In_775);
nor U4315 (N_4315,In_989,In_109);
and U4316 (N_4316,In_17,In_925);
and U4317 (N_4317,In_537,In_476);
nor U4318 (N_4318,In_947,In_518);
xnor U4319 (N_4319,In_262,In_737);
and U4320 (N_4320,In_58,In_622);
or U4321 (N_4321,In_272,In_342);
nor U4322 (N_4322,In_644,In_303);
nand U4323 (N_4323,In_75,In_74);
and U4324 (N_4324,In_526,In_401);
nor U4325 (N_4325,In_584,In_130);
nor U4326 (N_4326,In_590,In_157);
and U4327 (N_4327,In_197,In_180);
and U4328 (N_4328,In_844,In_766);
and U4329 (N_4329,In_86,In_949);
and U4330 (N_4330,In_338,In_889);
and U4331 (N_4331,In_152,In_853);
nor U4332 (N_4332,In_159,In_229);
nand U4333 (N_4333,In_728,In_985);
or U4334 (N_4334,In_49,In_903);
and U4335 (N_4335,In_51,In_379);
or U4336 (N_4336,In_944,In_165);
nor U4337 (N_4337,In_241,In_460);
nand U4338 (N_4338,In_299,In_523);
and U4339 (N_4339,In_906,In_486);
or U4340 (N_4340,In_921,In_101);
and U4341 (N_4341,In_317,In_815);
and U4342 (N_4342,In_633,In_373);
and U4343 (N_4343,In_40,In_680);
or U4344 (N_4344,In_32,In_263);
nand U4345 (N_4345,In_646,In_665);
and U4346 (N_4346,In_942,In_689);
or U4347 (N_4347,In_814,In_963);
nand U4348 (N_4348,In_855,In_930);
or U4349 (N_4349,In_480,In_255);
or U4350 (N_4350,In_412,In_240);
nand U4351 (N_4351,In_336,In_94);
and U4352 (N_4352,In_290,In_406);
xnor U4353 (N_4353,In_721,In_853);
nor U4354 (N_4354,In_340,In_879);
or U4355 (N_4355,In_787,In_263);
nor U4356 (N_4356,In_395,In_284);
xnor U4357 (N_4357,In_982,In_949);
nand U4358 (N_4358,In_102,In_130);
nand U4359 (N_4359,In_163,In_683);
and U4360 (N_4360,In_523,In_505);
or U4361 (N_4361,In_732,In_480);
and U4362 (N_4362,In_206,In_337);
and U4363 (N_4363,In_1,In_66);
xnor U4364 (N_4364,In_951,In_475);
or U4365 (N_4365,In_796,In_320);
or U4366 (N_4366,In_426,In_982);
nand U4367 (N_4367,In_103,In_127);
nand U4368 (N_4368,In_330,In_872);
and U4369 (N_4369,In_568,In_170);
nor U4370 (N_4370,In_719,In_961);
or U4371 (N_4371,In_642,In_486);
nor U4372 (N_4372,In_847,In_33);
nand U4373 (N_4373,In_984,In_139);
xnor U4374 (N_4374,In_281,In_923);
or U4375 (N_4375,In_586,In_242);
nand U4376 (N_4376,In_551,In_12);
and U4377 (N_4377,In_939,In_155);
or U4378 (N_4378,In_272,In_208);
nor U4379 (N_4379,In_871,In_72);
nor U4380 (N_4380,In_984,In_452);
nand U4381 (N_4381,In_2,In_273);
nand U4382 (N_4382,In_349,In_850);
nand U4383 (N_4383,In_296,In_538);
xnor U4384 (N_4384,In_132,In_20);
nand U4385 (N_4385,In_845,In_734);
nor U4386 (N_4386,In_292,In_728);
and U4387 (N_4387,In_241,In_28);
and U4388 (N_4388,In_637,In_405);
nor U4389 (N_4389,In_89,In_221);
and U4390 (N_4390,In_485,In_63);
or U4391 (N_4391,In_691,In_736);
nor U4392 (N_4392,In_294,In_642);
nand U4393 (N_4393,In_342,In_332);
xnor U4394 (N_4394,In_635,In_707);
or U4395 (N_4395,In_444,In_158);
nand U4396 (N_4396,In_832,In_161);
and U4397 (N_4397,In_193,In_98);
nor U4398 (N_4398,In_254,In_670);
or U4399 (N_4399,In_999,In_992);
nand U4400 (N_4400,In_268,In_236);
or U4401 (N_4401,In_482,In_844);
xnor U4402 (N_4402,In_614,In_481);
and U4403 (N_4403,In_19,In_302);
nor U4404 (N_4404,In_885,In_158);
xnor U4405 (N_4405,In_665,In_634);
nand U4406 (N_4406,In_133,In_468);
nand U4407 (N_4407,In_308,In_9);
or U4408 (N_4408,In_758,In_655);
or U4409 (N_4409,In_835,In_819);
xnor U4410 (N_4410,In_191,In_501);
nand U4411 (N_4411,In_613,In_841);
xnor U4412 (N_4412,In_551,In_188);
and U4413 (N_4413,In_487,In_512);
nand U4414 (N_4414,In_306,In_530);
nand U4415 (N_4415,In_430,In_972);
or U4416 (N_4416,In_851,In_116);
nand U4417 (N_4417,In_109,In_172);
nor U4418 (N_4418,In_680,In_49);
or U4419 (N_4419,In_721,In_90);
nand U4420 (N_4420,In_290,In_17);
nand U4421 (N_4421,In_995,In_996);
and U4422 (N_4422,In_503,In_395);
and U4423 (N_4423,In_183,In_639);
nor U4424 (N_4424,In_366,In_209);
or U4425 (N_4425,In_552,In_868);
nand U4426 (N_4426,In_936,In_330);
nand U4427 (N_4427,In_836,In_795);
and U4428 (N_4428,In_351,In_901);
or U4429 (N_4429,In_196,In_657);
or U4430 (N_4430,In_530,In_642);
or U4431 (N_4431,In_333,In_466);
nand U4432 (N_4432,In_952,In_605);
and U4433 (N_4433,In_328,In_711);
or U4434 (N_4434,In_292,In_969);
and U4435 (N_4435,In_762,In_178);
and U4436 (N_4436,In_382,In_717);
or U4437 (N_4437,In_662,In_242);
nor U4438 (N_4438,In_700,In_957);
nand U4439 (N_4439,In_780,In_186);
nand U4440 (N_4440,In_92,In_91);
and U4441 (N_4441,In_496,In_386);
nor U4442 (N_4442,In_938,In_556);
xnor U4443 (N_4443,In_90,In_697);
or U4444 (N_4444,In_769,In_831);
or U4445 (N_4445,In_456,In_136);
xor U4446 (N_4446,In_621,In_974);
nor U4447 (N_4447,In_613,In_800);
nand U4448 (N_4448,In_819,In_318);
xor U4449 (N_4449,In_153,In_163);
nand U4450 (N_4450,In_760,In_202);
or U4451 (N_4451,In_915,In_373);
or U4452 (N_4452,In_657,In_826);
nand U4453 (N_4453,In_218,In_444);
xor U4454 (N_4454,In_830,In_780);
or U4455 (N_4455,In_798,In_681);
nand U4456 (N_4456,In_258,In_495);
or U4457 (N_4457,In_20,In_611);
nand U4458 (N_4458,In_2,In_302);
nor U4459 (N_4459,In_794,In_1);
nand U4460 (N_4460,In_701,In_890);
nor U4461 (N_4461,In_190,In_978);
or U4462 (N_4462,In_158,In_69);
xor U4463 (N_4463,In_581,In_255);
nor U4464 (N_4464,In_599,In_941);
and U4465 (N_4465,In_38,In_943);
nor U4466 (N_4466,In_573,In_585);
and U4467 (N_4467,In_911,In_468);
nor U4468 (N_4468,In_302,In_637);
nor U4469 (N_4469,In_822,In_291);
nand U4470 (N_4470,In_772,In_629);
nand U4471 (N_4471,In_150,In_228);
nor U4472 (N_4472,In_565,In_690);
or U4473 (N_4473,In_76,In_458);
nand U4474 (N_4474,In_633,In_775);
nand U4475 (N_4475,In_232,In_451);
nand U4476 (N_4476,In_534,In_838);
or U4477 (N_4477,In_670,In_302);
xor U4478 (N_4478,In_374,In_379);
or U4479 (N_4479,In_110,In_639);
nand U4480 (N_4480,In_804,In_256);
or U4481 (N_4481,In_853,In_189);
nand U4482 (N_4482,In_372,In_572);
or U4483 (N_4483,In_879,In_757);
nor U4484 (N_4484,In_979,In_101);
nand U4485 (N_4485,In_178,In_737);
or U4486 (N_4486,In_585,In_145);
xnor U4487 (N_4487,In_929,In_359);
or U4488 (N_4488,In_278,In_839);
nand U4489 (N_4489,In_396,In_417);
nand U4490 (N_4490,In_535,In_774);
or U4491 (N_4491,In_702,In_475);
and U4492 (N_4492,In_811,In_169);
nor U4493 (N_4493,In_467,In_434);
xnor U4494 (N_4494,In_120,In_99);
nor U4495 (N_4495,In_593,In_706);
xnor U4496 (N_4496,In_280,In_320);
nand U4497 (N_4497,In_46,In_468);
nor U4498 (N_4498,In_603,In_910);
and U4499 (N_4499,In_531,In_466);
nor U4500 (N_4500,In_848,In_368);
nand U4501 (N_4501,In_629,In_270);
nand U4502 (N_4502,In_87,In_976);
nor U4503 (N_4503,In_343,In_85);
nand U4504 (N_4504,In_688,In_931);
xnor U4505 (N_4505,In_517,In_15);
or U4506 (N_4506,In_623,In_87);
or U4507 (N_4507,In_798,In_262);
or U4508 (N_4508,In_705,In_922);
or U4509 (N_4509,In_732,In_74);
xnor U4510 (N_4510,In_560,In_479);
nor U4511 (N_4511,In_301,In_670);
nor U4512 (N_4512,In_711,In_429);
nor U4513 (N_4513,In_195,In_982);
or U4514 (N_4514,In_635,In_574);
and U4515 (N_4515,In_366,In_129);
xnor U4516 (N_4516,In_138,In_527);
xnor U4517 (N_4517,In_577,In_397);
or U4518 (N_4518,In_711,In_875);
or U4519 (N_4519,In_566,In_70);
or U4520 (N_4520,In_38,In_45);
nand U4521 (N_4521,In_755,In_536);
nand U4522 (N_4522,In_521,In_141);
or U4523 (N_4523,In_683,In_919);
or U4524 (N_4524,In_927,In_642);
nand U4525 (N_4525,In_716,In_4);
nand U4526 (N_4526,In_777,In_584);
and U4527 (N_4527,In_912,In_323);
nand U4528 (N_4528,In_305,In_976);
nor U4529 (N_4529,In_937,In_307);
and U4530 (N_4530,In_611,In_542);
and U4531 (N_4531,In_521,In_49);
and U4532 (N_4532,In_328,In_645);
nor U4533 (N_4533,In_158,In_816);
or U4534 (N_4534,In_74,In_603);
nor U4535 (N_4535,In_492,In_370);
or U4536 (N_4536,In_120,In_762);
and U4537 (N_4537,In_597,In_169);
and U4538 (N_4538,In_503,In_648);
nand U4539 (N_4539,In_820,In_374);
nand U4540 (N_4540,In_488,In_371);
nor U4541 (N_4541,In_415,In_593);
or U4542 (N_4542,In_402,In_417);
nand U4543 (N_4543,In_911,In_125);
xnor U4544 (N_4544,In_391,In_126);
nand U4545 (N_4545,In_203,In_364);
nand U4546 (N_4546,In_171,In_511);
nor U4547 (N_4547,In_801,In_123);
or U4548 (N_4548,In_810,In_386);
and U4549 (N_4549,In_245,In_441);
or U4550 (N_4550,In_502,In_619);
or U4551 (N_4551,In_770,In_973);
nand U4552 (N_4552,In_114,In_581);
nor U4553 (N_4553,In_338,In_876);
nor U4554 (N_4554,In_105,In_428);
nand U4555 (N_4555,In_952,In_591);
nor U4556 (N_4556,In_682,In_443);
nand U4557 (N_4557,In_975,In_876);
or U4558 (N_4558,In_411,In_134);
and U4559 (N_4559,In_846,In_639);
nand U4560 (N_4560,In_509,In_988);
nand U4561 (N_4561,In_890,In_263);
and U4562 (N_4562,In_513,In_935);
or U4563 (N_4563,In_949,In_901);
nand U4564 (N_4564,In_17,In_613);
xnor U4565 (N_4565,In_367,In_174);
nor U4566 (N_4566,In_738,In_326);
nand U4567 (N_4567,In_890,In_731);
nand U4568 (N_4568,In_548,In_615);
nor U4569 (N_4569,In_618,In_629);
nand U4570 (N_4570,In_319,In_881);
nand U4571 (N_4571,In_85,In_199);
xor U4572 (N_4572,In_980,In_892);
xor U4573 (N_4573,In_953,In_135);
nand U4574 (N_4574,In_897,In_543);
and U4575 (N_4575,In_905,In_426);
nand U4576 (N_4576,In_888,In_885);
or U4577 (N_4577,In_920,In_549);
or U4578 (N_4578,In_28,In_910);
and U4579 (N_4579,In_780,In_45);
nand U4580 (N_4580,In_906,In_857);
nor U4581 (N_4581,In_157,In_488);
nor U4582 (N_4582,In_667,In_443);
and U4583 (N_4583,In_362,In_743);
and U4584 (N_4584,In_676,In_23);
xnor U4585 (N_4585,In_60,In_882);
and U4586 (N_4586,In_959,In_728);
and U4587 (N_4587,In_658,In_77);
nor U4588 (N_4588,In_972,In_1);
nand U4589 (N_4589,In_982,In_498);
xor U4590 (N_4590,In_63,In_591);
or U4591 (N_4591,In_819,In_858);
xnor U4592 (N_4592,In_658,In_798);
nand U4593 (N_4593,In_612,In_674);
nor U4594 (N_4594,In_618,In_871);
nor U4595 (N_4595,In_410,In_966);
or U4596 (N_4596,In_739,In_643);
and U4597 (N_4597,In_756,In_562);
xnor U4598 (N_4598,In_553,In_789);
nor U4599 (N_4599,In_101,In_638);
nor U4600 (N_4600,In_180,In_445);
nor U4601 (N_4601,In_249,In_979);
nand U4602 (N_4602,In_281,In_651);
nand U4603 (N_4603,In_825,In_287);
or U4604 (N_4604,In_782,In_903);
nor U4605 (N_4605,In_357,In_660);
nand U4606 (N_4606,In_873,In_648);
and U4607 (N_4607,In_855,In_969);
or U4608 (N_4608,In_150,In_356);
or U4609 (N_4609,In_98,In_880);
nand U4610 (N_4610,In_849,In_486);
and U4611 (N_4611,In_944,In_962);
and U4612 (N_4612,In_424,In_173);
nand U4613 (N_4613,In_53,In_83);
xor U4614 (N_4614,In_538,In_189);
nor U4615 (N_4615,In_374,In_332);
and U4616 (N_4616,In_125,In_126);
nand U4617 (N_4617,In_583,In_209);
or U4618 (N_4618,In_701,In_371);
nor U4619 (N_4619,In_229,In_993);
nor U4620 (N_4620,In_62,In_592);
nand U4621 (N_4621,In_143,In_197);
nor U4622 (N_4622,In_792,In_600);
nand U4623 (N_4623,In_925,In_788);
and U4624 (N_4624,In_787,In_111);
or U4625 (N_4625,In_161,In_10);
and U4626 (N_4626,In_21,In_5);
and U4627 (N_4627,In_529,In_151);
xor U4628 (N_4628,In_235,In_225);
nand U4629 (N_4629,In_432,In_141);
nor U4630 (N_4630,In_630,In_935);
xor U4631 (N_4631,In_473,In_863);
nand U4632 (N_4632,In_267,In_806);
and U4633 (N_4633,In_114,In_828);
nor U4634 (N_4634,In_63,In_227);
nor U4635 (N_4635,In_96,In_827);
or U4636 (N_4636,In_133,In_550);
nand U4637 (N_4637,In_35,In_580);
nand U4638 (N_4638,In_612,In_335);
nor U4639 (N_4639,In_988,In_680);
xor U4640 (N_4640,In_601,In_289);
xor U4641 (N_4641,In_889,In_703);
nand U4642 (N_4642,In_443,In_461);
nor U4643 (N_4643,In_237,In_368);
or U4644 (N_4644,In_920,In_509);
or U4645 (N_4645,In_460,In_692);
or U4646 (N_4646,In_272,In_171);
and U4647 (N_4647,In_372,In_597);
and U4648 (N_4648,In_640,In_470);
nand U4649 (N_4649,In_386,In_407);
and U4650 (N_4650,In_727,In_448);
or U4651 (N_4651,In_498,In_100);
nand U4652 (N_4652,In_948,In_264);
nand U4653 (N_4653,In_758,In_327);
or U4654 (N_4654,In_942,In_177);
xor U4655 (N_4655,In_509,In_174);
nand U4656 (N_4656,In_950,In_851);
nor U4657 (N_4657,In_463,In_318);
nand U4658 (N_4658,In_233,In_96);
or U4659 (N_4659,In_646,In_911);
nand U4660 (N_4660,In_848,In_924);
or U4661 (N_4661,In_282,In_722);
or U4662 (N_4662,In_577,In_972);
and U4663 (N_4663,In_712,In_629);
nor U4664 (N_4664,In_339,In_645);
xnor U4665 (N_4665,In_143,In_283);
nand U4666 (N_4666,In_238,In_825);
or U4667 (N_4667,In_703,In_621);
and U4668 (N_4668,In_123,In_697);
nor U4669 (N_4669,In_628,In_314);
nor U4670 (N_4670,In_428,In_814);
nand U4671 (N_4671,In_381,In_814);
and U4672 (N_4672,In_545,In_800);
or U4673 (N_4673,In_979,In_804);
and U4674 (N_4674,In_39,In_29);
or U4675 (N_4675,In_553,In_522);
or U4676 (N_4676,In_99,In_718);
nand U4677 (N_4677,In_839,In_13);
nor U4678 (N_4678,In_497,In_753);
or U4679 (N_4679,In_233,In_331);
nand U4680 (N_4680,In_949,In_802);
or U4681 (N_4681,In_609,In_719);
nor U4682 (N_4682,In_592,In_787);
xor U4683 (N_4683,In_181,In_142);
or U4684 (N_4684,In_155,In_895);
nor U4685 (N_4685,In_490,In_249);
nand U4686 (N_4686,In_655,In_520);
or U4687 (N_4687,In_458,In_493);
nor U4688 (N_4688,In_680,In_699);
xor U4689 (N_4689,In_99,In_640);
and U4690 (N_4690,In_825,In_607);
or U4691 (N_4691,In_735,In_286);
nand U4692 (N_4692,In_44,In_225);
and U4693 (N_4693,In_299,In_893);
nand U4694 (N_4694,In_369,In_411);
or U4695 (N_4695,In_17,In_493);
nand U4696 (N_4696,In_290,In_330);
nand U4697 (N_4697,In_800,In_409);
or U4698 (N_4698,In_759,In_705);
xor U4699 (N_4699,In_195,In_181);
or U4700 (N_4700,In_187,In_711);
and U4701 (N_4701,In_881,In_239);
nand U4702 (N_4702,In_39,In_480);
nor U4703 (N_4703,In_304,In_432);
and U4704 (N_4704,In_686,In_470);
and U4705 (N_4705,In_207,In_510);
and U4706 (N_4706,In_829,In_178);
or U4707 (N_4707,In_353,In_202);
xor U4708 (N_4708,In_751,In_383);
nor U4709 (N_4709,In_768,In_54);
nand U4710 (N_4710,In_576,In_427);
nand U4711 (N_4711,In_392,In_753);
and U4712 (N_4712,In_985,In_976);
nor U4713 (N_4713,In_151,In_704);
xor U4714 (N_4714,In_37,In_278);
and U4715 (N_4715,In_487,In_230);
nor U4716 (N_4716,In_699,In_550);
or U4717 (N_4717,In_933,In_353);
or U4718 (N_4718,In_718,In_63);
nor U4719 (N_4719,In_851,In_902);
nor U4720 (N_4720,In_774,In_101);
and U4721 (N_4721,In_765,In_250);
and U4722 (N_4722,In_259,In_941);
or U4723 (N_4723,In_911,In_596);
nor U4724 (N_4724,In_492,In_277);
or U4725 (N_4725,In_584,In_967);
or U4726 (N_4726,In_145,In_291);
or U4727 (N_4727,In_992,In_511);
xor U4728 (N_4728,In_766,In_821);
nor U4729 (N_4729,In_511,In_7);
nor U4730 (N_4730,In_976,In_990);
nor U4731 (N_4731,In_61,In_209);
nand U4732 (N_4732,In_888,In_155);
or U4733 (N_4733,In_730,In_782);
xor U4734 (N_4734,In_56,In_990);
and U4735 (N_4735,In_65,In_286);
nor U4736 (N_4736,In_823,In_51);
nor U4737 (N_4737,In_55,In_247);
nor U4738 (N_4738,In_330,In_508);
nand U4739 (N_4739,In_834,In_436);
or U4740 (N_4740,In_143,In_707);
nor U4741 (N_4741,In_180,In_701);
xor U4742 (N_4742,In_767,In_662);
xor U4743 (N_4743,In_630,In_686);
nand U4744 (N_4744,In_26,In_157);
nor U4745 (N_4745,In_842,In_846);
nand U4746 (N_4746,In_201,In_311);
xnor U4747 (N_4747,In_632,In_208);
and U4748 (N_4748,In_231,In_671);
nand U4749 (N_4749,In_147,In_705);
nand U4750 (N_4750,In_232,In_406);
nand U4751 (N_4751,In_71,In_381);
and U4752 (N_4752,In_975,In_166);
nand U4753 (N_4753,In_267,In_517);
and U4754 (N_4754,In_527,In_475);
and U4755 (N_4755,In_453,In_202);
and U4756 (N_4756,In_109,In_979);
or U4757 (N_4757,In_442,In_95);
or U4758 (N_4758,In_153,In_862);
nor U4759 (N_4759,In_70,In_974);
or U4760 (N_4760,In_811,In_384);
nand U4761 (N_4761,In_822,In_271);
nand U4762 (N_4762,In_759,In_475);
or U4763 (N_4763,In_178,In_989);
nor U4764 (N_4764,In_503,In_658);
or U4765 (N_4765,In_193,In_184);
nor U4766 (N_4766,In_287,In_546);
and U4767 (N_4767,In_311,In_183);
and U4768 (N_4768,In_880,In_489);
nand U4769 (N_4769,In_209,In_829);
nor U4770 (N_4770,In_676,In_400);
or U4771 (N_4771,In_782,In_14);
or U4772 (N_4772,In_876,In_687);
xor U4773 (N_4773,In_306,In_777);
nand U4774 (N_4774,In_313,In_57);
nand U4775 (N_4775,In_885,In_794);
nand U4776 (N_4776,In_787,In_151);
and U4777 (N_4777,In_743,In_95);
and U4778 (N_4778,In_757,In_159);
nand U4779 (N_4779,In_7,In_127);
or U4780 (N_4780,In_531,In_618);
and U4781 (N_4781,In_408,In_97);
or U4782 (N_4782,In_988,In_26);
or U4783 (N_4783,In_255,In_837);
nand U4784 (N_4784,In_268,In_214);
nand U4785 (N_4785,In_680,In_890);
and U4786 (N_4786,In_107,In_738);
nand U4787 (N_4787,In_942,In_350);
nand U4788 (N_4788,In_185,In_519);
nand U4789 (N_4789,In_601,In_454);
nand U4790 (N_4790,In_556,In_320);
nor U4791 (N_4791,In_973,In_361);
nor U4792 (N_4792,In_552,In_124);
nand U4793 (N_4793,In_620,In_237);
and U4794 (N_4794,In_862,In_314);
or U4795 (N_4795,In_290,In_974);
or U4796 (N_4796,In_958,In_289);
nor U4797 (N_4797,In_503,In_308);
nand U4798 (N_4798,In_450,In_550);
nor U4799 (N_4799,In_241,In_735);
nand U4800 (N_4800,In_642,In_363);
nor U4801 (N_4801,In_821,In_37);
and U4802 (N_4802,In_92,In_869);
nor U4803 (N_4803,In_638,In_962);
or U4804 (N_4804,In_691,In_302);
nor U4805 (N_4805,In_92,In_523);
and U4806 (N_4806,In_569,In_521);
and U4807 (N_4807,In_705,In_839);
nor U4808 (N_4808,In_264,In_609);
and U4809 (N_4809,In_353,In_954);
or U4810 (N_4810,In_262,In_990);
or U4811 (N_4811,In_934,In_998);
nor U4812 (N_4812,In_722,In_706);
xnor U4813 (N_4813,In_208,In_338);
xor U4814 (N_4814,In_418,In_163);
nand U4815 (N_4815,In_671,In_980);
nand U4816 (N_4816,In_488,In_429);
nor U4817 (N_4817,In_570,In_473);
or U4818 (N_4818,In_928,In_154);
nor U4819 (N_4819,In_273,In_672);
and U4820 (N_4820,In_22,In_205);
or U4821 (N_4821,In_251,In_996);
or U4822 (N_4822,In_524,In_781);
or U4823 (N_4823,In_104,In_284);
nand U4824 (N_4824,In_947,In_892);
nor U4825 (N_4825,In_370,In_522);
nor U4826 (N_4826,In_466,In_550);
nor U4827 (N_4827,In_336,In_585);
nand U4828 (N_4828,In_428,In_732);
or U4829 (N_4829,In_918,In_632);
or U4830 (N_4830,In_194,In_564);
or U4831 (N_4831,In_750,In_562);
nand U4832 (N_4832,In_368,In_883);
nor U4833 (N_4833,In_51,In_806);
or U4834 (N_4834,In_355,In_747);
nor U4835 (N_4835,In_69,In_527);
and U4836 (N_4836,In_675,In_982);
nor U4837 (N_4837,In_662,In_396);
nand U4838 (N_4838,In_609,In_305);
nor U4839 (N_4839,In_273,In_811);
and U4840 (N_4840,In_215,In_284);
or U4841 (N_4841,In_321,In_956);
nand U4842 (N_4842,In_454,In_470);
and U4843 (N_4843,In_792,In_165);
and U4844 (N_4844,In_55,In_126);
nand U4845 (N_4845,In_131,In_477);
nor U4846 (N_4846,In_294,In_960);
and U4847 (N_4847,In_121,In_625);
nor U4848 (N_4848,In_243,In_700);
or U4849 (N_4849,In_883,In_196);
nor U4850 (N_4850,In_603,In_89);
xnor U4851 (N_4851,In_603,In_936);
and U4852 (N_4852,In_128,In_90);
and U4853 (N_4853,In_14,In_224);
nor U4854 (N_4854,In_384,In_518);
nor U4855 (N_4855,In_151,In_491);
nor U4856 (N_4856,In_428,In_922);
and U4857 (N_4857,In_912,In_594);
nand U4858 (N_4858,In_638,In_909);
and U4859 (N_4859,In_482,In_177);
or U4860 (N_4860,In_258,In_673);
or U4861 (N_4861,In_824,In_550);
nand U4862 (N_4862,In_999,In_124);
nand U4863 (N_4863,In_968,In_764);
nand U4864 (N_4864,In_798,In_165);
or U4865 (N_4865,In_542,In_690);
nor U4866 (N_4866,In_128,In_264);
xor U4867 (N_4867,In_145,In_664);
nand U4868 (N_4868,In_180,In_199);
nand U4869 (N_4869,In_212,In_373);
or U4870 (N_4870,In_456,In_439);
nand U4871 (N_4871,In_527,In_388);
and U4872 (N_4872,In_667,In_709);
and U4873 (N_4873,In_716,In_148);
nor U4874 (N_4874,In_846,In_986);
or U4875 (N_4875,In_209,In_633);
nand U4876 (N_4876,In_356,In_343);
nor U4877 (N_4877,In_341,In_991);
nor U4878 (N_4878,In_445,In_361);
nand U4879 (N_4879,In_332,In_949);
or U4880 (N_4880,In_649,In_628);
xor U4881 (N_4881,In_905,In_878);
or U4882 (N_4882,In_607,In_756);
nand U4883 (N_4883,In_755,In_123);
or U4884 (N_4884,In_517,In_92);
nor U4885 (N_4885,In_378,In_242);
nand U4886 (N_4886,In_354,In_522);
xor U4887 (N_4887,In_617,In_267);
and U4888 (N_4888,In_539,In_546);
nand U4889 (N_4889,In_270,In_406);
nand U4890 (N_4890,In_296,In_24);
and U4891 (N_4891,In_348,In_779);
and U4892 (N_4892,In_507,In_451);
nor U4893 (N_4893,In_201,In_764);
nand U4894 (N_4894,In_991,In_601);
nor U4895 (N_4895,In_518,In_504);
nand U4896 (N_4896,In_787,In_349);
nand U4897 (N_4897,In_829,In_493);
and U4898 (N_4898,In_71,In_768);
or U4899 (N_4899,In_880,In_540);
xor U4900 (N_4900,In_981,In_572);
and U4901 (N_4901,In_810,In_342);
nand U4902 (N_4902,In_29,In_89);
and U4903 (N_4903,In_124,In_621);
xnor U4904 (N_4904,In_178,In_729);
nand U4905 (N_4905,In_688,In_954);
nand U4906 (N_4906,In_879,In_103);
xnor U4907 (N_4907,In_686,In_273);
nand U4908 (N_4908,In_342,In_378);
and U4909 (N_4909,In_770,In_178);
and U4910 (N_4910,In_796,In_478);
nor U4911 (N_4911,In_208,In_170);
or U4912 (N_4912,In_13,In_835);
nor U4913 (N_4913,In_570,In_910);
nor U4914 (N_4914,In_898,In_886);
xor U4915 (N_4915,In_445,In_592);
nor U4916 (N_4916,In_51,In_975);
or U4917 (N_4917,In_965,In_53);
or U4918 (N_4918,In_766,In_331);
and U4919 (N_4919,In_505,In_540);
nor U4920 (N_4920,In_407,In_719);
and U4921 (N_4921,In_593,In_963);
or U4922 (N_4922,In_574,In_732);
nor U4923 (N_4923,In_42,In_862);
nor U4924 (N_4924,In_642,In_547);
and U4925 (N_4925,In_83,In_788);
or U4926 (N_4926,In_716,In_516);
xnor U4927 (N_4927,In_749,In_21);
nand U4928 (N_4928,In_531,In_689);
nand U4929 (N_4929,In_939,In_386);
and U4930 (N_4930,In_14,In_130);
nand U4931 (N_4931,In_631,In_110);
nor U4932 (N_4932,In_166,In_411);
or U4933 (N_4933,In_900,In_759);
and U4934 (N_4934,In_435,In_676);
nand U4935 (N_4935,In_774,In_122);
nand U4936 (N_4936,In_22,In_43);
nor U4937 (N_4937,In_859,In_141);
nor U4938 (N_4938,In_666,In_474);
nor U4939 (N_4939,In_234,In_637);
and U4940 (N_4940,In_523,In_404);
and U4941 (N_4941,In_400,In_140);
and U4942 (N_4942,In_143,In_594);
and U4943 (N_4943,In_458,In_58);
and U4944 (N_4944,In_943,In_821);
or U4945 (N_4945,In_681,In_754);
nor U4946 (N_4946,In_349,In_93);
nor U4947 (N_4947,In_507,In_286);
nand U4948 (N_4948,In_669,In_223);
nand U4949 (N_4949,In_869,In_410);
nand U4950 (N_4950,In_137,In_617);
nor U4951 (N_4951,In_968,In_211);
xor U4952 (N_4952,In_804,In_779);
or U4953 (N_4953,In_876,In_906);
xor U4954 (N_4954,In_633,In_806);
nor U4955 (N_4955,In_786,In_201);
nor U4956 (N_4956,In_116,In_240);
nand U4957 (N_4957,In_188,In_230);
and U4958 (N_4958,In_824,In_169);
or U4959 (N_4959,In_967,In_683);
xnor U4960 (N_4960,In_650,In_1);
and U4961 (N_4961,In_8,In_195);
and U4962 (N_4962,In_979,In_274);
or U4963 (N_4963,In_19,In_700);
or U4964 (N_4964,In_327,In_133);
xnor U4965 (N_4965,In_311,In_223);
nand U4966 (N_4966,In_859,In_711);
nand U4967 (N_4967,In_70,In_859);
and U4968 (N_4968,In_129,In_879);
nor U4969 (N_4969,In_473,In_896);
xnor U4970 (N_4970,In_226,In_331);
and U4971 (N_4971,In_539,In_342);
nand U4972 (N_4972,In_434,In_652);
nor U4973 (N_4973,In_983,In_132);
or U4974 (N_4974,In_50,In_53);
or U4975 (N_4975,In_538,In_410);
or U4976 (N_4976,In_362,In_672);
and U4977 (N_4977,In_72,In_843);
and U4978 (N_4978,In_275,In_220);
nor U4979 (N_4979,In_816,In_729);
nor U4980 (N_4980,In_790,In_593);
or U4981 (N_4981,In_758,In_425);
nor U4982 (N_4982,In_190,In_54);
nand U4983 (N_4983,In_324,In_607);
and U4984 (N_4984,In_180,In_669);
or U4985 (N_4985,In_809,In_747);
nor U4986 (N_4986,In_777,In_687);
or U4987 (N_4987,In_293,In_362);
nand U4988 (N_4988,In_948,In_302);
nand U4989 (N_4989,In_113,In_640);
nand U4990 (N_4990,In_887,In_186);
nand U4991 (N_4991,In_43,In_692);
nor U4992 (N_4992,In_923,In_598);
nand U4993 (N_4993,In_247,In_520);
nor U4994 (N_4994,In_857,In_196);
nor U4995 (N_4995,In_747,In_926);
or U4996 (N_4996,In_870,In_447);
nor U4997 (N_4997,In_788,In_314);
and U4998 (N_4998,In_772,In_178);
nor U4999 (N_4999,In_189,In_787);
nor U5000 (N_5000,N_4300,N_3536);
nor U5001 (N_5001,N_825,N_2578);
nor U5002 (N_5002,N_66,N_3141);
xor U5003 (N_5003,N_4036,N_103);
xnor U5004 (N_5004,N_1620,N_1107);
nand U5005 (N_5005,N_4780,N_4314);
nor U5006 (N_5006,N_2840,N_4157);
or U5007 (N_5007,N_4202,N_4845);
nand U5008 (N_5008,N_2235,N_4915);
and U5009 (N_5009,N_4925,N_2271);
nor U5010 (N_5010,N_1284,N_2830);
and U5011 (N_5011,N_2947,N_2749);
or U5012 (N_5012,N_4909,N_4969);
nand U5013 (N_5013,N_2801,N_55);
and U5014 (N_5014,N_1964,N_4751);
and U5015 (N_5015,N_2706,N_2890);
nand U5016 (N_5016,N_3028,N_2435);
or U5017 (N_5017,N_2077,N_1338);
or U5018 (N_5018,N_2061,N_1318);
and U5019 (N_5019,N_4907,N_4930);
and U5020 (N_5020,N_4076,N_683);
or U5021 (N_5021,N_119,N_1669);
nor U5022 (N_5022,N_3009,N_1151);
and U5023 (N_5023,N_2392,N_433);
nand U5024 (N_5024,N_4298,N_4114);
xnor U5025 (N_5025,N_1981,N_243);
and U5026 (N_5026,N_3645,N_1659);
and U5027 (N_5027,N_960,N_2754);
nor U5028 (N_5028,N_1008,N_2227);
or U5029 (N_5029,N_2680,N_740);
nand U5030 (N_5030,N_2695,N_1883);
or U5031 (N_5031,N_3820,N_4272);
xor U5032 (N_5032,N_4978,N_4492);
nand U5033 (N_5033,N_3755,N_4828);
and U5034 (N_5034,N_1242,N_2218);
nor U5035 (N_5035,N_3867,N_4107);
and U5036 (N_5036,N_1900,N_4830);
or U5037 (N_5037,N_2582,N_3802);
xnor U5038 (N_5038,N_298,N_981);
and U5039 (N_5039,N_859,N_478);
nor U5040 (N_5040,N_841,N_809);
or U5041 (N_5041,N_141,N_2849);
xor U5042 (N_5042,N_4123,N_2716);
nand U5043 (N_5043,N_3231,N_1511);
nand U5044 (N_5044,N_1878,N_4186);
nand U5045 (N_5045,N_2318,N_2779);
nor U5046 (N_5046,N_4769,N_4678);
nor U5047 (N_5047,N_2389,N_3853);
nor U5048 (N_5048,N_3881,N_4718);
and U5049 (N_5049,N_2599,N_336);
or U5050 (N_5050,N_1592,N_1279);
nand U5051 (N_5051,N_308,N_1481);
and U5052 (N_5052,N_705,N_1798);
nor U5053 (N_5053,N_768,N_2675);
and U5054 (N_5054,N_1618,N_515);
xor U5055 (N_5055,N_4180,N_914);
nand U5056 (N_5056,N_3520,N_2222);
nand U5057 (N_5057,N_2597,N_1321);
and U5058 (N_5058,N_4367,N_3087);
and U5059 (N_5059,N_2642,N_3830);
xor U5060 (N_5060,N_4928,N_4343);
and U5061 (N_5061,N_3162,N_2751);
or U5062 (N_5062,N_2100,N_3457);
or U5063 (N_5063,N_1055,N_3551);
nand U5064 (N_5064,N_588,N_164);
nor U5065 (N_5065,N_1624,N_1771);
nand U5066 (N_5066,N_4619,N_1577);
xor U5067 (N_5067,N_3003,N_48);
nor U5068 (N_5068,N_3968,N_4248);
xnor U5069 (N_5069,N_2797,N_647);
or U5070 (N_5070,N_4998,N_1498);
or U5071 (N_5071,N_2044,N_4420);
nor U5072 (N_5072,N_871,N_12);
and U5073 (N_5073,N_1012,N_4456);
and U5074 (N_5074,N_3217,N_3743);
and U5075 (N_5075,N_2027,N_4785);
or U5076 (N_5076,N_2478,N_310);
nor U5077 (N_5077,N_1038,N_2861);
nor U5078 (N_5078,N_4699,N_3390);
nor U5079 (N_5079,N_1475,N_1575);
and U5080 (N_5080,N_3490,N_4220);
or U5081 (N_5081,N_2062,N_4446);
nor U5082 (N_5082,N_3796,N_4439);
xnor U5083 (N_5083,N_3602,N_701);
xnor U5084 (N_5084,N_3074,N_4084);
nor U5085 (N_5085,N_2055,N_2626);
nor U5086 (N_5086,N_4233,N_4745);
and U5087 (N_5087,N_2732,N_189);
or U5088 (N_5088,N_4566,N_1422);
and U5089 (N_5089,N_74,N_2750);
and U5090 (N_5090,N_2358,N_3903);
nand U5091 (N_5091,N_681,N_4245);
and U5092 (N_5092,N_4029,N_4074);
and U5093 (N_5093,N_96,N_4861);
nor U5094 (N_5094,N_3303,N_1786);
or U5095 (N_5095,N_1921,N_2829);
nor U5096 (N_5096,N_1464,N_542);
nor U5097 (N_5097,N_338,N_4093);
nor U5098 (N_5098,N_3666,N_88);
xor U5099 (N_5099,N_3173,N_673);
xor U5100 (N_5100,N_3384,N_679);
nand U5101 (N_5101,N_2878,N_659);
or U5102 (N_5102,N_709,N_3203);
or U5103 (N_5103,N_4708,N_180);
xor U5104 (N_5104,N_3160,N_3764);
or U5105 (N_5105,N_3437,N_3077);
nand U5106 (N_5106,N_2004,N_885);
or U5107 (N_5107,N_1500,N_2333);
and U5108 (N_5108,N_4646,N_2494);
nand U5109 (N_5109,N_4428,N_1846);
and U5110 (N_5110,N_3569,N_2303);
and U5111 (N_5111,N_75,N_3603);
or U5112 (N_5112,N_1101,N_2408);
nor U5113 (N_5113,N_2980,N_2361);
nor U5114 (N_5114,N_3516,N_1104);
and U5115 (N_5115,N_4473,N_3783);
and U5116 (N_5116,N_3326,N_64);
or U5117 (N_5117,N_1065,N_4696);
or U5118 (N_5118,N_735,N_4421);
or U5119 (N_5119,N_4673,N_1587);
or U5120 (N_5120,N_3518,N_100);
xnor U5121 (N_5121,N_1303,N_2451);
or U5122 (N_5122,N_1427,N_2356);
nor U5123 (N_5123,N_3115,N_4020);
xor U5124 (N_5124,N_2773,N_4972);
nand U5125 (N_5125,N_778,N_585);
or U5126 (N_5126,N_4787,N_1120);
nand U5127 (N_5127,N_3492,N_1354);
nor U5128 (N_5128,N_2782,N_2531);
xnor U5129 (N_5129,N_961,N_2199);
and U5130 (N_5130,N_4382,N_1632);
and U5131 (N_5131,N_2638,N_221);
nand U5132 (N_5132,N_34,N_566);
nand U5133 (N_5133,N_2817,N_2762);
and U5134 (N_5134,N_1257,N_3543);
or U5135 (N_5135,N_3133,N_3715);
or U5136 (N_5136,N_3404,N_4395);
nor U5137 (N_5137,N_1619,N_3273);
and U5138 (N_5138,N_2121,N_4803);
nand U5139 (N_5139,N_1488,N_1424);
or U5140 (N_5140,N_4565,N_1175);
and U5141 (N_5141,N_3910,N_574);
nand U5142 (N_5142,N_1829,N_1789);
nor U5143 (N_5143,N_4752,N_4539);
or U5144 (N_5144,N_4135,N_3630);
or U5145 (N_5145,N_2264,N_986);
xor U5146 (N_5146,N_3675,N_3729);
or U5147 (N_5147,N_1081,N_3546);
nor U5148 (N_5148,N_3294,N_2288);
nand U5149 (N_5149,N_1368,N_3271);
nor U5150 (N_5150,N_1899,N_4410);
xor U5151 (N_5151,N_1979,N_2009);
nor U5152 (N_5152,N_3264,N_1409);
and U5153 (N_5153,N_2988,N_3894);
or U5154 (N_5154,N_155,N_3926);
and U5155 (N_5155,N_4003,N_3387);
or U5156 (N_5156,N_2050,N_4683);
xor U5157 (N_5157,N_4187,N_2180);
and U5158 (N_5158,N_4797,N_3613);
or U5159 (N_5159,N_4130,N_2761);
nand U5160 (N_5160,N_280,N_3928);
nor U5161 (N_5161,N_4090,N_995);
and U5162 (N_5162,N_3989,N_3493);
and U5163 (N_5163,N_4488,N_2804);
nand U5164 (N_5164,N_2034,N_3459);
or U5165 (N_5165,N_2606,N_3506);
xor U5166 (N_5166,N_1664,N_2129);
nor U5167 (N_5167,N_2322,N_2882);
xnor U5168 (N_5168,N_4618,N_2542);
xnor U5169 (N_5169,N_4838,N_600);
xor U5170 (N_5170,N_2313,N_219);
nand U5171 (N_5171,N_4945,N_1485);
nand U5172 (N_5172,N_1643,N_117);
nor U5173 (N_5173,N_1429,N_4481);
or U5174 (N_5174,N_4217,N_983);
nand U5175 (N_5175,N_3904,N_229);
or U5176 (N_5176,N_1689,N_4363);
or U5177 (N_5177,N_2336,N_804);
and U5178 (N_5178,N_651,N_3931);
and U5179 (N_5179,N_370,N_822);
or U5180 (N_5180,N_4124,N_1646);
or U5181 (N_5181,N_1755,N_2390);
nor U5182 (N_5182,N_4760,N_1902);
xnor U5183 (N_5183,N_1513,N_1336);
xor U5184 (N_5184,N_3727,N_3447);
or U5185 (N_5185,N_2427,N_3611);
nor U5186 (N_5186,N_1987,N_2268);
nor U5187 (N_5187,N_4538,N_10);
and U5188 (N_5188,N_3591,N_1521);
or U5189 (N_5189,N_1613,N_2753);
and U5190 (N_5190,N_2039,N_4564);
nand U5191 (N_5191,N_2848,N_4424);
or U5192 (N_5192,N_1199,N_4598);
nor U5193 (N_5193,N_2431,N_1074);
and U5194 (N_5194,N_739,N_4772);
or U5195 (N_5195,N_4811,N_1732);
and U5196 (N_5196,N_1770,N_4281);
or U5197 (N_5197,N_2790,N_4562);
nand U5198 (N_5198,N_2473,N_3251);
xnor U5199 (N_5199,N_447,N_3892);
and U5200 (N_5200,N_1070,N_2700);
nand U5201 (N_5201,N_948,N_3138);
and U5202 (N_5202,N_3348,N_4523);
and U5203 (N_5203,N_3161,N_3239);
nand U5204 (N_5204,N_4170,N_1041);
nor U5205 (N_5205,N_1538,N_4094);
nor U5206 (N_5206,N_837,N_4019);
or U5207 (N_5207,N_704,N_1092);
nand U5208 (N_5208,N_3011,N_1911);
xor U5209 (N_5209,N_20,N_3572);
or U5210 (N_5210,N_3915,N_248);
xnor U5211 (N_5211,N_3062,N_3131);
nor U5212 (N_5212,N_1,N_213);
nand U5213 (N_5213,N_2933,N_95);
nor U5214 (N_5214,N_4137,N_3396);
nand U5215 (N_5215,N_76,N_2438);
or U5216 (N_5216,N_776,N_1989);
or U5217 (N_5217,N_874,N_4905);
nor U5218 (N_5218,N_2065,N_2331);
or U5219 (N_5219,N_388,N_138);
and U5220 (N_5220,N_3866,N_953);
or U5221 (N_5221,N_4415,N_350);
or U5222 (N_5222,N_4471,N_4832);
or U5223 (N_5223,N_4406,N_2622);
and U5224 (N_5224,N_4489,N_2654);
and U5225 (N_5225,N_156,N_1774);
or U5226 (N_5226,N_2735,N_1130);
nand U5227 (N_5227,N_1119,N_2202);
nand U5228 (N_5228,N_2673,N_431);
nand U5229 (N_5229,N_4364,N_3500);
xnor U5230 (N_5230,N_2902,N_2784);
nor U5231 (N_5231,N_1332,N_603);
nor U5232 (N_5232,N_254,N_4666);
nor U5233 (N_5233,N_183,N_2080);
nor U5234 (N_5234,N_3746,N_2175);
nand U5235 (N_5235,N_246,N_2592);
and U5236 (N_5236,N_3091,N_937);
nand U5237 (N_5237,N_4041,N_4937);
or U5238 (N_5238,N_3697,N_4596);
nor U5239 (N_5239,N_3609,N_3412);
nor U5240 (N_5240,N_1502,N_4606);
nand U5241 (N_5241,N_1398,N_1723);
or U5242 (N_5242,N_777,N_3884);
nor U5243 (N_5243,N_589,N_207);
and U5244 (N_5244,N_3106,N_1173);
and U5245 (N_5245,N_662,N_621);
nand U5246 (N_5246,N_576,N_4691);
nor U5247 (N_5247,N_4150,N_2049);
nand U5248 (N_5248,N_907,N_167);
or U5249 (N_5249,N_2704,N_3982);
and U5250 (N_5250,N_1423,N_4740);
or U5251 (N_5251,N_3125,N_2772);
or U5252 (N_5252,N_4502,N_4262);
nor U5253 (N_5253,N_4639,N_3973);
nor U5254 (N_5254,N_3403,N_4286);
and U5255 (N_5255,N_2748,N_1458);
and U5256 (N_5256,N_1048,N_2411);
and U5257 (N_5257,N_1831,N_4112);
and U5258 (N_5258,N_340,N_4008);
xnor U5259 (N_5259,N_2418,N_3810);
nand U5260 (N_5260,N_2153,N_3004);
or U5261 (N_5261,N_1684,N_2041);
and U5262 (N_5262,N_3799,N_65);
nor U5263 (N_5263,N_3248,N_928);
or U5264 (N_5264,N_4269,N_4109);
or U5265 (N_5265,N_3886,N_4843);
nand U5266 (N_5266,N_3128,N_2724);
nor U5267 (N_5267,N_1054,N_3332);
and U5268 (N_5268,N_1016,N_4818);
nand U5269 (N_5269,N_4503,N_4764);
nor U5270 (N_5270,N_1061,N_2926);
xnor U5271 (N_5271,N_611,N_3013);
nand U5272 (N_5272,N_2688,N_1761);
and U5273 (N_5273,N_1383,N_35);
or U5274 (N_5274,N_1133,N_1713);
or U5275 (N_5275,N_2628,N_2396);
nand U5276 (N_5276,N_4403,N_3455);
or U5277 (N_5277,N_2170,N_4700);
nand U5278 (N_5278,N_1790,N_4743);
xnor U5279 (N_5279,N_3998,N_4999);
nor U5280 (N_5280,N_1030,N_3537);
nor U5281 (N_5281,N_2279,N_3379);
xnor U5282 (N_5282,N_4080,N_2526);
xor U5283 (N_5283,N_1071,N_374);
and U5284 (N_5284,N_4354,N_3045);
nand U5285 (N_5285,N_1014,N_4859);
xor U5286 (N_5286,N_2831,N_1394);
nand U5287 (N_5287,N_4432,N_1180);
and U5288 (N_5288,N_2629,N_2160);
or U5289 (N_5289,N_251,N_2646);
nand U5290 (N_5290,N_2737,N_4579);
nand U5291 (N_5291,N_1589,N_3357);
or U5292 (N_5292,N_2037,N_3834);
and U5293 (N_5293,N_1265,N_1088);
nor U5294 (N_5294,N_3535,N_2904);
and U5295 (N_5295,N_538,N_4345);
and U5296 (N_5296,N_4814,N_1859);
and U5297 (N_5297,N_1652,N_2480);
or U5298 (N_5298,N_3556,N_2777);
nor U5299 (N_5299,N_372,N_1706);
or U5300 (N_5300,N_4973,N_2021);
nand U5301 (N_5301,N_2856,N_17);
and U5302 (N_5302,N_4512,N_3777);
or U5303 (N_5303,N_1693,N_3132);
nand U5304 (N_5304,N_1904,N_2962);
or U5305 (N_5305,N_1748,N_583);
or U5306 (N_5306,N_2569,N_2419);
nand U5307 (N_5307,N_2945,N_1200);
nor U5308 (N_5308,N_4440,N_2108);
nand U5309 (N_5309,N_800,N_3078);
and U5310 (N_5310,N_2891,N_4813);
and U5311 (N_5311,N_2920,N_3519);
nand U5312 (N_5312,N_3021,N_1945);
nor U5313 (N_5313,N_2138,N_972);
or U5314 (N_5314,N_556,N_2449);
nor U5315 (N_5315,N_362,N_429);
nor U5316 (N_5316,N_214,N_1600);
xor U5317 (N_5317,N_792,N_911);
nand U5318 (N_5318,N_3615,N_2415);
and U5319 (N_5319,N_2457,N_4060);
or U5320 (N_5320,N_326,N_3598);
and U5321 (N_5321,N_2959,N_1611);
nand U5322 (N_5322,N_2059,N_2566);
nand U5323 (N_5323,N_1740,N_965);
or U5324 (N_5324,N_4480,N_1949);
or U5325 (N_5325,N_4891,N_3210);
or U5326 (N_5326,N_1416,N_411);
or U5327 (N_5327,N_4274,N_1157);
and U5328 (N_5328,N_1868,N_3147);
nor U5329 (N_5329,N_1305,N_2917);
or U5330 (N_5330,N_268,N_504);
xnor U5331 (N_5331,N_263,N_2583);
nand U5332 (N_5332,N_4347,N_4111);
xnor U5333 (N_5333,N_820,N_3056);
and U5334 (N_5334,N_2354,N_945);
and U5335 (N_5335,N_3552,N_4950);
nor U5336 (N_5336,N_2952,N_4352);
nor U5337 (N_5337,N_3135,N_1818);
nand U5338 (N_5338,N_4848,N_771);
xor U5339 (N_5339,N_3568,N_2019);
and U5340 (N_5340,N_4253,N_3737);
nor U5341 (N_5341,N_4311,N_3891);
or U5342 (N_5342,N_2212,N_4321);
and U5343 (N_5343,N_2384,N_2922);
and U5344 (N_5344,N_618,N_1298);
or U5345 (N_5345,N_3902,N_1596);
and U5346 (N_5346,N_1391,N_3564);
or U5347 (N_5347,N_876,N_1780);
and U5348 (N_5348,N_4990,N_1308);
or U5349 (N_5349,N_667,N_3143);
xnor U5350 (N_5350,N_2052,N_79);
and U5351 (N_5351,N_4318,N_32);
nor U5352 (N_5352,N_1544,N_4851);
or U5353 (N_5353,N_3880,N_3649);
or U5354 (N_5354,N_1626,N_3157);
and U5355 (N_5355,N_456,N_3084);
nor U5356 (N_5356,N_3213,N_2176);
nor U5357 (N_5357,N_4301,N_4603);
nand U5358 (N_5358,N_743,N_40);
nor U5359 (N_5359,N_1349,N_4510);
or U5360 (N_5360,N_2293,N_368);
nand U5361 (N_5361,N_4991,N_1374);
xor U5362 (N_5362,N_2247,N_3607);
or U5363 (N_5363,N_4337,N_4534);
xnor U5364 (N_5364,N_135,N_2819);
nand U5365 (N_5365,N_307,N_1466);
or U5366 (N_5366,N_1816,N_657);
or U5367 (N_5367,N_2672,N_3789);
nand U5368 (N_5368,N_2366,N_4936);
or U5369 (N_5369,N_81,N_1648);
nand U5370 (N_5370,N_787,N_4864);
or U5371 (N_5371,N_969,N_3751);
or U5372 (N_5372,N_1205,N_325);
and U5373 (N_5373,N_2679,N_3662);
or U5374 (N_5374,N_3495,N_3585);
or U5375 (N_5375,N_3408,N_2066);
or U5376 (N_5376,N_639,N_3150);
nor U5377 (N_5377,N_2107,N_4374);
and U5378 (N_5378,N_4667,N_3494);
or U5379 (N_5379,N_2444,N_2346);
nor U5380 (N_5380,N_3193,N_3024);
or U5381 (N_5381,N_4784,N_3612);
or U5382 (N_5382,N_4616,N_4079);
nor U5383 (N_5383,N_567,N_4684);
nand U5384 (N_5384,N_2181,N_1275);
or U5385 (N_5385,N_1559,N_2025);
or U5386 (N_5386,N_4874,N_4887);
nand U5387 (N_5387,N_2368,N_554);
xor U5388 (N_5388,N_2728,N_1845);
nor U5389 (N_5389,N_3320,N_1033);
or U5390 (N_5390,N_1627,N_3824);
or U5391 (N_5391,N_966,N_199);
and U5392 (N_5392,N_2868,N_1395);
xnor U5393 (N_5393,N_4983,N_4569);
and U5394 (N_5394,N_2490,N_185);
or U5395 (N_5395,N_1389,N_1467);
xnor U5396 (N_5396,N_1941,N_2571);
or U5397 (N_5397,N_3686,N_1884);
or U5398 (N_5398,N_3323,N_2375);
and U5399 (N_5399,N_4230,N_4108);
nor U5400 (N_5400,N_4445,N_3184);
nand U5401 (N_5401,N_4641,N_4899);
nor U5402 (N_5402,N_4712,N_2854);
nor U5403 (N_5403,N_3502,N_3855);
or U5404 (N_5404,N_1834,N_118);
and U5405 (N_5405,N_1730,N_2452);
and U5406 (N_5406,N_3907,N_4304);
xnor U5407 (N_5407,N_606,N_4372);
nor U5408 (N_5408,N_4017,N_1892);
or U5409 (N_5409,N_3345,N_2095);
xor U5410 (N_5410,N_4576,N_3792);
nand U5411 (N_5411,N_3971,N_4654);
xor U5412 (N_5412,N_3767,N_2953);
nand U5413 (N_5413,N_1929,N_2506);
and U5414 (N_5414,N_1714,N_2570);
xnor U5415 (N_5415,N_4102,N_3095);
xnor U5416 (N_5416,N_430,N_46);
nand U5417 (N_5417,N_2832,N_3623);
and U5418 (N_5418,N_3626,N_828);
xor U5419 (N_5419,N_1810,N_2696);
or U5420 (N_5420,N_4185,N_3875);
or U5421 (N_5421,N_2230,N_2267);
or U5422 (N_5422,N_3822,N_4160);
xor U5423 (N_5423,N_3139,N_755);
nor U5424 (N_5424,N_3680,N_198);
and U5425 (N_5425,N_3298,N_1348);
and U5426 (N_5426,N_730,N_1392);
nor U5427 (N_5427,N_292,N_2200);
nand U5428 (N_5428,N_2443,N_240);
nand U5429 (N_5429,N_1742,N_4279);
or U5430 (N_5430,N_4496,N_3547);
nor U5431 (N_5431,N_1472,N_819);
or U5432 (N_5432,N_139,N_210);
or U5433 (N_5433,N_3334,N_2927);
nand U5434 (N_5434,N_2984,N_507);
nand U5435 (N_5435,N_3672,N_1253);
and U5436 (N_5436,N_3532,N_3807);
nor U5437 (N_5437,N_1123,N_967);
or U5438 (N_5438,N_3090,N_327);
xor U5439 (N_5439,N_2585,N_3436);
and U5440 (N_5440,N_2360,N_4179);
xnor U5441 (N_5441,N_4283,N_250);
nand U5442 (N_5442,N_4633,N_1499);
and U5443 (N_5443,N_2717,N_2971);
nand U5444 (N_5444,N_1489,N_4097);
and U5445 (N_5445,N_4910,N_1089);
or U5446 (N_5446,N_1696,N_3050);
and U5447 (N_5447,N_3513,N_2844);
nand U5448 (N_5448,N_3301,N_85);
nand U5449 (N_5449,N_1222,N_3683);
nand U5450 (N_5450,N_2224,N_4886);
and U5451 (N_5451,N_1042,N_3905);
or U5452 (N_5452,N_4419,N_3274);
xor U5453 (N_5453,N_2404,N_3719);
xor U5454 (N_5454,N_4296,N_4357);
nor U5455 (N_5455,N_342,N_3043);
or U5456 (N_5456,N_614,N_3951);
or U5457 (N_5457,N_1719,N_1982);
and U5458 (N_5458,N_2765,N_4571);
and U5459 (N_5459,N_2263,N_3589);
or U5460 (N_5460,N_4710,N_2796);
xnor U5461 (N_5461,N_4054,N_15);
xnor U5462 (N_5462,N_3716,N_3965);
nor U5463 (N_5463,N_4776,N_1324);
xor U5464 (N_5464,N_1137,N_168);
nor U5465 (N_5465,N_4922,N_3828);
nor U5466 (N_5466,N_1148,N_293);
and U5467 (N_5467,N_691,N_2311);
xnor U5468 (N_5468,N_4935,N_477);
and U5469 (N_5469,N_3453,N_3460);
and U5470 (N_5470,N_145,N_3454);
and U5471 (N_5471,N_880,N_2338);
nor U5472 (N_5472,N_916,N_3218);
or U5473 (N_5473,N_1192,N_3642);
nand U5474 (N_5474,N_3307,N_1271);
nor U5475 (N_5475,N_4584,N_1344);
nand U5476 (N_5476,N_2213,N_3841);
nand U5477 (N_5477,N_1728,N_2476);
and U5478 (N_5478,N_3648,N_2069);
xor U5479 (N_5479,N_605,N_463);
or U5480 (N_5480,N_1948,N_3465);
or U5481 (N_5481,N_3625,N_1183);
xor U5482 (N_5482,N_225,N_752);
nand U5483 (N_5483,N_1082,N_4402);
xnor U5484 (N_5484,N_4721,N_2307);
nor U5485 (N_5485,N_2944,N_2579);
or U5486 (N_5486,N_3922,N_3963);
nor U5487 (N_5487,N_1817,N_2671);
and U5488 (N_5488,N_494,N_255);
and U5489 (N_5489,N_3076,N_4329);
xnor U5490 (N_5490,N_4405,N_3382);
and U5491 (N_5491,N_349,N_1535);
nand U5492 (N_5492,N_524,N_2875);
xnor U5493 (N_5493,N_4749,N_1970);
and U5494 (N_5494,N_711,N_1760);
or U5495 (N_5495,N_2332,N_2504);
nor U5496 (N_5496,N_90,N_4145);
xnor U5497 (N_5497,N_2821,N_333);
nor U5498 (N_5498,N_773,N_4530);
nor U5499 (N_5499,N_4866,N_3864);
nand U5500 (N_5500,N_1449,N_4064);
nor U5501 (N_5501,N_3299,N_4653);
nor U5502 (N_5502,N_3126,N_1286);
or U5503 (N_5503,N_2656,N_806);
and U5504 (N_5504,N_964,N_3722);
xor U5505 (N_5505,N_4004,N_1425);
nor U5506 (N_5506,N_27,N_527);
nand U5507 (N_5507,N_3185,N_3485);
nand U5508 (N_5508,N_2530,N_3944);
nand U5509 (N_5509,N_4686,N_4804);
xor U5510 (N_5510,N_4083,N_2562);
xnor U5511 (N_5511,N_650,N_4177);
nand U5512 (N_5512,N_4209,N_4273);
and U5513 (N_5513,N_2635,N_842);
nand U5514 (N_5514,N_4173,N_2177);
or U5515 (N_5515,N_1260,N_1830);
and U5516 (N_5516,N_2122,N_2352);
or U5517 (N_5517,N_798,N_2031);
and U5518 (N_5518,N_2365,N_4555);
and U5519 (N_5519,N_3383,N_4781);
xor U5520 (N_5520,N_1630,N_4110);
and U5521 (N_5521,N_3283,N_2791);
xor U5522 (N_5522,N_3790,N_4475);
nor U5523 (N_5523,N_4065,N_2369);
nor U5524 (N_5524,N_186,N_593);
nand U5525 (N_5525,N_4487,N_3163);
nor U5526 (N_5526,N_3461,N_1835);
nand U5527 (N_5527,N_586,N_4184);
xnor U5528 (N_5528,N_4989,N_1530);
nor U5529 (N_5529,N_4192,N_1247);
nor U5530 (N_5530,N_796,N_3763);
nor U5531 (N_5531,N_2083,N_2347);
nand U5532 (N_5532,N_2747,N_4733);
and U5533 (N_5533,N_815,N_3688);
and U5534 (N_5534,N_30,N_3936);
nor U5535 (N_5535,N_2977,N_4266);
nor U5536 (N_5536,N_3843,N_4455);
or U5537 (N_5537,N_979,N_1311);
nand U5538 (N_5538,N_42,N_3491);
or U5539 (N_5539,N_220,N_4889);
nor U5540 (N_5540,N_4016,N_177);
and U5541 (N_5541,N_649,N_1453);
and U5542 (N_5542,N_3137,N_4836);
nand U5543 (N_5543,N_4871,N_2523);
and U5544 (N_5544,N_2150,N_2008);
nand U5545 (N_5545,N_3724,N_1051);
and U5546 (N_5546,N_4849,N_453);
nor U5547 (N_5547,N_1967,N_3063);
nand U5548 (N_5548,N_686,N_2521);
and U5549 (N_5549,N_1231,N_1350);
nor U5550 (N_5550,N_1687,N_2188);
or U5551 (N_5551,N_3265,N_1520);
and U5552 (N_5552,N_363,N_1094);
and U5553 (N_5553,N_1522,N_3565);
nor U5554 (N_5554,N_128,N_412);
or U5555 (N_5555,N_2558,N_900);
and U5556 (N_5556,N_2607,N_1091);
or U5557 (N_5557,N_467,N_557);
nor U5558 (N_5558,N_4702,N_2556);
nor U5559 (N_5559,N_3640,N_2687);
nor U5560 (N_5560,N_4193,N_1023);
or U5561 (N_5561,N_3469,N_2099);
nor U5562 (N_5562,N_1751,N_939);
or U5563 (N_5563,N_373,N_905);
nor U5564 (N_5564,N_2056,N_2220);
nand U5565 (N_5565,N_1571,N_3873);
or U5566 (N_5566,N_2022,N_4391);
nand U5567 (N_5567,N_3634,N_4149);
or U5568 (N_5568,N_4518,N_1641);
nor U5569 (N_5569,N_3438,N_339);
nor U5570 (N_5570,N_1504,N_2234);
and U5571 (N_5571,N_1905,N_2243);
and U5572 (N_5572,N_2367,N_1754);
or U5573 (N_5573,N_4247,N_3578);
nor U5574 (N_5574,N_286,N_1470);
nor U5575 (N_5575,N_604,N_3819);
nor U5576 (N_5576,N_692,N_888);
nor U5577 (N_5577,N_3563,N_4474);
or U5578 (N_5578,N_4844,N_9);
nor U5579 (N_5579,N_2938,N_2662);
nand U5580 (N_5580,N_1953,N_1758);
nor U5581 (N_5581,N_1842,N_1738);
and U5582 (N_5582,N_3152,N_4375);
nand U5583 (N_5583,N_4590,N_3190);
nor U5584 (N_5584,N_1115,N_4006);
or U5585 (N_5585,N_61,N_1049);
or U5586 (N_5586,N_466,N_2553);
xor U5587 (N_5587,N_2510,N_4517);
nor U5588 (N_5588,N_4586,N_2632);
nand U5589 (N_5589,N_716,N_1182);
nand U5590 (N_5590,N_2843,N_4544);
nand U5591 (N_5591,N_947,N_4551);
xor U5592 (N_5592,N_2820,N_132);
nand U5593 (N_5593,N_3343,N_4680);
or U5594 (N_5594,N_2098,N_1203);
or U5595 (N_5595,N_4239,N_4433);
nor U5596 (N_5596,N_2690,N_4541);
nor U5597 (N_5597,N_4742,N_1887);
and U5598 (N_5598,N_2337,N_4161);
and U5599 (N_5599,N_2385,N_4508);
nor U5600 (N_5600,N_4582,N_2381);
nand U5601 (N_5601,N_577,N_695);
or U5602 (N_5602,N_2663,N_2403);
or U5603 (N_5603,N_2516,N_4365);
nand U5604 (N_5604,N_3893,N_275);
nand U5605 (N_5605,N_3879,N_491);
nand U5606 (N_5606,N_2304,N_1444);
and U5607 (N_5607,N_3425,N_4241);
nor U5608 (N_5608,N_160,N_2631);
and U5609 (N_5609,N_98,N_1011);
or U5610 (N_5610,N_2329,N_765);
or U5611 (N_5611,N_1456,N_3527);
nor U5612 (N_5612,N_1230,N_3001);
or U5613 (N_5613,N_2867,N_94);
nor U5614 (N_5614,N_1570,N_3756);
xor U5615 (N_5615,N_674,N_4464);
or U5616 (N_5616,N_1197,N_1787);
xnor U5617 (N_5617,N_3741,N_147);
or U5618 (N_5618,N_4821,N_4924);
xnor U5619 (N_5619,N_4482,N_663);
nand U5620 (N_5620,N_3407,N_3930);
nor U5621 (N_5621,N_3848,N_1805);
nand U5622 (N_5622,N_4416,N_1105);
or U5623 (N_5623,N_449,N_209);
or U5624 (N_5624,N_3275,N_4734);
nand U5625 (N_5625,N_1207,N_3577);
nand U5626 (N_5626,N_400,N_4059);
nor U5627 (N_5627,N_1838,N_3813);
nor U5628 (N_5628,N_4511,N_2439);
or U5629 (N_5629,N_3129,N_4578);
nor U5630 (N_5630,N_630,N_2968);
nand U5631 (N_5631,N_1019,N_1259);
and U5632 (N_5632,N_3654,N_1797);
or U5633 (N_5633,N_392,N_481);
nor U5634 (N_5634,N_2908,N_3112);
and U5635 (N_5635,N_1121,N_4472);
and U5636 (N_5636,N_3069,N_573);
and U5637 (N_5637,N_3202,N_2895);
or U5638 (N_5638,N_615,N_4501);
nand U5639 (N_5639,N_744,N_4438);
or U5640 (N_5640,N_2173,N_2725);
nor U5641 (N_5641,N_3575,N_3151);
or U5642 (N_5642,N_2705,N_1341);
xnor U5643 (N_5643,N_1158,N_86);
nor U5644 (N_5644,N_718,N_2306);
nor U5645 (N_5645,N_2371,N_3413);
nor U5646 (N_5646,N_1501,N_2998);
and U5647 (N_5647,N_1077,N_4450);
nor U5648 (N_5648,N_2144,N_4291);
nand U5649 (N_5649,N_2258,N_4454);
xnor U5650 (N_5650,N_2216,N_1753);
or U5651 (N_5651,N_2105,N_3523);
or U5652 (N_5652,N_3837,N_3793);
and U5653 (N_5653,N_1027,N_3361);
xnor U5654 (N_5654,N_1708,N_3212);
xnor U5655 (N_5655,N_2159,N_4426);
or U5656 (N_5656,N_814,N_1443);
nor U5657 (N_5657,N_2740,N_852);
and U5658 (N_5658,N_2330,N_1926);
nand U5659 (N_5659,N_1512,N_178);
and U5660 (N_5660,N_1933,N_641);
and U5661 (N_5661,N_3635,N_3795);
nor U5662 (N_5662,N_4235,N_2376);
or U5663 (N_5663,N_4168,N_4047);
nand U5664 (N_5664,N_324,N_4313);
xor U5665 (N_5665,N_4587,N_3079);
and U5666 (N_5666,N_4996,N_627);
and U5667 (N_5667,N_2864,N_3329);
nor U5668 (N_5668,N_1828,N_3690);
and U5669 (N_5669,N_4834,N_1822);
xor U5670 (N_5670,N_3020,N_1806);
and U5671 (N_5671,N_4768,N_3300);
nand U5672 (N_5672,N_2084,N_3714);
and U5673 (N_5673,N_4351,N_1433);
xor U5674 (N_5674,N_846,N_3731);
and U5675 (N_5675,N_4275,N_501);
nor U5676 (N_5676,N_697,N_665);
xor U5677 (N_5677,N_2465,N_3811);
nor U5678 (N_5678,N_3015,N_810);
or U5679 (N_5679,N_438,N_278);
or U5680 (N_5680,N_480,N_1138);
or U5681 (N_5681,N_3032,N_108);
and U5682 (N_5682,N_2918,N_281);
nand U5683 (N_5683,N_2815,N_1007);
nand U5684 (N_5684,N_857,N_4466);
xor U5685 (N_5685,N_4032,N_2532);
nand U5686 (N_5686,N_2283,N_3806);
xnor U5687 (N_5687,N_2117,N_782);
nor U5688 (N_5688,N_73,N_862);
nor U5689 (N_5689,N_3696,N_873);
nor U5690 (N_5690,N_3805,N_2282);
nor U5691 (N_5691,N_2468,N_4088);
nor U5692 (N_5692,N_4504,N_2722);
or U5693 (N_5693,N_3949,N_3912);
nor U5694 (N_5694,N_1895,N_726);
or U5695 (N_5695,N_770,N_3124);
or U5696 (N_5696,N_4890,N_1037);
and U5697 (N_5697,N_551,N_3371);
nor U5698 (N_5698,N_1612,N_4285);
nor U5699 (N_5699,N_2987,N_1316);
nand U5700 (N_5700,N_2463,N_2341);
and U5701 (N_5701,N_2169,N_69);
xor U5702 (N_5702,N_749,N_3104);
and U5703 (N_5703,N_3620,N_3670);
nand U5704 (N_5704,N_2455,N_3854);
nand U5705 (N_5705,N_6,N_3346);
and U5706 (N_5706,N_2763,N_3832);
nand U5707 (N_5707,N_3660,N_1634);
xnor U5708 (N_5708,N_2742,N_4011);
xnor U5709 (N_5709,N_3327,N_2097);
nor U5710 (N_5710,N_2076,N_4593);
nor U5711 (N_5711,N_3277,N_2620);
nand U5712 (N_5712,N_3099,N_2163);
nand U5713 (N_5713,N_3858,N_3443);
nor U5714 (N_5714,N_1583,N_4852);
nand U5715 (N_5715,N_2005,N_2484);
or U5716 (N_5716,N_625,N_4753);
nor U5717 (N_5717,N_1788,N_1557);
nand U5718 (N_5718,N_758,N_4997);
xor U5719 (N_5719,N_4178,N_3594);
nor U5720 (N_5720,N_1217,N_425);
xor U5721 (N_5721,N_423,N_3221);
nor U5722 (N_5722,N_1210,N_1682);
or U5723 (N_5723,N_4547,N_3966);
xnor U5724 (N_5724,N_2694,N_235);
nand U5725 (N_5725,N_2559,N_944);
or U5726 (N_5726,N_1135,N_111);
or U5727 (N_5727,N_4623,N_1283);
nand U5728 (N_5728,N_2651,N_4793);
nand U5729 (N_5729,N_1195,N_732);
nor U5730 (N_5730,N_2888,N_1650);
xnor U5731 (N_5731,N_1479,N_1517);
nor U5732 (N_5732,N_4791,N_4515);
nor U5733 (N_5733,N_1725,N_4159);
or U5734 (N_5734,N_1031,N_546);
and U5735 (N_5735,N_343,N_959);
nand U5736 (N_5736,N_4939,N_1694);
nor U5737 (N_5737,N_2233,N_555);
nand U5738 (N_5738,N_4228,N_4817);
nor U5739 (N_5739,N_4344,N_3586);
nand U5740 (N_5740,N_1168,N_385);
or U5741 (N_5741,N_3052,N_4715);
nor U5742 (N_5742,N_2970,N_124);
and U5743 (N_5743,N_2091,N_1690);
nand U5744 (N_5744,N_3482,N_4325);
or U5745 (N_5745,N_154,N_3226);
or U5746 (N_5746,N_2911,N_2866);
nand U5747 (N_5747,N_4657,N_3375);
and U5748 (N_5748,N_2669,N_737);
or U5749 (N_5749,N_4302,N_2697);
xnor U5750 (N_5750,N_2081,N_151);
or U5751 (N_5751,N_1411,N_3549);
nand U5752 (N_5752,N_3847,N_1068);
and U5753 (N_5753,N_4810,N_4792);
nand U5754 (N_5754,N_2225,N_1666);
and U5755 (N_5755,N_3059,N_4023);
nand U5756 (N_5756,N_4139,N_1882);
nand U5757 (N_5757,N_3096,N_1543);
or U5758 (N_5758,N_882,N_712);
and U5759 (N_5759,N_1322,N_2850);
nor U5760 (N_5760,N_2130,N_4865);
nor U5761 (N_5761,N_713,N_1837);
and U5762 (N_5762,N_4549,N_492);
nand U5763 (N_5763,N_4570,N_2300);
nor U5764 (N_5764,N_2103,N_1766);
nor U5765 (N_5765,N_2492,N_4323);
or U5766 (N_5766,N_974,N_766);
xnor U5767 (N_5767,N_4968,N_1441);
nand U5768 (N_5768,N_2308,N_3336);
nor U5769 (N_5769,N_3414,N_637);
or U5770 (N_5770,N_2007,N_454);
nand U5771 (N_5771,N_2881,N_850);
or U5772 (N_5772,N_2778,N_223);
or U5773 (N_5773,N_3177,N_3684);
nand U5774 (N_5774,N_3424,N_3996);
nor U5775 (N_5775,N_2101,N_169);
nor U5776 (N_5776,N_868,N_2514);
nand U5777 (N_5777,N_2239,N_2146);
nand U5778 (N_5778,N_1095,N_3140);
nand U5779 (N_5779,N_3528,N_1067);
or U5780 (N_5780,N_3198,N_4164);
or U5781 (N_5781,N_925,N_1057);
nor U5782 (N_5782,N_4305,N_3985);
xor U5783 (N_5783,N_4435,N_2197);
or U5784 (N_5784,N_3860,N_1861);
xnor U5785 (N_5785,N_759,N_106);
and U5786 (N_5786,N_3899,N_4526);
nand U5787 (N_5787,N_1977,N_1747);
nand U5788 (N_5788,N_3956,N_406);
nor U5789 (N_5789,N_540,N_1268);
and U5790 (N_5790,N_1525,N_545);
nor U5791 (N_5791,N_4031,N_4341);
and U5792 (N_5792,N_2520,N_3446);
nand U5793 (N_5793,N_763,N_2757);
nand U5794 (N_5794,N_1406,N_3787);
nand U5795 (N_5795,N_2916,N_4589);
xor U5796 (N_5796,N_1695,N_2889);
nor U5797 (N_5797,N_455,N_1963);
nor U5798 (N_5798,N_3010,N_1773);
or U5799 (N_5799,N_764,N_975);
nor U5800 (N_5800,N_535,N_2780);
xor U5801 (N_5801,N_4401,N_3869);
nand U5802 (N_5802,N_329,N_923);
xnor U5803 (N_5803,N_1190,N_2151);
and U5804 (N_5804,N_4929,N_834);
nand U5805 (N_5805,N_413,N_3047);
or U5806 (N_5806,N_2018,N_4101);
and U5807 (N_5807,N_2548,N_1541);
nor U5808 (N_5808,N_451,N_4966);
nand U5809 (N_5809,N_341,N_133);
or U5810 (N_5810,N_4267,N_3353);
or U5811 (N_5811,N_2350,N_353);
xor U5812 (N_5812,N_1361,N_4319);
nor U5813 (N_5813,N_2270,N_4115);
and U5814 (N_5814,N_2846,N_2702);
or U5815 (N_5815,N_1333,N_4660);
nand U5816 (N_5816,N_1971,N_59);
nor U5817 (N_5817,N_3468,N_561);
or U5818 (N_5818,N_3768,N_4944);
nor U5819 (N_5819,N_2575,N_563);
nor U5820 (N_5820,N_4265,N_1640);
and U5821 (N_5821,N_424,N_522);
nand U5822 (N_5822,N_906,N_4775);
and U5823 (N_5823,N_3601,N_2132);
or U5824 (N_5824,N_4034,N_4624);
and U5825 (N_5825,N_4163,N_3410);
or U5826 (N_5826,N_4893,N_1978);
nand U5827 (N_5827,N_14,N_497);
nor U5828 (N_5828,N_2807,N_4920);
nand U5829 (N_5829,N_2727,N_1794);
nand U5830 (N_5830,N_505,N_3913);
and U5831 (N_5831,N_0,N_1597);
or U5832 (N_5832,N_2485,N_1784);
and U5833 (N_5833,N_3168,N_2810);
xor U5834 (N_5834,N_1746,N_1460);
and U5835 (N_5835,N_1140,N_658);
xnor U5836 (N_5836,N_1915,N_4882);
and U5837 (N_5837,N_1241,N_4213);
nand U5838 (N_5838,N_1874,N_262);
nor U5839 (N_5839,N_2828,N_3216);
nor U5840 (N_5840,N_4194,N_3984);
or U5841 (N_5841,N_1997,N_3574);
nor U5842 (N_5842,N_2195,N_1744);
or U5843 (N_5843,N_3025,N_4317);
and U5844 (N_5844,N_2223,N_968);
nor U5845 (N_5845,N_2764,N_793);
nor U5846 (N_5846,N_902,N_1006);
xor U5847 (N_5847,N_2327,N_3610);
or U5848 (N_5848,N_377,N_1999);
nand U5849 (N_5849,N_3863,N_16);
xor U5850 (N_5850,N_1586,N_3800);
and U5851 (N_5851,N_4133,N_550);
xnor U5852 (N_5852,N_890,N_1440);
or U5853 (N_5853,N_4662,N_3861);
and U5854 (N_5854,N_2539,N_4730);
nor U5855 (N_5855,N_2568,N_3006);
xor U5856 (N_5856,N_1493,N_2030);
or U5857 (N_5857,N_2914,N_3098);
or U5858 (N_5858,N_4801,N_4819);
nor U5859 (N_5859,N_4888,N_3652);
nor U5860 (N_5860,N_1056,N_3992);
nand U5861 (N_5861,N_949,N_4225);
and U5862 (N_5862,N_3330,N_4729);
and U5863 (N_5863,N_2191,N_4001);
and U5864 (N_5864,N_4436,N_1114);
or U5865 (N_5865,N_2374,N_562);
and U5866 (N_5866,N_4152,N_4490);
and U5867 (N_5867,N_4627,N_4649);
xor U5868 (N_5868,N_93,N_394);
nor U5869 (N_5869,N_2941,N_149);
and U5870 (N_5870,N_4451,N_2869);
and U5871 (N_5871,N_1639,N_2060);
nand U5872 (N_5872,N_1017,N_2565);
or U5873 (N_5873,N_1079,N_1090);
and U5874 (N_5874,N_3954,N_4465);
or U5875 (N_5875,N_239,N_3953);
xor U5876 (N_5876,N_1250,N_446);
or U5877 (N_5877,N_1607,N_1886);
nor U5878 (N_5878,N_3538,N_4066);
nand U5879 (N_5879,N_3048,N_3705);
nand U5880 (N_5880,N_1515,N_3142);
nand U5881 (N_5881,N_3896,N_3938);
or U5882 (N_5882,N_4728,N_4506);
nand U5883 (N_5883,N_4332,N_3445);
nand U5884 (N_5884,N_3480,N_3359);
nor U5885 (N_5885,N_4967,N_2873);
or U5886 (N_5886,N_3988,N_4682);
xor U5887 (N_5887,N_3254,N_4704);
nor U5888 (N_5888,N_3779,N_3744);
or U5889 (N_5889,N_4675,N_4833);
or U5890 (N_5890,N_2816,N_4461);
nand U5891 (N_5891,N_689,N_1938);
nor U5892 (N_5892,N_1353,N_2092);
nand U5893 (N_5893,N_2469,N_2281);
nand U5894 (N_5894,N_4940,N_946);
nor U5895 (N_5895,N_2275,N_4655);
nor U5896 (N_5896,N_2710,N_3766);
and U5897 (N_5897,N_731,N_668);
xor U5898 (N_5898,N_2124,N_2919);
nor U5899 (N_5899,N_309,N_1802);
and U5900 (N_5900,N_4645,N_3397);
nor U5901 (N_5901,N_675,N_4984);
nand U5902 (N_5902,N_3733,N_1950);
or U5903 (N_5903,N_4647,N_1315);
nor U5904 (N_5904,N_1972,N_1556);
nor U5905 (N_5905,N_3364,N_2161);
and U5906 (N_5906,N_1262,N_358);
or U5907 (N_5907,N_2057,N_3797);
nor U5908 (N_5908,N_439,N_137);
nand U5909 (N_5909,N_559,N_36);
or U5910 (N_5910,N_3590,N_3761);
nor U5911 (N_5911,N_3752,N_131);
nand U5912 (N_5912,N_1629,N_4476);
xor U5913 (N_5913,N_2133,N_3219);
xor U5914 (N_5914,N_2079,N_3278);
nor U5915 (N_5915,N_4278,N_3786);
nand U5916 (N_5916,N_3318,N_196);
nand U5917 (N_5917,N_426,N_432);
nand U5918 (N_5918,N_1942,N_1947);
and U5919 (N_5919,N_3835,N_3304);
or U5920 (N_5920,N_2529,N_669);
nand U5921 (N_5921,N_140,N_2434);
and U5922 (N_5922,N_3027,N_3253);
or U5923 (N_5923,N_1269,N_4183);
xnor U5924 (N_5924,N_3677,N_3037);
nor U5925 (N_5925,N_2343,N_3758);
nor U5926 (N_5926,N_311,N_2561);
nand U5927 (N_5927,N_71,N_441);
nor U5928 (N_5928,N_1866,N_511);
xnor U5929 (N_5929,N_2135,N_2287);
or U5930 (N_5930,N_1145,N_3100);
nor U5931 (N_5931,N_3292,N_2201);
nor U5932 (N_5932,N_4820,N_3845);
or U5933 (N_5933,N_3172,N_3701);
and U5934 (N_5934,N_2715,N_3246);
and U5935 (N_5935,N_619,N_1066);
nand U5936 (N_5936,N_3117,N_3297);
nor U5937 (N_5937,N_2073,N_2909);
and U5938 (N_5938,N_2372,N_1854);
and U5939 (N_5939,N_2589,N_523);
nand U5940 (N_5940,N_2291,N_570);
and U5941 (N_5941,N_1328,N_2612);
nor U5942 (N_5942,N_2664,N_2811);
nand U5943 (N_5943,N_702,N_3391);
xnor U5944 (N_5944,N_833,N_4854);
nand U5945 (N_5945,N_3687,N_1676);
nor U5946 (N_5946,N_376,N_1108);
and U5947 (N_5947,N_3497,N_3704);
nand U5948 (N_5948,N_1782,N_4007);
nor U5949 (N_5949,N_807,N_396);
and U5950 (N_5950,N_1136,N_4671);
xnor U5951 (N_5951,N_2661,N_790);
nor U5952 (N_5952,N_264,N_39);
nand U5953 (N_5953,N_2112,N_192);
or U5954 (N_5954,N_2689,N_2900);
and U5955 (N_5955,N_3999,N_1871);
xor U5956 (N_5956,N_3957,N_126);
nor U5957 (N_5957,N_1212,N_269);
nand U5958 (N_5958,N_2872,N_1482);
nand U5959 (N_5959,N_493,N_628);
nand U5960 (N_5960,N_386,N_4018);
or U5961 (N_5961,N_622,N_3478);
and U5962 (N_5962,N_980,N_4546);
nand U5963 (N_5963,N_134,N_437);
nand U5964 (N_5964,N_1858,N_1110);
and U5965 (N_5965,N_2685,N_1400);
nand U5966 (N_5966,N_4155,N_4650);
nand U5967 (N_5967,N_2334,N_469);
xnor U5968 (N_5968,N_1777,N_2942);
nor U5969 (N_5969,N_2006,N_2719);
or U5970 (N_5970,N_590,N_4411);
and U5971 (N_5971,N_1164,N_784);
nand U5972 (N_5972,N_4553,N_3249);
and U5973 (N_5973,N_1863,N_2410);
nor U5974 (N_5974,N_122,N_4885);
or U5975 (N_5975,N_2886,N_4370);
nand U5976 (N_5976,N_2106,N_4789);
xnor U5977 (N_5977,N_1968,N_3599);
nor U5978 (N_5978,N_2261,N_4014);
and U5979 (N_5979,N_2963,N_1913);
xnor U5980 (N_5980,N_767,N_3352);
and U5981 (N_5981,N_2517,N_1326);
nor U5982 (N_5982,N_299,N_3258);
or U5983 (N_5983,N_2974,N_245);
and U5984 (N_5984,N_1734,N_3814);
or U5985 (N_5985,N_3507,N_4898);
nand U5986 (N_5986,N_3068,N_1459);
and U5987 (N_5987,N_4692,N_2405);
nor U5988 (N_5988,N_2524,N_4290);
and U5989 (N_5989,N_2540,N_2214);
nand U5990 (N_5990,N_1623,N_290);
nor U5991 (N_5991,N_1131,N_4959);
and U5992 (N_5992,N_4400,N_2986);
nor U5993 (N_5993,N_1906,N_2254);
nand U5994 (N_5994,N_2979,N_1010);
or U5995 (N_5995,N_1503,N_4223);
and U5996 (N_5996,N_1327,N_3321);
nand U5997 (N_5997,N_4182,N_1551);
and U5998 (N_5998,N_3816,N_2903);
or U5999 (N_5999,N_3498,N_1134);
nor U6000 (N_6000,N_929,N_4005);
xor U6001 (N_6001,N_4056,N_1756);
and U6002 (N_6002,N_2536,N_3284);
and U6003 (N_6003,N_3656,N_4701);
nand U6004 (N_6004,N_2991,N_927);
nand U6005 (N_6005,N_3072,N_4025);
or U6006 (N_6006,N_3481,N_328);
and U6007 (N_6007,N_881,N_4078);
or U6008 (N_6008,N_2755,N_1718);
or U6009 (N_6009,N_2609,N_633);
xnor U6010 (N_6010,N_2491,N_1447);
nor U6011 (N_6011,N_1803,N_261);
or U6012 (N_6012,N_1163,N_4377);
nor U6013 (N_6013,N_3114,N_3711);
and U6014 (N_6014,N_4394,N_416);
and U6015 (N_6015,N_184,N_4507);
nor U6016 (N_6016,N_3542,N_462);
nor U6017 (N_6017,N_3183,N_3627);
nor U6018 (N_6018,N_484,N_3123);
nor U6019 (N_6019,N_3753,N_1143);
or U6020 (N_6020,N_2847,N_1401);
and U6021 (N_6021,N_3456,N_2905);
nand U6022 (N_6022,N_3659,N_2720);
and U6023 (N_6023,N_2420,N_1939);
or U6024 (N_6024,N_4895,N_1127);
nand U6025 (N_6025,N_926,N_715);
or U6026 (N_6026,N_2289,N_3462);
and U6027 (N_6027,N_2893,N_1860);
nor U6028 (N_6028,N_1093,N_3092);
or U6029 (N_6029,N_3600,N_3189);
and U6030 (N_6030,N_729,N_988);
and U6031 (N_6031,N_450,N_1211);
nand U6032 (N_6032,N_3471,N_3773);
nor U6033 (N_6033,N_4479,N_3526);
or U6034 (N_6034,N_2259,N_1295);
and U6035 (N_6035,N_4386,N_2110);
nor U6036 (N_6036,N_51,N_774);
and U6037 (N_6037,N_1434,N_4175);
nand U6038 (N_6038,N_1919,N_1927);
or U6039 (N_6039,N_1386,N_3676);
nor U6040 (N_6040,N_2863,N_1277);
and U6041 (N_6041,N_1772,N_3735);
nor U6042 (N_6042,N_3145,N_1436);
xnor U6043 (N_6043,N_4765,N_3643);
or U6044 (N_6044,N_4574,N_3505);
or U6045 (N_6045,N_1198,N_4353);
nor U6046 (N_6046,N_2497,N_1494);
and U6047 (N_6047,N_1840,N_296);
or U6048 (N_6048,N_4270,N_4608);
and U6049 (N_6049,N_3941,N_2321);
nor U6050 (N_6050,N_3362,N_3344);
xnor U6051 (N_6051,N_277,N_3900);
nand U6052 (N_6052,N_1879,N_409);
nor U6053 (N_6053,N_2512,N_289);
and U6054 (N_6054,N_3736,N_3368);
nand U6055 (N_6055,N_2743,N_4554);
nand U6056 (N_6056,N_442,N_123);
nand U6057 (N_6057,N_2940,N_2351);
or U6058 (N_6058,N_1375,N_1452);
nor U6059 (N_6059,N_2245,N_786);
or U6060 (N_6060,N_4174,N_1480);
nor U6061 (N_6061,N_4685,N_3281);
or U6062 (N_6062,N_2897,N_2344);
or U6063 (N_6063,N_1636,N_2424);
and U6064 (N_6064,N_4695,N_2406);
nor U6065 (N_6065,N_4735,N_2708);
nor U6066 (N_6066,N_4413,N_3639);
or U6067 (N_6067,N_3089,N_2379);
xnor U6068 (N_6068,N_1585,N_4815);
nand U6069 (N_6069,N_3338,N_4548);
or U6070 (N_6070,N_68,N_2446);
and U6071 (N_6071,N_2983,N_1867);
nand U6072 (N_6072,N_4802,N_2244);
or U6073 (N_6073,N_161,N_2096);
nor U6074 (N_6074,N_2126,N_4575);
nand U6075 (N_6075,N_2488,N_1404);
nor U6076 (N_6076,N_4468,N_3862);
or U6077 (N_6077,N_1661,N_3633);
and U6078 (N_6078,N_3280,N_2733);
or U6079 (N_6079,N_4495,N_3486);
nor U6080 (N_6080,N_738,N_3754);
and U6081 (N_6081,N_2142,N_4033);
or U6082 (N_6082,N_1317,N_1985);
and U6083 (N_6083,N_987,N_4719);
xor U6084 (N_6084,N_2602,N_4607);
and U6085 (N_6085,N_4467,N_1179);
nor U6086 (N_6086,N_4894,N_4513);
nor U6087 (N_6087,N_2152,N_4044);
or U6088 (N_6088,N_2428,N_3337);
xnor U6089 (N_6089,N_908,N_4316);
nor U6090 (N_6090,N_4943,N_4648);
and U6091 (N_6091,N_4389,N_3788);
and U6092 (N_6092,N_1807,N_3313);
nand U6093 (N_6093,N_2912,N_403);
or U6094 (N_6094,N_2211,N_3728);
or U6095 (N_6095,N_1881,N_1958);
nor U6096 (N_6096,N_1799,N_4509);
and U6097 (N_6097,N_3508,N_746);
or U6098 (N_6098,N_1679,N_680);
nor U6099 (N_6099,N_2851,N_2147);
xor U6100 (N_6100,N_4268,N_4600);
or U6101 (N_6101,N_3693,N_1491);
xor U6102 (N_6102,N_2528,N_38);
or U6103 (N_6103,N_3282,N_1865);
and U6104 (N_6104,N_2250,N_2573);
nor U6105 (N_6105,N_4739,N_63);
and U6106 (N_6106,N_548,N_1847);
and U6107 (N_6107,N_4140,N_2422);
or U6108 (N_6108,N_943,N_1155);
nand U6109 (N_6109,N_568,N_282);
nand U6110 (N_6110,N_2174,N_3950);
and U6111 (N_6111,N_4958,N_4790);
and U6112 (N_6112,N_2973,N_2618);
nor U6113 (N_6113,N_750,N_4457);
and U6114 (N_6114,N_2472,N_2442);
and U6115 (N_6115,N_476,N_4846);
or U6116 (N_6116,N_3101,N_3882);
nor U6117 (N_6117,N_2511,N_2738);
nand U6118 (N_6118,N_4498,N_2613);
or U6119 (N_6119,N_4380,N_2158);
xnor U6120 (N_6120,N_4237,N_1273);
and U6121 (N_6121,N_1750,N_241);
and U6122 (N_6122,N_4460,N_725);
xor U6123 (N_6123,N_4206,N_4722);
or U6124 (N_6124,N_757,N_4315);
and U6125 (N_6125,N_4215,N_2746);
and U6126 (N_6126,N_1599,N_4469);
nor U6127 (N_6127,N_3983,N_113);
xor U6128 (N_6128,N_4543,N_83);
nand U6129 (N_6129,N_1649,N_3057);
and U6130 (N_6130,N_1710,N_2215);
nand U6131 (N_6131,N_1028,N_2614);
nor U6132 (N_6132,N_2936,N_4750);
nand U6133 (N_6133,N_1129,N_2950);
or U6134 (N_6134,N_4113,N_4484);
or U6135 (N_6135,N_3942,N_4067);
nand U6136 (N_6136,N_4200,N_2426);
nand U6137 (N_6137,N_748,N_3877);
or U6138 (N_6138,N_1726,N_2155);
xnor U6139 (N_6139,N_4099,N_4392);
and U6140 (N_6140,N_4308,N_4982);
or U6141 (N_6141,N_2676,N_4759);
and U6142 (N_6142,N_3972,N_445);
nand U6143 (N_6143,N_2292,N_2430);
xnor U6144 (N_6144,N_2932,N_1254);
or U6145 (N_6145,N_4383,N_1531);
xor U6146 (N_6146,N_4009,N_334);
or U6147 (N_6147,N_1767,N_4320);
xor U6148 (N_6148,N_1990,N_4599);
xnor U6149 (N_6149,N_1576,N_4942);
or U6150 (N_6150,N_3702,N_1996);
xor U6151 (N_6151,N_4236,N_845);
nand U6152 (N_6152,N_696,N_1098);
nor U6153 (N_6153,N_331,N_1800);
nor U6154 (N_6154,N_2805,N_389);
nand U6155 (N_6155,N_2992,N_3242);
and U6156 (N_6156,N_1355,N_4378);
nor U6157 (N_6157,N_4628,N_1366);
and U6158 (N_6158,N_244,N_3180);
and U6159 (N_6159,N_204,N_661);
xor U6160 (N_6160,N_2028,N_1186);
or U6161 (N_6161,N_4057,N_3159);
and U6162 (N_6162,N_3395,N_1060);
and U6163 (N_6163,N_3007,N_1457);
nand U6164 (N_6164,N_3555,N_1894);
or U6165 (N_6165,N_4447,N_1984);
or U6166 (N_6166,N_3419,N_3166);
nor U6167 (N_6167,N_2397,N_830);
or U6168 (N_6168,N_4425,N_4954);
and U6169 (N_6169,N_978,N_3582);
or U6170 (N_6170,N_2421,N_1783);
nand U6171 (N_6171,N_3541,N_2496);
or U6172 (N_6172,N_2501,N_912);
and U6173 (N_6173,N_3081,N_4271);
nand U6174 (N_6174,N_3641,N_3285);
nand U6175 (N_6175,N_1628,N_3108);
nor U6176 (N_6176,N_1764,N_2357);
xor U6177 (N_6177,N_4037,N_1855);
xnor U6178 (N_6178,N_252,N_734);
xnor U6179 (N_6179,N_4602,N_3631);
nor U6180 (N_6180,N_3876,N_1936);
nand U6181 (N_6181,N_2425,N_3587);
or U6182 (N_6182,N_597,N_2317);
nand U6183 (N_6183,N_3689,N_1188);
nor U6184 (N_6184,N_1251,N_318);
and U6185 (N_6185,N_1573,N_1053);
and U6186 (N_6186,N_4491,N_1287);
nand U6187 (N_6187,N_2228,N_3110);
nor U6188 (N_6188,N_2894,N_4000);
nand U6189 (N_6189,N_865,N_4585);
nand U6190 (N_6190,N_1331,N_4881);
or U6191 (N_6191,N_2712,N_1853);
xnor U6192 (N_6192,N_1974,N_2935);
nand U6193 (N_6193,N_428,N_193);
xnor U6194 (N_6194,N_4724,N_4134);
and U6195 (N_6195,N_1240,N_703);
and U6196 (N_6196,N_1849,N_3760);
nor U6197 (N_6197,N_2093,N_4568);
or U6198 (N_6198,N_4204,N_3933);
nand U6199 (N_6199,N_3289,N_2229);
nand U6200 (N_6200,N_1312,N_664);
or U6201 (N_6201,N_2634,N_1181);
and U6202 (N_6202,N_4953,N_3934);
nor U6203 (N_6203,N_4988,N_474);
nand U6204 (N_6204,N_2120,N_4976);
xor U6205 (N_6205,N_1492,N_4767);
or U6206 (N_6206,N_1000,N_1408);
or U6207 (N_6207,N_3745,N_3279);
nand U6208 (N_6208,N_2692,N_187);
and U6209 (N_6209,N_1087,N_1671);
and U6210 (N_6210,N_3358,N_1762);
or U6211 (N_6211,N_1154,N_4573);
and U6212 (N_6212,N_436,N_4674);
xnor U6213 (N_6213,N_483,N_201);
nor U6214 (N_6214,N_4073,N_2297);
or U6215 (N_6215,N_4533,N_2781);
and U6216 (N_6216,N_1590,N_3064);
nor U6217 (N_6217,N_3857,N_4778);
nand U6218 (N_6218,N_1920,N_2502);
and U6219 (N_6219,N_575,N_3515);
nand U6220 (N_6220,N_849,N_1602);
and U6221 (N_6221,N_4720,N_4858);
and U6222 (N_6222,N_1334,N_3386);
or U6223 (N_6223,N_721,N_417);
nand U6224 (N_6224,N_1293,N_4494);
nand U6225 (N_6225,N_422,N_4322);
and U6226 (N_6226,N_2391,N_1451);
or U6227 (N_6227,N_996,N_897);
and U6228 (N_6228,N_4346,N_3545);
xor U6229 (N_6229,N_3889,N_4561);
and U6230 (N_6230,N_1178,N_4709);
and U6231 (N_6231,N_3451,N_303);
nor U6232 (N_6232,N_894,N_1329);
or U6233 (N_6233,N_1085,N_3405);
or U6234 (N_6234,N_2603,N_3646);
nand U6235 (N_6235,N_2134,N_4604);
or U6236 (N_6236,N_3512,N_581);
and U6237 (N_6237,N_56,N_2960);
and U6238 (N_6238,N_1862,N_1160);
xnor U6239 (N_6239,N_4957,N_232);
and U6240 (N_6240,N_1013,N_1564);
xnor U6241 (N_6241,N_500,N_2966);
nor U6242 (N_6242,N_3605,N_2489);
and U6243 (N_6243,N_4444,N_419);
and U6244 (N_6244,N_971,N_4782);
nor U6245 (N_6245,N_4199,N_1075);
xnor U6246 (N_6246,N_2876,N_2584);
or U6247 (N_6247,N_3055,N_1486);
xor U6248 (N_6248,N_1165,N_742);
nor U6249 (N_6249,N_2587,N_2915);
xor U6250 (N_6250,N_1850,N_4717);
nand U6251 (N_6251,N_360,N_2401);
or U6252 (N_6252,N_4521,N_1801);
and U6253 (N_6253,N_867,N_4360);
nor U6254 (N_6254,N_107,N_565);
or U6255 (N_6255,N_3235,N_754);
or U6256 (N_6256,N_3224,N_2993);
nor U6257 (N_6257,N_4284,N_2802);
nand U6258 (N_6258,N_2906,N_2929);
nand U6259 (N_6259,N_1319,N_794);
and U6260 (N_6260,N_4328,N_903);
nor U6261 (N_6261,N_3023,N_4141);
and U6262 (N_6262,N_2925,N_3997);
and U6263 (N_6263,N_375,N_795);
nand U6264 (N_6264,N_1567,N_1534);
nor U6265 (N_6265,N_4580,N_838);
and U6266 (N_6266,N_1058,N_613);
nor U6267 (N_6267,N_4902,N_2879);
or U6268 (N_6268,N_4072,N_2440);
or U6269 (N_6269,N_2554,N_2505);
or U6270 (N_6270,N_1005,N_4892);
nand U6271 (N_6271,N_1040,N_799);
nand U6272 (N_6272,N_3401,N_2978);
or U6273 (N_6273,N_4723,N_2207);
and U6274 (N_6274,N_2433,N_3053);
or U6275 (N_6275,N_2088,N_4560);
and U6276 (N_6276,N_4259,N_950);
xnor U6277 (N_6277,N_2048,N_1809);
xnor U6278 (N_6278,N_1292,N_2290);
nand U6279 (N_6279,N_472,N_626);
and U6280 (N_6280,N_2756,N_3374);
xor U6281 (N_6281,N_3839,N_560);
xnor U6282 (N_6282,N_3243,N_402);
and U6283 (N_6283,N_1473,N_1169);
nor U6284 (N_6284,N_2834,N_3270);
and U6285 (N_6285,N_693,N_2276);
or U6286 (N_6286,N_2855,N_3393);
or U6287 (N_6287,N_1533,N_335);
nand U6288 (N_6288,N_3718,N_435);
and U6289 (N_6289,N_2394,N_4361);
nor U6290 (N_6290,N_3061,N_3441);
and U6291 (N_6291,N_1637,N_4430);
and U6292 (N_6292,N_769,N_4583);
and U6293 (N_6293,N_33,N_1566);
nand U6294 (N_6294,N_3708,N_2253);
nand U6295 (N_6295,N_3354,N_4625);
nor U6296 (N_6296,N_4690,N_1554);
xnor U6297 (N_6297,N_1214,N_3182);
nand U6298 (N_6298,N_1064,N_1946);
or U6299 (N_6299,N_2652,N_4519);
or U6300 (N_6300,N_4788,N_4306);
and U6301 (N_6301,N_4197,N_4340);
xor U6302 (N_6302,N_909,N_3411);
nand U6303 (N_6303,N_2546,N_1215);
and U6304 (N_6304,N_818,N_2714);
or U6305 (N_6305,N_1004,N_1961);
nor U6306 (N_6306,N_3195,N_2808);
or U6307 (N_6307,N_4166,N_3423);
xnor U6308 (N_6308,N_3237,N_677);
and U6309 (N_6309,N_21,N_4459);
or U6310 (N_6310,N_1668,N_1581);
or U6311 (N_6311,N_3208,N_4853);
nand U6312 (N_6312,N_3734,N_3955);
or U6313 (N_6313,N_1405,N_2319);
or U6314 (N_6314,N_2448,N_707);
nor U6315 (N_6315,N_1925,N_1980);
nand U6316 (N_6316,N_4911,N_4961);
nor U6317 (N_6317,N_3261,N_4663);
and U6318 (N_6318,N_496,N_1371);
nor U6319 (N_6319,N_3174,N_1769);
nand U6320 (N_6320,N_638,N_1731);
nand U6321 (N_6321,N_2042,N_1885);
nor U6322 (N_6322,N_3347,N_4336);
nand U6323 (N_6323,N_813,N_2186);
nor U6324 (N_6324,N_4165,N_3801);
or U6325 (N_6325,N_401,N_2255);
or U6326 (N_6326,N_2611,N_4219);
and U6327 (N_6327,N_1841,N_300);
xor U6328 (N_6328,N_694,N_2462);
nor U6329 (N_6329,N_2538,N_348);
and U6330 (N_6330,N_1680,N_1593);
nand U6331 (N_6331,N_4368,N_1381);
or U6332 (N_6332,N_840,N_1387);
nand U6333 (N_6333,N_997,N_1869);
xor U6334 (N_6334,N_1026,N_3267);
or U6335 (N_6335,N_2838,N_2739);
and U6336 (N_6336,N_1069,N_1524);
nor U6337 (N_6337,N_1909,N_4362);
nor U6338 (N_6338,N_756,N_2168);
and U6339 (N_6339,N_4567,N_1126);
or U6340 (N_6340,N_153,N_4331);
nor U6341 (N_6341,N_3923,N_690);
and U6342 (N_6342,N_3236,N_2595);
xnor U6343 (N_6343,N_733,N_3342);
and U6344 (N_6344,N_3842,N_4840);
or U6345 (N_6345,N_1527,N_24);
nand U6346 (N_6346,N_3852,N_2795);
and U6347 (N_6347,N_762,N_1167);
nor U6348 (N_6348,N_506,N_4528);
nor U6349 (N_6349,N_1229,N_855);
nor U6350 (N_6350,N_3721,N_2770);
nand U6351 (N_6351,N_3488,N_2776);
nand U6352 (N_6352,N_827,N_1249);
xor U6353 (N_6353,N_4658,N_3372);
and U6354 (N_6354,N_3759,N_1539);
nor U6355 (N_6355,N_642,N_3909);
or U6356 (N_6356,N_870,N_4862);
nor U6357 (N_6357,N_1039,N_4956);
and U6358 (N_6358,N_2074,N_503);
nand U6359 (N_6359,N_1820,N_1560);
nor U6360 (N_6360,N_4679,N_2788);
and U6361 (N_6361,N_4867,N_114);
nand U6362 (N_6362,N_2248,N_2596);
xnor U6363 (N_6363,N_4609,N_954);
and U6364 (N_6364,N_1727,N_3102);
and U6365 (N_6365,N_3325,N_4208);
and U6366 (N_6366,N_1574,N_142);
nor U6367 (N_6367,N_3916,N_4118);
nand U6368 (N_6368,N_4171,N_2001);
or U6369 (N_6369,N_1814,N_4744);
and U6370 (N_6370,N_4955,N_4249);
xnor U6371 (N_6371,N_4835,N_1873);
xor U6372 (N_6372,N_1983,N_1516);
xor U6373 (N_6373,N_4379,N_886);
xnor U6374 (N_6374,N_13,N_1235);
nand U6375 (N_6375,N_3650,N_3257);
or U6376 (N_6376,N_3826,N_3319);
nor U6377 (N_6377,N_1819,N_1172);
nor U6378 (N_6378,N_1588,N_2615);
and U6379 (N_6379,N_2997,N_3046);
or U6380 (N_6380,N_1109,N_1219);
and U6381 (N_6381,N_591,N_2621);
nand U6382 (N_6382,N_4869,N_4816);
nor U6383 (N_6383,N_4588,N_4975);
nor U6384 (N_6384,N_4443,N_1875);
and U6385 (N_6385,N_312,N_2114);
or U6386 (N_6386,N_2789,N_714);
nor U6387 (N_6387,N_4986,N_2913);
and U6388 (N_6388,N_4974,N_2731);
or U6389 (N_6389,N_3389,N_4127);
and U6390 (N_6390,N_1839,N_3473);
and U6391 (N_6391,N_1582,N_612);
or U6392 (N_6392,N_2691,N_1660);
and U6393 (N_6393,N_2674,N_434);
nand U6394 (N_6394,N_3651,N_4615);
nand U6395 (N_6395,N_1745,N_3458);
nor U6396 (N_6396,N_4458,N_1477);
nand U6397 (N_6397,N_1888,N_1523);
and U6398 (N_6398,N_4366,N_4931);
xnor U6399 (N_6399,N_3229,N_645);
and U6400 (N_6400,N_1692,N_49);
nand U6401 (N_6401,N_1604,N_896);
or U6402 (N_6402,N_2975,N_4652);
and U6403 (N_6403,N_672,N_1796);
and U6404 (N_6404,N_832,N_259);
nor U6405 (N_6405,N_4807,N_3272);
nor U6406 (N_6406,N_4860,N_4831);
nand U6407 (N_6407,N_720,N_2907);
and U6408 (N_6408,N_1826,N_3341);
nand U6409 (N_6409,N_1705,N_1890);
and U6410 (N_6410,N_2859,N_3288);
and U6411 (N_6411,N_2094,N_3153);
nand U6412 (N_6412,N_4774,N_1084);
xnor U6413 (N_6413,N_4850,N_4050);
nor U6414 (N_6414,N_3250,N_3511);
and U6415 (N_6415,N_322,N_4221);
or U6416 (N_6416,N_3803,N_3167);
and U6417 (N_6417,N_549,N_1291);
nor U6418 (N_6418,N_2956,N_2185);
or U6419 (N_6419,N_378,N_994);
nor U6420 (N_6420,N_217,N_2841);
xnor U6421 (N_6421,N_3113,N_72);
nand U6422 (N_6422,N_1812,N_1609);
or U6423 (N_6423,N_835,N_2183);
or U6424 (N_6424,N_2931,N_719);
xnor U6425 (N_6425,N_4222,N_228);
or U6426 (N_6426,N_486,N_913);
nand U6427 (N_6427,N_2564,N_4462);
nand U6428 (N_6428,N_3234,N_2324);
nand U6429 (N_6429,N_2537,N_791);
xor U6430 (N_6430,N_1478,N_2460);
or U6431 (N_6431,N_517,N_1034);
or U6432 (N_6432,N_532,N_1340);
or U6433 (N_6433,N_4732,N_273);
or U6434 (N_6434,N_4581,N_2608);
and U6435 (N_6435,N_4238,N_2466);
nand U6436 (N_6436,N_2232,N_8);
xnor U6437 (N_6437,N_105,N_3030);
xnor U6438 (N_6438,N_1552,N_3679);
nand U6439 (N_6439,N_933,N_2686);
nor U6440 (N_6440,N_4994,N_2315);
nand U6441 (N_6441,N_1047,N_1701);
or U6442 (N_6442,N_4224,N_1112);
nor U6443 (N_6443,N_3636,N_1957);
and U6444 (N_6444,N_1598,N_58);
and U6445 (N_6445,N_3014,N_4055);
nand U6446 (N_6446,N_4148,N_2899);
or U6447 (N_6447,N_3703,N_4550);
nor U6448 (N_6448,N_993,N_53);
nand U6449 (N_6449,N_62,N_2839);
or U6450 (N_6450,N_1272,N_2650);
nor U6451 (N_6451,N_1966,N_4522);
xor U6452 (N_6452,N_1448,N_1663);
nor U6453 (N_6453,N_537,N_4053);
nand U6454 (N_6454,N_4039,N_552);
nor U6455 (N_6455,N_4676,N_4142);
nand U6456 (N_6456,N_666,N_4800);
and U6457 (N_6457,N_3914,N_1396);
and U6458 (N_6458,N_4917,N_2835);
xor U6459 (N_6459,N_1224,N_2017);
xor U6460 (N_6460,N_283,N_2407);
or U6461 (N_6461,N_4342,N_165);
nor U6462 (N_6462,N_1791,N_2320);
nor U6463 (N_6463,N_1986,N_699);
nor U6464 (N_6464,N_4288,N_1662);
xor U6465 (N_6465,N_1553,N_4880);
nand U6466 (N_6466,N_1792,N_1380);
or U6467 (N_6467,N_4711,N_404);
or U6468 (N_6468,N_1015,N_285);
and U6469 (N_6469,N_1360,N_3244);
or U6470 (N_6470,N_4045,N_182);
or U6471 (N_6471,N_4312,N_3742);
or U6472 (N_6472,N_4303,N_2051);
and U6473 (N_6473,N_2072,N_4333);
or U6474 (N_6474,N_1651,N_3521);
and U6475 (N_6475,N_1209,N_2814);
or U6476 (N_6476,N_274,N_2071);
or U6477 (N_6477,N_3302,N_1194);
nor U6478 (N_6478,N_2450,N_3890);
and U6479 (N_6479,N_1704,N_2892);
nor U6480 (N_6480,N_2242,N_2167);
nor U6481 (N_6481,N_4453,N_2623);
or U6482 (N_6482,N_3291,N_2665);
and U6483 (N_6483,N_1020,N_2310);
nand U6484 (N_6484,N_236,N_2649);
and U6485 (N_6485,N_1403,N_2698);
nand U6486 (N_6486,N_3448,N_1940);
and U6487 (N_6487,N_2240,N_1150);
nand U6488 (N_6488,N_1998,N_4839);
nand U6489 (N_6489,N_698,N_4442);
xor U6490 (N_6490,N_1595,N_2043);
xnor U6491 (N_6491,N_3617,N_2272);
xnor U6492 (N_6492,N_2681,N_3169);
nor U6493 (N_6493,N_60,N_1476);
xor U6494 (N_6494,N_4162,N_4098);
xor U6495 (N_6495,N_1711,N_1208);
nor U6496 (N_6496,N_4012,N_1304);
nor U6497 (N_6497,N_4640,N_302);
nand U6498 (N_6498,N_930,N_2604);
or U6499 (N_6499,N_3769,N_129);
nand U6500 (N_6500,N_4310,N_2837);
xor U6501 (N_6501,N_3036,N_4592);
or U6502 (N_6502,N_847,N_166);
nand U6503 (N_6503,N_1804,N_2928);
nand U6504 (N_6504,N_934,N_3450);
nand U6505 (N_6505,N_3829,N_2246);
nor U6506 (N_6506,N_3154,N_1547);
and U6507 (N_6507,N_2178,N_4773);
or U6508 (N_6508,N_19,N_460);
xnor U6509 (N_6509,N_2269,N_82);
and U6510 (N_6510,N_3470,N_344);
nor U6511 (N_6511,N_2312,N_1518);
xor U6512 (N_6512,N_2339,N_2774);
and U6513 (N_6513,N_1931,N_1073);
and U6514 (N_6514,N_2995,N_4755);
nand U6515 (N_6515,N_1258,N_3416);
nand U6516 (N_6516,N_4040,N_1035);
or U6517 (N_6517,N_1954,N_1390);
and U6518 (N_6518,N_3475,N_884);
and U6519 (N_6519,N_3489,N_3240);
and U6520 (N_6520,N_858,N_1159);
nand U6521 (N_6521,N_2349,N_1385);
and U6522 (N_6522,N_1550,N_4201);
or U6523 (N_6523,N_4418,N_1579);
nor U6524 (N_6524,N_1621,N_580);
and U6525 (N_6525,N_4637,N_418);
nand U6526 (N_6526,N_97,N_4746);
or U6527 (N_6527,N_359,N_917);
nand U6528 (N_6528,N_1700,N_2033);
and U6529 (N_6529,N_1096,N_623);
or U6530 (N_6530,N_265,N_3503);
or U6531 (N_6531,N_4725,N_3351);
nand U6532 (N_6532,N_1674,N_499);
and U6533 (N_6533,N_3252,N_4906);
and U6534 (N_6534,N_87,N_2981);
nor U6535 (N_6535,N_4483,N_3921);
nor U6536 (N_6536,N_4048,N_836);
nor U6537 (N_6537,N_4264,N_382);
or U6538 (N_6538,N_1227,N_1715);
nor U6539 (N_6539,N_1102,N_1364);
nor U6540 (N_6540,N_3187,N_3812);
and U6541 (N_6541,N_3365,N_7);
or U6542 (N_6542,N_3706,N_3287);
nand U6543 (N_6543,N_3947,N_970);
or U6544 (N_6544,N_3144,N_1080);
nor U6545 (N_6545,N_284,N_238);
nand U6546 (N_6546,N_4577,N_1307);
nand U6547 (N_6547,N_367,N_547);
nor U6548 (N_6548,N_2647,N_1264);
nand U6549 (N_6549,N_91,N_4158);
and U6550 (N_6550,N_646,N_25);
or U6551 (N_6551,N_116,N_3002);
and U6552 (N_6552,N_1893,N_2522);
nor U6553 (N_6553,N_2996,N_485);
nor U6554 (N_6554,N_2803,N_2792);
or U6555 (N_6555,N_1072,N_2693);
and U6556 (N_6556,N_4196,N_2285);
nor U6557 (N_6557,N_4398,N_1930);
nand U6558 (N_6558,N_2518,N_2493);
or U6559 (N_6559,N_1189,N_578);
and U6560 (N_6560,N_1864,N_1644);
nand U6561 (N_6561,N_3049,N_4244);
nor U6562 (N_6562,N_531,N_2486);
and U6563 (N_6563,N_4605,N_1741);
or U6564 (N_6564,N_4128,N_1709);
and U6565 (N_6565,N_4282,N_1962);
or U6566 (N_6566,N_584,N_518);
and U6567 (N_6567,N_3466,N_3558);
xor U6568 (N_6568,N_3695,N_4703);
or U6569 (N_6569,N_1337,N_3315);
and U6570 (N_6570,N_3606,N_2104);
and U6571 (N_6571,N_1876,N_3533);
nand U6572 (N_6572,N_4326,N_443);
and U6573 (N_6573,N_1465,N_2577);
nor U6574 (N_6574,N_41,N_1667);
and U6575 (N_6575,N_2340,N_2387);
and U6576 (N_6576,N_3363,N_3725);
or U6577 (N_6577,N_3039,N_3260);
nand U6578 (N_6578,N_1568,N_653);
and U6579 (N_6579,N_3312,N_3464);
and U6580 (N_6580,N_4595,N_1497);
and U6581 (N_6581,N_1431,N_3952);
nand U6582 (N_6582,N_4144,N_2741);
and U6583 (N_6583,N_1642,N_1994);
nor U6584 (N_6584,N_1022,N_519);
nor U6585 (N_6585,N_872,N_2481);
or U6586 (N_6586,N_2038,N_4563);
and U6587 (N_6587,N_3220,N_1402);
nand U6588 (N_6588,N_1851,N_4738);
nor U6589 (N_6589,N_2003,N_1297);
and U6590 (N_6590,N_3366,N_2787);
and U6591 (N_6591,N_3422,N_631);
nor U6592 (N_6592,N_4556,N_922);
and U6593 (N_6593,N_2010,N_2826);
nor U6594 (N_6594,N_3559,N_3067);
and U6595 (N_6595,N_1614,N_347);
nor U6596 (N_6596,N_4527,N_112);
nand U6597 (N_6597,N_2543,N_3339);
nor U6598 (N_6598,N_2527,N_4449);
or U6599 (N_6599,N_3584,N_520);
nor U6600 (N_6600,N_174,N_1245);
xor U6601 (N_6601,N_3155,N_1236);
and U6602 (N_6602,N_1024,N_1813);
nand U6603 (N_6603,N_2432,N_1255);
nand U6604 (N_6604,N_4096,N_2204);
nor U6605 (N_6605,N_2238,N_3116);
and U6606 (N_6606,N_1752,N_330);
nand U6607 (N_6607,N_459,N_676);
nor U6608 (N_6608,N_3314,N_2544);
or U6609 (N_6609,N_1036,N_753);
and U6610 (N_6610,N_3878,N_2459);
nand U6611 (N_6611,N_1908,N_2924);
xor U6612 (N_6612,N_2853,N_616);
nand U6613 (N_6613,N_4514,N_4951);
nor U6614 (N_6614,N_3664,N_3804);
xnor U6615 (N_6615,N_1223,N_2939);
or U6616 (N_6616,N_4043,N_3960);
nand U6617 (N_6617,N_3958,N_1608);
and U6618 (N_6618,N_610,N_4525);
nand U6619 (N_6619,N_516,N_3791);
and U6620 (N_6620,N_3618,N_1399);
or U6621 (N_6621,N_4358,N_1896);
or U6622 (N_6622,N_3215,N_3573);
and U6623 (N_6623,N_2937,N_4254);
and U6624 (N_6624,N_3255,N_4713);
and U6625 (N_6625,N_2723,N_257);
and U6626 (N_6626,N_1739,N_1153);
nand U6627 (N_6627,N_4349,N_1376);
or U6628 (N_6628,N_2880,N_3653);
and U6629 (N_6629,N_3031,N_821);
xor U6630 (N_6630,N_2989,N_4863);
nor U6631 (N_6631,N_2012,N_45);
nor U6632 (N_6632,N_2000,N_2047);
nand U6633 (N_6633,N_4125,N_579);
or U6634 (N_6634,N_899,N_1824);
nand U6635 (N_6635,N_3681,N_2113);
and U6636 (N_6636,N_3293,N_1496);
or U6637 (N_6637,N_2273,N_4211);
and U6638 (N_6638,N_1956,N_4536);
nand U6639 (N_6639,N_471,N_2454);
or U6640 (N_6640,N_305,N_644);
and U6641 (N_6641,N_2241,N_2684);
nor U6642 (N_6642,N_3442,N_2015);
nor U6643 (N_6643,N_2141,N_1580);
nor U6644 (N_6644,N_502,N_2342);
nand U6645 (N_6645,N_3747,N_3097);
nand U6646 (N_6646,N_80,N_1083);
or U6647 (N_6647,N_1827,N_951);
nor U6648 (N_6648,N_3991,N_3316);
nor U6649 (N_6649,N_2148,N_4992);
xor U6650 (N_6650,N_1923,N_4758);
or U6651 (N_6651,N_3041,N_4232);
and U6652 (N_6652,N_4635,N_2075);
or U6653 (N_6653,N_4747,N_3317);
nor U6654 (N_6654,N_915,N_3669);
or U6655 (N_6655,N_1678,N_4531);
or U6656 (N_6656,N_3856,N_2870);
nor U6657 (N_6657,N_2024,N_887);
or U6658 (N_6658,N_2316,N_4630);
and U6659 (N_6659,N_3908,N_1171);
nand U6660 (N_6660,N_1526,N_4613);
nor U6661 (N_6661,N_2729,N_2645);
or U6662 (N_6662,N_1025,N_495);
nand U6663 (N_6663,N_1735,N_2758);
or U6664 (N_6664,N_351,N_785);
nor U6665 (N_6665,N_1495,N_2934);
or U6666 (N_6666,N_2395,N_3825);
nand U6667 (N_6667,N_2961,N_3581);
or U6668 (N_6668,N_805,N_2305);
and U6669 (N_6669,N_1736,N_2437);
or U6670 (N_6670,N_4169,N_4965);
nand U6671 (N_6671,N_3268,N_1951);
nor U6672 (N_6672,N_1688,N_270);
and U6673 (N_6673,N_2767,N_1891);
xor U6674 (N_6674,N_427,N_3937);
nor U6675 (N_6675,N_4151,N_498);
xor U6676 (N_6676,N_2766,N_200);
or U6677 (N_6677,N_1712,N_4106);
xnor U6678 (N_6678,N_369,N_3017);
or U6679 (N_6679,N_2946,N_2601);
and U6680 (N_6680,N_3071,N_4923);
and U6681 (N_6681,N_1698,N_4783);
nand U6682 (N_6682,N_4756,N_4636);
xnor U6683 (N_6683,N_1263,N_1435);
and U6684 (N_6684,N_488,N_2576);
nor U6685 (N_6685,N_3467,N_1238);
and U6686 (N_6686,N_4015,N_688);
or U6687 (N_6687,N_1300,N_4897);
nand U6688 (N_6688,N_3369,N_2957);
nand U6689 (N_6689,N_205,N_2206);
nor U6690 (N_6690,N_919,N_143);
and U6691 (N_6691,N_3222,N_258);
nor U6692 (N_6692,N_727,N_4529);
nor U6693 (N_6693,N_3554,N_3370);
nand U6694 (N_6694,N_4242,N_4824);
or U6695 (N_6695,N_3529,N_1901);
and U6696 (N_6696,N_775,N_266);
or U6697 (N_6697,N_1675,N_635);
nand U6698 (N_6698,N_817,N_4500);
nand U6699 (N_6699,N_1177,N_4132);
or U6700 (N_6700,N_1044,N_4095);
xnor U6701 (N_6701,N_1490,N_4626);
nor U6702 (N_6702,N_3827,N_889);
nor U6703 (N_6703,N_1417,N_1419);
nor U6704 (N_6704,N_4407,N_4);
nor U6705 (N_6705,N_489,N_208);
and U6706 (N_6706,N_1124,N_2898);
and U6707 (N_6707,N_4156,N_4841);
nand U6708 (N_6708,N_3360,N_2137);
nor U6709 (N_6709,N_4659,N_1976);
nor U6710 (N_6710,N_3726,N_2617);
nand U6711 (N_6711,N_4121,N_831);
or U6712 (N_6712,N_1420,N_4091);
and U6713 (N_6713,N_1469,N_3978);
or U6714 (N_6714,N_3557,N_1811);
or U6715 (N_6715,N_4448,N_1729);
nand U6716 (N_6716,N_2388,N_2139);
nand U6717 (N_6717,N_321,N_789);
nand U6718 (N_6718,N_4918,N_4914);
nand U6719 (N_6719,N_1009,N_4105);
and U6720 (N_6720,N_3308,N_2668);
nor U6721 (N_6721,N_2118,N_643);
nor U6722 (N_6722,N_1430,N_4373);
and U6723 (N_6723,N_4634,N_2818);
nand U6724 (N_6724,N_848,N_487);
or U6725 (N_6725,N_3539,N_3713);
nor U6726 (N_6726,N_3233,N_1445);
and U6727 (N_6727,N_992,N_1111);
nand U6728 (N_6728,N_84,N_3107);
nor U6729 (N_6729,N_2364,N_380);
xor U6730 (N_6730,N_1216,N_1421);
and U6731 (N_6731,N_3776,N_4927);
nor U6732 (N_6732,N_4049,N_3597);
nand U6733 (N_6733,N_2474,N_3771);
or U6734 (N_6734,N_1468,N_3421);
nand U6735 (N_6735,N_2179,N_1563);
nor U6736 (N_6736,N_3400,N_4309);
and U6737 (N_6737,N_3306,N_844);
and U6738 (N_6738,N_390,N_853);
or U6739 (N_6739,N_4058,N_4829);
nor U6740 (N_6740,N_3426,N_2586);
and U6741 (N_6741,N_3897,N_387);
nand U6742 (N_6742,N_2335,N_4779);
nor U6743 (N_6743,N_3016,N_3823);
nor U6744 (N_6744,N_1584,N_3429);
nor U6745 (N_6745,N_3730,N_2149);
nor U6746 (N_6746,N_687,N_2581);
or U6747 (N_6747,N_4297,N_3175);
or U6748 (N_6748,N_4189,N_829);
nand U6749 (N_6749,N_3990,N_921);
nand U6750 (N_6750,N_2857,N_3238);
or U6751 (N_6751,N_1697,N_405);
or U6752 (N_6752,N_1603,N_2640);
nand U6753 (N_6753,N_4231,N_2294);
and U6754 (N_6754,N_2769,N_3197);
nor U6755 (N_6755,N_355,N_4086);
nor U6756 (N_6756,N_741,N_2445);
or U6757 (N_6757,N_1922,N_1244);
and U6758 (N_6758,N_1306,N_4294);
and U6759 (N_6759,N_652,N_536);
nor U6760 (N_6760,N_4348,N_803);
nand U6761 (N_6761,N_3540,N_393);
and U6762 (N_6762,N_1407,N_3484);
nand U6763 (N_6763,N_2657,N_1063);
or U6764 (N_6764,N_314,N_4191);
nor U6765 (N_6765,N_3171,N_963);
or U6766 (N_6766,N_4172,N_1174);
or U6767 (N_6767,N_4388,N_1078);
or U6768 (N_6768,N_2409,N_3309);
nor U6769 (N_6769,N_1462,N_410);
nand U6770 (N_6770,N_2630,N_760);
nand U6771 (N_6771,N_181,N_3739);
xor U6772 (N_6772,N_4826,N_2555);
nor U6773 (N_6773,N_4934,N_4104);
nor U6774 (N_6774,N_78,N_4825);
nor U6775 (N_6775,N_3418,N_4837);
nor U6776 (N_6776,N_4946,N_4075);
nor U6777 (N_6777,N_942,N_1166);
and U6778 (N_6778,N_2256,N_2064);
and U6779 (N_6779,N_632,N_3638);
or U6780 (N_6780,N_420,N_3868);
and U6781 (N_6781,N_3628,N_863);
nor U6782 (N_6782,N_4638,N_4727);
nor U6783 (N_6783,N_2624,N_3588);
and U6784 (N_6784,N_2734,N_1781);
and U6785 (N_6785,N_399,N_2413);
and U6786 (N_6786,N_924,N_2014);
nand U6787 (N_6787,N_851,N_1507);
or U6788 (N_6788,N_158,N_1221);
or U6789 (N_6789,N_4412,N_553);
nand U6790 (N_6790,N_414,N_4013);
nand U6791 (N_6791,N_1372,N_526);
nor U6792 (N_6792,N_408,N_1239);
nand U6793 (N_6793,N_1018,N_1914);
nor U6794 (N_6794,N_3833,N_4226);
or U6795 (N_6795,N_364,N_3821);
nor U6796 (N_6796,N_366,N_1562);
nor U6797 (N_6797,N_3874,N_2217);
nand U6798 (N_6798,N_1352,N_1546);
nand U6799 (N_6799,N_2380,N_3165);
xor U6800 (N_6800,N_2383,N_1246);
or U6801 (N_6801,N_4339,N_4478);
or U6802 (N_6802,N_3962,N_2252);
and U6803 (N_6803,N_1397,N_23);
and U6804 (N_6804,N_3256,N_1561);
nand U6805 (N_6805,N_3276,N_1086);
nand U6806 (N_6806,N_3977,N_2887);
nor U6807 (N_6807,N_3566,N_1565);
nor U6808 (N_6808,N_4100,N_4190);
xor U6809 (N_6809,N_4441,N_3663);
nor U6810 (N_6810,N_202,N_3888);
xor U6811 (N_6811,N_3553,N_1029);
nand U6812 (N_6812,N_3356,N_3230);
nand U6813 (N_6813,N_2298,N_582);
nand U6814 (N_6814,N_3367,N_1529);
and U6815 (N_6815,N_592,N_2162);
or U6816 (N_6816,N_4857,N_935);
xnor U6817 (N_6817,N_1917,N_1045);
and U6818 (N_6818,N_3029,N_2799);
or U6819 (N_6819,N_2500,N_352);
xor U6820 (N_6820,N_162,N_1302);
nor U6821 (N_6821,N_3381,N_130);
nor U6822 (N_6822,N_2172,N_1276);
nand U6823 (N_6823,N_407,N_2416);
xor U6824 (N_6824,N_306,N_4390);
nand U6825 (N_6825,N_1672,N_2196);
or U6826 (N_6826,N_3290,N_1617);
and U6827 (N_6827,N_3340,N_4941);
and U6828 (N_6828,N_3831,N_938);
nand U6829 (N_6829,N_2477,N_176);
nand U6830 (N_6830,N_700,N_4856);
nor U6831 (N_6831,N_4417,N_2745);
nand U6832 (N_6832,N_383,N_3176);
xor U6833 (N_6833,N_1415,N_4656);
and U6834 (N_6834,N_1256,N_2760);
or U6835 (N_6835,N_1280,N_2541);
xnor U6836 (N_6836,N_3622,N_2499);
or U6837 (N_6837,N_4706,N_2667);
and U6838 (N_6838,N_2023,N_747);
and U6839 (N_6839,N_3548,N_1823);
nor U6840 (N_6840,N_1059,N_4921);
nor U6841 (N_6841,N_365,N_4681);
or U6842 (N_6842,N_4299,N_2325);
nor U6843 (N_6843,N_2377,N_1959);
and U6844 (N_6844,N_3655,N_1872);
nor U6845 (N_6845,N_877,N_724);
and U6846 (N_6846,N_4545,N_4879);
and U6847 (N_6847,N_4669,N_316);
nor U6848 (N_6848,N_2921,N_4129);
xnor U6849 (N_6849,N_3927,N_2370);
xnor U6850 (N_6850,N_159,N_2266);
and U6851 (N_6851,N_2111,N_452);
and U6852 (N_6852,N_1325,N_211);
nor U6853 (N_6853,N_2551,N_3022);
nand U6854 (N_6854,N_3207,N_1439);
or U6855 (N_6855,N_1578,N_2967);
nand U6856 (N_6856,N_2999,N_3335);
nand U6857 (N_6857,N_4061,N_3784);
or U6858 (N_6858,N_295,N_2054);
nand U6859 (N_6859,N_4434,N_1549);
xor U6860 (N_6860,N_513,N_976);
nor U6861 (N_6861,N_671,N_3849);
or U6862 (N_6862,N_4594,N_898);
nand U6863 (N_6863,N_4621,N_3895);
or U6864 (N_6864,N_1377,N_3534);
nand U6865 (N_6865,N_3979,N_2182);
and U6866 (N_6866,N_4614,N_1633);
nand U6867 (N_6867,N_2659,N_4572);
nand U6868 (N_6868,N_4731,N_3980);
or U6869 (N_6869,N_475,N_3296);
xnor U6870 (N_6870,N_28,N_1232);
nand U6871 (N_6871,N_2572,N_1184);
xnor U6872 (N_6872,N_891,N_892);
nor U6873 (N_6873,N_4153,N_2165);
or U6874 (N_6874,N_1358,N_1779);
nand U6875 (N_6875,N_533,N_1691);
nor U6876 (N_6876,N_109,N_1474);
nor U6877 (N_6877,N_272,N_1097);
nor U6878 (N_6878,N_2775,N_1426);
and U6879 (N_6879,N_3614,N_973);
nor U6880 (N_6880,N_2157,N_1365);
xnor U6881 (N_6881,N_1202,N_1393);
or U6882 (N_6882,N_4277,N_2145);
or U6883 (N_6883,N_736,N_1944);
nand U6884 (N_6884,N_684,N_2087);
nor U6885 (N_6885,N_2314,N_4757);
or U6886 (N_6886,N_4737,N_1825);
nor U6887 (N_6887,N_1903,N_990);
nor U6888 (N_6888,N_3872,N_816);
nor U6889 (N_6889,N_654,N_3018);
nor U6890 (N_6890,N_608,N_2123);
nor U6891 (N_6891,N_216,N_4422);
and U6892 (N_6892,N_4035,N_3075);
and U6893 (N_6893,N_26,N_3762);
nor U6894 (N_6894,N_2824,N_3608);
or U6895 (N_6895,N_1347,N_2636);
or U6896 (N_6896,N_2707,N_2498);
or U6897 (N_6897,N_4470,N_3192);
and U6898 (N_6898,N_4698,N_3449);
nor U6899 (N_6899,N_448,N_3871);
nor U6900 (N_6900,N_4932,N_1808);
nand U6901 (N_6901,N_1844,N_2759);
or U6902 (N_6902,N_1370,N_2552);
nor U6903 (N_6903,N_3415,N_4948);
nand U6904 (N_6904,N_2453,N_2125);
nand U6905 (N_6905,N_3712,N_1099);
or U6906 (N_6906,N_4799,N_2456);
and U6907 (N_6907,N_4809,N_1228);
nand U6908 (N_6908,N_2461,N_4085);
and U6909 (N_6909,N_957,N_3008);
and U6910 (N_6910,N_313,N_31);
nor U6911 (N_6911,N_708,N_1635);
nand U6912 (N_6912,N_2475,N_3373);
or U6913 (N_6913,N_2923,N_1196);
and U6914 (N_6914,N_4024,N_2382);
xor U6915 (N_6915,N_989,N_179);
or U6916 (N_6916,N_2670,N_3474);
nor U6917 (N_6917,N_121,N_2194);
or U6918 (N_6918,N_2985,N_4643);
xor U6919 (N_6919,N_464,N_1418);
nand U6920 (N_6920,N_1681,N_4908);
nand U6921 (N_6921,N_4540,N_194);
or U6922 (N_6922,N_70,N_879);
nand U6923 (N_6923,N_2128,N_2666);
and U6924 (N_6924,N_514,N_1122);
and U6925 (N_6925,N_940,N_3196);
or U6926 (N_6926,N_3080,N_812);
xnor U6927 (N_6927,N_4705,N_3214);
and U6928 (N_6928,N_780,N_2619);
or U6929 (N_6929,N_1656,N_3948);
nand U6930 (N_6930,N_2035,N_3086);
and U6931 (N_6931,N_50,N_931);
nor U6932 (N_6932,N_3885,N_3188);
nor U6933 (N_6933,N_4597,N_2210);
nand U6934 (N_6934,N_4611,N_826);
xor U6935 (N_6935,N_1508,N_3483);
nor U6936 (N_6936,N_864,N_4051);
nand U6937 (N_6937,N_2495,N_4010);
nand U6938 (N_6938,N_1243,N_2447);
or U6939 (N_6939,N_4981,N_1843);
or U6940 (N_6940,N_4499,N_3200);
and U6941 (N_6941,N_297,N_2362);
xnor U6942 (N_6942,N_571,N_2862);
nor U6943 (N_6943,N_301,N_18);
and U6944 (N_6944,N_2955,N_4505);
nand U6945 (N_6945,N_2633,N_856);
or U6946 (N_6946,N_2274,N_4629);
or U6947 (N_6947,N_2257,N_1294);
and U6948 (N_6948,N_1683,N_89);
or U6949 (N_6949,N_479,N_2699);
and U6950 (N_6950,N_3504,N_421);
nand U6951 (N_6951,N_1969,N_4642);
nor U6952 (N_6952,N_2192,N_1932);
or U6953 (N_6953,N_1062,N_2328);
nand U6954 (N_6954,N_4535,N_2116);
nor U6955 (N_6955,N_2515,N_2525);
or U6956 (N_6956,N_2594,N_1463);
nand U6957 (N_6957,N_4030,N_3111);
nand U6958 (N_6958,N_222,N_3428);
nand U6959 (N_6959,N_2842,N_230);
or U6960 (N_6960,N_1910,N_2353);
nor U6961 (N_6961,N_1170,N_723);
and U6962 (N_6962,N_3269,N_1301);
and U6963 (N_6963,N_2726,N_3772);
nor U6964 (N_6964,N_2910,N_660);
nor U6965 (N_6965,N_1973,N_444);
and U6966 (N_6966,N_3355,N_4847);
xor U6967 (N_6967,N_710,N_3932);
nor U6968 (N_6968,N_2533,N_3026);
nand U6969 (N_6969,N_2949,N_170);
or U6970 (N_6970,N_1548,N_218);
and U6971 (N_6971,N_1506,N_4071);
nand U6972 (N_6972,N_4246,N_247);
and U6973 (N_6973,N_3476,N_1139);
and U6974 (N_6974,N_3994,N_2885);
nor U6975 (N_6975,N_1113,N_4903);
nand U6976 (N_6976,N_1937,N_457);
and U6977 (N_6977,N_4261,N_1877);
nor U6978 (N_6978,N_2648,N_3738);
nand U6979 (N_6979,N_3514,N_4949);
nand U6980 (N_6980,N_2883,N_136);
or U6981 (N_6981,N_4617,N_1654);
or U6982 (N_6982,N_315,N_146);
xnor U6983 (N_6983,N_3060,N_4532);
nand U6984 (N_6984,N_1916,N_4429);
or U6985 (N_6985,N_4612,N_2535);
or U6986 (N_6986,N_4136,N_3051);
nand U6987 (N_6987,N_4827,N_4255);
or U6988 (N_6988,N_3785,N_3127);
and U6989 (N_6989,N_901,N_3324);
xor U6990 (N_6990,N_4904,N_2301);
or U6991 (N_6991,N_4770,N_163);
or U6992 (N_6992,N_3859,N_3781);
nand U6993 (N_6993,N_1702,N_215);
or U6994 (N_6994,N_323,N_3717);
or U6995 (N_6995,N_1605,N_4771);
or U6996 (N_6996,N_509,N_3579);
nand U6997 (N_6997,N_4714,N_4665);
or U6998 (N_6998,N_3975,N_4335);
or U6999 (N_6999,N_2078,N_1367);
and U7000 (N_7000,N_2,N_3241);
nor U7001 (N_7001,N_4970,N_521);
nor U7002 (N_7002,N_2994,N_4693);
and U7003 (N_7003,N_3392,N_2164);
and U7004 (N_7004,N_4408,N_2046);
and U7005 (N_7005,N_1716,N_2736);
or U7006 (N_7006,N_54,N_3682);
and U7007 (N_7007,N_3158,N_4327);
and U7008 (N_7008,N_4963,N_1519);
nand U7009 (N_7009,N_92,N_3305);
nor U7010 (N_7010,N_1330,N_2771);
or U7011 (N_7011,N_337,N_1285);
nand U7012 (N_7012,N_3550,N_4960);
nor U7013 (N_7013,N_3122,N_2836);
or U7014 (N_7014,N_99,N_2591);
and U7015 (N_7015,N_3435,N_2262);
nor U7016 (N_7016,N_1144,N_2326);
and U7017 (N_7017,N_3775,N_4644);
nand U7018 (N_7018,N_607,N_3925);
or U7019 (N_7019,N_3066,N_4873);
nand U7020 (N_7020,N_3178,N_237);
or U7021 (N_7021,N_2588,N_1897);
and U7022 (N_7022,N_2563,N_3692);
and U7023 (N_7023,N_224,N_3817);
nand U7024 (N_7024,N_4761,N_4397);
nor U7025 (N_7025,N_1446,N_4028);
or U7026 (N_7026,N_2423,N_3986);
nand U7027 (N_7027,N_3444,N_3595);
nor U7028 (N_7028,N_3846,N_4622);
or U7029 (N_7029,N_3035,N_678);
nor U7030 (N_7030,N_101,N_2265);
nand U7031 (N_7031,N_4138,N_4805);
xnor U7032 (N_7032,N_3911,N_2557);
and U7033 (N_7033,N_279,N_4022);
and U7034 (N_7034,N_3058,N_1412);
xnor U7035 (N_7035,N_525,N_2483);
nand U7036 (N_7036,N_3000,N_1261);
and U7037 (N_7037,N_354,N_2209);
and U7038 (N_7038,N_3993,N_1149);
and U7039 (N_7039,N_3331,N_4610);
nand U7040 (N_7040,N_2089,N_233);
nor U7041 (N_7041,N_4243,N_3531);
nor U7042 (N_7042,N_3,N_4350);
nor U7043 (N_7043,N_2965,N_4766);
or U7044 (N_7044,N_3501,N_2813);
or U7045 (N_7045,N_1631,N_2414);
nand U7046 (N_7046,N_1721,N_3388);
nor U7047 (N_7047,N_287,N_569);
or U7048 (N_7048,N_640,N_3399);
or U7049 (N_7049,N_2277,N_2323);
nand U7050 (N_7050,N_3385,N_4359);
nand U7051 (N_7051,N_2221,N_1832);
nand U7052 (N_7052,N_4393,N_242);
and U7053 (N_7053,N_1432,N_3311);
xor U7054 (N_7054,N_3522,N_4257);
xnor U7055 (N_7055,N_4068,N_1487);
nand U7056 (N_7056,N_883,N_4070);
nand U7057 (N_7057,N_1274,N_4952);
and U7058 (N_7058,N_3038,N_3619);
or U7059 (N_7059,N_1193,N_2976);
xnor U7060 (N_7060,N_195,N_4414);
nand U7061 (N_7061,N_2593,N_4823);
and U7062 (N_7062,N_3181,N_648);
nor U7063 (N_7063,N_4214,N_2547);
nor U7064 (N_7064,N_2070,N_1991);
or U7065 (N_7065,N_4736,N_4542);
and U7066 (N_7066,N_1532,N_1601);
nand U7067 (N_7067,N_2513,N_4938);
or U7068 (N_7068,N_4672,N_2682);
and U7069 (N_7069,N_1313,N_2131);
and U7070 (N_7070,N_2251,N_234);
nor U7071 (N_7071,N_3477,N_4620);
and U7072 (N_7072,N_172,N_2441);
and U7073 (N_7073,N_2678,N_3929);
and U7074 (N_7074,N_1610,N_4081);
nand U7075 (N_7075,N_2806,N_4212);
and U7076 (N_7076,N_212,N_4280);
and U7077 (N_7077,N_22,N_1907);
nor U7078 (N_7078,N_587,N_4376);
or U7079 (N_7079,N_1733,N_3671);
nor U7080 (N_7080,N_797,N_1848);
xnor U7081 (N_7081,N_3995,N_3709);
nor U7082 (N_7082,N_2655,N_2677);
xor U7083 (N_7083,N_2874,N_717);
nor U7084 (N_7084,N_152,N_144);
and U7085 (N_7085,N_4872,N_4985);
xor U7086 (N_7086,N_3604,N_991);
nand U7087 (N_7087,N_3698,N_3094);
nor U7088 (N_7088,N_4324,N_1357);
nor U7089 (N_7089,N_357,N_4933);
nand U7090 (N_7090,N_4077,N_3431);
and U7091 (N_7091,N_3691,N_3228);
or U7092 (N_7092,N_3901,N_3798);
nor U7093 (N_7093,N_3987,N_2053);
and U7094 (N_7094,N_4396,N_878);
and U7095 (N_7095,N_4295,N_1622);
nand U7096 (N_7096,N_4962,N_2823);
nand U7097 (N_7097,N_4806,N_1645);
and U7098 (N_7098,N_3119,N_3917);
xnor U7099 (N_7099,N_52,N_4205);
and U7100 (N_7100,N_3525,N_783);
or U7101 (N_7101,N_320,N_3263);
nand U7102 (N_7102,N_2487,N_1220);
and U7103 (N_7103,N_1100,N_2029);
nand U7104 (N_7104,N_319,N_728);
nand U7105 (N_7105,N_2205,N_1320);
and U7106 (N_7106,N_1296,N_2641);
or U7107 (N_7107,N_2299,N_1237);
or U7108 (N_7108,N_1428,N_2730);
and U7109 (N_7109,N_956,N_2507);
and U7110 (N_7110,N_2616,N_4964);
or U7111 (N_7111,N_4252,N_1594);
nor U7112 (N_7112,N_3616,N_4822);
or U7113 (N_7113,N_1206,N_4808);
nand U7114 (N_7114,N_4855,N_2752);
or U7115 (N_7115,N_1363,N_346);
nor U7116 (N_7116,N_2398,N_4122);
nand U7117 (N_7117,N_3223,N_2825);
nand U7118 (N_7118,N_3266,N_2187);
nor U7119 (N_7119,N_4664,N_2231);
nor U7120 (N_7120,N_304,N_3887);
or U7121 (N_7121,N_3164,N_2140);
nor U7122 (N_7122,N_2658,N_1384);
nand U7123 (N_7123,N_2082,N_2309);
xor U7124 (N_7124,N_2637,N_1763);
and U7125 (N_7125,N_2058,N_802);
nand U7126 (N_7126,N_1310,N_3836);
and U7127 (N_7127,N_3019,N_1935);
xnor U7128 (N_7128,N_761,N_1314);
and U7129 (N_7129,N_2534,N_985);
and U7130 (N_7130,N_3479,N_1616);
nand U7131 (N_7131,N_5,N_1510);
nand U7132 (N_7132,N_1142,N_104);
xor U7133 (N_7133,N_3310,N_2363);
xnor U7134 (N_7134,N_4687,N_44);
xnor U7135 (N_7135,N_3262,N_4287);
and U7136 (N_7136,N_1484,N_3976);
or U7137 (N_7137,N_3005,N_4993);
nand U7138 (N_7138,N_227,N_3844);
xnor U7139 (N_7139,N_4292,N_3544);
xnor U7140 (N_7140,N_1722,N_1625);
nor U7141 (N_7141,N_866,N_125);
or U7142 (N_7142,N_397,N_1379);
nor U7143 (N_7143,N_4052,N_4796);
and U7144 (N_7144,N_3073,N_3286);
nand U7145 (N_7145,N_2171,N_1281);
xnor U7146 (N_7146,N_3870,N_3417);
nor U7147 (N_7147,N_127,N_2860);
or U7148 (N_7148,N_4147,N_2783);
or U7149 (N_7149,N_594,N_4227);
nand U7150 (N_7150,N_2550,N_490);
and U7151 (N_7151,N_2464,N_4026);
or U7152 (N_7152,N_2090,N_3109);
xnor U7153 (N_7153,N_2560,N_2184);
or U7154 (N_7154,N_4977,N_2948);
or U7155 (N_7155,N_1856,N_157);
nor U7156 (N_7156,N_4477,N_1795);
nand U7157 (N_7157,N_510,N_745);
nor U7158 (N_7158,N_4371,N_4557);
nor U7159 (N_7159,N_4198,N_2809);
or U7160 (N_7160,N_2800,N_1934);
nand U7161 (N_7161,N_4181,N_3774);
nor U7162 (N_7162,N_2865,N_3674);
xor U7163 (N_7163,N_2718,N_1943);
nand U7164 (N_7164,N_1686,N_2085);
xor U7165 (N_7165,N_4063,N_3225);
xnor U7166 (N_7166,N_470,N_1776);
nand U7167 (N_7167,N_3583,N_4631);
nor U7168 (N_7168,N_371,N_670);
xor U7169 (N_7169,N_482,N_4437);
nor U7170 (N_7170,N_3964,N_2115);
and U7171 (N_7171,N_3170,N_3699);
or U7172 (N_7172,N_3120,N_1414);
xor U7173 (N_7173,N_2972,N_4884);
nor U7174 (N_7174,N_1615,N_3571);
and U7175 (N_7175,N_3850,N_1928);
and U7176 (N_7176,N_4524,N_1572);
nor U7177 (N_7177,N_2822,N_2503);
and U7178 (N_7178,N_4896,N_2348);
nand U7179 (N_7179,N_4195,N_3070);
xor U7180 (N_7180,N_4463,N_2067);
or U7181 (N_7181,N_1373,N_1309);
nor U7182 (N_7182,N_2203,N_102);
nand U7183 (N_7183,N_860,N_1768);
or U7184 (N_7184,N_2109,N_3398);
and U7185 (N_7185,N_256,N_3377);
or U7186 (N_7186,N_999,N_1528);
and U7187 (N_7187,N_191,N_1880);
xor U7188 (N_7188,N_4381,N_2020);
and U7189 (N_7189,N_3818,N_4812);
xor U7190 (N_7190,N_4038,N_1176);
nor U7191 (N_7191,N_1106,N_1737);
xor U7192 (N_7192,N_3562,N_801);
xnor U7193 (N_7193,N_3380,N_3149);
nand U7194 (N_7194,N_4234,N_3409);
or U7195 (N_7195,N_3350,N_4188);
and U7196 (N_7196,N_4021,N_2119);
and U7197 (N_7197,N_1924,N_4979);
nor U7198 (N_7198,N_2302,N_962);
xor U7199 (N_7199,N_4670,N_294);
and U7200 (N_7200,N_529,N_2284);
or U7201 (N_7201,N_4307,N_685);
nand U7202 (N_7202,N_4870,N_379);
xnor U7203 (N_7203,N_4900,N_3576);
xor U7204 (N_7204,N_2002,N_3510);
xnor U7205 (N_7205,N_1213,N_4409);
or U7206 (N_7206,N_1339,N_2040);
and U7207 (N_7207,N_1749,N_3199);
nor U7208 (N_7208,N_4404,N_893);
nand U7209 (N_7209,N_1461,N_2127);
nor U7210 (N_7210,N_2237,N_634);
nor U7211 (N_7211,N_808,N_2393);
and U7212 (N_7212,N_3201,N_3808);
and U7213 (N_7213,N_3118,N_1146);
nor U7214 (N_7214,N_3148,N_1278);
nand U7215 (N_7215,N_267,N_3981);
and U7216 (N_7216,N_173,N_1778);
and U7217 (N_7217,N_473,N_1509);
or U7218 (N_7218,N_3227,N_1141);
and U7219 (N_7219,N_3083,N_4632);
and U7220 (N_7220,N_4842,N_3809);
and U7221 (N_7221,N_2189,N_3580);
nand U7222 (N_7222,N_2032,N_875);
xor U7223 (N_7223,N_1670,N_260);
nor U7224 (N_7224,N_2793,N_3209);
and U7225 (N_7225,N_3943,N_4452);
and U7226 (N_7226,N_175,N_4355);
or U7227 (N_7227,N_788,N_3130);
and U7228 (N_7228,N_148,N_1362);
or U7229 (N_7229,N_3794,N_918);
nor U7230 (N_7230,N_1233,N_4385);
nand U7231 (N_7231,N_3146,N_3838);
nand U7232 (N_7232,N_904,N_2400);
and U7233 (N_7233,N_601,N_4167);
xor U7234 (N_7234,N_3970,N_1992);
or U7235 (N_7235,N_381,N_2625);
and U7236 (N_7236,N_37,N_4082);
nor U7237 (N_7237,N_2296,N_4062);
xor U7238 (N_7238,N_998,N_4694);
or U7239 (N_7239,N_150,N_3967);
and U7240 (N_7240,N_1290,N_2845);
xor U7241 (N_7241,N_1438,N_461);
nand U7242 (N_7242,N_3560,N_197);
nor U7243 (N_7243,N_1685,N_1356);
or U7244 (N_7244,N_1540,N_440);
and U7245 (N_7245,N_2063,N_2703);
xor U7246 (N_7246,N_3920,N_2598);
or U7247 (N_7247,N_2036,N_2016);
nor U7248 (N_7248,N_1288,N_1343);
and U7249 (N_7249,N_115,N_4256);
and U7250 (N_7250,N_3780,N_3247);
nand U7251 (N_7251,N_936,N_3707);
nor U7252 (N_7252,N_3134,N_2600);
nor U7253 (N_7253,N_2701,N_2798);
nor U7254 (N_7254,N_564,N_1267);
nor U7255 (N_7255,N_1665,N_1076);
and U7256 (N_7256,N_2068,N_3939);
or U7257 (N_7257,N_1116,N_2359);
nor U7258 (N_7258,N_3782,N_2458);
or U7259 (N_7259,N_4207,N_1021);
nor U7260 (N_7260,N_3103,N_4741);
and U7261 (N_7261,N_512,N_3624);
nor U7262 (N_7262,N_620,N_3211);
or U7263 (N_7263,N_2969,N_2249);
nor U7264 (N_7264,N_249,N_530);
nand U7265 (N_7265,N_2896,N_2627);
and U7266 (N_7266,N_4601,N_1638);
nand U7267 (N_7267,N_3472,N_2402);
or U7268 (N_7268,N_4154,N_3524);
nor U7269 (N_7269,N_544,N_3959);
nand U7270 (N_7270,N_4668,N_602);
nand U7271 (N_7271,N_1995,N_2399);
nor U7272 (N_7272,N_3420,N_2785);
and U7273 (N_7273,N_332,N_1785);
xor U7274 (N_7274,N_4901,N_4120);
nor U7275 (N_7275,N_4384,N_3394);
or U7276 (N_7276,N_2590,N_2519);
nand U7277 (N_7277,N_1156,N_2711);
and U7278 (N_7278,N_1117,N_1162);
and U7279 (N_7279,N_2260,N_3328);
and U7280 (N_7280,N_171,N_4431);
nor U7281 (N_7281,N_3757,N_3033);
nand U7282 (N_7282,N_2190,N_3040);
or U7283 (N_7283,N_1870,N_4330);
and U7284 (N_7284,N_4883,N_1342);
nand U7285 (N_7285,N_3732,N_1335);
nand U7286 (N_7286,N_1952,N_3463);
nand U7287 (N_7287,N_4293,N_2958);
or U7288 (N_7288,N_4338,N_4131);
nor U7289 (N_7289,N_2286,N_2345);
and U7290 (N_7290,N_2954,N_458);
nor U7291 (N_7291,N_3678,N_1359);
and U7292 (N_7292,N_3924,N_1032);
xnor U7293 (N_7293,N_4002,N_977);
or U7294 (N_7294,N_4176,N_3592);
or U7295 (N_7295,N_958,N_2610);
and U7296 (N_7296,N_869,N_843);
nand U7297 (N_7297,N_2653,N_3156);
or U7298 (N_7298,N_2721,N_3865);
and U7299 (N_7299,N_824,N_1161);
or U7300 (N_7300,N_2943,N_291);
nand U7301 (N_7301,N_2990,N_2045);
or U7302 (N_7302,N_2412,N_2574);
and U7303 (N_7303,N_722,N_3378);
and U7304 (N_7304,N_3065,N_596);
or U7305 (N_7305,N_3935,N_3851);
xor U7306 (N_7306,N_3206,N_982);
and U7307 (N_7307,N_2198,N_4980);
nor U7308 (N_7308,N_2355,N_4763);
nor U7309 (N_7309,N_3723,N_465);
or U7310 (N_7310,N_541,N_4777);
and U7311 (N_7311,N_1743,N_2436);
nor U7312 (N_7312,N_2378,N_4092);
or U7313 (N_7313,N_4591,N_955);
or U7314 (N_7314,N_595,N_3658);
xor U7315 (N_7315,N_2982,N_188);
and U7316 (N_7316,N_1717,N_4875);
nor U7317 (N_7317,N_1505,N_1724);
xor U7318 (N_7318,N_4552,N_2208);
nor U7319 (N_7319,N_682,N_4661);
xor U7320 (N_7320,N_384,N_1001);
and U7321 (N_7321,N_4995,N_2744);
or U7322 (N_7322,N_2086,N_3815);
nor U7323 (N_7323,N_1703,N_2549);
nand U7324 (N_7324,N_3906,N_1606);
nand U7325 (N_7325,N_1673,N_1569);
nand U7326 (N_7326,N_3632,N_226);
nor U7327 (N_7327,N_2226,N_3621);
nand U7328 (N_7328,N_4276,N_231);
or U7329 (N_7329,N_1653,N_3433);
nor U7330 (N_7330,N_67,N_4119);
nand U7331 (N_7331,N_4143,N_3685);
and U7332 (N_7332,N_4987,N_941);
nand U7333 (N_7333,N_1191,N_2429);
nand U7334 (N_7334,N_4216,N_4356);
or U7335 (N_7335,N_2011,N_1536);
or U7336 (N_7336,N_572,N_2471);
nor U7337 (N_7337,N_3940,N_3487);
nor U7338 (N_7338,N_2479,N_4263);
xnor U7339 (N_7339,N_3665,N_1815);
or U7340 (N_7340,N_952,N_1388);
and U7341 (N_7341,N_1821,N_1759);
nand U7342 (N_7342,N_57,N_2877);
nand U7343 (N_7343,N_3969,N_4289);
and U7344 (N_7344,N_636,N_706);
nor U7345 (N_7345,N_4087,N_29);
and U7346 (N_7346,N_4103,N_1185);
and U7347 (N_7347,N_1252,N_3530);
and U7348 (N_7348,N_910,N_3439);
nand U7349 (N_7349,N_3434,N_2373);
or U7350 (N_7350,N_3082,N_1757);
or U7351 (N_7351,N_2417,N_2644);
and U7352 (N_7352,N_3042,N_2827);
and U7353 (N_7353,N_3452,N_1857);
and U7354 (N_7354,N_4876,N_1558);
or U7355 (N_7355,N_2102,N_4427);
nor U7356 (N_7356,N_3430,N_2768);
nor U7357 (N_7357,N_4707,N_2858);
xor U7358 (N_7358,N_3496,N_3644);
nor U7359 (N_7359,N_2833,N_1002);
or U7360 (N_7360,N_3432,N_3961);
nand U7361 (N_7361,N_3085,N_3567);
and U7362 (N_7362,N_3593,N_1542);
and U7363 (N_7363,N_811,N_4258);
nand U7364 (N_7364,N_3105,N_599);
or U7365 (N_7365,N_4486,N_3406);
and U7366 (N_7366,N_4947,N_4046);
and U7367 (N_7367,N_4754,N_1234);
or U7368 (N_7368,N_4877,N_1043);
nor U7369 (N_7369,N_4913,N_3295);
nor U7370 (N_7370,N_2278,N_2871);
xnor U7371 (N_7371,N_624,N_1299);
and U7372 (N_7372,N_468,N_3191);
nand U7373 (N_7373,N_4485,N_3054);
nand U7374 (N_7374,N_1955,N_3088);
nand U7375 (N_7375,N_543,N_2794);
xnor U7376 (N_7376,N_2013,N_110);
or U7377 (N_7377,N_3121,N_2580);
and U7378 (N_7378,N_3778,N_3499);
xnor U7379 (N_7379,N_3740,N_528);
or U7380 (N_7380,N_3919,N_3427);
nor U7381 (N_7381,N_2236,N_4251);
and U7382 (N_7382,N_4716,N_1647);
or U7383 (N_7383,N_288,N_4069);
or U7384 (N_7384,N_3232,N_4689);
nor U7385 (N_7385,N_4795,N_1345);
nand U7386 (N_7386,N_1225,N_4558);
nor U7387 (N_7387,N_4971,N_4240);
nor U7388 (N_7388,N_1248,N_4399);
nand U7389 (N_7389,N_1699,N_3204);
or U7390 (N_7390,N_4794,N_2709);
nand U7391 (N_7391,N_1975,N_2567);
nand U7392 (N_7392,N_4423,N_1918);
nor U7393 (N_7393,N_1655,N_2901);
or U7394 (N_7394,N_2884,N_4250);
nor U7395 (N_7395,N_3673,N_2386);
nor U7396 (N_7396,N_4537,N_3205);
nand U7397 (N_7397,N_2812,N_2470);
xor U7398 (N_7398,N_4146,N_120);
nor U7399 (N_7399,N_617,N_4210);
nand U7400 (N_7400,N_190,N_4497);
and U7401 (N_7401,N_4117,N_1677);
nor U7402 (N_7402,N_3034,N_4369);
nor U7403 (N_7403,N_4919,N_4677);
xor U7404 (N_7404,N_1147,N_534);
or U7405 (N_7405,N_3245,N_1128);
nand U7406 (N_7406,N_1658,N_3440);
and U7407 (N_7407,N_271,N_3376);
nand U7408 (N_7408,N_1455,N_4786);
nor U7409 (N_7409,N_895,N_3668);
or U7410 (N_7410,N_3637,N_1351);
nor U7411 (N_7411,N_3259,N_1282);
nor U7412 (N_7412,N_3657,N_4916);
xor U7413 (N_7413,N_1836,N_932);
or U7414 (N_7414,N_1410,N_1775);
xnor U7415 (N_7415,N_3179,N_2508);
or U7416 (N_7416,N_4798,N_3322);
nand U7417 (N_7417,N_3840,N_4027);
xnor U7418 (N_7418,N_1993,N_4218);
nand U7419 (N_7419,N_4559,N_206);
nor U7420 (N_7420,N_751,N_3517);
nor U7421 (N_7421,N_598,N_3194);
and U7422 (N_7422,N_1218,N_4868);
nor U7423 (N_7423,N_3661,N_1793);
and U7424 (N_7424,N_1118,N_11);
nor U7425 (N_7425,N_1152,N_1369);
nand U7426 (N_7426,N_2951,N_854);
xnor U7427 (N_7427,N_1226,N_203);
and U7428 (N_7428,N_3667,N_1591);
or U7429 (N_7429,N_317,N_629);
nand U7430 (N_7430,N_1720,N_3093);
xnor U7431 (N_7431,N_3044,N_2683);
nand U7432 (N_7432,N_2545,N_1204);
and U7433 (N_7433,N_3974,N_3561);
nor U7434 (N_7434,N_1765,N_3898);
nor U7435 (N_7435,N_3710,N_4334);
nand U7436 (N_7436,N_2964,N_609);
nand U7437 (N_7437,N_839,N_823);
nor U7438 (N_7438,N_3918,N_4089);
and U7439 (N_7439,N_4260,N_1555);
nor U7440 (N_7440,N_1201,N_2852);
xnor U7441 (N_7441,N_4878,N_2154);
nor U7442 (N_7442,N_3596,N_1471);
nand U7443 (N_7443,N_2605,N_1052);
xor U7444 (N_7444,N_2482,N_4762);
nor U7445 (N_7445,N_391,N_1454);
or U7446 (N_7446,N_1450,N_4387);
nor U7447 (N_7447,N_1707,N_3333);
nor U7448 (N_7448,N_3945,N_1046);
nand U7449 (N_7449,N_2280,N_4516);
and U7450 (N_7450,N_361,N_2166);
xor U7451 (N_7451,N_2639,N_3694);
and U7452 (N_7452,N_1898,N_920);
and U7453 (N_7453,N_43,N_539);
and U7454 (N_7454,N_1483,N_2026);
nor U7455 (N_7455,N_1960,N_4688);
or U7456 (N_7456,N_1289,N_1833);
and U7457 (N_7457,N_1545,N_2156);
or U7458 (N_7458,N_4116,N_4229);
or U7459 (N_7459,N_1912,N_781);
and U7460 (N_7460,N_2143,N_1132);
and U7461 (N_7461,N_1442,N_3136);
and U7462 (N_7462,N_2713,N_4126);
and U7463 (N_7463,N_395,N_3748);
and U7464 (N_7464,N_2930,N_4493);
xor U7465 (N_7465,N_655,N_861);
nor U7466 (N_7466,N_47,N_1003);
nand U7467 (N_7467,N_253,N_4748);
xnor U7468 (N_7468,N_3765,N_3186);
and U7469 (N_7469,N_1378,N_1050);
and U7470 (N_7470,N_2295,N_2660);
xor U7471 (N_7471,N_558,N_4726);
nand U7472 (N_7472,N_1852,N_1413);
nand U7473 (N_7473,N_984,N_3402);
nand U7474 (N_7474,N_4203,N_3570);
nand U7475 (N_7475,N_1988,N_1889);
xnor U7476 (N_7476,N_1103,N_3750);
or U7477 (N_7477,N_2193,N_3720);
nand U7478 (N_7478,N_1323,N_276);
xnor U7479 (N_7479,N_4651,N_2786);
nor U7480 (N_7480,N_1965,N_1187);
nor U7481 (N_7481,N_398,N_1657);
nor U7482 (N_7482,N_3700,N_4697);
nand U7483 (N_7483,N_77,N_1514);
and U7484 (N_7484,N_4042,N_3509);
and U7485 (N_7485,N_1437,N_1346);
nand U7486 (N_7486,N_415,N_345);
or U7487 (N_7487,N_3349,N_3883);
nor U7488 (N_7488,N_2219,N_3647);
nand U7489 (N_7489,N_508,N_1537);
or U7490 (N_7490,N_1270,N_1382);
nand U7491 (N_7491,N_2509,N_656);
nor U7492 (N_7492,N_2467,N_3012);
or U7493 (N_7493,N_772,N_4912);
or U7494 (N_7494,N_3629,N_2643);
nand U7495 (N_7495,N_1125,N_3946);
or U7496 (N_7496,N_3749,N_2136);
nor U7497 (N_7497,N_4520,N_356);
nor U7498 (N_7498,N_779,N_3770);
nor U7499 (N_7499,N_1266,N_4926);
and U7500 (N_7500,N_3902,N_1208);
nor U7501 (N_7501,N_4310,N_4708);
nand U7502 (N_7502,N_2691,N_2162);
or U7503 (N_7503,N_1062,N_4127);
or U7504 (N_7504,N_4993,N_2063);
or U7505 (N_7505,N_97,N_4336);
nand U7506 (N_7506,N_4683,N_2233);
nand U7507 (N_7507,N_1290,N_2219);
xor U7508 (N_7508,N_1813,N_4736);
or U7509 (N_7509,N_1689,N_3193);
xnor U7510 (N_7510,N_1093,N_1031);
nor U7511 (N_7511,N_2646,N_1061);
nand U7512 (N_7512,N_725,N_3904);
and U7513 (N_7513,N_643,N_3224);
and U7514 (N_7514,N_346,N_3762);
and U7515 (N_7515,N_4480,N_1842);
or U7516 (N_7516,N_1096,N_1659);
xnor U7517 (N_7517,N_4603,N_3465);
nor U7518 (N_7518,N_1150,N_1037);
and U7519 (N_7519,N_577,N_3969);
nand U7520 (N_7520,N_3407,N_393);
nor U7521 (N_7521,N_2386,N_1469);
or U7522 (N_7522,N_4093,N_1697);
and U7523 (N_7523,N_1563,N_4807);
and U7524 (N_7524,N_3317,N_100);
and U7525 (N_7525,N_389,N_4537);
and U7526 (N_7526,N_776,N_926);
nand U7527 (N_7527,N_1264,N_3277);
nand U7528 (N_7528,N_3556,N_2897);
nor U7529 (N_7529,N_2903,N_2182);
or U7530 (N_7530,N_870,N_1681);
nand U7531 (N_7531,N_1393,N_1345);
nor U7532 (N_7532,N_4803,N_3156);
nand U7533 (N_7533,N_457,N_4996);
nor U7534 (N_7534,N_529,N_3254);
and U7535 (N_7535,N_2743,N_628);
nor U7536 (N_7536,N_2230,N_2805);
nand U7537 (N_7537,N_95,N_2271);
xor U7538 (N_7538,N_3274,N_3631);
and U7539 (N_7539,N_4232,N_2931);
and U7540 (N_7540,N_4473,N_1942);
and U7541 (N_7541,N_2589,N_4852);
or U7542 (N_7542,N_217,N_389);
nor U7543 (N_7543,N_2004,N_4448);
or U7544 (N_7544,N_11,N_4634);
nor U7545 (N_7545,N_2517,N_2002);
and U7546 (N_7546,N_3887,N_3085);
xnor U7547 (N_7547,N_4634,N_2897);
and U7548 (N_7548,N_2048,N_1390);
nand U7549 (N_7549,N_3527,N_469);
nand U7550 (N_7550,N_2974,N_3612);
or U7551 (N_7551,N_3739,N_4506);
and U7552 (N_7552,N_100,N_2476);
nor U7553 (N_7553,N_1670,N_4744);
or U7554 (N_7554,N_1207,N_3164);
xor U7555 (N_7555,N_2547,N_4310);
nor U7556 (N_7556,N_416,N_2608);
xnor U7557 (N_7557,N_3311,N_3641);
xnor U7558 (N_7558,N_499,N_3992);
nor U7559 (N_7559,N_2468,N_4060);
and U7560 (N_7560,N_4349,N_1733);
nand U7561 (N_7561,N_158,N_2402);
or U7562 (N_7562,N_1801,N_3544);
and U7563 (N_7563,N_4168,N_3413);
and U7564 (N_7564,N_3912,N_2183);
and U7565 (N_7565,N_2244,N_4317);
nor U7566 (N_7566,N_2790,N_2663);
nand U7567 (N_7567,N_286,N_4140);
nand U7568 (N_7568,N_1497,N_418);
and U7569 (N_7569,N_3460,N_10);
and U7570 (N_7570,N_4988,N_2095);
nand U7571 (N_7571,N_1568,N_1107);
and U7572 (N_7572,N_4911,N_4219);
and U7573 (N_7573,N_3230,N_4288);
or U7574 (N_7574,N_845,N_1969);
and U7575 (N_7575,N_1662,N_2932);
or U7576 (N_7576,N_3887,N_38);
nor U7577 (N_7577,N_3457,N_1150);
or U7578 (N_7578,N_1824,N_1479);
and U7579 (N_7579,N_4838,N_1831);
or U7580 (N_7580,N_4658,N_2615);
or U7581 (N_7581,N_2279,N_1830);
nand U7582 (N_7582,N_977,N_3031);
and U7583 (N_7583,N_1401,N_391);
nand U7584 (N_7584,N_890,N_968);
and U7585 (N_7585,N_3408,N_4268);
and U7586 (N_7586,N_3440,N_3304);
and U7587 (N_7587,N_593,N_1265);
nor U7588 (N_7588,N_3489,N_2249);
and U7589 (N_7589,N_3730,N_1491);
nor U7590 (N_7590,N_4522,N_2963);
or U7591 (N_7591,N_3404,N_2931);
nor U7592 (N_7592,N_1783,N_412);
nand U7593 (N_7593,N_4590,N_4918);
xnor U7594 (N_7594,N_2503,N_4881);
nor U7595 (N_7595,N_980,N_1454);
nand U7596 (N_7596,N_3730,N_1532);
or U7597 (N_7597,N_3370,N_525);
and U7598 (N_7598,N_4941,N_4561);
or U7599 (N_7599,N_464,N_4618);
nor U7600 (N_7600,N_2591,N_1195);
nor U7601 (N_7601,N_3091,N_4265);
nand U7602 (N_7602,N_2903,N_926);
nor U7603 (N_7603,N_646,N_4154);
or U7604 (N_7604,N_641,N_920);
nand U7605 (N_7605,N_3499,N_3771);
and U7606 (N_7606,N_1934,N_2621);
and U7607 (N_7607,N_4091,N_1467);
nor U7608 (N_7608,N_1485,N_1408);
and U7609 (N_7609,N_3143,N_4738);
nor U7610 (N_7610,N_412,N_2402);
nor U7611 (N_7611,N_698,N_35);
or U7612 (N_7612,N_1807,N_1015);
nand U7613 (N_7613,N_2380,N_489);
and U7614 (N_7614,N_2724,N_1339);
nor U7615 (N_7615,N_657,N_756);
nor U7616 (N_7616,N_2755,N_2567);
or U7617 (N_7617,N_791,N_969);
nand U7618 (N_7618,N_378,N_1645);
nand U7619 (N_7619,N_2441,N_1540);
nor U7620 (N_7620,N_4373,N_2672);
nor U7621 (N_7621,N_3681,N_1401);
xnor U7622 (N_7622,N_3199,N_3406);
and U7623 (N_7623,N_1854,N_4158);
nor U7624 (N_7624,N_2335,N_3612);
or U7625 (N_7625,N_1043,N_1837);
and U7626 (N_7626,N_3377,N_1675);
xnor U7627 (N_7627,N_1899,N_2377);
nand U7628 (N_7628,N_3766,N_672);
or U7629 (N_7629,N_1480,N_1859);
and U7630 (N_7630,N_415,N_748);
nor U7631 (N_7631,N_53,N_128);
and U7632 (N_7632,N_887,N_2174);
nor U7633 (N_7633,N_4456,N_3939);
nand U7634 (N_7634,N_429,N_941);
or U7635 (N_7635,N_2785,N_217);
or U7636 (N_7636,N_1980,N_4846);
nand U7637 (N_7637,N_1076,N_744);
nor U7638 (N_7638,N_4594,N_549);
and U7639 (N_7639,N_3894,N_4858);
nand U7640 (N_7640,N_4730,N_4142);
or U7641 (N_7641,N_3762,N_4941);
and U7642 (N_7642,N_4,N_943);
nor U7643 (N_7643,N_2575,N_2362);
and U7644 (N_7644,N_2387,N_2163);
or U7645 (N_7645,N_71,N_2539);
and U7646 (N_7646,N_453,N_2006);
xor U7647 (N_7647,N_3361,N_1804);
nor U7648 (N_7648,N_4657,N_318);
or U7649 (N_7649,N_1279,N_2035);
nand U7650 (N_7650,N_3989,N_1473);
nand U7651 (N_7651,N_2984,N_1192);
nor U7652 (N_7652,N_925,N_4749);
xor U7653 (N_7653,N_2153,N_3724);
nor U7654 (N_7654,N_549,N_765);
nor U7655 (N_7655,N_3789,N_3336);
or U7656 (N_7656,N_120,N_1392);
nand U7657 (N_7657,N_4903,N_1941);
nor U7658 (N_7658,N_3075,N_2506);
or U7659 (N_7659,N_664,N_2647);
or U7660 (N_7660,N_1003,N_1034);
or U7661 (N_7661,N_176,N_1405);
or U7662 (N_7662,N_3065,N_995);
and U7663 (N_7663,N_435,N_1260);
xor U7664 (N_7664,N_985,N_3672);
or U7665 (N_7665,N_1610,N_4142);
nand U7666 (N_7666,N_2454,N_3034);
or U7667 (N_7667,N_1735,N_3143);
or U7668 (N_7668,N_457,N_1176);
and U7669 (N_7669,N_3583,N_4008);
nor U7670 (N_7670,N_1555,N_4367);
nor U7671 (N_7671,N_1831,N_3716);
nor U7672 (N_7672,N_4727,N_3833);
or U7673 (N_7673,N_563,N_918);
nor U7674 (N_7674,N_3247,N_4186);
or U7675 (N_7675,N_892,N_276);
and U7676 (N_7676,N_4159,N_2867);
or U7677 (N_7677,N_2708,N_980);
and U7678 (N_7678,N_3184,N_4752);
or U7679 (N_7679,N_4206,N_2351);
nor U7680 (N_7680,N_34,N_1844);
nand U7681 (N_7681,N_4494,N_2688);
nor U7682 (N_7682,N_2469,N_3189);
nor U7683 (N_7683,N_1147,N_2058);
or U7684 (N_7684,N_189,N_1449);
nand U7685 (N_7685,N_2317,N_589);
and U7686 (N_7686,N_1198,N_1227);
nand U7687 (N_7687,N_2877,N_4631);
or U7688 (N_7688,N_2643,N_459);
nand U7689 (N_7689,N_4532,N_841);
or U7690 (N_7690,N_690,N_1679);
xor U7691 (N_7691,N_3219,N_1419);
xor U7692 (N_7692,N_4046,N_2359);
and U7693 (N_7693,N_4895,N_1294);
or U7694 (N_7694,N_522,N_4450);
or U7695 (N_7695,N_831,N_4486);
or U7696 (N_7696,N_392,N_3073);
nand U7697 (N_7697,N_2402,N_1568);
xor U7698 (N_7698,N_3094,N_4709);
and U7699 (N_7699,N_2376,N_2028);
and U7700 (N_7700,N_2778,N_833);
nor U7701 (N_7701,N_4527,N_2555);
nor U7702 (N_7702,N_2100,N_220);
nand U7703 (N_7703,N_1831,N_3311);
xor U7704 (N_7704,N_3426,N_3535);
nor U7705 (N_7705,N_3109,N_2472);
and U7706 (N_7706,N_2335,N_3143);
and U7707 (N_7707,N_2458,N_3141);
nor U7708 (N_7708,N_4177,N_904);
and U7709 (N_7709,N_4118,N_880);
and U7710 (N_7710,N_1569,N_3210);
and U7711 (N_7711,N_3866,N_623);
nor U7712 (N_7712,N_922,N_3632);
and U7713 (N_7713,N_3510,N_3927);
nor U7714 (N_7714,N_4795,N_370);
nand U7715 (N_7715,N_1762,N_2226);
nor U7716 (N_7716,N_2081,N_2343);
and U7717 (N_7717,N_4769,N_1331);
nor U7718 (N_7718,N_4310,N_2492);
xnor U7719 (N_7719,N_2730,N_1055);
and U7720 (N_7720,N_3861,N_2718);
and U7721 (N_7721,N_4336,N_2902);
and U7722 (N_7722,N_925,N_4888);
or U7723 (N_7723,N_4235,N_859);
or U7724 (N_7724,N_4231,N_779);
nand U7725 (N_7725,N_265,N_4511);
nor U7726 (N_7726,N_4967,N_4524);
or U7727 (N_7727,N_187,N_1550);
nor U7728 (N_7728,N_3650,N_1235);
and U7729 (N_7729,N_1062,N_1267);
nand U7730 (N_7730,N_1291,N_2974);
or U7731 (N_7731,N_1518,N_2480);
nor U7732 (N_7732,N_3800,N_1058);
nand U7733 (N_7733,N_616,N_4664);
or U7734 (N_7734,N_4088,N_2297);
or U7735 (N_7735,N_1370,N_3803);
and U7736 (N_7736,N_3368,N_468);
or U7737 (N_7737,N_1131,N_4064);
and U7738 (N_7738,N_1317,N_1953);
nor U7739 (N_7739,N_2005,N_647);
xor U7740 (N_7740,N_1512,N_1445);
and U7741 (N_7741,N_4047,N_4079);
xor U7742 (N_7742,N_3758,N_2426);
nor U7743 (N_7743,N_4490,N_17);
nand U7744 (N_7744,N_4183,N_3746);
nand U7745 (N_7745,N_4057,N_4962);
nor U7746 (N_7746,N_3065,N_903);
nand U7747 (N_7747,N_3128,N_4193);
and U7748 (N_7748,N_1191,N_1269);
nand U7749 (N_7749,N_1737,N_4631);
and U7750 (N_7750,N_2596,N_4250);
and U7751 (N_7751,N_3345,N_3096);
nor U7752 (N_7752,N_2385,N_1573);
nor U7753 (N_7753,N_4276,N_116);
xnor U7754 (N_7754,N_2553,N_4358);
and U7755 (N_7755,N_1041,N_2850);
and U7756 (N_7756,N_2159,N_2415);
nand U7757 (N_7757,N_229,N_1264);
nor U7758 (N_7758,N_1645,N_4216);
or U7759 (N_7759,N_3521,N_2595);
nor U7760 (N_7760,N_2731,N_3648);
nand U7761 (N_7761,N_420,N_951);
or U7762 (N_7762,N_2093,N_2357);
or U7763 (N_7763,N_1104,N_630);
nand U7764 (N_7764,N_4192,N_1092);
and U7765 (N_7765,N_4176,N_1347);
and U7766 (N_7766,N_2917,N_2605);
nand U7767 (N_7767,N_3450,N_102);
nor U7768 (N_7768,N_4626,N_1641);
nor U7769 (N_7769,N_4435,N_4762);
or U7770 (N_7770,N_4256,N_2407);
and U7771 (N_7771,N_4540,N_3793);
nand U7772 (N_7772,N_206,N_3336);
or U7773 (N_7773,N_362,N_2364);
nand U7774 (N_7774,N_4178,N_3379);
or U7775 (N_7775,N_3347,N_3910);
and U7776 (N_7776,N_3655,N_2134);
and U7777 (N_7777,N_4934,N_1271);
xnor U7778 (N_7778,N_1199,N_1201);
or U7779 (N_7779,N_4047,N_3739);
or U7780 (N_7780,N_3910,N_2932);
nand U7781 (N_7781,N_4305,N_2773);
or U7782 (N_7782,N_1785,N_2855);
nor U7783 (N_7783,N_261,N_526);
or U7784 (N_7784,N_4385,N_2947);
nor U7785 (N_7785,N_1149,N_3913);
and U7786 (N_7786,N_2197,N_3844);
xnor U7787 (N_7787,N_3248,N_270);
nand U7788 (N_7788,N_2113,N_3938);
nand U7789 (N_7789,N_4325,N_4879);
and U7790 (N_7790,N_3505,N_4593);
and U7791 (N_7791,N_1635,N_1577);
nor U7792 (N_7792,N_4442,N_2371);
or U7793 (N_7793,N_4990,N_4219);
and U7794 (N_7794,N_896,N_3611);
nand U7795 (N_7795,N_4940,N_4167);
nand U7796 (N_7796,N_2722,N_3103);
nor U7797 (N_7797,N_1468,N_3133);
or U7798 (N_7798,N_4853,N_2078);
or U7799 (N_7799,N_285,N_205);
nor U7800 (N_7800,N_587,N_839);
and U7801 (N_7801,N_4600,N_2268);
xnor U7802 (N_7802,N_2027,N_2492);
or U7803 (N_7803,N_1817,N_3596);
nand U7804 (N_7804,N_1755,N_3795);
xnor U7805 (N_7805,N_1789,N_2353);
or U7806 (N_7806,N_1437,N_3430);
and U7807 (N_7807,N_700,N_1122);
and U7808 (N_7808,N_1403,N_2404);
and U7809 (N_7809,N_2278,N_3245);
xnor U7810 (N_7810,N_3562,N_3785);
and U7811 (N_7811,N_2566,N_3564);
nor U7812 (N_7812,N_1125,N_3757);
nor U7813 (N_7813,N_1643,N_71);
nand U7814 (N_7814,N_4939,N_1755);
nand U7815 (N_7815,N_3899,N_3051);
nand U7816 (N_7816,N_1050,N_214);
xnor U7817 (N_7817,N_4606,N_1486);
nand U7818 (N_7818,N_4265,N_3829);
nand U7819 (N_7819,N_2305,N_2898);
and U7820 (N_7820,N_3402,N_4294);
nand U7821 (N_7821,N_1007,N_3515);
and U7822 (N_7822,N_2493,N_2247);
xor U7823 (N_7823,N_2784,N_3356);
nand U7824 (N_7824,N_4808,N_1211);
nor U7825 (N_7825,N_890,N_3492);
nor U7826 (N_7826,N_4810,N_1332);
nand U7827 (N_7827,N_128,N_3535);
xnor U7828 (N_7828,N_3998,N_1259);
or U7829 (N_7829,N_2823,N_1979);
and U7830 (N_7830,N_3001,N_2446);
nor U7831 (N_7831,N_1040,N_3066);
and U7832 (N_7832,N_4518,N_4176);
or U7833 (N_7833,N_2339,N_268);
nor U7834 (N_7834,N_2847,N_582);
and U7835 (N_7835,N_1447,N_4850);
and U7836 (N_7836,N_4617,N_4548);
or U7837 (N_7837,N_1215,N_2740);
xor U7838 (N_7838,N_3796,N_1480);
or U7839 (N_7839,N_3326,N_2549);
or U7840 (N_7840,N_198,N_1932);
or U7841 (N_7841,N_48,N_865);
nor U7842 (N_7842,N_4154,N_3168);
or U7843 (N_7843,N_3537,N_1233);
and U7844 (N_7844,N_206,N_181);
or U7845 (N_7845,N_2365,N_2355);
nand U7846 (N_7846,N_3,N_769);
nand U7847 (N_7847,N_1885,N_3471);
nor U7848 (N_7848,N_1201,N_2873);
nand U7849 (N_7849,N_4705,N_3076);
nor U7850 (N_7850,N_225,N_4009);
nor U7851 (N_7851,N_2572,N_3945);
and U7852 (N_7852,N_2230,N_3704);
nor U7853 (N_7853,N_2465,N_2457);
and U7854 (N_7854,N_1220,N_4108);
nand U7855 (N_7855,N_1987,N_2641);
and U7856 (N_7856,N_4403,N_4027);
nand U7857 (N_7857,N_3365,N_4649);
or U7858 (N_7858,N_837,N_1593);
nand U7859 (N_7859,N_779,N_3875);
and U7860 (N_7860,N_3020,N_1081);
or U7861 (N_7861,N_4026,N_3456);
nor U7862 (N_7862,N_3756,N_2701);
and U7863 (N_7863,N_1754,N_401);
or U7864 (N_7864,N_1855,N_988);
or U7865 (N_7865,N_2478,N_42);
or U7866 (N_7866,N_45,N_168);
and U7867 (N_7867,N_2385,N_4012);
or U7868 (N_7868,N_1338,N_4127);
or U7869 (N_7869,N_4642,N_3069);
nor U7870 (N_7870,N_1943,N_4032);
and U7871 (N_7871,N_1342,N_97);
and U7872 (N_7872,N_3008,N_1555);
nor U7873 (N_7873,N_661,N_3765);
or U7874 (N_7874,N_4405,N_39);
nor U7875 (N_7875,N_2932,N_4909);
and U7876 (N_7876,N_4352,N_3083);
or U7877 (N_7877,N_1237,N_3636);
nor U7878 (N_7878,N_1512,N_2425);
nand U7879 (N_7879,N_4031,N_3143);
nand U7880 (N_7880,N_4724,N_2824);
nor U7881 (N_7881,N_2342,N_4419);
nand U7882 (N_7882,N_693,N_1628);
nand U7883 (N_7883,N_3006,N_645);
xor U7884 (N_7884,N_2333,N_3253);
nand U7885 (N_7885,N_1006,N_1557);
nand U7886 (N_7886,N_3340,N_3419);
or U7887 (N_7887,N_1984,N_4690);
nand U7888 (N_7888,N_3946,N_3835);
nand U7889 (N_7889,N_2145,N_1423);
and U7890 (N_7890,N_2381,N_2362);
and U7891 (N_7891,N_3062,N_3360);
and U7892 (N_7892,N_3508,N_3547);
nand U7893 (N_7893,N_3725,N_521);
and U7894 (N_7894,N_15,N_2029);
and U7895 (N_7895,N_783,N_2069);
nor U7896 (N_7896,N_4696,N_2707);
nor U7897 (N_7897,N_2907,N_3044);
and U7898 (N_7898,N_4492,N_3325);
or U7899 (N_7899,N_2983,N_2104);
xnor U7900 (N_7900,N_2223,N_3486);
nor U7901 (N_7901,N_142,N_38);
nor U7902 (N_7902,N_1099,N_2089);
and U7903 (N_7903,N_4727,N_2629);
or U7904 (N_7904,N_1079,N_1161);
nor U7905 (N_7905,N_4386,N_2283);
nor U7906 (N_7906,N_3026,N_632);
nor U7907 (N_7907,N_288,N_1417);
or U7908 (N_7908,N_3525,N_3927);
and U7909 (N_7909,N_2998,N_2085);
or U7910 (N_7910,N_1033,N_2989);
or U7911 (N_7911,N_4130,N_3762);
nor U7912 (N_7912,N_522,N_2674);
xnor U7913 (N_7913,N_466,N_2402);
nand U7914 (N_7914,N_3172,N_2464);
or U7915 (N_7915,N_4885,N_2934);
xor U7916 (N_7916,N_723,N_3988);
or U7917 (N_7917,N_4036,N_169);
xnor U7918 (N_7918,N_3709,N_410);
nor U7919 (N_7919,N_3193,N_671);
xor U7920 (N_7920,N_3702,N_220);
and U7921 (N_7921,N_1831,N_1948);
and U7922 (N_7922,N_1208,N_3290);
nand U7923 (N_7923,N_1032,N_2868);
or U7924 (N_7924,N_2384,N_1319);
nand U7925 (N_7925,N_2557,N_428);
nor U7926 (N_7926,N_1789,N_610);
xor U7927 (N_7927,N_1040,N_3639);
nor U7928 (N_7928,N_1571,N_4419);
nor U7929 (N_7929,N_4302,N_4629);
and U7930 (N_7930,N_117,N_1510);
xor U7931 (N_7931,N_3769,N_4395);
and U7932 (N_7932,N_2173,N_586);
xor U7933 (N_7933,N_220,N_4650);
nand U7934 (N_7934,N_1022,N_3758);
or U7935 (N_7935,N_4867,N_3673);
or U7936 (N_7936,N_4298,N_4326);
nor U7937 (N_7937,N_4476,N_4960);
nor U7938 (N_7938,N_2477,N_2568);
nor U7939 (N_7939,N_1230,N_4352);
and U7940 (N_7940,N_2909,N_1147);
and U7941 (N_7941,N_2750,N_1462);
nor U7942 (N_7942,N_4279,N_1912);
and U7943 (N_7943,N_1612,N_3314);
nor U7944 (N_7944,N_3354,N_1852);
and U7945 (N_7945,N_2352,N_3911);
nor U7946 (N_7946,N_2173,N_1865);
or U7947 (N_7947,N_3563,N_1482);
nand U7948 (N_7948,N_3939,N_4321);
and U7949 (N_7949,N_4409,N_2767);
or U7950 (N_7950,N_3075,N_1214);
and U7951 (N_7951,N_2860,N_140);
xnor U7952 (N_7952,N_1013,N_3272);
nand U7953 (N_7953,N_4985,N_2208);
nand U7954 (N_7954,N_4980,N_1488);
nand U7955 (N_7955,N_3210,N_665);
or U7956 (N_7956,N_2843,N_3222);
xnor U7957 (N_7957,N_4589,N_3255);
and U7958 (N_7958,N_762,N_1586);
xnor U7959 (N_7959,N_2213,N_3588);
or U7960 (N_7960,N_4073,N_774);
nor U7961 (N_7961,N_3573,N_2043);
nor U7962 (N_7962,N_4087,N_3653);
nor U7963 (N_7963,N_1649,N_4049);
or U7964 (N_7964,N_4299,N_198);
xnor U7965 (N_7965,N_4157,N_1006);
or U7966 (N_7966,N_3021,N_3346);
nand U7967 (N_7967,N_347,N_773);
nand U7968 (N_7968,N_2255,N_2163);
and U7969 (N_7969,N_1682,N_49);
nand U7970 (N_7970,N_2318,N_4466);
nand U7971 (N_7971,N_4874,N_4768);
or U7972 (N_7972,N_2371,N_4741);
and U7973 (N_7973,N_4707,N_4580);
nor U7974 (N_7974,N_922,N_1695);
or U7975 (N_7975,N_4385,N_493);
xor U7976 (N_7976,N_1803,N_4980);
xor U7977 (N_7977,N_3815,N_4776);
and U7978 (N_7978,N_2048,N_4638);
nand U7979 (N_7979,N_3789,N_2237);
nor U7980 (N_7980,N_2054,N_3598);
nor U7981 (N_7981,N_2568,N_251);
and U7982 (N_7982,N_3598,N_2407);
nor U7983 (N_7983,N_2383,N_1054);
nor U7984 (N_7984,N_4714,N_4257);
or U7985 (N_7985,N_1007,N_1122);
nand U7986 (N_7986,N_3464,N_736);
nand U7987 (N_7987,N_1565,N_482);
nor U7988 (N_7988,N_1186,N_159);
nor U7989 (N_7989,N_4907,N_3041);
nand U7990 (N_7990,N_1317,N_3393);
or U7991 (N_7991,N_3941,N_604);
nand U7992 (N_7992,N_2737,N_3872);
nor U7993 (N_7993,N_4148,N_424);
nand U7994 (N_7994,N_2871,N_2862);
and U7995 (N_7995,N_3656,N_3727);
and U7996 (N_7996,N_3075,N_1491);
and U7997 (N_7997,N_936,N_222);
xor U7998 (N_7998,N_4793,N_3024);
nor U7999 (N_7999,N_4631,N_3242);
nor U8000 (N_8000,N_1290,N_3213);
and U8001 (N_8001,N_664,N_1986);
nand U8002 (N_8002,N_4110,N_782);
xor U8003 (N_8003,N_2635,N_4974);
nor U8004 (N_8004,N_1270,N_3103);
or U8005 (N_8005,N_1906,N_1892);
nand U8006 (N_8006,N_4921,N_1227);
or U8007 (N_8007,N_1512,N_798);
and U8008 (N_8008,N_125,N_2419);
nand U8009 (N_8009,N_1605,N_3586);
nor U8010 (N_8010,N_1070,N_1337);
nand U8011 (N_8011,N_384,N_4788);
nor U8012 (N_8012,N_849,N_4003);
nand U8013 (N_8013,N_2279,N_1380);
nand U8014 (N_8014,N_3992,N_569);
nor U8015 (N_8015,N_4100,N_753);
nand U8016 (N_8016,N_242,N_1717);
nand U8017 (N_8017,N_2993,N_2652);
nand U8018 (N_8018,N_2723,N_4335);
and U8019 (N_8019,N_648,N_2358);
or U8020 (N_8020,N_1981,N_2151);
nand U8021 (N_8021,N_4730,N_1027);
and U8022 (N_8022,N_3083,N_4389);
nor U8023 (N_8023,N_3698,N_2225);
and U8024 (N_8024,N_3353,N_1983);
xnor U8025 (N_8025,N_1511,N_3072);
xnor U8026 (N_8026,N_1965,N_206);
or U8027 (N_8027,N_4576,N_1214);
nand U8028 (N_8028,N_499,N_1740);
xor U8029 (N_8029,N_458,N_3094);
or U8030 (N_8030,N_4154,N_43);
nand U8031 (N_8031,N_501,N_2235);
or U8032 (N_8032,N_1171,N_4915);
and U8033 (N_8033,N_816,N_1337);
nand U8034 (N_8034,N_1188,N_3607);
nand U8035 (N_8035,N_4437,N_4617);
or U8036 (N_8036,N_2874,N_2054);
nor U8037 (N_8037,N_3586,N_4492);
nand U8038 (N_8038,N_1954,N_4754);
nor U8039 (N_8039,N_729,N_4303);
nor U8040 (N_8040,N_131,N_2816);
nand U8041 (N_8041,N_3099,N_181);
and U8042 (N_8042,N_1469,N_2405);
nor U8043 (N_8043,N_3596,N_1232);
nor U8044 (N_8044,N_4920,N_1604);
or U8045 (N_8045,N_4868,N_198);
nand U8046 (N_8046,N_2024,N_2364);
and U8047 (N_8047,N_3407,N_565);
nand U8048 (N_8048,N_2477,N_3863);
or U8049 (N_8049,N_349,N_3656);
and U8050 (N_8050,N_785,N_4523);
nor U8051 (N_8051,N_2738,N_4820);
nand U8052 (N_8052,N_3101,N_534);
and U8053 (N_8053,N_543,N_2454);
xnor U8054 (N_8054,N_2492,N_1409);
or U8055 (N_8055,N_3125,N_134);
or U8056 (N_8056,N_415,N_2162);
and U8057 (N_8057,N_4183,N_3295);
nand U8058 (N_8058,N_1599,N_4494);
or U8059 (N_8059,N_4604,N_3619);
nand U8060 (N_8060,N_2577,N_3978);
nand U8061 (N_8061,N_4766,N_2734);
and U8062 (N_8062,N_4583,N_392);
nand U8063 (N_8063,N_2023,N_2655);
nor U8064 (N_8064,N_2189,N_2956);
and U8065 (N_8065,N_2250,N_4913);
and U8066 (N_8066,N_2963,N_4397);
nand U8067 (N_8067,N_4482,N_1848);
or U8068 (N_8068,N_3188,N_3602);
nand U8069 (N_8069,N_1259,N_1076);
nand U8070 (N_8070,N_3718,N_2784);
nor U8071 (N_8071,N_596,N_2788);
and U8072 (N_8072,N_4325,N_2574);
and U8073 (N_8073,N_3961,N_2897);
and U8074 (N_8074,N_2174,N_975);
xnor U8075 (N_8075,N_2092,N_1773);
and U8076 (N_8076,N_1545,N_2798);
and U8077 (N_8077,N_1325,N_1373);
xor U8078 (N_8078,N_1600,N_1344);
or U8079 (N_8079,N_1777,N_4893);
or U8080 (N_8080,N_69,N_213);
and U8081 (N_8081,N_4223,N_878);
and U8082 (N_8082,N_428,N_3008);
or U8083 (N_8083,N_2329,N_555);
and U8084 (N_8084,N_4928,N_3350);
nor U8085 (N_8085,N_4631,N_862);
or U8086 (N_8086,N_4844,N_2734);
nor U8087 (N_8087,N_1136,N_4549);
or U8088 (N_8088,N_1483,N_1894);
nand U8089 (N_8089,N_4501,N_460);
nor U8090 (N_8090,N_3172,N_3258);
and U8091 (N_8091,N_1999,N_3433);
and U8092 (N_8092,N_74,N_388);
and U8093 (N_8093,N_4983,N_738);
nand U8094 (N_8094,N_4024,N_2365);
or U8095 (N_8095,N_1702,N_450);
and U8096 (N_8096,N_1388,N_3157);
xnor U8097 (N_8097,N_43,N_640);
nor U8098 (N_8098,N_981,N_4121);
nand U8099 (N_8099,N_1188,N_2507);
nor U8100 (N_8100,N_1964,N_440);
nand U8101 (N_8101,N_1622,N_3786);
or U8102 (N_8102,N_723,N_2203);
and U8103 (N_8103,N_2192,N_3450);
nor U8104 (N_8104,N_4363,N_1036);
or U8105 (N_8105,N_3285,N_4362);
or U8106 (N_8106,N_992,N_3398);
nor U8107 (N_8107,N_3459,N_2540);
and U8108 (N_8108,N_146,N_4342);
xnor U8109 (N_8109,N_4105,N_1853);
nor U8110 (N_8110,N_1846,N_270);
nand U8111 (N_8111,N_1608,N_622);
and U8112 (N_8112,N_2870,N_173);
and U8113 (N_8113,N_4453,N_1353);
xor U8114 (N_8114,N_2656,N_4455);
nor U8115 (N_8115,N_4323,N_4833);
and U8116 (N_8116,N_2835,N_291);
nand U8117 (N_8117,N_1719,N_2739);
nor U8118 (N_8118,N_4642,N_4182);
nor U8119 (N_8119,N_4415,N_2569);
nand U8120 (N_8120,N_2373,N_3797);
nor U8121 (N_8121,N_1769,N_3214);
nor U8122 (N_8122,N_3612,N_2442);
nor U8123 (N_8123,N_1586,N_3765);
nor U8124 (N_8124,N_174,N_392);
or U8125 (N_8125,N_3837,N_2084);
nor U8126 (N_8126,N_4385,N_2493);
and U8127 (N_8127,N_4518,N_4703);
or U8128 (N_8128,N_1022,N_421);
and U8129 (N_8129,N_3832,N_4853);
xnor U8130 (N_8130,N_3709,N_2212);
nand U8131 (N_8131,N_3832,N_78);
or U8132 (N_8132,N_121,N_3615);
xnor U8133 (N_8133,N_2957,N_4765);
nor U8134 (N_8134,N_2423,N_3161);
nor U8135 (N_8135,N_826,N_1307);
xnor U8136 (N_8136,N_967,N_1406);
nor U8137 (N_8137,N_3044,N_4334);
or U8138 (N_8138,N_1784,N_2269);
nand U8139 (N_8139,N_3537,N_1951);
nor U8140 (N_8140,N_4591,N_4370);
or U8141 (N_8141,N_4839,N_4933);
or U8142 (N_8142,N_982,N_412);
or U8143 (N_8143,N_994,N_267);
and U8144 (N_8144,N_4366,N_3550);
nand U8145 (N_8145,N_2248,N_4950);
nand U8146 (N_8146,N_3782,N_4658);
nand U8147 (N_8147,N_1089,N_2999);
or U8148 (N_8148,N_4084,N_2213);
and U8149 (N_8149,N_2678,N_2333);
and U8150 (N_8150,N_2170,N_1056);
nor U8151 (N_8151,N_1041,N_1976);
and U8152 (N_8152,N_1055,N_3647);
and U8153 (N_8153,N_4794,N_3155);
nor U8154 (N_8154,N_4589,N_1230);
or U8155 (N_8155,N_4557,N_2300);
nand U8156 (N_8156,N_1043,N_544);
and U8157 (N_8157,N_781,N_247);
xnor U8158 (N_8158,N_210,N_980);
nand U8159 (N_8159,N_2871,N_3318);
nor U8160 (N_8160,N_1330,N_4949);
nor U8161 (N_8161,N_912,N_1298);
or U8162 (N_8162,N_1889,N_2131);
nand U8163 (N_8163,N_759,N_2518);
nand U8164 (N_8164,N_1336,N_3788);
and U8165 (N_8165,N_1019,N_2299);
nand U8166 (N_8166,N_3824,N_4725);
or U8167 (N_8167,N_4518,N_2088);
nor U8168 (N_8168,N_4336,N_4988);
and U8169 (N_8169,N_646,N_523);
and U8170 (N_8170,N_3315,N_4862);
nand U8171 (N_8171,N_1178,N_1986);
nand U8172 (N_8172,N_3572,N_2354);
nor U8173 (N_8173,N_3970,N_590);
and U8174 (N_8174,N_2857,N_1761);
or U8175 (N_8175,N_3430,N_278);
and U8176 (N_8176,N_4047,N_4400);
nand U8177 (N_8177,N_2264,N_1508);
nand U8178 (N_8178,N_2183,N_1124);
nand U8179 (N_8179,N_165,N_331);
xor U8180 (N_8180,N_3625,N_3631);
nand U8181 (N_8181,N_2504,N_4841);
nand U8182 (N_8182,N_984,N_450);
nor U8183 (N_8183,N_496,N_4752);
nand U8184 (N_8184,N_1717,N_3355);
or U8185 (N_8185,N_2205,N_2931);
or U8186 (N_8186,N_4351,N_348);
nand U8187 (N_8187,N_1932,N_825);
xor U8188 (N_8188,N_2895,N_2974);
xor U8189 (N_8189,N_3089,N_4026);
and U8190 (N_8190,N_3058,N_2539);
or U8191 (N_8191,N_4713,N_3322);
or U8192 (N_8192,N_1155,N_2434);
nor U8193 (N_8193,N_4075,N_3488);
nor U8194 (N_8194,N_1369,N_4135);
and U8195 (N_8195,N_1231,N_3994);
or U8196 (N_8196,N_3285,N_4541);
or U8197 (N_8197,N_4889,N_3222);
nor U8198 (N_8198,N_2470,N_4202);
or U8199 (N_8199,N_1358,N_2405);
and U8200 (N_8200,N_1790,N_4461);
nor U8201 (N_8201,N_2933,N_1978);
and U8202 (N_8202,N_1862,N_3900);
nor U8203 (N_8203,N_1498,N_1375);
or U8204 (N_8204,N_1938,N_3646);
nand U8205 (N_8205,N_572,N_4206);
nand U8206 (N_8206,N_530,N_2070);
nor U8207 (N_8207,N_3742,N_1716);
and U8208 (N_8208,N_2517,N_2133);
or U8209 (N_8209,N_250,N_3397);
nand U8210 (N_8210,N_4838,N_3675);
nor U8211 (N_8211,N_687,N_3214);
nor U8212 (N_8212,N_3970,N_2198);
or U8213 (N_8213,N_2185,N_1260);
nor U8214 (N_8214,N_855,N_190);
and U8215 (N_8215,N_49,N_2624);
and U8216 (N_8216,N_2512,N_4420);
and U8217 (N_8217,N_2533,N_1981);
and U8218 (N_8218,N_1547,N_4959);
or U8219 (N_8219,N_4692,N_4392);
nor U8220 (N_8220,N_4777,N_2882);
nor U8221 (N_8221,N_3728,N_4616);
and U8222 (N_8222,N_4167,N_2724);
nor U8223 (N_8223,N_1046,N_1829);
and U8224 (N_8224,N_3193,N_579);
nand U8225 (N_8225,N_3658,N_1038);
nor U8226 (N_8226,N_309,N_752);
nor U8227 (N_8227,N_809,N_3631);
or U8228 (N_8228,N_838,N_4923);
nor U8229 (N_8229,N_1900,N_1846);
and U8230 (N_8230,N_4232,N_2504);
or U8231 (N_8231,N_4145,N_4180);
nand U8232 (N_8232,N_4434,N_3974);
nand U8233 (N_8233,N_1922,N_2570);
nor U8234 (N_8234,N_1889,N_4236);
or U8235 (N_8235,N_2688,N_3231);
and U8236 (N_8236,N_3861,N_3740);
and U8237 (N_8237,N_3993,N_2828);
xor U8238 (N_8238,N_4219,N_1148);
nand U8239 (N_8239,N_2379,N_842);
nor U8240 (N_8240,N_4393,N_2577);
nand U8241 (N_8241,N_3623,N_1116);
or U8242 (N_8242,N_2803,N_4467);
or U8243 (N_8243,N_3420,N_3930);
nor U8244 (N_8244,N_4170,N_338);
nor U8245 (N_8245,N_4300,N_2709);
nor U8246 (N_8246,N_1995,N_908);
nand U8247 (N_8247,N_4144,N_2950);
nor U8248 (N_8248,N_4844,N_4740);
and U8249 (N_8249,N_410,N_4026);
and U8250 (N_8250,N_4450,N_2722);
or U8251 (N_8251,N_3518,N_2272);
nand U8252 (N_8252,N_2411,N_242);
xor U8253 (N_8253,N_4555,N_775);
nor U8254 (N_8254,N_2136,N_3109);
nor U8255 (N_8255,N_3384,N_4601);
nand U8256 (N_8256,N_2419,N_2071);
xnor U8257 (N_8257,N_1568,N_1394);
nand U8258 (N_8258,N_2489,N_2263);
nand U8259 (N_8259,N_2820,N_947);
or U8260 (N_8260,N_1886,N_1600);
nand U8261 (N_8261,N_1413,N_2469);
and U8262 (N_8262,N_3746,N_3350);
and U8263 (N_8263,N_2284,N_2214);
nor U8264 (N_8264,N_778,N_4793);
or U8265 (N_8265,N_502,N_2676);
and U8266 (N_8266,N_3420,N_4930);
nor U8267 (N_8267,N_70,N_732);
xnor U8268 (N_8268,N_2303,N_4189);
or U8269 (N_8269,N_2657,N_4165);
and U8270 (N_8270,N_3581,N_1353);
and U8271 (N_8271,N_3056,N_1281);
or U8272 (N_8272,N_504,N_3733);
xnor U8273 (N_8273,N_3218,N_305);
or U8274 (N_8274,N_2961,N_1961);
nor U8275 (N_8275,N_2534,N_4617);
and U8276 (N_8276,N_322,N_1418);
nand U8277 (N_8277,N_4347,N_0);
or U8278 (N_8278,N_3238,N_4622);
nor U8279 (N_8279,N_1252,N_2182);
xnor U8280 (N_8280,N_4345,N_4445);
and U8281 (N_8281,N_256,N_3068);
xor U8282 (N_8282,N_2253,N_3937);
xnor U8283 (N_8283,N_3020,N_1545);
nor U8284 (N_8284,N_4140,N_1618);
nor U8285 (N_8285,N_4810,N_4482);
or U8286 (N_8286,N_4743,N_1173);
and U8287 (N_8287,N_2971,N_4322);
or U8288 (N_8288,N_3598,N_535);
and U8289 (N_8289,N_1166,N_4682);
nor U8290 (N_8290,N_4726,N_1850);
or U8291 (N_8291,N_4230,N_1878);
nand U8292 (N_8292,N_380,N_1118);
nand U8293 (N_8293,N_1224,N_4455);
and U8294 (N_8294,N_3970,N_2618);
nor U8295 (N_8295,N_74,N_152);
or U8296 (N_8296,N_4467,N_482);
xor U8297 (N_8297,N_1973,N_170);
nand U8298 (N_8298,N_2437,N_4179);
and U8299 (N_8299,N_2774,N_4715);
or U8300 (N_8300,N_1406,N_629);
nor U8301 (N_8301,N_4582,N_1489);
and U8302 (N_8302,N_3022,N_3057);
or U8303 (N_8303,N_3283,N_2761);
nor U8304 (N_8304,N_1677,N_3736);
nor U8305 (N_8305,N_4387,N_3829);
or U8306 (N_8306,N_3268,N_842);
nor U8307 (N_8307,N_2345,N_746);
xnor U8308 (N_8308,N_602,N_153);
xor U8309 (N_8309,N_3129,N_995);
or U8310 (N_8310,N_392,N_3343);
nand U8311 (N_8311,N_3048,N_4452);
or U8312 (N_8312,N_4243,N_4293);
or U8313 (N_8313,N_3647,N_923);
and U8314 (N_8314,N_2311,N_2577);
xnor U8315 (N_8315,N_2395,N_4264);
nand U8316 (N_8316,N_1298,N_3808);
and U8317 (N_8317,N_2850,N_1170);
nor U8318 (N_8318,N_3658,N_3866);
xnor U8319 (N_8319,N_2922,N_4856);
nand U8320 (N_8320,N_2671,N_4616);
or U8321 (N_8321,N_4673,N_3742);
xor U8322 (N_8322,N_728,N_2511);
nand U8323 (N_8323,N_161,N_4279);
or U8324 (N_8324,N_2230,N_3295);
and U8325 (N_8325,N_4176,N_2900);
xnor U8326 (N_8326,N_4047,N_608);
or U8327 (N_8327,N_4198,N_2149);
and U8328 (N_8328,N_1954,N_3333);
nor U8329 (N_8329,N_3672,N_3206);
nand U8330 (N_8330,N_1517,N_1547);
and U8331 (N_8331,N_2929,N_2471);
nor U8332 (N_8332,N_1723,N_2685);
nor U8333 (N_8333,N_4306,N_1942);
nand U8334 (N_8334,N_717,N_4559);
nor U8335 (N_8335,N_505,N_2178);
xor U8336 (N_8336,N_2269,N_4944);
and U8337 (N_8337,N_2343,N_4988);
xor U8338 (N_8338,N_4125,N_4005);
nor U8339 (N_8339,N_4381,N_3816);
or U8340 (N_8340,N_1861,N_2224);
xor U8341 (N_8341,N_1781,N_3729);
or U8342 (N_8342,N_2505,N_2484);
nor U8343 (N_8343,N_430,N_37);
nor U8344 (N_8344,N_4597,N_137);
nand U8345 (N_8345,N_2086,N_2986);
nand U8346 (N_8346,N_4355,N_425);
nand U8347 (N_8347,N_3222,N_2370);
nor U8348 (N_8348,N_1195,N_1981);
nand U8349 (N_8349,N_1486,N_1542);
nor U8350 (N_8350,N_838,N_1630);
and U8351 (N_8351,N_1477,N_2671);
nand U8352 (N_8352,N_4066,N_2088);
and U8353 (N_8353,N_248,N_1565);
or U8354 (N_8354,N_2060,N_2186);
or U8355 (N_8355,N_4409,N_2812);
or U8356 (N_8356,N_2646,N_729);
or U8357 (N_8357,N_1832,N_4255);
or U8358 (N_8358,N_4768,N_4254);
nor U8359 (N_8359,N_4503,N_976);
or U8360 (N_8360,N_2555,N_1908);
or U8361 (N_8361,N_2848,N_1818);
or U8362 (N_8362,N_3513,N_361);
nor U8363 (N_8363,N_3998,N_3028);
and U8364 (N_8364,N_188,N_3074);
and U8365 (N_8365,N_4546,N_4405);
nand U8366 (N_8366,N_3512,N_4379);
nand U8367 (N_8367,N_214,N_1601);
nand U8368 (N_8368,N_1148,N_3578);
nor U8369 (N_8369,N_3692,N_3041);
nor U8370 (N_8370,N_8,N_2185);
nor U8371 (N_8371,N_847,N_4687);
xor U8372 (N_8372,N_3591,N_450);
or U8373 (N_8373,N_3462,N_2484);
or U8374 (N_8374,N_3515,N_3660);
and U8375 (N_8375,N_4562,N_3507);
or U8376 (N_8376,N_2496,N_563);
and U8377 (N_8377,N_3565,N_1815);
or U8378 (N_8378,N_4095,N_2240);
and U8379 (N_8379,N_3122,N_3398);
nor U8380 (N_8380,N_3461,N_2750);
nor U8381 (N_8381,N_448,N_1724);
and U8382 (N_8382,N_898,N_748);
nor U8383 (N_8383,N_1834,N_3495);
nand U8384 (N_8384,N_1478,N_2142);
and U8385 (N_8385,N_3738,N_4722);
and U8386 (N_8386,N_3071,N_4691);
nor U8387 (N_8387,N_1960,N_4464);
xor U8388 (N_8388,N_1997,N_3743);
or U8389 (N_8389,N_4208,N_2212);
or U8390 (N_8390,N_2380,N_792);
nor U8391 (N_8391,N_3229,N_3040);
nand U8392 (N_8392,N_41,N_2966);
nand U8393 (N_8393,N_2427,N_669);
nor U8394 (N_8394,N_409,N_1389);
nor U8395 (N_8395,N_1648,N_3924);
or U8396 (N_8396,N_2609,N_1677);
nor U8397 (N_8397,N_442,N_386);
and U8398 (N_8398,N_4123,N_2516);
xor U8399 (N_8399,N_160,N_4162);
and U8400 (N_8400,N_207,N_1923);
nand U8401 (N_8401,N_1966,N_2854);
nor U8402 (N_8402,N_128,N_2080);
and U8403 (N_8403,N_4412,N_2373);
and U8404 (N_8404,N_3120,N_3687);
and U8405 (N_8405,N_3552,N_4033);
nand U8406 (N_8406,N_117,N_3725);
and U8407 (N_8407,N_1470,N_4011);
nand U8408 (N_8408,N_3983,N_2810);
or U8409 (N_8409,N_1311,N_1363);
xnor U8410 (N_8410,N_2876,N_4966);
or U8411 (N_8411,N_3077,N_766);
and U8412 (N_8412,N_2569,N_3202);
or U8413 (N_8413,N_3511,N_731);
or U8414 (N_8414,N_4323,N_4397);
xnor U8415 (N_8415,N_4083,N_4259);
or U8416 (N_8416,N_1917,N_4342);
or U8417 (N_8417,N_977,N_3817);
nor U8418 (N_8418,N_3541,N_1949);
nand U8419 (N_8419,N_2284,N_4675);
or U8420 (N_8420,N_867,N_1587);
or U8421 (N_8421,N_2437,N_3518);
or U8422 (N_8422,N_4333,N_2912);
nor U8423 (N_8423,N_2151,N_3590);
nor U8424 (N_8424,N_2841,N_2265);
nand U8425 (N_8425,N_4146,N_2746);
or U8426 (N_8426,N_3825,N_3017);
and U8427 (N_8427,N_3152,N_591);
xnor U8428 (N_8428,N_942,N_3461);
nand U8429 (N_8429,N_1291,N_115);
and U8430 (N_8430,N_1669,N_762);
nand U8431 (N_8431,N_2541,N_4954);
nor U8432 (N_8432,N_1125,N_1878);
nand U8433 (N_8433,N_4155,N_2815);
nor U8434 (N_8434,N_1806,N_4208);
or U8435 (N_8435,N_3824,N_107);
or U8436 (N_8436,N_2848,N_2999);
nand U8437 (N_8437,N_3197,N_516);
nand U8438 (N_8438,N_1066,N_3685);
nor U8439 (N_8439,N_3528,N_3764);
nor U8440 (N_8440,N_1186,N_3362);
or U8441 (N_8441,N_3968,N_828);
nor U8442 (N_8442,N_615,N_4752);
nor U8443 (N_8443,N_4680,N_1254);
and U8444 (N_8444,N_616,N_1161);
and U8445 (N_8445,N_2234,N_3641);
or U8446 (N_8446,N_1205,N_540);
and U8447 (N_8447,N_2189,N_4856);
nor U8448 (N_8448,N_401,N_3277);
nor U8449 (N_8449,N_1671,N_556);
or U8450 (N_8450,N_1871,N_236);
or U8451 (N_8451,N_1631,N_4483);
or U8452 (N_8452,N_4557,N_1704);
nand U8453 (N_8453,N_4532,N_645);
and U8454 (N_8454,N_2747,N_818);
or U8455 (N_8455,N_2745,N_3452);
and U8456 (N_8456,N_1050,N_2366);
xnor U8457 (N_8457,N_4292,N_201);
and U8458 (N_8458,N_603,N_1696);
xor U8459 (N_8459,N_4033,N_321);
xor U8460 (N_8460,N_980,N_1901);
nand U8461 (N_8461,N_2009,N_3682);
and U8462 (N_8462,N_3024,N_992);
or U8463 (N_8463,N_3692,N_4467);
nor U8464 (N_8464,N_3661,N_3962);
nand U8465 (N_8465,N_2135,N_4021);
nor U8466 (N_8466,N_870,N_4422);
and U8467 (N_8467,N_2252,N_2836);
nor U8468 (N_8468,N_3142,N_1738);
and U8469 (N_8469,N_1023,N_4221);
nand U8470 (N_8470,N_3833,N_673);
or U8471 (N_8471,N_3135,N_2544);
nand U8472 (N_8472,N_1993,N_528);
and U8473 (N_8473,N_3588,N_3939);
xor U8474 (N_8474,N_4237,N_2377);
xor U8475 (N_8475,N_4758,N_2310);
nor U8476 (N_8476,N_1050,N_4483);
or U8477 (N_8477,N_408,N_3566);
and U8478 (N_8478,N_812,N_3749);
and U8479 (N_8479,N_3327,N_310);
xor U8480 (N_8480,N_2639,N_2419);
and U8481 (N_8481,N_4475,N_17);
nor U8482 (N_8482,N_2062,N_2035);
and U8483 (N_8483,N_2220,N_4878);
or U8484 (N_8484,N_2859,N_2710);
xor U8485 (N_8485,N_3129,N_1552);
and U8486 (N_8486,N_1088,N_1712);
or U8487 (N_8487,N_2477,N_4604);
xor U8488 (N_8488,N_1891,N_476);
nor U8489 (N_8489,N_113,N_443);
nand U8490 (N_8490,N_3129,N_4248);
and U8491 (N_8491,N_761,N_2389);
nor U8492 (N_8492,N_3112,N_3883);
xnor U8493 (N_8493,N_401,N_2699);
or U8494 (N_8494,N_1873,N_2238);
nand U8495 (N_8495,N_4554,N_1332);
or U8496 (N_8496,N_2334,N_3495);
or U8497 (N_8497,N_4493,N_1387);
and U8498 (N_8498,N_2398,N_2171);
or U8499 (N_8499,N_4968,N_2520);
or U8500 (N_8500,N_3544,N_2759);
nor U8501 (N_8501,N_1335,N_1648);
nand U8502 (N_8502,N_439,N_4529);
and U8503 (N_8503,N_2451,N_426);
and U8504 (N_8504,N_1959,N_3876);
nor U8505 (N_8505,N_2358,N_1876);
nand U8506 (N_8506,N_4320,N_3093);
and U8507 (N_8507,N_1924,N_3744);
nor U8508 (N_8508,N_4880,N_4736);
and U8509 (N_8509,N_2927,N_686);
nand U8510 (N_8510,N_3753,N_3247);
nor U8511 (N_8511,N_2088,N_3313);
nor U8512 (N_8512,N_3796,N_714);
nand U8513 (N_8513,N_1174,N_4491);
or U8514 (N_8514,N_950,N_1319);
and U8515 (N_8515,N_2663,N_1061);
nand U8516 (N_8516,N_1550,N_442);
or U8517 (N_8517,N_3643,N_2185);
nand U8518 (N_8518,N_4667,N_1221);
and U8519 (N_8519,N_4602,N_346);
xor U8520 (N_8520,N_4089,N_406);
nor U8521 (N_8521,N_2635,N_1652);
and U8522 (N_8522,N_3925,N_1167);
xnor U8523 (N_8523,N_2771,N_339);
nand U8524 (N_8524,N_3865,N_883);
nor U8525 (N_8525,N_1832,N_2784);
nor U8526 (N_8526,N_3790,N_4596);
and U8527 (N_8527,N_194,N_2000);
xor U8528 (N_8528,N_4809,N_3825);
or U8529 (N_8529,N_4277,N_2138);
or U8530 (N_8530,N_1433,N_2292);
nand U8531 (N_8531,N_4682,N_4057);
and U8532 (N_8532,N_3746,N_1250);
nand U8533 (N_8533,N_3602,N_595);
nand U8534 (N_8534,N_3959,N_394);
and U8535 (N_8535,N_1921,N_2752);
or U8536 (N_8536,N_2996,N_4819);
nand U8537 (N_8537,N_4025,N_2624);
nor U8538 (N_8538,N_204,N_2278);
and U8539 (N_8539,N_3988,N_2469);
or U8540 (N_8540,N_850,N_2354);
nor U8541 (N_8541,N_758,N_1409);
nor U8542 (N_8542,N_2638,N_999);
or U8543 (N_8543,N_315,N_1544);
and U8544 (N_8544,N_2484,N_3278);
and U8545 (N_8545,N_4853,N_289);
xnor U8546 (N_8546,N_4879,N_4249);
nor U8547 (N_8547,N_1974,N_2810);
nor U8548 (N_8548,N_2916,N_3647);
or U8549 (N_8549,N_4143,N_2899);
or U8550 (N_8550,N_1951,N_3974);
or U8551 (N_8551,N_3978,N_2733);
or U8552 (N_8552,N_313,N_1984);
nand U8553 (N_8553,N_1419,N_3311);
xnor U8554 (N_8554,N_3159,N_3177);
xnor U8555 (N_8555,N_2759,N_4680);
or U8556 (N_8556,N_501,N_1658);
nand U8557 (N_8557,N_3057,N_3961);
nand U8558 (N_8558,N_1952,N_2525);
xnor U8559 (N_8559,N_484,N_2841);
or U8560 (N_8560,N_4447,N_2321);
or U8561 (N_8561,N_1221,N_2584);
and U8562 (N_8562,N_4840,N_557);
or U8563 (N_8563,N_3425,N_1068);
nand U8564 (N_8564,N_2239,N_2267);
nor U8565 (N_8565,N_3122,N_1531);
nor U8566 (N_8566,N_4669,N_160);
and U8567 (N_8567,N_642,N_3088);
xor U8568 (N_8568,N_4234,N_1875);
or U8569 (N_8569,N_4887,N_3268);
nor U8570 (N_8570,N_681,N_261);
and U8571 (N_8571,N_3528,N_4235);
nand U8572 (N_8572,N_3075,N_4624);
or U8573 (N_8573,N_3151,N_1919);
nor U8574 (N_8574,N_1862,N_4645);
or U8575 (N_8575,N_411,N_2164);
nand U8576 (N_8576,N_1977,N_2902);
nor U8577 (N_8577,N_4387,N_1807);
xor U8578 (N_8578,N_1458,N_621);
nor U8579 (N_8579,N_4107,N_3586);
xnor U8580 (N_8580,N_2412,N_3716);
or U8581 (N_8581,N_3642,N_4979);
nand U8582 (N_8582,N_1751,N_1547);
nor U8583 (N_8583,N_3650,N_3038);
or U8584 (N_8584,N_135,N_1620);
and U8585 (N_8585,N_2184,N_1228);
nand U8586 (N_8586,N_3605,N_1431);
and U8587 (N_8587,N_3294,N_3558);
or U8588 (N_8588,N_940,N_4424);
and U8589 (N_8589,N_357,N_4875);
nand U8590 (N_8590,N_4276,N_2127);
and U8591 (N_8591,N_848,N_1905);
nand U8592 (N_8592,N_1973,N_1533);
nor U8593 (N_8593,N_3439,N_4688);
nor U8594 (N_8594,N_3647,N_3522);
nand U8595 (N_8595,N_2190,N_682);
nand U8596 (N_8596,N_4822,N_1166);
nand U8597 (N_8597,N_3915,N_997);
or U8598 (N_8598,N_989,N_2454);
and U8599 (N_8599,N_3592,N_1127);
xnor U8600 (N_8600,N_3800,N_1911);
nand U8601 (N_8601,N_275,N_356);
nor U8602 (N_8602,N_4477,N_3443);
nand U8603 (N_8603,N_2386,N_3578);
nand U8604 (N_8604,N_2704,N_3604);
and U8605 (N_8605,N_4694,N_4092);
nand U8606 (N_8606,N_2756,N_4181);
nor U8607 (N_8607,N_553,N_3241);
nor U8608 (N_8608,N_1735,N_2306);
and U8609 (N_8609,N_1323,N_783);
or U8610 (N_8610,N_355,N_1133);
xnor U8611 (N_8611,N_4571,N_2622);
nor U8612 (N_8612,N_2722,N_54);
nand U8613 (N_8613,N_1314,N_1005);
and U8614 (N_8614,N_2798,N_1615);
and U8615 (N_8615,N_4977,N_3274);
nand U8616 (N_8616,N_1659,N_1027);
or U8617 (N_8617,N_4000,N_4361);
and U8618 (N_8618,N_2315,N_989);
xnor U8619 (N_8619,N_655,N_4586);
or U8620 (N_8620,N_4389,N_3886);
and U8621 (N_8621,N_4285,N_1446);
nand U8622 (N_8622,N_3072,N_3109);
and U8623 (N_8623,N_595,N_615);
or U8624 (N_8624,N_4541,N_1449);
nor U8625 (N_8625,N_3676,N_2994);
and U8626 (N_8626,N_1352,N_1514);
nor U8627 (N_8627,N_2965,N_4279);
nand U8628 (N_8628,N_3377,N_2266);
xnor U8629 (N_8629,N_4879,N_3185);
and U8630 (N_8630,N_1697,N_3071);
or U8631 (N_8631,N_3221,N_2992);
nor U8632 (N_8632,N_2950,N_836);
and U8633 (N_8633,N_4042,N_1051);
xor U8634 (N_8634,N_107,N_63);
or U8635 (N_8635,N_3757,N_2168);
and U8636 (N_8636,N_4451,N_729);
and U8637 (N_8637,N_720,N_2002);
nor U8638 (N_8638,N_1,N_529);
and U8639 (N_8639,N_1755,N_730);
nand U8640 (N_8640,N_1167,N_4738);
or U8641 (N_8641,N_3123,N_770);
and U8642 (N_8642,N_4297,N_4784);
nor U8643 (N_8643,N_349,N_4868);
nor U8644 (N_8644,N_2618,N_3824);
and U8645 (N_8645,N_1502,N_4815);
and U8646 (N_8646,N_4510,N_384);
and U8647 (N_8647,N_3642,N_1014);
or U8648 (N_8648,N_4007,N_3118);
or U8649 (N_8649,N_4787,N_2983);
xor U8650 (N_8650,N_833,N_3123);
and U8651 (N_8651,N_1007,N_1318);
and U8652 (N_8652,N_4018,N_3070);
and U8653 (N_8653,N_851,N_6);
or U8654 (N_8654,N_4522,N_2691);
and U8655 (N_8655,N_560,N_2093);
nand U8656 (N_8656,N_3732,N_2274);
nand U8657 (N_8657,N_987,N_4705);
and U8658 (N_8658,N_2842,N_941);
nor U8659 (N_8659,N_1964,N_3711);
nand U8660 (N_8660,N_1238,N_3128);
nor U8661 (N_8661,N_1428,N_190);
or U8662 (N_8662,N_1816,N_3014);
or U8663 (N_8663,N_3525,N_4677);
and U8664 (N_8664,N_2948,N_3103);
nand U8665 (N_8665,N_2450,N_2119);
and U8666 (N_8666,N_2081,N_1768);
nor U8667 (N_8667,N_1693,N_1472);
and U8668 (N_8668,N_958,N_1514);
nand U8669 (N_8669,N_1000,N_4296);
nand U8670 (N_8670,N_4758,N_3267);
or U8671 (N_8671,N_2945,N_1071);
nor U8672 (N_8672,N_3879,N_2750);
and U8673 (N_8673,N_1767,N_3107);
nor U8674 (N_8674,N_2911,N_1208);
xor U8675 (N_8675,N_380,N_4883);
and U8676 (N_8676,N_4313,N_2016);
or U8677 (N_8677,N_3149,N_4873);
and U8678 (N_8678,N_3046,N_2766);
nand U8679 (N_8679,N_884,N_3512);
nor U8680 (N_8680,N_1649,N_2039);
nor U8681 (N_8681,N_980,N_4960);
and U8682 (N_8682,N_557,N_1014);
and U8683 (N_8683,N_860,N_4336);
or U8684 (N_8684,N_291,N_87);
or U8685 (N_8685,N_1059,N_1920);
xor U8686 (N_8686,N_3908,N_59);
or U8687 (N_8687,N_121,N_2175);
nand U8688 (N_8688,N_1565,N_4895);
or U8689 (N_8689,N_3927,N_1023);
nand U8690 (N_8690,N_922,N_2855);
nand U8691 (N_8691,N_4179,N_3713);
nor U8692 (N_8692,N_3739,N_4315);
nor U8693 (N_8693,N_1788,N_2149);
or U8694 (N_8694,N_3946,N_2742);
nand U8695 (N_8695,N_4614,N_2099);
and U8696 (N_8696,N_4494,N_4304);
nand U8697 (N_8697,N_2186,N_4677);
nor U8698 (N_8698,N_430,N_82);
nor U8699 (N_8699,N_1784,N_3598);
nor U8700 (N_8700,N_3622,N_1722);
and U8701 (N_8701,N_4639,N_4004);
or U8702 (N_8702,N_4394,N_842);
nand U8703 (N_8703,N_3076,N_675);
and U8704 (N_8704,N_4015,N_3325);
xor U8705 (N_8705,N_1092,N_4368);
nand U8706 (N_8706,N_4702,N_4995);
nand U8707 (N_8707,N_1657,N_2478);
nor U8708 (N_8708,N_4241,N_3803);
nand U8709 (N_8709,N_2791,N_325);
or U8710 (N_8710,N_1326,N_4712);
nand U8711 (N_8711,N_1667,N_1385);
nor U8712 (N_8712,N_1305,N_626);
and U8713 (N_8713,N_2811,N_2948);
and U8714 (N_8714,N_2989,N_3648);
nor U8715 (N_8715,N_131,N_4118);
and U8716 (N_8716,N_3869,N_3856);
nand U8717 (N_8717,N_1513,N_2477);
and U8718 (N_8718,N_289,N_474);
nor U8719 (N_8719,N_4308,N_3322);
or U8720 (N_8720,N_2814,N_4247);
nand U8721 (N_8721,N_4670,N_70);
and U8722 (N_8722,N_4444,N_2318);
nor U8723 (N_8723,N_4734,N_4394);
nor U8724 (N_8724,N_3036,N_600);
and U8725 (N_8725,N_4804,N_485);
nand U8726 (N_8726,N_4571,N_1498);
and U8727 (N_8727,N_1480,N_275);
or U8728 (N_8728,N_2299,N_615);
xnor U8729 (N_8729,N_3255,N_4778);
nand U8730 (N_8730,N_3861,N_2485);
and U8731 (N_8731,N_4660,N_3624);
or U8732 (N_8732,N_2859,N_385);
or U8733 (N_8733,N_2015,N_3079);
nand U8734 (N_8734,N_3507,N_1488);
nor U8735 (N_8735,N_3060,N_435);
nand U8736 (N_8736,N_3871,N_1312);
nand U8737 (N_8737,N_601,N_664);
and U8738 (N_8738,N_600,N_1443);
and U8739 (N_8739,N_3416,N_2018);
and U8740 (N_8740,N_3918,N_1238);
xor U8741 (N_8741,N_2275,N_3589);
nor U8742 (N_8742,N_2858,N_4929);
or U8743 (N_8743,N_4992,N_1502);
and U8744 (N_8744,N_328,N_1589);
nand U8745 (N_8745,N_3067,N_1184);
nor U8746 (N_8746,N_2353,N_3591);
nand U8747 (N_8747,N_249,N_2344);
and U8748 (N_8748,N_4628,N_116);
xor U8749 (N_8749,N_1279,N_2939);
nor U8750 (N_8750,N_1921,N_1300);
or U8751 (N_8751,N_950,N_4323);
nor U8752 (N_8752,N_3542,N_2250);
or U8753 (N_8753,N_1593,N_2781);
and U8754 (N_8754,N_2644,N_3004);
or U8755 (N_8755,N_1760,N_3030);
xor U8756 (N_8756,N_3298,N_4952);
nor U8757 (N_8757,N_3654,N_2505);
nor U8758 (N_8758,N_4332,N_4086);
nand U8759 (N_8759,N_363,N_2282);
and U8760 (N_8760,N_3893,N_3105);
or U8761 (N_8761,N_210,N_3282);
nor U8762 (N_8762,N_2265,N_3228);
and U8763 (N_8763,N_1415,N_2529);
nor U8764 (N_8764,N_4408,N_1484);
nor U8765 (N_8765,N_1155,N_1043);
and U8766 (N_8766,N_2475,N_3836);
or U8767 (N_8767,N_3041,N_1137);
nand U8768 (N_8768,N_24,N_1138);
and U8769 (N_8769,N_4090,N_1883);
and U8770 (N_8770,N_4671,N_2391);
or U8771 (N_8771,N_805,N_2427);
nor U8772 (N_8772,N_3041,N_4141);
and U8773 (N_8773,N_3327,N_3990);
and U8774 (N_8774,N_4827,N_2438);
nor U8775 (N_8775,N_2503,N_1697);
nand U8776 (N_8776,N_2224,N_7);
xor U8777 (N_8777,N_4935,N_406);
nor U8778 (N_8778,N_4177,N_4389);
and U8779 (N_8779,N_2572,N_2117);
nand U8780 (N_8780,N_1501,N_4943);
or U8781 (N_8781,N_4724,N_3438);
nand U8782 (N_8782,N_384,N_137);
nor U8783 (N_8783,N_711,N_4782);
and U8784 (N_8784,N_423,N_435);
and U8785 (N_8785,N_402,N_2897);
or U8786 (N_8786,N_4137,N_4517);
xnor U8787 (N_8787,N_1412,N_4725);
and U8788 (N_8788,N_83,N_4835);
and U8789 (N_8789,N_234,N_2638);
nor U8790 (N_8790,N_4949,N_3776);
nand U8791 (N_8791,N_3076,N_4766);
nor U8792 (N_8792,N_1299,N_2275);
nor U8793 (N_8793,N_3967,N_2888);
or U8794 (N_8794,N_332,N_3124);
and U8795 (N_8795,N_1724,N_3830);
and U8796 (N_8796,N_4888,N_3980);
nor U8797 (N_8797,N_4648,N_1932);
nand U8798 (N_8798,N_1373,N_2787);
nand U8799 (N_8799,N_3957,N_1492);
xor U8800 (N_8800,N_860,N_3200);
xnor U8801 (N_8801,N_889,N_1051);
nor U8802 (N_8802,N_455,N_3163);
and U8803 (N_8803,N_1240,N_4881);
nand U8804 (N_8804,N_2700,N_1747);
xnor U8805 (N_8805,N_4308,N_4657);
xor U8806 (N_8806,N_2340,N_1279);
xor U8807 (N_8807,N_3249,N_2916);
nand U8808 (N_8808,N_3758,N_3968);
nand U8809 (N_8809,N_1822,N_797);
or U8810 (N_8810,N_4886,N_2515);
and U8811 (N_8811,N_2512,N_4585);
and U8812 (N_8812,N_4457,N_777);
nand U8813 (N_8813,N_3492,N_1690);
and U8814 (N_8814,N_1110,N_4344);
nand U8815 (N_8815,N_4381,N_5);
nor U8816 (N_8816,N_3928,N_2484);
nand U8817 (N_8817,N_794,N_4618);
xnor U8818 (N_8818,N_4814,N_4063);
nor U8819 (N_8819,N_1539,N_2359);
or U8820 (N_8820,N_3366,N_3520);
nor U8821 (N_8821,N_4687,N_474);
nor U8822 (N_8822,N_473,N_680);
nor U8823 (N_8823,N_4819,N_1563);
nor U8824 (N_8824,N_3575,N_4187);
or U8825 (N_8825,N_4469,N_3205);
nand U8826 (N_8826,N_4903,N_1304);
and U8827 (N_8827,N_2372,N_2431);
nor U8828 (N_8828,N_4847,N_1084);
and U8829 (N_8829,N_1917,N_3654);
nor U8830 (N_8830,N_4688,N_4521);
or U8831 (N_8831,N_1544,N_1849);
nor U8832 (N_8832,N_976,N_1255);
xor U8833 (N_8833,N_2311,N_1683);
nor U8834 (N_8834,N_3134,N_2669);
nor U8835 (N_8835,N_650,N_2108);
or U8836 (N_8836,N_4770,N_29);
nor U8837 (N_8837,N_3103,N_3988);
and U8838 (N_8838,N_3224,N_2429);
nand U8839 (N_8839,N_4151,N_1820);
and U8840 (N_8840,N_1825,N_4256);
or U8841 (N_8841,N_936,N_348);
xnor U8842 (N_8842,N_400,N_2434);
nor U8843 (N_8843,N_4216,N_25);
and U8844 (N_8844,N_1109,N_704);
and U8845 (N_8845,N_3566,N_1027);
or U8846 (N_8846,N_4614,N_1906);
nor U8847 (N_8847,N_28,N_4217);
or U8848 (N_8848,N_4772,N_439);
and U8849 (N_8849,N_1959,N_3442);
and U8850 (N_8850,N_377,N_1848);
and U8851 (N_8851,N_608,N_2065);
and U8852 (N_8852,N_1948,N_1631);
or U8853 (N_8853,N_4406,N_3786);
or U8854 (N_8854,N_4471,N_4994);
nor U8855 (N_8855,N_1464,N_1124);
xor U8856 (N_8856,N_886,N_687);
and U8857 (N_8857,N_3968,N_916);
nand U8858 (N_8858,N_3742,N_1961);
nor U8859 (N_8859,N_2730,N_698);
and U8860 (N_8860,N_3030,N_4457);
nand U8861 (N_8861,N_4844,N_825);
and U8862 (N_8862,N_3630,N_4898);
or U8863 (N_8863,N_3788,N_3848);
nor U8864 (N_8864,N_3455,N_3016);
nand U8865 (N_8865,N_4835,N_1712);
nor U8866 (N_8866,N_1973,N_2884);
and U8867 (N_8867,N_4705,N_887);
nand U8868 (N_8868,N_909,N_748);
nor U8869 (N_8869,N_748,N_2028);
nand U8870 (N_8870,N_1849,N_2649);
nor U8871 (N_8871,N_4940,N_2890);
nor U8872 (N_8872,N_4054,N_3889);
nand U8873 (N_8873,N_1309,N_3334);
and U8874 (N_8874,N_3535,N_3500);
nand U8875 (N_8875,N_5,N_3644);
and U8876 (N_8876,N_559,N_2154);
nand U8877 (N_8877,N_4425,N_4000);
nor U8878 (N_8878,N_716,N_2957);
nor U8879 (N_8879,N_2768,N_4779);
and U8880 (N_8880,N_4750,N_3276);
and U8881 (N_8881,N_1735,N_3009);
or U8882 (N_8882,N_463,N_2088);
xor U8883 (N_8883,N_3302,N_1557);
xnor U8884 (N_8884,N_3728,N_1273);
xnor U8885 (N_8885,N_4272,N_4993);
xnor U8886 (N_8886,N_2798,N_4073);
and U8887 (N_8887,N_2482,N_2185);
nor U8888 (N_8888,N_514,N_2936);
nand U8889 (N_8889,N_2832,N_206);
xnor U8890 (N_8890,N_3016,N_3491);
or U8891 (N_8891,N_4876,N_496);
nor U8892 (N_8892,N_1842,N_3072);
xnor U8893 (N_8893,N_335,N_1705);
or U8894 (N_8894,N_1956,N_1686);
xor U8895 (N_8895,N_4277,N_4545);
or U8896 (N_8896,N_4603,N_2814);
nor U8897 (N_8897,N_1152,N_2594);
and U8898 (N_8898,N_417,N_1900);
nand U8899 (N_8899,N_2654,N_3679);
nor U8900 (N_8900,N_155,N_1361);
nor U8901 (N_8901,N_3862,N_3527);
nand U8902 (N_8902,N_3759,N_3158);
nor U8903 (N_8903,N_4560,N_666);
and U8904 (N_8904,N_2341,N_3409);
nand U8905 (N_8905,N_993,N_1329);
nand U8906 (N_8906,N_2557,N_1539);
nor U8907 (N_8907,N_210,N_4294);
or U8908 (N_8908,N_3178,N_2405);
and U8909 (N_8909,N_3274,N_2465);
nand U8910 (N_8910,N_425,N_3230);
xnor U8911 (N_8911,N_3697,N_3846);
nor U8912 (N_8912,N_4799,N_703);
or U8913 (N_8913,N_3729,N_2338);
nor U8914 (N_8914,N_4874,N_1767);
nor U8915 (N_8915,N_1515,N_2468);
nor U8916 (N_8916,N_1732,N_4059);
nor U8917 (N_8917,N_3092,N_4426);
and U8918 (N_8918,N_4796,N_2929);
nor U8919 (N_8919,N_3017,N_3773);
xor U8920 (N_8920,N_978,N_733);
nand U8921 (N_8921,N_4872,N_744);
nor U8922 (N_8922,N_1326,N_2089);
nor U8923 (N_8923,N_2718,N_4963);
nor U8924 (N_8924,N_4483,N_941);
and U8925 (N_8925,N_1186,N_2984);
nand U8926 (N_8926,N_3138,N_88);
xnor U8927 (N_8927,N_665,N_3850);
or U8928 (N_8928,N_3158,N_4224);
nor U8929 (N_8929,N_3750,N_1982);
or U8930 (N_8930,N_2899,N_2179);
nand U8931 (N_8931,N_135,N_3497);
nor U8932 (N_8932,N_4778,N_35);
and U8933 (N_8933,N_612,N_196);
xor U8934 (N_8934,N_4742,N_558);
nand U8935 (N_8935,N_939,N_1149);
nand U8936 (N_8936,N_4404,N_2307);
nor U8937 (N_8937,N_4933,N_397);
xnor U8938 (N_8938,N_856,N_3730);
nand U8939 (N_8939,N_4364,N_1035);
xnor U8940 (N_8940,N_246,N_3471);
nor U8941 (N_8941,N_2342,N_4651);
nand U8942 (N_8942,N_3102,N_1083);
and U8943 (N_8943,N_3363,N_2519);
xnor U8944 (N_8944,N_4142,N_1953);
nand U8945 (N_8945,N_3809,N_4135);
and U8946 (N_8946,N_606,N_3905);
xor U8947 (N_8947,N_882,N_2440);
nor U8948 (N_8948,N_2539,N_3130);
and U8949 (N_8949,N_3751,N_2970);
nand U8950 (N_8950,N_4712,N_1223);
or U8951 (N_8951,N_690,N_4468);
and U8952 (N_8952,N_4505,N_4775);
or U8953 (N_8953,N_306,N_3189);
nor U8954 (N_8954,N_3830,N_28);
or U8955 (N_8955,N_3331,N_2098);
nor U8956 (N_8956,N_1358,N_4040);
or U8957 (N_8957,N_2364,N_2983);
xnor U8958 (N_8958,N_4404,N_4719);
xor U8959 (N_8959,N_768,N_2579);
nor U8960 (N_8960,N_3355,N_2642);
nand U8961 (N_8961,N_1858,N_3770);
or U8962 (N_8962,N_1926,N_2504);
nor U8963 (N_8963,N_2360,N_859);
nor U8964 (N_8964,N_2599,N_2864);
xnor U8965 (N_8965,N_1758,N_4747);
or U8966 (N_8966,N_3732,N_99);
or U8967 (N_8967,N_458,N_1209);
xnor U8968 (N_8968,N_3928,N_775);
nand U8969 (N_8969,N_815,N_4081);
or U8970 (N_8970,N_3422,N_1740);
or U8971 (N_8971,N_4145,N_4556);
and U8972 (N_8972,N_2935,N_709);
nand U8973 (N_8973,N_3912,N_213);
or U8974 (N_8974,N_923,N_3927);
nand U8975 (N_8975,N_4000,N_4098);
nand U8976 (N_8976,N_1760,N_1649);
nor U8977 (N_8977,N_1857,N_2734);
nand U8978 (N_8978,N_4383,N_3241);
nand U8979 (N_8979,N_810,N_583);
nor U8980 (N_8980,N_2329,N_2641);
nor U8981 (N_8981,N_4392,N_1572);
nand U8982 (N_8982,N_2037,N_1685);
or U8983 (N_8983,N_1832,N_893);
or U8984 (N_8984,N_3216,N_3690);
nor U8985 (N_8985,N_4437,N_3279);
nor U8986 (N_8986,N_4971,N_577);
nor U8987 (N_8987,N_1329,N_3772);
nor U8988 (N_8988,N_2497,N_4166);
nor U8989 (N_8989,N_1130,N_2764);
nor U8990 (N_8990,N_600,N_422);
and U8991 (N_8991,N_3721,N_1392);
or U8992 (N_8992,N_2033,N_2032);
nand U8993 (N_8993,N_3488,N_2297);
xnor U8994 (N_8994,N_897,N_2976);
and U8995 (N_8995,N_2264,N_4561);
and U8996 (N_8996,N_4508,N_975);
xor U8997 (N_8997,N_1001,N_7);
nor U8998 (N_8998,N_4021,N_1038);
or U8999 (N_8999,N_4600,N_2774);
or U9000 (N_9000,N_791,N_3322);
xnor U9001 (N_9001,N_3799,N_82);
nor U9002 (N_9002,N_3650,N_399);
nor U9003 (N_9003,N_2321,N_117);
nand U9004 (N_9004,N_3397,N_3120);
and U9005 (N_9005,N_1639,N_4650);
nand U9006 (N_9006,N_639,N_2260);
or U9007 (N_9007,N_1800,N_705);
nor U9008 (N_9008,N_1440,N_45);
nor U9009 (N_9009,N_3232,N_2778);
and U9010 (N_9010,N_3238,N_563);
and U9011 (N_9011,N_2490,N_3256);
nor U9012 (N_9012,N_2615,N_4846);
nor U9013 (N_9013,N_4111,N_4362);
or U9014 (N_9014,N_4553,N_1588);
xnor U9015 (N_9015,N_4358,N_657);
and U9016 (N_9016,N_2654,N_40);
nand U9017 (N_9017,N_1385,N_4332);
and U9018 (N_9018,N_90,N_544);
or U9019 (N_9019,N_1328,N_1920);
nor U9020 (N_9020,N_3838,N_264);
nor U9021 (N_9021,N_909,N_861);
nand U9022 (N_9022,N_2842,N_1917);
and U9023 (N_9023,N_4831,N_599);
nor U9024 (N_9024,N_623,N_383);
and U9025 (N_9025,N_1511,N_4762);
nor U9026 (N_9026,N_4969,N_567);
or U9027 (N_9027,N_2328,N_1420);
and U9028 (N_9028,N_597,N_1249);
nand U9029 (N_9029,N_3516,N_868);
nand U9030 (N_9030,N_1247,N_4104);
and U9031 (N_9031,N_2614,N_3059);
or U9032 (N_9032,N_1476,N_3475);
and U9033 (N_9033,N_3858,N_1098);
and U9034 (N_9034,N_4231,N_2490);
and U9035 (N_9035,N_728,N_749);
and U9036 (N_9036,N_2861,N_3653);
or U9037 (N_9037,N_1923,N_3426);
xor U9038 (N_9038,N_1376,N_2629);
and U9039 (N_9039,N_288,N_3209);
nand U9040 (N_9040,N_2000,N_720);
or U9041 (N_9041,N_1661,N_4144);
nor U9042 (N_9042,N_4759,N_896);
nor U9043 (N_9043,N_4260,N_4379);
xnor U9044 (N_9044,N_3705,N_587);
or U9045 (N_9045,N_57,N_2988);
nand U9046 (N_9046,N_1893,N_2836);
and U9047 (N_9047,N_777,N_1487);
nand U9048 (N_9048,N_3600,N_2848);
nand U9049 (N_9049,N_4142,N_2056);
nand U9050 (N_9050,N_4241,N_2107);
and U9051 (N_9051,N_2302,N_4380);
nor U9052 (N_9052,N_4697,N_4346);
nand U9053 (N_9053,N_3001,N_2680);
or U9054 (N_9054,N_3877,N_1714);
nor U9055 (N_9055,N_3273,N_3440);
or U9056 (N_9056,N_1034,N_2678);
and U9057 (N_9057,N_2931,N_3486);
and U9058 (N_9058,N_2656,N_4875);
nor U9059 (N_9059,N_3348,N_2673);
and U9060 (N_9060,N_3470,N_3252);
and U9061 (N_9061,N_1673,N_1526);
nand U9062 (N_9062,N_1250,N_1619);
nand U9063 (N_9063,N_3533,N_2218);
and U9064 (N_9064,N_123,N_2267);
xor U9065 (N_9065,N_420,N_856);
nand U9066 (N_9066,N_4419,N_3109);
nor U9067 (N_9067,N_2896,N_518);
nand U9068 (N_9068,N_3295,N_3527);
nor U9069 (N_9069,N_3765,N_16);
nand U9070 (N_9070,N_2022,N_1603);
nor U9071 (N_9071,N_3455,N_1313);
nor U9072 (N_9072,N_817,N_3677);
and U9073 (N_9073,N_4347,N_729);
or U9074 (N_9074,N_3131,N_28);
or U9075 (N_9075,N_2337,N_2013);
and U9076 (N_9076,N_4826,N_4989);
or U9077 (N_9077,N_1950,N_3935);
and U9078 (N_9078,N_3528,N_2053);
or U9079 (N_9079,N_59,N_3552);
or U9080 (N_9080,N_473,N_444);
nor U9081 (N_9081,N_3080,N_2687);
and U9082 (N_9082,N_1459,N_1513);
or U9083 (N_9083,N_4429,N_3373);
or U9084 (N_9084,N_2704,N_4588);
nand U9085 (N_9085,N_1383,N_1833);
nand U9086 (N_9086,N_1636,N_4957);
and U9087 (N_9087,N_2225,N_3627);
nand U9088 (N_9088,N_4640,N_2419);
or U9089 (N_9089,N_1251,N_263);
and U9090 (N_9090,N_3608,N_700);
and U9091 (N_9091,N_2329,N_4049);
or U9092 (N_9092,N_1329,N_3275);
and U9093 (N_9093,N_2955,N_2767);
or U9094 (N_9094,N_1772,N_1499);
xor U9095 (N_9095,N_3249,N_4109);
nor U9096 (N_9096,N_4101,N_2370);
nand U9097 (N_9097,N_3338,N_1483);
or U9098 (N_9098,N_2404,N_2461);
nor U9099 (N_9099,N_188,N_3280);
or U9100 (N_9100,N_4220,N_4776);
or U9101 (N_9101,N_4042,N_257);
and U9102 (N_9102,N_1181,N_3537);
or U9103 (N_9103,N_3712,N_1304);
or U9104 (N_9104,N_3250,N_3400);
nor U9105 (N_9105,N_2536,N_2250);
and U9106 (N_9106,N_4914,N_2765);
xor U9107 (N_9107,N_2940,N_1085);
nand U9108 (N_9108,N_603,N_4397);
nand U9109 (N_9109,N_4248,N_3322);
nor U9110 (N_9110,N_1325,N_1648);
nand U9111 (N_9111,N_4616,N_3617);
and U9112 (N_9112,N_3259,N_2923);
or U9113 (N_9113,N_3944,N_899);
nor U9114 (N_9114,N_3641,N_721);
and U9115 (N_9115,N_3708,N_3139);
and U9116 (N_9116,N_325,N_4988);
xnor U9117 (N_9117,N_1186,N_2247);
nor U9118 (N_9118,N_3015,N_1841);
and U9119 (N_9119,N_2064,N_1636);
or U9120 (N_9120,N_2655,N_1924);
nand U9121 (N_9121,N_3460,N_759);
or U9122 (N_9122,N_25,N_1778);
or U9123 (N_9123,N_1434,N_3595);
nor U9124 (N_9124,N_4013,N_2292);
or U9125 (N_9125,N_109,N_3769);
nand U9126 (N_9126,N_1765,N_4244);
xor U9127 (N_9127,N_4224,N_1919);
and U9128 (N_9128,N_1878,N_895);
xor U9129 (N_9129,N_1104,N_3756);
nor U9130 (N_9130,N_857,N_3770);
and U9131 (N_9131,N_3497,N_1503);
or U9132 (N_9132,N_3232,N_3475);
nand U9133 (N_9133,N_1831,N_4752);
xnor U9134 (N_9134,N_4216,N_2811);
and U9135 (N_9135,N_3790,N_3911);
or U9136 (N_9136,N_1728,N_174);
xnor U9137 (N_9137,N_1598,N_1184);
and U9138 (N_9138,N_3415,N_231);
and U9139 (N_9139,N_541,N_1412);
and U9140 (N_9140,N_2935,N_4797);
nor U9141 (N_9141,N_4024,N_493);
or U9142 (N_9142,N_783,N_601);
or U9143 (N_9143,N_2622,N_1770);
or U9144 (N_9144,N_1203,N_2178);
and U9145 (N_9145,N_248,N_3869);
nor U9146 (N_9146,N_2276,N_2704);
and U9147 (N_9147,N_2336,N_679);
nor U9148 (N_9148,N_259,N_2870);
or U9149 (N_9149,N_3707,N_2791);
nor U9150 (N_9150,N_3455,N_2277);
nor U9151 (N_9151,N_4830,N_1123);
xnor U9152 (N_9152,N_4419,N_3128);
nor U9153 (N_9153,N_183,N_545);
nand U9154 (N_9154,N_2347,N_2884);
nand U9155 (N_9155,N_964,N_1295);
nand U9156 (N_9156,N_1944,N_3978);
nor U9157 (N_9157,N_816,N_1686);
and U9158 (N_9158,N_4876,N_3719);
and U9159 (N_9159,N_428,N_4384);
nor U9160 (N_9160,N_3456,N_1371);
nand U9161 (N_9161,N_2595,N_4925);
nor U9162 (N_9162,N_4152,N_4154);
or U9163 (N_9163,N_8,N_4098);
or U9164 (N_9164,N_3166,N_4415);
or U9165 (N_9165,N_1835,N_1043);
or U9166 (N_9166,N_834,N_1925);
or U9167 (N_9167,N_3380,N_4321);
and U9168 (N_9168,N_3575,N_3278);
nand U9169 (N_9169,N_4820,N_2935);
nor U9170 (N_9170,N_3105,N_3621);
xnor U9171 (N_9171,N_1041,N_4733);
xor U9172 (N_9172,N_4196,N_1673);
or U9173 (N_9173,N_827,N_15);
nand U9174 (N_9174,N_3825,N_3399);
or U9175 (N_9175,N_4678,N_1032);
or U9176 (N_9176,N_3897,N_2318);
nand U9177 (N_9177,N_4103,N_4304);
nand U9178 (N_9178,N_770,N_1386);
or U9179 (N_9179,N_4265,N_3276);
and U9180 (N_9180,N_3381,N_3583);
or U9181 (N_9181,N_1749,N_407);
nand U9182 (N_9182,N_3381,N_4678);
nand U9183 (N_9183,N_2737,N_170);
nand U9184 (N_9184,N_505,N_2416);
and U9185 (N_9185,N_4586,N_2043);
and U9186 (N_9186,N_3646,N_1759);
xor U9187 (N_9187,N_487,N_2082);
nor U9188 (N_9188,N_1115,N_256);
and U9189 (N_9189,N_458,N_4123);
nor U9190 (N_9190,N_3183,N_3350);
or U9191 (N_9191,N_3408,N_3421);
and U9192 (N_9192,N_529,N_3744);
nand U9193 (N_9193,N_4667,N_2973);
nor U9194 (N_9194,N_2268,N_1211);
nor U9195 (N_9195,N_3803,N_4904);
or U9196 (N_9196,N_2966,N_219);
nor U9197 (N_9197,N_2602,N_3934);
or U9198 (N_9198,N_2988,N_2890);
or U9199 (N_9199,N_2733,N_757);
and U9200 (N_9200,N_1154,N_2558);
nor U9201 (N_9201,N_769,N_2140);
or U9202 (N_9202,N_2110,N_4165);
or U9203 (N_9203,N_1574,N_72);
or U9204 (N_9204,N_4656,N_4836);
nand U9205 (N_9205,N_4760,N_2210);
xnor U9206 (N_9206,N_1484,N_1989);
nor U9207 (N_9207,N_4217,N_1378);
and U9208 (N_9208,N_1816,N_665);
nor U9209 (N_9209,N_1660,N_1364);
nor U9210 (N_9210,N_4094,N_4782);
nor U9211 (N_9211,N_4378,N_3534);
and U9212 (N_9212,N_3456,N_3847);
and U9213 (N_9213,N_4056,N_4979);
nor U9214 (N_9214,N_4865,N_3992);
nand U9215 (N_9215,N_2972,N_2667);
and U9216 (N_9216,N_2148,N_1600);
nor U9217 (N_9217,N_10,N_1275);
nand U9218 (N_9218,N_3914,N_2178);
and U9219 (N_9219,N_3864,N_2371);
or U9220 (N_9220,N_443,N_2318);
nand U9221 (N_9221,N_4891,N_424);
or U9222 (N_9222,N_913,N_1286);
and U9223 (N_9223,N_4873,N_1451);
nor U9224 (N_9224,N_4620,N_2089);
nand U9225 (N_9225,N_4260,N_4504);
nor U9226 (N_9226,N_324,N_1265);
xnor U9227 (N_9227,N_1895,N_3945);
xor U9228 (N_9228,N_4338,N_749);
nor U9229 (N_9229,N_0,N_1064);
xnor U9230 (N_9230,N_741,N_681);
nand U9231 (N_9231,N_4631,N_2830);
nor U9232 (N_9232,N_3806,N_1598);
or U9233 (N_9233,N_2988,N_3847);
or U9234 (N_9234,N_3677,N_807);
nand U9235 (N_9235,N_2427,N_3693);
and U9236 (N_9236,N_4751,N_3255);
or U9237 (N_9237,N_1493,N_2716);
xor U9238 (N_9238,N_4937,N_459);
nor U9239 (N_9239,N_3418,N_4509);
nor U9240 (N_9240,N_970,N_3032);
and U9241 (N_9241,N_3156,N_2686);
nor U9242 (N_9242,N_25,N_3081);
and U9243 (N_9243,N_4618,N_2568);
and U9244 (N_9244,N_1014,N_4246);
or U9245 (N_9245,N_1328,N_3372);
nand U9246 (N_9246,N_3638,N_2861);
and U9247 (N_9247,N_3802,N_121);
nor U9248 (N_9248,N_3803,N_2087);
nand U9249 (N_9249,N_4784,N_3248);
xor U9250 (N_9250,N_1001,N_29);
nand U9251 (N_9251,N_343,N_1903);
or U9252 (N_9252,N_293,N_4865);
nor U9253 (N_9253,N_991,N_4332);
xnor U9254 (N_9254,N_4471,N_4121);
nor U9255 (N_9255,N_3365,N_485);
xnor U9256 (N_9256,N_930,N_3051);
nand U9257 (N_9257,N_4034,N_1919);
or U9258 (N_9258,N_695,N_4447);
and U9259 (N_9259,N_4352,N_4380);
and U9260 (N_9260,N_1369,N_87);
nor U9261 (N_9261,N_3009,N_802);
nand U9262 (N_9262,N_2966,N_1585);
or U9263 (N_9263,N_202,N_923);
nor U9264 (N_9264,N_3121,N_1231);
nor U9265 (N_9265,N_1781,N_3307);
nand U9266 (N_9266,N_514,N_1670);
nor U9267 (N_9267,N_2122,N_3062);
nor U9268 (N_9268,N_2781,N_945);
nor U9269 (N_9269,N_3337,N_4847);
and U9270 (N_9270,N_4289,N_2640);
or U9271 (N_9271,N_941,N_4495);
xor U9272 (N_9272,N_2691,N_1473);
nand U9273 (N_9273,N_363,N_4537);
or U9274 (N_9274,N_100,N_1595);
nor U9275 (N_9275,N_2727,N_4907);
and U9276 (N_9276,N_367,N_14);
nand U9277 (N_9277,N_984,N_3929);
or U9278 (N_9278,N_3669,N_804);
nor U9279 (N_9279,N_2952,N_3725);
nor U9280 (N_9280,N_1810,N_181);
nand U9281 (N_9281,N_1123,N_302);
and U9282 (N_9282,N_2504,N_4568);
xor U9283 (N_9283,N_279,N_1860);
nor U9284 (N_9284,N_3412,N_1802);
and U9285 (N_9285,N_1368,N_3606);
nand U9286 (N_9286,N_2732,N_580);
nor U9287 (N_9287,N_4257,N_1002);
xnor U9288 (N_9288,N_3918,N_4324);
xnor U9289 (N_9289,N_3439,N_4546);
or U9290 (N_9290,N_41,N_2689);
or U9291 (N_9291,N_1347,N_4544);
and U9292 (N_9292,N_3433,N_4277);
nor U9293 (N_9293,N_946,N_2981);
nand U9294 (N_9294,N_4210,N_4943);
and U9295 (N_9295,N_2214,N_189);
nor U9296 (N_9296,N_2743,N_2069);
nor U9297 (N_9297,N_4630,N_2767);
or U9298 (N_9298,N_4315,N_3720);
nand U9299 (N_9299,N_2801,N_164);
or U9300 (N_9300,N_4569,N_3299);
nand U9301 (N_9301,N_4249,N_312);
nor U9302 (N_9302,N_1571,N_3789);
and U9303 (N_9303,N_3417,N_2548);
or U9304 (N_9304,N_637,N_4640);
or U9305 (N_9305,N_270,N_1276);
and U9306 (N_9306,N_672,N_2198);
xor U9307 (N_9307,N_3377,N_3667);
and U9308 (N_9308,N_4783,N_2404);
and U9309 (N_9309,N_3313,N_1272);
and U9310 (N_9310,N_2080,N_548);
nand U9311 (N_9311,N_1757,N_2903);
nor U9312 (N_9312,N_1485,N_2308);
xor U9313 (N_9313,N_2580,N_3335);
or U9314 (N_9314,N_3745,N_2764);
or U9315 (N_9315,N_3295,N_662);
nand U9316 (N_9316,N_1043,N_1061);
or U9317 (N_9317,N_4367,N_3986);
or U9318 (N_9318,N_4785,N_2455);
or U9319 (N_9319,N_4402,N_449);
and U9320 (N_9320,N_4044,N_4271);
xnor U9321 (N_9321,N_2152,N_4023);
or U9322 (N_9322,N_510,N_3585);
xor U9323 (N_9323,N_3690,N_3165);
or U9324 (N_9324,N_2174,N_1371);
nor U9325 (N_9325,N_4651,N_3157);
nand U9326 (N_9326,N_2616,N_2350);
and U9327 (N_9327,N_3374,N_4667);
nand U9328 (N_9328,N_4706,N_2270);
xor U9329 (N_9329,N_4940,N_6);
or U9330 (N_9330,N_4603,N_4104);
and U9331 (N_9331,N_2849,N_2671);
and U9332 (N_9332,N_3459,N_452);
or U9333 (N_9333,N_2179,N_534);
and U9334 (N_9334,N_4864,N_146);
or U9335 (N_9335,N_4055,N_2437);
nor U9336 (N_9336,N_2437,N_555);
nand U9337 (N_9337,N_596,N_3692);
nand U9338 (N_9338,N_4063,N_647);
nand U9339 (N_9339,N_2229,N_425);
and U9340 (N_9340,N_2393,N_4840);
nand U9341 (N_9341,N_4879,N_2321);
and U9342 (N_9342,N_39,N_3990);
nor U9343 (N_9343,N_2410,N_3088);
and U9344 (N_9344,N_2662,N_3515);
xor U9345 (N_9345,N_2962,N_3452);
nand U9346 (N_9346,N_976,N_2408);
or U9347 (N_9347,N_2760,N_1386);
and U9348 (N_9348,N_2381,N_105);
nand U9349 (N_9349,N_678,N_391);
nor U9350 (N_9350,N_2122,N_20);
nand U9351 (N_9351,N_169,N_4167);
or U9352 (N_9352,N_1701,N_2149);
nor U9353 (N_9353,N_203,N_4311);
nand U9354 (N_9354,N_4956,N_3149);
or U9355 (N_9355,N_4523,N_3100);
nand U9356 (N_9356,N_2879,N_445);
and U9357 (N_9357,N_1972,N_593);
nand U9358 (N_9358,N_3642,N_3744);
nor U9359 (N_9359,N_1738,N_2298);
nor U9360 (N_9360,N_2268,N_4531);
or U9361 (N_9361,N_1351,N_2329);
and U9362 (N_9362,N_2874,N_1580);
nor U9363 (N_9363,N_943,N_34);
nor U9364 (N_9364,N_2616,N_3259);
nand U9365 (N_9365,N_2509,N_4201);
and U9366 (N_9366,N_1077,N_1801);
xor U9367 (N_9367,N_1585,N_4704);
nor U9368 (N_9368,N_1357,N_2387);
and U9369 (N_9369,N_1821,N_2281);
and U9370 (N_9370,N_78,N_2300);
nand U9371 (N_9371,N_4340,N_1559);
and U9372 (N_9372,N_1975,N_3941);
nand U9373 (N_9373,N_2751,N_3725);
and U9374 (N_9374,N_3331,N_2636);
or U9375 (N_9375,N_3996,N_4296);
and U9376 (N_9376,N_4429,N_4532);
nor U9377 (N_9377,N_4401,N_352);
xnor U9378 (N_9378,N_4514,N_1002);
and U9379 (N_9379,N_217,N_830);
xnor U9380 (N_9380,N_2981,N_2355);
or U9381 (N_9381,N_2230,N_2600);
xnor U9382 (N_9382,N_1794,N_1494);
or U9383 (N_9383,N_910,N_3071);
and U9384 (N_9384,N_164,N_2469);
nor U9385 (N_9385,N_4611,N_502);
nor U9386 (N_9386,N_3138,N_909);
nand U9387 (N_9387,N_4935,N_2224);
xor U9388 (N_9388,N_3773,N_2632);
nor U9389 (N_9389,N_1571,N_3540);
nor U9390 (N_9390,N_414,N_983);
nand U9391 (N_9391,N_1626,N_2480);
nor U9392 (N_9392,N_2113,N_1458);
nand U9393 (N_9393,N_1889,N_2743);
nor U9394 (N_9394,N_2233,N_946);
and U9395 (N_9395,N_4845,N_87);
nand U9396 (N_9396,N_768,N_2879);
and U9397 (N_9397,N_3777,N_679);
nand U9398 (N_9398,N_590,N_2581);
nor U9399 (N_9399,N_4721,N_4695);
or U9400 (N_9400,N_3911,N_2127);
or U9401 (N_9401,N_3989,N_529);
nand U9402 (N_9402,N_1642,N_4424);
nor U9403 (N_9403,N_4914,N_2449);
nor U9404 (N_9404,N_4177,N_1555);
nor U9405 (N_9405,N_699,N_4085);
nor U9406 (N_9406,N_4112,N_4871);
and U9407 (N_9407,N_3618,N_4822);
or U9408 (N_9408,N_4448,N_4683);
nand U9409 (N_9409,N_2690,N_4993);
nor U9410 (N_9410,N_4363,N_3247);
nand U9411 (N_9411,N_282,N_3939);
nand U9412 (N_9412,N_4990,N_3552);
nand U9413 (N_9413,N_3043,N_3366);
or U9414 (N_9414,N_219,N_2004);
or U9415 (N_9415,N_4430,N_3806);
or U9416 (N_9416,N_4603,N_4897);
and U9417 (N_9417,N_4335,N_3327);
nor U9418 (N_9418,N_3143,N_3897);
and U9419 (N_9419,N_3703,N_3532);
nor U9420 (N_9420,N_1917,N_859);
nand U9421 (N_9421,N_3888,N_819);
nand U9422 (N_9422,N_2115,N_4431);
nand U9423 (N_9423,N_4935,N_902);
or U9424 (N_9424,N_3566,N_4467);
nor U9425 (N_9425,N_4447,N_2895);
xnor U9426 (N_9426,N_3443,N_882);
nor U9427 (N_9427,N_417,N_3182);
or U9428 (N_9428,N_3260,N_2312);
or U9429 (N_9429,N_234,N_2075);
xor U9430 (N_9430,N_2617,N_2911);
or U9431 (N_9431,N_3468,N_690);
nor U9432 (N_9432,N_1512,N_2557);
and U9433 (N_9433,N_2034,N_172);
or U9434 (N_9434,N_1694,N_2381);
nor U9435 (N_9435,N_2153,N_2432);
nand U9436 (N_9436,N_2968,N_1656);
and U9437 (N_9437,N_463,N_51);
and U9438 (N_9438,N_751,N_50);
or U9439 (N_9439,N_1400,N_3223);
and U9440 (N_9440,N_4350,N_1495);
or U9441 (N_9441,N_3901,N_4120);
or U9442 (N_9442,N_4739,N_1973);
nand U9443 (N_9443,N_1352,N_2184);
nor U9444 (N_9444,N_4655,N_4599);
or U9445 (N_9445,N_3801,N_2273);
nor U9446 (N_9446,N_3315,N_928);
nor U9447 (N_9447,N_953,N_3992);
and U9448 (N_9448,N_1682,N_4124);
and U9449 (N_9449,N_2972,N_2313);
nand U9450 (N_9450,N_1596,N_4315);
or U9451 (N_9451,N_2206,N_1183);
nor U9452 (N_9452,N_1897,N_3782);
and U9453 (N_9453,N_2533,N_2187);
nor U9454 (N_9454,N_2423,N_2400);
nor U9455 (N_9455,N_4277,N_1686);
xor U9456 (N_9456,N_1455,N_2143);
and U9457 (N_9457,N_4413,N_3247);
or U9458 (N_9458,N_4988,N_4262);
nand U9459 (N_9459,N_4348,N_4774);
nor U9460 (N_9460,N_3756,N_69);
and U9461 (N_9461,N_3175,N_54);
nand U9462 (N_9462,N_4329,N_2722);
or U9463 (N_9463,N_2236,N_126);
and U9464 (N_9464,N_3841,N_4468);
nor U9465 (N_9465,N_2511,N_3773);
nor U9466 (N_9466,N_3213,N_1720);
and U9467 (N_9467,N_2729,N_260);
and U9468 (N_9468,N_2709,N_2027);
nor U9469 (N_9469,N_4386,N_2834);
and U9470 (N_9470,N_1725,N_4790);
nor U9471 (N_9471,N_2674,N_2245);
or U9472 (N_9472,N_1480,N_444);
and U9473 (N_9473,N_1496,N_3612);
nor U9474 (N_9474,N_3243,N_4227);
nor U9475 (N_9475,N_4546,N_2108);
and U9476 (N_9476,N_3981,N_3360);
nor U9477 (N_9477,N_4328,N_1597);
nor U9478 (N_9478,N_82,N_4151);
and U9479 (N_9479,N_879,N_2152);
nand U9480 (N_9480,N_1778,N_2977);
nand U9481 (N_9481,N_3719,N_2109);
nand U9482 (N_9482,N_1135,N_3659);
or U9483 (N_9483,N_4756,N_938);
or U9484 (N_9484,N_1362,N_4059);
nor U9485 (N_9485,N_3049,N_1109);
nor U9486 (N_9486,N_1849,N_367);
nor U9487 (N_9487,N_378,N_2233);
or U9488 (N_9488,N_4761,N_3177);
or U9489 (N_9489,N_415,N_4999);
nor U9490 (N_9490,N_2374,N_2169);
and U9491 (N_9491,N_1428,N_354);
nand U9492 (N_9492,N_2706,N_1127);
nor U9493 (N_9493,N_1704,N_421);
nor U9494 (N_9494,N_2217,N_83);
or U9495 (N_9495,N_4878,N_22);
nor U9496 (N_9496,N_2818,N_3948);
or U9497 (N_9497,N_2299,N_4372);
or U9498 (N_9498,N_1855,N_2610);
and U9499 (N_9499,N_2578,N_4665);
nand U9500 (N_9500,N_2050,N_2826);
xor U9501 (N_9501,N_1573,N_2811);
nor U9502 (N_9502,N_4159,N_1243);
nand U9503 (N_9503,N_886,N_1369);
and U9504 (N_9504,N_4400,N_4784);
nor U9505 (N_9505,N_629,N_4014);
and U9506 (N_9506,N_3071,N_4980);
or U9507 (N_9507,N_3372,N_1724);
nor U9508 (N_9508,N_4469,N_1265);
nand U9509 (N_9509,N_4522,N_4787);
nor U9510 (N_9510,N_3764,N_4487);
nor U9511 (N_9511,N_824,N_4675);
xnor U9512 (N_9512,N_335,N_2348);
xor U9513 (N_9513,N_2152,N_3308);
and U9514 (N_9514,N_906,N_2358);
or U9515 (N_9515,N_4555,N_2430);
nor U9516 (N_9516,N_4721,N_4673);
nor U9517 (N_9517,N_902,N_4882);
or U9518 (N_9518,N_608,N_3661);
or U9519 (N_9519,N_4263,N_4912);
nand U9520 (N_9520,N_1455,N_3320);
xor U9521 (N_9521,N_4900,N_3841);
nand U9522 (N_9522,N_4185,N_880);
and U9523 (N_9523,N_324,N_2634);
or U9524 (N_9524,N_761,N_3524);
nor U9525 (N_9525,N_1608,N_4263);
or U9526 (N_9526,N_3699,N_2308);
nand U9527 (N_9527,N_1517,N_3770);
and U9528 (N_9528,N_1595,N_2732);
or U9529 (N_9529,N_2732,N_3693);
or U9530 (N_9530,N_4453,N_1590);
nor U9531 (N_9531,N_709,N_4253);
nor U9532 (N_9532,N_2590,N_4212);
and U9533 (N_9533,N_2338,N_3449);
nor U9534 (N_9534,N_152,N_1534);
xor U9535 (N_9535,N_1172,N_3408);
and U9536 (N_9536,N_1076,N_2162);
or U9537 (N_9537,N_2253,N_2901);
xnor U9538 (N_9538,N_595,N_1550);
and U9539 (N_9539,N_4099,N_844);
nand U9540 (N_9540,N_68,N_4622);
and U9541 (N_9541,N_3373,N_925);
nor U9542 (N_9542,N_4166,N_2646);
nand U9543 (N_9543,N_1120,N_4436);
xnor U9544 (N_9544,N_123,N_2760);
nor U9545 (N_9545,N_1968,N_1220);
or U9546 (N_9546,N_2311,N_2290);
or U9547 (N_9547,N_3669,N_4415);
or U9548 (N_9548,N_236,N_436);
nand U9549 (N_9549,N_1892,N_671);
nand U9550 (N_9550,N_1326,N_362);
and U9551 (N_9551,N_97,N_733);
or U9552 (N_9552,N_2842,N_7);
and U9553 (N_9553,N_573,N_2621);
and U9554 (N_9554,N_1320,N_1196);
xor U9555 (N_9555,N_1889,N_1951);
nor U9556 (N_9556,N_1051,N_1803);
nand U9557 (N_9557,N_282,N_2447);
nand U9558 (N_9558,N_3840,N_631);
xnor U9559 (N_9559,N_4958,N_2949);
nor U9560 (N_9560,N_1909,N_2497);
and U9561 (N_9561,N_2191,N_2433);
and U9562 (N_9562,N_1499,N_3650);
xor U9563 (N_9563,N_3772,N_2604);
nand U9564 (N_9564,N_1394,N_4298);
nand U9565 (N_9565,N_2595,N_4556);
or U9566 (N_9566,N_4225,N_2949);
nor U9567 (N_9567,N_1139,N_4770);
or U9568 (N_9568,N_2307,N_2937);
and U9569 (N_9569,N_740,N_2722);
nand U9570 (N_9570,N_1467,N_1400);
and U9571 (N_9571,N_3482,N_3091);
or U9572 (N_9572,N_2180,N_2215);
nand U9573 (N_9573,N_2516,N_2784);
or U9574 (N_9574,N_827,N_2414);
nor U9575 (N_9575,N_1620,N_559);
or U9576 (N_9576,N_3452,N_2996);
and U9577 (N_9577,N_3677,N_1718);
or U9578 (N_9578,N_4785,N_1821);
or U9579 (N_9579,N_543,N_4391);
or U9580 (N_9580,N_4939,N_2523);
nor U9581 (N_9581,N_1396,N_2678);
and U9582 (N_9582,N_4769,N_3458);
nor U9583 (N_9583,N_4090,N_873);
nor U9584 (N_9584,N_1784,N_3849);
nor U9585 (N_9585,N_3207,N_3251);
nand U9586 (N_9586,N_4467,N_23);
or U9587 (N_9587,N_4025,N_940);
xnor U9588 (N_9588,N_1495,N_3577);
nor U9589 (N_9589,N_341,N_1186);
nor U9590 (N_9590,N_3026,N_4286);
and U9591 (N_9591,N_3179,N_3919);
or U9592 (N_9592,N_1616,N_913);
xnor U9593 (N_9593,N_2178,N_642);
or U9594 (N_9594,N_3728,N_4871);
nand U9595 (N_9595,N_1848,N_2620);
or U9596 (N_9596,N_2679,N_2384);
nand U9597 (N_9597,N_1722,N_4783);
xor U9598 (N_9598,N_4227,N_3052);
nand U9599 (N_9599,N_4472,N_3635);
xor U9600 (N_9600,N_2706,N_3612);
nor U9601 (N_9601,N_4881,N_1529);
or U9602 (N_9602,N_1338,N_1155);
nor U9603 (N_9603,N_160,N_3165);
nand U9604 (N_9604,N_667,N_2226);
nor U9605 (N_9605,N_520,N_521);
nand U9606 (N_9606,N_4470,N_4994);
or U9607 (N_9607,N_3434,N_2535);
and U9608 (N_9608,N_472,N_1886);
nor U9609 (N_9609,N_973,N_2376);
or U9610 (N_9610,N_1564,N_3274);
or U9611 (N_9611,N_194,N_2192);
or U9612 (N_9612,N_3989,N_4470);
and U9613 (N_9613,N_1317,N_1574);
nor U9614 (N_9614,N_1829,N_3981);
and U9615 (N_9615,N_3575,N_2277);
nor U9616 (N_9616,N_864,N_2362);
and U9617 (N_9617,N_3237,N_1025);
nor U9618 (N_9618,N_3743,N_4407);
or U9619 (N_9619,N_286,N_4574);
or U9620 (N_9620,N_1051,N_4038);
or U9621 (N_9621,N_2137,N_1558);
xnor U9622 (N_9622,N_4050,N_2648);
nand U9623 (N_9623,N_391,N_3979);
nand U9624 (N_9624,N_3840,N_2606);
xnor U9625 (N_9625,N_1775,N_4471);
or U9626 (N_9626,N_1686,N_4861);
or U9627 (N_9627,N_3274,N_2369);
xnor U9628 (N_9628,N_3519,N_4153);
xnor U9629 (N_9629,N_3766,N_3998);
xnor U9630 (N_9630,N_140,N_4620);
nor U9631 (N_9631,N_1132,N_3506);
or U9632 (N_9632,N_883,N_1088);
nand U9633 (N_9633,N_609,N_1559);
or U9634 (N_9634,N_84,N_4547);
nand U9635 (N_9635,N_3050,N_2294);
or U9636 (N_9636,N_2,N_2953);
nor U9637 (N_9637,N_3080,N_4305);
nand U9638 (N_9638,N_1582,N_3509);
and U9639 (N_9639,N_270,N_4121);
nor U9640 (N_9640,N_3214,N_688);
or U9641 (N_9641,N_4220,N_2820);
nor U9642 (N_9642,N_1819,N_2057);
nor U9643 (N_9643,N_1277,N_201);
nor U9644 (N_9644,N_4918,N_4621);
and U9645 (N_9645,N_1429,N_2125);
nor U9646 (N_9646,N_3563,N_3607);
nand U9647 (N_9647,N_4141,N_2302);
nor U9648 (N_9648,N_2153,N_3709);
and U9649 (N_9649,N_3526,N_4054);
nor U9650 (N_9650,N_605,N_3955);
or U9651 (N_9651,N_213,N_4178);
or U9652 (N_9652,N_4909,N_18);
nand U9653 (N_9653,N_3632,N_2011);
xor U9654 (N_9654,N_1356,N_4073);
nor U9655 (N_9655,N_1262,N_3675);
xor U9656 (N_9656,N_3173,N_1926);
nand U9657 (N_9657,N_3691,N_1019);
or U9658 (N_9658,N_3159,N_2108);
xnor U9659 (N_9659,N_2535,N_612);
and U9660 (N_9660,N_1191,N_2005);
xor U9661 (N_9661,N_3265,N_3044);
nor U9662 (N_9662,N_3369,N_2518);
and U9663 (N_9663,N_4021,N_507);
or U9664 (N_9664,N_2792,N_2631);
nor U9665 (N_9665,N_4291,N_1455);
or U9666 (N_9666,N_3283,N_1368);
nor U9667 (N_9667,N_2798,N_2519);
nand U9668 (N_9668,N_139,N_2379);
and U9669 (N_9669,N_1939,N_511);
xor U9670 (N_9670,N_4302,N_1175);
and U9671 (N_9671,N_3684,N_2071);
nor U9672 (N_9672,N_4386,N_601);
nor U9673 (N_9673,N_493,N_2195);
and U9674 (N_9674,N_1452,N_4244);
nor U9675 (N_9675,N_4192,N_4120);
nand U9676 (N_9676,N_330,N_1840);
or U9677 (N_9677,N_2875,N_4226);
xor U9678 (N_9678,N_2330,N_4003);
nand U9679 (N_9679,N_3125,N_4483);
or U9680 (N_9680,N_1706,N_4046);
nor U9681 (N_9681,N_2553,N_2379);
and U9682 (N_9682,N_395,N_4233);
nor U9683 (N_9683,N_636,N_947);
nand U9684 (N_9684,N_2949,N_4390);
or U9685 (N_9685,N_2035,N_222);
and U9686 (N_9686,N_3620,N_2971);
nand U9687 (N_9687,N_2088,N_4679);
or U9688 (N_9688,N_3236,N_1520);
or U9689 (N_9689,N_3776,N_3544);
nand U9690 (N_9690,N_2348,N_2180);
xnor U9691 (N_9691,N_4554,N_485);
nor U9692 (N_9692,N_4145,N_303);
nand U9693 (N_9693,N_734,N_3228);
nand U9694 (N_9694,N_4565,N_3020);
xnor U9695 (N_9695,N_198,N_2039);
nand U9696 (N_9696,N_4911,N_2599);
nand U9697 (N_9697,N_950,N_1054);
and U9698 (N_9698,N_1573,N_1404);
nand U9699 (N_9699,N_1995,N_4973);
and U9700 (N_9700,N_697,N_2418);
nand U9701 (N_9701,N_414,N_619);
or U9702 (N_9702,N_1736,N_870);
or U9703 (N_9703,N_3362,N_1781);
xnor U9704 (N_9704,N_1744,N_901);
nor U9705 (N_9705,N_3186,N_3987);
xnor U9706 (N_9706,N_4855,N_3737);
and U9707 (N_9707,N_807,N_422);
nand U9708 (N_9708,N_1657,N_4219);
and U9709 (N_9709,N_3306,N_2997);
nor U9710 (N_9710,N_2767,N_974);
and U9711 (N_9711,N_1916,N_4253);
nand U9712 (N_9712,N_536,N_1608);
or U9713 (N_9713,N_3930,N_3090);
nor U9714 (N_9714,N_4093,N_2462);
or U9715 (N_9715,N_4693,N_3908);
and U9716 (N_9716,N_3035,N_1438);
or U9717 (N_9717,N_1172,N_4393);
and U9718 (N_9718,N_1154,N_1943);
or U9719 (N_9719,N_751,N_2858);
or U9720 (N_9720,N_3969,N_4082);
nor U9721 (N_9721,N_3459,N_3028);
nand U9722 (N_9722,N_3954,N_53);
and U9723 (N_9723,N_3745,N_2475);
nor U9724 (N_9724,N_2692,N_1173);
nor U9725 (N_9725,N_644,N_3762);
or U9726 (N_9726,N_3171,N_485);
nor U9727 (N_9727,N_4726,N_3056);
and U9728 (N_9728,N_1718,N_1756);
nor U9729 (N_9729,N_2382,N_2716);
nor U9730 (N_9730,N_4106,N_4487);
and U9731 (N_9731,N_1878,N_2333);
nand U9732 (N_9732,N_3650,N_3466);
nand U9733 (N_9733,N_1359,N_3155);
and U9734 (N_9734,N_4780,N_134);
xor U9735 (N_9735,N_3749,N_4671);
and U9736 (N_9736,N_194,N_1076);
nor U9737 (N_9737,N_2831,N_3168);
xnor U9738 (N_9738,N_3366,N_305);
nand U9739 (N_9739,N_4631,N_2135);
xnor U9740 (N_9740,N_2519,N_3821);
and U9741 (N_9741,N_558,N_3146);
and U9742 (N_9742,N_4131,N_3521);
nor U9743 (N_9743,N_2405,N_4006);
and U9744 (N_9744,N_876,N_1445);
nand U9745 (N_9745,N_158,N_1798);
nor U9746 (N_9746,N_335,N_1935);
xor U9747 (N_9747,N_2806,N_1694);
and U9748 (N_9748,N_2723,N_3488);
and U9749 (N_9749,N_4096,N_129);
or U9750 (N_9750,N_74,N_2942);
or U9751 (N_9751,N_1150,N_4952);
and U9752 (N_9752,N_3417,N_657);
and U9753 (N_9753,N_4304,N_2331);
nand U9754 (N_9754,N_3867,N_514);
xnor U9755 (N_9755,N_3606,N_3915);
nand U9756 (N_9756,N_685,N_3132);
or U9757 (N_9757,N_90,N_688);
or U9758 (N_9758,N_911,N_3414);
xor U9759 (N_9759,N_2473,N_3560);
and U9760 (N_9760,N_1445,N_1094);
or U9761 (N_9761,N_537,N_2951);
xor U9762 (N_9762,N_2299,N_4403);
or U9763 (N_9763,N_3924,N_2926);
and U9764 (N_9764,N_3229,N_4174);
nand U9765 (N_9765,N_1839,N_3691);
and U9766 (N_9766,N_3093,N_76);
xnor U9767 (N_9767,N_1354,N_550);
nor U9768 (N_9768,N_262,N_587);
xnor U9769 (N_9769,N_877,N_2700);
and U9770 (N_9770,N_3102,N_2046);
xor U9771 (N_9771,N_875,N_1832);
nor U9772 (N_9772,N_2356,N_1297);
nand U9773 (N_9773,N_2830,N_3629);
nand U9774 (N_9774,N_3595,N_3445);
and U9775 (N_9775,N_2796,N_1462);
nor U9776 (N_9776,N_2114,N_2691);
or U9777 (N_9777,N_2126,N_1391);
and U9778 (N_9778,N_1996,N_819);
and U9779 (N_9779,N_4595,N_3518);
and U9780 (N_9780,N_2780,N_619);
and U9781 (N_9781,N_4000,N_2336);
and U9782 (N_9782,N_1997,N_757);
xor U9783 (N_9783,N_67,N_2351);
nor U9784 (N_9784,N_354,N_3723);
nand U9785 (N_9785,N_3877,N_3565);
or U9786 (N_9786,N_4251,N_250);
nor U9787 (N_9787,N_4021,N_2935);
nor U9788 (N_9788,N_768,N_1299);
xnor U9789 (N_9789,N_4248,N_765);
and U9790 (N_9790,N_3879,N_1250);
and U9791 (N_9791,N_2273,N_3390);
nand U9792 (N_9792,N_2127,N_4585);
or U9793 (N_9793,N_1251,N_3886);
nor U9794 (N_9794,N_1819,N_1764);
nor U9795 (N_9795,N_2343,N_2385);
nor U9796 (N_9796,N_2015,N_2429);
or U9797 (N_9797,N_1878,N_2424);
nor U9798 (N_9798,N_2804,N_3271);
or U9799 (N_9799,N_1710,N_1834);
nand U9800 (N_9800,N_969,N_3475);
or U9801 (N_9801,N_2412,N_4437);
and U9802 (N_9802,N_38,N_2161);
nor U9803 (N_9803,N_2468,N_2152);
nor U9804 (N_9804,N_2777,N_3637);
or U9805 (N_9805,N_4412,N_2400);
xnor U9806 (N_9806,N_1300,N_2472);
or U9807 (N_9807,N_2653,N_2104);
nand U9808 (N_9808,N_1238,N_4996);
or U9809 (N_9809,N_3192,N_1606);
nand U9810 (N_9810,N_2106,N_1485);
and U9811 (N_9811,N_2933,N_3246);
nand U9812 (N_9812,N_4364,N_3262);
nor U9813 (N_9813,N_269,N_3955);
or U9814 (N_9814,N_4835,N_1041);
and U9815 (N_9815,N_563,N_1050);
nand U9816 (N_9816,N_907,N_3063);
nor U9817 (N_9817,N_2857,N_480);
or U9818 (N_9818,N_1881,N_956);
or U9819 (N_9819,N_4580,N_1499);
or U9820 (N_9820,N_3703,N_2912);
nor U9821 (N_9821,N_1958,N_380);
and U9822 (N_9822,N_666,N_665);
nor U9823 (N_9823,N_2325,N_1);
nand U9824 (N_9824,N_4064,N_2716);
xnor U9825 (N_9825,N_1985,N_626);
nor U9826 (N_9826,N_4680,N_4189);
nor U9827 (N_9827,N_4093,N_807);
or U9828 (N_9828,N_4111,N_3457);
and U9829 (N_9829,N_2756,N_3138);
nor U9830 (N_9830,N_4375,N_1109);
or U9831 (N_9831,N_4807,N_2078);
nor U9832 (N_9832,N_1408,N_1224);
or U9833 (N_9833,N_2912,N_709);
nor U9834 (N_9834,N_1216,N_4249);
nand U9835 (N_9835,N_979,N_2215);
nand U9836 (N_9836,N_4259,N_1745);
and U9837 (N_9837,N_3159,N_2537);
nor U9838 (N_9838,N_3402,N_685);
nand U9839 (N_9839,N_816,N_298);
and U9840 (N_9840,N_2749,N_4371);
nand U9841 (N_9841,N_4391,N_2148);
nor U9842 (N_9842,N_2063,N_1039);
and U9843 (N_9843,N_1253,N_2290);
or U9844 (N_9844,N_95,N_1673);
xor U9845 (N_9845,N_2372,N_2178);
xnor U9846 (N_9846,N_4843,N_1648);
nand U9847 (N_9847,N_2420,N_3204);
or U9848 (N_9848,N_4678,N_4470);
and U9849 (N_9849,N_1499,N_2928);
nand U9850 (N_9850,N_4683,N_1293);
and U9851 (N_9851,N_70,N_4047);
xor U9852 (N_9852,N_3167,N_4579);
nor U9853 (N_9853,N_1179,N_3634);
or U9854 (N_9854,N_2624,N_3150);
nand U9855 (N_9855,N_2121,N_1699);
or U9856 (N_9856,N_1163,N_359);
nor U9857 (N_9857,N_1295,N_1111);
nand U9858 (N_9858,N_1410,N_404);
and U9859 (N_9859,N_2629,N_3683);
and U9860 (N_9860,N_4568,N_4441);
nor U9861 (N_9861,N_62,N_4000);
and U9862 (N_9862,N_719,N_1130);
and U9863 (N_9863,N_1174,N_178);
nand U9864 (N_9864,N_1209,N_1153);
nor U9865 (N_9865,N_637,N_1362);
nand U9866 (N_9866,N_3766,N_2053);
nor U9867 (N_9867,N_1358,N_3593);
or U9868 (N_9868,N_3211,N_4573);
nand U9869 (N_9869,N_1380,N_916);
nand U9870 (N_9870,N_2093,N_916);
nor U9871 (N_9871,N_3190,N_2990);
nand U9872 (N_9872,N_4803,N_995);
or U9873 (N_9873,N_3989,N_1730);
and U9874 (N_9874,N_2387,N_2022);
and U9875 (N_9875,N_4120,N_939);
nand U9876 (N_9876,N_4927,N_252);
or U9877 (N_9877,N_3665,N_654);
xnor U9878 (N_9878,N_3740,N_2492);
nor U9879 (N_9879,N_4852,N_2857);
nor U9880 (N_9880,N_1374,N_1074);
nand U9881 (N_9881,N_4528,N_1286);
nor U9882 (N_9882,N_3364,N_352);
nor U9883 (N_9883,N_2245,N_3831);
nor U9884 (N_9884,N_25,N_1139);
and U9885 (N_9885,N_3072,N_4132);
nand U9886 (N_9886,N_3013,N_4633);
and U9887 (N_9887,N_4402,N_2314);
nand U9888 (N_9888,N_1985,N_1575);
and U9889 (N_9889,N_3655,N_1874);
nand U9890 (N_9890,N_2170,N_3757);
and U9891 (N_9891,N_1225,N_437);
nor U9892 (N_9892,N_4620,N_968);
nor U9893 (N_9893,N_1365,N_2004);
or U9894 (N_9894,N_493,N_4690);
and U9895 (N_9895,N_784,N_651);
nor U9896 (N_9896,N_2549,N_2568);
or U9897 (N_9897,N_2089,N_1296);
xor U9898 (N_9898,N_2843,N_2827);
and U9899 (N_9899,N_598,N_2661);
nand U9900 (N_9900,N_4988,N_958);
nand U9901 (N_9901,N_964,N_2146);
and U9902 (N_9902,N_891,N_4473);
or U9903 (N_9903,N_1658,N_996);
or U9904 (N_9904,N_1794,N_1206);
nor U9905 (N_9905,N_1334,N_750);
nand U9906 (N_9906,N_3995,N_2518);
nand U9907 (N_9907,N_3181,N_1534);
nand U9908 (N_9908,N_3366,N_1276);
nor U9909 (N_9909,N_4855,N_3065);
nand U9910 (N_9910,N_2651,N_881);
nor U9911 (N_9911,N_1246,N_2624);
and U9912 (N_9912,N_2678,N_98);
nand U9913 (N_9913,N_303,N_275);
nand U9914 (N_9914,N_1589,N_1460);
nand U9915 (N_9915,N_2076,N_3649);
nor U9916 (N_9916,N_405,N_615);
nor U9917 (N_9917,N_721,N_1610);
and U9918 (N_9918,N_1010,N_2808);
xor U9919 (N_9919,N_1251,N_3401);
and U9920 (N_9920,N_1846,N_3927);
nor U9921 (N_9921,N_1335,N_4644);
nor U9922 (N_9922,N_2026,N_1044);
nor U9923 (N_9923,N_2692,N_1896);
nand U9924 (N_9924,N_3955,N_3012);
nand U9925 (N_9925,N_4876,N_1941);
nor U9926 (N_9926,N_2876,N_4608);
nand U9927 (N_9927,N_4984,N_2122);
and U9928 (N_9928,N_4420,N_1179);
nand U9929 (N_9929,N_326,N_1802);
or U9930 (N_9930,N_4391,N_304);
nand U9931 (N_9931,N_3037,N_2066);
and U9932 (N_9932,N_89,N_2052);
xnor U9933 (N_9933,N_3992,N_1839);
nand U9934 (N_9934,N_2204,N_3642);
xnor U9935 (N_9935,N_520,N_4732);
and U9936 (N_9936,N_3024,N_3888);
or U9937 (N_9937,N_4014,N_2827);
or U9938 (N_9938,N_250,N_2531);
and U9939 (N_9939,N_900,N_501);
xor U9940 (N_9940,N_2174,N_3916);
and U9941 (N_9941,N_506,N_109);
nor U9942 (N_9942,N_3396,N_1449);
nand U9943 (N_9943,N_2813,N_4409);
xnor U9944 (N_9944,N_4038,N_1972);
xnor U9945 (N_9945,N_1641,N_1154);
nor U9946 (N_9946,N_3314,N_2656);
nand U9947 (N_9947,N_2634,N_923);
xor U9948 (N_9948,N_2699,N_4599);
nor U9949 (N_9949,N_3393,N_4222);
nand U9950 (N_9950,N_4332,N_3080);
and U9951 (N_9951,N_54,N_4448);
nand U9952 (N_9952,N_4463,N_2846);
and U9953 (N_9953,N_3020,N_2099);
or U9954 (N_9954,N_2917,N_2475);
nor U9955 (N_9955,N_3221,N_106);
nand U9956 (N_9956,N_3174,N_4532);
nand U9957 (N_9957,N_3308,N_4433);
nand U9958 (N_9958,N_3851,N_3664);
or U9959 (N_9959,N_3540,N_1142);
or U9960 (N_9960,N_1602,N_2519);
nor U9961 (N_9961,N_2646,N_1943);
or U9962 (N_9962,N_1789,N_2904);
xnor U9963 (N_9963,N_4431,N_2670);
or U9964 (N_9964,N_3900,N_4332);
and U9965 (N_9965,N_2034,N_1110);
and U9966 (N_9966,N_1255,N_2358);
or U9967 (N_9967,N_1317,N_4326);
nand U9968 (N_9968,N_1264,N_4398);
nor U9969 (N_9969,N_2707,N_2170);
nor U9970 (N_9970,N_3815,N_4301);
nor U9971 (N_9971,N_2907,N_4874);
xor U9972 (N_9972,N_22,N_1210);
xor U9973 (N_9973,N_657,N_4537);
or U9974 (N_9974,N_2757,N_1248);
nand U9975 (N_9975,N_1379,N_3330);
nand U9976 (N_9976,N_3194,N_4421);
or U9977 (N_9977,N_622,N_3040);
nor U9978 (N_9978,N_4886,N_388);
and U9979 (N_9979,N_3363,N_978);
nor U9980 (N_9980,N_4778,N_2566);
nor U9981 (N_9981,N_2635,N_2746);
nand U9982 (N_9982,N_4047,N_715);
or U9983 (N_9983,N_4504,N_563);
or U9984 (N_9984,N_613,N_2159);
and U9985 (N_9985,N_1349,N_3239);
and U9986 (N_9986,N_4314,N_173);
or U9987 (N_9987,N_3167,N_4778);
xnor U9988 (N_9988,N_3016,N_571);
nand U9989 (N_9989,N_3282,N_2342);
nand U9990 (N_9990,N_360,N_4358);
or U9991 (N_9991,N_1140,N_771);
and U9992 (N_9992,N_3532,N_357);
or U9993 (N_9993,N_1773,N_3540);
or U9994 (N_9994,N_2164,N_3680);
nand U9995 (N_9995,N_3894,N_1868);
or U9996 (N_9996,N_3335,N_217);
xnor U9997 (N_9997,N_3776,N_4587);
or U9998 (N_9998,N_4533,N_2386);
nor U9999 (N_9999,N_1689,N_3371);
or UO_0 (O_0,N_7573,N_9592);
nor UO_1 (O_1,N_6576,N_9412);
nand UO_2 (O_2,N_5773,N_7355);
xnor UO_3 (O_3,N_5466,N_9844);
nor UO_4 (O_4,N_5980,N_5560);
nand UO_5 (O_5,N_5549,N_7463);
or UO_6 (O_6,N_8580,N_6293);
or UO_7 (O_7,N_6303,N_8966);
nand UO_8 (O_8,N_7228,N_5403);
xor UO_9 (O_9,N_5639,N_8815);
nor UO_10 (O_10,N_6540,N_5760);
and UO_11 (O_11,N_9362,N_8456);
and UO_12 (O_12,N_8292,N_5534);
and UO_13 (O_13,N_6212,N_5424);
nor UO_14 (O_14,N_8732,N_7434);
nor UO_15 (O_15,N_6799,N_7557);
or UO_16 (O_16,N_9021,N_7691);
nor UO_17 (O_17,N_7665,N_9519);
or UO_18 (O_18,N_5201,N_5046);
nand UO_19 (O_19,N_7795,N_8858);
or UO_20 (O_20,N_8667,N_9901);
nand UO_21 (O_21,N_6294,N_5766);
nor UO_22 (O_22,N_7874,N_9690);
nor UO_23 (O_23,N_9753,N_8984);
nand UO_24 (O_24,N_7252,N_7366);
or UO_25 (O_25,N_6397,N_6705);
or UO_26 (O_26,N_6048,N_5938);
nor UO_27 (O_27,N_9577,N_9777);
nand UO_28 (O_28,N_8268,N_7596);
and UO_29 (O_29,N_6913,N_6845);
or UO_30 (O_30,N_6331,N_9167);
nand UO_31 (O_31,N_9434,N_8397);
or UO_32 (O_32,N_6472,N_9672);
and UO_33 (O_33,N_8560,N_6876);
nor UO_34 (O_34,N_9758,N_7696);
nand UO_35 (O_35,N_8626,N_8242);
and UO_36 (O_36,N_6569,N_5790);
or UO_37 (O_37,N_5241,N_9032);
and UO_38 (O_38,N_8431,N_6762);
nand UO_39 (O_39,N_5693,N_8440);
nor UO_40 (O_40,N_5996,N_7266);
nand UO_41 (O_41,N_6050,N_9963);
xnor UO_42 (O_42,N_8131,N_9416);
nor UO_43 (O_43,N_8750,N_5956);
or UO_44 (O_44,N_7818,N_8552);
xnor UO_45 (O_45,N_8880,N_6942);
and UO_46 (O_46,N_8518,N_8155);
and UO_47 (O_47,N_6579,N_5574);
and UO_48 (O_48,N_8150,N_5284);
or UO_49 (O_49,N_7002,N_8374);
and UO_50 (O_50,N_9917,N_7808);
xnor UO_51 (O_51,N_8078,N_5465);
nand UO_52 (O_52,N_7896,N_8490);
or UO_53 (O_53,N_5145,N_7230);
xor UO_54 (O_54,N_9875,N_9841);
or UO_55 (O_55,N_7381,N_8970);
nand UO_56 (O_56,N_6730,N_8668);
and UO_57 (O_57,N_7531,N_7423);
nor UO_58 (O_58,N_5249,N_7607);
xnor UO_59 (O_59,N_6284,N_9809);
or UO_60 (O_60,N_8583,N_7673);
or UO_61 (O_61,N_5017,N_5669);
or UO_62 (O_62,N_5304,N_5985);
or UO_63 (O_63,N_7922,N_7858);
and UO_64 (O_64,N_9092,N_6073);
and UO_65 (O_65,N_5454,N_8915);
and UO_66 (O_66,N_5666,N_6884);
nor UO_67 (O_67,N_5504,N_9977);
nor UO_68 (O_68,N_9517,N_5372);
and UO_69 (O_69,N_8751,N_8376);
nor UO_70 (O_70,N_5271,N_9569);
xor UO_71 (O_71,N_8383,N_5353);
nor UO_72 (O_72,N_7444,N_8158);
nand UO_73 (O_73,N_9624,N_9198);
or UO_74 (O_74,N_7403,N_6153);
and UO_75 (O_75,N_9242,N_6800);
nand UO_76 (O_76,N_7625,N_6249);
nand UO_77 (O_77,N_6451,N_9575);
nand UO_78 (O_78,N_8843,N_6424);
xnor UO_79 (O_79,N_8344,N_6588);
xor UO_80 (O_80,N_7130,N_9546);
nand UO_81 (O_81,N_9216,N_7387);
and UO_82 (O_82,N_6492,N_6128);
nand UO_83 (O_83,N_6805,N_7420);
and UO_84 (O_84,N_7297,N_7905);
and UO_85 (O_85,N_6826,N_6182);
nor UO_86 (O_86,N_9587,N_8914);
nor UO_87 (O_87,N_9573,N_8845);
and UO_88 (O_88,N_8188,N_5675);
xor UO_89 (O_89,N_9541,N_5858);
nor UO_90 (O_90,N_9887,N_6644);
and UO_91 (O_91,N_5463,N_8982);
xnor UO_92 (O_92,N_6046,N_7008);
and UO_93 (O_93,N_6109,N_7658);
and UO_94 (O_94,N_6785,N_8405);
nand UO_95 (O_95,N_8128,N_8076);
or UO_96 (O_96,N_5100,N_6161);
and UO_97 (O_97,N_5570,N_8235);
and UO_98 (O_98,N_6621,N_5280);
or UO_99 (O_99,N_7452,N_5678);
or UO_100 (O_100,N_9561,N_7789);
or UO_101 (O_101,N_7532,N_6803);
and UO_102 (O_102,N_8800,N_9655);
or UO_103 (O_103,N_8233,N_9469);
and UO_104 (O_104,N_5195,N_9181);
and UO_105 (O_105,N_7398,N_9872);
xor UO_106 (O_106,N_7097,N_7271);
nand UO_107 (O_107,N_5116,N_9568);
nand UO_108 (O_108,N_8429,N_8752);
or UO_109 (O_109,N_9554,N_5761);
and UO_110 (O_110,N_8247,N_9123);
nand UO_111 (O_111,N_9124,N_6502);
or UO_112 (O_112,N_6598,N_8735);
or UO_113 (O_113,N_5544,N_6572);
or UO_114 (O_114,N_8253,N_7268);
nor UO_115 (O_115,N_9421,N_6666);
and UO_116 (O_116,N_7346,N_7904);
nor UO_117 (O_117,N_7357,N_8399);
nor UO_118 (O_118,N_9333,N_5878);
nand UO_119 (O_119,N_8336,N_7809);
nor UO_120 (O_120,N_8491,N_7273);
and UO_121 (O_121,N_8236,N_6707);
or UO_122 (O_122,N_7305,N_7556);
xor UO_123 (O_123,N_7251,N_7016);
xor UO_124 (O_124,N_9090,N_7383);
or UO_125 (O_125,N_5419,N_6748);
xor UO_126 (O_126,N_5697,N_8756);
nand UO_127 (O_127,N_9368,N_9154);
xnor UO_128 (O_128,N_7920,N_9492);
nor UO_129 (O_129,N_9526,N_6524);
nor UO_130 (O_130,N_5876,N_7421);
nor UO_131 (O_131,N_6361,N_9889);
or UO_132 (O_132,N_7830,N_5112);
or UO_133 (O_133,N_8093,N_8838);
nor UO_134 (O_134,N_7000,N_7248);
and UO_135 (O_135,N_6980,N_6699);
nor UO_136 (O_136,N_8266,N_9023);
nand UO_137 (O_137,N_8444,N_9865);
nor UO_138 (O_138,N_5070,N_7616);
nand UO_139 (O_139,N_5684,N_5621);
xor UO_140 (O_140,N_8115,N_5422);
nor UO_141 (O_141,N_9497,N_9044);
xnor UO_142 (O_142,N_9941,N_9419);
nand UO_143 (O_143,N_9952,N_6671);
nor UO_144 (O_144,N_5873,N_9629);
or UO_145 (O_145,N_9811,N_5257);
xnor UO_146 (O_146,N_8390,N_9418);
nor UO_147 (O_147,N_7453,N_9539);
nor UO_148 (O_148,N_5486,N_9449);
or UO_149 (O_149,N_8103,N_9328);
and UO_150 (O_150,N_8010,N_8563);
or UO_151 (O_151,N_5740,N_9009);
or UO_152 (O_152,N_6947,N_8711);
nand UO_153 (O_153,N_8156,N_9504);
xor UO_154 (O_154,N_7354,N_6896);
and UO_155 (O_155,N_6774,N_8946);
nor UO_156 (O_156,N_7688,N_5916);
xnor UO_157 (O_157,N_8492,N_6861);
and UO_158 (O_158,N_5964,N_5412);
nor UO_159 (O_159,N_9191,N_9454);
nand UO_160 (O_160,N_7635,N_6713);
xnor UO_161 (O_161,N_9398,N_6647);
and UO_162 (O_162,N_8738,N_8195);
nor UO_163 (O_163,N_7497,N_5700);
or UO_164 (O_164,N_7417,N_9475);
and UO_165 (O_165,N_8484,N_9354);
nand UO_166 (O_166,N_8960,N_6346);
or UO_167 (O_167,N_9357,N_7860);
and UO_168 (O_168,N_8544,N_9289);
nor UO_169 (O_169,N_6304,N_5126);
nand UO_170 (O_170,N_9894,N_5138);
xor UO_171 (O_171,N_5188,N_5521);
nor UO_172 (O_172,N_9721,N_6696);
nor UO_173 (O_173,N_9282,N_7265);
and UO_174 (O_174,N_5437,N_6464);
or UO_175 (O_175,N_6404,N_7154);
or UO_176 (O_176,N_5727,N_7773);
nor UO_177 (O_177,N_8923,N_7027);
nand UO_178 (O_178,N_8486,N_9177);
nor UO_179 (O_179,N_8203,N_8455);
nand UO_180 (O_180,N_7917,N_7060);
nand UO_181 (O_181,N_5459,N_9819);
or UO_182 (O_182,N_8113,N_7745);
nand UO_183 (O_183,N_8574,N_8039);
nand UO_184 (O_184,N_6963,N_8004);
nand UO_185 (O_185,N_8821,N_5871);
or UO_186 (O_186,N_9866,N_8092);
and UO_187 (O_187,N_5345,N_8650);
xnor UO_188 (O_188,N_7024,N_9430);
nor UO_189 (O_189,N_6401,N_5842);
nor UO_190 (O_190,N_8331,N_5900);
or UO_191 (O_191,N_5680,N_6801);
or UO_192 (O_192,N_8187,N_9004);
xor UO_193 (O_193,N_8290,N_8833);
or UO_194 (O_194,N_6120,N_6151);
or UO_195 (O_195,N_7173,N_5452);
or UO_196 (O_196,N_9468,N_8931);
xnor UO_197 (O_197,N_6454,N_6243);
nand UO_198 (O_198,N_9765,N_9869);
nor UO_199 (O_199,N_9516,N_6829);
nand UO_200 (O_200,N_6717,N_8197);
or UO_201 (O_201,N_5154,N_7065);
or UO_202 (O_202,N_8505,N_7469);
or UO_203 (O_203,N_9604,N_9807);
and UO_204 (O_204,N_9723,N_7361);
and UO_205 (O_205,N_5067,N_8927);
nand UO_206 (O_206,N_9850,N_7036);
nor UO_207 (O_207,N_8066,N_9296);
or UO_208 (O_208,N_5069,N_5969);
nand UO_209 (O_209,N_6751,N_8214);
and UO_210 (O_210,N_5519,N_7327);
or UO_211 (O_211,N_7992,N_6652);
and UO_212 (O_212,N_7648,N_6733);
nand UO_213 (O_213,N_6635,N_9729);
xor UO_214 (O_214,N_9020,N_6378);
xor UO_215 (O_215,N_8705,N_5009);
or UO_216 (O_216,N_5782,N_7059);
nand UO_217 (O_217,N_9543,N_5594);
and UO_218 (O_218,N_7956,N_8285);
nor UO_219 (O_219,N_7140,N_9073);
and UO_220 (O_220,N_9520,N_7736);
xnor UO_221 (O_221,N_9613,N_5494);
or UO_222 (O_222,N_9898,N_7316);
or UO_223 (O_223,N_5614,N_9037);
nand UO_224 (O_224,N_5984,N_5897);
nor UO_225 (O_225,N_6993,N_9332);
nand UO_226 (O_226,N_5142,N_5894);
nand UO_227 (O_227,N_6849,N_7261);
or UO_228 (O_228,N_7334,N_7516);
or UO_229 (O_229,N_9472,N_5475);
or UO_230 (O_230,N_5895,N_8703);
nor UO_231 (O_231,N_9523,N_6069);
nand UO_232 (O_232,N_6405,N_7149);
xnor UO_233 (O_233,N_9771,N_5240);
nor UO_234 (O_234,N_6836,N_5840);
and UO_235 (O_235,N_6247,N_6632);
nor UO_236 (O_236,N_9265,N_5268);
or UO_237 (O_237,N_5690,N_7982);
or UO_238 (O_238,N_9638,N_7239);
nor UO_239 (O_239,N_8812,N_9432);
or UO_240 (O_240,N_9698,N_7602);
and UO_241 (O_241,N_8787,N_9025);
or UO_242 (O_242,N_6515,N_7600);
nand UO_243 (O_243,N_7178,N_5137);
nor UO_244 (O_244,N_7284,N_9040);
and UO_245 (O_245,N_5714,N_8325);
or UO_246 (O_246,N_9433,N_9578);
or UO_247 (O_247,N_6633,N_7037);
and UO_248 (O_248,N_5342,N_6364);
xor UO_249 (O_249,N_5397,N_9682);
nand UO_250 (O_250,N_5904,N_9708);
nand UO_251 (O_251,N_8428,N_8322);
or UO_252 (O_252,N_6608,N_6692);
and UO_253 (O_253,N_6535,N_5883);
xor UO_254 (O_254,N_6140,N_5815);
nor UO_255 (O_255,N_6710,N_8863);
or UO_256 (O_256,N_6289,N_7610);
nand UO_257 (O_257,N_7462,N_7219);
nor UO_258 (O_258,N_8291,N_8170);
nand UO_259 (O_259,N_6606,N_9784);
xnor UO_260 (O_260,N_6352,N_5538);
nor UO_261 (O_261,N_7539,N_8145);
or UO_262 (O_262,N_5363,N_7898);
or UO_263 (O_263,N_6139,N_9895);
nor UO_264 (O_264,N_8001,N_6010);
and UO_265 (O_265,N_5355,N_6573);
xnor UO_266 (O_266,N_7916,N_9770);
nor UO_267 (O_267,N_9407,N_9864);
or UO_268 (O_268,N_5712,N_8938);
and UO_269 (O_269,N_5183,N_9923);
and UO_270 (O_270,N_8656,N_7427);
or UO_271 (O_271,N_6125,N_8301);
xor UO_272 (O_272,N_7519,N_7805);
or UO_273 (O_273,N_7985,N_8709);
or UO_274 (O_274,N_5705,N_9046);
and UO_275 (O_275,N_8987,N_5857);
nor UO_276 (O_276,N_5741,N_8245);
and UO_277 (O_277,N_8745,N_9813);
and UO_278 (O_278,N_8141,N_5199);
nor UO_279 (O_279,N_8215,N_7363);
or UO_280 (O_280,N_5434,N_7225);
nor UO_281 (O_281,N_8388,N_8925);
and UO_282 (O_282,N_9944,N_7578);
or UO_283 (O_283,N_7994,N_8171);
and UO_284 (O_284,N_9462,N_7548);
or UO_285 (O_285,N_8442,N_5331);
and UO_286 (O_286,N_8207,N_8201);
nor UO_287 (O_287,N_7437,N_9590);
nor UO_288 (O_288,N_8252,N_7416);
nor UO_289 (O_289,N_9661,N_6037);
xnor UO_290 (O_290,N_8597,N_8144);
xnor UO_291 (O_291,N_6879,N_5719);
or UO_292 (O_292,N_6034,N_8133);
nor UO_293 (O_293,N_5512,N_6366);
nor UO_294 (O_294,N_8448,N_9217);
and UO_295 (O_295,N_6316,N_9769);
and UO_296 (O_296,N_5503,N_9755);
or UO_297 (O_297,N_9063,N_7522);
nor UO_298 (O_298,N_7972,N_6886);
nand UO_299 (O_299,N_6827,N_7472);
and UO_300 (O_300,N_5523,N_6484);
nor UO_301 (O_301,N_8818,N_5367);
nor UO_302 (O_302,N_8269,N_7496);
and UO_303 (O_303,N_9065,N_7201);
nand UO_304 (O_304,N_7717,N_9616);
nor UO_305 (O_305,N_5843,N_8157);
xor UO_306 (O_306,N_7580,N_8083);
nor UO_307 (O_307,N_8657,N_8166);
xor UO_308 (O_308,N_6994,N_6015);
xor UO_309 (O_309,N_6816,N_8808);
and UO_310 (O_310,N_9609,N_8872);
or UO_311 (O_311,N_7103,N_5561);
or UO_312 (O_312,N_7598,N_7957);
nand UO_313 (O_313,N_7570,N_9294);
nand UO_314 (O_314,N_8515,N_9318);
or UO_315 (O_315,N_9350,N_9595);
and UO_316 (O_316,N_7095,N_9269);
or UO_317 (O_317,N_8953,N_6244);
or UO_318 (O_318,N_9696,N_7618);
nand UO_319 (O_319,N_7353,N_6967);
nor UO_320 (O_320,N_9082,N_5979);
or UO_321 (O_321,N_5730,N_6757);
and UO_322 (O_322,N_8708,N_6081);
or UO_323 (O_323,N_7202,N_7442);
xor UO_324 (O_324,N_9766,N_5636);
nand UO_325 (O_325,N_6866,N_7200);
or UO_326 (O_326,N_6074,N_6216);
or UO_327 (O_327,N_7128,N_9319);
nor UO_328 (O_328,N_7685,N_7198);
xor UO_329 (O_329,N_8878,N_6523);
or UO_330 (O_330,N_5432,N_8786);
xor UO_331 (O_331,N_6900,N_9501);
xnor UO_332 (O_332,N_5168,N_7571);
nor UO_333 (O_333,N_7350,N_7919);
and UO_334 (O_334,N_6122,N_9972);
xnor UO_335 (O_335,N_8571,N_9863);
or UO_336 (O_336,N_6097,N_5299);
nand UO_337 (O_337,N_9103,N_5307);
or UO_338 (O_338,N_5094,N_9165);
and UO_339 (O_339,N_6927,N_7788);
nand UO_340 (O_340,N_6204,N_9626);
and UO_341 (O_341,N_6152,N_9104);
nand UO_342 (O_342,N_5706,N_8487);
nand UO_343 (O_343,N_6475,N_7454);
nor UO_344 (O_344,N_5735,N_9584);
and UO_345 (O_345,N_9600,N_6077);
nand UO_346 (O_346,N_5943,N_9618);
nand UO_347 (O_347,N_5566,N_6334);
nand UO_348 (O_348,N_7689,N_6257);
nor UO_349 (O_349,N_6237,N_6144);
and UO_350 (O_350,N_5767,N_8606);
or UO_351 (O_351,N_9994,N_5357);
nor UO_352 (O_352,N_8387,N_5295);
nor UO_353 (O_353,N_9078,N_5877);
or UO_354 (O_354,N_7647,N_8741);
nor UO_355 (O_355,N_6301,N_5598);
and UO_356 (O_356,N_6426,N_5568);
and UO_357 (O_357,N_5071,N_6400);
nand UO_358 (O_358,N_6670,N_5011);
or UO_359 (O_359,N_6483,N_5981);
nand UO_360 (O_360,N_5186,N_5948);
or UO_361 (O_361,N_9947,N_8476);
nor UO_362 (O_362,N_9936,N_8189);
or UO_363 (O_363,N_7599,N_7033);
or UO_364 (O_364,N_7400,N_5388);
and UO_365 (O_365,N_7976,N_7915);
or UO_366 (O_366,N_5132,N_7303);
xor UO_367 (O_367,N_7123,N_9463);
and UO_368 (O_368,N_9133,N_6350);
and UO_369 (O_369,N_5844,N_5202);
and UO_370 (O_370,N_7500,N_5149);
nand UO_371 (O_371,N_5772,N_8485);
or UO_372 (O_372,N_9137,N_6558);
nor UO_373 (O_373,N_6488,N_5276);
xor UO_374 (O_374,N_5330,N_6353);
and UO_375 (O_375,N_7545,N_7295);
nor UO_376 (O_376,N_6834,N_8542);
or UO_377 (O_377,N_7164,N_8805);
nand UO_378 (O_378,N_7465,N_9843);
and UO_379 (O_379,N_6051,N_6888);
and UO_380 (O_380,N_8177,N_7953);
nor UO_381 (O_381,N_8934,N_9744);
nor UO_382 (O_382,N_9635,N_5516);
nand UO_383 (O_383,N_5286,N_8472);
nor UO_384 (O_384,N_7755,N_6663);
nand UO_385 (O_385,N_7166,N_9387);
nand UO_386 (O_386,N_5525,N_9695);
nand UO_387 (O_387,N_5370,N_6170);
xnor UO_388 (O_388,N_9234,N_8666);
or UO_389 (O_389,N_8883,N_6448);
or UO_390 (O_390,N_9808,N_5489);
and UO_391 (O_391,N_7241,N_5151);
nand UO_392 (O_392,N_7418,N_8308);
and UO_393 (O_393,N_6675,N_6700);
nor UO_394 (O_394,N_6466,N_8416);
nand UO_395 (O_395,N_5128,N_7006);
nand UO_396 (O_396,N_8225,N_9852);
or UO_397 (O_397,N_8949,N_7478);
or UO_398 (O_398,N_7209,N_7988);
nor UO_399 (O_399,N_6683,N_9127);
and UO_400 (O_400,N_6597,N_8964);
xor UO_401 (O_401,N_8641,N_6593);
nand UO_402 (O_402,N_9916,N_7924);
and UO_403 (O_403,N_9185,N_5415);
nand UO_404 (O_404,N_7388,N_6842);
nor UO_405 (O_405,N_6920,N_5477);
xnor UO_406 (O_406,N_8935,N_6937);
and UO_407 (O_407,N_7111,N_8605);
and UO_408 (O_408,N_6735,N_8817);
and UO_409 (O_409,N_6808,N_9417);
nor UO_410 (O_410,N_6681,N_9679);
and UO_411 (O_411,N_8495,N_8098);
nand UO_412 (O_412,N_9288,N_8993);
nor UO_413 (O_413,N_7391,N_9444);
or UO_414 (O_414,N_8299,N_7009);
and UO_415 (O_415,N_7018,N_5034);
or UO_416 (O_416,N_7608,N_8768);
and UO_417 (O_417,N_9344,N_9161);
nand UO_418 (O_418,N_5165,N_9945);
or UO_419 (O_419,N_5292,N_7526);
or UO_420 (O_420,N_9759,N_8613);
or UO_421 (O_421,N_8856,N_5492);
nand UO_422 (O_422,N_8697,N_5309);
xor UO_423 (O_423,N_5234,N_7812);
nor UO_424 (O_424,N_8929,N_6299);
or UO_425 (O_425,N_8226,N_6324);
and UO_426 (O_426,N_5927,N_8704);
nor UO_427 (O_427,N_9183,N_9612);
nor UO_428 (O_428,N_7412,N_5421);
xor UO_429 (O_429,N_6601,N_5708);
nand UO_430 (O_430,N_8355,N_8223);
and UO_431 (O_431,N_8955,N_8579);
and UO_432 (O_432,N_5449,N_9839);
nor UO_433 (O_433,N_9408,N_9663);
or UO_434 (O_434,N_7029,N_9173);
nand UO_435 (O_435,N_7096,N_6714);
or UO_436 (O_436,N_6636,N_7969);
xor UO_437 (O_437,N_8734,N_6848);
nor UO_438 (O_438,N_6004,N_9622);
or UO_439 (O_439,N_6242,N_7550);
and UO_440 (O_440,N_9607,N_6723);
and UO_441 (O_441,N_8213,N_5796);
nand UO_442 (O_442,N_7214,N_8576);
nor UO_443 (O_443,N_5721,N_5395);
nor UO_444 (O_444,N_9231,N_9488);
and UO_445 (O_445,N_6877,N_7072);
nor UO_446 (O_446,N_5798,N_7101);
nand UO_447 (O_447,N_6038,N_6755);
nand UO_448 (O_448,N_5929,N_8210);
nand UO_449 (O_449,N_8680,N_8632);
and UO_450 (O_450,N_7039,N_7410);
or UO_451 (O_451,N_9473,N_6371);
nand UO_452 (O_452,N_5349,N_8413);
or UO_453 (O_453,N_5317,N_6337);
nand UO_454 (O_454,N_5170,N_8452);
nand UO_455 (O_455,N_7504,N_6889);
and UO_456 (O_456,N_6473,N_9693);
nand UO_457 (O_457,N_7160,N_7893);
and UO_458 (O_458,N_9598,N_9404);
nand UO_459 (O_459,N_7035,N_8143);
and UO_460 (O_460,N_6115,N_8531);
or UO_461 (O_461,N_9837,N_6129);
nor UO_462 (O_462,N_7141,N_6689);
or UO_463 (O_463,N_5599,N_9658);
and UO_464 (O_464,N_5264,N_9971);
xor UO_465 (O_465,N_9712,N_9779);
or UO_466 (O_466,N_7306,N_6162);
nor UO_467 (O_467,N_5113,N_8204);
nand UO_468 (O_468,N_7369,N_6163);
or UO_469 (O_469,N_5676,N_5756);
nand UO_470 (O_470,N_6266,N_9527);
nor UO_471 (O_471,N_8081,N_9995);
or UO_472 (O_472,N_7576,N_5872);
xor UO_473 (O_473,N_6584,N_9532);
nor UO_474 (O_474,N_7014,N_9414);
and UO_475 (O_475,N_9716,N_7856);
or UO_476 (O_476,N_7901,N_6042);
and UO_477 (O_477,N_6190,N_7380);
or UO_478 (O_478,N_7188,N_9534);
nor UO_479 (O_479,N_7840,N_6894);
or UO_480 (O_480,N_7834,N_5385);
xnor UO_481 (O_481,N_7884,N_9495);
and UO_482 (O_482,N_7950,N_5972);
nor UO_483 (O_483,N_7182,N_6096);
xor UO_484 (O_484,N_7585,N_8241);
or UO_485 (O_485,N_8148,N_7433);
nor UO_486 (O_486,N_7311,N_5665);
nor UO_487 (O_487,N_8271,N_9684);
xor UO_488 (O_488,N_8694,N_9876);
nand UO_489 (O_489,N_7070,N_9209);
nand UO_490 (O_490,N_8988,N_9425);
xnor UO_491 (O_491,N_5273,N_8603);
or UO_492 (O_492,N_8086,N_5414);
and UO_493 (O_493,N_9564,N_7010);
nor UO_494 (O_494,N_5051,N_7837);
and UO_495 (O_495,N_5040,N_8628);
or UO_496 (O_496,N_7312,N_9279);
nand UO_497 (O_497,N_9509,N_6505);
nand UO_498 (O_498,N_8229,N_8159);
nor UO_499 (O_499,N_6750,N_5572);
nand UO_500 (O_500,N_9670,N_9126);
and UO_501 (O_501,N_9438,N_9118);
nand UO_502 (O_502,N_5319,N_5335);
or UO_503 (O_503,N_7171,N_7011);
nor UO_504 (O_504,N_7744,N_8018);
and UO_505 (O_505,N_9010,N_6267);
nor UO_506 (O_506,N_6462,N_5266);
xnor UO_507 (O_507,N_6099,N_8330);
nand UO_508 (O_508,N_8071,N_5832);
and UO_509 (O_509,N_7032,N_7175);
and UO_510 (O_510,N_7921,N_5812);
and UO_511 (O_511,N_7786,N_7158);
or UO_512 (O_512,N_6246,N_5230);
and UO_513 (O_513,N_9232,N_6604);
or UO_514 (O_514,N_6185,N_8875);
nand UO_515 (O_515,N_7280,N_5944);
and UO_516 (O_516,N_9899,N_6315);
and UO_517 (O_517,N_9178,N_9145);
xor UO_518 (O_518,N_8023,N_9033);
or UO_519 (O_519,N_9928,N_7944);
or UO_520 (O_520,N_5068,N_6905);
nand UO_521 (O_521,N_6915,N_8995);
nor UO_522 (O_522,N_5461,N_8974);
and UO_523 (O_523,N_8395,N_5737);
or UO_524 (O_524,N_6066,N_5323);
nor UO_525 (O_525,N_6560,N_9979);
nor UO_526 (O_526,N_7778,N_6919);
and UO_527 (O_527,N_7933,N_6698);
nand UO_528 (O_528,N_5048,N_7399);
and UO_529 (O_529,N_9560,N_5750);
xnor UO_530 (O_530,N_9486,N_9576);
or UO_531 (O_531,N_6667,N_5846);
and UO_532 (O_532,N_7117,N_9311);
nand UO_533 (O_533,N_9305,N_6147);
or UO_534 (O_534,N_7811,N_7753);
nand UO_535 (O_535,N_5674,N_5887);
and UO_536 (O_536,N_8517,N_5303);
nor UO_537 (O_537,N_7674,N_6520);
or UO_538 (O_538,N_9641,N_7872);
nor UO_539 (O_539,N_7099,N_9938);
or UO_540 (O_540,N_5886,N_8227);
and UO_541 (O_541,N_7159,N_6989);
or UO_542 (O_542,N_5947,N_8933);
xnor UO_543 (O_543,N_9440,N_5628);
nand UO_544 (O_544,N_9822,N_5915);
nand UO_545 (O_545,N_7393,N_6873);
nor UO_546 (O_546,N_7996,N_9694);
nor UO_547 (O_547,N_9297,N_7370);
or UO_548 (O_548,N_9039,N_6221);
or UO_549 (O_549,N_7426,N_9445);
or UO_550 (O_550,N_7977,N_8403);
nand UO_551 (O_551,N_9112,N_7034);
or UO_552 (O_552,N_7485,N_6702);
xnor UO_553 (O_553,N_8032,N_9331);
nor UO_554 (O_554,N_7680,N_8064);
and UO_555 (O_555,N_9918,N_8958);
nor UO_556 (O_556,N_5066,N_5366);
xor UO_557 (O_557,N_6668,N_5851);
xnor UO_558 (O_558,N_8791,N_9788);
xnor UO_559 (O_559,N_8903,N_8588);
or UO_560 (O_560,N_7870,N_9775);
nand UO_561 (O_561,N_5093,N_9687);
nor UO_562 (O_562,N_5027,N_9719);
or UO_563 (O_563,N_8033,N_7492);
or UO_564 (O_564,N_8778,N_7836);
nor UO_565 (O_565,N_8014,N_7782);
nand UO_566 (O_566,N_9646,N_9254);
and UO_567 (O_567,N_9630,N_8598);
or UO_568 (O_568,N_9699,N_6036);
or UO_569 (O_569,N_8575,N_8779);
and UO_570 (O_570,N_9321,N_9200);
nand UO_571 (O_571,N_5031,N_6388);
and UO_572 (O_572,N_5775,N_5413);
nand UO_573 (O_573,N_8820,N_6728);
nor UO_574 (O_574,N_8499,N_5327);
nand UO_575 (O_575,N_7970,N_8616);
or UO_576 (O_576,N_6414,N_7126);
nor UO_577 (O_577,N_7204,N_8649);
and UO_578 (O_578,N_5864,N_8168);
xnor UO_579 (O_579,N_8332,N_9706);
nand UO_580 (O_580,N_9975,N_9940);
xor UO_581 (O_581,N_7208,N_7087);
xor UO_582 (O_582,N_7606,N_6600);
xnor UO_583 (O_583,N_5880,N_6883);
nand UO_584 (O_584,N_5799,N_9583);
xnor UO_585 (O_585,N_6438,N_5192);
and UO_586 (O_586,N_8208,N_6892);
nor UO_587 (O_587,N_8345,N_8937);
nand UO_588 (O_588,N_8700,N_6851);
or UO_589 (O_589,N_8414,N_6425);
or UO_590 (O_590,N_5625,N_7430);
nor UO_591 (O_591,N_8826,N_5441);
and UO_592 (O_592,N_5748,N_6177);
and UO_593 (O_593,N_6575,N_6559);
or UO_594 (O_594,N_8920,N_9170);
and UO_595 (O_595,N_6211,N_9422);
and UO_596 (O_596,N_7636,N_6281);
nor UO_597 (O_597,N_8830,N_9651);
nor UO_598 (O_598,N_7236,N_6155);
nor UO_599 (O_599,N_9817,N_5428);
nor UO_600 (O_600,N_9739,N_5752);
and UO_601 (O_601,N_8590,N_9358);
and UO_602 (O_602,N_8851,N_8294);
nand UO_603 (O_603,N_5096,N_6463);
or UO_604 (O_604,N_9997,N_6312);
and UO_605 (O_605,N_6716,N_6270);
nor UO_606 (O_606,N_7679,N_5528);
and UO_607 (O_607,N_9703,N_8706);
or UO_608 (O_608,N_9840,N_8315);
nand UO_609 (O_609,N_8813,N_8621);
and UO_610 (O_610,N_8462,N_8334);
nor UO_611 (O_611,N_8910,N_5018);
nand UO_612 (O_612,N_8015,N_6519);
nor UO_613 (O_613,N_9664,N_7547);
or UO_614 (O_614,N_7645,N_7999);
nand UO_615 (O_615,N_5134,N_6745);
nand UO_616 (O_616,N_9101,N_7359);
nor UO_617 (O_617,N_8912,N_7590);
and UO_618 (O_618,N_7584,N_6022);
or UO_619 (O_619,N_9828,N_7637);
nor UO_620 (O_620,N_8832,N_8402);
nand UO_621 (O_621,N_5181,N_8473);
nor UO_622 (O_622,N_6727,N_6175);
nor UO_623 (O_623,N_9351,N_6117);
or UO_624 (O_624,N_7001,N_7709);
or UO_625 (O_625,N_5227,N_9686);
or UO_626 (O_626,N_6040,N_7258);
xnor UO_627 (O_627,N_5577,N_9163);
xor UO_628 (O_628,N_5117,N_5076);
and UO_629 (O_629,N_5130,N_7855);
xor UO_630 (O_630,N_7511,N_6105);
nand UO_631 (O_631,N_7134,N_5671);
or UO_632 (O_632,N_6367,N_7707);
and UO_633 (O_633,N_7181,N_6567);
nand UO_634 (O_634,N_6328,N_7233);
or UO_635 (O_635,N_9308,N_7572);
or UO_636 (O_636,N_5033,N_7119);
nor UO_637 (O_637,N_7890,N_6956);
or UO_638 (O_638,N_6538,N_7211);
and UO_639 (O_639,N_8550,N_9474);
and UO_640 (O_640,N_7819,N_5447);
nor UO_641 (O_641,N_5114,N_5718);
and UO_642 (O_642,N_7521,N_7854);
and UO_643 (O_643,N_7170,N_6674);
and UO_644 (O_644,N_6985,N_7395);
xor UO_645 (O_645,N_6060,N_6854);
and UO_646 (O_646,N_9801,N_9218);
nor UO_647 (O_647,N_8760,N_9671);
and UO_648 (O_648,N_9386,N_9513);
and UO_649 (O_649,N_7187,N_6797);
or UO_650 (O_650,N_6867,N_8372);
or UO_651 (O_651,N_5553,N_5060);
xor UO_652 (O_652,N_6928,N_5265);
or UO_653 (O_653,N_6775,N_5653);
nand UO_654 (O_654,N_6885,N_6296);
and UO_655 (O_655,N_6768,N_8743);
xnor UO_656 (O_656,N_7483,N_7165);
and UO_657 (O_657,N_8837,N_9142);
nor UO_658 (O_658,N_8311,N_9984);
nand UO_659 (O_659,N_8609,N_7653);
nor UO_660 (O_660,N_7443,N_7231);
nor UO_661 (O_661,N_9804,N_7378);
or UO_662 (O_662,N_8897,N_6703);
nor UO_663 (O_663,N_5757,N_8112);
nand UO_664 (O_664,N_7215,N_7062);
nand UO_665 (O_665,N_6273,N_7458);
and UO_666 (O_666,N_6056,N_6311);
and UO_667 (O_667,N_8660,N_7218);
nand UO_668 (O_668,N_5016,N_6030);
or UO_669 (O_669,N_9734,N_7980);
nand UO_670 (O_670,N_8435,N_5178);
or UO_671 (O_671,N_8304,N_9764);
and UO_672 (O_672,N_9974,N_5722);
nand UO_673 (O_673,N_8107,N_7135);
nor UO_674 (O_674,N_9276,N_5491);
and UO_675 (O_675,N_8276,N_5629);
nand UO_676 (O_676,N_9858,N_9075);
or UO_677 (O_677,N_6594,N_9164);
xnor UO_678 (O_678,N_5633,N_6200);
xor UO_679 (O_679,N_5361,N_6664);
nor UO_680 (O_680,N_5742,N_6490);
nand UO_681 (O_681,N_8265,N_8165);
nor UO_682 (O_682,N_6738,N_8549);
and UO_683 (O_683,N_7843,N_6882);
or UO_684 (O_684,N_9312,N_9500);
xor UO_685 (O_685,N_9337,N_9230);
nand UO_686 (O_686,N_9410,N_6261);
nor UO_687 (O_687,N_8965,N_6168);
or UO_688 (O_688,N_8853,N_5077);
xor UO_689 (O_689,N_6173,N_6521);
xor UO_690 (O_690,N_9709,N_5946);
nand UO_691 (O_691,N_6330,N_9904);
nand UO_692 (O_692,N_7445,N_5970);
xor UO_693 (O_693,N_7581,N_8377);
nor UO_694 (O_694,N_5508,N_6432);
nor UO_695 (O_695,N_7749,N_6283);
nor UO_696 (O_696,N_5875,N_9913);
nor UO_697 (O_697,N_7120,N_5021);
xor UO_698 (O_698,N_7686,N_6708);
or UO_699 (O_699,N_8980,N_6868);
or UO_700 (O_700,N_7738,N_7044);
or UO_701 (O_701,N_7643,N_7787);
and UO_702 (O_702,N_9081,N_7595);
xnor UO_703 (O_703,N_5210,N_9054);
and UO_704 (O_704,N_7551,N_8257);
nor UO_705 (O_705,N_6996,N_5350);
and UO_706 (O_706,N_7263,N_6376);
nor UO_707 (O_707,N_7301,N_7628);
and UO_708 (O_708,N_9100,N_6720);
or UO_709 (O_709,N_6039,N_9774);
nand UO_710 (O_710,N_6198,N_5260);
or UO_711 (O_711,N_6595,N_6236);
and UO_712 (O_712,N_8061,N_5121);
nor UO_713 (O_713,N_6219,N_5739);
xor UO_714 (O_714,N_9749,N_7832);
nand UO_715 (O_715,N_7802,N_8825);
and UO_716 (O_716,N_9785,N_7364);
nand UO_717 (O_717,N_9553,N_8893);
or UO_718 (O_718,N_6306,N_7206);
nand UO_719 (O_719,N_5704,N_6174);
or UO_720 (O_720,N_5586,N_7642);
or UO_721 (O_721,N_7394,N_9227);
nor UO_722 (O_722,N_6231,N_5836);
nor UO_723 (O_723,N_8401,N_8418);
nor UO_724 (O_724,N_9760,N_9780);
or UO_725 (O_725,N_9605,N_8249);
and UO_726 (O_726,N_8684,N_5343);
nor UO_727 (O_727,N_8342,N_6570);
and UO_728 (O_728,N_7143,N_6944);
nor UO_729 (O_729,N_7510,N_7431);
nand UO_730 (O_730,N_5047,N_7262);
or UO_731 (O_731,N_9202,N_7615);
or UO_732 (O_732,N_7880,N_7948);
nor UO_733 (O_733,N_5120,N_9371);
nor UO_734 (O_734,N_6230,N_6859);
and UO_735 (O_735,N_6103,N_9968);
nor UO_736 (O_736,N_8481,N_8524);
and UO_737 (O_737,N_9080,N_9705);
and UO_738 (O_738,N_7730,N_8358);
xnor UO_739 (O_739,N_6661,N_5529);
xnor UO_740 (O_740,N_6697,N_7057);
nand UO_741 (O_741,N_6729,N_7092);
nor UO_742 (O_742,N_6166,N_8114);
nand UO_743 (O_743,N_9867,N_6627);
or UO_744 (O_744,N_9147,N_7331);
nor UO_745 (O_745,N_9018,N_5314);
or UO_746 (O_746,N_9518,N_7984);
nor UO_747 (O_747,N_9873,N_5450);
xor UO_748 (O_748,N_9847,N_8307);
or UO_749 (O_749,N_9330,N_9055);
or UO_750 (O_750,N_7555,N_9581);
and UO_751 (O_751,N_7683,N_7719);
nand UO_752 (O_752,N_5211,N_9394);
and UO_753 (O_753,N_8072,N_5942);
and UO_754 (O_754,N_5856,N_5511);
or UO_755 (O_755,N_6706,N_7731);
and UO_756 (O_756,N_9797,N_5660);
or UO_757 (O_757,N_8690,N_7987);
xnor UO_758 (O_758,N_5326,N_7906);
xor UO_759 (O_759,N_8119,N_5907);
and UO_760 (O_760,N_8421,N_7997);
and UO_761 (O_761,N_7012,N_7597);
nor UO_762 (O_762,N_6912,N_6526);
or UO_763 (O_763,N_8707,N_8142);
nand UO_764 (O_764,N_7232,N_5558);
nand UO_765 (O_765,N_8508,N_7212);
and UO_766 (O_766,N_9757,N_5474);
nand UO_767 (O_767,N_6734,N_7850);
or UO_768 (O_768,N_9464,N_5443);
and UO_769 (O_769,N_5717,N_6902);
nand UO_770 (O_770,N_5957,N_6971);
nor UO_771 (O_771,N_6806,N_9115);
nand UO_772 (O_772,N_9363,N_5694);
nand UO_773 (O_773,N_7540,N_6693);
nor UO_774 (O_774,N_8124,N_7857);
and UO_775 (O_775,N_6305,N_9038);
xor UO_776 (O_776,N_8357,N_9692);
and UO_777 (O_777,N_9399,N_9155);
xor UO_778 (O_778,N_6565,N_5515);
nor UO_779 (O_779,N_7205,N_8313);
nand UO_780 (O_780,N_9932,N_8288);
nand UO_781 (O_781,N_9778,N_6003);
or UO_782 (O_782,N_5902,N_9213);
or UO_783 (O_783,N_6976,N_5107);
and UO_784 (O_784,N_8297,N_9427);
nand UO_785 (O_785,N_7641,N_9502);
or UO_786 (O_786,N_9570,N_7605);
nor UO_787 (O_787,N_5179,N_7612);
xor UO_788 (O_788,N_9053,N_5332);
and UO_789 (O_789,N_9713,N_6648);
nand UO_790 (O_790,N_8854,N_5672);
or UO_791 (O_791,N_6427,N_5281);
nor UO_792 (O_792,N_8763,N_8464);
and UO_793 (O_793,N_9106,N_6428);
and UO_794 (O_794,N_9067,N_9726);
nor UO_795 (O_795,N_6180,N_8138);
or UO_796 (O_796,N_5404,N_5609);
nand UO_797 (O_797,N_9985,N_5774);
nand UO_798 (O_798,N_5600,N_5259);
nor UO_799 (O_799,N_9162,N_8482);
nand UO_800 (O_800,N_9029,N_6413);
or UO_801 (O_801,N_6314,N_6389);
xor UO_802 (O_802,N_8720,N_9599);
and UO_803 (O_803,N_6961,N_7777);
nand UO_804 (O_804,N_7544,N_5865);
nor UO_805 (O_805,N_8205,N_8200);
nand UO_806 (O_806,N_6000,N_9654);
and UO_807 (O_807,N_5399,N_8679);
or UO_808 (O_808,N_5487,N_6949);
and UO_809 (O_809,N_5351,N_9827);
or UO_810 (O_810,N_7934,N_9620);
or UO_811 (O_811,N_6763,N_8724);
and UO_812 (O_812,N_6825,N_7766);
and UO_813 (O_813,N_8765,N_8541);
nand UO_814 (O_814,N_7264,N_8539);
and UO_815 (O_815,N_9392,N_7514);
and UO_816 (O_816,N_7711,N_8424);
or UO_817 (O_817,N_7925,N_9890);
and UO_818 (O_818,N_7347,N_6824);
or UO_819 (O_819,N_8533,N_9786);
nor UO_820 (O_820,N_7242,N_9854);
xor UO_821 (O_821,N_5821,N_8324);
xnor UO_822 (O_822,N_8945,N_7321);
or UO_823 (O_823,N_8316,N_8420);
or UO_824 (O_824,N_5396,N_5644);
nand UO_825 (O_825,N_7105,N_9193);
nor UO_826 (O_826,N_9415,N_5338);
nor UO_827 (O_827,N_8511,N_5213);
or UO_828 (O_828,N_5012,N_7438);
nor UO_829 (O_829,N_9467,N_6580);
and UO_830 (O_830,N_9028,N_8173);
or UO_831 (O_831,N_6068,N_9919);
or UO_832 (O_832,N_9856,N_8622);
nor UO_833 (O_833,N_5579,N_8019);
and UO_834 (O_834,N_7269,N_7362);
xor UO_835 (O_835,N_6686,N_6953);
nand UO_836 (O_836,N_7894,N_8167);
and UO_837 (O_837,N_7792,N_5057);
xor UO_838 (O_838,N_6517,N_5253);
nand UO_839 (O_839,N_8037,N_5869);
nor UO_840 (O_840,N_6951,N_8493);
xnor UO_841 (O_841,N_5251,N_6035);
and UO_842 (O_842,N_9257,N_6631);
nor UO_843 (O_843,N_9821,N_5967);
nor UO_844 (O_844,N_5828,N_9885);
xor UO_845 (O_845,N_5545,N_8573);
and UO_846 (O_846,N_8672,N_6308);
or UO_847 (O_847,N_7052,N_9222);
and UO_848 (O_848,N_9283,N_8683);
nand UO_849 (O_849,N_5983,N_9818);
and UO_850 (O_850,N_6981,N_6537);
nand UO_851 (O_851,N_6437,N_5187);
or UO_852 (O_852,N_9195,N_9711);
xor UO_853 (O_853,N_6512,N_6149);
or UO_854 (O_854,N_7411,N_9954);
nand UO_855 (O_855,N_9948,N_8407);
and UO_856 (O_856,N_8184,N_5296);
nor UO_857 (O_857,N_9285,N_6506);
and UO_858 (O_858,N_8410,N_5405);
or UO_859 (O_859,N_5365,N_6857);
nand UO_860 (O_860,N_6907,N_7216);
nand UO_861 (O_861,N_7705,N_6384);
or UO_862 (O_862,N_8394,N_8329);
and UO_863 (O_863,N_8669,N_8618);
or UO_864 (O_864,N_8381,N_5668);
and UO_865 (O_865,N_7756,N_9241);
and UO_866 (O_866,N_9260,N_5686);
nand UO_867 (O_867,N_8983,N_5854);
nor UO_868 (O_868,N_6406,N_8710);
and UO_869 (O_869,N_6772,N_5457);
or UO_870 (O_870,N_8035,N_6864);
and UO_871 (O_871,N_8557,N_6685);
or UO_872 (O_872,N_8891,N_8163);
and UO_873 (O_873,N_5982,N_8586);
nor UO_874 (O_874,N_7903,N_8454);
nor UO_875 (O_875,N_5993,N_7814);
and UO_876 (O_876,N_8178,N_6148);
xnor UO_877 (O_877,N_9240,N_7118);
and UO_878 (O_878,N_5431,N_5892);
nand UO_879 (O_879,N_6071,N_5334);
nor UO_880 (O_880,N_8693,N_7538);
nand UO_881 (O_881,N_8088,N_7929);
and UO_882 (O_882,N_6548,N_9957);
and UO_883 (O_883,N_6160,N_9182);
or UO_884 (O_884,N_7732,N_8739);
or UO_885 (O_885,N_5649,N_7220);
nor UO_886 (O_886,N_7530,N_7360);
or UO_887 (O_887,N_5912,N_5244);
xor UO_888 (O_888,N_7509,N_7457);
nand UO_889 (O_889,N_6946,N_9268);
or UO_890 (O_890,N_9922,N_9925);
nor UO_891 (O_891,N_6922,N_5348);
xnor UO_892 (O_892,N_8209,N_5406);
or UO_893 (O_893,N_8568,N_8453);
and UO_894 (O_894,N_7865,N_8561);
and UO_895 (O_895,N_9139,N_5226);
or UO_896 (O_896,N_6020,N_8281);
nand UO_897 (O_897,N_8793,N_9636);
and UO_898 (O_898,N_7174,N_6625);
or UO_899 (O_899,N_6008,N_9426);
nor UO_900 (O_900,N_6167,N_6278);
nor UO_901 (O_901,N_9939,N_9306);
and UO_902 (O_902,N_9747,N_7223);
and UO_903 (O_903,N_9402,N_5356);
and UO_904 (O_904,N_8267,N_9180);
and UO_905 (O_905,N_6045,N_9083);
and UO_906 (O_906,N_8828,N_9505);
xor UO_907 (O_907,N_5688,N_7784);
and UO_908 (O_908,N_6422,N_9102);
and UO_909 (O_909,N_5507,N_7989);
nor UO_910 (O_910,N_7729,N_9443);
and UO_911 (O_911,N_5998,N_8082);
or UO_912 (O_912,N_5652,N_9483);
or UO_913 (O_913,N_9650,N_7293);
nor UO_914 (O_914,N_8451,N_6690);
or UO_915 (O_915,N_7852,N_6088);
or UO_916 (O_916,N_5030,N_7807);
nor UO_917 (O_917,N_6016,N_7633);
and UO_918 (O_918,N_8979,N_5787);
nand UO_919 (O_919,N_7481,N_5223);
nor UO_920 (O_920,N_8101,N_5905);
xor UO_921 (O_921,N_5922,N_6187);
nor UO_922 (O_922,N_6789,N_6322);
nor UO_923 (O_923,N_9116,N_8327);
nand UO_924 (O_924,N_6248,N_7199);
or UO_925 (O_925,N_6164,N_8067);
and UO_926 (O_926,N_5622,N_5278);
and UO_927 (O_927,N_9369,N_8909);
nand UO_928 (O_928,N_5218,N_7568);
or UO_929 (O_929,N_6176,N_6345);
and UO_930 (O_930,N_6062,N_9717);
or UO_931 (O_931,N_7414,N_8976);
and UO_932 (O_932,N_5986,N_9339);
or UO_933 (O_933,N_6722,N_8425);
or UO_934 (O_934,N_9284,N_8545);
xnor UO_935 (O_935,N_8636,N_8488);
nor UO_936 (O_936,N_5608,N_8049);
nor UO_937 (O_937,N_5375,N_9150);
nor UO_938 (O_938,N_8602,N_6969);
or UO_939 (O_939,N_9017,N_7864);
nand UO_940 (O_940,N_6798,N_6760);
xor UO_941 (O_941,N_5147,N_8723);
nor UO_942 (O_942,N_5346,N_7693);
nor UO_943 (O_943,N_7413,N_9991);
nor UO_944 (O_944,N_7639,N_6898);
or UO_945 (O_945,N_6966,N_7938);
or UO_946 (O_946,N_5853,N_5939);
nor UO_947 (O_947,N_6429,N_7759);
and UO_948 (O_948,N_7382,N_7229);
and UO_949 (O_949,N_6461,N_6802);
nor UO_950 (O_950,N_9565,N_7487);
nor UO_951 (O_951,N_6795,N_5198);
or UO_952 (O_952,N_9627,N_9701);
nand UO_953 (O_953,N_8351,N_8600);
nand UO_954 (O_954,N_6665,N_9990);
nor UO_955 (O_955,N_9524,N_9970);
and UO_956 (O_956,N_8807,N_5820);
or UO_957 (O_957,N_6659,N_7853);
and UO_958 (O_958,N_7084,N_8896);
nand UO_959 (O_959,N_7017,N_9156);
xor UO_960 (O_960,N_8359,N_9465);
nor UO_961 (O_961,N_8443,N_9642);
nor UO_962 (O_962,N_5906,N_8286);
or UO_963 (O_963,N_9643,N_9435);
nand UO_964 (O_964,N_6141,N_7163);
or UO_965 (O_965,N_6138,N_8022);
nand UO_966 (O_966,N_6309,N_9403);
or UO_967 (O_967,N_6532,N_7184);
and UO_968 (O_968,N_6983,N_5713);
nand UO_969 (O_969,N_5143,N_6280);
nor UO_970 (O_970,N_6645,N_6653);
or UO_971 (O_971,N_5391,N_5146);
and UO_972 (O_972,N_7804,N_6704);
or UO_973 (O_973,N_8615,N_6341);
and UO_974 (O_974,N_7764,N_7488);
or UO_975 (O_975,N_6011,N_5297);
and UO_976 (O_976,N_9832,N_5378);
nand UO_977 (O_977,N_5611,N_9324);
nor UO_978 (O_978,N_6226,N_5612);
and UO_979 (O_979,N_6179,N_7806);
or UO_980 (O_980,N_7282,N_8695);
and UO_981 (O_981,N_5156,N_7965);
or UO_982 (O_982,N_7567,N_5565);
or UO_983 (O_983,N_7726,N_5909);
or UO_984 (O_984,N_7952,N_8469);
or UO_985 (O_985,N_7839,N_8744);
xnor UO_986 (O_986,N_5747,N_8899);
and UO_987 (O_987,N_9007,N_7245);
nand UO_988 (O_988,N_7918,N_7594);
nand UO_989 (O_989,N_8972,N_8951);
and UO_990 (O_990,N_8692,N_6234);
nand UO_991 (O_991,N_8433,N_9484);
nor UO_992 (O_992,N_8675,N_6049);
nor UO_993 (O_993,N_9662,N_8783);
xor UO_994 (O_994,N_8232,N_9585);
nor UO_995 (O_995,N_9988,N_7937);
xor UO_996 (O_996,N_8943,N_8806);
or UO_997 (O_997,N_5539,N_6958);
and UO_998 (O_998,N_7772,N_7335);
nor UO_999 (O_999,N_9888,N_6370);
or UO_1000 (O_1000,N_8644,N_7527);
nor UO_1001 (O_1001,N_7365,N_7640);
nor UO_1002 (O_1002,N_5696,N_9011);
nor UO_1003 (O_1003,N_7314,N_7868);
nand UO_1004 (O_1004,N_6817,N_8564);
nor UO_1005 (O_1005,N_7793,N_9667);
and UO_1006 (O_1006,N_9714,N_9076);
nor UO_1007 (O_1007,N_6725,N_5548);
xor UO_1008 (O_1008,N_9781,N_7467);
nand UO_1009 (O_1009,N_6914,N_6984);
nand UO_1010 (O_1010,N_8190,N_8062);
xor UO_1011 (O_1011,N_7664,N_9250);
and UO_1012 (O_1012,N_8323,N_6694);
nor UO_1013 (O_1013,N_6998,N_9400);
or UO_1014 (O_1014,N_8840,N_9176);
nor UO_1015 (O_1015,N_6581,N_9493);
xnor UO_1016 (O_1016,N_9190,N_5975);
xnor UO_1017 (O_1017,N_9907,N_9996);
nand UO_1018 (O_1018,N_5038,N_8719);
and UO_1019 (O_1019,N_9515,N_7978);
xor UO_1020 (O_1020,N_8459,N_7286);
and UO_1021 (O_1021,N_8585,N_9251);
or UO_1022 (O_1022,N_5833,N_8186);
or UO_1023 (O_1023,N_8497,N_6622);
nand UO_1024 (O_1024,N_8343,N_8474);
nand UO_1025 (O_1025,N_6637,N_8643);
xor UO_1026 (O_1026,N_7962,N_8116);
and UO_1027 (O_1027,N_7964,N_8577);
or UO_1028 (O_1028,N_7945,N_9697);
or UO_1029 (O_1029,N_6972,N_5973);
nand UO_1030 (O_1030,N_9964,N_8468);
nor UO_1031 (O_1031,N_7554,N_8831);
nor UO_1032 (O_1032,N_6090,N_7508);
nand UO_1033 (O_1033,N_5310,N_6592);
xnor UO_1034 (O_1034,N_7177,N_9390);
and UO_1035 (O_1035,N_8231,N_7667);
and UO_1036 (O_1036,N_5530,N_6418);
and UO_1037 (O_1037,N_9580,N_5991);
and UO_1038 (O_1038,N_7131,N_9676);
nand UO_1039 (O_1039,N_6339,N_5848);
nand UO_1040 (O_1040,N_6880,N_9077);
nor UO_1041 (O_1041,N_9446,N_5751);
nand UO_1042 (O_1042,N_8065,N_8882);
and UO_1043 (O_1043,N_5324,N_9211);
nand UO_1044 (O_1044,N_7986,N_5587);
and UO_1045 (O_1045,N_9329,N_9237);
nor UO_1046 (O_1046,N_9491,N_9345);
or UO_1047 (O_1047,N_7882,N_9724);
xor UO_1048 (O_1048,N_6782,N_6787);
xor UO_1049 (O_1049,N_8824,N_5913);
and UO_1050 (O_1050,N_8079,N_7441);
nand UO_1051 (O_1051,N_5870,N_7586);
and UO_1052 (O_1052,N_8529,N_6044);
and UO_1053 (O_1053,N_7881,N_7690);
or UO_1054 (O_1054,N_5400,N_7758);
nor UO_1055 (O_1055,N_8911,N_5495);
and UO_1056 (O_1056,N_9277,N_5896);
nor UO_1057 (O_1057,N_9956,N_9533);
nand UO_1058 (O_1058,N_6057,N_5122);
nor UO_1059 (O_1059,N_9258,N_7246);
nand UO_1060 (O_1060,N_7698,N_8136);
or UO_1061 (O_1061,N_7063,N_9481);
and UO_1062 (O_1062,N_6372,N_9043);
nand UO_1063 (O_1063,N_8570,N_8172);
nand UO_1064 (O_1064,N_6292,N_6434);
and UO_1065 (O_1065,N_9871,N_9594);
nor UO_1066 (O_1066,N_8199,N_7408);
nand UO_1067 (O_1067,N_7435,N_9489);
or UO_1068 (O_1068,N_5890,N_8339);
nor UO_1069 (O_1069,N_7943,N_9503);
nor UO_1070 (O_1070,N_6583,N_7296);
nor UO_1071 (O_1071,N_6809,N_5043);
nor UO_1072 (O_1072,N_5354,N_5081);
and UO_1073 (O_1073,N_7019,N_9631);
and UO_1074 (O_1074,N_8772,N_9002);
nor UO_1075 (O_1075,N_7456,N_8687);
or UO_1076 (O_1076,N_7023,N_8582);
or UO_1077 (O_1077,N_5243,N_7650);
or UO_1078 (O_1078,N_6899,N_8780);
xor UO_1079 (O_1079,N_8986,N_5813);
and UO_1080 (O_1080,N_6076,N_8466);
and UO_1081 (O_1081,N_5209,N_8918);
nor UO_1082 (O_1082,N_5601,N_8691);
nand UO_1083 (O_1083,N_7356,N_8614);
and UO_1084 (O_1084,N_7704,N_5502);
nand UO_1085 (O_1085,N_8194,N_7951);
nand UO_1086 (O_1086,N_5605,N_6054);
and UO_1087 (O_1087,N_9619,N_9792);
nor UO_1088 (O_1088,N_6394,N_6197);
or UO_1089 (O_1089,N_5949,N_5825);
nor UO_1090 (O_1090,N_6962,N_8181);
and UO_1091 (O_1091,N_7678,N_9507);
nor UO_1092 (O_1092,N_7604,N_7842);
nor UO_1093 (O_1093,N_6075,N_8317);
nand UO_1094 (O_1094,N_8888,N_9659);
or UO_1095 (O_1095,N_5379,N_8814);
xnor UO_1096 (O_1096,N_8333,N_6402);
nor UO_1097 (O_1097,N_9019,N_7197);
or UO_1098 (O_1098,N_5464,N_9870);
and UO_1099 (O_1099,N_5834,N_5173);
or UO_1100 (O_1100,N_8775,N_5921);
nor UO_1101 (O_1101,N_9720,N_8559);
or UO_1102 (O_1102,N_5822,N_9383);
xor UO_1103 (O_1103,N_7993,N_6493);
or UO_1104 (O_1104,N_5446,N_8534);
or UO_1105 (O_1105,N_6395,N_7470);
or UO_1106 (O_1106,N_9255,N_9395);
nor UO_1107 (O_1107,N_5025,N_7288);
and UO_1108 (O_1108,N_9498,N_8766);
nand UO_1109 (O_1109,N_5056,N_6531);
nand UO_1110 (O_1110,N_8318,N_5054);
or UO_1111 (O_1111,N_6832,N_8326);
or UO_1112 (O_1112,N_8864,N_6095);
nand UO_1113 (O_1113,N_5546,N_5994);
nor UO_1114 (O_1114,N_6543,N_8439);
nor UO_1115 (O_1115,N_7169,N_5841);
nand UO_1116 (O_1116,N_7888,N_9287);
and UO_1117 (O_1117,N_9199,N_5427);
and UO_1118 (O_1118,N_7960,N_8610);
nand UO_1119 (O_1119,N_9423,N_6373);
xnor UO_1120 (O_1120,N_7501,N_8118);
and UO_1121 (O_1121,N_9567,N_7543);
or UO_1122 (O_1122,N_5918,N_7313);
or UO_1123 (O_1123,N_9499,N_8467);
or UO_1124 (O_1124,N_8127,N_6591);
and UO_1125 (O_1125,N_8992,N_8132);
nor UO_1126 (O_1126,N_8985,N_7845);
nand UO_1127 (O_1127,N_5641,N_7196);
nand UO_1128 (O_1128,N_7104,N_9447);
xnor UO_1129 (O_1129,N_8855,N_8594);
and UO_1130 (O_1130,N_8535,N_8393);
or UO_1131 (O_1131,N_8126,N_6029);
and UO_1132 (O_1132,N_8161,N_7907);
or UO_1133 (O_1133,N_5990,N_7582);
nand UO_1134 (O_1134,N_8038,N_8997);
nand UO_1135 (O_1135,N_6256,N_9223);
and UO_1136 (O_1136,N_6420,N_8321);
nor UO_1137 (O_1137,N_7577,N_6225);
or UO_1138 (O_1138,N_9702,N_9228);
nand UO_1139 (O_1139,N_9138,N_5627);
nor UO_1140 (O_1140,N_7151,N_9571);
and UO_1141 (O_1141,N_9272,N_8753);
nor UO_1142 (O_1142,N_7257,N_5685);
or UO_1143 (O_1143,N_8411,N_6412);
and UO_1144 (O_1144,N_6063,N_6443);
or UO_1145 (O_1145,N_7155,N_6487);
nand UO_1146 (O_1146,N_7373,N_7127);
xnor UO_1147 (O_1147,N_6124,N_6254);
or UO_1148 (O_1148,N_6753,N_7771);
or UO_1149 (O_1149,N_9768,N_8353);
nor UO_1150 (O_1150,N_9062,N_9680);
nand UO_1151 (O_1151,N_7324,N_8842);
and UO_1152 (O_1152,N_7377,N_8716);
nand UO_1153 (O_1153,N_8302,N_5966);
and UO_1154 (O_1154,N_7776,N_6072);
nor UO_1155 (O_1155,N_8396,N_6410);
or UO_1156 (O_1156,N_8108,N_6858);
xor UO_1157 (O_1157,N_7108,N_7367);
xor UO_1158 (O_1158,N_5557,N_7990);
nor UO_1159 (O_1159,N_5015,N_6251);
nor UO_1160 (O_1160,N_9830,N_9683);
or UO_1161 (O_1161,N_8762,N_5440);
nand UO_1162 (O_1162,N_6043,N_5160);
nand UO_1163 (O_1163,N_9496,N_7869);
nand UO_1164 (O_1164,N_8975,N_6676);
nand UO_1165 (O_1165,N_9437,N_7800);
nand UO_1166 (O_1166,N_9393,N_8876);
and UO_1167 (O_1167,N_7253,N_9908);
or UO_1168 (O_1168,N_9514,N_5115);
and UO_1169 (O_1169,N_9207,N_7507);
or UO_1170 (O_1170,N_6620,N_9247);
nand UO_1171 (O_1171,N_5564,N_8479);
nor UO_1172 (O_1172,N_9480,N_9108);
and UO_1173 (O_1173,N_9024,N_8522);
or UO_1174 (O_1174,N_5884,N_5333);
nand UO_1175 (O_1175,N_5312,N_9588);
or UO_1176 (O_1176,N_9121,N_7973);
and UO_1177 (O_1177,N_9239,N_7783);
nand UO_1178 (O_1178,N_6263,N_9973);
or UO_1179 (O_1179,N_5384,N_7661);
nor UO_1180 (O_1180,N_5256,N_7371);
or UO_1181 (O_1181,N_8477,N_5358);
and UO_1182 (O_1182,N_9861,N_8665);
or UO_1183 (O_1183,N_6791,N_7534);
or UO_1184 (O_1184,N_9563,N_5386);
nand UO_1185 (O_1185,N_6804,N_7040);
nor UO_1186 (O_1186,N_8391,N_8287);
or UO_1187 (O_1187,N_6812,N_8458);
nor UO_1188 (O_1188,N_6358,N_5786);
and UO_1189 (O_1189,N_5662,N_6500);
or UO_1190 (O_1190,N_6457,N_8135);
or UO_1191 (O_1191,N_5664,N_6908);
nand UO_1192 (O_1192,N_8677,N_5583);
xor UO_1193 (O_1193,N_5893,N_5085);
and UO_1194 (O_1194,N_6276,N_6275);
or UO_1195 (O_1195,N_8193,N_9756);
nand UO_1196 (O_1196,N_6687,N_9273);
nand UO_1197 (O_1197,N_7939,N_5527);
nand UO_1198 (O_1198,N_6975,N_5316);
or UO_1199 (O_1199,N_7238,N_8547);
and UO_1200 (O_1200,N_8593,N_8470);
nor UO_1201 (O_1201,N_5995,N_9035);
xnor UO_1202 (O_1202,N_7474,N_5526);
or UO_1203 (O_1203,N_9738,N_9742);
or UO_1204 (O_1204,N_5597,N_8871);
nor UO_1205 (O_1205,N_5248,N_5083);
and UO_1206 (O_1206,N_9299,N_7192);
or UO_1207 (O_1207,N_8152,N_8109);
or UO_1208 (O_1208,N_7076,N_7763);
or UO_1209 (O_1209,N_8627,N_5926);
nor UO_1210 (O_1210,N_7859,N_8569);
xor UO_1211 (O_1211,N_7998,N_9266);
nand UO_1212 (O_1212,N_8623,N_6987);
and UO_1213 (O_1213,N_5861,N_6756);
and UO_1214 (O_1214,N_6737,N_8969);
nand UO_1215 (O_1215,N_5275,N_8729);
nand UO_1216 (O_1216,N_5473,N_5098);
and UO_1217 (O_1217,N_8449,N_5233);
or UO_1218 (O_1218,N_8000,N_8423);
or UO_1219 (O_1219,N_8378,N_5496);
or UO_1220 (O_1220,N_9405,N_5874);
nand UO_1221 (O_1221,N_5933,N_6796);
or UO_1222 (O_1222,N_9685,N_5004);
nand UO_1223 (O_1223,N_7067,N_8498);
xnor UO_1224 (O_1224,N_8844,N_7464);
nor UO_1225 (O_1225,N_5078,N_5818);
nand UO_1226 (O_1226,N_6344,N_7240);
and UO_1227 (O_1227,N_9365,N_7372);
nor UO_1228 (O_1228,N_5780,N_7974);
nand UO_1229 (O_1229,N_9290,N_9478);
nand UO_1230 (O_1230,N_9782,N_8895);
and UO_1231 (O_1231,N_8389,N_9309);
nor UO_1232 (O_1232,N_7728,N_9006);
nor UO_1233 (O_1233,N_7237,N_6116);
nand UO_1234 (O_1234,N_9900,N_5418);
nand UO_1235 (O_1235,N_8375,N_9069);
nand UO_1236 (O_1236,N_9591,N_6086);
or UO_1237 (O_1237,N_9352,N_8850);
and UO_1238 (O_1238,N_6233,N_7114);
nand UO_1239 (O_1239,N_8721,N_8565);
or UO_1240 (O_1240,N_9380,N_9980);
nor UO_1241 (O_1241,N_6282,N_5127);
nand UO_1242 (O_1242,N_5086,N_8246);
xor UO_1243 (O_1243,N_6409,N_5509);
or UO_1244 (O_1244,N_7820,N_6191);
or UO_1245 (O_1245,N_6498,N_5920);
nor UO_1246 (O_1246,N_8284,N_8238);
or UO_1247 (O_1247,N_7677,N_9892);
and UO_1248 (O_1248,N_5736,N_8968);
xnor UO_1249 (O_1249,N_8558,N_6268);
nand UO_1250 (O_1250,N_7343,N_6758);
nand UO_1251 (O_1251,N_9673,N_6127);
or UO_1252 (O_1252,N_6957,N_8280);
or UO_1253 (O_1253,N_8005,N_5640);
and UO_1254 (O_1254,N_8733,N_9732);
or UO_1255 (O_1255,N_6669,N_6938);
and UO_1256 (O_1256,N_9783,N_8243);
or UO_1257 (O_1257,N_7791,N_5318);
nand UO_1258 (O_1258,N_7326,N_7056);
nor UO_1259 (O_1259,N_6835,N_7895);
nor UO_1260 (O_1260,N_7517,N_7910);
nand UO_1261 (O_1261,N_5520,N_8898);
nand UO_1262 (O_1262,N_7684,N_8230);
or UO_1263 (O_1263,N_8147,N_7292);
nor UO_1264 (O_1264,N_9157,N_5651);
nand UO_1265 (O_1265,N_8810,N_6721);
and UO_1266 (O_1266,N_9016,N_7623);
and UO_1267 (O_1267,N_8589,N_8278);
nand UO_1268 (O_1268,N_6411,N_8360);
nand UO_1269 (O_1269,N_8149,N_8328);
and UO_1270 (O_1270,N_8373,N_9342);
and UO_1271 (O_1271,N_9547,N_8309);
nand UO_1272 (O_1272,N_5300,N_9014);
and UO_1273 (O_1273,N_9998,N_5603);
or UO_1274 (O_1274,N_7574,N_6287);
nor UO_1275 (O_1275,N_5698,N_5732);
and UO_1276 (O_1276,N_9989,N_5123);
and UO_1277 (O_1277,N_7081,N_7147);
nand UO_1278 (O_1278,N_7505,N_5308);
nor UO_1279 (O_1279,N_7439,N_6973);
nand UO_1280 (O_1280,N_5493,N_5955);
or UO_1281 (O_1281,N_9204,N_7817);
and UO_1282 (O_1282,N_5290,N_5460);
or UO_1283 (O_1283,N_5339,N_7983);
or UO_1284 (O_1284,N_9245,N_9946);
or UO_1285 (O_1285,N_6865,N_6460);
nor UO_1286 (O_1286,N_8746,N_6223);
nor UO_1287 (O_1287,N_5997,N_9140);
and UO_1288 (O_1288,N_8674,N_8865);
xor UO_1289 (O_1289,N_6988,N_7712);
nand UO_1290 (O_1290,N_7329,N_5765);
nand UO_1291 (O_1291,N_8370,N_9981);
or UO_1292 (O_1292,N_9281,N_9110);
nand UO_1293 (O_1293,N_8300,N_7325);
nand UO_1294 (O_1294,N_5184,N_8816);
xnor UO_1295 (O_1295,N_6936,N_6354);
nor UO_1296 (O_1296,N_7936,N_6555);
nand UO_1297 (O_1297,N_6145,N_8924);
or UO_1298 (O_1298,N_6365,N_6651);
or UO_1299 (O_1299,N_9256,N_9530);
nand UO_1300 (O_1300,N_5716,N_8338);
or UO_1301 (O_1301,N_9878,N_6255);
nor UO_1302 (O_1302,N_8051,N_7028);
nor UO_1303 (O_1303,N_9041,N_8283);
nor UO_1304 (O_1304,N_5879,N_5383);
and UO_1305 (O_1305,N_7876,N_8846);
nor UO_1306 (O_1306,N_6349,N_6298);
nor UO_1307 (O_1307,N_5347,N_6830);
or UO_1308 (O_1308,N_5172,N_6486);
and UO_1309 (O_1309,N_5793,N_7183);
xor UO_1310 (O_1310,N_8777,N_5469);
and UO_1311 (O_1311,N_5531,N_5458);
nor UO_1312 (O_1312,N_5961,N_7137);
nand UO_1313 (O_1313,N_6542,N_6374);
xnor UO_1314 (O_1314,N_8085,N_8886);
and UO_1315 (O_1315,N_9307,N_5180);
and UO_1316 (O_1316,N_8686,N_6930);
or UO_1317 (O_1317,N_7716,N_5630);
nand UO_1318 (O_1318,N_5005,N_5837);
and UO_1319 (O_1319,N_8303,N_5252);
and UO_1320 (O_1320,N_8463,N_9153);
nor UO_1321 (O_1321,N_9910,N_5724);
or UO_1322 (O_1322,N_5293,N_9013);
or UO_1323 (O_1323,N_5433,N_6869);
nand UO_1324 (O_1324,N_9298,N_7013);
or UO_1325 (O_1325,N_8296,N_5914);
nor UO_1326 (O_1326,N_6295,N_5315);
nand UO_1327 (O_1327,N_5468,N_9253);
or UO_1328 (O_1328,N_6169,N_6557);
nor UO_1329 (O_1329,N_9660,N_5028);
nor UO_1330 (O_1330,N_9874,N_6672);
nand UO_1331 (O_1331,N_8653,N_9375);
or UO_1332 (O_1332,N_5749,N_7513);
nand UO_1333 (O_1333,N_9424,N_6082);
nor UO_1334 (O_1334,N_6494,N_7748);
nor UO_1335 (O_1335,N_6662,N_6813);
or UO_1336 (O_1336,N_5613,N_5683);
or UO_1337 (O_1337,N_5569,N_8939);
nand UO_1338 (O_1338,N_8634,N_7638);
nand UO_1339 (O_1339,N_7466,N_8587);
and UO_1340 (O_1340,N_9950,N_8748);
nor UO_1341 (O_1341,N_7152,N_8164);
nor UO_1342 (O_1342,N_5726,N_5097);
xor UO_1343 (O_1343,N_5231,N_5604);
nor UO_1344 (O_1344,N_8021,N_8504);
nand UO_1345 (O_1345,N_5376,N_6770);
or UO_1346 (O_1346,N_9537,N_7575);
nand UO_1347 (O_1347,N_6779,N_9335);
nor UO_1348 (O_1348,N_7448,N_7167);
nand UO_1349 (O_1349,N_7515,N_8406);
nand UO_1350 (O_1350,N_8228,N_8385);
or UO_1351 (O_1351,N_7058,N_5779);
and UO_1352 (O_1352,N_8917,N_7476);
and UO_1353 (O_1353,N_8179,N_9586);
and UO_1354 (O_1354,N_6822,N_6467);
nand UO_1355 (O_1355,N_6333,N_5788);
nor UO_1356 (O_1356,N_7621,N_5755);
or UO_1357 (O_1357,N_7157,N_8712);
and UO_1358 (O_1358,N_5807,N_5003);
nor UO_1359 (O_1359,N_5084,N_6613);
or UO_1360 (O_1360,N_5655,N_7375);
and UO_1361 (O_1361,N_9208,N_6871);
nand UO_1362 (O_1362,N_8957,N_7949);
xnor UO_1363 (O_1363,N_6465,N_6551);
or UO_1364 (O_1364,N_9927,N_8298);
and UO_1365 (O_1365,N_6786,N_8673);
and UO_1366 (O_1366,N_5866,N_8554);
or UO_1367 (O_1367,N_8902,N_6878);
xnor UO_1368 (O_1368,N_9275,N_6355);
or UO_1369 (O_1369,N_9601,N_9710);
nand UO_1370 (O_1370,N_9926,N_7168);
nand UO_1371 (O_1371,N_9205,N_6012);
nand UO_1372 (O_1372,N_9482,N_9058);
and UO_1373 (O_1373,N_8802,N_8894);
and UO_1374 (O_1374,N_9353,N_9557);
nor UO_1375 (O_1375,N_9117,N_7848);
or UO_1376 (O_1376,N_6146,N_6238);
nand UO_1377 (O_1377,N_5222,N_5575);
nor UO_1378 (O_1378,N_6018,N_7021);
or UO_1379 (O_1379,N_6218,N_8629);
or UO_1380 (O_1380,N_5272,N_9302);
or UO_1381 (O_1381,N_9144,N_8352);
or UO_1382 (O_1382,N_6482,N_8532);
xor UO_1383 (O_1383,N_9280,N_8584);
or UO_1384 (O_1384,N_9999,N_5483);
or UO_1385 (O_1385,N_5221,N_7207);
and UO_1386 (O_1386,N_8234,N_7374);
nor UO_1387 (O_1387,N_5352,N_8437);
or UO_1388 (O_1388,N_5940,N_6468);
xor UO_1389 (O_1389,N_6568,N_9829);
or UO_1390 (O_1390,N_6385,N_9772);
or UO_1391 (O_1391,N_9675,N_5026);
or UO_1392 (O_1392,N_7045,N_8480);
nand UO_1393 (O_1393,N_6765,N_9452);
xor UO_1394 (O_1394,N_5194,N_9815);
and UO_1395 (O_1395,N_7961,N_5037);
and UO_1396 (O_1396,N_6017,N_6106);
or UO_1397 (O_1397,N_9220,N_7847);
nor UO_1398 (O_1398,N_7486,N_5390);
nand UO_1399 (O_1399,N_9377,N_6359);
and UO_1400 (O_1400,N_8612,N_9442);
or UO_1401 (O_1401,N_7675,N_8881);
nor UO_1402 (O_1402,N_6195,N_8961);
nor UO_1403 (O_1403,N_8834,N_9456);
nand UO_1404 (O_1404,N_5908,N_7344);
nand UO_1405 (O_1405,N_9233,N_5169);
or UO_1406 (O_1406,N_5777,N_7867);
nor UO_1407 (O_1407,N_8320,N_8526);
and UO_1408 (O_1408,N_6794,N_5591);
xor UO_1409 (O_1409,N_9494,N_9229);
and UO_1410 (O_1410,N_6241,N_7447);
nor UO_1411 (O_1411,N_8926,N_6852);
or UO_1412 (O_1412,N_6612,N_7290);
xor UO_1413 (O_1413,N_7669,N_9094);
or UO_1414 (O_1414,N_6253,N_7506);
and UO_1415 (O_1415,N_5102,N_5654);
nand UO_1416 (O_1416,N_6658,N_8043);
and UO_1417 (O_1417,N_9511,N_6761);
or UO_1418 (O_1418,N_6213,N_6646);
or UO_1419 (O_1419,N_7912,N_7523);
and UO_1420 (O_1420,N_7015,N_7007);
nand UO_1421 (O_1421,N_7769,N_5745);
or UO_1422 (O_1422,N_5524,N_6495);
nand UO_1423 (O_1423,N_5645,N_9748);
or UO_1424 (O_1424,N_6332,N_5161);
or UO_1425 (O_1425,N_6999,N_7668);
xor UO_1426 (O_1426,N_9143,N_6680);
and UO_1427 (O_1427,N_6194,N_9614);
or UO_1428 (O_1428,N_7396,N_6496);
nor UO_1429 (O_1429,N_6974,N_6925);
or UO_1430 (O_1430,N_5153,N_7298);
nand UO_1431 (O_1431,N_6874,N_6641);
nor UO_1432 (O_1432,N_7100,N_9189);
or UO_1433 (O_1433,N_8624,N_5074);
nand UO_1434 (O_1434,N_7093,N_7815);
nand UO_1435 (O_1435,N_6909,N_9921);
and UO_1436 (O_1436,N_5670,N_9574);
or UO_1437 (O_1437,N_9943,N_8736);
nor UO_1438 (O_1438,N_9812,N_5470);
nand UO_1439 (O_1439,N_6965,N_5217);
nand UO_1440 (O_1440,N_5236,N_9034);
nand UO_1441 (O_1441,N_7338,N_7425);
nor UO_1442 (O_1442,N_6143,N_5163);
or UO_1443 (O_1443,N_6743,N_7340);
or UO_1444 (O_1444,N_8270,N_8952);
nor UO_1445 (O_1445,N_7047,N_9572);
nand UO_1446 (O_1446,N_7191,N_6571);
and UO_1447 (O_1447,N_8503,N_8398);
or UO_1448 (O_1448,N_6078,N_8024);
or UO_1449 (O_1449,N_5485,N_5533);
nand UO_1450 (O_1450,N_7627,N_6587);
and UO_1451 (O_1451,N_5109,N_5937);
nor UO_1452 (O_1452,N_7926,N_7482);
and UO_1453 (O_1453,N_6407,N_8120);
nor UO_1454 (O_1454,N_6135,N_7781);
or UO_1455 (O_1455,N_6300,N_8305);
and UO_1456 (O_1456,N_5164,N_8962);
nor UO_1457 (O_1457,N_6272,N_9730);
or UO_1458 (O_1458,N_8562,N_8380);
nor UO_1459 (O_1459,N_8596,N_7831);
nor UO_1460 (O_1460,N_6940,N_9264);
and UO_1461 (O_1461,N_9880,N_8206);
xnor UO_1462 (O_1462,N_5148,N_5274);
nand UO_1463 (O_1463,N_7256,N_8017);
nand UO_1464 (O_1464,N_7813,N_6321);
nor UO_1465 (O_1465,N_8664,N_5917);
nand UO_1466 (O_1466,N_9639,N_5430);
nor UO_1467 (O_1467,N_6574,N_5288);
or UO_1468 (O_1468,N_6206,N_8496);
or UO_1469 (O_1469,N_8160,N_5110);
nor UO_1470 (O_1470,N_9093,N_8877);
and UO_1471 (O_1471,N_7614,N_5393);
and UO_1472 (O_1472,N_7109,N_5371);
or UO_1473 (O_1473,N_8415,N_8130);
xor UO_1474 (O_1474,N_9457,N_5185);
xor UO_1475 (O_1475,N_9008,N_9893);
xor UO_1476 (O_1476,N_9862,N_8620);
xor UO_1477 (O_1477,N_8211,N_8041);
or UO_1478 (O_1478,N_6456,N_6754);
or UO_1479 (O_1479,N_8640,N_9348);
and UO_1480 (O_1480,N_5759,N_9396);
nor UO_1481 (O_1481,N_8090,N_9179);
or UO_1482 (O_1482,N_9930,N_9993);
nand UO_1483 (O_1483,N_5344,N_6369);
nand UO_1484 (O_1484,N_5642,N_5584);
and UO_1485 (O_1485,N_8852,N_7304);
or UO_1486 (O_1486,N_8289,N_7624);
and UO_1487 (O_1487,N_7877,N_9902);
or UO_1488 (O_1488,N_7591,N_7404);
nor UO_1489 (O_1489,N_5197,N_7133);
nand UO_1490 (O_1490,N_8978,N_7053);
and UO_1491 (O_1491,N_5451,N_8794);
nor UO_1492 (O_1492,N_5829,N_7734);
or UO_1493 (O_1493,N_9132,N_6108);
nor UO_1494 (O_1494,N_5950,N_9214);
xor UO_1495 (O_1495,N_8981,N_9833);
nor UO_1496 (O_1496,N_5910,N_9555);
xnor UO_1497 (O_1497,N_9149,N_5963);
and UO_1498 (O_1498,N_7844,N_8759);
xnor UO_1499 (O_1499,N_8796,N_5835);
endmodule