module basic_2000_20000_2500_5_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_317,In_1114);
nor U1 (N_1,In_179,In_1597);
or U2 (N_2,In_1475,In_1433);
nand U3 (N_3,In_455,In_1363);
or U4 (N_4,In_1467,In_993);
or U5 (N_5,In_234,In_912);
nand U6 (N_6,In_1659,In_753);
nor U7 (N_7,In_1343,In_1281);
or U8 (N_8,In_1660,In_1270);
or U9 (N_9,In_1350,In_1360);
nor U10 (N_10,In_1760,In_1596);
xor U11 (N_11,In_1489,In_1492);
or U12 (N_12,In_1330,In_1058);
nand U13 (N_13,In_1059,In_1653);
nor U14 (N_14,In_1549,In_1412);
xor U15 (N_15,In_1570,In_1924);
nand U16 (N_16,In_1101,In_383);
nor U17 (N_17,In_903,In_1126);
nor U18 (N_18,In_88,In_798);
and U19 (N_19,In_23,In_1121);
nor U20 (N_20,In_118,In_123);
nand U21 (N_21,In_565,In_896);
nand U22 (N_22,In_1553,In_771);
and U23 (N_23,In_814,In_1030);
xor U24 (N_24,In_794,In_1217);
nand U25 (N_25,In_1190,In_209);
nand U26 (N_26,In_174,In_757);
and U27 (N_27,In_1630,In_1605);
and U28 (N_28,In_1174,In_508);
nand U29 (N_29,In_1451,In_1119);
nor U30 (N_30,In_1536,In_951);
xor U31 (N_31,In_297,In_1505);
and U32 (N_32,In_1872,In_342);
xnor U33 (N_33,In_458,In_572);
nor U34 (N_34,In_1538,In_1168);
nand U35 (N_35,In_779,In_167);
and U36 (N_36,In_1001,In_799);
nand U37 (N_37,In_635,In_1818);
or U38 (N_38,In_990,In_1007);
and U39 (N_39,In_1312,In_1714);
xor U40 (N_40,In_1045,In_1838);
and U41 (N_41,In_597,In_1942);
xor U42 (N_42,In_1500,In_269);
xnor U43 (N_43,In_874,In_302);
and U44 (N_44,In_1098,In_760);
nor U45 (N_45,In_1669,In_1725);
and U46 (N_46,In_228,In_644);
nand U47 (N_47,In_1971,In_950);
nand U48 (N_48,In_1140,In_1930);
xor U49 (N_49,In_414,In_92);
and U50 (N_50,In_1026,In_1895);
and U51 (N_51,In_1850,In_955);
and U52 (N_52,In_974,In_62);
or U53 (N_53,In_578,In_1667);
and U54 (N_54,In_1399,In_926);
nand U55 (N_55,In_1210,In_1532);
xor U56 (N_56,In_556,In_1198);
nor U57 (N_57,In_1994,In_493);
and U58 (N_58,In_1237,In_7);
or U59 (N_59,In_1263,In_134);
xor U60 (N_60,In_17,In_223);
nand U61 (N_61,In_1652,In_411);
nor U62 (N_62,In_720,In_1072);
and U63 (N_63,In_1783,In_322);
xor U64 (N_64,In_1046,In_312);
nor U65 (N_65,In_1593,In_1321);
xnor U66 (N_66,In_1458,In_1191);
and U67 (N_67,In_396,In_294);
nand U68 (N_68,In_1426,In_1948);
or U69 (N_69,In_1718,In_1841);
and U70 (N_70,In_830,In_1671);
or U71 (N_71,In_552,In_519);
nor U72 (N_72,In_1441,In_773);
and U73 (N_73,In_1133,In_1512);
xnor U74 (N_74,In_605,In_1209);
nand U75 (N_75,In_978,In_1583);
and U76 (N_76,In_1918,In_9);
nand U77 (N_77,In_249,In_98);
or U78 (N_78,In_1116,In_1762);
or U79 (N_79,In_1131,In_73);
xor U80 (N_80,In_1914,In_626);
nand U81 (N_81,In_1925,In_1063);
and U82 (N_82,In_1158,In_924);
or U83 (N_83,In_1529,In_1461);
or U84 (N_84,In_326,In_464);
nor U85 (N_85,In_1770,In_1787);
and U86 (N_86,In_332,In_936);
and U87 (N_87,In_283,In_106);
or U88 (N_88,In_1146,In_65);
nor U89 (N_89,In_1346,In_1581);
nand U90 (N_90,In_774,In_751);
nand U91 (N_91,In_148,In_767);
or U92 (N_92,In_1904,In_51);
or U93 (N_93,In_1956,In_1736);
nand U94 (N_94,In_178,In_1648);
and U95 (N_95,In_1229,In_1590);
nand U96 (N_96,In_1632,In_350);
nor U97 (N_97,In_1071,In_109);
and U98 (N_98,In_1528,In_1054);
or U99 (N_99,In_1917,In_660);
xnor U100 (N_100,In_1043,In_4);
nor U101 (N_101,In_369,In_1389);
nor U102 (N_102,In_226,In_1953);
or U103 (N_103,In_547,In_777);
nand U104 (N_104,In_1643,In_1662);
nor U105 (N_105,In_41,In_492);
and U106 (N_106,In_575,In_920);
nand U107 (N_107,In_522,In_1265);
nand U108 (N_108,In_1535,In_338);
nor U109 (N_109,In_1254,In_89);
and U110 (N_110,In_967,In_1816);
xnor U111 (N_111,In_207,In_314);
and U112 (N_112,In_689,In_107);
nand U113 (N_113,In_1639,In_1285);
nor U114 (N_114,In_1743,In_59);
or U115 (N_115,In_138,In_1413);
and U116 (N_116,In_393,In_275);
and U117 (N_117,In_699,In_740);
or U118 (N_118,In_169,In_186);
nor U119 (N_119,In_531,In_583);
or U120 (N_120,In_1482,In_1753);
nor U121 (N_121,In_1073,In_1738);
nor U122 (N_122,In_423,In_1393);
nor U123 (N_123,In_1913,In_797);
nor U124 (N_124,In_212,In_504);
or U125 (N_125,In_1747,In_1151);
nor U126 (N_126,In_1871,In_1849);
nand U127 (N_127,In_126,In_1852);
nand U128 (N_128,In_1523,In_888);
or U129 (N_129,In_518,In_506);
nor U130 (N_130,In_1654,In_112);
and U131 (N_131,In_1411,In_680);
and U132 (N_132,In_618,In_449);
and U133 (N_133,In_253,In_1960);
and U134 (N_134,In_282,In_1222);
xor U135 (N_135,In_673,In_1201);
or U136 (N_136,In_918,In_219);
xnor U137 (N_137,In_1839,In_1866);
nor U138 (N_138,In_1235,In_1507);
nand U139 (N_139,In_152,In_36);
and U140 (N_140,In_40,In_1641);
nor U141 (N_141,In_945,In_1349);
nor U142 (N_142,In_940,In_630);
nor U143 (N_143,In_1272,In_1701);
nor U144 (N_144,In_1796,In_1587);
nand U145 (N_145,In_1069,In_1820);
and U146 (N_146,In_70,In_1031);
xor U147 (N_147,In_239,In_670);
nor U148 (N_148,In_860,In_783);
and U149 (N_149,In_452,In_1894);
and U150 (N_150,In_588,In_1585);
xnor U151 (N_151,In_1759,In_1407);
xor U152 (N_152,In_1189,In_1092);
or U153 (N_153,In_1162,In_946);
and U154 (N_154,In_459,In_354);
nor U155 (N_155,In_1418,In_67);
nor U156 (N_156,In_1955,In_1398);
and U157 (N_157,In_574,In_1873);
xor U158 (N_158,In_1427,In_1728);
and U159 (N_159,In_410,In_966);
or U160 (N_160,In_739,In_1384);
and U161 (N_161,In_1689,In_1920);
nand U162 (N_162,In_166,In_894);
or U163 (N_163,In_272,In_1806);
and U164 (N_164,In_1685,In_127);
or U165 (N_165,In_1979,In_1315);
nand U166 (N_166,In_1809,In_1322);
nand U167 (N_167,In_1861,In_1862);
and U168 (N_168,In_1620,In_420);
nor U169 (N_169,In_1415,In_579);
nor U170 (N_170,In_535,In_1203);
and U171 (N_171,In_1491,In_346);
nand U172 (N_172,In_476,In_415);
xor U173 (N_173,In_516,In_1881);
and U174 (N_174,In_847,In_533);
nand U175 (N_175,In_840,In_1037);
nand U176 (N_176,In_1014,In_1992);
nor U177 (N_177,In_274,In_443);
nand U178 (N_178,In_745,In_215);
nand U179 (N_179,In_1288,In_560);
or U180 (N_180,In_1167,In_1338);
nand U181 (N_181,In_1601,In_996);
and U182 (N_182,In_1025,In_781);
and U183 (N_183,In_1608,In_48);
and U184 (N_184,In_204,In_1172);
or U185 (N_185,In_241,In_478);
or U186 (N_186,In_1927,In_513);
nor U187 (N_187,In_374,In_505);
nor U188 (N_188,In_1776,In_879);
nor U189 (N_189,In_431,In_378);
nor U190 (N_190,In_453,In_948);
nor U191 (N_191,In_1163,In_1661);
and U192 (N_192,In_1137,In_216);
nand U193 (N_193,In_1694,In_729);
or U194 (N_194,In_820,In_1483);
nor U195 (N_195,In_707,In_730);
nor U196 (N_196,In_1749,In_979);
or U197 (N_197,In_1291,In_975);
and U198 (N_198,In_388,In_836);
and U199 (N_199,In_5,In_1262);
and U200 (N_200,In_1958,In_614);
and U201 (N_201,In_653,In_633);
nand U202 (N_202,In_880,In_844);
nor U203 (N_203,In_1945,In_719);
nor U204 (N_204,In_1110,In_1181);
and U205 (N_205,In_698,In_1255);
nand U206 (N_206,In_1822,In_1693);
nand U207 (N_207,In_304,In_1497);
and U208 (N_208,In_1260,In_260);
nor U209 (N_209,In_1306,In_49);
nand U210 (N_210,In_617,In_684);
nand U211 (N_211,In_240,In_1637);
nand U212 (N_212,In_1865,In_1345);
and U213 (N_213,In_1365,In_538);
or U214 (N_214,In_1390,In_171);
nor U215 (N_215,In_1598,In_103);
nand U216 (N_216,In_1863,In_710);
xor U217 (N_217,In_502,In_678);
xnor U218 (N_218,In_1786,In_1604);
nor U219 (N_219,In_1655,In_746);
nand U220 (N_220,In_542,In_1323);
nor U221 (N_221,In_1253,In_532);
or U222 (N_222,In_140,In_1983);
nand U223 (N_223,In_489,In_232);
or U224 (N_224,In_1290,In_1455);
and U225 (N_225,In_1545,In_1444);
and U226 (N_226,In_79,In_922);
and U227 (N_227,In_1810,In_1353);
nor U228 (N_228,In_1859,In_733);
and U229 (N_229,In_1827,In_994);
nand U230 (N_230,In_116,In_1864);
nor U231 (N_231,In_1589,In_1594);
nand U232 (N_232,In_1831,In_1954);
and U233 (N_233,In_157,In_16);
nor U234 (N_234,In_1,In_1943);
and U235 (N_235,In_1052,In_843);
or U236 (N_236,In_1740,In_1981);
nand U237 (N_237,In_61,In_390);
and U238 (N_238,In_377,In_191);
or U239 (N_239,In_380,In_31);
and U240 (N_240,In_1554,In_1877);
and U241 (N_241,In_1664,In_984);
and U242 (N_242,In_1814,In_1846);
and U243 (N_243,In_1870,In_934);
or U244 (N_244,In_1666,In_1099);
nand U245 (N_245,In_927,In_1577);
nand U246 (N_246,In_1771,In_1261);
nand U247 (N_247,In_418,In_1949);
or U248 (N_248,In_1763,In_437);
nand U249 (N_249,In_1300,In_12);
xor U250 (N_250,In_1518,In_970);
and U251 (N_251,In_601,In_1367);
and U252 (N_252,In_756,In_1339);
and U253 (N_253,In_1517,In_1978);
xor U254 (N_254,In_1106,In_1111);
and U255 (N_255,In_1926,In_1506);
nand U256 (N_256,In_636,In_1561);
nand U257 (N_257,In_382,In_907);
nand U258 (N_258,In_355,In_463);
or U259 (N_259,In_1672,In_242);
nor U260 (N_260,In_1607,In_184);
or U261 (N_261,In_1515,In_1318);
nor U262 (N_262,In_1773,In_1085);
xnor U263 (N_263,In_1055,In_1252);
nor U264 (N_264,In_986,In_1266);
nand U265 (N_265,In_1303,In_54);
or U266 (N_266,In_567,In_663);
nor U267 (N_267,In_1094,In_192);
and U268 (N_268,In_890,In_1702);
and U269 (N_269,In_158,In_691);
nor U270 (N_270,In_99,In_982);
nor U271 (N_271,In_1813,In_1154);
and U272 (N_272,In_1298,In_938);
or U273 (N_273,In_949,In_1902);
and U274 (N_274,In_782,In_1213);
nand U275 (N_275,In_359,In_754);
nor U276 (N_276,In_858,In_24);
or U277 (N_277,In_784,In_1756);
nor U278 (N_278,In_1699,In_1020);
nand U279 (N_279,In_902,In_1478);
or U280 (N_280,In_1688,In_146);
nand U281 (N_281,In_1606,In_1023);
nand U282 (N_282,In_563,In_1774);
nand U283 (N_283,In_1991,In_941);
nor U284 (N_284,In_835,In_436);
nor U285 (N_285,In_187,In_1793);
and U286 (N_286,In_1721,In_998);
or U287 (N_287,In_473,In_743);
nor U288 (N_288,In_1004,In_392);
and U289 (N_289,In_1034,In_1205);
nand U290 (N_290,In_1680,In_1690);
nand U291 (N_291,In_457,In_1449);
or U292 (N_292,In_873,In_1892);
nand U293 (N_293,In_1980,In_1531);
and U294 (N_294,In_1769,In_884);
nor U295 (N_295,In_1602,In_251);
nor U296 (N_296,In_515,In_1388);
and U297 (N_297,In_1644,In_335);
nand U298 (N_298,In_1223,In_952);
nor U299 (N_299,In_386,In_803);
nand U300 (N_300,In_702,In_34);
nand U301 (N_301,In_1490,In_424);
nor U302 (N_302,In_685,In_1022);
and U303 (N_303,In_68,In_1086);
and U304 (N_304,In_173,In_1788);
nand U305 (N_305,In_465,In_268);
nor U306 (N_306,In_829,In_868);
nand U307 (N_307,In_1887,In_365);
nand U308 (N_308,In_1764,In_1286);
nor U309 (N_309,In_726,In_1999);
nand U310 (N_310,In_399,In_400);
nand U311 (N_311,In_105,In_641);
nand U312 (N_312,In_75,In_885);
and U313 (N_313,In_168,In_227);
or U314 (N_314,In_1469,In_557);
and U315 (N_315,In_1921,In_1567);
nand U316 (N_316,In_748,In_1432);
nand U317 (N_317,In_1867,In_1599);
and U318 (N_318,In_855,In_682);
xor U319 (N_319,In_1334,In_1293);
nor U320 (N_320,In_1546,In_724);
nor U321 (N_321,In_1362,In_247);
nand U322 (N_322,In_637,In_1000);
xnor U323 (N_323,In_429,In_1784);
nand U324 (N_324,In_992,In_1485);
xnor U325 (N_325,In_577,In_706);
and U326 (N_326,In_1778,In_1647);
nand U327 (N_327,In_1898,In_183);
and U328 (N_328,In_1963,In_143);
or U329 (N_329,In_159,In_1275);
xnor U330 (N_330,In_1615,In_1143);
nor U331 (N_331,In_156,In_1132);
nand U332 (N_332,In_133,In_1805);
or U333 (N_333,In_276,In_1910);
or U334 (N_334,In_401,In_703);
nand U335 (N_335,In_1215,In_82);
nand U336 (N_336,In_839,In_363);
nand U337 (N_337,In_1424,In_715);
or U338 (N_338,In_1170,In_737);
nand U339 (N_339,In_91,In_46);
or U340 (N_340,In_1193,In_1501);
or U341 (N_341,In_1468,In_1595);
or U342 (N_342,In_1611,In_1442);
nor U343 (N_343,In_687,In_14);
xor U344 (N_344,In_122,In_1840);
nand U345 (N_345,In_664,In_600);
nor U346 (N_346,In_1320,In_819);
nand U347 (N_347,In_1027,In_1618);
or U348 (N_348,In_433,In_701);
or U349 (N_349,In_182,In_408);
nor U350 (N_350,In_915,In_944);
xnor U351 (N_351,In_1988,In_370);
or U352 (N_352,In_877,In_1516);
and U353 (N_353,In_288,In_1123);
and U354 (N_354,In_1640,In_86);
nor U355 (N_355,In_499,In_1387);
and U356 (N_356,In_1800,In_1421);
nor U357 (N_357,In_278,In_1480);
or U358 (N_358,In_307,In_395);
xor U359 (N_359,In_1136,In_435);
or U360 (N_360,In_235,In_765);
and U361 (N_361,In_570,In_1259);
nor U362 (N_362,In_980,In_988);
or U363 (N_363,In_1161,In_1541);
nand U364 (N_364,In_149,In_805);
or U365 (N_365,In_202,In_717);
nand U366 (N_366,In_1856,In_1066);
or U367 (N_367,In_898,In_1206);
and U368 (N_368,In_1834,In_1155);
nand U369 (N_369,In_576,In_1623);
or U370 (N_370,In_1445,In_284);
nand U371 (N_371,In_199,In_1473);
nand U372 (N_372,In_1704,In_1488);
and U373 (N_373,In_1804,In_658);
or U374 (N_374,In_971,In_872);
or U375 (N_375,In_336,In_554);
nand U376 (N_376,In_1931,In_1588);
nand U377 (N_377,In_190,In_1765);
or U378 (N_378,In_325,In_1208);
nor U379 (N_379,In_806,In_1038);
and U380 (N_380,In_1571,In_18);
nand U381 (N_381,In_841,In_1893);
and U382 (N_382,In_1896,In_609);
nand U383 (N_383,In_1200,In_1417);
and U384 (N_384,In_366,In_1044);
nand U385 (N_385,In_1267,In_1651);
or U386 (N_386,In_968,In_1157);
nor U387 (N_387,In_1295,In_1354);
or U388 (N_388,In_645,In_1533);
or U389 (N_389,In_1646,In_1876);
or U390 (N_390,In_863,In_709);
xor U391 (N_391,In_900,In_1083);
nand U392 (N_392,In_56,In_195);
nor U393 (N_393,In_323,In_571);
and U394 (N_394,In_104,In_889);
and U395 (N_395,In_875,In_813);
nand U396 (N_396,In_842,In_521);
or U397 (N_397,In_947,In_1744);
nand U398 (N_398,In_921,In_1745);
nor U399 (N_399,In_1269,In_1720);
and U400 (N_400,In_237,In_705);
xnor U401 (N_401,In_1150,In_1499);
and U402 (N_402,In_1629,In_1122);
or U403 (N_403,In_1544,In_120);
nand U404 (N_404,In_1368,In_1068);
xor U405 (N_405,In_1974,In_150);
or U406 (N_406,In_1177,In_624);
or U407 (N_407,In_1730,In_77);
and U408 (N_408,In_965,In_1657);
or U409 (N_409,In_1767,In_1803);
nor U410 (N_410,In_1186,In_320);
or U411 (N_411,In_481,In_1821);
and U412 (N_412,In_44,In_591);
and U413 (N_413,In_1328,In_1591);
and U414 (N_414,In_1246,In_1359);
nand U415 (N_415,In_511,In_1957);
xor U416 (N_416,In_1586,In_80);
xor U417 (N_417,In_1837,In_1542);
and U418 (N_418,In_50,In_160);
and U419 (N_419,In_1732,In_356);
and U420 (N_420,In_1946,In_914);
nor U421 (N_421,In_1982,In_594);
and U422 (N_422,In_662,In_931);
and U423 (N_423,In_826,In_727);
nor U424 (N_424,In_389,In_1279);
nor U425 (N_425,In_527,In_238);
nand U426 (N_426,In_1224,In_486);
nor U427 (N_427,In_211,In_642);
or U428 (N_428,In_1551,In_1975);
nor U429 (N_429,In_1755,In_52);
nor U430 (N_430,In_95,In_1450);
and U431 (N_431,In_290,In_1335);
xnor U432 (N_432,In_891,In_593);
or U433 (N_433,In_1324,In_289);
and U434 (N_434,In_1997,In_1088);
and U435 (N_435,In_1080,In_913);
nand U436 (N_436,In_744,In_1479);
and U437 (N_437,In_1232,In_677);
xor U438 (N_438,In_1051,In_280);
nor U439 (N_439,In_1248,In_1722);
and U440 (N_440,In_1989,In_1560);
nor U441 (N_441,In_259,In_291);
or U442 (N_442,In_1204,In_1076);
or U443 (N_443,In_544,In_964);
xnor U444 (N_444,In_1698,In_1860);
or U445 (N_445,In_1453,In_1886);
and U446 (N_446,In_582,In_1668);
nand U447 (N_447,In_1405,In_1011);
nor U448 (N_448,In_419,In_1337);
and U449 (N_449,In_611,In_295);
and U450 (N_450,In_1264,In_66);
and U451 (N_451,In_845,In_960);
xor U452 (N_452,In_758,In_1679);
nand U453 (N_453,In_1798,In_1302);
nor U454 (N_454,In_848,In_1711);
and U455 (N_455,In_1716,In_1525);
and U456 (N_456,In_1178,In_1826);
nand U457 (N_457,In_1683,In_585);
nor U458 (N_458,In_1018,In_517);
xnor U459 (N_459,In_1152,In_1401);
nor U460 (N_460,In_1195,In_1230);
or U461 (N_461,In_1416,In_460);
and U462 (N_462,In_243,In_1304);
or U463 (N_463,In_1127,In_904);
or U464 (N_464,In_1642,In_1187);
and U465 (N_465,In_1677,In_57);
or U466 (N_466,In_1117,In_1100);
nor U467 (N_467,In_1289,In_808);
nand U468 (N_468,In_590,In_1906);
nand U469 (N_469,In_222,In_221);
or U470 (N_470,In_824,In_524);
nand U471 (N_471,In_1364,In_1105);
or U472 (N_472,In_541,In_318);
nor U473 (N_473,In_22,In_1638);
nand U474 (N_474,In_1656,In_1658);
and U475 (N_475,In_1142,In_732);
nor U476 (N_476,In_1096,In_1258);
nand U477 (N_477,In_333,In_749);
and U478 (N_478,In_1282,In_1236);
xnor U479 (N_479,In_634,In_1169);
and U480 (N_480,In_244,In_1240);
nor U481 (N_481,In_8,In_1568);
nor U482 (N_482,In_1875,In_804);
nor U483 (N_483,In_200,In_1373);
or U484 (N_484,In_1292,In_19);
nand U485 (N_485,In_876,In_1268);
nand U486 (N_486,In_1294,In_387);
or U487 (N_487,In_612,In_456);
and U488 (N_488,In_113,In_321);
or U489 (N_489,In_1890,In_1634);
or U490 (N_490,In_831,In_997);
nand U491 (N_491,In_1428,In_1251);
xnor U492 (N_492,In_654,In_925);
nand U493 (N_493,In_53,In_853);
nand U494 (N_494,In_397,In_287);
and U495 (N_495,In_621,In_1650);
nor U496 (N_496,In_257,In_514);
and U497 (N_497,In_1029,In_33);
or U498 (N_498,In_1496,In_859);
nor U499 (N_499,In_164,In_1392);
and U500 (N_500,In_716,In_1884);
xnor U501 (N_501,In_752,In_1211);
xnor U502 (N_502,In_647,In_769);
or U503 (N_503,In_1508,In_627);
nand U504 (N_504,In_483,In_327);
and U505 (N_505,In_1278,In_728);
nor U506 (N_506,In_1357,In_1848);
nand U507 (N_507,In_638,In_85);
nand U508 (N_508,In_1919,In_1218);
nand U509 (N_509,In_650,In_543);
nand U510 (N_510,In_755,In_38);
nor U511 (N_511,In_973,In_405);
nor U512 (N_512,In_1868,In_115);
or U513 (N_513,In_181,In_1514);
and U514 (N_514,In_602,In_163);
nor U515 (N_515,In_1998,In_1002);
or U516 (N_516,In_1828,In_683);
nand U517 (N_517,In_1574,In_250);
or U518 (N_518,In_1443,In_1534);
and U519 (N_519,In_1234,In_629);
nor U520 (N_520,In_1673,In_428);
nor U521 (N_521,In_137,In_1422);
nand U522 (N_522,In_675,In_151);
nor U523 (N_523,In_766,In_1336);
nor U524 (N_524,In_610,In_1527);
and U525 (N_525,In_549,In_265);
and U526 (N_526,In_1352,In_1436);
nor U527 (N_527,In_1737,In_1340);
or U528 (N_528,In_1437,In_398);
nand U529 (N_529,In_1703,In_296);
xnor U530 (N_530,In_1857,In_787);
and U531 (N_531,In_1273,In_26);
nor U532 (N_532,In_895,In_1179);
xor U533 (N_533,In_792,In_1039);
or U534 (N_534,In_1792,In_1062);
nor U535 (N_535,In_991,In_281);
and U536 (N_536,In_529,In_1880);
nor U537 (N_537,In_1325,In_110);
and U538 (N_538,In_1540,In_1103);
or U539 (N_539,In_1844,In_339);
nand U540 (N_540,In_1274,In_1410);
nor U541 (N_541,In_1802,In_1299);
nand U542 (N_542,In_679,In_1015);
nor U543 (N_543,In_484,In_987);
and U544 (N_544,In_362,In_1462);
or U545 (N_545,In_1610,In_248);
nor U546 (N_546,In_1874,In_1090);
or U547 (N_547,In_1612,In_775);
nor U548 (N_548,In_1510,In_1681);
nor U549 (N_549,In_451,In_1952);
nor U550 (N_550,In_796,In_1125);
nor U551 (N_551,In_1724,In_81);
and U552 (N_552,In_738,In_285);
nand U553 (N_553,In_555,In_919);
or U554 (N_554,In_871,In_1056);
or U555 (N_555,In_580,In_933);
and U556 (N_556,In_1735,In_343);
xnor U557 (N_557,In_1907,In_210);
and U558 (N_558,In_1696,In_194);
and U559 (N_559,In_1326,In_1909);
nand U560 (N_560,In_640,In_330);
nand U561 (N_561,In_1276,In_213);
xnor U562 (N_562,In_1041,In_1130);
xnor U563 (N_563,In_1556,In_381);
xor U564 (N_564,In_1021,In_334);
or U565 (N_565,In_932,In_1578);
nor U566 (N_566,In_1959,In_1562);
nor U567 (N_567,In_1042,In_25);
or U568 (N_568,In_1375,In_537);
and U569 (N_569,In_1040,In_1242);
nor U570 (N_570,In_1341,In_929);
xor U571 (N_571,In_1727,In_1145);
and U572 (N_572,In_1635,In_1962);
or U573 (N_573,In_1391,In_1329);
nor U574 (N_574,In_1897,In_862);
nor U575 (N_575,In_669,In_1513);
and U576 (N_576,In_1751,In_1032);
nand U577 (N_577,In_957,In_1383);
nand U578 (N_578,In_293,In_185);
or U579 (N_579,In_1082,In_488);
or U580 (N_580,In_731,In_1148);
nor U581 (N_581,In_1617,In_64);
or U582 (N_582,In_309,In_801);
and U583 (N_583,In_963,In_1385);
nand U584 (N_584,In_1616,In_1366);
nand U585 (N_585,In_1879,In_1457);
or U586 (N_586,In_692,In_1511);
and U587 (N_587,In_1757,In_1790);
and U588 (N_588,In_1456,In_1710);
and U589 (N_589,In_1582,In_1627);
and U590 (N_590,In_656,In_1081);
and U591 (N_591,In_1319,In_1214);
nor U592 (N_592,In_1951,In_1882);
or U593 (N_593,In_972,In_214);
xnor U594 (N_594,In_292,In_651);
or U595 (N_595,In_208,In_426);
or U596 (N_596,In_1091,In_909);
or U597 (N_597,In_1746,In_1067);
nor U598 (N_598,In_131,In_407);
nand U599 (N_599,In_1915,In_661);
nand U600 (N_600,In_1579,In_1376);
nor U601 (N_601,In_416,In_1309);
xnor U602 (N_602,In_1471,In_1280);
nand U603 (N_603,In_300,In_1853);
nand U604 (N_604,In_1645,In_599);
nand U605 (N_605,In_1878,In_795);
and U606 (N_606,In_316,In_6);
and U607 (N_607,In_121,In_534);
and U608 (N_608,In_220,In_911);
xnor U609 (N_609,In_1079,In_72);
or U610 (N_610,In_1128,In_956);
xor U611 (N_611,In_1719,In_849);
nand U612 (N_612,In_1316,In_646);
nand U613 (N_613,In_1928,In_1372);
nand U614 (N_614,In_135,In_434);
or U615 (N_615,In_1912,In_1308);
or U616 (N_616,In_595,In_403);
nor U617 (N_617,In_1521,In_1761);
or U618 (N_618,In_800,In_1937);
and U619 (N_619,In_319,In_180);
nor U620 (N_620,In_84,In_1207);
xnor U621 (N_621,In_937,In_1939);
or U622 (N_622,In_1048,In_832);
or U623 (N_623,In_1519,In_613);
xnor U624 (N_624,In_114,In_1271);
and U625 (N_625,In_1386,In_856);
and U626 (N_626,In_1903,In_1494);
or U627 (N_627,In_1563,In_1592);
or U628 (N_628,In_551,In_1228);
nand U629 (N_629,In_1758,In_1734);
xnor U630 (N_630,In_1972,In_141);
and U631 (N_631,In_1369,In_1819);
and U632 (N_632,In_1687,In_1183);
xor U633 (N_633,In_21,In_1911);
nand U634 (N_634,In_1970,In_976);
and U635 (N_635,In_1219,In_144);
or U636 (N_636,In_1194,In_1074);
nand U637 (N_637,In_1923,In_850);
nand U638 (N_638,In_203,In_943);
and U639 (N_639,In_1922,In_604);
xor U640 (N_640,In_286,In_893);
xnor U641 (N_641,In_422,In_596);
nor U642 (N_642,In_768,In_1481);
nor U643 (N_643,In_1397,In_545);
nor U644 (N_644,In_353,In_1284);
nand U645 (N_645,In_802,In_111);
nor U646 (N_646,In_495,In_1509);
nand U647 (N_647,In_1631,In_1564);
or U648 (N_648,In_759,In_550);
and U649 (N_649,In_119,In_480);
or U650 (N_650,In_1739,In_1869);
nor U651 (N_651,In_477,In_1750);
nor U652 (N_652,In_1394,In_1305);
xor U653 (N_653,In_854,In_252);
or U654 (N_654,In_1371,In_1768);
nand U655 (N_655,In_245,In_461);
and U656 (N_656,In_1192,In_1414);
nor U657 (N_657,In_1486,In_197);
nor U658 (N_658,In_357,In_261);
nand U659 (N_659,In_985,In_899);
and U660 (N_660,In_1573,In_867);
and U661 (N_661,In_29,In_1139);
and U662 (N_662,In_175,In_977);
nor U663 (N_663,In_466,In_1257);
nor U664 (N_664,In_1916,In_823);
nand U665 (N_665,In_553,In_1985);
or U666 (N_666,In_468,In_812);
or U667 (N_667,In_1377,In_35);
or U668 (N_668,In_1780,In_45);
nand U669 (N_669,In_1692,In_1019);
xnor U670 (N_670,In_643,In_1093);
nor U671 (N_671,In_995,In_1212);
nand U672 (N_672,In_0,In_470);
nor U673 (N_673,In_1855,In_1256);
nor U674 (N_674,In_712,In_1754);
or U675 (N_675,In_87,In_1695);
and U676 (N_676,In_454,In_983);
nand U677 (N_677,In_1811,In_1966);
and U678 (N_678,In_901,In_402);
and U679 (N_679,In_368,In_345);
and U680 (N_680,In_562,In_540);
and U681 (N_681,In_625,In_1547);
or U682 (N_682,In_791,In_1842);
xor U683 (N_683,In_1995,In_421);
xor U684 (N_684,In_1166,In_1682);
nor U685 (N_685,In_1008,In_676);
nor U686 (N_686,In_1171,In_564);
or U687 (N_687,In_1459,In_818);
nand U688 (N_688,In_1188,In_1454);
and U689 (N_689,In_1439,In_189);
nor U690 (N_690,In_721,In_432);
nand U691 (N_691,In_1057,In_1824);
nor U692 (N_692,In_1565,In_1539);
nand U693 (N_693,In_1566,In_1815);
and U694 (N_694,In_878,In_1996);
and U695 (N_695,In_1987,In_816);
and U696 (N_696,In_1580,In_263);
or U697 (N_697,In_865,In_404);
or U698 (N_698,In_916,In_303);
nor U699 (N_699,In_217,In_828);
nor U700 (N_700,In_711,In_1708);
nand U701 (N_701,In_11,In_1107);
nor U702 (N_702,In_1470,In_623);
nand U703 (N_703,In_1314,In_1944);
and U704 (N_704,In_1498,In_267);
xor U705 (N_705,In_1231,In_1900);
or U706 (N_706,In_1141,In_1851);
and U707 (N_707,In_747,In_559);
or U708 (N_708,In_905,In_1452);
or U709 (N_709,In_1466,In_693);
nand U710 (N_710,In_1726,In_236);
and U711 (N_711,In_1569,In_581);
and U712 (N_712,In_1986,In_1609);
or U713 (N_713,In_1238,In_101);
nor U714 (N_714,In_1408,In_1173);
nand U715 (N_715,In_1526,In_1197);
and U716 (N_716,In_546,In_1670);
xnor U717 (N_717,In_1016,In_1239);
or U718 (N_718,In_1147,In_311);
nor U719 (N_719,In_231,In_1164);
nand U720 (N_720,In_20,In_1313);
and U721 (N_721,In_1835,In_526);
xor U722 (N_722,In_1003,In_352);
xor U723 (N_723,In_1120,In_1036);
or U724 (N_724,In_1403,In_681);
and U725 (N_725,In_851,In_1938);
or U726 (N_726,In_439,In_1794);
or U727 (N_727,In_30,In_1487);
and U728 (N_728,In_385,In_1296);
xnor U729 (N_729,In_1005,In_652);
nand U730 (N_730,In_999,In_1358);
and U731 (N_731,In_1775,In_351);
nand U732 (N_732,In_358,In_445);
nor U733 (N_733,In_379,In_1138);
xor U734 (N_734,In_373,In_1785);
nor U735 (N_735,In_1446,In_628);
nand U736 (N_736,In_1250,In_723);
xnor U737 (N_737,In_349,In_615);
xnor U738 (N_738,In_908,In_881);
nand U739 (N_739,In_1572,In_224);
nor U740 (N_740,In_954,In_60);
nand U741 (N_741,In_258,In_1676);
nand U742 (N_742,In_299,In_128);
nand U743 (N_743,In_935,In_742);
nor U744 (N_744,In_1817,In_132);
xnor U745 (N_745,In_472,In_376);
and U746 (N_746,In_736,In_97);
nor U747 (N_747,In_1899,In_1176);
or U748 (N_748,In_923,In_15);
and U749 (N_749,In_942,In_1115);
or U750 (N_750,In_1060,In_1012);
or U751 (N_751,In_273,In_530);
or U752 (N_752,In_1748,In_1713);
or U753 (N_753,In_427,In_384);
or U754 (N_754,In_1216,In_866);
nand U755 (N_755,In_498,In_469);
nand U756 (N_756,In_145,In_1409);
nor U757 (N_757,In_1400,In_485);
or U758 (N_758,In_308,In_1182);
or U759 (N_759,In_1976,In_827);
and U760 (N_760,In_1477,In_1777);
nand U761 (N_761,In_1752,In_1889);
and U762 (N_762,In_474,In_1244);
xnor U763 (N_763,In_1050,In_76);
and U764 (N_764,In_1932,In_409);
nand U765 (N_765,In_558,In_930);
nor U766 (N_766,In_1493,In_1520);
or U767 (N_767,In_838,In_1883);
nor U768 (N_768,In_1077,In_1124);
xnor U769 (N_769,In_310,In_587);
nor U770 (N_770,In_1772,In_603);
and U771 (N_771,In_83,In_32);
or U772 (N_772,In_667,In_266);
and U773 (N_773,In_1782,In_1965);
nand U774 (N_774,In_1557,In_1287);
nor U775 (N_775,In_188,In_989);
nor U776 (N_776,In_479,In_1307);
nand U777 (N_777,In_10,In_1552);
nand U778 (N_778,In_704,In_1731);
or U779 (N_779,In_1331,In_834);
and U780 (N_780,In_1700,In_1064);
nand U781 (N_781,In_1355,In_1382);
nand U782 (N_782,In_1799,In_833);
or U783 (N_783,In_510,In_1984);
and U784 (N_784,In_569,In_837);
or U785 (N_785,In_1430,In_1543);
nand U786 (N_786,In_1901,In_1614);
or U787 (N_787,In_655,In_1344);
xor U788 (N_788,In_1075,In_1706);
nand U789 (N_789,In_139,In_776);
and U790 (N_790,In_298,In_1404);
xnor U791 (N_791,In_153,In_1440);
nor U792 (N_792,In_674,In_1283);
and U793 (N_793,In_807,In_1626);
nand U794 (N_794,In_1277,In_1061);
nor U795 (N_795,In_525,In_697);
or U796 (N_796,In_1102,In_1327);
nor U797 (N_797,In_1600,In_1435);
and U798 (N_798,In_406,In_1812);
nand U799 (N_799,In_1709,In_566);
nor U800 (N_800,In_93,In_1797);
nor U801 (N_801,In_1808,In_198);
and U802 (N_802,In_136,In_616);
nand U803 (N_803,In_620,In_28);
nor U804 (N_804,In_1829,In_969);
or U805 (N_805,In_607,In_1396);
nor U806 (N_806,In_1245,In_1636);
nor U807 (N_807,In_361,In_1233);
or U808 (N_808,In_959,In_1220);
nand U809 (N_809,In_1613,In_344);
nand U810 (N_810,In_1625,In_864);
nor U811 (N_811,In_255,In_1993);
and U812 (N_812,In_447,In_785);
nor U813 (N_813,In_1947,In_55);
nor U814 (N_814,In_962,In_1537);
xnor U815 (N_815,In_1049,In_718);
nand U816 (N_816,In_225,In_1463);
and U817 (N_817,In_1108,In_869);
and U818 (N_818,In_196,In_1033);
xnor U819 (N_819,In_78,In_1584);
and U820 (N_820,In_825,In_649);
nand U821 (N_821,In_1503,In_1196);
and U822 (N_822,In_1144,In_47);
xor U823 (N_823,In_857,In_130);
nor U824 (N_824,In_1202,In_1933);
or U825 (N_825,In_1941,In_573);
or U826 (N_826,In_665,In_500);
and U827 (N_827,In_817,In_561);
or U828 (N_828,In_391,In_1495);
or U829 (N_829,In_301,In_1833);
nand U830 (N_830,In_1185,In_1502);
or U831 (N_831,In_124,In_1665);
and U832 (N_832,In_1789,In_1697);
or U833 (N_833,In_981,In_176);
or U834 (N_834,In_441,In_1830);
or U835 (N_835,In_786,In_846);
nand U836 (N_836,In_1379,In_1097);
and U837 (N_837,In_446,In_1447);
or U838 (N_838,In_341,In_939);
nand U839 (N_839,In_230,In_165);
and U840 (N_840,In_1741,In_1576);
or U841 (N_841,In_622,In_1402);
nor U842 (N_842,In_958,In_793);
nor U843 (N_843,In_1301,In_1766);
and U844 (N_844,In_1973,In_328);
nand U845 (N_845,In_1065,In_1156);
nor U846 (N_846,In_467,In_100);
and U847 (N_847,In_1950,In_1429);
and U848 (N_848,In_1622,In_1929);
nand U849 (N_849,In_1675,In_1243);
or U850 (N_850,In_490,In_725);
nand U851 (N_851,In_1089,In_735);
and U852 (N_852,In_367,In_440);
xnor U853 (N_853,In_598,In_523);
and U854 (N_854,In_1686,In_1420);
nand U855 (N_855,In_1836,In_425);
or U856 (N_856,In_619,In_1791);
nor U857 (N_857,In_694,In_394);
or U858 (N_858,In_13,In_58);
nand U859 (N_859,In_74,In_1555);
nor U860 (N_860,In_741,In_471);
nor U861 (N_861,In_917,In_1153);
and U862 (N_862,In_1425,In_1180);
and U863 (N_863,In_444,In_501);
nand U864 (N_864,In_539,In_313);
xor U865 (N_865,In_448,In_1715);
xor U866 (N_866,In_1964,In_375);
or U867 (N_867,In_331,In_1548);
or U868 (N_868,In_1227,In_1832);
or U869 (N_869,In_883,In_659);
and U870 (N_870,In_708,In_360);
and U871 (N_871,In_206,In_1843);
and U872 (N_872,In_1522,In_329);
nor U873 (N_873,In_155,In_1333);
or U874 (N_874,In_700,In_102);
xor U875 (N_875,In_347,In_306);
or U876 (N_876,In_1717,In_1225);
or U877 (N_877,In_372,In_1199);
nand U878 (N_878,In_1524,In_1504);
or U879 (N_879,In_1013,In_1342);
nor U880 (N_880,In_1370,In_1129);
xnor U881 (N_881,In_1633,In_27);
and U882 (N_882,In_277,In_1035);
or U883 (N_883,In_170,In_475);
or U884 (N_884,In_1559,In_348);
or U885 (N_885,In_690,In_1484);
nor U886 (N_886,In_1807,In_509);
nor U887 (N_887,In_1084,In_1112);
or U888 (N_888,In_1530,In_695);
nand U889 (N_889,In_906,In_897);
nand U890 (N_890,In_1460,In_1977);
nor U891 (N_891,In_1221,In_305);
xor U892 (N_892,In_1165,In_1712);
or U893 (N_893,In_1311,In_1801);
nor U894 (N_894,In_1705,In_71);
nor U895 (N_895,In_1474,In_1184);
nand U896 (N_896,In_672,In_442);
and U897 (N_897,In_1135,In_668);
nor U898 (N_898,In_928,In_1347);
nor U899 (N_899,In_1047,In_1649);
xnor U900 (N_900,In_686,In_688);
nand U901 (N_901,In_90,In_494);
and U902 (N_902,In_1723,In_666);
or U903 (N_903,In_790,In_1226);
and U904 (N_904,In_1348,In_910);
nor U905 (N_905,In_315,In_584);
and U906 (N_906,In_772,In_496);
nand U907 (N_907,In_1053,In_172);
nand U908 (N_908,In_1908,In_271);
and U909 (N_909,In_608,In_1619);
nand U910 (N_910,In_770,In_254);
nand U911 (N_911,In_125,In_671);
nor U912 (N_912,In_1476,In_1159);
nor U913 (N_913,In_512,In_780);
nand U914 (N_914,In_1017,In_788);
and U915 (N_915,In_1009,In_1885);
or U916 (N_916,In_507,In_1678);
or U917 (N_917,In_94,In_1663);
nor U918 (N_918,In_1380,In_37);
xnor U919 (N_919,In_337,In_43);
nor U920 (N_920,In_3,In_1472);
or U921 (N_921,In_632,In_1733);
nand U922 (N_922,In_63,In_810);
nor U923 (N_923,In_1742,In_568);
or U924 (N_924,In_887,In_1078);
nor U925 (N_925,In_364,In_734);
and U926 (N_926,In_1558,In_108);
nand U927 (N_927,In_696,In_592);
and U928 (N_928,In_1448,In_1940);
or U929 (N_929,In_1550,In_482);
nor U930 (N_930,In_861,In_417);
nand U931 (N_931,In_1113,In_1781);
or U932 (N_932,In_892,In_69);
nor U933 (N_933,In_1104,In_1935);
xor U934 (N_934,In_1351,In_1825);
and U935 (N_935,In_487,In_450);
and U936 (N_936,In_1241,In_1028);
xor U937 (N_937,In_1006,In_1575);
or U938 (N_938,In_1149,In_1674);
nor U939 (N_939,In_229,In_961);
and U940 (N_940,In_177,In_1024);
nand U941 (N_941,In_39,In_1374);
nand U942 (N_942,In_1419,In_1967);
nand U943 (N_943,In_1888,In_648);
nand U944 (N_944,In_1332,In_1464);
nand U945 (N_945,In_1823,In_1691);
and U946 (N_946,In_201,In_1779);
or U947 (N_947,In_520,In_714);
xnor U948 (N_948,In_42,In_1356);
or U949 (N_949,In_497,In_1684);
or U950 (N_950,In_96,In_882);
nand U951 (N_951,In_1905,In_1990);
nand U952 (N_952,In_142,In_536);
and U953 (N_953,In_870,In_953);
or U954 (N_954,In_606,In_162);
nor U955 (N_955,In_270,In_1406);
or U956 (N_956,In_503,In_1628);
nand U957 (N_957,In_279,In_256);
or U958 (N_958,In_1118,In_815);
nand U959 (N_959,In_639,In_1729);
and U960 (N_960,In_1795,In_246);
or U961 (N_961,In_811,In_1095);
nor U962 (N_962,In_1624,In_761);
nand U963 (N_963,In_1247,In_430);
nor U964 (N_964,In_822,In_218);
nand U965 (N_965,In_589,In_1317);
nor U966 (N_966,In_1936,In_1423);
nand U967 (N_967,In_548,In_1361);
and U968 (N_968,In_1381,In_809);
or U969 (N_969,In_1465,In_1707);
nand U970 (N_970,In_324,In_750);
nand U971 (N_971,In_2,In_657);
nor U972 (N_972,In_722,In_1845);
and U973 (N_973,In_1010,In_154);
nand U974 (N_974,In_161,In_886);
nor U975 (N_975,In_264,In_1969);
and U976 (N_976,In_821,In_1891);
and U977 (N_977,In_528,In_1621);
nand U978 (N_978,In_1070,In_205);
nand U979 (N_979,In_1378,In_129);
nand U980 (N_980,In_1175,In_1854);
xor U981 (N_981,In_1934,In_412);
or U982 (N_982,In_1310,In_491);
nor U983 (N_983,In_233,In_1847);
nor U984 (N_984,In_764,In_789);
or U985 (N_985,In_1961,In_1160);
nand U986 (N_986,In_631,In_1134);
and U987 (N_987,In_778,In_762);
and U988 (N_988,In_713,In_413);
nand U989 (N_989,In_1109,In_1603);
or U990 (N_990,In_1858,In_1968);
and U991 (N_991,In_1249,In_438);
or U992 (N_992,In_1434,In_586);
nor U993 (N_993,In_462,In_1431);
or U994 (N_994,In_147,In_1087);
nor U995 (N_995,In_117,In_1395);
nand U996 (N_996,In_340,In_1297);
nand U997 (N_997,In_371,In_1438);
nand U998 (N_998,In_193,In_852);
nor U999 (N_999,In_763,In_262);
and U1000 (N_1000,In_1608,In_1992);
xor U1001 (N_1001,In_851,In_958);
nor U1002 (N_1002,In_42,In_254);
or U1003 (N_1003,In_1941,In_392);
and U1004 (N_1004,In_307,In_773);
or U1005 (N_1005,In_990,In_1432);
and U1006 (N_1006,In_549,In_980);
and U1007 (N_1007,In_753,In_592);
and U1008 (N_1008,In_1898,In_1476);
or U1009 (N_1009,In_1594,In_1123);
xnor U1010 (N_1010,In_1078,In_1937);
nand U1011 (N_1011,In_715,In_1856);
or U1012 (N_1012,In_270,In_1291);
and U1013 (N_1013,In_1587,In_879);
and U1014 (N_1014,In_297,In_516);
nand U1015 (N_1015,In_1497,In_1097);
and U1016 (N_1016,In_858,In_296);
or U1017 (N_1017,In_1816,In_514);
nor U1018 (N_1018,In_420,In_142);
or U1019 (N_1019,In_1405,In_540);
or U1020 (N_1020,In_1535,In_101);
and U1021 (N_1021,In_1836,In_826);
or U1022 (N_1022,In_1775,In_850);
nand U1023 (N_1023,In_778,In_349);
nand U1024 (N_1024,In_63,In_1116);
or U1025 (N_1025,In_1698,In_1378);
or U1026 (N_1026,In_1256,In_928);
nor U1027 (N_1027,In_1129,In_819);
and U1028 (N_1028,In_818,In_544);
and U1029 (N_1029,In_1971,In_633);
xor U1030 (N_1030,In_1836,In_362);
nand U1031 (N_1031,In_20,In_1281);
or U1032 (N_1032,In_335,In_481);
nor U1033 (N_1033,In_660,In_581);
and U1034 (N_1034,In_292,In_547);
nor U1035 (N_1035,In_1344,In_1636);
xnor U1036 (N_1036,In_1627,In_519);
nand U1037 (N_1037,In_561,In_791);
or U1038 (N_1038,In_310,In_951);
or U1039 (N_1039,In_1227,In_1339);
nand U1040 (N_1040,In_1894,In_553);
or U1041 (N_1041,In_1832,In_628);
and U1042 (N_1042,In_153,In_1036);
nand U1043 (N_1043,In_554,In_238);
and U1044 (N_1044,In_961,In_822);
nand U1045 (N_1045,In_1577,In_609);
and U1046 (N_1046,In_786,In_639);
and U1047 (N_1047,In_220,In_301);
or U1048 (N_1048,In_277,In_1403);
xor U1049 (N_1049,In_1746,In_460);
and U1050 (N_1050,In_298,In_615);
nand U1051 (N_1051,In_1867,In_1978);
nand U1052 (N_1052,In_1901,In_508);
and U1053 (N_1053,In_1590,In_1045);
and U1054 (N_1054,In_1243,In_1317);
and U1055 (N_1055,In_724,In_1587);
xor U1056 (N_1056,In_1925,In_149);
nand U1057 (N_1057,In_1209,In_658);
or U1058 (N_1058,In_1397,In_804);
nand U1059 (N_1059,In_926,In_1896);
or U1060 (N_1060,In_1651,In_419);
nor U1061 (N_1061,In_667,In_1594);
and U1062 (N_1062,In_336,In_742);
or U1063 (N_1063,In_843,In_1976);
nor U1064 (N_1064,In_1232,In_417);
or U1065 (N_1065,In_311,In_589);
or U1066 (N_1066,In_1829,In_1699);
xnor U1067 (N_1067,In_623,In_1659);
nor U1068 (N_1068,In_1821,In_1257);
nor U1069 (N_1069,In_1843,In_1873);
and U1070 (N_1070,In_678,In_410);
xor U1071 (N_1071,In_1541,In_82);
or U1072 (N_1072,In_243,In_1516);
and U1073 (N_1073,In_354,In_399);
and U1074 (N_1074,In_232,In_1738);
nor U1075 (N_1075,In_1080,In_1794);
and U1076 (N_1076,In_974,In_682);
or U1077 (N_1077,In_1618,In_1977);
nor U1078 (N_1078,In_1130,In_435);
nor U1079 (N_1079,In_1077,In_1145);
nor U1080 (N_1080,In_1532,In_680);
nand U1081 (N_1081,In_1432,In_740);
and U1082 (N_1082,In_1274,In_458);
nor U1083 (N_1083,In_1083,In_334);
nor U1084 (N_1084,In_409,In_637);
nor U1085 (N_1085,In_77,In_902);
nor U1086 (N_1086,In_260,In_1772);
and U1087 (N_1087,In_713,In_564);
nor U1088 (N_1088,In_1970,In_1285);
or U1089 (N_1089,In_962,In_348);
nor U1090 (N_1090,In_1225,In_467);
nor U1091 (N_1091,In_1130,In_193);
and U1092 (N_1092,In_54,In_147);
or U1093 (N_1093,In_1254,In_1022);
nor U1094 (N_1094,In_1980,In_419);
xor U1095 (N_1095,In_1999,In_1634);
and U1096 (N_1096,In_1424,In_1445);
or U1097 (N_1097,In_583,In_616);
and U1098 (N_1098,In_1332,In_985);
xnor U1099 (N_1099,In_1610,In_728);
and U1100 (N_1100,In_13,In_1308);
xor U1101 (N_1101,In_386,In_792);
nor U1102 (N_1102,In_1237,In_1827);
nand U1103 (N_1103,In_1896,In_587);
xnor U1104 (N_1104,In_1163,In_466);
and U1105 (N_1105,In_873,In_389);
nor U1106 (N_1106,In_1009,In_842);
and U1107 (N_1107,In_395,In_200);
and U1108 (N_1108,In_1251,In_639);
or U1109 (N_1109,In_281,In_1493);
or U1110 (N_1110,In_1691,In_815);
nand U1111 (N_1111,In_1390,In_1336);
or U1112 (N_1112,In_894,In_1332);
or U1113 (N_1113,In_1120,In_988);
nor U1114 (N_1114,In_1517,In_714);
nand U1115 (N_1115,In_1631,In_1239);
and U1116 (N_1116,In_1092,In_1041);
and U1117 (N_1117,In_1597,In_1578);
nor U1118 (N_1118,In_191,In_216);
nand U1119 (N_1119,In_1803,In_1646);
nor U1120 (N_1120,In_1715,In_1119);
nor U1121 (N_1121,In_1956,In_1898);
and U1122 (N_1122,In_212,In_1261);
and U1123 (N_1123,In_152,In_485);
nand U1124 (N_1124,In_1525,In_1363);
nand U1125 (N_1125,In_1492,In_162);
nor U1126 (N_1126,In_1956,In_761);
or U1127 (N_1127,In_1716,In_1778);
nand U1128 (N_1128,In_1782,In_1830);
and U1129 (N_1129,In_1060,In_362);
xnor U1130 (N_1130,In_569,In_990);
and U1131 (N_1131,In_1853,In_992);
xor U1132 (N_1132,In_1597,In_1331);
or U1133 (N_1133,In_1478,In_1718);
and U1134 (N_1134,In_1007,In_245);
and U1135 (N_1135,In_523,In_594);
and U1136 (N_1136,In_1376,In_92);
nor U1137 (N_1137,In_69,In_670);
and U1138 (N_1138,In_985,In_863);
nand U1139 (N_1139,In_1746,In_182);
nand U1140 (N_1140,In_558,In_1855);
nand U1141 (N_1141,In_805,In_117);
and U1142 (N_1142,In_1537,In_977);
nor U1143 (N_1143,In_1192,In_448);
nand U1144 (N_1144,In_395,In_1465);
nand U1145 (N_1145,In_1529,In_589);
nand U1146 (N_1146,In_171,In_1867);
or U1147 (N_1147,In_322,In_1469);
and U1148 (N_1148,In_733,In_886);
and U1149 (N_1149,In_932,In_195);
nand U1150 (N_1150,In_1070,In_1411);
and U1151 (N_1151,In_340,In_489);
and U1152 (N_1152,In_1510,In_1930);
nand U1153 (N_1153,In_1799,In_1122);
nor U1154 (N_1154,In_697,In_1836);
nand U1155 (N_1155,In_1400,In_975);
nor U1156 (N_1156,In_327,In_403);
or U1157 (N_1157,In_555,In_1530);
xnor U1158 (N_1158,In_1355,In_1646);
nand U1159 (N_1159,In_78,In_336);
nand U1160 (N_1160,In_1796,In_1727);
xnor U1161 (N_1161,In_900,In_382);
and U1162 (N_1162,In_1781,In_174);
and U1163 (N_1163,In_512,In_1657);
and U1164 (N_1164,In_142,In_124);
or U1165 (N_1165,In_722,In_29);
nand U1166 (N_1166,In_1786,In_554);
and U1167 (N_1167,In_1270,In_226);
and U1168 (N_1168,In_984,In_244);
or U1169 (N_1169,In_1331,In_1928);
nand U1170 (N_1170,In_526,In_1455);
nor U1171 (N_1171,In_538,In_1016);
nand U1172 (N_1172,In_1535,In_593);
or U1173 (N_1173,In_1,In_1149);
and U1174 (N_1174,In_1440,In_1108);
nor U1175 (N_1175,In_1919,In_396);
nor U1176 (N_1176,In_1267,In_1716);
and U1177 (N_1177,In_1562,In_1814);
or U1178 (N_1178,In_626,In_68);
and U1179 (N_1179,In_1160,In_492);
xor U1180 (N_1180,In_304,In_1829);
or U1181 (N_1181,In_1157,In_1231);
nor U1182 (N_1182,In_829,In_1868);
nand U1183 (N_1183,In_515,In_1178);
or U1184 (N_1184,In_677,In_62);
or U1185 (N_1185,In_404,In_1134);
xnor U1186 (N_1186,In_1301,In_696);
and U1187 (N_1187,In_1633,In_805);
or U1188 (N_1188,In_262,In_224);
and U1189 (N_1189,In_580,In_911);
or U1190 (N_1190,In_1741,In_1184);
or U1191 (N_1191,In_1893,In_37);
or U1192 (N_1192,In_1606,In_491);
xor U1193 (N_1193,In_1304,In_100);
nand U1194 (N_1194,In_0,In_624);
or U1195 (N_1195,In_416,In_69);
nand U1196 (N_1196,In_293,In_1414);
and U1197 (N_1197,In_654,In_1785);
nor U1198 (N_1198,In_244,In_1917);
nor U1199 (N_1199,In_1547,In_20);
or U1200 (N_1200,In_1647,In_1906);
nor U1201 (N_1201,In_1149,In_301);
or U1202 (N_1202,In_944,In_782);
and U1203 (N_1203,In_1033,In_1779);
and U1204 (N_1204,In_1681,In_255);
nand U1205 (N_1205,In_195,In_215);
nor U1206 (N_1206,In_1727,In_447);
or U1207 (N_1207,In_192,In_730);
xor U1208 (N_1208,In_1406,In_1747);
and U1209 (N_1209,In_362,In_634);
and U1210 (N_1210,In_1416,In_721);
nand U1211 (N_1211,In_1952,In_1162);
and U1212 (N_1212,In_1636,In_1987);
nor U1213 (N_1213,In_471,In_376);
or U1214 (N_1214,In_1646,In_1075);
and U1215 (N_1215,In_211,In_113);
nor U1216 (N_1216,In_1587,In_711);
xor U1217 (N_1217,In_222,In_1566);
and U1218 (N_1218,In_440,In_56);
xnor U1219 (N_1219,In_710,In_1808);
or U1220 (N_1220,In_744,In_1926);
nor U1221 (N_1221,In_1470,In_122);
xnor U1222 (N_1222,In_1394,In_1768);
or U1223 (N_1223,In_257,In_1166);
and U1224 (N_1224,In_1973,In_992);
nor U1225 (N_1225,In_400,In_1214);
or U1226 (N_1226,In_1806,In_1433);
nor U1227 (N_1227,In_1717,In_1012);
nor U1228 (N_1228,In_48,In_313);
xor U1229 (N_1229,In_1687,In_212);
or U1230 (N_1230,In_307,In_339);
and U1231 (N_1231,In_1477,In_173);
or U1232 (N_1232,In_1916,In_728);
and U1233 (N_1233,In_1815,In_895);
xnor U1234 (N_1234,In_1236,In_1258);
and U1235 (N_1235,In_1921,In_685);
nor U1236 (N_1236,In_1903,In_389);
and U1237 (N_1237,In_338,In_1382);
nor U1238 (N_1238,In_857,In_23);
and U1239 (N_1239,In_1338,In_1719);
and U1240 (N_1240,In_853,In_202);
nor U1241 (N_1241,In_1485,In_453);
nand U1242 (N_1242,In_1407,In_1196);
and U1243 (N_1243,In_1224,In_1378);
or U1244 (N_1244,In_1048,In_936);
or U1245 (N_1245,In_1083,In_712);
nand U1246 (N_1246,In_803,In_1302);
nand U1247 (N_1247,In_53,In_1840);
or U1248 (N_1248,In_1142,In_1966);
nor U1249 (N_1249,In_5,In_1922);
and U1250 (N_1250,In_965,In_1589);
or U1251 (N_1251,In_1449,In_1003);
nand U1252 (N_1252,In_897,In_1773);
and U1253 (N_1253,In_937,In_1717);
xor U1254 (N_1254,In_898,In_659);
nor U1255 (N_1255,In_1436,In_317);
or U1256 (N_1256,In_289,In_602);
nor U1257 (N_1257,In_1637,In_533);
nand U1258 (N_1258,In_1129,In_536);
and U1259 (N_1259,In_263,In_1792);
nor U1260 (N_1260,In_1744,In_883);
nor U1261 (N_1261,In_108,In_60);
or U1262 (N_1262,In_276,In_543);
nor U1263 (N_1263,In_1336,In_131);
or U1264 (N_1264,In_1809,In_1613);
nor U1265 (N_1265,In_1227,In_655);
and U1266 (N_1266,In_1091,In_1843);
nor U1267 (N_1267,In_1539,In_773);
xnor U1268 (N_1268,In_1920,In_947);
nor U1269 (N_1269,In_1391,In_1726);
nand U1270 (N_1270,In_1987,In_257);
xor U1271 (N_1271,In_548,In_657);
nand U1272 (N_1272,In_1912,In_701);
nand U1273 (N_1273,In_1965,In_1177);
xor U1274 (N_1274,In_435,In_1230);
nand U1275 (N_1275,In_1293,In_1002);
nand U1276 (N_1276,In_1933,In_144);
and U1277 (N_1277,In_30,In_494);
and U1278 (N_1278,In_539,In_1087);
nor U1279 (N_1279,In_299,In_1062);
and U1280 (N_1280,In_1627,In_108);
or U1281 (N_1281,In_1786,In_1108);
nor U1282 (N_1282,In_1474,In_1495);
nor U1283 (N_1283,In_113,In_1103);
nor U1284 (N_1284,In_617,In_996);
and U1285 (N_1285,In_540,In_1456);
nand U1286 (N_1286,In_1007,In_742);
nand U1287 (N_1287,In_604,In_343);
and U1288 (N_1288,In_238,In_1663);
or U1289 (N_1289,In_1147,In_53);
nor U1290 (N_1290,In_542,In_735);
nand U1291 (N_1291,In_1926,In_341);
or U1292 (N_1292,In_736,In_959);
nand U1293 (N_1293,In_1924,In_184);
xnor U1294 (N_1294,In_864,In_122);
nand U1295 (N_1295,In_1258,In_1499);
nand U1296 (N_1296,In_1075,In_391);
or U1297 (N_1297,In_1539,In_253);
nor U1298 (N_1298,In_1694,In_1356);
nand U1299 (N_1299,In_1717,In_1851);
and U1300 (N_1300,In_1356,In_1099);
nand U1301 (N_1301,In_1912,In_1956);
and U1302 (N_1302,In_1673,In_1566);
xnor U1303 (N_1303,In_1879,In_1596);
nor U1304 (N_1304,In_960,In_553);
nor U1305 (N_1305,In_163,In_703);
nand U1306 (N_1306,In_43,In_1943);
and U1307 (N_1307,In_589,In_313);
nor U1308 (N_1308,In_960,In_819);
xnor U1309 (N_1309,In_1655,In_224);
xnor U1310 (N_1310,In_1367,In_1375);
or U1311 (N_1311,In_1697,In_1580);
and U1312 (N_1312,In_1482,In_221);
nor U1313 (N_1313,In_1896,In_1215);
or U1314 (N_1314,In_1740,In_1710);
nor U1315 (N_1315,In_1612,In_1157);
nand U1316 (N_1316,In_1341,In_445);
or U1317 (N_1317,In_812,In_1432);
nand U1318 (N_1318,In_665,In_401);
xor U1319 (N_1319,In_343,In_1916);
nor U1320 (N_1320,In_512,In_570);
or U1321 (N_1321,In_1003,In_595);
nand U1322 (N_1322,In_1940,In_1892);
nand U1323 (N_1323,In_857,In_657);
and U1324 (N_1324,In_1426,In_515);
and U1325 (N_1325,In_1085,In_1592);
and U1326 (N_1326,In_1324,In_66);
nor U1327 (N_1327,In_1788,In_1930);
and U1328 (N_1328,In_179,In_1617);
and U1329 (N_1329,In_1548,In_1975);
or U1330 (N_1330,In_1939,In_1865);
xnor U1331 (N_1331,In_1,In_1856);
and U1332 (N_1332,In_786,In_654);
or U1333 (N_1333,In_1565,In_104);
nor U1334 (N_1334,In_1871,In_1379);
or U1335 (N_1335,In_1280,In_599);
and U1336 (N_1336,In_710,In_1458);
xnor U1337 (N_1337,In_110,In_1476);
and U1338 (N_1338,In_838,In_1151);
and U1339 (N_1339,In_1919,In_367);
nor U1340 (N_1340,In_288,In_430);
nand U1341 (N_1341,In_201,In_1008);
or U1342 (N_1342,In_919,In_1577);
and U1343 (N_1343,In_1629,In_1571);
xnor U1344 (N_1344,In_172,In_1661);
or U1345 (N_1345,In_55,In_521);
nor U1346 (N_1346,In_1538,In_1836);
and U1347 (N_1347,In_27,In_1518);
nor U1348 (N_1348,In_1864,In_1322);
and U1349 (N_1349,In_560,In_483);
xnor U1350 (N_1350,In_493,In_1624);
nand U1351 (N_1351,In_1042,In_79);
and U1352 (N_1352,In_1142,In_1371);
or U1353 (N_1353,In_1777,In_830);
or U1354 (N_1354,In_1669,In_1497);
nand U1355 (N_1355,In_48,In_1258);
xnor U1356 (N_1356,In_1823,In_717);
or U1357 (N_1357,In_1567,In_947);
nand U1358 (N_1358,In_213,In_1575);
nor U1359 (N_1359,In_1928,In_1821);
nand U1360 (N_1360,In_658,In_1317);
or U1361 (N_1361,In_1828,In_1263);
nor U1362 (N_1362,In_1284,In_51);
nand U1363 (N_1363,In_1391,In_1062);
and U1364 (N_1364,In_558,In_1684);
or U1365 (N_1365,In_1119,In_1853);
nor U1366 (N_1366,In_1760,In_933);
nor U1367 (N_1367,In_1220,In_1110);
xor U1368 (N_1368,In_803,In_1792);
and U1369 (N_1369,In_1022,In_1688);
xor U1370 (N_1370,In_1440,In_58);
nand U1371 (N_1371,In_922,In_297);
and U1372 (N_1372,In_294,In_1920);
nor U1373 (N_1373,In_1600,In_1538);
nand U1374 (N_1374,In_927,In_149);
nor U1375 (N_1375,In_1853,In_637);
nor U1376 (N_1376,In_1642,In_1814);
xnor U1377 (N_1377,In_484,In_1481);
xor U1378 (N_1378,In_833,In_1706);
and U1379 (N_1379,In_1218,In_1180);
nor U1380 (N_1380,In_1134,In_365);
or U1381 (N_1381,In_174,In_315);
or U1382 (N_1382,In_322,In_1621);
nor U1383 (N_1383,In_1812,In_55);
and U1384 (N_1384,In_1235,In_1138);
or U1385 (N_1385,In_192,In_1393);
and U1386 (N_1386,In_746,In_1018);
nand U1387 (N_1387,In_1188,In_258);
nand U1388 (N_1388,In_1293,In_609);
xnor U1389 (N_1389,In_1905,In_989);
nor U1390 (N_1390,In_1548,In_1978);
nor U1391 (N_1391,In_312,In_1345);
xnor U1392 (N_1392,In_846,In_1663);
nand U1393 (N_1393,In_1401,In_859);
and U1394 (N_1394,In_1737,In_1069);
xnor U1395 (N_1395,In_1798,In_770);
or U1396 (N_1396,In_1189,In_1458);
nor U1397 (N_1397,In_1593,In_1067);
xor U1398 (N_1398,In_1879,In_77);
nand U1399 (N_1399,In_471,In_1552);
nand U1400 (N_1400,In_1983,In_1997);
and U1401 (N_1401,In_646,In_740);
xor U1402 (N_1402,In_633,In_1350);
nor U1403 (N_1403,In_836,In_1005);
nor U1404 (N_1404,In_115,In_1802);
and U1405 (N_1405,In_1268,In_1930);
and U1406 (N_1406,In_1976,In_907);
nand U1407 (N_1407,In_732,In_1274);
nor U1408 (N_1408,In_772,In_1692);
nor U1409 (N_1409,In_426,In_1909);
xor U1410 (N_1410,In_775,In_1341);
nor U1411 (N_1411,In_1341,In_65);
nand U1412 (N_1412,In_1167,In_758);
and U1413 (N_1413,In_1188,In_502);
nand U1414 (N_1414,In_634,In_264);
nor U1415 (N_1415,In_2,In_80);
or U1416 (N_1416,In_1673,In_1648);
nand U1417 (N_1417,In_291,In_516);
or U1418 (N_1418,In_1980,In_788);
nor U1419 (N_1419,In_879,In_1320);
nor U1420 (N_1420,In_1983,In_262);
xnor U1421 (N_1421,In_610,In_399);
and U1422 (N_1422,In_1970,In_390);
nor U1423 (N_1423,In_1017,In_916);
and U1424 (N_1424,In_1126,In_1375);
xnor U1425 (N_1425,In_929,In_368);
nor U1426 (N_1426,In_1194,In_271);
nor U1427 (N_1427,In_1762,In_1);
nand U1428 (N_1428,In_248,In_1826);
nor U1429 (N_1429,In_1008,In_1389);
nand U1430 (N_1430,In_349,In_499);
or U1431 (N_1431,In_1622,In_232);
or U1432 (N_1432,In_1964,In_1835);
and U1433 (N_1433,In_1204,In_1389);
and U1434 (N_1434,In_1182,In_1609);
nand U1435 (N_1435,In_744,In_42);
xor U1436 (N_1436,In_378,In_856);
nand U1437 (N_1437,In_1960,In_1863);
and U1438 (N_1438,In_1726,In_858);
or U1439 (N_1439,In_680,In_649);
nor U1440 (N_1440,In_719,In_1083);
nor U1441 (N_1441,In_735,In_1554);
nor U1442 (N_1442,In_400,In_539);
nor U1443 (N_1443,In_1105,In_40);
or U1444 (N_1444,In_1064,In_234);
and U1445 (N_1445,In_1802,In_1237);
nor U1446 (N_1446,In_617,In_243);
nand U1447 (N_1447,In_1720,In_266);
nor U1448 (N_1448,In_1620,In_1235);
and U1449 (N_1449,In_288,In_1222);
xnor U1450 (N_1450,In_794,In_1533);
nor U1451 (N_1451,In_1497,In_1338);
and U1452 (N_1452,In_1766,In_1544);
xnor U1453 (N_1453,In_1268,In_1004);
and U1454 (N_1454,In_365,In_1313);
xnor U1455 (N_1455,In_1049,In_1137);
nor U1456 (N_1456,In_347,In_1788);
nand U1457 (N_1457,In_19,In_1485);
or U1458 (N_1458,In_1757,In_1772);
nor U1459 (N_1459,In_1049,In_848);
and U1460 (N_1460,In_1536,In_1280);
and U1461 (N_1461,In_201,In_1541);
or U1462 (N_1462,In_98,In_1943);
nand U1463 (N_1463,In_189,In_1525);
or U1464 (N_1464,In_1746,In_145);
or U1465 (N_1465,In_1465,In_603);
and U1466 (N_1466,In_730,In_158);
nand U1467 (N_1467,In_108,In_404);
or U1468 (N_1468,In_1548,In_1821);
nand U1469 (N_1469,In_538,In_152);
nor U1470 (N_1470,In_1298,In_1433);
xnor U1471 (N_1471,In_1896,In_18);
or U1472 (N_1472,In_213,In_189);
nor U1473 (N_1473,In_905,In_1031);
xor U1474 (N_1474,In_1746,In_474);
nand U1475 (N_1475,In_1819,In_172);
and U1476 (N_1476,In_1366,In_758);
or U1477 (N_1477,In_120,In_547);
and U1478 (N_1478,In_261,In_1059);
nor U1479 (N_1479,In_323,In_653);
xor U1480 (N_1480,In_414,In_271);
nand U1481 (N_1481,In_1816,In_521);
nor U1482 (N_1482,In_887,In_632);
or U1483 (N_1483,In_393,In_1781);
or U1484 (N_1484,In_1642,In_1840);
xor U1485 (N_1485,In_319,In_51);
or U1486 (N_1486,In_1364,In_1904);
or U1487 (N_1487,In_1939,In_1680);
nor U1488 (N_1488,In_1711,In_1346);
or U1489 (N_1489,In_64,In_681);
nor U1490 (N_1490,In_1074,In_1445);
and U1491 (N_1491,In_84,In_1225);
nor U1492 (N_1492,In_754,In_1503);
and U1493 (N_1493,In_1688,In_1);
nor U1494 (N_1494,In_1004,In_30);
xor U1495 (N_1495,In_333,In_1915);
and U1496 (N_1496,In_787,In_615);
and U1497 (N_1497,In_742,In_46);
nor U1498 (N_1498,In_118,In_144);
nor U1499 (N_1499,In_981,In_605);
xor U1500 (N_1500,In_477,In_695);
nand U1501 (N_1501,In_1683,In_887);
and U1502 (N_1502,In_1191,In_518);
and U1503 (N_1503,In_1437,In_1091);
nor U1504 (N_1504,In_1342,In_1456);
xor U1505 (N_1505,In_387,In_1388);
and U1506 (N_1506,In_1986,In_1292);
and U1507 (N_1507,In_1871,In_1233);
nand U1508 (N_1508,In_98,In_1947);
xnor U1509 (N_1509,In_430,In_1144);
nand U1510 (N_1510,In_463,In_1536);
nand U1511 (N_1511,In_92,In_1004);
and U1512 (N_1512,In_639,In_368);
nand U1513 (N_1513,In_1944,In_1557);
or U1514 (N_1514,In_1093,In_1942);
nor U1515 (N_1515,In_67,In_827);
nand U1516 (N_1516,In_98,In_740);
or U1517 (N_1517,In_101,In_657);
and U1518 (N_1518,In_1808,In_456);
nand U1519 (N_1519,In_104,In_384);
nand U1520 (N_1520,In_1739,In_687);
or U1521 (N_1521,In_1398,In_156);
and U1522 (N_1522,In_1998,In_1141);
or U1523 (N_1523,In_137,In_1697);
or U1524 (N_1524,In_1587,In_755);
xnor U1525 (N_1525,In_509,In_1903);
nand U1526 (N_1526,In_1038,In_1307);
and U1527 (N_1527,In_313,In_202);
or U1528 (N_1528,In_1218,In_1797);
or U1529 (N_1529,In_1826,In_524);
or U1530 (N_1530,In_350,In_968);
or U1531 (N_1531,In_1643,In_854);
and U1532 (N_1532,In_334,In_1);
and U1533 (N_1533,In_433,In_26);
nand U1534 (N_1534,In_488,In_1168);
nor U1535 (N_1535,In_1514,In_1608);
nand U1536 (N_1536,In_515,In_402);
or U1537 (N_1537,In_1859,In_333);
and U1538 (N_1538,In_1225,In_800);
or U1539 (N_1539,In_79,In_195);
and U1540 (N_1540,In_77,In_1955);
nor U1541 (N_1541,In_1436,In_487);
nand U1542 (N_1542,In_964,In_379);
nand U1543 (N_1543,In_1520,In_603);
nand U1544 (N_1544,In_1707,In_1334);
nor U1545 (N_1545,In_732,In_1109);
and U1546 (N_1546,In_991,In_947);
nand U1547 (N_1547,In_364,In_245);
or U1548 (N_1548,In_1933,In_1511);
and U1549 (N_1549,In_559,In_1187);
and U1550 (N_1550,In_457,In_1809);
and U1551 (N_1551,In_1273,In_1250);
and U1552 (N_1552,In_1518,In_786);
nand U1553 (N_1553,In_1436,In_980);
nor U1554 (N_1554,In_70,In_717);
nor U1555 (N_1555,In_1502,In_1917);
nand U1556 (N_1556,In_436,In_1847);
and U1557 (N_1557,In_942,In_1506);
nor U1558 (N_1558,In_1151,In_1298);
xor U1559 (N_1559,In_978,In_1221);
or U1560 (N_1560,In_1668,In_1165);
nor U1561 (N_1561,In_1843,In_534);
xnor U1562 (N_1562,In_1477,In_1736);
or U1563 (N_1563,In_905,In_706);
and U1564 (N_1564,In_1119,In_252);
and U1565 (N_1565,In_1645,In_752);
nand U1566 (N_1566,In_352,In_702);
nor U1567 (N_1567,In_1561,In_298);
and U1568 (N_1568,In_1308,In_736);
xnor U1569 (N_1569,In_1309,In_1901);
nor U1570 (N_1570,In_1923,In_1260);
nand U1571 (N_1571,In_429,In_1266);
nand U1572 (N_1572,In_1436,In_70);
xnor U1573 (N_1573,In_67,In_184);
and U1574 (N_1574,In_448,In_576);
nand U1575 (N_1575,In_646,In_1954);
and U1576 (N_1576,In_229,In_1748);
or U1577 (N_1577,In_853,In_118);
or U1578 (N_1578,In_1413,In_304);
xnor U1579 (N_1579,In_37,In_1285);
nor U1580 (N_1580,In_28,In_609);
nor U1581 (N_1581,In_916,In_412);
or U1582 (N_1582,In_861,In_1352);
and U1583 (N_1583,In_906,In_853);
and U1584 (N_1584,In_1861,In_1842);
or U1585 (N_1585,In_1855,In_1423);
xor U1586 (N_1586,In_1721,In_296);
xnor U1587 (N_1587,In_1963,In_54);
or U1588 (N_1588,In_867,In_618);
nand U1589 (N_1589,In_1039,In_231);
or U1590 (N_1590,In_914,In_1550);
nand U1591 (N_1591,In_1940,In_1833);
or U1592 (N_1592,In_1465,In_280);
nand U1593 (N_1593,In_1025,In_1057);
and U1594 (N_1594,In_1212,In_444);
nand U1595 (N_1595,In_924,In_88);
nand U1596 (N_1596,In_40,In_1339);
or U1597 (N_1597,In_1834,In_999);
xor U1598 (N_1598,In_238,In_544);
xor U1599 (N_1599,In_1886,In_1759);
nand U1600 (N_1600,In_667,In_980);
nor U1601 (N_1601,In_486,In_366);
nand U1602 (N_1602,In_1409,In_1798);
nor U1603 (N_1603,In_964,In_426);
nor U1604 (N_1604,In_1305,In_1693);
or U1605 (N_1605,In_1029,In_1944);
nand U1606 (N_1606,In_1774,In_472);
xnor U1607 (N_1607,In_1628,In_82);
or U1608 (N_1608,In_792,In_1718);
and U1609 (N_1609,In_516,In_966);
or U1610 (N_1610,In_209,In_1419);
and U1611 (N_1611,In_952,In_140);
or U1612 (N_1612,In_1106,In_1522);
and U1613 (N_1613,In_80,In_3);
nand U1614 (N_1614,In_759,In_1958);
nor U1615 (N_1615,In_1028,In_711);
and U1616 (N_1616,In_217,In_932);
and U1617 (N_1617,In_1693,In_1629);
or U1618 (N_1618,In_197,In_1940);
nor U1619 (N_1619,In_149,In_1803);
and U1620 (N_1620,In_1577,In_647);
nor U1621 (N_1621,In_543,In_1218);
xor U1622 (N_1622,In_317,In_179);
nand U1623 (N_1623,In_820,In_1657);
and U1624 (N_1624,In_1360,In_1363);
nand U1625 (N_1625,In_1066,In_661);
nor U1626 (N_1626,In_1105,In_881);
nor U1627 (N_1627,In_972,In_535);
and U1628 (N_1628,In_229,In_1272);
nor U1629 (N_1629,In_516,In_760);
nand U1630 (N_1630,In_74,In_1225);
nor U1631 (N_1631,In_1950,In_82);
nand U1632 (N_1632,In_1829,In_1205);
nor U1633 (N_1633,In_1876,In_962);
or U1634 (N_1634,In_697,In_1150);
nor U1635 (N_1635,In_1924,In_132);
and U1636 (N_1636,In_626,In_1301);
nor U1637 (N_1637,In_434,In_809);
nor U1638 (N_1638,In_1350,In_133);
nor U1639 (N_1639,In_281,In_1428);
xor U1640 (N_1640,In_1261,In_256);
or U1641 (N_1641,In_309,In_1645);
nor U1642 (N_1642,In_1813,In_1285);
or U1643 (N_1643,In_1280,In_978);
and U1644 (N_1644,In_946,In_962);
nand U1645 (N_1645,In_1916,In_786);
nand U1646 (N_1646,In_933,In_1831);
nand U1647 (N_1647,In_421,In_1596);
and U1648 (N_1648,In_659,In_1269);
or U1649 (N_1649,In_713,In_1379);
nand U1650 (N_1650,In_1825,In_1339);
nor U1651 (N_1651,In_1545,In_713);
nor U1652 (N_1652,In_756,In_1591);
or U1653 (N_1653,In_149,In_1699);
or U1654 (N_1654,In_487,In_610);
or U1655 (N_1655,In_387,In_1350);
nor U1656 (N_1656,In_720,In_1826);
nand U1657 (N_1657,In_863,In_1592);
xnor U1658 (N_1658,In_747,In_420);
or U1659 (N_1659,In_1424,In_7);
and U1660 (N_1660,In_1015,In_1441);
nor U1661 (N_1661,In_482,In_1339);
or U1662 (N_1662,In_1131,In_603);
or U1663 (N_1663,In_324,In_1650);
nor U1664 (N_1664,In_881,In_507);
nand U1665 (N_1665,In_1801,In_686);
nor U1666 (N_1666,In_404,In_818);
and U1667 (N_1667,In_966,In_1602);
nor U1668 (N_1668,In_59,In_169);
and U1669 (N_1669,In_538,In_1775);
and U1670 (N_1670,In_1791,In_1236);
nand U1671 (N_1671,In_1921,In_1429);
nor U1672 (N_1672,In_1200,In_1198);
nand U1673 (N_1673,In_589,In_1329);
and U1674 (N_1674,In_1420,In_395);
nand U1675 (N_1675,In_656,In_423);
nor U1676 (N_1676,In_990,In_1695);
and U1677 (N_1677,In_632,In_498);
and U1678 (N_1678,In_777,In_440);
nor U1679 (N_1679,In_423,In_903);
nand U1680 (N_1680,In_941,In_1952);
nand U1681 (N_1681,In_1558,In_1992);
nor U1682 (N_1682,In_1860,In_510);
and U1683 (N_1683,In_914,In_169);
xor U1684 (N_1684,In_1512,In_496);
and U1685 (N_1685,In_665,In_766);
nand U1686 (N_1686,In_442,In_420);
and U1687 (N_1687,In_1368,In_197);
or U1688 (N_1688,In_1582,In_570);
nand U1689 (N_1689,In_1781,In_1153);
and U1690 (N_1690,In_307,In_1725);
and U1691 (N_1691,In_1224,In_1147);
nor U1692 (N_1692,In_1062,In_591);
xor U1693 (N_1693,In_161,In_523);
and U1694 (N_1694,In_94,In_524);
and U1695 (N_1695,In_471,In_1058);
nor U1696 (N_1696,In_1127,In_957);
nand U1697 (N_1697,In_1057,In_228);
or U1698 (N_1698,In_1939,In_1112);
or U1699 (N_1699,In_1037,In_1703);
xnor U1700 (N_1700,In_42,In_1322);
or U1701 (N_1701,In_1013,In_869);
nor U1702 (N_1702,In_952,In_1748);
nand U1703 (N_1703,In_1209,In_1050);
xnor U1704 (N_1704,In_409,In_535);
nand U1705 (N_1705,In_1783,In_1100);
nand U1706 (N_1706,In_1911,In_1293);
xnor U1707 (N_1707,In_1384,In_1073);
nand U1708 (N_1708,In_689,In_834);
nand U1709 (N_1709,In_1716,In_1916);
nor U1710 (N_1710,In_999,In_1727);
or U1711 (N_1711,In_315,In_785);
nand U1712 (N_1712,In_1399,In_1448);
nand U1713 (N_1713,In_1103,In_1593);
nand U1714 (N_1714,In_1800,In_429);
or U1715 (N_1715,In_702,In_798);
nor U1716 (N_1716,In_1906,In_1517);
and U1717 (N_1717,In_678,In_1559);
nand U1718 (N_1718,In_947,In_275);
and U1719 (N_1719,In_1779,In_1843);
nand U1720 (N_1720,In_1982,In_1892);
xor U1721 (N_1721,In_885,In_1868);
or U1722 (N_1722,In_1304,In_1210);
nand U1723 (N_1723,In_1450,In_235);
xnor U1724 (N_1724,In_1422,In_1394);
nor U1725 (N_1725,In_1618,In_663);
xnor U1726 (N_1726,In_1987,In_1543);
or U1727 (N_1727,In_179,In_755);
nor U1728 (N_1728,In_1043,In_1334);
and U1729 (N_1729,In_1276,In_997);
and U1730 (N_1730,In_1555,In_14);
or U1731 (N_1731,In_689,In_1832);
or U1732 (N_1732,In_1223,In_477);
nand U1733 (N_1733,In_776,In_1060);
or U1734 (N_1734,In_559,In_1404);
nor U1735 (N_1735,In_312,In_784);
nor U1736 (N_1736,In_1440,In_1188);
nor U1737 (N_1737,In_1163,In_46);
nand U1738 (N_1738,In_1052,In_1995);
nor U1739 (N_1739,In_519,In_1907);
and U1740 (N_1740,In_206,In_601);
and U1741 (N_1741,In_1442,In_661);
nor U1742 (N_1742,In_1681,In_648);
and U1743 (N_1743,In_1440,In_1748);
xnor U1744 (N_1744,In_62,In_461);
nor U1745 (N_1745,In_969,In_1366);
nand U1746 (N_1746,In_225,In_584);
nor U1747 (N_1747,In_549,In_922);
xnor U1748 (N_1748,In_204,In_16);
nand U1749 (N_1749,In_1384,In_1688);
or U1750 (N_1750,In_1328,In_1636);
nor U1751 (N_1751,In_1604,In_26);
nor U1752 (N_1752,In_317,In_164);
and U1753 (N_1753,In_562,In_862);
nor U1754 (N_1754,In_399,In_214);
or U1755 (N_1755,In_780,In_560);
nand U1756 (N_1756,In_1633,In_11);
nor U1757 (N_1757,In_1603,In_1495);
nor U1758 (N_1758,In_1376,In_1432);
xor U1759 (N_1759,In_31,In_1841);
or U1760 (N_1760,In_554,In_560);
or U1761 (N_1761,In_1675,In_1032);
nand U1762 (N_1762,In_712,In_64);
nor U1763 (N_1763,In_1471,In_112);
or U1764 (N_1764,In_95,In_1928);
and U1765 (N_1765,In_19,In_539);
or U1766 (N_1766,In_361,In_1205);
or U1767 (N_1767,In_1305,In_702);
or U1768 (N_1768,In_277,In_163);
nor U1769 (N_1769,In_125,In_22);
nand U1770 (N_1770,In_515,In_1832);
or U1771 (N_1771,In_753,In_413);
or U1772 (N_1772,In_1267,In_1058);
nor U1773 (N_1773,In_672,In_1471);
xor U1774 (N_1774,In_64,In_443);
nor U1775 (N_1775,In_165,In_1637);
and U1776 (N_1776,In_1597,In_1294);
nor U1777 (N_1777,In_1582,In_1510);
and U1778 (N_1778,In_1037,In_364);
nand U1779 (N_1779,In_289,In_74);
or U1780 (N_1780,In_711,In_126);
or U1781 (N_1781,In_1902,In_460);
nor U1782 (N_1782,In_965,In_757);
or U1783 (N_1783,In_1886,In_1604);
or U1784 (N_1784,In_1482,In_1198);
and U1785 (N_1785,In_1436,In_1741);
or U1786 (N_1786,In_985,In_1699);
and U1787 (N_1787,In_1298,In_1866);
nor U1788 (N_1788,In_770,In_933);
or U1789 (N_1789,In_1300,In_933);
or U1790 (N_1790,In_1486,In_896);
and U1791 (N_1791,In_306,In_671);
xnor U1792 (N_1792,In_1735,In_654);
or U1793 (N_1793,In_1367,In_967);
xor U1794 (N_1794,In_1010,In_1557);
xnor U1795 (N_1795,In_1176,In_595);
nor U1796 (N_1796,In_1455,In_1626);
nor U1797 (N_1797,In_434,In_23);
xor U1798 (N_1798,In_1943,In_1321);
nor U1799 (N_1799,In_115,In_1984);
nor U1800 (N_1800,In_695,In_497);
nand U1801 (N_1801,In_940,In_292);
or U1802 (N_1802,In_1015,In_438);
nor U1803 (N_1803,In_956,In_1944);
nor U1804 (N_1804,In_1388,In_392);
xor U1805 (N_1805,In_1233,In_815);
xnor U1806 (N_1806,In_1715,In_1149);
or U1807 (N_1807,In_485,In_444);
and U1808 (N_1808,In_1545,In_901);
nand U1809 (N_1809,In_324,In_1542);
and U1810 (N_1810,In_1568,In_1502);
nand U1811 (N_1811,In_497,In_372);
and U1812 (N_1812,In_5,In_1234);
and U1813 (N_1813,In_586,In_505);
nor U1814 (N_1814,In_1246,In_939);
nor U1815 (N_1815,In_1175,In_9);
xor U1816 (N_1816,In_963,In_1389);
nand U1817 (N_1817,In_1159,In_1792);
and U1818 (N_1818,In_494,In_608);
nor U1819 (N_1819,In_956,In_1986);
or U1820 (N_1820,In_23,In_758);
or U1821 (N_1821,In_362,In_336);
or U1822 (N_1822,In_1212,In_1545);
or U1823 (N_1823,In_1977,In_1346);
or U1824 (N_1824,In_1691,In_1844);
and U1825 (N_1825,In_744,In_313);
and U1826 (N_1826,In_620,In_787);
and U1827 (N_1827,In_357,In_1688);
or U1828 (N_1828,In_1182,In_705);
nand U1829 (N_1829,In_878,In_1305);
xnor U1830 (N_1830,In_974,In_678);
and U1831 (N_1831,In_1165,In_1999);
xnor U1832 (N_1832,In_426,In_673);
and U1833 (N_1833,In_1251,In_1509);
nand U1834 (N_1834,In_1301,In_1367);
and U1835 (N_1835,In_873,In_180);
and U1836 (N_1836,In_624,In_1111);
and U1837 (N_1837,In_851,In_638);
nor U1838 (N_1838,In_886,In_425);
and U1839 (N_1839,In_388,In_1547);
or U1840 (N_1840,In_765,In_1382);
or U1841 (N_1841,In_1607,In_190);
or U1842 (N_1842,In_508,In_132);
and U1843 (N_1843,In_379,In_963);
nor U1844 (N_1844,In_1232,In_1130);
nand U1845 (N_1845,In_1771,In_341);
xor U1846 (N_1846,In_1491,In_1043);
nor U1847 (N_1847,In_1657,In_1569);
or U1848 (N_1848,In_926,In_874);
or U1849 (N_1849,In_1864,In_990);
nor U1850 (N_1850,In_257,In_867);
nand U1851 (N_1851,In_1367,In_1328);
nand U1852 (N_1852,In_1836,In_6);
nor U1853 (N_1853,In_1326,In_980);
nand U1854 (N_1854,In_56,In_336);
or U1855 (N_1855,In_261,In_1929);
nor U1856 (N_1856,In_266,In_47);
or U1857 (N_1857,In_439,In_1221);
nor U1858 (N_1858,In_135,In_170);
nor U1859 (N_1859,In_1246,In_868);
nand U1860 (N_1860,In_888,In_1574);
nor U1861 (N_1861,In_325,In_864);
or U1862 (N_1862,In_1589,In_1288);
and U1863 (N_1863,In_1297,In_1548);
nand U1864 (N_1864,In_401,In_1257);
and U1865 (N_1865,In_1292,In_1456);
nand U1866 (N_1866,In_344,In_30);
xnor U1867 (N_1867,In_1743,In_722);
xnor U1868 (N_1868,In_891,In_931);
or U1869 (N_1869,In_1960,In_1266);
or U1870 (N_1870,In_420,In_510);
nor U1871 (N_1871,In_1044,In_161);
nor U1872 (N_1872,In_64,In_1817);
or U1873 (N_1873,In_1472,In_93);
or U1874 (N_1874,In_1381,In_1291);
nand U1875 (N_1875,In_675,In_424);
nor U1876 (N_1876,In_891,In_1973);
nor U1877 (N_1877,In_1077,In_69);
nor U1878 (N_1878,In_294,In_712);
nor U1879 (N_1879,In_45,In_1444);
xnor U1880 (N_1880,In_477,In_265);
or U1881 (N_1881,In_1748,In_745);
nand U1882 (N_1882,In_1334,In_1289);
and U1883 (N_1883,In_579,In_135);
nand U1884 (N_1884,In_1233,In_976);
and U1885 (N_1885,In_947,In_369);
nor U1886 (N_1886,In_732,In_1298);
and U1887 (N_1887,In_162,In_107);
nor U1888 (N_1888,In_1256,In_448);
nor U1889 (N_1889,In_843,In_1075);
nand U1890 (N_1890,In_1214,In_208);
and U1891 (N_1891,In_1614,In_115);
and U1892 (N_1892,In_447,In_454);
and U1893 (N_1893,In_580,In_1435);
xnor U1894 (N_1894,In_1412,In_1313);
nand U1895 (N_1895,In_1120,In_784);
nor U1896 (N_1896,In_927,In_1213);
nor U1897 (N_1897,In_66,In_1730);
nor U1898 (N_1898,In_915,In_1052);
or U1899 (N_1899,In_1994,In_1495);
or U1900 (N_1900,In_1546,In_1302);
nor U1901 (N_1901,In_1502,In_1643);
or U1902 (N_1902,In_438,In_1510);
nor U1903 (N_1903,In_858,In_1984);
nor U1904 (N_1904,In_1061,In_839);
nand U1905 (N_1905,In_557,In_1851);
and U1906 (N_1906,In_869,In_924);
nand U1907 (N_1907,In_1703,In_559);
nor U1908 (N_1908,In_781,In_1375);
nand U1909 (N_1909,In_706,In_1570);
nor U1910 (N_1910,In_1096,In_639);
nor U1911 (N_1911,In_588,In_1464);
nor U1912 (N_1912,In_979,In_1486);
xnor U1913 (N_1913,In_1073,In_1670);
nor U1914 (N_1914,In_1605,In_984);
and U1915 (N_1915,In_1655,In_575);
and U1916 (N_1916,In_1055,In_1298);
and U1917 (N_1917,In_706,In_1285);
nor U1918 (N_1918,In_1261,In_863);
and U1919 (N_1919,In_67,In_1313);
xor U1920 (N_1920,In_361,In_526);
or U1921 (N_1921,In_95,In_1014);
or U1922 (N_1922,In_1438,In_640);
and U1923 (N_1923,In_641,In_1159);
nand U1924 (N_1924,In_1680,In_1517);
and U1925 (N_1925,In_1145,In_1706);
nand U1926 (N_1926,In_1079,In_302);
or U1927 (N_1927,In_47,In_576);
nor U1928 (N_1928,In_1145,In_258);
nor U1929 (N_1929,In_202,In_574);
nor U1930 (N_1930,In_1755,In_818);
nor U1931 (N_1931,In_456,In_1920);
nor U1932 (N_1932,In_720,In_313);
nor U1933 (N_1933,In_1208,In_435);
or U1934 (N_1934,In_1463,In_326);
or U1935 (N_1935,In_772,In_1458);
and U1936 (N_1936,In_718,In_1127);
and U1937 (N_1937,In_1219,In_776);
and U1938 (N_1938,In_243,In_1451);
nor U1939 (N_1939,In_432,In_810);
nand U1940 (N_1940,In_1655,In_333);
and U1941 (N_1941,In_985,In_1524);
and U1942 (N_1942,In_1308,In_1982);
nand U1943 (N_1943,In_1062,In_164);
and U1944 (N_1944,In_412,In_58);
nor U1945 (N_1945,In_605,In_323);
and U1946 (N_1946,In_724,In_1819);
nand U1947 (N_1947,In_1738,In_1857);
nand U1948 (N_1948,In_1914,In_1642);
and U1949 (N_1949,In_527,In_45);
and U1950 (N_1950,In_943,In_1334);
nor U1951 (N_1951,In_726,In_584);
nor U1952 (N_1952,In_1134,In_1619);
xor U1953 (N_1953,In_196,In_1708);
or U1954 (N_1954,In_7,In_1940);
or U1955 (N_1955,In_1903,In_222);
nor U1956 (N_1956,In_408,In_1845);
or U1957 (N_1957,In_729,In_282);
nand U1958 (N_1958,In_362,In_1580);
nand U1959 (N_1959,In_1540,In_1632);
xor U1960 (N_1960,In_1418,In_984);
or U1961 (N_1961,In_57,In_739);
nand U1962 (N_1962,In_1317,In_314);
and U1963 (N_1963,In_1890,In_987);
nand U1964 (N_1964,In_13,In_1276);
nor U1965 (N_1965,In_1129,In_85);
nand U1966 (N_1966,In_1781,In_865);
xor U1967 (N_1967,In_1996,In_1858);
xor U1968 (N_1968,In_755,In_1504);
or U1969 (N_1969,In_174,In_615);
nand U1970 (N_1970,In_1731,In_617);
nor U1971 (N_1971,In_1674,In_264);
or U1972 (N_1972,In_252,In_490);
and U1973 (N_1973,In_425,In_895);
nand U1974 (N_1974,In_1274,In_562);
and U1975 (N_1975,In_876,In_446);
or U1976 (N_1976,In_715,In_1464);
nand U1977 (N_1977,In_596,In_875);
nor U1978 (N_1978,In_972,In_1448);
or U1979 (N_1979,In_1993,In_1184);
nand U1980 (N_1980,In_127,In_404);
and U1981 (N_1981,In_1608,In_1412);
and U1982 (N_1982,In_805,In_99);
xor U1983 (N_1983,In_456,In_1148);
or U1984 (N_1984,In_618,In_409);
and U1985 (N_1985,In_156,In_333);
nor U1986 (N_1986,In_1756,In_843);
nor U1987 (N_1987,In_1419,In_1645);
and U1988 (N_1988,In_1398,In_26);
and U1989 (N_1989,In_1486,In_1194);
or U1990 (N_1990,In_395,In_239);
or U1991 (N_1991,In_250,In_1838);
nor U1992 (N_1992,In_1204,In_578);
and U1993 (N_1993,In_1266,In_961);
nand U1994 (N_1994,In_680,In_1128);
and U1995 (N_1995,In_1173,In_722);
nand U1996 (N_1996,In_1361,In_1084);
and U1997 (N_1997,In_782,In_937);
or U1998 (N_1998,In_892,In_273);
or U1999 (N_1999,In_93,In_1708);
nand U2000 (N_2000,In_1485,In_412);
nor U2001 (N_2001,In_712,In_393);
nor U2002 (N_2002,In_673,In_903);
xnor U2003 (N_2003,In_902,In_631);
xor U2004 (N_2004,In_1485,In_1600);
and U2005 (N_2005,In_1443,In_1194);
nand U2006 (N_2006,In_446,In_1406);
or U2007 (N_2007,In_1220,In_1855);
or U2008 (N_2008,In_854,In_919);
nand U2009 (N_2009,In_1563,In_1784);
and U2010 (N_2010,In_1626,In_1571);
and U2011 (N_2011,In_1948,In_1535);
and U2012 (N_2012,In_1940,In_952);
or U2013 (N_2013,In_1732,In_1752);
or U2014 (N_2014,In_489,In_957);
and U2015 (N_2015,In_1969,In_703);
nor U2016 (N_2016,In_1627,In_998);
nor U2017 (N_2017,In_1267,In_1946);
nor U2018 (N_2018,In_632,In_1263);
and U2019 (N_2019,In_5,In_1779);
nand U2020 (N_2020,In_1903,In_798);
and U2021 (N_2021,In_1041,In_1279);
nand U2022 (N_2022,In_1137,In_480);
nand U2023 (N_2023,In_784,In_1632);
or U2024 (N_2024,In_690,In_8);
and U2025 (N_2025,In_724,In_164);
and U2026 (N_2026,In_591,In_1248);
nand U2027 (N_2027,In_204,In_1911);
and U2028 (N_2028,In_1974,In_268);
or U2029 (N_2029,In_1153,In_832);
and U2030 (N_2030,In_335,In_966);
and U2031 (N_2031,In_960,In_596);
and U2032 (N_2032,In_1286,In_1390);
xor U2033 (N_2033,In_839,In_25);
and U2034 (N_2034,In_811,In_1405);
and U2035 (N_2035,In_756,In_374);
or U2036 (N_2036,In_1300,In_35);
or U2037 (N_2037,In_1106,In_436);
nand U2038 (N_2038,In_712,In_1778);
and U2039 (N_2039,In_107,In_1468);
nand U2040 (N_2040,In_1683,In_1535);
nand U2041 (N_2041,In_1729,In_1574);
xor U2042 (N_2042,In_875,In_852);
nor U2043 (N_2043,In_1593,In_1559);
nor U2044 (N_2044,In_337,In_808);
xnor U2045 (N_2045,In_612,In_1163);
nor U2046 (N_2046,In_424,In_24);
and U2047 (N_2047,In_249,In_60);
nor U2048 (N_2048,In_86,In_564);
or U2049 (N_2049,In_361,In_765);
nor U2050 (N_2050,In_220,In_1824);
and U2051 (N_2051,In_1065,In_613);
nand U2052 (N_2052,In_1693,In_1446);
nand U2053 (N_2053,In_1922,In_446);
and U2054 (N_2054,In_1895,In_514);
nor U2055 (N_2055,In_1759,In_206);
or U2056 (N_2056,In_707,In_814);
nor U2057 (N_2057,In_313,In_439);
nor U2058 (N_2058,In_1078,In_1849);
nand U2059 (N_2059,In_1444,In_704);
or U2060 (N_2060,In_478,In_1671);
xor U2061 (N_2061,In_509,In_1661);
nor U2062 (N_2062,In_647,In_933);
xnor U2063 (N_2063,In_485,In_73);
nor U2064 (N_2064,In_309,In_1470);
nand U2065 (N_2065,In_894,In_389);
nor U2066 (N_2066,In_282,In_1383);
nor U2067 (N_2067,In_773,In_127);
or U2068 (N_2068,In_1031,In_1116);
nand U2069 (N_2069,In_1151,In_516);
and U2070 (N_2070,In_1960,In_1525);
nor U2071 (N_2071,In_1817,In_984);
and U2072 (N_2072,In_1615,In_486);
or U2073 (N_2073,In_939,In_608);
or U2074 (N_2074,In_1252,In_1553);
nand U2075 (N_2075,In_1395,In_1981);
nor U2076 (N_2076,In_1764,In_1811);
and U2077 (N_2077,In_805,In_1850);
nand U2078 (N_2078,In_287,In_211);
nor U2079 (N_2079,In_1476,In_1808);
nor U2080 (N_2080,In_163,In_601);
xor U2081 (N_2081,In_1095,In_1218);
nor U2082 (N_2082,In_87,In_1196);
nand U2083 (N_2083,In_754,In_1581);
nand U2084 (N_2084,In_1127,In_1879);
nand U2085 (N_2085,In_1531,In_1604);
nand U2086 (N_2086,In_180,In_1020);
xor U2087 (N_2087,In_405,In_1293);
xnor U2088 (N_2088,In_942,In_1637);
nand U2089 (N_2089,In_609,In_1379);
nand U2090 (N_2090,In_941,In_981);
or U2091 (N_2091,In_1979,In_1971);
nor U2092 (N_2092,In_390,In_496);
nand U2093 (N_2093,In_1449,In_198);
or U2094 (N_2094,In_1152,In_177);
or U2095 (N_2095,In_724,In_964);
nor U2096 (N_2096,In_1084,In_1845);
or U2097 (N_2097,In_1260,In_1949);
nor U2098 (N_2098,In_463,In_1174);
xnor U2099 (N_2099,In_1840,In_1519);
or U2100 (N_2100,In_904,In_1903);
nand U2101 (N_2101,In_121,In_1805);
or U2102 (N_2102,In_927,In_1872);
nor U2103 (N_2103,In_1946,In_54);
nor U2104 (N_2104,In_227,In_893);
xor U2105 (N_2105,In_1608,In_137);
and U2106 (N_2106,In_42,In_1780);
nor U2107 (N_2107,In_1273,In_1438);
nand U2108 (N_2108,In_1039,In_953);
xnor U2109 (N_2109,In_1630,In_1835);
and U2110 (N_2110,In_917,In_1321);
and U2111 (N_2111,In_1049,In_1767);
and U2112 (N_2112,In_1518,In_1987);
and U2113 (N_2113,In_747,In_1371);
or U2114 (N_2114,In_197,In_627);
or U2115 (N_2115,In_388,In_1148);
nand U2116 (N_2116,In_1271,In_208);
and U2117 (N_2117,In_127,In_468);
or U2118 (N_2118,In_1213,In_614);
xnor U2119 (N_2119,In_1853,In_680);
or U2120 (N_2120,In_1695,In_189);
nor U2121 (N_2121,In_245,In_988);
nand U2122 (N_2122,In_1163,In_1746);
nor U2123 (N_2123,In_574,In_102);
nor U2124 (N_2124,In_840,In_1229);
xor U2125 (N_2125,In_1267,In_879);
or U2126 (N_2126,In_286,In_252);
and U2127 (N_2127,In_439,In_1735);
or U2128 (N_2128,In_1473,In_382);
and U2129 (N_2129,In_1287,In_551);
and U2130 (N_2130,In_1871,In_1074);
nor U2131 (N_2131,In_140,In_1790);
nand U2132 (N_2132,In_833,In_1829);
and U2133 (N_2133,In_307,In_743);
or U2134 (N_2134,In_1601,In_469);
nand U2135 (N_2135,In_124,In_231);
or U2136 (N_2136,In_393,In_1180);
nor U2137 (N_2137,In_1330,In_526);
or U2138 (N_2138,In_743,In_588);
or U2139 (N_2139,In_551,In_454);
and U2140 (N_2140,In_1282,In_17);
and U2141 (N_2141,In_1794,In_542);
and U2142 (N_2142,In_1378,In_66);
nor U2143 (N_2143,In_630,In_1257);
and U2144 (N_2144,In_1708,In_128);
nor U2145 (N_2145,In_1824,In_1131);
or U2146 (N_2146,In_110,In_542);
and U2147 (N_2147,In_511,In_1587);
and U2148 (N_2148,In_991,In_732);
nand U2149 (N_2149,In_1682,In_659);
and U2150 (N_2150,In_1559,In_442);
nor U2151 (N_2151,In_1836,In_551);
xor U2152 (N_2152,In_1065,In_669);
nor U2153 (N_2153,In_1361,In_34);
nor U2154 (N_2154,In_782,In_1339);
or U2155 (N_2155,In_1090,In_1083);
nand U2156 (N_2156,In_130,In_1000);
nor U2157 (N_2157,In_1381,In_202);
or U2158 (N_2158,In_779,In_729);
or U2159 (N_2159,In_1792,In_410);
and U2160 (N_2160,In_1328,In_80);
or U2161 (N_2161,In_1692,In_123);
nor U2162 (N_2162,In_1073,In_313);
or U2163 (N_2163,In_1291,In_511);
nand U2164 (N_2164,In_310,In_1903);
nor U2165 (N_2165,In_1708,In_896);
or U2166 (N_2166,In_746,In_1852);
nor U2167 (N_2167,In_1170,In_1408);
nor U2168 (N_2168,In_565,In_95);
nor U2169 (N_2169,In_857,In_1288);
xnor U2170 (N_2170,In_35,In_1635);
nand U2171 (N_2171,In_905,In_120);
or U2172 (N_2172,In_1910,In_563);
and U2173 (N_2173,In_772,In_499);
and U2174 (N_2174,In_1102,In_1648);
nand U2175 (N_2175,In_1556,In_553);
or U2176 (N_2176,In_1655,In_215);
nor U2177 (N_2177,In_798,In_1676);
xor U2178 (N_2178,In_1773,In_53);
and U2179 (N_2179,In_247,In_86);
or U2180 (N_2180,In_1412,In_1213);
nand U2181 (N_2181,In_878,In_892);
nor U2182 (N_2182,In_1399,In_733);
nand U2183 (N_2183,In_1503,In_1951);
and U2184 (N_2184,In_1616,In_1951);
and U2185 (N_2185,In_1019,In_1204);
or U2186 (N_2186,In_1236,In_1622);
xor U2187 (N_2187,In_1299,In_1968);
or U2188 (N_2188,In_1051,In_1197);
nor U2189 (N_2189,In_653,In_1506);
and U2190 (N_2190,In_1180,In_107);
nand U2191 (N_2191,In_847,In_506);
nor U2192 (N_2192,In_1225,In_703);
and U2193 (N_2193,In_1256,In_239);
nand U2194 (N_2194,In_1843,In_1022);
and U2195 (N_2195,In_301,In_669);
nor U2196 (N_2196,In_510,In_409);
or U2197 (N_2197,In_1113,In_1411);
or U2198 (N_2198,In_1804,In_1204);
nor U2199 (N_2199,In_45,In_646);
or U2200 (N_2200,In_1238,In_563);
or U2201 (N_2201,In_1327,In_1016);
or U2202 (N_2202,In_1768,In_1440);
nand U2203 (N_2203,In_1161,In_746);
or U2204 (N_2204,In_1453,In_480);
nor U2205 (N_2205,In_703,In_1037);
or U2206 (N_2206,In_1504,In_801);
nand U2207 (N_2207,In_576,In_224);
nand U2208 (N_2208,In_1965,In_1305);
or U2209 (N_2209,In_819,In_1805);
or U2210 (N_2210,In_948,In_1664);
nand U2211 (N_2211,In_929,In_1540);
nand U2212 (N_2212,In_989,In_1931);
nor U2213 (N_2213,In_358,In_1285);
nor U2214 (N_2214,In_214,In_1363);
or U2215 (N_2215,In_685,In_814);
and U2216 (N_2216,In_1155,In_1255);
or U2217 (N_2217,In_1341,In_579);
or U2218 (N_2218,In_366,In_1680);
nor U2219 (N_2219,In_946,In_189);
nand U2220 (N_2220,In_1631,In_238);
or U2221 (N_2221,In_1413,In_931);
nor U2222 (N_2222,In_158,In_1054);
nor U2223 (N_2223,In_1385,In_412);
or U2224 (N_2224,In_1412,In_183);
or U2225 (N_2225,In_316,In_1910);
nor U2226 (N_2226,In_922,In_183);
or U2227 (N_2227,In_233,In_908);
nor U2228 (N_2228,In_160,In_1358);
and U2229 (N_2229,In_396,In_312);
nor U2230 (N_2230,In_1329,In_321);
nor U2231 (N_2231,In_1107,In_1934);
nand U2232 (N_2232,In_1842,In_569);
nand U2233 (N_2233,In_769,In_1694);
and U2234 (N_2234,In_116,In_808);
or U2235 (N_2235,In_1358,In_394);
and U2236 (N_2236,In_1333,In_766);
or U2237 (N_2237,In_211,In_636);
and U2238 (N_2238,In_473,In_1898);
or U2239 (N_2239,In_188,In_921);
nor U2240 (N_2240,In_1942,In_1132);
and U2241 (N_2241,In_1588,In_884);
and U2242 (N_2242,In_516,In_405);
and U2243 (N_2243,In_1469,In_593);
nand U2244 (N_2244,In_1022,In_648);
and U2245 (N_2245,In_1380,In_1897);
nand U2246 (N_2246,In_1830,In_161);
or U2247 (N_2247,In_1283,In_1153);
nand U2248 (N_2248,In_706,In_1336);
and U2249 (N_2249,In_1280,In_942);
xnor U2250 (N_2250,In_425,In_1286);
and U2251 (N_2251,In_1718,In_1847);
nand U2252 (N_2252,In_1208,In_1417);
xor U2253 (N_2253,In_101,In_69);
nand U2254 (N_2254,In_528,In_1427);
xnor U2255 (N_2255,In_191,In_1666);
and U2256 (N_2256,In_9,In_1143);
or U2257 (N_2257,In_365,In_1519);
and U2258 (N_2258,In_56,In_1937);
or U2259 (N_2259,In_1306,In_1796);
and U2260 (N_2260,In_863,In_471);
or U2261 (N_2261,In_1250,In_282);
nor U2262 (N_2262,In_1999,In_1493);
nor U2263 (N_2263,In_869,In_282);
and U2264 (N_2264,In_77,In_814);
nand U2265 (N_2265,In_713,In_221);
or U2266 (N_2266,In_1224,In_1957);
or U2267 (N_2267,In_529,In_153);
nand U2268 (N_2268,In_955,In_566);
nor U2269 (N_2269,In_1380,In_1050);
nand U2270 (N_2270,In_293,In_1114);
xnor U2271 (N_2271,In_457,In_103);
nor U2272 (N_2272,In_1095,In_970);
and U2273 (N_2273,In_1265,In_1143);
or U2274 (N_2274,In_1871,In_645);
nand U2275 (N_2275,In_1670,In_667);
nand U2276 (N_2276,In_938,In_1766);
xor U2277 (N_2277,In_1055,In_659);
xor U2278 (N_2278,In_1446,In_448);
nand U2279 (N_2279,In_762,In_135);
or U2280 (N_2280,In_341,In_1572);
or U2281 (N_2281,In_307,In_662);
and U2282 (N_2282,In_797,In_123);
or U2283 (N_2283,In_913,In_1961);
or U2284 (N_2284,In_223,In_1282);
or U2285 (N_2285,In_400,In_1396);
or U2286 (N_2286,In_1428,In_1703);
nand U2287 (N_2287,In_736,In_603);
xor U2288 (N_2288,In_1731,In_279);
xnor U2289 (N_2289,In_677,In_1234);
xnor U2290 (N_2290,In_675,In_629);
nor U2291 (N_2291,In_193,In_125);
or U2292 (N_2292,In_1774,In_1339);
and U2293 (N_2293,In_1583,In_1749);
or U2294 (N_2294,In_1902,In_831);
nor U2295 (N_2295,In_387,In_199);
nand U2296 (N_2296,In_1333,In_379);
nor U2297 (N_2297,In_1178,In_1896);
and U2298 (N_2298,In_27,In_202);
nor U2299 (N_2299,In_1755,In_1396);
nand U2300 (N_2300,In_1141,In_1927);
or U2301 (N_2301,In_1102,In_168);
nor U2302 (N_2302,In_1512,In_199);
and U2303 (N_2303,In_1224,In_1778);
xnor U2304 (N_2304,In_1264,In_1100);
and U2305 (N_2305,In_1200,In_858);
nor U2306 (N_2306,In_1213,In_1406);
nand U2307 (N_2307,In_1371,In_997);
and U2308 (N_2308,In_7,In_146);
xor U2309 (N_2309,In_119,In_1115);
or U2310 (N_2310,In_770,In_1176);
and U2311 (N_2311,In_1806,In_965);
nand U2312 (N_2312,In_1036,In_207);
nand U2313 (N_2313,In_505,In_358);
or U2314 (N_2314,In_1493,In_1663);
nor U2315 (N_2315,In_1623,In_1077);
or U2316 (N_2316,In_1446,In_1762);
nor U2317 (N_2317,In_342,In_697);
and U2318 (N_2318,In_1893,In_545);
and U2319 (N_2319,In_1251,In_497);
or U2320 (N_2320,In_84,In_1469);
nor U2321 (N_2321,In_1032,In_1191);
nand U2322 (N_2322,In_855,In_1784);
nand U2323 (N_2323,In_1090,In_1207);
nor U2324 (N_2324,In_190,In_1116);
and U2325 (N_2325,In_1213,In_954);
or U2326 (N_2326,In_532,In_839);
or U2327 (N_2327,In_635,In_1481);
nand U2328 (N_2328,In_1953,In_1190);
nand U2329 (N_2329,In_1164,In_280);
xnor U2330 (N_2330,In_1991,In_277);
and U2331 (N_2331,In_1380,In_1102);
and U2332 (N_2332,In_483,In_1974);
nor U2333 (N_2333,In_838,In_212);
nor U2334 (N_2334,In_364,In_583);
nor U2335 (N_2335,In_496,In_848);
or U2336 (N_2336,In_643,In_64);
and U2337 (N_2337,In_1055,In_1617);
nand U2338 (N_2338,In_1397,In_1323);
xor U2339 (N_2339,In_920,In_356);
and U2340 (N_2340,In_1212,In_603);
nand U2341 (N_2341,In_81,In_1818);
nor U2342 (N_2342,In_1903,In_900);
nor U2343 (N_2343,In_902,In_1577);
nor U2344 (N_2344,In_719,In_1655);
and U2345 (N_2345,In_403,In_1963);
and U2346 (N_2346,In_649,In_221);
or U2347 (N_2347,In_102,In_448);
and U2348 (N_2348,In_455,In_286);
or U2349 (N_2349,In_466,In_691);
nand U2350 (N_2350,In_1791,In_1841);
or U2351 (N_2351,In_1,In_1392);
or U2352 (N_2352,In_454,In_148);
nand U2353 (N_2353,In_334,In_1877);
nand U2354 (N_2354,In_684,In_1610);
nor U2355 (N_2355,In_1484,In_137);
nor U2356 (N_2356,In_1783,In_415);
nand U2357 (N_2357,In_150,In_440);
or U2358 (N_2358,In_375,In_1484);
and U2359 (N_2359,In_1085,In_678);
or U2360 (N_2360,In_478,In_1160);
nor U2361 (N_2361,In_1780,In_530);
nand U2362 (N_2362,In_32,In_1993);
or U2363 (N_2363,In_18,In_1258);
or U2364 (N_2364,In_322,In_445);
xnor U2365 (N_2365,In_1757,In_531);
or U2366 (N_2366,In_401,In_1005);
nand U2367 (N_2367,In_1591,In_75);
and U2368 (N_2368,In_1096,In_672);
nor U2369 (N_2369,In_773,In_1822);
or U2370 (N_2370,In_336,In_1607);
nand U2371 (N_2371,In_1745,In_1838);
or U2372 (N_2372,In_1191,In_1064);
nand U2373 (N_2373,In_871,In_1829);
nand U2374 (N_2374,In_1728,In_109);
nor U2375 (N_2375,In_1777,In_1949);
nand U2376 (N_2376,In_116,In_14);
nand U2377 (N_2377,In_819,In_1316);
and U2378 (N_2378,In_929,In_242);
nor U2379 (N_2379,In_1779,In_804);
and U2380 (N_2380,In_162,In_1583);
nand U2381 (N_2381,In_633,In_1719);
and U2382 (N_2382,In_1672,In_330);
and U2383 (N_2383,In_1636,In_1353);
nor U2384 (N_2384,In_83,In_710);
or U2385 (N_2385,In_1928,In_1337);
nand U2386 (N_2386,In_618,In_1301);
xnor U2387 (N_2387,In_712,In_323);
nand U2388 (N_2388,In_70,In_365);
nand U2389 (N_2389,In_1979,In_1042);
and U2390 (N_2390,In_1316,In_1722);
nor U2391 (N_2391,In_1755,In_673);
nand U2392 (N_2392,In_713,In_570);
or U2393 (N_2393,In_955,In_1471);
xor U2394 (N_2394,In_1350,In_1186);
nand U2395 (N_2395,In_445,In_1263);
nand U2396 (N_2396,In_1446,In_15);
and U2397 (N_2397,In_282,In_454);
nand U2398 (N_2398,In_939,In_1607);
and U2399 (N_2399,In_919,In_482);
or U2400 (N_2400,In_121,In_328);
nand U2401 (N_2401,In_774,In_220);
nand U2402 (N_2402,In_490,In_1113);
and U2403 (N_2403,In_1147,In_1740);
nand U2404 (N_2404,In_779,In_612);
and U2405 (N_2405,In_1292,In_1495);
nand U2406 (N_2406,In_1902,In_1282);
and U2407 (N_2407,In_1582,In_1602);
nor U2408 (N_2408,In_1094,In_535);
nand U2409 (N_2409,In_810,In_1708);
xnor U2410 (N_2410,In_1914,In_837);
xnor U2411 (N_2411,In_549,In_546);
nand U2412 (N_2412,In_1185,In_346);
nor U2413 (N_2413,In_462,In_1770);
nand U2414 (N_2414,In_1975,In_690);
xor U2415 (N_2415,In_689,In_739);
nand U2416 (N_2416,In_676,In_1902);
and U2417 (N_2417,In_1850,In_1947);
nor U2418 (N_2418,In_745,In_1470);
and U2419 (N_2419,In_1360,In_313);
xnor U2420 (N_2420,In_1075,In_1120);
nor U2421 (N_2421,In_1493,In_1044);
and U2422 (N_2422,In_1389,In_696);
and U2423 (N_2423,In_1254,In_167);
and U2424 (N_2424,In_244,In_1074);
nand U2425 (N_2425,In_1723,In_1498);
or U2426 (N_2426,In_129,In_673);
nor U2427 (N_2427,In_535,In_407);
nor U2428 (N_2428,In_1203,In_1436);
and U2429 (N_2429,In_1154,In_2);
nand U2430 (N_2430,In_1007,In_1452);
and U2431 (N_2431,In_588,In_1852);
and U2432 (N_2432,In_65,In_1224);
nor U2433 (N_2433,In_1131,In_1181);
or U2434 (N_2434,In_616,In_1409);
and U2435 (N_2435,In_1978,In_1459);
nor U2436 (N_2436,In_1656,In_1221);
nand U2437 (N_2437,In_230,In_1525);
nor U2438 (N_2438,In_1065,In_1674);
nand U2439 (N_2439,In_526,In_28);
or U2440 (N_2440,In_885,In_875);
nor U2441 (N_2441,In_1995,In_58);
nand U2442 (N_2442,In_145,In_1606);
and U2443 (N_2443,In_1601,In_771);
nand U2444 (N_2444,In_1149,In_270);
nand U2445 (N_2445,In_1992,In_627);
or U2446 (N_2446,In_376,In_362);
nor U2447 (N_2447,In_1846,In_1383);
nor U2448 (N_2448,In_1743,In_183);
or U2449 (N_2449,In_1502,In_1127);
xnor U2450 (N_2450,In_1404,In_137);
and U2451 (N_2451,In_458,In_1799);
nor U2452 (N_2452,In_898,In_1689);
nand U2453 (N_2453,In_1014,In_1405);
nor U2454 (N_2454,In_1932,In_1631);
nor U2455 (N_2455,In_1891,In_897);
and U2456 (N_2456,In_1723,In_63);
and U2457 (N_2457,In_291,In_1765);
nand U2458 (N_2458,In_571,In_164);
nor U2459 (N_2459,In_683,In_1959);
and U2460 (N_2460,In_969,In_1980);
and U2461 (N_2461,In_669,In_992);
nor U2462 (N_2462,In_355,In_1791);
nand U2463 (N_2463,In_1842,In_730);
xor U2464 (N_2464,In_1724,In_302);
nor U2465 (N_2465,In_1428,In_395);
and U2466 (N_2466,In_1968,In_1760);
or U2467 (N_2467,In_343,In_865);
and U2468 (N_2468,In_1244,In_85);
or U2469 (N_2469,In_1054,In_768);
nor U2470 (N_2470,In_92,In_1942);
nor U2471 (N_2471,In_1550,In_306);
nor U2472 (N_2472,In_1559,In_450);
nand U2473 (N_2473,In_787,In_1164);
and U2474 (N_2474,In_1172,In_241);
or U2475 (N_2475,In_369,In_1858);
or U2476 (N_2476,In_1730,In_40);
or U2477 (N_2477,In_1768,In_635);
xnor U2478 (N_2478,In_1461,In_1576);
or U2479 (N_2479,In_240,In_1872);
and U2480 (N_2480,In_432,In_726);
xor U2481 (N_2481,In_51,In_997);
nor U2482 (N_2482,In_280,In_1996);
and U2483 (N_2483,In_74,In_1479);
nand U2484 (N_2484,In_863,In_543);
or U2485 (N_2485,In_270,In_1028);
xor U2486 (N_2486,In_1400,In_837);
or U2487 (N_2487,In_610,In_1288);
and U2488 (N_2488,In_1029,In_1522);
and U2489 (N_2489,In_836,In_354);
and U2490 (N_2490,In_468,In_1638);
or U2491 (N_2491,In_1727,In_1231);
nand U2492 (N_2492,In_648,In_493);
nand U2493 (N_2493,In_1933,In_301);
nor U2494 (N_2494,In_874,In_770);
and U2495 (N_2495,In_625,In_1543);
nand U2496 (N_2496,In_142,In_1021);
and U2497 (N_2497,In_608,In_195);
and U2498 (N_2498,In_1176,In_1591);
or U2499 (N_2499,In_190,In_1834);
nand U2500 (N_2500,In_1556,In_1177);
and U2501 (N_2501,In_968,In_1102);
and U2502 (N_2502,In_1198,In_825);
or U2503 (N_2503,In_1817,In_182);
nand U2504 (N_2504,In_731,In_778);
xnor U2505 (N_2505,In_1809,In_1899);
nand U2506 (N_2506,In_592,In_417);
nor U2507 (N_2507,In_1355,In_1823);
xnor U2508 (N_2508,In_1292,In_767);
or U2509 (N_2509,In_181,In_1512);
and U2510 (N_2510,In_1788,In_1383);
nor U2511 (N_2511,In_630,In_819);
and U2512 (N_2512,In_1140,In_1496);
or U2513 (N_2513,In_1661,In_1228);
nand U2514 (N_2514,In_311,In_704);
nand U2515 (N_2515,In_546,In_1430);
nand U2516 (N_2516,In_359,In_1340);
or U2517 (N_2517,In_1076,In_1426);
xor U2518 (N_2518,In_1962,In_1495);
or U2519 (N_2519,In_11,In_16);
and U2520 (N_2520,In_155,In_1412);
and U2521 (N_2521,In_1411,In_718);
nand U2522 (N_2522,In_613,In_1252);
and U2523 (N_2523,In_460,In_1758);
xor U2524 (N_2524,In_1095,In_786);
and U2525 (N_2525,In_491,In_1801);
xnor U2526 (N_2526,In_1857,In_1370);
xnor U2527 (N_2527,In_146,In_1285);
or U2528 (N_2528,In_1589,In_1747);
and U2529 (N_2529,In_529,In_975);
nor U2530 (N_2530,In_1744,In_100);
or U2531 (N_2531,In_580,In_677);
and U2532 (N_2532,In_1399,In_1655);
or U2533 (N_2533,In_149,In_1979);
or U2534 (N_2534,In_28,In_445);
nand U2535 (N_2535,In_1798,In_859);
or U2536 (N_2536,In_544,In_246);
or U2537 (N_2537,In_261,In_1806);
nand U2538 (N_2538,In_458,In_983);
or U2539 (N_2539,In_1387,In_1728);
nor U2540 (N_2540,In_1820,In_1557);
nor U2541 (N_2541,In_662,In_970);
and U2542 (N_2542,In_834,In_1133);
or U2543 (N_2543,In_1454,In_1835);
or U2544 (N_2544,In_843,In_1304);
or U2545 (N_2545,In_683,In_1577);
nand U2546 (N_2546,In_1304,In_1467);
or U2547 (N_2547,In_537,In_1917);
nand U2548 (N_2548,In_628,In_45);
or U2549 (N_2549,In_1770,In_1711);
nand U2550 (N_2550,In_1128,In_1071);
nor U2551 (N_2551,In_964,In_1678);
nor U2552 (N_2552,In_120,In_1371);
nor U2553 (N_2553,In_420,In_1533);
nand U2554 (N_2554,In_1469,In_990);
nand U2555 (N_2555,In_233,In_1866);
nor U2556 (N_2556,In_135,In_1753);
nor U2557 (N_2557,In_1840,In_1536);
nor U2558 (N_2558,In_1131,In_489);
or U2559 (N_2559,In_1633,In_1910);
nor U2560 (N_2560,In_621,In_49);
nand U2561 (N_2561,In_1604,In_1611);
or U2562 (N_2562,In_495,In_677);
or U2563 (N_2563,In_1225,In_1095);
nor U2564 (N_2564,In_790,In_194);
and U2565 (N_2565,In_1175,In_564);
and U2566 (N_2566,In_1822,In_1107);
xor U2567 (N_2567,In_1485,In_1469);
or U2568 (N_2568,In_469,In_840);
or U2569 (N_2569,In_1435,In_1378);
nand U2570 (N_2570,In_1279,In_1296);
or U2571 (N_2571,In_807,In_1761);
nor U2572 (N_2572,In_221,In_176);
nand U2573 (N_2573,In_1046,In_178);
nand U2574 (N_2574,In_37,In_1111);
nor U2575 (N_2575,In_245,In_581);
nand U2576 (N_2576,In_1155,In_607);
xor U2577 (N_2577,In_585,In_1945);
or U2578 (N_2578,In_596,In_1623);
or U2579 (N_2579,In_14,In_74);
nand U2580 (N_2580,In_179,In_346);
and U2581 (N_2581,In_1410,In_597);
nor U2582 (N_2582,In_478,In_1574);
nor U2583 (N_2583,In_1396,In_854);
or U2584 (N_2584,In_1114,In_374);
nor U2585 (N_2585,In_442,In_1435);
and U2586 (N_2586,In_1900,In_1372);
nand U2587 (N_2587,In_1126,In_81);
nor U2588 (N_2588,In_480,In_1424);
nor U2589 (N_2589,In_810,In_1704);
nand U2590 (N_2590,In_240,In_1134);
or U2591 (N_2591,In_988,In_898);
or U2592 (N_2592,In_1072,In_122);
nor U2593 (N_2593,In_681,In_1457);
nor U2594 (N_2594,In_1601,In_228);
or U2595 (N_2595,In_365,In_1837);
or U2596 (N_2596,In_1853,In_1174);
or U2597 (N_2597,In_1708,In_925);
nand U2598 (N_2598,In_261,In_1853);
nand U2599 (N_2599,In_1597,In_1684);
or U2600 (N_2600,In_1180,In_552);
nor U2601 (N_2601,In_1494,In_982);
xnor U2602 (N_2602,In_37,In_1191);
nor U2603 (N_2603,In_1357,In_89);
or U2604 (N_2604,In_1822,In_470);
nand U2605 (N_2605,In_1739,In_1089);
and U2606 (N_2606,In_1915,In_1577);
and U2607 (N_2607,In_157,In_1997);
nand U2608 (N_2608,In_1272,In_1546);
and U2609 (N_2609,In_978,In_1151);
or U2610 (N_2610,In_1080,In_553);
nor U2611 (N_2611,In_1084,In_1942);
or U2612 (N_2612,In_1082,In_455);
nand U2613 (N_2613,In_1375,In_800);
nor U2614 (N_2614,In_563,In_279);
and U2615 (N_2615,In_1034,In_1832);
xnor U2616 (N_2616,In_1667,In_839);
and U2617 (N_2617,In_916,In_1732);
or U2618 (N_2618,In_31,In_259);
or U2619 (N_2619,In_1093,In_1192);
nand U2620 (N_2620,In_262,In_366);
or U2621 (N_2621,In_899,In_992);
nor U2622 (N_2622,In_634,In_401);
nand U2623 (N_2623,In_1668,In_528);
nor U2624 (N_2624,In_42,In_503);
nand U2625 (N_2625,In_457,In_44);
nand U2626 (N_2626,In_833,In_398);
nor U2627 (N_2627,In_917,In_641);
nand U2628 (N_2628,In_1653,In_1075);
or U2629 (N_2629,In_90,In_573);
nor U2630 (N_2630,In_913,In_1102);
nor U2631 (N_2631,In_1575,In_1766);
or U2632 (N_2632,In_1840,In_1058);
nor U2633 (N_2633,In_406,In_70);
nor U2634 (N_2634,In_1017,In_220);
xnor U2635 (N_2635,In_1718,In_1084);
or U2636 (N_2636,In_340,In_547);
xnor U2637 (N_2637,In_379,In_544);
or U2638 (N_2638,In_1035,In_503);
xor U2639 (N_2639,In_659,In_1896);
nand U2640 (N_2640,In_652,In_1414);
nand U2641 (N_2641,In_851,In_1524);
or U2642 (N_2642,In_404,In_1742);
or U2643 (N_2643,In_594,In_291);
or U2644 (N_2644,In_1007,In_1465);
or U2645 (N_2645,In_1691,In_271);
or U2646 (N_2646,In_1844,In_566);
and U2647 (N_2647,In_686,In_1687);
or U2648 (N_2648,In_1936,In_930);
nand U2649 (N_2649,In_1720,In_898);
nor U2650 (N_2650,In_1439,In_454);
nor U2651 (N_2651,In_1472,In_974);
or U2652 (N_2652,In_372,In_897);
nor U2653 (N_2653,In_518,In_1201);
and U2654 (N_2654,In_693,In_1519);
or U2655 (N_2655,In_537,In_1531);
nor U2656 (N_2656,In_990,In_519);
nand U2657 (N_2657,In_1735,In_736);
or U2658 (N_2658,In_1612,In_587);
nor U2659 (N_2659,In_1268,In_31);
or U2660 (N_2660,In_808,In_1056);
nand U2661 (N_2661,In_1939,In_307);
xnor U2662 (N_2662,In_1433,In_1243);
nor U2663 (N_2663,In_1683,In_1366);
xnor U2664 (N_2664,In_762,In_1858);
or U2665 (N_2665,In_57,In_1091);
or U2666 (N_2666,In_880,In_1637);
nand U2667 (N_2667,In_881,In_1608);
or U2668 (N_2668,In_1268,In_982);
or U2669 (N_2669,In_1791,In_1729);
and U2670 (N_2670,In_1217,In_1055);
nand U2671 (N_2671,In_557,In_1771);
nor U2672 (N_2672,In_912,In_1219);
nor U2673 (N_2673,In_405,In_1978);
xor U2674 (N_2674,In_1112,In_1259);
nand U2675 (N_2675,In_1772,In_1574);
nor U2676 (N_2676,In_1299,In_927);
nand U2677 (N_2677,In_470,In_733);
nor U2678 (N_2678,In_1936,In_1166);
and U2679 (N_2679,In_1369,In_303);
nand U2680 (N_2680,In_363,In_396);
nor U2681 (N_2681,In_427,In_1832);
nor U2682 (N_2682,In_1482,In_637);
and U2683 (N_2683,In_101,In_1866);
and U2684 (N_2684,In_1557,In_83);
nor U2685 (N_2685,In_1005,In_1346);
nand U2686 (N_2686,In_1858,In_1335);
and U2687 (N_2687,In_1780,In_823);
nand U2688 (N_2688,In_1658,In_1050);
nand U2689 (N_2689,In_1952,In_1845);
nand U2690 (N_2690,In_1133,In_303);
nand U2691 (N_2691,In_620,In_1670);
or U2692 (N_2692,In_1758,In_348);
and U2693 (N_2693,In_87,In_331);
and U2694 (N_2694,In_535,In_432);
or U2695 (N_2695,In_1513,In_473);
nor U2696 (N_2696,In_1409,In_1328);
and U2697 (N_2697,In_469,In_1783);
xnor U2698 (N_2698,In_886,In_681);
nand U2699 (N_2699,In_676,In_130);
nor U2700 (N_2700,In_1366,In_1959);
nor U2701 (N_2701,In_1854,In_1329);
nor U2702 (N_2702,In_1570,In_1631);
nor U2703 (N_2703,In_381,In_1587);
or U2704 (N_2704,In_1689,In_1999);
xnor U2705 (N_2705,In_1162,In_1234);
nor U2706 (N_2706,In_99,In_1030);
and U2707 (N_2707,In_1005,In_349);
nand U2708 (N_2708,In_1497,In_1394);
nor U2709 (N_2709,In_781,In_1219);
and U2710 (N_2710,In_831,In_337);
or U2711 (N_2711,In_89,In_150);
and U2712 (N_2712,In_669,In_1198);
nor U2713 (N_2713,In_457,In_57);
or U2714 (N_2714,In_1543,In_883);
nor U2715 (N_2715,In_302,In_1039);
or U2716 (N_2716,In_497,In_314);
nand U2717 (N_2717,In_475,In_1270);
nor U2718 (N_2718,In_1353,In_155);
nand U2719 (N_2719,In_1528,In_1285);
nor U2720 (N_2720,In_354,In_1686);
xor U2721 (N_2721,In_567,In_1068);
nor U2722 (N_2722,In_1175,In_1070);
and U2723 (N_2723,In_939,In_1636);
or U2724 (N_2724,In_1109,In_524);
xnor U2725 (N_2725,In_1815,In_239);
nand U2726 (N_2726,In_1827,In_624);
nand U2727 (N_2727,In_166,In_458);
nand U2728 (N_2728,In_117,In_1693);
nor U2729 (N_2729,In_735,In_45);
nor U2730 (N_2730,In_914,In_1205);
xor U2731 (N_2731,In_529,In_813);
and U2732 (N_2732,In_1052,In_1078);
nand U2733 (N_2733,In_1024,In_1252);
and U2734 (N_2734,In_206,In_1785);
nand U2735 (N_2735,In_868,In_1118);
nand U2736 (N_2736,In_540,In_66);
and U2737 (N_2737,In_304,In_373);
nand U2738 (N_2738,In_646,In_67);
or U2739 (N_2739,In_1507,In_369);
nor U2740 (N_2740,In_1721,In_846);
nand U2741 (N_2741,In_404,In_1611);
xnor U2742 (N_2742,In_748,In_1348);
xnor U2743 (N_2743,In_579,In_849);
and U2744 (N_2744,In_325,In_1679);
and U2745 (N_2745,In_446,In_202);
or U2746 (N_2746,In_1911,In_1309);
and U2747 (N_2747,In_380,In_1030);
and U2748 (N_2748,In_822,In_580);
and U2749 (N_2749,In_766,In_955);
nor U2750 (N_2750,In_861,In_946);
nor U2751 (N_2751,In_127,In_1783);
and U2752 (N_2752,In_221,In_1301);
or U2753 (N_2753,In_1115,In_228);
nand U2754 (N_2754,In_131,In_1184);
or U2755 (N_2755,In_952,In_892);
and U2756 (N_2756,In_1324,In_473);
or U2757 (N_2757,In_135,In_1109);
and U2758 (N_2758,In_150,In_129);
or U2759 (N_2759,In_653,In_173);
and U2760 (N_2760,In_1874,In_711);
nand U2761 (N_2761,In_450,In_1018);
or U2762 (N_2762,In_1756,In_576);
or U2763 (N_2763,In_560,In_1129);
nand U2764 (N_2764,In_1087,In_475);
or U2765 (N_2765,In_357,In_242);
or U2766 (N_2766,In_958,In_685);
or U2767 (N_2767,In_1226,In_1946);
or U2768 (N_2768,In_1663,In_1781);
nor U2769 (N_2769,In_1178,In_1988);
or U2770 (N_2770,In_761,In_1126);
nand U2771 (N_2771,In_1204,In_4);
nor U2772 (N_2772,In_1653,In_406);
xor U2773 (N_2773,In_1015,In_1647);
and U2774 (N_2774,In_422,In_186);
nor U2775 (N_2775,In_1060,In_912);
nand U2776 (N_2776,In_619,In_1376);
and U2777 (N_2777,In_822,In_73);
nand U2778 (N_2778,In_1668,In_1989);
and U2779 (N_2779,In_1080,In_1767);
and U2780 (N_2780,In_436,In_11);
and U2781 (N_2781,In_1958,In_602);
nor U2782 (N_2782,In_1191,In_1584);
nor U2783 (N_2783,In_1809,In_236);
and U2784 (N_2784,In_0,In_1986);
nor U2785 (N_2785,In_1382,In_1846);
and U2786 (N_2786,In_1384,In_1250);
and U2787 (N_2787,In_1339,In_1776);
nor U2788 (N_2788,In_967,In_470);
or U2789 (N_2789,In_56,In_1291);
or U2790 (N_2790,In_788,In_936);
or U2791 (N_2791,In_1014,In_987);
or U2792 (N_2792,In_1955,In_1774);
nor U2793 (N_2793,In_187,In_513);
nand U2794 (N_2794,In_192,In_1750);
or U2795 (N_2795,In_833,In_1347);
nand U2796 (N_2796,In_309,In_1024);
or U2797 (N_2797,In_1919,In_1359);
xnor U2798 (N_2798,In_1851,In_398);
and U2799 (N_2799,In_585,In_939);
nor U2800 (N_2800,In_1442,In_1657);
or U2801 (N_2801,In_1346,In_1051);
and U2802 (N_2802,In_812,In_957);
nor U2803 (N_2803,In_1424,In_1840);
nand U2804 (N_2804,In_1385,In_41);
or U2805 (N_2805,In_1284,In_1403);
xor U2806 (N_2806,In_44,In_989);
or U2807 (N_2807,In_1765,In_15);
or U2808 (N_2808,In_1828,In_1096);
or U2809 (N_2809,In_1161,In_54);
nand U2810 (N_2810,In_849,In_813);
nand U2811 (N_2811,In_457,In_1620);
and U2812 (N_2812,In_192,In_728);
xor U2813 (N_2813,In_80,In_449);
xnor U2814 (N_2814,In_1003,In_316);
nor U2815 (N_2815,In_151,In_1515);
nor U2816 (N_2816,In_46,In_703);
xnor U2817 (N_2817,In_34,In_1880);
nor U2818 (N_2818,In_512,In_1992);
and U2819 (N_2819,In_1042,In_126);
or U2820 (N_2820,In_1144,In_1606);
nor U2821 (N_2821,In_1618,In_1696);
and U2822 (N_2822,In_1499,In_1762);
or U2823 (N_2823,In_1795,In_1707);
or U2824 (N_2824,In_1342,In_1391);
nand U2825 (N_2825,In_412,In_965);
and U2826 (N_2826,In_231,In_923);
or U2827 (N_2827,In_812,In_1843);
or U2828 (N_2828,In_1772,In_176);
nand U2829 (N_2829,In_1372,In_453);
and U2830 (N_2830,In_848,In_352);
nand U2831 (N_2831,In_1718,In_1187);
or U2832 (N_2832,In_1306,In_702);
and U2833 (N_2833,In_1326,In_1295);
and U2834 (N_2834,In_425,In_1977);
or U2835 (N_2835,In_1116,In_307);
or U2836 (N_2836,In_559,In_491);
and U2837 (N_2837,In_171,In_844);
nor U2838 (N_2838,In_1388,In_1952);
or U2839 (N_2839,In_1950,In_746);
nand U2840 (N_2840,In_311,In_7);
nor U2841 (N_2841,In_1418,In_1529);
nor U2842 (N_2842,In_1554,In_1340);
nand U2843 (N_2843,In_263,In_123);
nor U2844 (N_2844,In_931,In_1400);
and U2845 (N_2845,In_765,In_1480);
and U2846 (N_2846,In_101,In_1891);
nand U2847 (N_2847,In_699,In_588);
xnor U2848 (N_2848,In_1422,In_736);
nor U2849 (N_2849,In_307,In_127);
nand U2850 (N_2850,In_864,In_57);
or U2851 (N_2851,In_220,In_640);
and U2852 (N_2852,In_480,In_1608);
or U2853 (N_2853,In_694,In_415);
nor U2854 (N_2854,In_298,In_1640);
or U2855 (N_2855,In_697,In_1454);
nor U2856 (N_2856,In_161,In_1690);
nor U2857 (N_2857,In_1463,In_906);
nand U2858 (N_2858,In_1869,In_679);
xnor U2859 (N_2859,In_4,In_1620);
or U2860 (N_2860,In_1089,In_871);
nand U2861 (N_2861,In_1355,In_1964);
nor U2862 (N_2862,In_1238,In_416);
or U2863 (N_2863,In_1013,In_1475);
or U2864 (N_2864,In_1753,In_1781);
or U2865 (N_2865,In_497,In_926);
nor U2866 (N_2866,In_1530,In_1050);
nor U2867 (N_2867,In_121,In_1839);
nor U2868 (N_2868,In_1502,In_1907);
or U2869 (N_2869,In_1147,In_29);
nand U2870 (N_2870,In_673,In_402);
or U2871 (N_2871,In_240,In_792);
nand U2872 (N_2872,In_1517,In_1010);
and U2873 (N_2873,In_1663,In_12);
and U2874 (N_2874,In_1145,In_349);
or U2875 (N_2875,In_876,In_1226);
nand U2876 (N_2876,In_1661,In_274);
nand U2877 (N_2877,In_1413,In_1820);
and U2878 (N_2878,In_1365,In_1284);
or U2879 (N_2879,In_1401,In_192);
or U2880 (N_2880,In_461,In_1378);
and U2881 (N_2881,In_76,In_1308);
xor U2882 (N_2882,In_1279,In_621);
or U2883 (N_2883,In_64,In_1242);
or U2884 (N_2884,In_1240,In_648);
or U2885 (N_2885,In_89,In_504);
nand U2886 (N_2886,In_269,In_1624);
or U2887 (N_2887,In_254,In_66);
nand U2888 (N_2888,In_320,In_1588);
nand U2889 (N_2889,In_946,In_1513);
and U2890 (N_2890,In_1729,In_398);
nor U2891 (N_2891,In_678,In_1687);
or U2892 (N_2892,In_1734,In_757);
nand U2893 (N_2893,In_1808,In_891);
or U2894 (N_2894,In_473,In_867);
or U2895 (N_2895,In_1937,In_705);
nand U2896 (N_2896,In_513,In_205);
and U2897 (N_2897,In_456,In_219);
or U2898 (N_2898,In_1883,In_1307);
or U2899 (N_2899,In_1799,In_1659);
or U2900 (N_2900,In_894,In_1697);
or U2901 (N_2901,In_786,In_1486);
xnor U2902 (N_2902,In_612,In_1859);
and U2903 (N_2903,In_462,In_1874);
and U2904 (N_2904,In_475,In_1384);
nor U2905 (N_2905,In_744,In_1804);
nand U2906 (N_2906,In_399,In_1964);
or U2907 (N_2907,In_1607,In_684);
and U2908 (N_2908,In_1943,In_1668);
or U2909 (N_2909,In_820,In_1534);
and U2910 (N_2910,In_944,In_1872);
nor U2911 (N_2911,In_1073,In_474);
nor U2912 (N_2912,In_293,In_1013);
nor U2913 (N_2913,In_682,In_966);
xor U2914 (N_2914,In_490,In_1199);
nand U2915 (N_2915,In_1523,In_720);
nand U2916 (N_2916,In_1912,In_1320);
and U2917 (N_2917,In_1401,In_1327);
and U2918 (N_2918,In_1793,In_879);
nor U2919 (N_2919,In_960,In_1053);
nor U2920 (N_2920,In_1191,In_490);
nor U2921 (N_2921,In_1429,In_1826);
nand U2922 (N_2922,In_1329,In_1780);
nand U2923 (N_2923,In_254,In_233);
and U2924 (N_2924,In_1927,In_180);
nand U2925 (N_2925,In_347,In_1846);
and U2926 (N_2926,In_1491,In_1434);
or U2927 (N_2927,In_67,In_308);
or U2928 (N_2928,In_462,In_1692);
or U2929 (N_2929,In_1638,In_1894);
or U2930 (N_2930,In_773,In_140);
nor U2931 (N_2931,In_714,In_1413);
nand U2932 (N_2932,In_825,In_1520);
nand U2933 (N_2933,In_578,In_1446);
or U2934 (N_2934,In_1299,In_1497);
or U2935 (N_2935,In_1708,In_1930);
and U2936 (N_2936,In_139,In_576);
and U2937 (N_2937,In_362,In_1033);
and U2938 (N_2938,In_142,In_98);
and U2939 (N_2939,In_1685,In_215);
or U2940 (N_2940,In_840,In_200);
xnor U2941 (N_2941,In_1428,In_1012);
nand U2942 (N_2942,In_1124,In_569);
nand U2943 (N_2943,In_1073,In_1652);
and U2944 (N_2944,In_586,In_1771);
and U2945 (N_2945,In_382,In_1358);
and U2946 (N_2946,In_770,In_419);
nand U2947 (N_2947,In_1819,In_275);
or U2948 (N_2948,In_1068,In_1172);
or U2949 (N_2949,In_1661,In_193);
nor U2950 (N_2950,In_185,In_213);
nor U2951 (N_2951,In_1786,In_646);
nor U2952 (N_2952,In_1765,In_1556);
xnor U2953 (N_2953,In_1564,In_541);
or U2954 (N_2954,In_585,In_1024);
or U2955 (N_2955,In_1593,In_1514);
xor U2956 (N_2956,In_1737,In_1152);
nor U2957 (N_2957,In_125,In_826);
nor U2958 (N_2958,In_276,In_319);
or U2959 (N_2959,In_1086,In_463);
nand U2960 (N_2960,In_670,In_1819);
or U2961 (N_2961,In_578,In_708);
or U2962 (N_2962,In_1074,In_141);
and U2963 (N_2963,In_1419,In_839);
nor U2964 (N_2964,In_254,In_1246);
and U2965 (N_2965,In_344,In_955);
nand U2966 (N_2966,In_130,In_1719);
xor U2967 (N_2967,In_1897,In_1587);
nand U2968 (N_2968,In_1387,In_50);
xor U2969 (N_2969,In_729,In_1593);
xor U2970 (N_2970,In_1078,In_1108);
or U2971 (N_2971,In_821,In_759);
nand U2972 (N_2972,In_978,In_145);
nand U2973 (N_2973,In_359,In_123);
nor U2974 (N_2974,In_1983,In_984);
and U2975 (N_2975,In_1680,In_512);
nor U2976 (N_2976,In_1921,In_1525);
nand U2977 (N_2977,In_1772,In_1982);
or U2978 (N_2978,In_293,In_1652);
or U2979 (N_2979,In_32,In_29);
and U2980 (N_2980,In_1615,In_295);
xor U2981 (N_2981,In_877,In_539);
or U2982 (N_2982,In_1657,In_1414);
and U2983 (N_2983,In_1785,In_348);
or U2984 (N_2984,In_802,In_1869);
xor U2985 (N_2985,In_1382,In_980);
nand U2986 (N_2986,In_334,In_1359);
or U2987 (N_2987,In_1689,In_241);
nand U2988 (N_2988,In_52,In_213);
xor U2989 (N_2989,In_756,In_944);
nor U2990 (N_2990,In_916,In_1877);
nor U2991 (N_2991,In_1254,In_997);
nor U2992 (N_2992,In_1172,In_501);
nor U2993 (N_2993,In_1849,In_1334);
or U2994 (N_2994,In_1585,In_211);
or U2995 (N_2995,In_1985,In_38);
nor U2996 (N_2996,In_1010,In_363);
nor U2997 (N_2997,In_231,In_1215);
xor U2998 (N_2998,In_1539,In_430);
and U2999 (N_2999,In_1143,In_1969);
and U3000 (N_3000,In_192,In_582);
or U3001 (N_3001,In_970,In_1561);
nand U3002 (N_3002,In_741,In_1448);
nand U3003 (N_3003,In_705,In_912);
or U3004 (N_3004,In_1452,In_1697);
nand U3005 (N_3005,In_490,In_216);
and U3006 (N_3006,In_1330,In_507);
nand U3007 (N_3007,In_1870,In_460);
nor U3008 (N_3008,In_163,In_1800);
and U3009 (N_3009,In_888,In_871);
or U3010 (N_3010,In_336,In_317);
or U3011 (N_3011,In_625,In_1631);
nand U3012 (N_3012,In_1376,In_30);
and U3013 (N_3013,In_795,In_1691);
nand U3014 (N_3014,In_538,In_740);
or U3015 (N_3015,In_301,In_151);
nand U3016 (N_3016,In_753,In_1163);
and U3017 (N_3017,In_1739,In_1385);
xnor U3018 (N_3018,In_1368,In_465);
and U3019 (N_3019,In_45,In_1403);
nand U3020 (N_3020,In_124,In_1849);
or U3021 (N_3021,In_747,In_1939);
and U3022 (N_3022,In_1323,In_573);
xnor U3023 (N_3023,In_1815,In_104);
and U3024 (N_3024,In_1546,In_1376);
and U3025 (N_3025,In_1365,In_1340);
xnor U3026 (N_3026,In_835,In_1659);
nor U3027 (N_3027,In_576,In_1328);
and U3028 (N_3028,In_416,In_1544);
and U3029 (N_3029,In_1532,In_1520);
nor U3030 (N_3030,In_969,In_1091);
nand U3031 (N_3031,In_482,In_721);
nand U3032 (N_3032,In_1269,In_1475);
or U3033 (N_3033,In_344,In_1140);
and U3034 (N_3034,In_1856,In_1314);
or U3035 (N_3035,In_704,In_729);
and U3036 (N_3036,In_201,In_1647);
nor U3037 (N_3037,In_787,In_558);
and U3038 (N_3038,In_1669,In_1118);
or U3039 (N_3039,In_1643,In_819);
nor U3040 (N_3040,In_101,In_365);
or U3041 (N_3041,In_355,In_1944);
nand U3042 (N_3042,In_5,In_83);
nor U3043 (N_3043,In_815,In_1676);
nor U3044 (N_3044,In_956,In_1744);
or U3045 (N_3045,In_1742,In_1738);
and U3046 (N_3046,In_1400,In_1742);
and U3047 (N_3047,In_793,In_1968);
or U3048 (N_3048,In_1067,In_5);
or U3049 (N_3049,In_67,In_618);
or U3050 (N_3050,In_206,In_1728);
or U3051 (N_3051,In_74,In_653);
and U3052 (N_3052,In_1008,In_153);
or U3053 (N_3053,In_938,In_671);
nor U3054 (N_3054,In_472,In_712);
or U3055 (N_3055,In_1391,In_380);
nor U3056 (N_3056,In_178,In_1152);
nand U3057 (N_3057,In_1867,In_1912);
xnor U3058 (N_3058,In_1950,In_1448);
nor U3059 (N_3059,In_1443,In_1530);
nand U3060 (N_3060,In_253,In_702);
nand U3061 (N_3061,In_1993,In_1013);
or U3062 (N_3062,In_453,In_1465);
or U3063 (N_3063,In_1743,In_1527);
nand U3064 (N_3064,In_880,In_924);
or U3065 (N_3065,In_1810,In_194);
xnor U3066 (N_3066,In_511,In_1670);
or U3067 (N_3067,In_1764,In_325);
nor U3068 (N_3068,In_1407,In_946);
or U3069 (N_3069,In_746,In_1682);
and U3070 (N_3070,In_1271,In_85);
nand U3071 (N_3071,In_173,In_854);
xnor U3072 (N_3072,In_780,In_658);
nor U3073 (N_3073,In_496,In_1980);
or U3074 (N_3074,In_125,In_767);
xor U3075 (N_3075,In_501,In_1096);
or U3076 (N_3076,In_1274,In_1107);
and U3077 (N_3077,In_1518,In_1339);
or U3078 (N_3078,In_306,In_1058);
and U3079 (N_3079,In_1330,In_695);
or U3080 (N_3080,In_592,In_66);
and U3081 (N_3081,In_525,In_207);
and U3082 (N_3082,In_491,In_1921);
nand U3083 (N_3083,In_1533,In_1283);
or U3084 (N_3084,In_1669,In_1687);
nor U3085 (N_3085,In_400,In_1925);
or U3086 (N_3086,In_390,In_890);
or U3087 (N_3087,In_824,In_306);
nor U3088 (N_3088,In_1073,In_685);
and U3089 (N_3089,In_551,In_1493);
nand U3090 (N_3090,In_1788,In_1366);
xnor U3091 (N_3091,In_45,In_983);
nor U3092 (N_3092,In_1817,In_1561);
xnor U3093 (N_3093,In_1217,In_932);
nor U3094 (N_3094,In_1177,In_949);
or U3095 (N_3095,In_167,In_490);
or U3096 (N_3096,In_80,In_917);
or U3097 (N_3097,In_1038,In_402);
and U3098 (N_3098,In_738,In_1680);
nor U3099 (N_3099,In_1428,In_880);
nor U3100 (N_3100,In_1220,In_745);
nor U3101 (N_3101,In_1768,In_965);
and U3102 (N_3102,In_1775,In_1868);
nor U3103 (N_3103,In_236,In_1626);
nand U3104 (N_3104,In_1881,In_805);
and U3105 (N_3105,In_226,In_316);
nor U3106 (N_3106,In_1496,In_560);
nor U3107 (N_3107,In_1738,In_823);
nor U3108 (N_3108,In_922,In_287);
or U3109 (N_3109,In_1733,In_1848);
or U3110 (N_3110,In_1636,In_351);
nor U3111 (N_3111,In_613,In_1224);
and U3112 (N_3112,In_1154,In_1356);
nor U3113 (N_3113,In_143,In_657);
or U3114 (N_3114,In_116,In_1063);
or U3115 (N_3115,In_181,In_1078);
nor U3116 (N_3116,In_161,In_464);
nand U3117 (N_3117,In_1134,In_1349);
or U3118 (N_3118,In_895,In_1977);
nor U3119 (N_3119,In_730,In_1123);
and U3120 (N_3120,In_1099,In_294);
nand U3121 (N_3121,In_1234,In_846);
nor U3122 (N_3122,In_1025,In_1450);
or U3123 (N_3123,In_1304,In_1297);
or U3124 (N_3124,In_1516,In_1768);
nor U3125 (N_3125,In_1030,In_1119);
xor U3126 (N_3126,In_550,In_308);
and U3127 (N_3127,In_444,In_1378);
and U3128 (N_3128,In_1804,In_354);
or U3129 (N_3129,In_249,In_1268);
and U3130 (N_3130,In_854,In_478);
nor U3131 (N_3131,In_846,In_1562);
xor U3132 (N_3132,In_640,In_602);
nand U3133 (N_3133,In_1165,In_708);
or U3134 (N_3134,In_1280,In_115);
and U3135 (N_3135,In_1749,In_838);
nor U3136 (N_3136,In_31,In_1901);
nor U3137 (N_3137,In_842,In_1145);
nor U3138 (N_3138,In_146,In_1146);
and U3139 (N_3139,In_1500,In_1895);
or U3140 (N_3140,In_564,In_589);
nand U3141 (N_3141,In_1367,In_1531);
and U3142 (N_3142,In_1857,In_1821);
and U3143 (N_3143,In_1955,In_294);
nand U3144 (N_3144,In_433,In_1859);
xor U3145 (N_3145,In_201,In_285);
and U3146 (N_3146,In_949,In_1920);
or U3147 (N_3147,In_407,In_1361);
or U3148 (N_3148,In_393,In_682);
nor U3149 (N_3149,In_329,In_1434);
nor U3150 (N_3150,In_1085,In_1788);
or U3151 (N_3151,In_1420,In_342);
nor U3152 (N_3152,In_665,In_1917);
xnor U3153 (N_3153,In_962,In_972);
nor U3154 (N_3154,In_278,In_1731);
nor U3155 (N_3155,In_75,In_1178);
nor U3156 (N_3156,In_1270,In_1063);
nand U3157 (N_3157,In_1434,In_1849);
nor U3158 (N_3158,In_1477,In_303);
nor U3159 (N_3159,In_436,In_1680);
and U3160 (N_3160,In_20,In_1862);
nand U3161 (N_3161,In_314,In_820);
xnor U3162 (N_3162,In_746,In_1713);
and U3163 (N_3163,In_656,In_482);
and U3164 (N_3164,In_904,In_980);
or U3165 (N_3165,In_1229,In_550);
xnor U3166 (N_3166,In_159,In_1488);
nand U3167 (N_3167,In_57,In_1332);
or U3168 (N_3168,In_1113,In_513);
or U3169 (N_3169,In_1905,In_1154);
nor U3170 (N_3170,In_1402,In_296);
or U3171 (N_3171,In_372,In_1026);
nand U3172 (N_3172,In_30,In_95);
or U3173 (N_3173,In_583,In_543);
nor U3174 (N_3174,In_564,In_1606);
nor U3175 (N_3175,In_328,In_869);
xnor U3176 (N_3176,In_1735,In_655);
nor U3177 (N_3177,In_1817,In_1074);
or U3178 (N_3178,In_1846,In_126);
nor U3179 (N_3179,In_431,In_377);
nor U3180 (N_3180,In_1267,In_1777);
and U3181 (N_3181,In_1042,In_1353);
nand U3182 (N_3182,In_953,In_836);
and U3183 (N_3183,In_536,In_280);
xor U3184 (N_3184,In_1045,In_1664);
nand U3185 (N_3185,In_218,In_549);
xnor U3186 (N_3186,In_1430,In_1472);
nor U3187 (N_3187,In_775,In_1642);
and U3188 (N_3188,In_674,In_1398);
or U3189 (N_3189,In_1612,In_1092);
and U3190 (N_3190,In_638,In_1909);
and U3191 (N_3191,In_874,In_1243);
or U3192 (N_3192,In_1554,In_114);
or U3193 (N_3193,In_289,In_930);
or U3194 (N_3194,In_1819,In_35);
or U3195 (N_3195,In_221,In_1352);
and U3196 (N_3196,In_1428,In_1620);
and U3197 (N_3197,In_799,In_1490);
or U3198 (N_3198,In_1691,In_689);
nand U3199 (N_3199,In_435,In_1579);
and U3200 (N_3200,In_584,In_1371);
and U3201 (N_3201,In_1255,In_1887);
nor U3202 (N_3202,In_423,In_562);
or U3203 (N_3203,In_240,In_1187);
xor U3204 (N_3204,In_1726,In_1783);
nand U3205 (N_3205,In_179,In_1665);
or U3206 (N_3206,In_1210,In_766);
xor U3207 (N_3207,In_1662,In_1854);
or U3208 (N_3208,In_1091,In_415);
nand U3209 (N_3209,In_1232,In_1202);
or U3210 (N_3210,In_387,In_1600);
nor U3211 (N_3211,In_1345,In_1565);
nor U3212 (N_3212,In_997,In_329);
nor U3213 (N_3213,In_564,In_1509);
nand U3214 (N_3214,In_1448,In_288);
or U3215 (N_3215,In_1489,In_1485);
xor U3216 (N_3216,In_1778,In_1823);
nand U3217 (N_3217,In_1948,In_1778);
nor U3218 (N_3218,In_957,In_638);
nand U3219 (N_3219,In_1749,In_1696);
nand U3220 (N_3220,In_1114,In_1848);
nand U3221 (N_3221,In_839,In_964);
or U3222 (N_3222,In_768,In_1176);
nor U3223 (N_3223,In_901,In_1975);
nand U3224 (N_3224,In_775,In_814);
nand U3225 (N_3225,In_495,In_852);
or U3226 (N_3226,In_1345,In_1982);
or U3227 (N_3227,In_116,In_159);
xor U3228 (N_3228,In_192,In_1174);
and U3229 (N_3229,In_886,In_1904);
or U3230 (N_3230,In_994,In_43);
or U3231 (N_3231,In_127,In_573);
or U3232 (N_3232,In_1723,In_843);
nand U3233 (N_3233,In_1320,In_1974);
and U3234 (N_3234,In_767,In_946);
and U3235 (N_3235,In_1754,In_656);
or U3236 (N_3236,In_414,In_1548);
or U3237 (N_3237,In_1242,In_1616);
nor U3238 (N_3238,In_1811,In_1163);
xnor U3239 (N_3239,In_983,In_906);
nand U3240 (N_3240,In_479,In_23);
or U3241 (N_3241,In_1503,In_506);
nand U3242 (N_3242,In_122,In_1042);
or U3243 (N_3243,In_1417,In_74);
nand U3244 (N_3244,In_1338,In_300);
nor U3245 (N_3245,In_701,In_486);
nand U3246 (N_3246,In_757,In_1878);
nor U3247 (N_3247,In_1735,In_432);
nand U3248 (N_3248,In_1446,In_1690);
and U3249 (N_3249,In_638,In_1627);
nor U3250 (N_3250,In_1106,In_1669);
nand U3251 (N_3251,In_113,In_1097);
and U3252 (N_3252,In_1153,In_653);
nor U3253 (N_3253,In_1839,In_1663);
nor U3254 (N_3254,In_327,In_766);
nand U3255 (N_3255,In_1635,In_1815);
xnor U3256 (N_3256,In_1163,In_537);
nor U3257 (N_3257,In_782,In_1760);
or U3258 (N_3258,In_1913,In_737);
and U3259 (N_3259,In_1638,In_1477);
or U3260 (N_3260,In_1888,In_1585);
nand U3261 (N_3261,In_833,In_1512);
nor U3262 (N_3262,In_168,In_60);
nand U3263 (N_3263,In_553,In_1565);
and U3264 (N_3264,In_1645,In_1487);
nor U3265 (N_3265,In_1022,In_47);
or U3266 (N_3266,In_1705,In_962);
nor U3267 (N_3267,In_1963,In_893);
and U3268 (N_3268,In_225,In_1018);
and U3269 (N_3269,In_1660,In_903);
nand U3270 (N_3270,In_853,In_806);
or U3271 (N_3271,In_559,In_1642);
or U3272 (N_3272,In_815,In_730);
and U3273 (N_3273,In_762,In_1753);
xor U3274 (N_3274,In_994,In_307);
or U3275 (N_3275,In_1608,In_1793);
nand U3276 (N_3276,In_1041,In_181);
or U3277 (N_3277,In_805,In_929);
nor U3278 (N_3278,In_1369,In_1676);
nor U3279 (N_3279,In_1456,In_1119);
and U3280 (N_3280,In_1532,In_220);
nand U3281 (N_3281,In_309,In_69);
and U3282 (N_3282,In_1722,In_1281);
nor U3283 (N_3283,In_812,In_1335);
or U3284 (N_3284,In_273,In_372);
nor U3285 (N_3285,In_717,In_220);
xor U3286 (N_3286,In_1166,In_251);
or U3287 (N_3287,In_1063,In_1730);
or U3288 (N_3288,In_39,In_1156);
and U3289 (N_3289,In_1965,In_988);
or U3290 (N_3290,In_508,In_1236);
nand U3291 (N_3291,In_335,In_1540);
xnor U3292 (N_3292,In_408,In_371);
nor U3293 (N_3293,In_1370,In_962);
and U3294 (N_3294,In_1347,In_1629);
and U3295 (N_3295,In_111,In_1218);
nand U3296 (N_3296,In_860,In_196);
nand U3297 (N_3297,In_714,In_915);
and U3298 (N_3298,In_1103,In_968);
or U3299 (N_3299,In_1093,In_251);
nor U3300 (N_3300,In_947,In_1504);
nor U3301 (N_3301,In_53,In_1569);
nand U3302 (N_3302,In_1925,In_172);
nor U3303 (N_3303,In_188,In_1658);
or U3304 (N_3304,In_1278,In_596);
nor U3305 (N_3305,In_89,In_983);
or U3306 (N_3306,In_75,In_1839);
and U3307 (N_3307,In_1234,In_1922);
and U3308 (N_3308,In_1666,In_1854);
nor U3309 (N_3309,In_930,In_872);
nand U3310 (N_3310,In_10,In_1125);
nand U3311 (N_3311,In_1180,In_1832);
nor U3312 (N_3312,In_1661,In_1204);
and U3313 (N_3313,In_914,In_72);
xnor U3314 (N_3314,In_239,In_1711);
or U3315 (N_3315,In_574,In_1861);
and U3316 (N_3316,In_468,In_1149);
nor U3317 (N_3317,In_184,In_1700);
nand U3318 (N_3318,In_422,In_343);
and U3319 (N_3319,In_1049,In_405);
nand U3320 (N_3320,In_1866,In_666);
nand U3321 (N_3321,In_1163,In_1745);
nor U3322 (N_3322,In_1014,In_1467);
or U3323 (N_3323,In_1197,In_810);
or U3324 (N_3324,In_1650,In_153);
nor U3325 (N_3325,In_1677,In_582);
nor U3326 (N_3326,In_1990,In_1585);
nand U3327 (N_3327,In_1405,In_987);
or U3328 (N_3328,In_169,In_916);
nand U3329 (N_3329,In_1855,In_87);
xor U3330 (N_3330,In_1751,In_1042);
and U3331 (N_3331,In_625,In_1318);
or U3332 (N_3332,In_1727,In_1176);
and U3333 (N_3333,In_659,In_1459);
or U3334 (N_3334,In_113,In_1672);
nand U3335 (N_3335,In_193,In_580);
or U3336 (N_3336,In_1895,In_1657);
nand U3337 (N_3337,In_1613,In_488);
or U3338 (N_3338,In_1068,In_297);
nor U3339 (N_3339,In_950,In_1844);
or U3340 (N_3340,In_1740,In_272);
nor U3341 (N_3341,In_1314,In_1360);
or U3342 (N_3342,In_1730,In_774);
nor U3343 (N_3343,In_535,In_1161);
nand U3344 (N_3344,In_1700,In_598);
nand U3345 (N_3345,In_779,In_301);
nand U3346 (N_3346,In_1729,In_1314);
and U3347 (N_3347,In_1562,In_1015);
nor U3348 (N_3348,In_64,In_29);
and U3349 (N_3349,In_41,In_488);
or U3350 (N_3350,In_449,In_943);
or U3351 (N_3351,In_381,In_492);
and U3352 (N_3352,In_962,In_1830);
nor U3353 (N_3353,In_1036,In_882);
or U3354 (N_3354,In_771,In_71);
nor U3355 (N_3355,In_896,In_1261);
or U3356 (N_3356,In_357,In_1642);
or U3357 (N_3357,In_1454,In_474);
nand U3358 (N_3358,In_1360,In_1619);
and U3359 (N_3359,In_1489,In_221);
or U3360 (N_3360,In_1400,In_708);
nor U3361 (N_3361,In_1379,In_1797);
or U3362 (N_3362,In_468,In_585);
nor U3363 (N_3363,In_1886,In_1128);
and U3364 (N_3364,In_589,In_1201);
and U3365 (N_3365,In_48,In_1767);
or U3366 (N_3366,In_1995,In_1053);
and U3367 (N_3367,In_1887,In_1902);
nor U3368 (N_3368,In_805,In_1697);
nor U3369 (N_3369,In_1494,In_708);
and U3370 (N_3370,In_91,In_845);
nor U3371 (N_3371,In_1714,In_716);
and U3372 (N_3372,In_1959,In_173);
and U3373 (N_3373,In_689,In_1110);
and U3374 (N_3374,In_1928,In_1909);
and U3375 (N_3375,In_705,In_1722);
nor U3376 (N_3376,In_1629,In_749);
nor U3377 (N_3377,In_701,In_1122);
and U3378 (N_3378,In_436,In_1618);
and U3379 (N_3379,In_535,In_420);
nor U3380 (N_3380,In_205,In_40);
or U3381 (N_3381,In_444,In_604);
or U3382 (N_3382,In_1641,In_514);
xnor U3383 (N_3383,In_726,In_322);
nor U3384 (N_3384,In_633,In_1515);
or U3385 (N_3385,In_1498,In_936);
and U3386 (N_3386,In_345,In_1979);
xnor U3387 (N_3387,In_1287,In_1681);
nand U3388 (N_3388,In_1036,In_1510);
nand U3389 (N_3389,In_152,In_731);
xor U3390 (N_3390,In_1983,In_734);
or U3391 (N_3391,In_444,In_1424);
or U3392 (N_3392,In_1131,In_1529);
nor U3393 (N_3393,In_1522,In_131);
nand U3394 (N_3394,In_352,In_1798);
nor U3395 (N_3395,In_42,In_1033);
nand U3396 (N_3396,In_473,In_504);
or U3397 (N_3397,In_1618,In_1018);
nand U3398 (N_3398,In_1504,In_1436);
or U3399 (N_3399,In_149,In_818);
nor U3400 (N_3400,In_1121,In_369);
and U3401 (N_3401,In_879,In_536);
nand U3402 (N_3402,In_1737,In_650);
and U3403 (N_3403,In_1329,In_1711);
and U3404 (N_3404,In_1219,In_1988);
or U3405 (N_3405,In_42,In_927);
nor U3406 (N_3406,In_482,In_789);
or U3407 (N_3407,In_1438,In_1025);
and U3408 (N_3408,In_1455,In_114);
nor U3409 (N_3409,In_470,In_1090);
nor U3410 (N_3410,In_1723,In_263);
nand U3411 (N_3411,In_1174,In_19);
nor U3412 (N_3412,In_397,In_148);
or U3413 (N_3413,In_1209,In_73);
nor U3414 (N_3414,In_351,In_1038);
nand U3415 (N_3415,In_1581,In_1607);
or U3416 (N_3416,In_1053,In_326);
and U3417 (N_3417,In_1688,In_617);
nor U3418 (N_3418,In_758,In_488);
or U3419 (N_3419,In_897,In_1905);
and U3420 (N_3420,In_1667,In_572);
nor U3421 (N_3421,In_1494,In_1365);
xnor U3422 (N_3422,In_930,In_1048);
nand U3423 (N_3423,In_1408,In_60);
nand U3424 (N_3424,In_1890,In_1522);
or U3425 (N_3425,In_1150,In_1951);
nand U3426 (N_3426,In_285,In_1872);
nand U3427 (N_3427,In_531,In_1939);
nand U3428 (N_3428,In_570,In_438);
nor U3429 (N_3429,In_1156,In_1039);
nor U3430 (N_3430,In_1058,In_27);
xnor U3431 (N_3431,In_1313,In_1216);
nand U3432 (N_3432,In_47,In_1099);
or U3433 (N_3433,In_387,In_1016);
and U3434 (N_3434,In_753,In_321);
nor U3435 (N_3435,In_1196,In_1249);
and U3436 (N_3436,In_1233,In_850);
xnor U3437 (N_3437,In_881,In_1871);
or U3438 (N_3438,In_1205,In_1196);
xnor U3439 (N_3439,In_1159,In_1022);
or U3440 (N_3440,In_1349,In_1287);
nand U3441 (N_3441,In_864,In_1949);
and U3442 (N_3442,In_1995,In_1642);
or U3443 (N_3443,In_329,In_482);
or U3444 (N_3444,In_1362,In_1951);
or U3445 (N_3445,In_1067,In_1435);
nor U3446 (N_3446,In_1422,In_1818);
and U3447 (N_3447,In_376,In_568);
and U3448 (N_3448,In_1725,In_1928);
or U3449 (N_3449,In_861,In_791);
nor U3450 (N_3450,In_1802,In_1792);
nand U3451 (N_3451,In_1664,In_86);
nor U3452 (N_3452,In_1216,In_1041);
and U3453 (N_3453,In_1052,In_1732);
or U3454 (N_3454,In_1215,In_1196);
nand U3455 (N_3455,In_592,In_348);
nor U3456 (N_3456,In_1860,In_1437);
and U3457 (N_3457,In_43,In_1919);
and U3458 (N_3458,In_1570,In_1448);
or U3459 (N_3459,In_205,In_1006);
xnor U3460 (N_3460,In_115,In_757);
xnor U3461 (N_3461,In_1315,In_1805);
nor U3462 (N_3462,In_191,In_1936);
nor U3463 (N_3463,In_884,In_1280);
nor U3464 (N_3464,In_1975,In_1339);
and U3465 (N_3465,In_505,In_57);
nand U3466 (N_3466,In_863,In_1919);
nor U3467 (N_3467,In_1208,In_1693);
xor U3468 (N_3468,In_34,In_1928);
nand U3469 (N_3469,In_335,In_995);
xnor U3470 (N_3470,In_1173,In_1654);
or U3471 (N_3471,In_970,In_358);
nand U3472 (N_3472,In_1871,In_116);
or U3473 (N_3473,In_1992,In_286);
or U3474 (N_3474,In_331,In_752);
or U3475 (N_3475,In_1206,In_949);
nor U3476 (N_3476,In_1719,In_1133);
or U3477 (N_3477,In_416,In_1090);
nor U3478 (N_3478,In_238,In_1994);
or U3479 (N_3479,In_183,In_1818);
and U3480 (N_3480,In_546,In_1623);
nand U3481 (N_3481,In_1157,In_726);
nand U3482 (N_3482,In_714,In_1555);
nand U3483 (N_3483,In_1084,In_1211);
and U3484 (N_3484,In_1603,In_1775);
xnor U3485 (N_3485,In_969,In_24);
xnor U3486 (N_3486,In_1756,In_1746);
and U3487 (N_3487,In_1966,In_1408);
nor U3488 (N_3488,In_1876,In_1556);
and U3489 (N_3489,In_1789,In_87);
nand U3490 (N_3490,In_1958,In_1858);
nand U3491 (N_3491,In_1712,In_1609);
and U3492 (N_3492,In_246,In_1975);
nor U3493 (N_3493,In_1891,In_1333);
nand U3494 (N_3494,In_1736,In_1398);
or U3495 (N_3495,In_1854,In_1990);
or U3496 (N_3496,In_414,In_377);
or U3497 (N_3497,In_1992,In_1974);
or U3498 (N_3498,In_1716,In_1138);
nand U3499 (N_3499,In_1396,In_1517);
and U3500 (N_3500,In_1973,In_60);
nand U3501 (N_3501,In_1522,In_579);
or U3502 (N_3502,In_1320,In_43);
nand U3503 (N_3503,In_1994,In_1321);
and U3504 (N_3504,In_503,In_643);
and U3505 (N_3505,In_1870,In_1234);
nand U3506 (N_3506,In_991,In_1575);
nor U3507 (N_3507,In_1227,In_328);
nand U3508 (N_3508,In_1843,In_1427);
xnor U3509 (N_3509,In_1014,In_1658);
xnor U3510 (N_3510,In_1340,In_1650);
and U3511 (N_3511,In_1742,In_1252);
nand U3512 (N_3512,In_124,In_1042);
nand U3513 (N_3513,In_648,In_144);
and U3514 (N_3514,In_118,In_1491);
nor U3515 (N_3515,In_1999,In_958);
or U3516 (N_3516,In_1701,In_592);
nand U3517 (N_3517,In_1445,In_1118);
nand U3518 (N_3518,In_703,In_1838);
or U3519 (N_3519,In_1306,In_730);
or U3520 (N_3520,In_1112,In_410);
nand U3521 (N_3521,In_694,In_951);
or U3522 (N_3522,In_1078,In_1844);
xor U3523 (N_3523,In_872,In_247);
or U3524 (N_3524,In_1515,In_59);
nor U3525 (N_3525,In_1342,In_1026);
nor U3526 (N_3526,In_1898,In_756);
or U3527 (N_3527,In_1336,In_748);
xor U3528 (N_3528,In_1872,In_1921);
xor U3529 (N_3529,In_1573,In_1850);
nand U3530 (N_3530,In_268,In_1703);
xnor U3531 (N_3531,In_388,In_481);
nand U3532 (N_3532,In_1787,In_218);
nor U3533 (N_3533,In_191,In_405);
nand U3534 (N_3534,In_1568,In_988);
nor U3535 (N_3535,In_1804,In_1408);
or U3536 (N_3536,In_1802,In_1926);
and U3537 (N_3537,In_359,In_239);
xnor U3538 (N_3538,In_1296,In_854);
nand U3539 (N_3539,In_858,In_503);
or U3540 (N_3540,In_1483,In_567);
and U3541 (N_3541,In_73,In_941);
or U3542 (N_3542,In_1815,In_1978);
nand U3543 (N_3543,In_64,In_467);
nor U3544 (N_3544,In_269,In_755);
and U3545 (N_3545,In_1520,In_1445);
nor U3546 (N_3546,In_1567,In_374);
xor U3547 (N_3547,In_612,In_1829);
or U3548 (N_3548,In_1873,In_770);
nand U3549 (N_3549,In_1882,In_258);
nor U3550 (N_3550,In_1267,In_1205);
and U3551 (N_3551,In_656,In_809);
nor U3552 (N_3552,In_87,In_1626);
nand U3553 (N_3553,In_623,In_1194);
nor U3554 (N_3554,In_1683,In_102);
nor U3555 (N_3555,In_663,In_1948);
and U3556 (N_3556,In_891,In_182);
and U3557 (N_3557,In_1110,In_1132);
and U3558 (N_3558,In_1248,In_232);
xnor U3559 (N_3559,In_1570,In_1767);
and U3560 (N_3560,In_1987,In_172);
and U3561 (N_3561,In_580,In_798);
or U3562 (N_3562,In_52,In_579);
nor U3563 (N_3563,In_1820,In_1951);
or U3564 (N_3564,In_743,In_1795);
nand U3565 (N_3565,In_1721,In_1901);
nand U3566 (N_3566,In_650,In_1067);
nand U3567 (N_3567,In_753,In_9);
nor U3568 (N_3568,In_356,In_1579);
nor U3569 (N_3569,In_914,In_84);
xnor U3570 (N_3570,In_478,In_1870);
nand U3571 (N_3571,In_1497,In_1196);
nor U3572 (N_3572,In_1458,In_1607);
nor U3573 (N_3573,In_1388,In_1186);
nor U3574 (N_3574,In_1508,In_718);
or U3575 (N_3575,In_1979,In_893);
xnor U3576 (N_3576,In_180,In_1913);
and U3577 (N_3577,In_264,In_505);
nor U3578 (N_3578,In_1053,In_1893);
or U3579 (N_3579,In_437,In_136);
nor U3580 (N_3580,In_22,In_778);
nor U3581 (N_3581,In_1035,In_1005);
xnor U3582 (N_3582,In_855,In_1841);
nor U3583 (N_3583,In_805,In_925);
nand U3584 (N_3584,In_767,In_1503);
xor U3585 (N_3585,In_1641,In_304);
xor U3586 (N_3586,In_1159,In_1459);
nand U3587 (N_3587,In_851,In_1131);
nand U3588 (N_3588,In_1859,In_1290);
xor U3589 (N_3589,In_47,In_28);
and U3590 (N_3590,In_432,In_1026);
nand U3591 (N_3591,In_361,In_1506);
nand U3592 (N_3592,In_1472,In_1677);
nand U3593 (N_3593,In_1241,In_960);
nand U3594 (N_3594,In_1405,In_80);
or U3595 (N_3595,In_836,In_197);
and U3596 (N_3596,In_899,In_795);
nand U3597 (N_3597,In_1884,In_1768);
and U3598 (N_3598,In_290,In_712);
nand U3599 (N_3599,In_1347,In_883);
nor U3600 (N_3600,In_85,In_669);
nand U3601 (N_3601,In_200,In_696);
and U3602 (N_3602,In_1064,In_1583);
nor U3603 (N_3603,In_440,In_1823);
and U3604 (N_3604,In_244,In_1511);
and U3605 (N_3605,In_1933,In_760);
or U3606 (N_3606,In_911,In_693);
nand U3607 (N_3607,In_281,In_82);
nor U3608 (N_3608,In_1891,In_1366);
nor U3609 (N_3609,In_1828,In_1163);
nand U3610 (N_3610,In_1429,In_916);
or U3611 (N_3611,In_757,In_686);
or U3612 (N_3612,In_534,In_434);
and U3613 (N_3613,In_536,In_704);
and U3614 (N_3614,In_1893,In_718);
nand U3615 (N_3615,In_695,In_953);
nand U3616 (N_3616,In_1519,In_355);
nand U3617 (N_3617,In_1928,In_214);
or U3618 (N_3618,In_588,In_1641);
or U3619 (N_3619,In_921,In_895);
or U3620 (N_3620,In_779,In_1157);
and U3621 (N_3621,In_239,In_1852);
xor U3622 (N_3622,In_1367,In_1172);
or U3623 (N_3623,In_300,In_814);
nor U3624 (N_3624,In_1125,In_774);
or U3625 (N_3625,In_1778,In_322);
or U3626 (N_3626,In_342,In_1459);
and U3627 (N_3627,In_1700,In_1110);
xor U3628 (N_3628,In_1041,In_1695);
or U3629 (N_3629,In_1569,In_674);
nand U3630 (N_3630,In_32,In_1451);
nand U3631 (N_3631,In_699,In_1832);
nor U3632 (N_3632,In_1191,In_382);
nor U3633 (N_3633,In_137,In_626);
xnor U3634 (N_3634,In_1917,In_1761);
and U3635 (N_3635,In_1046,In_1715);
or U3636 (N_3636,In_1050,In_1742);
nand U3637 (N_3637,In_1974,In_1335);
and U3638 (N_3638,In_1641,In_1130);
and U3639 (N_3639,In_950,In_1450);
nor U3640 (N_3640,In_595,In_96);
and U3641 (N_3641,In_1878,In_1491);
nor U3642 (N_3642,In_341,In_632);
nand U3643 (N_3643,In_1258,In_796);
nor U3644 (N_3644,In_1610,In_444);
xnor U3645 (N_3645,In_1027,In_37);
nand U3646 (N_3646,In_1277,In_1727);
and U3647 (N_3647,In_708,In_640);
nand U3648 (N_3648,In_270,In_1478);
xor U3649 (N_3649,In_1833,In_1208);
nor U3650 (N_3650,In_108,In_1062);
xor U3651 (N_3651,In_1612,In_651);
nor U3652 (N_3652,In_807,In_467);
or U3653 (N_3653,In_1444,In_1699);
nor U3654 (N_3654,In_608,In_669);
and U3655 (N_3655,In_1108,In_565);
and U3656 (N_3656,In_164,In_627);
or U3657 (N_3657,In_1344,In_912);
and U3658 (N_3658,In_760,In_1635);
and U3659 (N_3659,In_1843,In_1957);
and U3660 (N_3660,In_305,In_1866);
nor U3661 (N_3661,In_1159,In_65);
nor U3662 (N_3662,In_1934,In_789);
and U3663 (N_3663,In_1156,In_1096);
or U3664 (N_3664,In_26,In_540);
and U3665 (N_3665,In_542,In_1011);
and U3666 (N_3666,In_317,In_1504);
nand U3667 (N_3667,In_522,In_1023);
nand U3668 (N_3668,In_816,In_260);
xnor U3669 (N_3669,In_1481,In_1831);
and U3670 (N_3670,In_414,In_1802);
and U3671 (N_3671,In_894,In_370);
xor U3672 (N_3672,In_1418,In_1720);
or U3673 (N_3673,In_707,In_1139);
nor U3674 (N_3674,In_1078,In_1319);
and U3675 (N_3675,In_606,In_362);
or U3676 (N_3676,In_1887,In_1096);
and U3677 (N_3677,In_1804,In_326);
nand U3678 (N_3678,In_824,In_1483);
nor U3679 (N_3679,In_1553,In_309);
or U3680 (N_3680,In_423,In_613);
and U3681 (N_3681,In_516,In_638);
xor U3682 (N_3682,In_157,In_1952);
nand U3683 (N_3683,In_1409,In_947);
nor U3684 (N_3684,In_1594,In_466);
or U3685 (N_3685,In_1164,In_649);
nand U3686 (N_3686,In_1003,In_235);
nor U3687 (N_3687,In_1535,In_794);
nor U3688 (N_3688,In_441,In_957);
or U3689 (N_3689,In_831,In_1043);
or U3690 (N_3690,In_444,In_1503);
xnor U3691 (N_3691,In_483,In_277);
nor U3692 (N_3692,In_144,In_1030);
nor U3693 (N_3693,In_385,In_607);
and U3694 (N_3694,In_1631,In_1488);
nor U3695 (N_3695,In_874,In_356);
and U3696 (N_3696,In_1271,In_1070);
nor U3697 (N_3697,In_765,In_722);
or U3698 (N_3698,In_1597,In_1790);
xnor U3699 (N_3699,In_894,In_618);
or U3700 (N_3700,In_681,In_1381);
or U3701 (N_3701,In_1641,In_1085);
xnor U3702 (N_3702,In_788,In_83);
xnor U3703 (N_3703,In_1649,In_903);
nand U3704 (N_3704,In_873,In_1807);
and U3705 (N_3705,In_783,In_1450);
xor U3706 (N_3706,In_1548,In_59);
or U3707 (N_3707,In_1810,In_1582);
and U3708 (N_3708,In_641,In_1041);
and U3709 (N_3709,In_1316,In_712);
nor U3710 (N_3710,In_719,In_701);
and U3711 (N_3711,In_1220,In_679);
or U3712 (N_3712,In_1710,In_1887);
and U3713 (N_3713,In_0,In_1857);
and U3714 (N_3714,In_626,In_557);
nand U3715 (N_3715,In_175,In_851);
and U3716 (N_3716,In_1854,In_205);
nor U3717 (N_3717,In_1308,In_1339);
or U3718 (N_3718,In_487,In_427);
and U3719 (N_3719,In_655,In_1359);
and U3720 (N_3720,In_1905,In_1570);
xor U3721 (N_3721,In_1680,In_1502);
nand U3722 (N_3722,In_1099,In_1347);
or U3723 (N_3723,In_1832,In_1269);
xnor U3724 (N_3724,In_788,In_1443);
nand U3725 (N_3725,In_430,In_1187);
and U3726 (N_3726,In_1295,In_217);
nor U3727 (N_3727,In_1212,In_746);
nor U3728 (N_3728,In_28,In_677);
and U3729 (N_3729,In_1567,In_252);
or U3730 (N_3730,In_954,In_1665);
nor U3731 (N_3731,In_1414,In_1326);
nor U3732 (N_3732,In_1390,In_1201);
nor U3733 (N_3733,In_1478,In_947);
nor U3734 (N_3734,In_723,In_778);
or U3735 (N_3735,In_1547,In_1841);
nor U3736 (N_3736,In_1484,In_1861);
or U3737 (N_3737,In_192,In_280);
and U3738 (N_3738,In_1984,In_1518);
nand U3739 (N_3739,In_72,In_996);
and U3740 (N_3740,In_1282,In_1974);
nor U3741 (N_3741,In_357,In_1128);
and U3742 (N_3742,In_1763,In_373);
and U3743 (N_3743,In_1324,In_849);
nand U3744 (N_3744,In_225,In_589);
and U3745 (N_3745,In_38,In_939);
and U3746 (N_3746,In_1773,In_1287);
and U3747 (N_3747,In_1940,In_109);
or U3748 (N_3748,In_455,In_442);
and U3749 (N_3749,In_1803,In_126);
or U3750 (N_3750,In_294,In_230);
nand U3751 (N_3751,In_1670,In_248);
and U3752 (N_3752,In_567,In_1693);
and U3753 (N_3753,In_925,In_609);
nor U3754 (N_3754,In_1855,In_192);
or U3755 (N_3755,In_1404,In_1487);
or U3756 (N_3756,In_1487,In_123);
nor U3757 (N_3757,In_1765,In_1553);
or U3758 (N_3758,In_1418,In_806);
or U3759 (N_3759,In_909,In_582);
nand U3760 (N_3760,In_1297,In_981);
nand U3761 (N_3761,In_1992,In_1835);
nand U3762 (N_3762,In_107,In_1961);
nor U3763 (N_3763,In_20,In_238);
nand U3764 (N_3764,In_669,In_442);
or U3765 (N_3765,In_744,In_1183);
nand U3766 (N_3766,In_1410,In_1764);
nor U3767 (N_3767,In_1597,In_1898);
nor U3768 (N_3768,In_868,In_1843);
nand U3769 (N_3769,In_1690,In_59);
and U3770 (N_3770,In_1141,In_484);
and U3771 (N_3771,In_1228,In_505);
and U3772 (N_3772,In_1136,In_414);
or U3773 (N_3773,In_1957,In_1755);
nand U3774 (N_3774,In_48,In_279);
xor U3775 (N_3775,In_334,In_1010);
nand U3776 (N_3776,In_1984,In_1931);
nand U3777 (N_3777,In_447,In_1395);
nor U3778 (N_3778,In_1314,In_1518);
nand U3779 (N_3779,In_986,In_1296);
or U3780 (N_3780,In_281,In_1113);
nand U3781 (N_3781,In_1596,In_1350);
or U3782 (N_3782,In_463,In_808);
and U3783 (N_3783,In_4,In_1113);
xor U3784 (N_3784,In_1738,In_1305);
nor U3785 (N_3785,In_391,In_831);
and U3786 (N_3786,In_266,In_930);
and U3787 (N_3787,In_1609,In_1772);
and U3788 (N_3788,In_404,In_574);
nor U3789 (N_3789,In_523,In_1650);
nand U3790 (N_3790,In_1505,In_1160);
nand U3791 (N_3791,In_1792,In_656);
nor U3792 (N_3792,In_512,In_623);
and U3793 (N_3793,In_25,In_281);
or U3794 (N_3794,In_1645,In_1625);
nor U3795 (N_3795,In_1402,In_966);
or U3796 (N_3796,In_1144,In_698);
nor U3797 (N_3797,In_515,In_1798);
nand U3798 (N_3798,In_1375,In_1260);
xnor U3799 (N_3799,In_509,In_1296);
nand U3800 (N_3800,In_713,In_344);
nand U3801 (N_3801,In_1414,In_981);
and U3802 (N_3802,In_1487,In_823);
nand U3803 (N_3803,In_1741,In_366);
nand U3804 (N_3804,In_1358,In_1143);
and U3805 (N_3805,In_318,In_1563);
nor U3806 (N_3806,In_1494,In_1798);
nor U3807 (N_3807,In_1448,In_366);
and U3808 (N_3808,In_372,In_998);
or U3809 (N_3809,In_720,In_1094);
or U3810 (N_3810,In_238,In_18);
and U3811 (N_3811,In_1538,In_232);
nand U3812 (N_3812,In_800,In_1271);
nor U3813 (N_3813,In_1494,In_4);
and U3814 (N_3814,In_142,In_1765);
nand U3815 (N_3815,In_1724,In_240);
nor U3816 (N_3816,In_1793,In_481);
or U3817 (N_3817,In_1739,In_621);
nand U3818 (N_3818,In_388,In_132);
xnor U3819 (N_3819,In_1332,In_1210);
nor U3820 (N_3820,In_987,In_390);
nor U3821 (N_3821,In_1623,In_1592);
or U3822 (N_3822,In_1727,In_1445);
xor U3823 (N_3823,In_154,In_1649);
or U3824 (N_3824,In_185,In_755);
xor U3825 (N_3825,In_1263,In_550);
nor U3826 (N_3826,In_8,In_1432);
nor U3827 (N_3827,In_1797,In_683);
and U3828 (N_3828,In_200,In_932);
and U3829 (N_3829,In_1598,In_1045);
nor U3830 (N_3830,In_1920,In_899);
nor U3831 (N_3831,In_3,In_1902);
nor U3832 (N_3832,In_235,In_844);
xor U3833 (N_3833,In_1441,In_1997);
nor U3834 (N_3834,In_102,In_720);
nor U3835 (N_3835,In_991,In_1412);
and U3836 (N_3836,In_1025,In_415);
or U3837 (N_3837,In_1978,In_1747);
and U3838 (N_3838,In_1585,In_1435);
nand U3839 (N_3839,In_298,In_1777);
nand U3840 (N_3840,In_1401,In_670);
nor U3841 (N_3841,In_429,In_1895);
nor U3842 (N_3842,In_1210,In_707);
and U3843 (N_3843,In_1970,In_1860);
nor U3844 (N_3844,In_1159,In_578);
and U3845 (N_3845,In_559,In_952);
xnor U3846 (N_3846,In_1232,In_300);
xnor U3847 (N_3847,In_1477,In_1349);
nand U3848 (N_3848,In_300,In_55);
nand U3849 (N_3849,In_1316,In_227);
nor U3850 (N_3850,In_1558,In_18);
xor U3851 (N_3851,In_1249,In_1284);
nor U3852 (N_3852,In_1252,In_842);
nor U3853 (N_3853,In_186,In_34);
nand U3854 (N_3854,In_630,In_1803);
or U3855 (N_3855,In_74,In_378);
or U3856 (N_3856,In_1579,In_1936);
nor U3857 (N_3857,In_841,In_1379);
and U3858 (N_3858,In_48,In_1557);
and U3859 (N_3859,In_99,In_1324);
nand U3860 (N_3860,In_1633,In_174);
and U3861 (N_3861,In_1515,In_798);
nor U3862 (N_3862,In_1668,In_1128);
or U3863 (N_3863,In_1248,In_1865);
nor U3864 (N_3864,In_18,In_1009);
nand U3865 (N_3865,In_1506,In_1507);
and U3866 (N_3866,In_147,In_1515);
and U3867 (N_3867,In_247,In_546);
nor U3868 (N_3868,In_564,In_1542);
or U3869 (N_3869,In_1371,In_873);
nor U3870 (N_3870,In_1394,In_1136);
nand U3871 (N_3871,In_102,In_1313);
or U3872 (N_3872,In_850,In_361);
and U3873 (N_3873,In_343,In_1629);
nand U3874 (N_3874,In_1551,In_1443);
nand U3875 (N_3875,In_958,In_740);
nor U3876 (N_3876,In_1641,In_1313);
nand U3877 (N_3877,In_1516,In_1223);
nor U3878 (N_3878,In_882,In_394);
nand U3879 (N_3879,In_786,In_842);
xor U3880 (N_3880,In_1821,In_57);
nor U3881 (N_3881,In_326,In_242);
or U3882 (N_3882,In_1628,In_563);
or U3883 (N_3883,In_747,In_320);
xor U3884 (N_3884,In_380,In_1638);
and U3885 (N_3885,In_1515,In_1124);
and U3886 (N_3886,In_401,In_1742);
and U3887 (N_3887,In_769,In_476);
nand U3888 (N_3888,In_148,In_786);
or U3889 (N_3889,In_249,In_541);
and U3890 (N_3890,In_1223,In_1008);
nor U3891 (N_3891,In_173,In_1848);
nor U3892 (N_3892,In_1825,In_1770);
nor U3893 (N_3893,In_450,In_1147);
nor U3894 (N_3894,In_446,In_1919);
or U3895 (N_3895,In_125,In_1967);
nand U3896 (N_3896,In_463,In_1378);
nor U3897 (N_3897,In_178,In_900);
and U3898 (N_3898,In_831,In_1461);
or U3899 (N_3899,In_1742,In_1134);
xnor U3900 (N_3900,In_1620,In_297);
nor U3901 (N_3901,In_90,In_984);
or U3902 (N_3902,In_919,In_238);
nand U3903 (N_3903,In_979,In_1434);
or U3904 (N_3904,In_412,In_514);
and U3905 (N_3905,In_579,In_438);
xnor U3906 (N_3906,In_1658,In_1971);
nand U3907 (N_3907,In_1988,In_811);
nand U3908 (N_3908,In_907,In_1855);
nand U3909 (N_3909,In_268,In_105);
or U3910 (N_3910,In_98,In_174);
and U3911 (N_3911,In_626,In_1923);
nor U3912 (N_3912,In_1460,In_100);
xnor U3913 (N_3913,In_513,In_1482);
and U3914 (N_3914,In_1698,In_17);
nand U3915 (N_3915,In_592,In_159);
and U3916 (N_3916,In_1506,In_1964);
or U3917 (N_3917,In_1078,In_1541);
or U3918 (N_3918,In_105,In_1600);
nand U3919 (N_3919,In_751,In_1050);
nand U3920 (N_3920,In_382,In_1445);
nor U3921 (N_3921,In_536,In_138);
nand U3922 (N_3922,In_1960,In_1574);
or U3923 (N_3923,In_1270,In_1792);
nor U3924 (N_3924,In_1314,In_174);
nand U3925 (N_3925,In_523,In_1503);
xor U3926 (N_3926,In_1159,In_1057);
or U3927 (N_3927,In_410,In_412);
nor U3928 (N_3928,In_1322,In_1441);
nor U3929 (N_3929,In_165,In_292);
nand U3930 (N_3930,In_1940,In_1816);
nor U3931 (N_3931,In_912,In_740);
nand U3932 (N_3932,In_149,In_612);
xor U3933 (N_3933,In_429,In_1336);
or U3934 (N_3934,In_686,In_1264);
xnor U3935 (N_3935,In_720,In_227);
nand U3936 (N_3936,In_866,In_456);
nand U3937 (N_3937,In_738,In_1233);
nand U3938 (N_3938,In_671,In_1005);
or U3939 (N_3939,In_1182,In_1929);
xor U3940 (N_3940,In_1265,In_968);
nand U3941 (N_3941,In_1767,In_219);
and U3942 (N_3942,In_953,In_1069);
nor U3943 (N_3943,In_1479,In_1904);
and U3944 (N_3944,In_379,In_1315);
and U3945 (N_3945,In_1886,In_507);
nor U3946 (N_3946,In_81,In_1412);
nor U3947 (N_3947,In_21,In_856);
nand U3948 (N_3948,In_1375,In_1933);
nor U3949 (N_3949,In_547,In_162);
or U3950 (N_3950,In_544,In_1205);
nand U3951 (N_3951,In_1322,In_1895);
or U3952 (N_3952,In_213,In_624);
xnor U3953 (N_3953,In_597,In_902);
or U3954 (N_3954,In_452,In_557);
nand U3955 (N_3955,In_1056,In_433);
or U3956 (N_3956,In_432,In_246);
or U3957 (N_3957,In_869,In_892);
nand U3958 (N_3958,In_1007,In_385);
nand U3959 (N_3959,In_1090,In_1831);
and U3960 (N_3960,In_1198,In_1596);
or U3961 (N_3961,In_204,In_57);
nor U3962 (N_3962,In_901,In_716);
nand U3963 (N_3963,In_1677,In_1251);
xnor U3964 (N_3964,In_1008,In_1930);
or U3965 (N_3965,In_214,In_568);
and U3966 (N_3966,In_1925,In_818);
and U3967 (N_3967,In_785,In_1937);
nand U3968 (N_3968,In_992,In_528);
nor U3969 (N_3969,In_505,In_758);
or U3970 (N_3970,In_192,In_1896);
or U3971 (N_3971,In_1686,In_783);
and U3972 (N_3972,In_663,In_1497);
or U3973 (N_3973,In_1947,In_592);
or U3974 (N_3974,In_594,In_355);
or U3975 (N_3975,In_440,In_1872);
xnor U3976 (N_3976,In_1407,In_399);
and U3977 (N_3977,In_357,In_190);
and U3978 (N_3978,In_142,In_1431);
xnor U3979 (N_3979,In_102,In_1375);
xnor U3980 (N_3980,In_561,In_1441);
nand U3981 (N_3981,In_63,In_502);
or U3982 (N_3982,In_384,In_685);
or U3983 (N_3983,In_1733,In_949);
nor U3984 (N_3984,In_1276,In_1852);
or U3985 (N_3985,In_1543,In_1683);
and U3986 (N_3986,In_798,In_176);
nor U3987 (N_3987,In_1840,In_554);
nand U3988 (N_3988,In_883,In_834);
nand U3989 (N_3989,In_1052,In_1785);
and U3990 (N_3990,In_1936,In_1854);
nand U3991 (N_3991,In_927,In_1857);
xor U3992 (N_3992,In_1118,In_1984);
nor U3993 (N_3993,In_1238,In_1245);
nand U3994 (N_3994,In_1549,In_1045);
nand U3995 (N_3995,In_812,In_244);
or U3996 (N_3996,In_1375,In_525);
nand U3997 (N_3997,In_492,In_808);
nor U3998 (N_3998,In_1937,In_1129);
nand U3999 (N_3999,In_1664,In_837);
nand U4000 (N_4000,N_562,N_1113);
and U4001 (N_4001,N_2643,N_1502);
nor U4002 (N_4002,N_3712,N_1648);
xor U4003 (N_4003,N_2322,N_35);
and U4004 (N_4004,N_3748,N_982);
nor U4005 (N_4005,N_1540,N_3006);
and U4006 (N_4006,N_2830,N_3980);
and U4007 (N_4007,N_702,N_2862);
nor U4008 (N_4008,N_3119,N_372);
nor U4009 (N_4009,N_229,N_1199);
nand U4010 (N_4010,N_2492,N_2432);
and U4011 (N_4011,N_944,N_2619);
or U4012 (N_4012,N_3796,N_61);
or U4013 (N_4013,N_2631,N_802);
and U4014 (N_4014,N_2968,N_3561);
and U4015 (N_4015,N_2034,N_654);
xor U4016 (N_4016,N_632,N_3637);
nor U4017 (N_4017,N_3328,N_2630);
or U4018 (N_4018,N_823,N_1618);
nand U4019 (N_4019,N_675,N_256);
and U4020 (N_4020,N_3440,N_2025);
xor U4021 (N_4021,N_1727,N_3351);
xnor U4022 (N_4022,N_886,N_2194);
nand U4023 (N_4023,N_3598,N_1320);
and U4024 (N_4024,N_2806,N_3989);
or U4025 (N_4025,N_3631,N_2);
or U4026 (N_4026,N_3145,N_2576);
and U4027 (N_4027,N_939,N_1840);
or U4028 (N_4028,N_3528,N_3397);
nor U4029 (N_4029,N_2129,N_717);
nand U4030 (N_4030,N_413,N_1243);
or U4031 (N_4031,N_3024,N_3965);
nand U4032 (N_4032,N_3572,N_1421);
nand U4033 (N_4033,N_1074,N_3698);
and U4034 (N_4034,N_3322,N_2161);
and U4035 (N_4035,N_3746,N_2735);
nand U4036 (N_4036,N_2902,N_48);
or U4037 (N_4037,N_1459,N_1955);
or U4038 (N_4038,N_1065,N_480);
or U4039 (N_4039,N_1439,N_214);
and U4040 (N_4040,N_2912,N_2731);
and U4041 (N_4041,N_2487,N_3009);
nor U4042 (N_4042,N_2627,N_350);
or U4043 (N_4043,N_3384,N_1341);
and U4044 (N_4044,N_1495,N_1147);
xor U4045 (N_4045,N_2182,N_196);
nand U4046 (N_4046,N_220,N_512);
and U4047 (N_4047,N_1822,N_3850);
or U4048 (N_4048,N_3043,N_2003);
and U4049 (N_4049,N_2148,N_793);
nor U4050 (N_4050,N_1474,N_1970);
or U4051 (N_4051,N_596,N_3793);
nor U4052 (N_4052,N_1482,N_3786);
nor U4053 (N_4053,N_1164,N_1914);
nor U4054 (N_4054,N_1333,N_3467);
or U4055 (N_4055,N_2197,N_2698);
nor U4056 (N_4056,N_73,N_1256);
or U4057 (N_4057,N_2573,N_3427);
and U4058 (N_4058,N_854,N_1782);
nor U4059 (N_4059,N_3608,N_3183);
nor U4060 (N_4060,N_348,N_129);
or U4061 (N_4061,N_3843,N_2589);
or U4062 (N_4062,N_820,N_2447);
and U4063 (N_4063,N_2469,N_565);
nor U4064 (N_4064,N_2337,N_3305);
nand U4065 (N_4065,N_663,N_1823);
or U4066 (N_4066,N_732,N_1275);
and U4067 (N_4067,N_438,N_1441);
or U4068 (N_4068,N_3299,N_1794);
nand U4069 (N_4069,N_1494,N_243);
nor U4070 (N_4070,N_2092,N_996);
nand U4071 (N_4071,N_2564,N_3184);
and U4072 (N_4072,N_1934,N_2345);
nand U4073 (N_4073,N_3066,N_1192);
or U4074 (N_4074,N_2470,N_3747);
or U4075 (N_4075,N_116,N_2036);
and U4076 (N_4076,N_2012,N_2821);
or U4077 (N_4077,N_1385,N_3563);
nand U4078 (N_4078,N_2227,N_1242);
nand U4079 (N_4079,N_1141,N_1774);
or U4080 (N_4080,N_3016,N_241);
and U4081 (N_4081,N_175,N_2050);
and U4082 (N_4082,N_1396,N_756);
nand U4083 (N_4083,N_314,N_113);
and U4084 (N_4084,N_2230,N_1738);
or U4085 (N_4085,N_1881,N_2645);
nand U4086 (N_4086,N_1852,N_1995);
nand U4087 (N_4087,N_2316,N_2325);
and U4088 (N_4088,N_1520,N_3863);
or U4089 (N_4089,N_3915,N_3599);
or U4090 (N_4090,N_3114,N_2008);
nand U4091 (N_4091,N_3679,N_3994);
nand U4092 (N_4092,N_2261,N_1077);
nor U4093 (N_4093,N_183,N_388);
and U4094 (N_4094,N_1829,N_2856);
nand U4095 (N_4095,N_2608,N_3671);
nand U4096 (N_4096,N_2370,N_3412);
nand U4097 (N_4097,N_3837,N_2499);
nor U4098 (N_4098,N_3073,N_2359);
and U4099 (N_4099,N_2905,N_2181);
and U4100 (N_4100,N_642,N_12);
or U4101 (N_4101,N_2247,N_3065);
and U4102 (N_4102,N_1041,N_2871);
or U4103 (N_4103,N_2449,N_2820);
and U4104 (N_4104,N_2880,N_2309);
nand U4105 (N_4105,N_2504,N_2314);
or U4106 (N_4106,N_3347,N_1231);
nor U4107 (N_4107,N_1045,N_743);
nand U4108 (N_4108,N_1317,N_2216);
nor U4109 (N_4109,N_2738,N_2157);
nor U4110 (N_4110,N_3870,N_1859);
nor U4111 (N_4111,N_3583,N_941);
nor U4112 (N_4112,N_3281,N_967);
and U4113 (N_4113,N_1454,N_2199);
or U4114 (N_4114,N_2524,N_2623);
and U4115 (N_4115,N_184,N_1527);
and U4116 (N_4116,N_3548,N_3873);
nand U4117 (N_4117,N_1958,N_3054);
and U4118 (N_4118,N_3929,N_3869);
nor U4119 (N_4119,N_3996,N_3271);
nand U4120 (N_4120,N_3042,N_3378);
nand U4121 (N_4121,N_1068,N_2693);
nor U4122 (N_4122,N_123,N_359);
and U4123 (N_4123,N_799,N_223);
or U4124 (N_4124,N_1665,N_3550);
or U4125 (N_4125,N_227,N_2975);
or U4126 (N_4126,N_940,N_3758);
or U4127 (N_4127,N_689,N_2486);
or U4128 (N_4128,N_1062,N_3590);
and U4129 (N_4129,N_1851,N_3532);
nand U4130 (N_4130,N_3576,N_1266);
or U4131 (N_4131,N_211,N_588);
or U4132 (N_4132,N_526,N_1625);
or U4133 (N_4133,N_1432,N_3382);
and U4134 (N_4134,N_534,N_788);
and U4135 (N_4135,N_1327,N_2707);
nor U4136 (N_4136,N_3275,N_155);
or U4137 (N_4137,N_2713,N_1127);
and U4138 (N_4138,N_3422,N_2768);
nand U4139 (N_4139,N_666,N_1388);
and U4140 (N_4140,N_1215,N_244);
and U4141 (N_4141,N_3824,N_444);
nand U4142 (N_4142,N_570,N_784);
nor U4143 (N_4143,N_3071,N_3567);
nor U4144 (N_4144,N_2037,N_1532);
nor U4145 (N_4145,N_2026,N_3015);
or U4146 (N_4146,N_3188,N_1673);
and U4147 (N_4147,N_898,N_1078);
nor U4148 (N_4148,N_3147,N_1438);
nor U4149 (N_4149,N_2750,N_1216);
or U4150 (N_4150,N_1060,N_1724);
xor U4151 (N_4151,N_3539,N_2391);
xor U4152 (N_4152,N_1095,N_1012);
and U4153 (N_4153,N_1966,N_3948);
or U4154 (N_4154,N_605,N_1050);
nor U4155 (N_4155,N_210,N_3256);
nor U4156 (N_4156,N_1815,N_3797);
or U4157 (N_4157,N_3922,N_569);
nor U4158 (N_4158,N_923,N_3137);
nand U4159 (N_4159,N_1945,N_490);
nor U4160 (N_4160,N_672,N_3955);
nand U4161 (N_4161,N_1098,N_1509);
nand U4162 (N_4162,N_3341,N_3151);
nand U4163 (N_4163,N_1337,N_3966);
nor U4164 (N_4164,N_2537,N_2150);
or U4165 (N_4165,N_3359,N_2833);
and U4166 (N_4166,N_1027,N_2393);
nand U4167 (N_4167,N_1884,N_3215);
or U4168 (N_4168,N_3686,N_3619);
or U4169 (N_4169,N_3925,N_1916);
nor U4170 (N_4170,N_2593,N_1401);
nor U4171 (N_4171,N_2403,N_2387);
and U4172 (N_4172,N_1947,N_1197);
xnor U4173 (N_4173,N_1671,N_455);
or U4174 (N_4174,N_2443,N_309);
and U4175 (N_4175,N_3983,N_369);
nand U4176 (N_4176,N_1226,N_1982);
and U4177 (N_4177,N_2616,N_771);
nor U4178 (N_4178,N_3033,N_772);
nand U4179 (N_4179,N_584,N_1225);
nand U4180 (N_4180,N_806,N_2584);
nand U4181 (N_4181,N_3160,N_2176);
nand U4182 (N_4182,N_60,N_1683);
nand U4183 (N_4183,N_197,N_3909);
or U4184 (N_4184,N_1725,N_1559);
nand U4185 (N_4185,N_3673,N_2895);
or U4186 (N_4186,N_3931,N_2217);
nor U4187 (N_4187,N_3834,N_2474);
and U4188 (N_4188,N_2172,N_74);
or U4189 (N_4189,N_1783,N_149);
nand U4190 (N_4190,N_2254,N_1332);
nor U4191 (N_4191,N_794,N_166);
or U4192 (N_4192,N_2045,N_1138);
nor U4193 (N_4193,N_2634,N_3798);
or U4194 (N_4194,N_208,N_3294);
and U4195 (N_4195,N_892,N_3064);
xnor U4196 (N_4196,N_961,N_1824);
xor U4197 (N_4197,N_2596,N_3193);
or U4198 (N_4198,N_1573,N_3441);
or U4199 (N_4199,N_894,N_3142);
nand U4200 (N_4200,N_224,N_2427);
and U4201 (N_4201,N_2746,N_2699);
nand U4202 (N_4202,N_1087,N_2030);
and U4203 (N_4203,N_1651,N_2444);
and U4204 (N_4204,N_288,N_1953);
and U4205 (N_4205,N_2581,N_1608);
nor U4206 (N_4206,N_1445,N_958);
and U4207 (N_4207,N_2467,N_259);
or U4208 (N_4208,N_2591,N_3239);
nand U4209 (N_4209,N_1892,N_1518);
nand U4210 (N_4210,N_2782,N_2859);
or U4211 (N_4211,N_3379,N_3836);
nand U4212 (N_4212,N_3404,N_375);
and U4213 (N_4213,N_1489,N_2389);
nor U4214 (N_4214,N_2369,N_847);
and U4215 (N_4215,N_1365,N_1239);
nor U4216 (N_4216,N_2670,N_3571);
and U4217 (N_4217,N_3725,N_1517);
and U4218 (N_4218,N_3987,N_3454);
and U4219 (N_4219,N_3968,N_2560);
or U4220 (N_4220,N_1100,N_1780);
xor U4221 (N_4221,N_3486,N_2233);
xor U4222 (N_4222,N_2689,N_2672);
and U4223 (N_4223,N_2915,N_946);
and U4224 (N_4224,N_1252,N_703);
and U4225 (N_4225,N_1775,N_3167);
and U4226 (N_4226,N_64,N_2722);
nand U4227 (N_4227,N_1771,N_1543);
or U4228 (N_4228,N_2588,N_89);
xnor U4229 (N_4229,N_1735,N_1580);
or U4230 (N_4230,N_1374,N_680);
nor U4231 (N_4231,N_2826,N_3484);
nor U4232 (N_4232,N_1922,N_2298);
nor U4233 (N_4233,N_2123,N_895);
xnor U4234 (N_4234,N_1654,N_2542);
nand U4235 (N_4235,N_1781,N_3990);
or U4236 (N_4236,N_1709,N_525);
nor U4237 (N_4237,N_1435,N_2759);
and U4238 (N_4238,N_263,N_2433);
nand U4239 (N_4239,N_1081,N_699);
or U4240 (N_4240,N_3287,N_2574);
nor U4241 (N_4241,N_720,N_3889);
or U4242 (N_4242,N_1854,N_1300);
nand U4243 (N_4243,N_1280,N_465);
nand U4244 (N_4244,N_2076,N_2002);
nand U4245 (N_4245,N_3506,N_1359);
or U4246 (N_4246,N_2151,N_298);
nand U4247 (N_4247,N_3757,N_3858);
nor U4248 (N_4248,N_189,N_585);
and U4249 (N_4249,N_3267,N_590);
xor U4250 (N_4250,N_1760,N_399);
nand U4251 (N_4251,N_606,N_3904);
or U4252 (N_4252,N_835,N_640);
nor U4253 (N_4253,N_3330,N_1528);
nor U4254 (N_4254,N_2603,N_2162);
and U4255 (N_4255,N_2484,N_99);
nor U4256 (N_4256,N_2018,N_627);
nor U4257 (N_4257,N_2855,N_2421);
and U4258 (N_4258,N_3888,N_3026);
nor U4259 (N_4259,N_1986,N_2801);
xor U4260 (N_4260,N_3315,N_3704);
nand U4261 (N_4261,N_376,N_93);
nor U4262 (N_4262,N_2005,N_832);
nor U4263 (N_4263,N_2411,N_3691);
or U4264 (N_4264,N_3639,N_1344);
nand U4265 (N_4265,N_3210,N_1057);
xor U4266 (N_4266,N_333,N_275);
or U4267 (N_4267,N_1299,N_2945);
nor U4268 (N_4268,N_910,N_1857);
nor U4269 (N_4269,N_2152,N_2897);
or U4270 (N_4270,N_266,N_1537);
nor U4271 (N_4271,N_3775,N_2347);
nand U4272 (N_4272,N_2877,N_908);
nand U4273 (N_4273,N_3876,N_942);
and U4274 (N_4274,N_1366,N_2927);
or U4275 (N_4275,N_1719,N_2223);
nor U4276 (N_4276,N_1550,N_1377);
or U4277 (N_4277,N_1515,N_158);
nand U4278 (N_4278,N_1981,N_2500);
nand U4279 (N_4279,N_3817,N_1467);
nand U4280 (N_4280,N_1563,N_2453);
nor U4281 (N_4281,N_434,N_2694);
and U4282 (N_4282,N_454,N_2536);
or U4283 (N_4283,N_3102,N_1898);
nor U4284 (N_4284,N_1777,N_3468);
and U4285 (N_4285,N_2088,N_392);
or U4286 (N_4286,N_3039,N_2562);
and U4287 (N_4287,N_13,N_308);
nor U4288 (N_4288,N_1860,N_2202);
nand U4289 (N_4289,N_3162,N_1909);
xnor U4290 (N_4290,N_3587,N_2349);
nor U4291 (N_4291,N_3135,N_2242);
nand U4292 (N_4292,N_3428,N_2684);
and U4293 (N_4293,N_3891,N_613);
or U4294 (N_4294,N_1716,N_501);
nor U4295 (N_4295,N_758,N_3010);
or U4296 (N_4296,N_3981,N_3616);
xnor U4297 (N_4297,N_3290,N_1265);
or U4298 (N_4298,N_3951,N_2983);
or U4299 (N_4299,N_1646,N_3603);
and U4300 (N_4300,N_2490,N_1075);
and U4301 (N_4301,N_2118,N_1714);
nor U4302 (N_4302,N_3985,N_2366);
or U4303 (N_4303,N_869,N_306);
or U4304 (N_4304,N_2650,N_594);
xnor U4305 (N_4305,N_1007,N_1832);
and U4306 (N_4306,N_57,N_3360);
xnor U4307 (N_4307,N_1624,N_3419);
xor U4308 (N_4308,N_2111,N_10);
or U4309 (N_4309,N_2131,N_1754);
or U4310 (N_4310,N_1734,N_2571);
and U4311 (N_4311,N_3722,N_861);
nor U4312 (N_4312,N_2060,N_2851);
nor U4313 (N_4313,N_2971,N_3091);
and U4314 (N_4314,N_102,N_620);
or U4315 (N_4315,N_1340,N_3005);
nor U4316 (N_4316,N_172,N_803);
nand U4317 (N_4317,N_2778,N_1162);
nand U4318 (N_4318,N_1921,N_2052);
nand U4319 (N_4319,N_112,N_2988);
nor U4320 (N_4320,N_3377,N_3920);
and U4321 (N_4321,N_3957,N_2710);
xnor U4322 (N_4322,N_2275,N_1996);
and U4323 (N_4323,N_779,N_3235);
or U4324 (N_4324,N_915,N_3736);
and U4325 (N_4325,N_474,N_3094);
nor U4326 (N_4326,N_2068,N_3217);
nand U4327 (N_4327,N_1336,N_1865);
nand U4328 (N_4328,N_631,N_2072);
or U4329 (N_4329,N_1311,N_2132);
nand U4330 (N_4330,N_3199,N_3317);
or U4331 (N_4331,N_1929,N_3866);
or U4332 (N_4332,N_3477,N_2256);
nor U4333 (N_4333,N_1507,N_1117);
and U4334 (N_4334,N_3662,N_192);
or U4335 (N_4335,N_955,N_1181);
nand U4336 (N_4336,N_2458,N_1497);
or U4337 (N_4337,N_529,N_738);
or U4338 (N_4338,N_1711,N_3895);
xnor U4339 (N_4339,N_1670,N_3614);
nor U4340 (N_4340,N_669,N_3783);
and U4341 (N_4341,N_3122,N_2064);
nand U4342 (N_4342,N_2953,N_151);
and U4343 (N_4343,N_3546,N_1353);
or U4344 (N_4344,N_3175,N_2662);
xnor U4345 (N_4345,N_124,N_906);
and U4346 (N_4346,N_609,N_842);
or U4347 (N_4347,N_2292,N_1911);
and U4348 (N_4348,N_1429,N_1577);
and U4349 (N_4349,N_2957,N_3911);
and U4350 (N_4350,N_714,N_3963);
nand U4351 (N_4351,N_104,N_1927);
and U4352 (N_4352,N_1593,N_69);
nor U4353 (N_4353,N_1967,N_2290);
xor U4354 (N_4354,N_2297,N_911);
nand U4355 (N_4355,N_3582,N_1620);
nand U4356 (N_4356,N_1685,N_320);
or U4357 (N_4357,N_2838,N_2919);
or U4358 (N_4358,N_3325,N_1133);
or U4359 (N_4359,N_888,N_2244);
nand U4360 (N_4360,N_2083,N_3597);
or U4361 (N_4361,N_1842,N_1667);
and U4362 (N_4362,N_499,N_2554);
and U4363 (N_4363,N_2402,N_398);
and U4364 (N_4364,N_3406,N_1490);
or U4365 (N_4365,N_3182,N_2405);
nand U4366 (N_4366,N_3237,N_3696);
nor U4367 (N_4367,N_2528,N_1188);
and U4368 (N_4368,N_1603,N_3128);
nor U4369 (N_4369,N_121,N_1574);
xnor U4370 (N_4370,N_3898,N_1013);
nor U4371 (N_4371,N_1586,N_3943);
or U4372 (N_4372,N_3314,N_2993);
or U4373 (N_4373,N_2201,N_960);
nand U4374 (N_4374,N_3855,N_1297);
and U4375 (N_4375,N_1157,N_2841);
and U4376 (N_4376,N_1814,N_3710);
nand U4377 (N_4377,N_3345,N_696);
and U4378 (N_4378,N_1839,N_3264);
nor U4379 (N_4379,N_95,N_1902);
nand U4380 (N_4380,N_3763,N_791);
or U4381 (N_4381,N_2488,N_3211);
nand U4382 (N_4382,N_2311,N_1161);
nor U4383 (N_4383,N_3297,N_2943);
or U4384 (N_4384,N_1599,N_2091);
nor U4385 (N_4385,N_177,N_443);
nand U4386 (N_4386,N_1129,N_2221);
and U4387 (N_4387,N_2512,N_2042);
nand U4388 (N_4388,N_579,N_2677);
and U4389 (N_4389,N_3103,N_2679);
and U4390 (N_4390,N_2107,N_3618);
or U4391 (N_4391,N_3472,N_2613);
and U4392 (N_4392,N_1640,N_3367);
nor U4393 (N_4393,N_382,N_1170);
and U4394 (N_4394,N_2455,N_1579);
or U4395 (N_4395,N_2465,N_2959);
and U4396 (N_4396,N_807,N_3672);
nand U4397 (N_4397,N_546,N_1669);
nor U4398 (N_4398,N_3740,N_2476);
and U4399 (N_4399,N_3827,N_2878);
and U4400 (N_4400,N_2480,N_1952);
and U4401 (N_4401,N_3840,N_1793);
nor U4402 (N_4402,N_1255,N_3070);
nor U4403 (N_4403,N_2675,N_3670);
and U4404 (N_4404,N_3212,N_1492);
nand U4405 (N_4405,N_2485,N_3390);
and U4406 (N_4406,N_2812,N_414);
nand U4407 (N_4407,N_2166,N_995);
xor U4408 (N_4408,N_511,N_134);
or U4409 (N_4409,N_1871,N_3201);
or U4410 (N_4410,N_2920,N_2867);
or U4411 (N_4411,N_1044,N_1469);
nor U4412 (N_4412,N_3003,N_3495);
nor U4413 (N_4413,N_2914,N_2509);
and U4414 (N_4414,N_3106,N_3079);
and U4415 (N_4415,N_478,N_2657);
xnor U4416 (N_4416,N_2348,N_1984);
nor U4417 (N_4417,N_2318,N_2543);
nand U4418 (N_4418,N_3659,N_366);
nor U4419 (N_4419,N_2991,N_1296);
and U4420 (N_4420,N_1739,N_246);
or U4421 (N_4421,N_507,N_1473);
nand U4422 (N_4422,N_1331,N_2028);
nand U4423 (N_4423,N_3971,N_2475);
nand U4424 (N_4424,N_2377,N_1283);
or U4425 (N_4425,N_3490,N_2113);
nand U4426 (N_4426,N_3737,N_2415);
or U4427 (N_4427,N_3007,N_530);
nor U4428 (N_4428,N_451,N_135);
or U4429 (N_4429,N_318,N_2893);
or U4430 (N_4430,N_762,N_765);
nand U4431 (N_4431,N_3092,N_670);
nor U4432 (N_4432,N_3534,N_2146);
nand U4433 (N_4433,N_437,N_363);
and U4434 (N_4434,N_2206,N_2695);
nor U4435 (N_4435,N_686,N_598);
and U4436 (N_4436,N_1318,N_1182);
nand U4437 (N_4437,N_1820,N_2872);
nor U4438 (N_4438,N_2279,N_984);
nand U4439 (N_4439,N_810,N_1430);
and U4440 (N_4440,N_2418,N_1416);
nor U4441 (N_4441,N_3914,N_824);
and U4442 (N_4442,N_646,N_2374);
nand U4443 (N_4443,N_2268,N_1362);
nor U4444 (N_4444,N_2013,N_3214);
and U4445 (N_4445,N_3683,N_3286);
or U4446 (N_4446,N_449,N_3335);
nor U4447 (N_4447,N_3560,N_757);
xnor U4448 (N_4448,N_3984,N_3650);
nor U4449 (N_4449,N_3084,N_117);
or U4450 (N_4450,N_336,N_1221);
and U4451 (N_4451,N_2653,N_494);
and U4452 (N_4452,N_834,N_3475);
nor U4453 (N_4453,N_3407,N_3832);
and U4454 (N_4454,N_22,N_2610);
xor U4455 (N_4455,N_1812,N_2135);
nor U4456 (N_4456,N_1034,N_3625);
or U4457 (N_4457,N_1792,N_1159);
or U4458 (N_4458,N_3905,N_2375);
and U4459 (N_4459,N_1604,N_1612);
nand U4460 (N_4460,N_2765,N_2997);
nand U4461 (N_4461,N_1072,N_432);
or U4462 (N_4462,N_1906,N_3735);
and U4463 (N_4463,N_539,N_1557);
nor U4464 (N_4464,N_851,N_905);
and U4465 (N_4465,N_798,N_3681);
xnor U4466 (N_4466,N_1185,N_976);
nor U4467 (N_4467,N_3306,N_3172);
or U4468 (N_4468,N_3265,N_2756);
nand U4469 (N_4469,N_354,N_3794);
and U4470 (N_4470,N_3324,N_805);
and U4471 (N_4471,N_1102,N_254);
and U4472 (N_4472,N_3730,N_3292);
and U4473 (N_4473,N_2070,N_1307);
and U4474 (N_4474,N_389,N_2436);
and U4475 (N_4475,N_3320,N_2930);
xor U4476 (N_4476,N_1622,N_2976);
nor U4477 (N_4477,N_2205,N_137);
xor U4478 (N_4478,N_357,N_1251);
or U4479 (N_4479,N_2674,N_3434);
and U4480 (N_4480,N_746,N_3236);
nor U4481 (N_4481,N_1219,N_1524);
nand U4482 (N_4482,N_3721,N_3370);
nand U4483 (N_4483,N_890,N_317);
nor U4484 (N_4484,N_2688,N_773);
or U4485 (N_4485,N_3165,N_120);
nor U4486 (N_4486,N_1103,N_145);
or U4487 (N_4487,N_1312,N_230);
xnor U4488 (N_4488,N_2141,N_1731);
and U4489 (N_4489,N_615,N_371);
nor U4490 (N_4490,N_2531,N_2046);
nor U4491 (N_4491,N_3076,N_1606);
xor U4492 (N_4492,N_1773,N_2745);
or U4493 (N_4493,N_3476,N_3385);
nand U4494 (N_4494,N_1346,N_1291);
nor U4495 (N_4495,N_2795,N_90);
nor U4496 (N_4496,N_2404,N_836);
nor U4497 (N_4497,N_1031,N_677);
nor U4498 (N_4498,N_3509,N_3962);
and U4499 (N_4499,N_209,N_761);
or U4500 (N_4500,N_1214,N_1298);
and U4501 (N_4501,N_2109,N_3323);
nand U4502 (N_4502,N_3204,N_637);
or U4503 (N_4503,N_3973,N_1611);
nor U4504 (N_4504,N_1761,N_2463);
or U4505 (N_4505,N_1381,N_3695);
and U4506 (N_4506,N_1634,N_2723);
or U4507 (N_4507,N_3713,N_1335);
and U4508 (N_4508,N_2825,N_1119);
or U4509 (N_4509,N_3556,N_1977);
nand U4510 (N_4510,N_453,N_983);
nor U4511 (N_4511,N_1002,N_595);
xor U4512 (N_4512,N_2572,N_1210);
or U4513 (N_4513,N_278,N_2601);
nand U4514 (N_4514,N_1841,N_1290);
or U4515 (N_4515,N_721,N_1609);
xnor U4516 (N_4516,N_2714,N_1691);
nand U4517 (N_4517,N_952,N_222);
and U4518 (N_4518,N_2815,N_3008);
or U4519 (N_4519,N_3537,N_3031);
or U4520 (N_4520,N_242,N_1903);
and U4521 (N_4521,N_3969,N_1016);
nor U4522 (N_4522,N_487,N_3706);
nand U4523 (N_4523,N_2887,N_2385);
and U4524 (N_4524,N_935,N_2980);
nor U4525 (N_4525,N_3533,N_1647);
or U4526 (N_4526,N_656,N_3241);
xor U4527 (N_4527,N_2456,N_3025);
nand U4528 (N_4528,N_1380,N_748);
and U4529 (N_4529,N_3874,N_3338);
or U4530 (N_4530,N_2364,N_1915);
nor U4531 (N_4531,N_3180,N_682);
or U4532 (N_4532,N_39,N_797);
or U4533 (N_4533,N_2342,N_593);
or U4534 (N_4534,N_447,N_3586);
nand U4535 (N_4535,N_945,N_3273);
or U4536 (N_4536,N_3714,N_2291);
or U4537 (N_4537,N_695,N_200);
nor U4538 (N_4538,N_3668,N_2125);
nand U4539 (N_4539,N_3882,N_1207);
or U4540 (N_4540,N_264,N_2108);
nor U4541 (N_4541,N_3329,N_2803);
xnor U4542 (N_4542,N_2963,N_2682);
or U4543 (N_4543,N_2719,N_2660);
or U4544 (N_4544,N_415,N_2119);
nand U4545 (N_4545,N_2724,N_1234);
or U4546 (N_4546,N_2493,N_3489);
nor U4547 (N_4547,N_752,N_901);
nand U4548 (N_4548,N_3085,N_1805);
nor U4549 (N_4549,N_846,N_1395);
and U4550 (N_4550,N_2294,N_3665);
nor U4551 (N_4551,N_560,N_330);
xnor U4552 (N_4552,N_217,N_1345);
nor U4553 (N_4553,N_3207,N_668);
xor U4554 (N_4554,N_186,N_3809);
and U4555 (N_4555,N_1090,N_1833);
xnor U4556 (N_4556,N_1621,N_235);
and U4557 (N_4557,N_884,N_3391);
or U4558 (N_4558,N_472,N_396);
nand U4559 (N_4559,N_3555,N_1519);
or U4560 (N_4560,N_1158,N_2355);
and U4561 (N_4561,N_517,N_431);
nand U4562 (N_4562,N_72,N_1942);
nand U4563 (N_4563,N_404,N_2538);
nor U4564 (N_4564,N_1240,N_2098);
or U4565 (N_4565,N_515,N_2154);
or U4566 (N_4566,N_1798,N_199);
nand U4567 (N_4567,N_324,N_718);
nand U4568 (N_4568,N_2910,N_167);
nor U4569 (N_4569,N_1339,N_1715);
xnor U4570 (N_4570,N_3463,N_1849);
nand U4571 (N_4571,N_378,N_1173);
nor U4572 (N_4572,N_114,N_251);
nor U4573 (N_4573,N_694,N_2096);
nor U4574 (N_4574,N_800,N_1939);
nor U4575 (N_4575,N_3233,N_3474);
nand U4576 (N_4576,N_2590,N_3774);
nor U4577 (N_4577,N_3749,N_20);
nand U4578 (N_4578,N_2854,N_269);
nor U4579 (N_4579,N_2004,N_2525);
or U4580 (N_4580,N_2934,N_1073);
nand U4581 (N_4581,N_1535,N_2769);
or U4582 (N_4582,N_3811,N_3998);
xnor U4583 (N_4583,N_182,N_417);
or U4584 (N_4584,N_1607,N_3549);
nand U4585 (N_4585,N_2622,N_3720);
nand U4586 (N_4586,N_3742,N_1079);
nor U4587 (N_4587,N_1009,N_3778);
nand U4588 (N_4588,N_2262,N_3607);
xnor U4589 (N_4589,N_1088,N_2792);
nor U4590 (N_4590,N_1309,N_1809);
nand U4591 (N_4591,N_2904,N_2295);
and U4592 (N_4592,N_1772,N_3127);
or U4593 (N_4593,N_1993,N_2358);
nand U4594 (N_4594,N_3956,N_3627);
nor U4595 (N_4595,N_2085,N_3664);
or U4596 (N_4596,N_3693,N_491);
and U4597 (N_4597,N_2267,N_2307);
and U4598 (N_4598,N_439,N_3865);
nor U4599 (N_4599,N_1548,N_1674);
nand U4600 (N_4600,N_489,N_1402);
nor U4601 (N_4601,N_287,N_2530);
and U4602 (N_4602,N_3481,N_1136);
nand U4603 (N_4603,N_386,N_3853);
or U4604 (N_4604,N_1811,N_2681);
nor U4605 (N_4605,N_1971,N_1064);
nor U4606 (N_4606,N_1657,N_2293);
and U4607 (N_4607,N_2102,N_1039);
nand U4608 (N_4608,N_1361,N_3296);
and U4609 (N_4609,N_1810,N_3936);
and U4610 (N_4610,N_3258,N_1011);
nand U4611 (N_4611,N_1169,N_725);
nor U4612 (N_4612,N_2383,N_3154);
xnor U4613 (N_4613,N_3892,N_3903);
or U4614 (N_4614,N_547,N_626);
and U4615 (N_4615,N_2898,N_1319);
or U4616 (N_4616,N_1245,N_1153);
nor U4617 (N_4617,N_1209,N_1150);
nor U4618 (N_4618,N_435,N_232);
xor U4619 (N_4619,N_1506,N_2219);
and U4620 (N_4620,N_1024,N_3372);
xnor U4621 (N_4621,N_535,N_2159);
nor U4622 (N_4622,N_831,N_362);
nor U4623 (N_4623,N_3821,N_2517);
and U4624 (N_4624,N_3164,N_3926);
nor U4625 (N_4625,N_2401,N_1457);
and U4626 (N_4626,N_161,N_1850);
nand U4627 (N_4627,N_3729,N_3221);
nand U4628 (N_4628,N_889,N_795);
nand U4629 (N_4629,N_3646,N_1690);
nor U4630 (N_4630,N_1644,N_342);
or U4631 (N_4631,N_566,N_3839);
and U4632 (N_4632,N_1655,N_1321);
and U4633 (N_4633,N_2416,N_550);
nor U4634 (N_4634,N_1542,N_1973);
nand U4635 (N_4635,N_1521,N_2029);
nor U4636 (N_4636,N_3253,N_2505);
and U4637 (N_4637,N_657,N_108);
nor U4638 (N_4638,N_2189,N_2180);
and U4639 (N_4639,N_2373,N_316);
or U4640 (N_4640,N_3769,N_3242);
nor U4641 (N_4641,N_274,N_2121);
or U4642 (N_4642,N_587,N_3021);
nor U4643 (N_4643,N_353,N_3902);
or U4644 (N_4644,N_3029,N_2394);
nand U4645 (N_4645,N_2565,N_3129);
or U4646 (N_4646,N_706,N_1126);
or U4647 (N_4647,N_548,N_3197);
or U4648 (N_4648,N_1510,N_3675);
or U4649 (N_4649,N_2646,N_1351);
and U4650 (N_4650,N_84,N_591);
nand U4651 (N_4651,N_1446,N_2678);
and U4652 (N_4652,N_1174,N_1877);
and U4653 (N_4653,N_1985,N_2690);
nand U4654 (N_4654,N_1084,N_2658);
and U4655 (N_4655,N_1334,N_2179);
nor U4656 (N_4656,N_3857,N_2243);
and U4657 (N_4657,N_1425,N_2648);
nor U4658 (N_4658,N_1534,N_379);
xnor U4659 (N_4659,N_3744,N_1749);
nand U4660 (N_4660,N_3711,N_1721);
nand U4661 (N_4661,N_956,N_873);
and U4662 (N_4662,N_3935,N_2668);
or U4663 (N_4663,N_3433,N_3964);
and U4664 (N_4664,N_850,N_2780);
nand U4665 (N_4665,N_2516,N_966);
nor U4666 (N_4666,N_55,N_2952);
or U4667 (N_4667,N_988,N_1516);
nor U4668 (N_4668,N_630,N_2406);
and U4669 (N_4669,N_2720,N_1750);
nand U4670 (N_4670,N_62,N_3232);
or U4671 (N_4671,N_2712,N_1706);
or U4672 (N_4672,N_2876,N_733);
or U4673 (N_4673,N_127,N_3348);
and U4674 (N_4674,N_1897,N_2691);
nor U4675 (N_4675,N_2353,N_904);
or U4676 (N_4676,N_621,N_41);
nand U4677 (N_4677,N_878,N_845);
nor U4678 (N_4678,N_2909,N_1397);
nand U4679 (N_4679,N_937,N_1329);
and U4680 (N_4680,N_2286,N_3488);
nand U4681 (N_4681,N_231,N_728);
and U4682 (N_4682,N_2200,N_3885);
nand U4683 (N_4683,N_421,N_2031);
nand U4684 (N_4684,N_3098,N_2947);
or U4685 (N_4685,N_2563,N_19);
or U4686 (N_4686,N_3741,N_56);
and U4687 (N_4687,N_3443,N_1664);
nand U4688 (N_4688,N_1566,N_2184);
or U4689 (N_4689,N_929,N_3396);
and U4690 (N_4690,N_2773,N_1736);
and U4691 (N_4691,N_162,N_786);
or U4692 (N_4692,N_1701,N_147);
and U4693 (N_4693,N_3694,N_483);
or U4694 (N_4694,N_533,N_1753);
and U4695 (N_4695,N_2755,N_2124);
nand U4696 (N_4696,N_3168,N_1448);
nand U4697 (N_4697,N_1752,N_2454);
and U4698 (N_4698,N_1367,N_2916);
or U4699 (N_4699,N_14,N_796);
or U4700 (N_4700,N_2624,N_2984);
or U4701 (N_4701,N_3805,N_1763);
and U4702 (N_4702,N_1601,N_2834);
nor U4703 (N_4703,N_2703,N_2644);
or U4704 (N_4704,N_1999,N_1023);
or U4705 (N_4705,N_383,N_1597);
nand U4706 (N_4706,N_3986,N_1697);
nand U4707 (N_4707,N_859,N_2300);
and U4708 (N_4708,N_1879,N_3633);
xnor U4709 (N_4709,N_493,N_1976);
and U4710 (N_4710,N_1422,N_3542);
nand U4711 (N_4711,N_649,N_3947);
and U4712 (N_4712,N_1020,N_3125);
nor U4713 (N_4713,N_881,N_1594);
or U4714 (N_4714,N_3465,N_2882);
nand U4715 (N_4715,N_1124,N_1878);
or U4716 (N_4716,N_739,N_3457);
xnor U4717 (N_4717,N_1198,N_769);
and U4718 (N_4718,N_1503,N_448);
and U4719 (N_4719,N_3636,N_2245);
xor U4720 (N_4720,N_3037,N_1369);
and U4721 (N_4721,N_3032,N_3678);
nand U4722 (N_4722,N_49,N_1354);
nor U4723 (N_4723,N_2911,N_3126);
or U4724 (N_4724,N_3386,N_2640);
or U4725 (N_4725,N_1414,N_2941);
xor U4726 (N_4726,N_3785,N_1109);
nor U4727 (N_4727,N_2317,N_573);
nor U4728 (N_4728,N_2519,N_2570);
or U4729 (N_4729,N_808,N_468);
and U4730 (N_4730,N_47,N_420);
xor U4731 (N_4731,N_3813,N_3594);
or U4732 (N_4732,N_2327,N_3403);
nand U4733 (N_4733,N_3295,N_2479);
nand U4734 (N_4734,N_1447,N_2924);
or U4735 (N_4735,N_3344,N_3449);
and U4736 (N_4736,N_3112,N_3584);
or U4737 (N_4737,N_2228,N_3771);
nand U4738 (N_4738,N_2115,N_1757);
and U4739 (N_4739,N_531,N_1910);
nand U4740 (N_4740,N_1187,N_218);
nor U4741 (N_4741,N_2027,N_2339);
or U4742 (N_4742,N_2744,N_2178);
xor U4743 (N_4743,N_692,N_2459);
or U4744 (N_4744,N_1642,N_2628);
xor U4745 (N_4745,N_1531,N_3610);
and U4746 (N_4746,N_2430,N_3884);
nand U4747 (N_4747,N_3381,N_1863);
nor U4748 (N_4748,N_674,N_1949);
nand U4749 (N_4749,N_713,N_2101);
nand U4750 (N_4750,N_1202,N_2213);
or U4751 (N_4751,N_1912,N_651);
and U4752 (N_4752,N_3030,N_3376);
nand U4753 (N_4753,N_975,N_3161);
nor U4754 (N_4754,N_3366,N_734);
nand U4755 (N_4755,N_3442,N_1917);
and U4756 (N_4756,N_2354,N_1569);
nor U4757 (N_4757,N_2439,N_253);
nand U4758 (N_4758,N_1628,N_2861);
or U4759 (N_4759,N_3591,N_1686);
and U4760 (N_4760,N_2529,N_2371);
nand U4761 (N_4761,N_2918,N_2960);
and U4762 (N_4762,N_3992,N_1028);
or U4763 (N_4763,N_1276,N_1211);
or U4764 (N_4764,N_2849,N_1870);
or U4765 (N_4765,N_2269,N_3409);
xnor U4766 (N_4766,N_3949,N_1680);
or U4767 (N_4767,N_1466,N_3353);
and U4768 (N_4768,N_3860,N_3343);
and U4769 (N_4769,N_3049,N_1137);
and U4770 (N_4770,N_3113,N_2276);
or U4771 (N_4771,N_3674,N_2398);
nand U4772 (N_4772,N_840,N_2789);
nand U4773 (N_4773,N_3500,N_2362);
and U4774 (N_4774,N_2235,N_394);
xnor U4775 (N_4775,N_1554,N_3099);
or U4776 (N_4776,N_2986,N_624);
xor U4777 (N_4777,N_2791,N_2313);
or U4778 (N_4778,N_3446,N_985);
nor U4779 (N_4779,N_3851,N_2133);
and U4780 (N_4780,N_3156,N_358);
and U4781 (N_4781,N_1091,N_1376);
nand U4782 (N_4782,N_2094,N_1862);
or U4783 (N_4783,N_938,N_1935);
nand U4784 (N_4784,N_2043,N_1630);
and U4785 (N_4785,N_3105,N_3520);
and U4786 (N_4786,N_508,N_2515);
nand U4787 (N_4787,N_2638,N_664);
and U4788 (N_4788,N_2686,N_736);
or U4789 (N_4789,N_518,N_1410);
nor U4790 (N_4790,N_3893,N_912);
or U4791 (N_4791,N_2066,N_2310);
nor U4792 (N_4792,N_2973,N_2040);
and U4793 (N_4793,N_3411,N_883);
nand U4794 (N_4794,N_1926,N_3349);
nand U4795 (N_4795,N_3408,N_2829);
nor U4796 (N_4796,N_148,N_3977);
nor U4797 (N_4797,N_2392,N_2057);
and U4798 (N_4798,N_2024,N_3176);
nor U4799 (N_4799,N_2363,N_1632);
and U4800 (N_4800,N_568,N_3760);
and U4801 (N_4801,N_1758,N_747);
nand U4802 (N_4802,N_2766,N_3731);
nor U4803 (N_4803,N_1217,N_2442);
and U4804 (N_4804,N_1005,N_142);
nor U4805 (N_4805,N_1522,N_3667);
or U4806 (N_4806,N_900,N_2793);
xnor U4807 (N_4807,N_2192,N_1471);
or U4808 (N_4808,N_986,N_549);
nand U4809 (N_4809,N_1099,N_347);
xor U4810 (N_4810,N_1383,N_2048);
or U4811 (N_4811,N_1762,N_868);
xnor U4812 (N_4812,N_3455,N_1561);
nor U4813 (N_4813,N_3093,N_3181);
and U4814 (N_4814,N_659,N_667);
nor U4815 (N_4815,N_2605,N_3788);
and U4816 (N_4816,N_2238,N_1702);
xnor U4817 (N_4817,N_3394,N_2080);
and U4818 (N_4818,N_2808,N_481);
or U4819 (N_4819,N_2280,N_326);
and U4820 (N_4820,N_1195,N_1026);
nor U4821 (N_4821,N_2303,N_2702);
nor U4822 (N_4822,N_3942,N_3854);
nor U4823 (N_4823,N_860,N_1145);
or U4824 (N_4824,N_2751,N_3522);
nor U4825 (N_4825,N_3958,N_1316);
and U4826 (N_4826,N_1356,N_1387);
and U4827 (N_4827,N_3057,N_559);
nand U4828 (N_4828,N_3782,N_1525);
or U4829 (N_4829,N_2649,N_3038);
xor U4830 (N_4830,N_3224,N_1848);
and U4831 (N_4831,N_2246,N_325);
xor U4832 (N_4832,N_790,N_2270);
and U4833 (N_4833,N_3439,N_648);
nand U4834 (N_4834,N_3279,N_78);
nor U4835 (N_4835,N_1567,N_3222);
nand U4836 (N_4836,N_971,N_2117);
xnor U4837 (N_4837,N_2095,N_440);
and U4838 (N_4838,N_1452,N_2676);
and U4839 (N_4839,N_118,N_1799);
nand U4840 (N_4840,N_1004,N_2143);
nand U4841 (N_4841,N_249,N_240);
and U4842 (N_4842,N_2618,N_1825);
nor U4843 (N_4843,N_2177,N_920);
or U4844 (N_4844,N_532,N_3918);
or U4845 (N_4845,N_2917,N_488);
nor U4846 (N_4846,N_1779,N_1006);
or U4847 (N_4847,N_3471,N_1843);
or U4848 (N_4848,N_3575,N_3723);
or U4849 (N_4849,N_2452,N_180);
or U4850 (N_4850,N_2062,N_3708);
nor U4851 (N_4851,N_132,N_3327);
nor U4852 (N_4852,N_1434,N_3562);
and U4853 (N_4853,N_261,N_2330);
nor U4854 (N_4854,N_3309,N_3531);
nand U4855 (N_4855,N_1238,N_1190);
or U4856 (N_4856,N_1152,N_3445);
nand U4857 (N_4857,N_2278,N_1203);
and U4858 (N_4858,N_3814,N_2908);
nand U4859 (N_4859,N_1572,N_1287);
nand U4860 (N_4860,N_3519,N_1544);
or U4861 (N_4861,N_307,N_1933);
nor U4862 (N_4862,N_1957,N_322);
nand U4863 (N_4863,N_1042,N_311);
or U4864 (N_4864,N_2784,N_3648);
and U4865 (N_4865,N_693,N_1436);
and U4866 (N_4866,N_1698,N_1123);
and U4867 (N_4867,N_281,N_422);
and U4868 (N_4868,N_1627,N_918);
nor U4869 (N_4869,N_1420,N_2839);
and U4870 (N_4870,N_1666,N_1001);
nor U4871 (N_4871,N_1740,N_2894);
and U4872 (N_4872,N_3950,N_2972);
or U4873 (N_4873,N_3035,N_3189);
or U4874 (N_4874,N_1305,N_818);
or U4875 (N_4875,N_2739,N_302);
nand U4876 (N_4876,N_623,N_1874);
nor U4877 (N_4877,N_238,N_373);
nand U4878 (N_4878,N_3585,N_3803);
nand U4879 (N_4879,N_76,N_638);
nand U4880 (N_4880,N_2597,N_2734);
xnor U4881 (N_4881,N_2845,N_2224);
and U4882 (N_4882,N_3661,N_3762);
or U4883 (N_4883,N_1160,N_2743);
or U4884 (N_4884,N_3553,N_3373);
and U4885 (N_4885,N_1048,N_581);
nor U4886 (N_4886,N_2609,N_1017);
nor U4887 (N_4887,N_2948,N_3768);
nor U4888 (N_4888,N_3579,N_3046);
or U4889 (N_4889,N_1128,N_2592);
or U4890 (N_4890,N_2555,N_3362);
and U4891 (N_4891,N_2473,N_1483);
nand U4892 (N_4892,N_3828,N_1895);
nor U4893 (N_4893,N_3185,N_2770);
and U4894 (N_4894,N_3196,N_125);
and U4895 (N_4895,N_1390,N_785);
xnor U4896 (N_4896,N_2933,N_267);
and U4897 (N_4897,N_3831,N_3932);
nor U4898 (N_4898,N_1479,N_1689);
nand U4899 (N_4899,N_2966,N_2762);
nor U4900 (N_4900,N_2397,N_1941);
nand U4901 (N_4901,N_387,N_3291);
and U4902 (N_4902,N_2462,N_2715);
nor U4903 (N_4903,N_228,N_950);
nor U4904 (N_4904,N_509,N_188);
nor U4905 (N_4905,N_2606,N_2457);
or U4906 (N_4906,N_2633,N_1308);
and U4907 (N_4907,N_3680,N_506);
nand U4908 (N_4908,N_1948,N_2764);
and U4909 (N_4909,N_1726,N_257);
nor U4910 (N_4910,N_3420,N_3848);
nor U4911 (N_4911,N_2170,N_3833);
nor U4912 (N_4912,N_1992,N_812);
nor U4913 (N_4913,N_2130,N_185);
and U4914 (N_4914,N_750,N_1708);
and U4915 (N_4915,N_1696,N_2814);
and U4916 (N_4916,N_3605,N_926);
and U4917 (N_4917,N_3157,N_828);
or U4918 (N_4918,N_3734,N_2477);
nand U4919 (N_4919,N_2340,N_1744);
and U4920 (N_4920,N_2836,N_3640);
and U4921 (N_4921,N_2907,N_3131);
or U4922 (N_4922,N_2116,N_2994);
nand U4923 (N_4923,N_866,N_1465);
and U4924 (N_4924,N_2082,N_381);
or U4925 (N_4925,N_1237,N_3004);
and U4926 (N_4926,N_1788,N_3756);
or U4927 (N_4927,N_2533,N_2632);
nand U4928 (N_4928,N_3178,N_1228);
nor U4929 (N_4929,N_2257,N_3173);
or U4930 (N_4930,N_601,N_1301);
and U4931 (N_4931,N_792,N_844);
nor U4932 (N_4932,N_2407,N_3387);
and U4933 (N_4933,N_1596,N_2078);
nor U4934 (N_4934,N_697,N_2153);
and U4935 (N_4935,N_3896,N_2567);
or U4936 (N_4936,N_475,N_2301);
nand U4937 (N_4937,N_523,N_3000);
nand U4938 (N_4938,N_3626,N_1030);
and U4939 (N_4939,N_2513,N_2482);
nor U4940 (N_4940,N_1315,N_1498);
and U4941 (N_4941,N_2441,N_3535);
nor U4942 (N_4942,N_979,N_29);
nand U4943 (N_4943,N_3612,N_1925);
or U4944 (N_4944,N_3497,N_67);
and U4945 (N_4945,N_1866,N_856);
xnor U4946 (N_4946,N_3975,N_1918);
nand U4947 (N_4947,N_2704,N_3143);
nand U4948 (N_4948,N_3361,N_3581);
nor U4949 (N_4949,N_1450,N_2883);
nand U4950 (N_4950,N_345,N_1861);
xor U4951 (N_4951,N_46,N_882);
nand U4952 (N_4952,N_3050,N_3288);
or U4953 (N_4953,N_3464,N_3430);
nand U4954 (N_4954,N_3727,N_2964);
and U4955 (N_4955,N_1827,N_1692);
and U4956 (N_4956,N_1787,N_597);
nand U4957 (N_4957,N_1998,N_370);
or U4958 (N_4958,N_2204,N_356);
nand U4959 (N_4959,N_622,N_3053);
nand U4960 (N_4960,N_3862,N_776);
xor U4961 (N_4961,N_2840,N_685);
and U4962 (N_4962,N_3166,N_2607);
and U4963 (N_4963,N_1343,N_2099);
nand U4964 (N_4964,N_1400,N_3159);
nand U4965 (N_4965,N_3595,N_3504);
nand U4966 (N_4966,N_1058,N_737);
and U4967 (N_4967,N_3067,N_272);
nor U4968 (N_4968,N_1248,N_2903);
nand U4969 (N_4969,N_545,N_2038);
nor U4970 (N_4970,N_578,N_425);
nor U4971 (N_4971,N_1770,N_3933);
xnor U4972 (N_4972,N_2022,N_2020);
or U4973 (N_4973,N_3569,N_3781);
and U4974 (N_4974,N_3392,N_1451);
or U4975 (N_4975,N_1204,N_2575);
nand U4976 (N_4976,N_987,N_424);
xnor U4977 (N_4977,N_925,N_1464);
or U4978 (N_4978,N_2104,N_1764);
and U4979 (N_4979,N_3,N_2852);
or U4980 (N_4980,N_1979,N_250);
xor U4981 (N_4981,N_3841,N_2190);
and U4982 (N_4982,N_2625,N_63);
nand U4983 (N_4983,N_2232,N_1268);
or U4984 (N_4984,N_2241,N_1262);
nor U4985 (N_4985,N_3709,N_1443);
or U4986 (N_4986,N_616,N_1575);
nand U4987 (N_4987,N_2656,N_1629);
nand U4988 (N_4988,N_1122,N_1493);
nor U4989 (N_4989,N_3090,N_2799);
nand U4990 (N_4990,N_3906,N_852);
nor U4991 (N_4991,N_1328,N_3247);
or U4992 (N_4992,N_1964,N_3191);
or U4993 (N_4993,N_3086,N_3516);
or U4994 (N_4994,N_726,N_2251);
or U4995 (N_4995,N_2786,N_1481);
and U4996 (N_4996,N_3529,N_715);
and U4997 (N_4997,N_2326,N_3460);
nor U4998 (N_4998,N_2729,N_1723);
or U4999 (N_4999,N_2319,N_2328);
nor U5000 (N_5000,N_1526,N_1653);
nand U5001 (N_5001,N_2578,N_830);
and U5002 (N_5002,N_3970,N_3939);
nor U5003 (N_5003,N_2015,N_3600);
or U5004 (N_5004,N_1796,N_3334);
or U5005 (N_5005,N_2598,N_1325);
or U5006 (N_5006,N_1759,N_1053);
xnor U5007 (N_5007,N_2938,N_3700);
or U5008 (N_5008,N_2831,N_708);
or U5009 (N_5009,N_2305,N_3512);
and U5010 (N_5010,N_2127,N_2777);
nor U5011 (N_5011,N_2215,N_3940);
nor U5012 (N_5012,N_2336,N_2979);
nor U5013 (N_5013,N_1658,N_337);
nor U5014 (N_5014,N_1304,N_951);
xnor U5015 (N_5015,N_789,N_3508);
and U5016 (N_5016,N_1360,N_258);
nor U5017 (N_5017,N_1035,N_2321);
or U5018 (N_5018,N_2011,N_2059);
nand U5019 (N_5019,N_1867,N_3899);
nor U5020 (N_5020,N_1370,N_143);
nand U5021 (N_5021,N_1789,N_3134);
nand U5022 (N_5022,N_2725,N_476);
xnor U5023 (N_5023,N_2138,N_1093);
nor U5024 (N_5024,N_574,N_2174);
and U5025 (N_5025,N_1440,N_2534);
or U5026 (N_5026,N_3437,N_2868);
and U5027 (N_5027,N_1755,N_778);
nand U5028 (N_5028,N_2069,N_2496);
or U5029 (N_5029,N_2122,N_1222);
nand U5030 (N_5030,N_1931,N_2835);
and U5031 (N_5031,N_1616,N_426);
nand U5032 (N_5032,N_933,N_2137);
nor U5033 (N_5033,N_466,N_1477);
nand U5034 (N_5034,N_3072,N_661);
nand U5035 (N_5035,N_1154,N_3613);
nand U5036 (N_5036,N_2754,N_1449);
nor U5037 (N_5037,N_3766,N_1349);
or U5038 (N_5038,N_2940,N_331);
nor U5039 (N_5039,N_3701,N_3967);
or U5040 (N_5040,N_1765,N_3272);
nand U5041 (N_5041,N_3545,N_3238);
nor U5042 (N_5042,N_1131,N_1886);
or U5043 (N_5043,N_1940,N_469);
nand U5044 (N_5044,N_3682,N_3830);
nor U5045 (N_5045,N_3543,N_3194);
nand U5046 (N_5046,N_992,N_3573);
nor U5047 (N_5047,N_1140,N_2320);
nor U5048 (N_5048,N_825,N_1263);
xor U5049 (N_5049,N_1052,N_2680);
nor U5050 (N_5050,N_2685,N_1484);
and U5051 (N_5051,N_1059,N_700);
nand U5052 (N_5052,N_3483,N_226);
xnor U5053 (N_5053,N_53,N_427);
xor U5054 (N_5054,N_3907,N_3622);
xnor U5055 (N_5055,N_2891,N_1539);
nor U5056 (N_5056,N_764,N_397);
nor U5057 (N_5057,N_589,N_2561);
nand U5058 (N_5058,N_2541,N_3540);
nor U5059 (N_5059,N_643,N_1180);
or U5060 (N_5060,N_2809,N_152);
nand U5061 (N_5061,N_2225,N_2539);
nor U5062 (N_5062,N_2231,N_1962);
or U5063 (N_5063,N_513,N_1786);
or U5064 (N_5064,N_3660,N_2445);
nor U5065 (N_5065,N_3470,N_604);
or U5066 (N_5066,N_3115,N_1923);
and U5067 (N_5067,N_2888,N_1821);
and U5068 (N_5068,N_2332,N_1070);
nand U5069 (N_5069,N_897,N_3812);
or U5070 (N_5070,N_2428,N_40);
or U5071 (N_5071,N_460,N_3326);
nand U5072 (N_5072,N_1206,N_3055);
nand U5073 (N_5073,N_3316,N_2260);
nor U5074 (N_5074,N_3663,N_3628);
nand U5075 (N_5075,N_1930,N_2620);
and U5076 (N_5076,N_436,N_3802);
nor U5077 (N_5077,N_2526,N_1819);
nor U5078 (N_5078,N_2520,N_3624);
nor U5079 (N_5079,N_3402,N_2271);
nor U5080 (N_5080,N_3620,N_2171);
xnor U5081 (N_5081,N_819,N_3415);
xor U5082 (N_5082,N_519,N_3200);
nand U5083 (N_5083,N_1382,N_1475);
or U5084 (N_5084,N_564,N_760);
xor U5085 (N_5085,N_496,N_2185);
and U5086 (N_5086,N_849,N_1864);
and U5087 (N_5087,N_1038,N_2860);
nand U5088 (N_5088,N_2253,N_79);
or U5089 (N_5089,N_1114,N_1555);
and U5090 (N_5090,N_2797,N_3699);
nand U5091 (N_5091,N_2708,N_1142);
and U5092 (N_5092,N_2929,N_101);
xor U5093 (N_5093,N_2546,N_2881);
or U5094 (N_5094,N_3564,N_332);
nor U5095 (N_5095,N_2817,N_544);
or U5096 (N_5096,N_1950,N_879);
xor U5097 (N_5097,N_3399,N_921);
xor U5098 (N_5098,N_3697,N_9);
xnor U5099 (N_5099,N_1681,N_1292);
nand U5100 (N_5100,N_3274,N_1894);
and U5101 (N_5101,N_380,N_1743);
nand U5102 (N_5102,N_3900,N_2535);
nor U5103 (N_5103,N_742,N_3243);
nand U5104 (N_5104,N_2802,N_3466);
and U5105 (N_5105,N_2426,N_1856);
xor U5106 (N_5106,N_1212,N_3124);
and U5107 (N_5107,N_3823,N_3753);
or U5108 (N_5108,N_1080,N_781);
and U5109 (N_5109,N_3779,N_3816);
nand U5110 (N_5110,N_3369,N_3331);
nand U5111 (N_5111,N_927,N_3835);
nor U5112 (N_5112,N_2306,N_2557);
and U5113 (N_5113,N_3108,N_2510);
or U5114 (N_5114,N_2423,N_1055);
or U5115 (N_5115,N_1818,N_3917);
or U5116 (N_5116,N_3861,N_1730);
xor U5117 (N_5117,N_1232,N_2950);
xnor U5118 (N_5118,N_1802,N_59);
nand U5119 (N_5119,N_1394,N_323);
and U5120 (N_5120,N_3864,N_2939);
and U5121 (N_5121,N_977,N_2438);
or U5122 (N_5122,N_292,N_3759);
nor U5123 (N_5123,N_650,N_3643);
xnor U5124 (N_5124,N_2220,N_3226);
or U5125 (N_5125,N_467,N_2863);
or U5126 (N_5126,N_2054,N_297);
nand U5127 (N_5127,N_3960,N_2885);
and U5128 (N_5128,N_3669,N_1896);
nor U5129 (N_5129,N_2696,N_775);
nand U5130 (N_5130,N_313,N_2079);
nand U5131 (N_5131,N_312,N_482);
nor U5132 (N_5132,N_2372,N_2956);
or U5133 (N_5133,N_2569,N_416);
xnor U5134 (N_5134,N_86,N_2483);
nand U5135 (N_5135,N_1728,N_3240);
or U5136 (N_5136,N_1274,N_391);
and U5137 (N_5137,N_2995,N_2420);
nor U5138 (N_5138,N_1386,N_1748);
xor U5139 (N_5139,N_1784,N_3047);
or U5140 (N_5140,N_3208,N_1872);
and U5141 (N_5141,N_2056,N_1978);
and U5142 (N_5142,N_1956,N_3732);
nor U5143 (N_5143,N_2023,N_3109);
or U5144 (N_5144,N_767,N_2471);
nor U5145 (N_5145,N_2944,N_3916);
and U5146 (N_5146,N_83,N_221);
xnor U5147 (N_5147,N_1363,N_2164);
nand U5148 (N_5148,N_2169,N_3218);
and U5149 (N_5149,N_2647,N_390);
or U5150 (N_5150,N_1067,N_3364);
and U5151 (N_5151,N_3405,N_839);
nor U5152 (N_5152,N_2547,N_2866);
nor U5153 (N_5153,N_1082,N_2577);
or U5154 (N_5154,N_2440,N_2700);
nand U5155 (N_5155,N_1104,N_3752);
nand U5156 (N_5156,N_3048,N_429);
nor U5157 (N_5157,N_1983,N_914);
and U5158 (N_5158,N_3937,N_3120);
nand U5159 (N_5159,N_2965,N_1054);
nor U5160 (N_5160,N_2250,N_1108);
xor U5161 (N_5161,N_1270,N_2360);
nor U5162 (N_5162,N_2936,N_1433);
xor U5163 (N_5163,N_3991,N_3745);
and U5164 (N_5164,N_1501,N_3890);
nand U5165 (N_5165,N_1101,N_3728);
or U5166 (N_5166,N_65,N_3118);
or U5167 (N_5167,N_641,N_2413);
nor U5168 (N_5168,N_1795,N_71);
xor U5169 (N_5169,N_255,N_2752);
and U5170 (N_5170,N_2010,N_3155);
nor U5171 (N_5171,N_105,N_3171);
nand U5172 (N_5172,N_1560,N_1965);
nand U5173 (N_5173,N_1487,N_32);
or U5174 (N_5174,N_479,N_3249);
or U5175 (N_5175,N_3518,N_3615);
or U5176 (N_5176,N_1155,N_1144);
xnor U5177 (N_5177,N_582,N_848);
nor U5178 (N_5178,N_782,N_843);
and U5179 (N_5179,N_1358,N_3262);
nand U5180 (N_5180,N_1040,N_419);
xor U5181 (N_5181,N_2771,N_2599);
or U5182 (N_5182,N_305,N_2508);
and U5183 (N_5183,N_3284,N_1813);
nor U5184 (N_5184,N_3954,N_1570);
xor U5185 (N_5185,N_3491,N_3820);
nor U5186 (N_5186,N_2992,N_16);
nand U5187 (N_5187,N_965,N_857);
and U5188 (N_5188,N_3289,N_1066);
and U5189 (N_5189,N_1974,N_1224);
xor U5190 (N_5190,N_2198,N_3011);
or U5191 (N_5191,N_1105,N_3082);
or U5192 (N_5192,N_978,N_887);
and U5193 (N_5193,N_3148,N_2641);
or U5194 (N_5194,N_3485,N_527);
and U5195 (N_5195,N_1946,N_3868);
nand U5196 (N_5196,N_1660,N_3250);
and U5197 (N_5197,N_1437,N_2796);
or U5198 (N_5198,N_885,N_751);
xor U5199 (N_5199,N_3787,N_1938);
nand U5200 (N_5200,N_1125,N_3371);
xor U5201 (N_5201,N_1717,N_1828);
nor U5202 (N_5202,N_3280,N_2208);
and U5203 (N_5203,N_3789,N_2857);
nand U5204 (N_5204,N_1116,N_3310);
xnor U5205 (N_5205,N_45,N_3780);
or U5206 (N_5206,N_2501,N_24);
nor U5207 (N_5207,N_2985,N_1288);
nor U5208 (N_5208,N_3492,N_3685);
xnor U5209 (N_5209,N_740,N_1191);
xnor U5210 (N_5210,N_3432,N_1988);
or U5211 (N_5211,N_1552,N_3346);
or U5212 (N_5212,N_2429,N_777);
or U5213 (N_5213,N_1247,N_402);
and U5214 (N_5214,N_3206,N_3190);
and U5215 (N_5215,N_3077,N_2669);
xor U5216 (N_5216,N_3557,N_1505);
xor U5217 (N_5217,N_159,N_1565);
or U5218 (N_5218,N_3380,N_2186);
xnor U5219 (N_5219,N_68,N_3601);
nor U5220 (N_5220,N_1605,N_1598);
nand U5221 (N_5221,N_0,N_1472);
nand U5222 (N_5222,N_2236,N_503);
nor U5223 (N_5223,N_612,N_1278);
and U5224 (N_5224,N_3938,N_617);
nand U5225 (N_5225,N_239,N_1249);
or U5226 (N_5226,N_327,N_3946);
and U5227 (N_5227,N_3589,N_293);
or U5228 (N_5228,N_1508,N_1808);
nand U5229 (N_5229,N_2334,N_3418);
or U5230 (N_5230,N_3074,N_902);
and U5231 (N_5231,N_2400,N_1707);
xnor U5232 (N_5232,N_2954,N_3784);
nand U5233 (N_5233,N_3311,N_191);
nand U5234 (N_5234,N_2367,N_3149);
and U5235 (N_5235,N_1176,N_3919);
and U5236 (N_5236,N_194,N_1868);
and U5237 (N_5237,N_2450,N_1936);
nor U5238 (N_5238,N_1406,N_1391);
or U5239 (N_5239,N_3130,N_2937);
nand U5240 (N_5240,N_50,N_1987);
and U5241 (N_5241,N_3773,N_2047);
xnor U5242 (N_5242,N_709,N_524);
or U5243 (N_5243,N_400,N_2595);
nand U5244 (N_5244,N_2864,N_170);
or U5245 (N_5245,N_3652,N_2511);
and U5246 (N_5246,N_198,N_2637);
nand U5247 (N_5247,N_2412,N_684);
or U5248 (N_5248,N_1816,N_3453);
or U5249 (N_5249,N_3089,N_109);
nor U5250 (N_5250,N_2683,N_1139);
xnor U5251 (N_5251,N_1663,N_744);
nor U5252 (N_5252,N_3140,N_1172);
nor U5253 (N_5253,N_688,N_131);
or U5254 (N_5254,N_3826,N_1845);
or U5255 (N_5255,N_3653,N_1882);
and U5256 (N_5256,N_1549,N_3220);
nand U5257 (N_5257,N_660,N_1200);
nand U5258 (N_5258,N_3293,N_3388);
nand U5259 (N_5259,N_2717,N_23);
nor U5260 (N_5260,N_3393,N_909);
nand U5261 (N_5261,N_2014,N_5);
and U5262 (N_5262,N_33,N_2120);
or U5263 (N_5263,N_339,N_2001);
nand U5264 (N_5264,N_3152,N_2196);
or U5265 (N_5265,N_1913,N_1112);
nor U5266 (N_5266,N_3153,N_3541);
nand U5267 (N_5267,N_17,N_1751);
and U5268 (N_5268,N_1617,N_2478);
nor U5269 (N_5269,N_2399,N_522);
and U5270 (N_5270,N_554,N_2842);
and U5271 (N_5271,N_1817,N_85);
or U5272 (N_5272,N_2335,N_2626);
nor U5273 (N_5273,N_1582,N_865);
or U5274 (N_5274,N_3934,N_2932);
and U5275 (N_5275,N_37,N_3435);
nand U5276 (N_5276,N_2061,N_2757);
or U5277 (N_5277,N_571,N_498);
and U5278 (N_5278,N_3602,N_411);
and U5279 (N_5279,N_2843,N_1889);
nor U5280 (N_5280,N_552,N_2451);
nand U5281 (N_5281,N_219,N_3111);
and U5282 (N_5282,N_2384,N_497);
nand U5283 (N_5283,N_1844,N_2007);
nand U5284 (N_5284,N_1015,N_1201);
nand U5285 (N_5285,N_1218,N_1094);
or U5286 (N_5286,N_1196,N_2788);
or U5287 (N_5287,N_1348,N_1277);
or U5288 (N_5288,N_2727,N_3510);
or U5289 (N_5289,N_139,N_3187);
nand U5290 (N_5290,N_340,N_3501);
nor U5291 (N_5291,N_754,N_3507);
and U5292 (N_5292,N_1720,N_296);
and U5293 (N_5293,N_1254,N_2776);
nand U5294 (N_5294,N_724,N_1076);
and U5295 (N_5295,N_462,N_1610);
and U5296 (N_5296,N_299,N_2382);
and U5297 (N_5297,N_3498,N_891);
nand U5298 (N_5298,N_2277,N_2203);
nor U5299 (N_5299,N_2351,N_858);
nor U5300 (N_5300,N_2687,N_521);
nand U5301 (N_5301,N_3263,N_2136);
and U5302 (N_5302,N_1000,N_3578);
and U5303 (N_5303,N_557,N_2875);
nand U5304 (N_5304,N_3846,N_1086);
nor U5305 (N_5305,N_1700,N_495);
xor U5306 (N_5306,N_2273,N_2497);
or U5307 (N_5307,N_234,N_154);
and U5308 (N_5308,N_136,N_126);
or U5309 (N_5309,N_2163,N_1442);
nand U5310 (N_5310,N_3645,N_1602);
nand U5311 (N_5311,N_658,N_3687);
and U5312 (N_5312,N_2006,N_1562);
or U5313 (N_5313,N_1399,N_2156);
and U5314 (N_5314,N_1899,N_3978);
xnor U5315 (N_5315,N_3248,N_51);
or U5316 (N_5316,N_763,N_3795);
or U5317 (N_5317,N_36,N_3521);
and U5318 (N_5318,N_1463,N_3496);
and U5319 (N_5319,N_2021,N_1954);
or U5320 (N_5320,N_349,N_3469);
or U5321 (N_5321,N_2063,N_1595);
nand U5322 (N_5322,N_1904,N_3776);
nor U5323 (N_5323,N_2167,N_395);
nor U5324 (N_5324,N_2962,N_2114);
nand U5325 (N_5325,N_968,N_3012);
nor U5326 (N_5326,N_1194,N_2692);
nor U5327 (N_5327,N_304,N_205);
or U5328 (N_5328,N_160,N_2229);
or U5329 (N_5329,N_2655,N_245);
nand U5330 (N_5330,N_2709,N_1695);
nor U5331 (N_5331,N_727,N_1132);
nor U5332 (N_5332,N_801,N_1590);
or U5333 (N_5333,N_2586,N_1920);
nand U5334 (N_5334,N_2134,N_577);
nand U5335 (N_5335,N_1412,N_1742);
and U5336 (N_5336,N_3536,N_2090);
or U5337 (N_5337,N_2448,N_3634);
nand U5338 (N_5338,N_2958,N_2329);
nor U5339 (N_5339,N_2285,N_3302);
and U5340 (N_5340,N_936,N_262);
nor U5341 (N_5341,N_173,N_321);
or U5342 (N_5342,N_3429,N_247);
and U5343 (N_5343,N_3913,N_3654);
or U5344 (N_5344,N_2263,N_3761);
nor U5345 (N_5345,N_2494,N_719);
xnor U5346 (N_5346,N_3139,N_1143);
or U5347 (N_5347,N_665,N_1025);
and U5348 (N_5348,N_1512,N_1797);
nor U5349 (N_5349,N_1732,N_3867);
and U5350 (N_5350,N_18,N_2726);
xnor U5351 (N_5351,N_1636,N_2249);
xor U5352 (N_5352,N_575,N_3019);
nor U5353 (N_5353,N_2787,N_2967);
or U5354 (N_5354,N_3413,N_1342);
xnor U5355 (N_5355,N_1178,N_2585);
or U5356 (N_5356,N_1286,N_364);
xnor U5357 (N_5357,N_3436,N_97);
and U5358 (N_5358,N_1790,N_974);
nand U5359 (N_5359,N_1491,N_3002);
nand U5360 (N_5360,N_3270,N_2935);
nor U5361 (N_5361,N_567,N_2775);
nand U5362 (N_5362,N_924,N_286);
and U5363 (N_5363,N_163,N_2642);
nor U5364 (N_5364,N_679,N_3425);
nand U5365 (N_5365,N_1257,N_190);
nor U5366 (N_5366,N_783,N_1943);
and U5367 (N_5367,N_3877,N_1488);
xor U5368 (N_5368,N_3574,N_213);
and U5369 (N_5369,N_551,N_3806);
or U5370 (N_5370,N_2264,N_855);
nor U5371 (N_5371,N_1046,N_3551);
nand U5372 (N_5372,N_2673,N_1530);
and U5373 (N_5373,N_384,N_2255);
nor U5374 (N_5374,N_452,N_3658);
nand U5375 (N_5375,N_853,N_3524);
or U5376 (N_5376,N_1907,N_1485);
nor U5377 (N_5377,N_2032,N_3423);
or U5378 (N_5378,N_3365,N_2781);
nor U5379 (N_5379,N_1975,N_1688);
nor U5380 (N_5380,N_3716,N_2977);
nor U5381 (N_5381,N_3141,N_1888);
and U5382 (N_5382,N_2356,N_2149);
or U5383 (N_5383,N_1110,N_3945);
and U5384 (N_5384,N_1504,N_3339);
and U5385 (N_5385,N_2361,N_2614);
and U5386 (N_5386,N_2705,N_206);
and U5387 (N_5387,N_3767,N_814);
nand U5388 (N_5388,N_629,N_3502);
nor U5389 (N_5389,N_174,N_662);
nor U5390 (N_5390,N_3352,N_1261);
nand U5391 (N_5391,N_30,N_2556);
nor U5392 (N_5392,N_2711,N_2870);
or U5393 (N_5393,N_144,N_3849);
nand U5394 (N_5394,N_276,N_181);
or U5395 (N_5395,N_1029,N_3651);
nor U5396 (N_5396,N_88,N_1322);
nand U5397 (N_5397,N_3101,N_1571);
nor U5398 (N_5398,N_2343,N_1036);
or U5399 (N_5399,N_2837,N_2160);
nand U5400 (N_5400,N_592,N_3479);
nor U5401 (N_5401,N_1411,N_1033);
nand U5402 (N_5402,N_1168,N_3363);
and U5403 (N_5403,N_2193,N_542);
xor U5404 (N_5404,N_1908,N_3912);
or U5405 (N_5405,N_3818,N_1269);
or U5406 (N_5406,N_1756,N_3883);
nand U5407 (N_5407,N_3526,N_2258);
or U5408 (N_5408,N_2730,N_636);
nor U5409 (N_5409,N_187,N_294);
nor U5410 (N_5410,N_485,N_365);
and U5411 (N_5411,N_418,N_3448);
and U5412 (N_5412,N_3044,N_1937);
nand U5413 (N_5413,N_1364,N_3719);
nand U5414 (N_5414,N_463,N_993);
nor U5415 (N_5415,N_409,N_2664);
and U5416 (N_5416,N_3063,N_2209);
nor U5417 (N_5417,N_2800,N_1846);
or U5418 (N_5418,N_1306,N_2873);
nor U5419 (N_5419,N_3928,N_2969);
nand U5420 (N_5420,N_319,N_3340);
nor U5421 (N_5421,N_1184,N_3417);
nand U5422 (N_5422,N_3632,N_634);
and U5423 (N_5423,N_1838,N_3058);
nor U5424 (N_5424,N_610,N_504);
or U5425 (N_5425,N_2019,N_2237);
nand U5426 (N_5426,N_2283,N_1626);
nand U5427 (N_5427,N_310,N_3847);
or U5428 (N_5428,N_2811,N_2218);
nand U5429 (N_5429,N_179,N_165);
xnor U5430 (N_5430,N_959,N_3458);
nand U5431 (N_5431,N_82,N_2097);
nor U5432 (N_5432,N_1419,N_1135);
or U5433 (N_5433,N_3880,N_1747);
nor U5434 (N_5434,N_1355,N_2388);
or U5435 (N_5435,N_1043,N_3205);
xor U5436 (N_5436,N_3040,N_1323);
nand U5437 (N_5437,N_676,N_3216);
or U5438 (N_5438,N_3301,N_2783);
nand U5439 (N_5439,N_633,N_2600);
or U5440 (N_5440,N_1687,N_3319);
nand U5441 (N_5441,N_176,N_2671);
nor U5442 (N_5442,N_58,N_270);
and U5443 (N_5443,N_826,N_652);
and U5444 (N_5444,N_896,N_3228);
and U5445 (N_5445,N_3924,N_1639);
nor U5446 (N_5446,N_15,N_1146);
and U5447 (N_5447,N_361,N_3158);
or U5448 (N_5448,N_3617,N_291);
and U5449 (N_5449,N_355,N_3023);
and U5450 (N_5450,N_1293,N_2659);
and U5451 (N_5451,N_645,N_809);
or U5452 (N_5452,N_2464,N_3908);
or U5453 (N_5453,N_1313,N_3558);
nor U5454 (N_5454,N_1932,N_459);
or U5455 (N_5455,N_433,N_1991);
and U5456 (N_5456,N_2818,N_3703);
nor U5457 (N_5457,N_1887,N_903);
nor U5458 (N_5458,N_21,N_608);
xnor U5459 (N_5459,N_3666,N_3993);
or U5460 (N_5460,N_1259,N_2126);
nand U5461 (N_5461,N_2805,N_289);
and U5462 (N_5462,N_1592,N_3104);
nor U5463 (N_5463,N_1745,N_133);
or U5464 (N_5464,N_2749,N_98);
or U5465 (N_5465,N_2654,N_2188);
nand U5466 (N_5466,N_3791,N_3515);
nor U5467 (N_5467,N_1564,N_3829);
nand U5468 (N_5468,N_1830,N_2879);
xor U5469 (N_5469,N_2737,N_2906);
or U5470 (N_5470,N_3799,N_893);
or U5471 (N_5471,N_492,N_1167);
xor U5472 (N_5472,N_103,N_315);
and U5473 (N_5473,N_867,N_2140);
or U5474 (N_5474,N_3318,N_1589);
and U5475 (N_5475,N_3100,N_3342);
or U5476 (N_5476,N_607,N_2502);
nor U5477 (N_5477,N_1969,N_932);
nor U5478 (N_5478,N_1233,N_3961);
nor U5479 (N_5479,N_3815,N_2252);
xnor U5480 (N_5480,N_106,N_3770);
nand U5481 (N_5481,N_2222,N_3959);
nand U5482 (N_5482,N_1453,N_385);
or U5483 (N_5483,N_2760,N_768);
nor U5484 (N_5484,N_3036,N_484);
or U5485 (N_5485,N_3738,N_2299);
and U5486 (N_5486,N_2951,N_999);
nand U5487 (N_5487,N_430,N_3800);
nand U5488 (N_5488,N_445,N_3022);
and U5489 (N_5489,N_2112,N_2822);
xnor U5490 (N_5490,N_618,N_583);
nand U5491 (N_5491,N_3116,N_2044);
nor U5492 (N_5492,N_3621,N_3647);
nand U5493 (N_5493,N_500,N_271);
or U5494 (N_5494,N_2460,N_1834);
and U5495 (N_5495,N_3313,N_753);
xnor U5496 (N_5496,N_2552,N_2896);
xnor U5497 (N_5497,N_368,N_2173);
nor U5498 (N_5498,N_1384,N_3527);
nand U5499 (N_5499,N_972,N_561);
nor U5500 (N_5500,N_2304,N_2461);
and U5501 (N_5501,N_2009,N_2214);
or U5502 (N_5502,N_3045,N_3478);
or U5503 (N_5503,N_2191,N_1511);
xor U5504 (N_5504,N_576,N_2288);
or U5505 (N_5505,N_2848,N_1418);
or U5506 (N_5506,N_3676,N_1712);
xnor U5507 (N_5507,N_374,N_2844);
nor U5508 (N_5508,N_2748,N_949);
or U5509 (N_5509,N_1803,N_410);
or U5510 (N_5510,N_822,N_2899);
nand U5511 (N_5511,N_164,N_3588);
nor U5512 (N_5512,N_3061,N_2381);
or U5513 (N_5513,N_628,N_335);
and U5514 (N_5514,N_3688,N_749);
and U5515 (N_5515,N_3881,N_3644);
or U5516 (N_5516,N_2890,N_203);
and U5517 (N_5517,N_3513,N_3350);
and U5518 (N_5518,N_2651,N_406);
nor U5519 (N_5519,N_815,N_1649);
nand U5520 (N_5520,N_3493,N_3997);
or U5521 (N_5521,N_4,N_2990);
nand U5522 (N_5522,N_3401,N_153);
xor U5523 (N_5523,N_171,N_2553);
nor U5524 (N_5524,N_87,N_283);
nand U5525 (N_5525,N_3027,N_233);
and U5526 (N_5526,N_2302,N_3001);
nor U5527 (N_5527,N_2338,N_2424);
nor U5528 (N_5528,N_1638,N_100);
and U5529 (N_5529,N_3230,N_2435);
nor U5530 (N_5530,N_3901,N_3941);
or U5531 (N_5531,N_1682,N_295);
and U5532 (N_5532,N_2210,N_639);
xnor U5533 (N_5533,N_2706,N_473);
nand U5534 (N_5534,N_3424,N_3976);
nand U5535 (N_5535,N_1424,N_755);
xnor U5536 (N_5536,N_3596,N_1693);
and U5537 (N_5537,N_811,N_1407);
or U5538 (N_5538,N_2272,N_871);
or U5539 (N_5539,N_2380,N_1405);
xnor U5540 (N_5540,N_3138,N_1478);
or U5541 (N_5541,N_1458,N_1003);
or U5542 (N_5542,N_1496,N_864);
or U5543 (N_5543,N_70,N_3400);
nor U5544 (N_5544,N_1703,N_2550);
or U5545 (N_5545,N_2523,N_2296);
and U5546 (N_5546,N_461,N_2823);
or U5547 (N_5547,N_2419,N_2466);
and U5548 (N_5548,N_745,N_3878);
or U5549 (N_5549,N_303,N_3702);
nand U5550 (N_5550,N_300,N_3570);
nand U5551 (N_5551,N_2617,N_3133);
and U5552 (N_5552,N_2621,N_3801);
or U5553 (N_5553,N_3234,N_3426);
or U5554 (N_5554,N_3298,N_2774);
and U5555 (N_5555,N_201,N_922);
or U5556 (N_5556,N_3568,N_580);
or U5557 (N_5557,N_1545,N_268);
nor U5558 (N_5558,N_1022,N_735);
or U5559 (N_5559,N_2886,N_1578);
nor U5560 (N_5560,N_3028,N_3689);
and U5561 (N_5561,N_1462,N_2772);
nor U5562 (N_5562,N_3606,N_948);
and U5563 (N_5563,N_2390,N_1614);
nor U5564 (N_5564,N_280,N_691);
nor U5565 (N_5565,N_1018,N_957);
nand U5566 (N_5566,N_3566,N_2495);
or U5567 (N_5567,N_3692,N_81);
nor U5568 (N_5568,N_2611,N_635);
nand U5569 (N_5569,N_3333,N_2144);
and U5570 (N_5570,N_367,N_157);
nor U5571 (N_5571,N_2379,N_3254);
or U5572 (N_5572,N_2921,N_2767);
and U5573 (N_5573,N_207,N_3017);
nand U5574 (N_5574,N_3251,N_502);
and U5575 (N_5575,N_3530,N_1097);
xor U5576 (N_5576,N_1069,N_1826);
nor U5577 (N_5577,N_2982,N_2832);
or U5578 (N_5578,N_7,N_1250);
nand U5579 (N_5579,N_1541,N_11);
nor U5580 (N_5580,N_3123,N_2165);
and U5581 (N_5581,N_1741,N_787);
nand U5582 (N_5582,N_2414,N_393);
nand U5583 (N_5583,N_1047,N_1213);
nand U5584 (N_5584,N_3717,N_553);
nand U5585 (N_5585,N_1785,N_2315);
nand U5586 (N_5586,N_1230,N_75);
or U5587 (N_5587,N_66,N_3096);
nor U5588 (N_5588,N_953,N_3525);
or U5589 (N_5589,N_3209,N_3649);
nand U5590 (N_5590,N_2847,N_1737);
nor U5591 (N_5591,N_1423,N_2697);
nor U5592 (N_5592,N_1460,N_1223);
nand U5593 (N_5593,N_2089,N_3268);
and U5594 (N_5594,N_1326,N_3336);
xor U5595 (N_5595,N_964,N_3715);
nand U5596 (N_5596,N_928,N_351);
and U5597 (N_5597,N_963,N_3514);
nor U5598 (N_5598,N_92,N_600);
nor U5599 (N_5599,N_2425,N_1470);
and U5600 (N_5600,N_27,N_969);
or U5601 (N_5601,N_1710,N_1875);
nor U5602 (N_5602,N_343,N_1273);
nand U5603 (N_5603,N_1426,N_1855);
and U5604 (N_5604,N_707,N_2874);
and U5605 (N_5605,N_1807,N_1166);
nand U5606 (N_5606,N_3655,N_2884);
nand U5607 (N_5607,N_248,N_1480);
nand U5608 (N_5608,N_34,N_1428);
nand U5609 (N_5609,N_2281,N_285);
or U5610 (N_5610,N_1085,N_94);
or U5611 (N_5611,N_3604,N_947);
nand U5612 (N_5612,N_1643,N_2187);
xnor U5613 (N_5613,N_3657,N_3988);
and U5614 (N_5614,N_3822,N_1375);
and U5615 (N_5615,N_215,N_3088);
nand U5616 (N_5616,N_2779,N_538);
or U5617 (N_5617,N_2145,N_1295);
and U5618 (N_5618,N_2667,N_3972);
nor U5619 (N_5619,N_3982,N_723);
or U5620 (N_5620,N_2721,N_3375);
and U5621 (N_5621,N_3355,N_195);
or U5622 (N_5622,N_2604,N_260);
and U5623 (N_5623,N_510,N_3642);
or U5624 (N_5624,N_2548,N_3051);
or U5625 (N_5625,N_3544,N_2521);
xor U5626 (N_5626,N_1513,N_3808);
and U5627 (N_5627,N_514,N_943);
and U5628 (N_5628,N_2946,N_3246);
and U5629 (N_5629,N_3307,N_2701);
xor U5630 (N_5630,N_1951,N_3724);
nand U5631 (N_5631,N_1220,N_973);
and U5632 (N_5632,N_2807,N_1880);
xor U5633 (N_5633,N_2081,N_2514);
or U5634 (N_5634,N_130,N_540);
and U5635 (N_5635,N_741,N_3764);
and U5636 (N_5636,N_1403,N_1427);
nor U5637 (N_5637,N_1990,N_2376);
xnor U5638 (N_5638,N_3844,N_1373);
nor U5639 (N_5639,N_3144,N_2652);
nor U5640 (N_5640,N_2434,N_407);
or U5641 (N_5641,N_1533,N_3777);
or U5642 (N_5642,N_3656,N_2055);
or U5643 (N_5643,N_2999,N_1746);
xnor U5644 (N_5644,N_671,N_1229);
nor U5645 (N_5645,N_77,N_1883);
and U5646 (N_5646,N_833,N_2067);
xnor U5647 (N_5647,N_1615,N_2422);
nor U5648 (N_5648,N_2740,N_1959);
nand U5649 (N_5649,N_3069,N_1847);
nand U5650 (N_5650,N_54,N_3013);
nor U5651 (N_5651,N_3897,N_3751);
and U5652 (N_5652,N_1778,N_766);
nor U5653 (N_5653,N_1963,N_837);
nand U5654 (N_5654,N_290,N_1032);
nand U5655 (N_5655,N_1972,N_1853);
nor U5656 (N_5656,N_2183,N_1289);
and U5657 (N_5657,N_1008,N_3081);
and U5658 (N_5658,N_556,N_3018);
and U5659 (N_5659,N_2352,N_2503);
nor U5660 (N_5660,N_3245,N_2718);
nand U5661 (N_5661,N_3223,N_3684);
nand U5662 (N_5662,N_8,N_3389);
nand U5663 (N_5663,N_1118,N_3705);
or U5664 (N_5664,N_338,N_3303);
or U5665 (N_5665,N_329,N_1989);
nor U5666 (N_5666,N_2234,N_1944);
or U5667 (N_5667,N_3559,N_1704);
xor U5668 (N_5668,N_1631,N_80);
nor U5669 (N_5669,N_528,N_3505);
nand U5670 (N_5670,N_3229,N_3810);
xnor U5671 (N_5671,N_875,N_1619);
nand U5672 (N_5672,N_2446,N_2981);
nand U5673 (N_5673,N_1186,N_403);
and U5674 (N_5674,N_1536,N_2365);
or U5675 (N_5675,N_2763,N_1165);
nand U5676 (N_5676,N_3447,N_1581);
xor U5677 (N_5677,N_212,N_2901);
or U5678 (N_5678,N_1675,N_1806);
nor U5679 (N_5679,N_3552,N_2308);
nor U5680 (N_5680,N_2350,N_3856);
xor U5681 (N_5681,N_2324,N_1568);
xnor U5682 (N_5682,N_3629,N_1584);
and U5683 (N_5683,N_644,N_25);
and U5684 (N_5684,N_2226,N_1633);
nor U5685 (N_5685,N_1968,N_2733);
and U5686 (N_5686,N_1379,N_3213);
or U5687 (N_5687,N_3431,N_1556);
or U5688 (N_5688,N_2039,N_3726);
or U5689 (N_5689,N_3150,N_1063);
or U5690 (N_5690,N_3261,N_3354);
and U5691 (N_5691,N_1130,N_1282);
nand U5692 (N_5692,N_2804,N_2758);
and U5693 (N_5693,N_1668,N_2549);
or U5694 (N_5694,N_423,N_2074);
or U5695 (N_5695,N_141,N_1713);
nand U5696 (N_5696,N_1980,N_2491);
or U5697 (N_5697,N_2207,N_1791);
and U5698 (N_5698,N_1156,N_204);
nor U5699 (N_5699,N_412,N_2506);
and U5700 (N_5700,N_3260,N_3357);
and U5701 (N_5701,N_3132,N_817);
nand U5702 (N_5702,N_3565,N_458);
or U5703 (N_5703,N_3163,N_1768);
and U5704 (N_5704,N_780,N_3452);
and U5705 (N_5705,N_759,N_3266);
and U5706 (N_5706,N_1499,N_2518);
xor U5707 (N_5707,N_2175,N_2168);
nor U5708 (N_5708,N_2741,N_2974);
nor U5709 (N_5709,N_2265,N_178);
and U5710 (N_5710,N_2410,N_2961);
xor U5711 (N_5711,N_168,N_1179);
and U5712 (N_5712,N_3358,N_3146);
and U5713 (N_5713,N_3052,N_2086);
nor U5714 (N_5714,N_3952,N_408);
nand U5715 (N_5715,N_3974,N_3304);
and U5716 (N_5716,N_3459,N_1960);
or U5717 (N_5717,N_2431,N_1431);
xor U5718 (N_5718,N_1310,N_405);
or U5719 (N_5719,N_140,N_931);
and U5720 (N_5720,N_2507,N_1107);
nor U5721 (N_5721,N_3886,N_731);
and U5722 (N_5722,N_3807,N_2579);
xor U5723 (N_5723,N_2850,N_1637);
and U5724 (N_5724,N_1177,N_2274);
or U5725 (N_5725,N_1800,N_2323);
or U5726 (N_5726,N_3707,N_3231);
or U5727 (N_5727,N_2000,N_614);
nor U5728 (N_5728,N_2093,N_1051);
or U5729 (N_5729,N_3083,N_989);
nor U5730 (N_5730,N_3765,N_3062);
and U5731 (N_5731,N_3547,N_998);
xor U5732 (N_5732,N_1635,N_470);
nand U5733 (N_5733,N_1677,N_471);
and U5734 (N_5734,N_3244,N_3227);
and U5735 (N_5735,N_2417,N_813);
xnor U5736 (N_5736,N_1523,N_2551);
nor U5737 (N_5737,N_1837,N_1258);
xor U5738 (N_5738,N_1585,N_2853);
nand U5739 (N_5739,N_690,N_3635);
and U5740 (N_5740,N_2075,N_3075);
or U5741 (N_5741,N_1538,N_1235);
or U5742 (N_5742,N_1061,N_1303);
nor U5743 (N_5743,N_1,N_2532);
or U5744 (N_5744,N_401,N_678);
xor U5745 (N_5745,N_1591,N_1171);
and U5746 (N_5746,N_284,N_1835);
nor U5747 (N_5747,N_3461,N_3255);
and U5748 (N_5748,N_2790,N_1672);
and U5749 (N_5749,N_907,N_1891);
nor U5750 (N_5750,N_1149,N_237);
nand U5751 (N_5751,N_3368,N_2077);
nand U5752 (N_5752,N_91,N_1417);
nand U5753 (N_5753,N_2540,N_477);
nor U5754 (N_5754,N_3107,N_2824);
or U5755 (N_5755,N_1831,N_6);
nand U5756 (N_5756,N_1151,N_2666);
nand U5757 (N_5757,N_1705,N_3252);
and U5758 (N_5758,N_1718,N_1120);
nor U5759 (N_5759,N_2892,N_344);
nand U5760 (N_5760,N_505,N_2612);
or U5761 (N_5761,N_962,N_3577);
nor U5762 (N_5762,N_3332,N_456);
or U5763 (N_5763,N_3499,N_2033);
nand U5764 (N_5764,N_2661,N_1404);
xor U5765 (N_5765,N_3842,N_28);
nand U5766 (N_5766,N_1873,N_1163);
nand U5767 (N_5767,N_829,N_1729);
nand U5768 (N_5768,N_3014,N_1587);
or U5769 (N_5769,N_3414,N_282);
nand U5770 (N_5770,N_919,N_1547);
nand U5771 (N_5771,N_997,N_3638);
and U5772 (N_5772,N_1408,N_2747);
or U5773 (N_5773,N_1389,N_774);
or U5774 (N_5774,N_1294,N_2810);
or U5775 (N_5775,N_770,N_3421);
nand U5776 (N_5776,N_841,N_3641);
or U5777 (N_5777,N_3277,N_1733);
nor U5778 (N_5778,N_1330,N_1551);
nand U5779 (N_5779,N_1378,N_2211);
or U5780 (N_5780,N_701,N_3225);
nor U5781 (N_5781,N_3059,N_2865);
nand U5782 (N_5782,N_3944,N_3852);
or U5783 (N_5783,N_44,N_279);
or U5784 (N_5784,N_2663,N_3690);
nor U5785 (N_5785,N_1271,N_3438);
or U5786 (N_5786,N_2594,N_377);
and U5787 (N_5787,N_2105,N_880);
xor U5788 (N_5788,N_1858,N_107);
nand U5789 (N_5789,N_150,N_119);
nand U5790 (N_5790,N_1121,N_360);
nor U5791 (N_5791,N_3269,N_516);
or U5792 (N_5792,N_1267,N_2742);
xnor U5793 (N_5793,N_3202,N_980);
nor U5794 (N_5794,N_3121,N_2084);
nand U5795 (N_5795,N_2481,N_917);
or U5796 (N_5796,N_1347,N_862);
nor U5797 (N_5797,N_2282,N_2344);
nor U5798 (N_5798,N_1684,N_3845);
or U5799 (N_5799,N_3790,N_2103);
nand U5800 (N_5800,N_1645,N_3930);
nand U5801 (N_5801,N_1244,N_3772);
or U5802 (N_5802,N_2017,N_2110);
xor U5803 (N_5803,N_1885,N_52);
nor U5804 (N_5804,N_1253,N_3192);
xnor U5805 (N_5805,N_3487,N_710);
nor U5806 (N_5806,N_1092,N_1576);
nand U5807 (N_5807,N_1468,N_2333);
and U5808 (N_5808,N_558,N_1010);
nor U5809 (N_5809,N_541,N_2378);
and U5810 (N_5810,N_3580,N_716);
nor U5811 (N_5811,N_3995,N_705);
and U5812 (N_5812,N_687,N_3068);
nor U5813 (N_5813,N_2970,N_730);
or U5814 (N_5814,N_2922,N_2582);
or U5815 (N_5815,N_2558,N_1324);
or U5816 (N_5816,N_3136,N_3179);
or U5817 (N_5817,N_1189,N_1083);
and U5818 (N_5818,N_3312,N_3677);
xor U5819 (N_5819,N_1659,N_1901);
and U5820 (N_5820,N_3337,N_2139);
nor U5821 (N_5821,N_2665,N_3203);
nor U5822 (N_5822,N_3927,N_3511);
xor U5823 (N_5823,N_3743,N_3494);
or U5824 (N_5824,N_625,N_1893);
nor U5825 (N_5825,N_1766,N_1115);
or U5826 (N_5826,N_146,N_2761);
and U5827 (N_5827,N_252,N_2544);
and U5828 (N_5828,N_2368,N_1049);
and U5829 (N_5829,N_1905,N_1613);
or U5830 (N_5830,N_3872,N_3078);
nand U5831 (N_5831,N_2545,N_2949);
or U5832 (N_5832,N_655,N_1679);
and U5833 (N_5833,N_428,N_1284);
nor U5834 (N_5834,N_536,N_138);
nor U5835 (N_5835,N_1641,N_1661);
or U5836 (N_5836,N_2386,N_712);
nor U5837 (N_5837,N_602,N_96);
or U5838 (N_5838,N_683,N_193);
nor U5839 (N_5839,N_1398,N_3095);
or U5840 (N_5840,N_2284,N_2240);
nor U5841 (N_5841,N_1314,N_1444);
nor U5842 (N_5842,N_1106,N_38);
xnor U5843 (N_5843,N_2212,N_3374);
nor U5844 (N_5844,N_563,N_673);
or U5845 (N_5845,N_486,N_2498);
or U5846 (N_5846,N_611,N_3739);
nand U5847 (N_5847,N_2813,N_3910);
or U5848 (N_5848,N_3792,N_2602);
and U5849 (N_5849,N_2195,N_3416);
or U5850 (N_5850,N_3356,N_599);
and U5851 (N_5851,N_2472,N_352);
nor U5852 (N_5852,N_2794,N_1546);
nor U5853 (N_5853,N_2312,N_3999);
and U5854 (N_5854,N_1241,N_2639);
xnor U5855 (N_5855,N_1134,N_3482);
and U5856 (N_5856,N_2900,N_2635);
nand U5857 (N_5857,N_2629,N_1662);
or U5858 (N_5858,N_1769,N_1193);
nand U5859 (N_5859,N_1801,N_301);
or U5860 (N_5860,N_2041,N_1836);
and U5861 (N_5861,N_2987,N_346);
and U5862 (N_5862,N_1227,N_970);
nor U5863 (N_5863,N_1071,N_994);
and U5864 (N_5864,N_1997,N_1694);
or U5865 (N_5865,N_981,N_110);
nand U5866 (N_5866,N_1476,N_1264);
nand U5867 (N_5867,N_2158,N_872);
or U5868 (N_5868,N_1352,N_555);
or U5869 (N_5869,N_520,N_2819);
or U5870 (N_5870,N_876,N_2489);
or U5871 (N_5871,N_1357,N_3282);
and U5872 (N_5872,N_1455,N_821);
nand U5873 (N_5873,N_954,N_442);
and U5874 (N_5874,N_3750,N_1208);
or U5875 (N_5875,N_1272,N_3921);
or U5876 (N_5876,N_3879,N_2289);
nand U5877 (N_5877,N_3219,N_1393);
nor U5878 (N_5878,N_1350,N_2437);
nor U5879 (N_5879,N_1021,N_827);
xor U5880 (N_5880,N_2926,N_3444);
nor U5881 (N_5881,N_1260,N_2147);
nand U5882 (N_5882,N_1678,N_2798);
xnor U5883 (N_5883,N_1148,N_3041);
nand U5884 (N_5884,N_216,N_1776);
or U5885 (N_5885,N_2913,N_1183);
and U5886 (N_5886,N_3450,N_1514);
and U5887 (N_5887,N_899,N_1281);
xnor U5888 (N_5888,N_3257,N_704);
or U5889 (N_5889,N_2527,N_1461);
nand U5890 (N_5890,N_572,N_2331);
nor U5891 (N_5891,N_3177,N_3923);
and U5892 (N_5892,N_3410,N_930);
and U5893 (N_5893,N_42,N_2942);
nand U5894 (N_5894,N_2395,N_202);
nand U5895 (N_5895,N_3169,N_2827);
or U5896 (N_5896,N_2716,N_3110);
nor U5897 (N_5897,N_1869,N_2049);
and U5898 (N_5898,N_2155,N_1529);
or U5899 (N_5899,N_3195,N_3034);
or U5900 (N_5900,N_1588,N_2828);
or U5901 (N_5901,N_3593,N_934);
or U5902 (N_5902,N_711,N_2636);
and U5903 (N_5903,N_916,N_111);
nand U5904 (N_5904,N_3538,N_3174);
nor U5905 (N_5905,N_3609,N_236);
and U5906 (N_5906,N_838,N_2998);
nand U5907 (N_5907,N_1600,N_3875);
and U5908 (N_5908,N_3383,N_3554);
xnor U5909 (N_5909,N_2065,N_586);
or U5910 (N_5910,N_2239,N_225);
nor U5911 (N_5911,N_3871,N_1413);
and U5912 (N_5912,N_3080,N_3321);
nor U5913 (N_5913,N_3517,N_1056);
nor U5914 (N_5914,N_2522,N_870);
nand U5915 (N_5915,N_2106,N_2925);
and U5916 (N_5916,N_328,N_1767);
or U5917 (N_5917,N_3278,N_681);
nand U5918 (N_5918,N_1652,N_1037);
nand U5919 (N_5919,N_464,N_3953);
xnor U5920 (N_5920,N_273,N_1014);
and U5921 (N_5921,N_1583,N_2846);
nand U5922 (N_5922,N_2753,N_2978);
and U5923 (N_5923,N_698,N_3859);
nand U5924 (N_5924,N_3117,N_913);
or U5925 (N_5925,N_1371,N_2732);
nor U5926 (N_5926,N_1302,N_3451);
nor U5927 (N_5927,N_2100,N_3718);
xor U5928 (N_5928,N_3097,N_653);
nand U5929 (N_5929,N_1924,N_26);
nand U5930 (N_5930,N_2409,N_3186);
and U5931 (N_5931,N_1415,N_450);
nand U5932 (N_5932,N_2889,N_169);
nand U5933 (N_5933,N_619,N_2869);
and U5934 (N_5934,N_2051,N_2580);
or U5935 (N_5935,N_3056,N_1175);
nor U5936 (N_5936,N_1019,N_1722);
nor U5937 (N_5937,N_122,N_729);
and U5938 (N_5938,N_3398,N_2128);
nor U5939 (N_5939,N_1089,N_3838);
and U5940 (N_5940,N_3887,N_1676);
and U5941 (N_5941,N_1500,N_1456);
and U5942 (N_5942,N_2468,N_2087);
nand U5943 (N_5943,N_1236,N_1623);
xnor U5944 (N_5944,N_457,N_863);
or U5945 (N_5945,N_2728,N_3979);
or U5946 (N_5946,N_1486,N_2396);
nand U5947 (N_5947,N_1368,N_1392);
xnor U5948 (N_5948,N_3395,N_2858);
nor U5949 (N_5949,N_2142,N_2357);
and U5950 (N_5950,N_1919,N_2071);
nand U5951 (N_5951,N_1246,N_1890);
or U5952 (N_5952,N_3283,N_3623);
nand U5953 (N_5953,N_990,N_3804);
or U5954 (N_5954,N_3523,N_3503);
nand U5955 (N_5955,N_1409,N_3733);
and U5956 (N_5956,N_1900,N_2816);
nand U5957 (N_5957,N_2035,N_2408);
or U5958 (N_5958,N_874,N_2287);
nor U5959 (N_5959,N_2266,N_1372);
nor U5960 (N_5960,N_2989,N_2341);
or U5961 (N_5961,N_816,N_1205);
or U5962 (N_5962,N_1994,N_1804);
or U5963 (N_5963,N_991,N_128);
nand U5964 (N_5964,N_3630,N_2073);
nand U5965 (N_5965,N_2931,N_1699);
nand U5966 (N_5966,N_722,N_2559);
or U5967 (N_5967,N_3611,N_603);
and U5968 (N_5968,N_1650,N_2928);
xnor U5969 (N_5969,N_1656,N_2053);
xnor U5970 (N_5970,N_3020,N_543);
and U5971 (N_5971,N_3894,N_3480);
nor U5972 (N_5972,N_3276,N_334);
xor U5973 (N_5973,N_2955,N_115);
nor U5974 (N_5974,N_1338,N_2736);
xor U5975 (N_5975,N_2785,N_877);
and U5976 (N_5976,N_2058,N_2346);
nand U5977 (N_5977,N_2615,N_2016);
or U5978 (N_5978,N_3087,N_1961);
nand U5979 (N_5979,N_1096,N_1279);
or U5980 (N_5980,N_3259,N_2566);
nand U5981 (N_5981,N_1285,N_341);
or U5982 (N_5982,N_3462,N_277);
and U5983 (N_5983,N_2587,N_804);
and U5984 (N_5984,N_2923,N_3592);
or U5985 (N_5985,N_2259,N_265);
and U5986 (N_5986,N_537,N_3308);
and U5987 (N_5987,N_43,N_1553);
nand U5988 (N_5988,N_3060,N_3456);
nand U5989 (N_5989,N_3825,N_3754);
or U5990 (N_5990,N_3473,N_446);
and U5991 (N_5991,N_3170,N_2568);
nand U5992 (N_5992,N_3755,N_3300);
xor U5993 (N_5993,N_31,N_1928);
nor U5994 (N_5994,N_1558,N_647);
xnor U5995 (N_5995,N_3198,N_3285);
and U5996 (N_5996,N_441,N_2583);
xnor U5997 (N_5997,N_1111,N_2248);
nor U5998 (N_5998,N_3819,N_2996);
or U5999 (N_5999,N_156,N_1876);
nand U6000 (N_6000,N_335,N_675);
nor U6001 (N_6001,N_2098,N_3985);
nand U6002 (N_6002,N_2530,N_204);
nand U6003 (N_6003,N_3110,N_2697);
xnor U6004 (N_6004,N_3984,N_1072);
nand U6005 (N_6005,N_3300,N_1610);
xnor U6006 (N_6006,N_394,N_2075);
nand U6007 (N_6007,N_3997,N_203);
nand U6008 (N_6008,N_1402,N_2206);
xnor U6009 (N_6009,N_605,N_1279);
or U6010 (N_6010,N_3157,N_3568);
nor U6011 (N_6011,N_2955,N_633);
or U6012 (N_6012,N_3602,N_1748);
and U6013 (N_6013,N_3668,N_135);
or U6014 (N_6014,N_861,N_1721);
or U6015 (N_6015,N_2574,N_1489);
or U6016 (N_6016,N_2658,N_270);
nand U6017 (N_6017,N_100,N_2211);
or U6018 (N_6018,N_1676,N_1947);
xnor U6019 (N_6019,N_1336,N_1281);
nor U6020 (N_6020,N_1727,N_1313);
nand U6021 (N_6021,N_566,N_3209);
or U6022 (N_6022,N_1554,N_1123);
nand U6023 (N_6023,N_2340,N_143);
nand U6024 (N_6024,N_1548,N_827);
nor U6025 (N_6025,N_2981,N_1718);
nor U6026 (N_6026,N_1331,N_1246);
or U6027 (N_6027,N_514,N_1558);
or U6028 (N_6028,N_3099,N_2502);
nand U6029 (N_6029,N_3613,N_1400);
and U6030 (N_6030,N_3814,N_135);
nand U6031 (N_6031,N_2800,N_988);
and U6032 (N_6032,N_2329,N_1642);
nor U6033 (N_6033,N_2609,N_2344);
or U6034 (N_6034,N_1862,N_1017);
or U6035 (N_6035,N_609,N_1635);
and U6036 (N_6036,N_660,N_427);
nor U6037 (N_6037,N_2735,N_1095);
nand U6038 (N_6038,N_3426,N_1039);
nand U6039 (N_6039,N_3495,N_3481);
nor U6040 (N_6040,N_3942,N_2239);
and U6041 (N_6041,N_263,N_2988);
or U6042 (N_6042,N_1231,N_1035);
nor U6043 (N_6043,N_2721,N_3632);
and U6044 (N_6044,N_1671,N_3323);
xor U6045 (N_6045,N_3467,N_1895);
nand U6046 (N_6046,N_1501,N_2108);
nand U6047 (N_6047,N_3512,N_3568);
nor U6048 (N_6048,N_1392,N_2328);
or U6049 (N_6049,N_2835,N_70);
nor U6050 (N_6050,N_2197,N_1121);
xor U6051 (N_6051,N_2428,N_1777);
and U6052 (N_6052,N_2373,N_3738);
or U6053 (N_6053,N_193,N_1691);
or U6054 (N_6054,N_2714,N_1615);
nand U6055 (N_6055,N_2932,N_3296);
or U6056 (N_6056,N_3872,N_3889);
or U6057 (N_6057,N_3498,N_2937);
nor U6058 (N_6058,N_2509,N_2797);
and U6059 (N_6059,N_1002,N_3366);
nand U6060 (N_6060,N_420,N_404);
nor U6061 (N_6061,N_124,N_2120);
or U6062 (N_6062,N_1591,N_1610);
nand U6063 (N_6063,N_1473,N_3309);
nor U6064 (N_6064,N_3518,N_2935);
and U6065 (N_6065,N_3557,N_3750);
or U6066 (N_6066,N_342,N_429);
nand U6067 (N_6067,N_3629,N_105);
and U6068 (N_6068,N_1986,N_268);
nand U6069 (N_6069,N_1100,N_3295);
or U6070 (N_6070,N_630,N_2512);
xnor U6071 (N_6071,N_606,N_2083);
xnor U6072 (N_6072,N_373,N_2963);
and U6073 (N_6073,N_3635,N_3747);
and U6074 (N_6074,N_70,N_1723);
or U6075 (N_6075,N_2660,N_3946);
xor U6076 (N_6076,N_308,N_2262);
or U6077 (N_6077,N_843,N_3211);
and U6078 (N_6078,N_3870,N_74);
and U6079 (N_6079,N_1619,N_2820);
nand U6080 (N_6080,N_2740,N_1790);
nand U6081 (N_6081,N_383,N_1080);
or U6082 (N_6082,N_1108,N_3701);
or U6083 (N_6083,N_2692,N_667);
or U6084 (N_6084,N_1351,N_3595);
nand U6085 (N_6085,N_1081,N_672);
xnor U6086 (N_6086,N_3031,N_1748);
or U6087 (N_6087,N_2493,N_62);
nand U6088 (N_6088,N_2055,N_2487);
nand U6089 (N_6089,N_2666,N_3732);
or U6090 (N_6090,N_2971,N_1055);
or U6091 (N_6091,N_3322,N_1248);
and U6092 (N_6092,N_790,N_2106);
nand U6093 (N_6093,N_3953,N_3325);
xnor U6094 (N_6094,N_3373,N_1622);
or U6095 (N_6095,N_930,N_953);
and U6096 (N_6096,N_3330,N_2945);
or U6097 (N_6097,N_1766,N_2675);
and U6098 (N_6098,N_2687,N_1453);
nor U6099 (N_6099,N_1759,N_223);
nor U6100 (N_6100,N_2012,N_2523);
or U6101 (N_6101,N_1991,N_762);
and U6102 (N_6102,N_1125,N_2304);
and U6103 (N_6103,N_2437,N_2171);
nand U6104 (N_6104,N_757,N_1702);
nand U6105 (N_6105,N_1090,N_2325);
nand U6106 (N_6106,N_60,N_965);
nor U6107 (N_6107,N_3504,N_1490);
nor U6108 (N_6108,N_3366,N_2624);
or U6109 (N_6109,N_2683,N_386);
and U6110 (N_6110,N_3118,N_488);
nor U6111 (N_6111,N_943,N_1098);
and U6112 (N_6112,N_2403,N_627);
nand U6113 (N_6113,N_1089,N_3956);
nor U6114 (N_6114,N_687,N_2730);
and U6115 (N_6115,N_477,N_3806);
or U6116 (N_6116,N_2470,N_2185);
and U6117 (N_6117,N_506,N_428);
xor U6118 (N_6118,N_2417,N_998);
and U6119 (N_6119,N_963,N_1361);
nor U6120 (N_6120,N_1368,N_1419);
and U6121 (N_6121,N_837,N_728);
nand U6122 (N_6122,N_3963,N_483);
nor U6123 (N_6123,N_2272,N_2402);
nor U6124 (N_6124,N_425,N_677);
nand U6125 (N_6125,N_1850,N_1569);
nor U6126 (N_6126,N_3781,N_2865);
or U6127 (N_6127,N_2803,N_3008);
nand U6128 (N_6128,N_2114,N_3744);
nor U6129 (N_6129,N_2009,N_692);
nand U6130 (N_6130,N_1175,N_1628);
nand U6131 (N_6131,N_141,N_1710);
nand U6132 (N_6132,N_124,N_1952);
or U6133 (N_6133,N_15,N_2929);
nand U6134 (N_6134,N_991,N_62);
and U6135 (N_6135,N_259,N_3172);
and U6136 (N_6136,N_192,N_1140);
and U6137 (N_6137,N_2282,N_1210);
nand U6138 (N_6138,N_2311,N_3006);
or U6139 (N_6139,N_3318,N_3756);
nor U6140 (N_6140,N_2259,N_3335);
or U6141 (N_6141,N_1877,N_3855);
and U6142 (N_6142,N_3699,N_1545);
nand U6143 (N_6143,N_983,N_3340);
nand U6144 (N_6144,N_2569,N_3906);
nand U6145 (N_6145,N_1029,N_1861);
and U6146 (N_6146,N_162,N_3042);
nand U6147 (N_6147,N_3296,N_973);
nand U6148 (N_6148,N_478,N_3902);
and U6149 (N_6149,N_808,N_1964);
and U6150 (N_6150,N_955,N_1465);
nor U6151 (N_6151,N_2088,N_2481);
nand U6152 (N_6152,N_2892,N_936);
or U6153 (N_6153,N_2745,N_1391);
or U6154 (N_6154,N_3063,N_3859);
nand U6155 (N_6155,N_1538,N_1595);
nor U6156 (N_6156,N_2824,N_2800);
or U6157 (N_6157,N_2605,N_3161);
and U6158 (N_6158,N_3519,N_899);
or U6159 (N_6159,N_1203,N_70);
nor U6160 (N_6160,N_1596,N_3731);
and U6161 (N_6161,N_2835,N_305);
or U6162 (N_6162,N_457,N_2802);
or U6163 (N_6163,N_1984,N_3976);
or U6164 (N_6164,N_2240,N_3982);
nor U6165 (N_6165,N_1580,N_3039);
xor U6166 (N_6166,N_3983,N_3017);
nor U6167 (N_6167,N_1718,N_2729);
nand U6168 (N_6168,N_1547,N_719);
nand U6169 (N_6169,N_1847,N_2851);
nor U6170 (N_6170,N_3450,N_2245);
nand U6171 (N_6171,N_76,N_1864);
or U6172 (N_6172,N_3970,N_1468);
nor U6173 (N_6173,N_3229,N_1856);
and U6174 (N_6174,N_1578,N_395);
or U6175 (N_6175,N_1930,N_2875);
nor U6176 (N_6176,N_3380,N_3332);
and U6177 (N_6177,N_1133,N_1819);
nand U6178 (N_6178,N_351,N_3254);
or U6179 (N_6179,N_832,N_1233);
and U6180 (N_6180,N_2865,N_2757);
nand U6181 (N_6181,N_1533,N_15);
or U6182 (N_6182,N_2544,N_2526);
xnor U6183 (N_6183,N_1757,N_1927);
and U6184 (N_6184,N_3153,N_1649);
or U6185 (N_6185,N_188,N_23);
nor U6186 (N_6186,N_1891,N_2811);
nand U6187 (N_6187,N_1986,N_1769);
nand U6188 (N_6188,N_1791,N_2818);
nor U6189 (N_6189,N_3160,N_2179);
nor U6190 (N_6190,N_348,N_331);
and U6191 (N_6191,N_2334,N_2173);
or U6192 (N_6192,N_2895,N_1608);
or U6193 (N_6193,N_2356,N_616);
or U6194 (N_6194,N_1654,N_3726);
or U6195 (N_6195,N_3660,N_2634);
or U6196 (N_6196,N_591,N_2263);
nor U6197 (N_6197,N_3209,N_998);
nand U6198 (N_6198,N_2310,N_2701);
and U6199 (N_6199,N_2928,N_1530);
nor U6200 (N_6200,N_2455,N_995);
or U6201 (N_6201,N_1665,N_3500);
nor U6202 (N_6202,N_339,N_2052);
and U6203 (N_6203,N_3492,N_2662);
and U6204 (N_6204,N_3637,N_2202);
and U6205 (N_6205,N_1354,N_1883);
and U6206 (N_6206,N_2743,N_711);
or U6207 (N_6207,N_1057,N_1499);
or U6208 (N_6208,N_3111,N_923);
nor U6209 (N_6209,N_3773,N_3917);
nand U6210 (N_6210,N_3294,N_2512);
or U6211 (N_6211,N_1513,N_511);
and U6212 (N_6212,N_1296,N_2810);
nor U6213 (N_6213,N_1656,N_1878);
xor U6214 (N_6214,N_2740,N_1807);
or U6215 (N_6215,N_3419,N_3410);
or U6216 (N_6216,N_1423,N_238);
xor U6217 (N_6217,N_443,N_2673);
and U6218 (N_6218,N_3816,N_320);
nor U6219 (N_6219,N_2651,N_2711);
and U6220 (N_6220,N_958,N_178);
or U6221 (N_6221,N_2660,N_2470);
nand U6222 (N_6222,N_2836,N_1890);
nand U6223 (N_6223,N_2549,N_3482);
xor U6224 (N_6224,N_2481,N_3837);
nor U6225 (N_6225,N_428,N_2336);
or U6226 (N_6226,N_2205,N_2930);
nand U6227 (N_6227,N_3898,N_1059);
and U6228 (N_6228,N_3566,N_3370);
or U6229 (N_6229,N_1244,N_2383);
or U6230 (N_6230,N_3713,N_2611);
nand U6231 (N_6231,N_3923,N_2136);
nand U6232 (N_6232,N_3249,N_3507);
nand U6233 (N_6233,N_2214,N_357);
and U6234 (N_6234,N_2689,N_2784);
or U6235 (N_6235,N_3919,N_1466);
xnor U6236 (N_6236,N_3939,N_2261);
or U6237 (N_6237,N_1912,N_1658);
or U6238 (N_6238,N_847,N_1024);
and U6239 (N_6239,N_1318,N_1468);
nor U6240 (N_6240,N_1303,N_3445);
nand U6241 (N_6241,N_1628,N_1996);
and U6242 (N_6242,N_909,N_1029);
and U6243 (N_6243,N_1697,N_3040);
nand U6244 (N_6244,N_2524,N_3828);
nor U6245 (N_6245,N_756,N_2503);
nor U6246 (N_6246,N_3140,N_3366);
nor U6247 (N_6247,N_3525,N_3116);
or U6248 (N_6248,N_3492,N_764);
or U6249 (N_6249,N_2958,N_3523);
nor U6250 (N_6250,N_866,N_3757);
nor U6251 (N_6251,N_3734,N_984);
xnor U6252 (N_6252,N_3293,N_1031);
nor U6253 (N_6253,N_1763,N_85);
or U6254 (N_6254,N_1598,N_1374);
nand U6255 (N_6255,N_401,N_3474);
nand U6256 (N_6256,N_2667,N_259);
nand U6257 (N_6257,N_3874,N_80);
nor U6258 (N_6258,N_2861,N_2404);
or U6259 (N_6259,N_849,N_1374);
or U6260 (N_6260,N_2793,N_569);
xnor U6261 (N_6261,N_881,N_22);
or U6262 (N_6262,N_3493,N_2457);
or U6263 (N_6263,N_156,N_3587);
nand U6264 (N_6264,N_1547,N_2163);
nand U6265 (N_6265,N_2555,N_1751);
or U6266 (N_6266,N_354,N_6);
and U6267 (N_6267,N_2167,N_2826);
nor U6268 (N_6268,N_1694,N_271);
or U6269 (N_6269,N_2844,N_3680);
xnor U6270 (N_6270,N_548,N_1353);
or U6271 (N_6271,N_1619,N_1612);
or U6272 (N_6272,N_3717,N_1271);
nor U6273 (N_6273,N_1523,N_2355);
or U6274 (N_6274,N_244,N_3326);
and U6275 (N_6275,N_79,N_2758);
nor U6276 (N_6276,N_1763,N_2104);
nand U6277 (N_6277,N_2832,N_1257);
xnor U6278 (N_6278,N_3276,N_2750);
or U6279 (N_6279,N_60,N_3980);
or U6280 (N_6280,N_803,N_3662);
nand U6281 (N_6281,N_744,N_12);
or U6282 (N_6282,N_3958,N_2376);
nor U6283 (N_6283,N_1225,N_1714);
or U6284 (N_6284,N_1668,N_2956);
and U6285 (N_6285,N_3279,N_2699);
and U6286 (N_6286,N_1756,N_416);
nand U6287 (N_6287,N_2683,N_189);
nand U6288 (N_6288,N_1519,N_2279);
nor U6289 (N_6289,N_3205,N_3865);
nand U6290 (N_6290,N_1225,N_3362);
xor U6291 (N_6291,N_33,N_3895);
xnor U6292 (N_6292,N_2134,N_1254);
and U6293 (N_6293,N_3114,N_2537);
nor U6294 (N_6294,N_3786,N_861);
and U6295 (N_6295,N_158,N_3292);
nand U6296 (N_6296,N_488,N_682);
nand U6297 (N_6297,N_3086,N_1569);
or U6298 (N_6298,N_2795,N_2646);
or U6299 (N_6299,N_3380,N_838);
and U6300 (N_6300,N_516,N_1283);
nand U6301 (N_6301,N_493,N_3030);
nand U6302 (N_6302,N_2507,N_2222);
and U6303 (N_6303,N_3098,N_3135);
and U6304 (N_6304,N_801,N_2956);
and U6305 (N_6305,N_1822,N_20);
nor U6306 (N_6306,N_1404,N_3373);
nand U6307 (N_6307,N_2577,N_2101);
nand U6308 (N_6308,N_790,N_3340);
nand U6309 (N_6309,N_3574,N_3013);
nor U6310 (N_6310,N_631,N_3420);
nand U6311 (N_6311,N_1120,N_1375);
nand U6312 (N_6312,N_2965,N_3191);
and U6313 (N_6313,N_394,N_2913);
and U6314 (N_6314,N_1121,N_1128);
xnor U6315 (N_6315,N_1734,N_856);
or U6316 (N_6316,N_3856,N_147);
and U6317 (N_6317,N_383,N_2003);
nor U6318 (N_6318,N_1670,N_921);
nand U6319 (N_6319,N_149,N_1180);
nand U6320 (N_6320,N_2272,N_1432);
and U6321 (N_6321,N_2041,N_669);
and U6322 (N_6322,N_3037,N_2742);
nor U6323 (N_6323,N_2284,N_115);
and U6324 (N_6324,N_3796,N_1960);
nand U6325 (N_6325,N_1987,N_2665);
xor U6326 (N_6326,N_2801,N_3409);
nand U6327 (N_6327,N_3743,N_3491);
and U6328 (N_6328,N_3833,N_3669);
or U6329 (N_6329,N_2512,N_342);
and U6330 (N_6330,N_1500,N_3641);
nand U6331 (N_6331,N_293,N_2325);
xnor U6332 (N_6332,N_2962,N_2694);
nor U6333 (N_6333,N_713,N_2276);
and U6334 (N_6334,N_1007,N_3796);
and U6335 (N_6335,N_1066,N_991);
or U6336 (N_6336,N_1320,N_3257);
xnor U6337 (N_6337,N_3905,N_3727);
and U6338 (N_6338,N_2490,N_2897);
nand U6339 (N_6339,N_2149,N_1757);
nand U6340 (N_6340,N_2587,N_3074);
nand U6341 (N_6341,N_1966,N_965);
or U6342 (N_6342,N_110,N_3807);
nor U6343 (N_6343,N_1667,N_3956);
nor U6344 (N_6344,N_1193,N_2118);
and U6345 (N_6345,N_2915,N_3642);
nor U6346 (N_6346,N_1329,N_3203);
nor U6347 (N_6347,N_83,N_642);
and U6348 (N_6348,N_1730,N_287);
xor U6349 (N_6349,N_3397,N_3679);
nand U6350 (N_6350,N_990,N_2404);
nand U6351 (N_6351,N_3489,N_130);
and U6352 (N_6352,N_3890,N_1517);
nand U6353 (N_6353,N_2927,N_2802);
nand U6354 (N_6354,N_1396,N_2266);
or U6355 (N_6355,N_1204,N_2831);
nor U6356 (N_6356,N_56,N_3080);
xnor U6357 (N_6357,N_2799,N_637);
or U6358 (N_6358,N_338,N_2285);
nor U6359 (N_6359,N_2696,N_3707);
and U6360 (N_6360,N_2886,N_1374);
and U6361 (N_6361,N_1113,N_2616);
xor U6362 (N_6362,N_194,N_887);
nand U6363 (N_6363,N_618,N_2147);
and U6364 (N_6364,N_2522,N_357);
nand U6365 (N_6365,N_1516,N_2393);
nand U6366 (N_6366,N_598,N_1945);
nor U6367 (N_6367,N_2981,N_29);
xnor U6368 (N_6368,N_3066,N_1091);
nand U6369 (N_6369,N_1416,N_3648);
nor U6370 (N_6370,N_2553,N_1054);
nor U6371 (N_6371,N_3812,N_2563);
nand U6372 (N_6372,N_1508,N_668);
or U6373 (N_6373,N_1263,N_1935);
nand U6374 (N_6374,N_2584,N_2217);
nor U6375 (N_6375,N_3250,N_164);
or U6376 (N_6376,N_2039,N_3880);
or U6377 (N_6377,N_730,N_305);
xnor U6378 (N_6378,N_447,N_305);
nand U6379 (N_6379,N_468,N_1554);
or U6380 (N_6380,N_3573,N_1940);
or U6381 (N_6381,N_361,N_97);
or U6382 (N_6382,N_572,N_2096);
and U6383 (N_6383,N_2038,N_1264);
and U6384 (N_6384,N_1068,N_753);
nand U6385 (N_6385,N_1123,N_3527);
and U6386 (N_6386,N_1086,N_2801);
nand U6387 (N_6387,N_1331,N_3637);
and U6388 (N_6388,N_3746,N_1169);
nor U6389 (N_6389,N_3197,N_3185);
or U6390 (N_6390,N_2233,N_2512);
nand U6391 (N_6391,N_3466,N_383);
or U6392 (N_6392,N_498,N_3135);
xnor U6393 (N_6393,N_3762,N_1161);
and U6394 (N_6394,N_547,N_1336);
xor U6395 (N_6395,N_289,N_3592);
nor U6396 (N_6396,N_1843,N_1533);
or U6397 (N_6397,N_1601,N_1029);
nor U6398 (N_6398,N_2843,N_1605);
and U6399 (N_6399,N_373,N_1246);
nand U6400 (N_6400,N_345,N_1386);
or U6401 (N_6401,N_2420,N_891);
or U6402 (N_6402,N_3405,N_1802);
nand U6403 (N_6403,N_2654,N_2426);
nand U6404 (N_6404,N_2772,N_1703);
xor U6405 (N_6405,N_3272,N_373);
nand U6406 (N_6406,N_866,N_3617);
and U6407 (N_6407,N_3567,N_461);
and U6408 (N_6408,N_2746,N_3077);
and U6409 (N_6409,N_1305,N_510);
nor U6410 (N_6410,N_2850,N_2364);
or U6411 (N_6411,N_1001,N_2121);
and U6412 (N_6412,N_1844,N_104);
nand U6413 (N_6413,N_3159,N_2431);
or U6414 (N_6414,N_1673,N_3307);
nand U6415 (N_6415,N_2463,N_2046);
and U6416 (N_6416,N_1525,N_3287);
nand U6417 (N_6417,N_1680,N_3022);
or U6418 (N_6418,N_3040,N_708);
and U6419 (N_6419,N_502,N_2589);
nand U6420 (N_6420,N_3007,N_1019);
nand U6421 (N_6421,N_169,N_1874);
or U6422 (N_6422,N_1257,N_1);
or U6423 (N_6423,N_1020,N_2778);
nor U6424 (N_6424,N_3501,N_2927);
and U6425 (N_6425,N_3145,N_2181);
and U6426 (N_6426,N_1143,N_74);
and U6427 (N_6427,N_931,N_1673);
nand U6428 (N_6428,N_3570,N_3002);
nand U6429 (N_6429,N_151,N_2889);
and U6430 (N_6430,N_1678,N_1831);
or U6431 (N_6431,N_748,N_3738);
nand U6432 (N_6432,N_2781,N_2133);
or U6433 (N_6433,N_3115,N_2905);
or U6434 (N_6434,N_2031,N_3997);
or U6435 (N_6435,N_2443,N_549);
or U6436 (N_6436,N_612,N_808);
or U6437 (N_6437,N_449,N_3155);
and U6438 (N_6438,N_2597,N_938);
and U6439 (N_6439,N_632,N_1696);
or U6440 (N_6440,N_1088,N_3972);
or U6441 (N_6441,N_3794,N_1472);
nand U6442 (N_6442,N_1910,N_2050);
nand U6443 (N_6443,N_243,N_380);
or U6444 (N_6444,N_2066,N_1597);
nand U6445 (N_6445,N_2073,N_2827);
nand U6446 (N_6446,N_37,N_1547);
nand U6447 (N_6447,N_2420,N_11);
or U6448 (N_6448,N_3918,N_1818);
and U6449 (N_6449,N_1577,N_1894);
and U6450 (N_6450,N_3367,N_1669);
xnor U6451 (N_6451,N_1533,N_134);
xor U6452 (N_6452,N_3949,N_3514);
nor U6453 (N_6453,N_1917,N_3925);
nand U6454 (N_6454,N_881,N_2972);
nor U6455 (N_6455,N_3134,N_1090);
nor U6456 (N_6456,N_2702,N_1535);
and U6457 (N_6457,N_3015,N_79);
nor U6458 (N_6458,N_319,N_1437);
and U6459 (N_6459,N_1076,N_1154);
xnor U6460 (N_6460,N_1293,N_3512);
or U6461 (N_6461,N_3135,N_2883);
xnor U6462 (N_6462,N_3491,N_3587);
or U6463 (N_6463,N_3988,N_1017);
nand U6464 (N_6464,N_574,N_690);
nor U6465 (N_6465,N_3019,N_3328);
and U6466 (N_6466,N_990,N_3234);
or U6467 (N_6467,N_3255,N_2843);
or U6468 (N_6468,N_1722,N_2152);
nor U6469 (N_6469,N_2503,N_186);
xnor U6470 (N_6470,N_1124,N_2698);
nand U6471 (N_6471,N_3946,N_503);
and U6472 (N_6472,N_403,N_476);
xor U6473 (N_6473,N_565,N_525);
or U6474 (N_6474,N_3670,N_1810);
nor U6475 (N_6475,N_3937,N_3980);
or U6476 (N_6476,N_805,N_2453);
and U6477 (N_6477,N_703,N_153);
nor U6478 (N_6478,N_2473,N_2895);
nor U6479 (N_6479,N_185,N_2827);
or U6480 (N_6480,N_3343,N_3934);
or U6481 (N_6481,N_3681,N_3298);
or U6482 (N_6482,N_2020,N_881);
nor U6483 (N_6483,N_2588,N_408);
or U6484 (N_6484,N_647,N_1155);
nand U6485 (N_6485,N_431,N_870);
and U6486 (N_6486,N_2971,N_2838);
nor U6487 (N_6487,N_2015,N_3100);
nor U6488 (N_6488,N_1114,N_3085);
and U6489 (N_6489,N_1726,N_3115);
and U6490 (N_6490,N_1291,N_1303);
xor U6491 (N_6491,N_1932,N_2649);
nand U6492 (N_6492,N_2546,N_677);
nor U6493 (N_6493,N_2297,N_3342);
or U6494 (N_6494,N_3265,N_2067);
or U6495 (N_6495,N_237,N_2920);
or U6496 (N_6496,N_2115,N_1526);
and U6497 (N_6497,N_1626,N_1894);
xnor U6498 (N_6498,N_2882,N_465);
and U6499 (N_6499,N_1508,N_720);
xor U6500 (N_6500,N_715,N_3778);
and U6501 (N_6501,N_1191,N_3947);
or U6502 (N_6502,N_3149,N_471);
and U6503 (N_6503,N_2103,N_770);
or U6504 (N_6504,N_1250,N_1350);
or U6505 (N_6505,N_906,N_3281);
and U6506 (N_6506,N_527,N_2513);
or U6507 (N_6507,N_1738,N_1818);
and U6508 (N_6508,N_2037,N_3097);
nand U6509 (N_6509,N_1104,N_1684);
or U6510 (N_6510,N_26,N_3915);
and U6511 (N_6511,N_317,N_2707);
and U6512 (N_6512,N_3748,N_2859);
or U6513 (N_6513,N_1842,N_2335);
or U6514 (N_6514,N_2605,N_2222);
nor U6515 (N_6515,N_971,N_2533);
nor U6516 (N_6516,N_2435,N_3437);
or U6517 (N_6517,N_2326,N_2114);
or U6518 (N_6518,N_3104,N_1932);
nand U6519 (N_6519,N_376,N_1573);
or U6520 (N_6520,N_3007,N_1401);
or U6521 (N_6521,N_2547,N_379);
and U6522 (N_6522,N_2555,N_1511);
nand U6523 (N_6523,N_1998,N_356);
nand U6524 (N_6524,N_2882,N_626);
xor U6525 (N_6525,N_1372,N_3517);
nand U6526 (N_6526,N_1309,N_999);
and U6527 (N_6527,N_2447,N_1557);
xor U6528 (N_6528,N_3797,N_2693);
and U6529 (N_6529,N_2370,N_2728);
and U6530 (N_6530,N_1422,N_2705);
or U6531 (N_6531,N_3227,N_3163);
xor U6532 (N_6532,N_2369,N_1125);
nand U6533 (N_6533,N_2364,N_3208);
and U6534 (N_6534,N_272,N_1403);
or U6535 (N_6535,N_2223,N_374);
nor U6536 (N_6536,N_183,N_2724);
nand U6537 (N_6537,N_1036,N_763);
or U6538 (N_6538,N_1442,N_3877);
nand U6539 (N_6539,N_2863,N_1058);
and U6540 (N_6540,N_3359,N_3975);
nand U6541 (N_6541,N_1923,N_2469);
nor U6542 (N_6542,N_154,N_3774);
nor U6543 (N_6543,N_1095,N_1200);
and U6544 (N_6544,N_1202,N_2585);
or U6545 (N_6545,N_3696,N_2709);
nor U6546 (N_6546,N_3247,N_1887);
or U6547 (N_6547,N_714,N_3902);
nand U6548 (N_6548,N_1068,N_2325);
and U6549 (N_6549,N_321,N_3196);
nor U6550 (N_6550,N_359,N_2600);
or U6551 (N_6551,N_731,N_1532);
xnor U6552 (N_6552,N_359,N_3146);
nor U6553 (N_6553,N_2391,N_2054);
and U6554 (N_6554,N_2147,N_3472);
and U6555 (N_6555,N_2255,N_134);
and U6556 (N_6556,N_913,N_2643);
nand U6557 (N_6557,N_1924,N_1693);
or U6558 (N_6558,N_892,N_1185);
or U6559 (N_6559,N_54,N_257);
nand U6560 (N_6560,N_3165,N_1438);
nand U6561 (N_6561,N_1270,N_2518);
or U6562 (N_6562,N_1726,N_2864);
and U6563 (N_6563,N_767,N_2982);
or U6564 (N_6564,N_1411,N_1912);
or U6565 (N_6565,N_3761,N_39);
and U6566 (N_6566,N_3935,N_3199);
nand U6567 (N_6567,N_400,N_2540);
or U6568 (N_6568,N_469,N_2179);
and U6569 (N_6569,N_3613,N_3721);
nand U6570 (N_6570,N_3734,N_2382);
nor U6571 (N_6571,N_3389,N_351);
nor U6572 (N_6572,N_1542,N_3228);
or U6573 (N_6573,N_2594,N_3964);
nand U6574 (N_6574,N_617,N_3477);
xor U6575 (N_6575,N_3854,N_180);
nor U6576 (N_6576,N_1486,N_3338);
and U6577 (N_6577,N_3332,N_78);
xnor U6578 (N_6578,N_3997,N_3466);
and U6579 (N_6579,N_3831,N_3075);
or U6580 (N_6580,N_2694,N_2100);
nand U6581 (N_6581,N_3672,N_1085);
nand U6582 (N_6582,N_1569,N_3088);
nor U6583 (N_6583,N_3518,N_1395);
or U6584 (N_6584,N_2931,N_266);
nor U6585 (N_6585,N_2487,N_3501);
nor U6586 (N_6586,N_2422,N_3364);
xor U6587 (N_6587,N_2565,N_1180);
or U6588 (N_6588,N_2847,N_2135);
nand U6589 (N_6589,N_1395,N_684);
nor U6590 (N_6590,N_1601,N_1365);
nand U6591 (N_6591,N_3399,N_2210);
or U6592 (N_6592,N_1266,N_2760);
or U6593 (N_6593,N_207,N_955);
or U6594 (N_6594,N_1382,N_458);
nand U6595 (N_6595,N_2232,N_553);
nand U6596 (N_6596,N_1140,N_2336);
or U6597 (N_6597,N_181,N_2869);
and U6598 (N_6598,N_82,N_1057);
xor U6599 (N_6599,N_53,N_1259);
and U6600 (N_6600,N_3190,N_674);
nand U6601 (N_6601,N_2040,N_3422);
nand U6602 (N_6602,N_1463,N_842);
or U6603 (N_6603,N_3150,N_2561);
xnor U6604 (N_6604,N_822,N_3321);
and U6605 (N_6605,N_975,N_1880);
nand U6606 (N_6606,N_3615,N_717);
and U6607 (N_6607,N_1793,N_841);
nor U6608 (N_6608,N_2894,N_360);
or U6609 (N_6609,N_605,N_3566);
nor U6610 (N_6610,N_810,N_1439);
and U6611 (N_6611,N_838,N_3726);
or U6612 (N_6612,N_1960,N_1937);
or U6613 (N_6613,N_1123,N_1179);
nand U6614 (N_6614,N_3205,N_974);
nand U6615 (N_6615,N_3104,N_1709);
or U6616 (N_6616,N_3596,N_44);
nand U6617 (N_6617,N_133,N_155);
xnor U6618 (N_6618,N_2787,N_1519);
nor U6619 (N_6619,N_1764,N_2432);
nand U6620 (N_6620,N_748,N_1492);
and U6621 (N_6621,N_1528,N_2498);
or U6622 (N_6622,N_2208,N_2335);
and U6623 (N_6623,N_362,N_1045);
nand U6624 (N_6624,N_3998,N_3679);
and U6625 (N_6625,N_252,N_2164);
nand U6626 (N_6626,N_3712,N_2717);
or U6627 (N_6627,N_3975,N_3213);
nor U6628 (N_6628,N_1183,N_2452);
and U6629 (N_6629,N_2290,N_2);
and U6630 (N_6630,N_835,N_1163);
nor U6631 (N_6631,N_3366,N_3002);
nand U6632 (N_6632,N_1260,N_1821);
or U6633 (N_6633,N_1648,N_3505);
or U6634 (N_6634,N_3482,N_3037);
nand U6635 (N_6635,N_3625,N_476);
nand U6636 (N_6636,N_3111,N_2754);
or U6637 (N_6637,N_2298,N_1318);
or U6638 (N_6638,N_402,N_405);
nor U6639 (N_6639,N_3753,N_2125);
or U6640 (N_6640,N_2930,N_274);
nand U6641 (N_6641,N_822,N_2219);
xnor U6642 (N_6642,N_1165,N_3453);
nand U6643 (N_6643,N_3596,N_2819);
nand U6644 (N_6644,N_1255,N_226);
nand U6645 (N_6645,N_376,N_993);
or U6646 (N_6646,N_836,N_1136);
nand U6647 (N_6647,N_1829,N_2244);
nor U6648 (N_6648,N_2468,N_2634);
xor U6649 (N_6649,N_1886,N_1328);
xnor U6650 (N_6650,N_162,N_1723);
nor U6651 (N_6651,N_1563,N_2427);
xnor U6652 (N_6652,N_1109,N_3176);
and U6653 (N_6653,N_635,N_2954);
nor U6654 (N_6654,N_3154,N_414);
xor U6655 (N_6655,N_3943,N_2170);
and U6656 (N_6656,N_2736,N_3006);
nand U6657 (N_6657,N_811,N_1301);
or U6658 (N_6658,N_3635,N_908);
nor U6659 (N_6659,N_2956,N_2298);
xor U6660 (N_6660,N_3764,N_3809);
nor U6661 (N_6661,N_305,N_3136);
xnor U6662 (N_6662,N_2434,N_2501);
nor U6663 (N_6663,N_2222,N_2051);
and U6664 (N_6664,N_470,N_1641);
nor U6665 (N_6665,N_3409,N_980);
or U6666 (N_6666,N_1451,N_1868);
or U6667 (N_6667,N_1588,N_3615);
and U6668 (N_6668,N_3958,N_3471);
nor U6669 (N_6669,N_1407,N_2243);
and U6670 (N_6670,N_3765,N_16);
nor U6671 (N_6671,N_372,N_2662);
nor U6672 (N_6672,N_2168,N_580);
nor U6673 (N_6673,N_3284,N_1078);
nand U6674 (N_6674,N_1680,N_1805);
and U6675 (N_6675,N_606,N_3731);
and U6676 (N_6676,N_2704,N_207);
and U6677 (N_6677,N_3794,N_1389);
xnor U6678 (N_6678,N_3718,N_2406);
and U6679 (N_6679,N_61,N_165);
or U6680 (N_6680,N_545,N_2954);
and U6681 (N_6681,N_3281,N_2704);
nand U6682 (N_6682,N_606,N_3662);
and U6683 (N_6683,N_2522,N_3558);
nand U6684 (N_6684,N_1154,N_1961);
nand U6685 (N_6685,N_2035,N_3305);
or U6686 (N_6686,N_79,N_3724);
nor U6687 (N_6687,N_2571,N_1909);
nand U6688 (N_6688,N_1857,N_1099);
and U6689 (N_6689,N_3573,N_2142);
or U6690 (N_6690,N_3752,N_1771);
nor U6691 (N_6691,N_2391,N_2393);
nand U6692 (N_6692,N_3368,N_2125);
or U6693 (N_6693,N_2622,N_3575);
and U6694 (N_6694,N_1045,N_926);
xnor U6695 (N_6695,N_3379,N_1089);
nand U6696 (N_6696,N_2109,N_262);
and U6697 (N_6697,N_3257,N_3750);
nor U6698 (N_6698,N_3299,N_1397);
nand U6699 (N_6699,N_2737,N_474);
and U6700 (N_6700,N_647,N_1256);
nor U6701 (N_6701,N_148,N_982);
nand U6702 (N_6702,N_1557,N_238);
or U6703 (N_6703,N_895,N_2815);
or U6704 (N_6704,N_559,N_860);
nor U6705 (N_6705,N_3973,N_2284);
nor U6706 (N_6706,N_2083,N_1928);
and U6707 (N_6707,N_3445,N_374);
nor U6708 (N_6708,N_1058,N_3727);
nand U6709 (N_6709,N_3155,N_2455);
nor U6710 (N_6710,N_1193,N_659);
or U6711 (N_6711,N_3004,N_1332);
and U6712 (N_6712,N_1757,N_1180);
and U6713 (N_6713,N_2672,N_3378);
or U6714 (N_6714,N_3323,N_3280);
nor U6715 (N_6715,N_97,N_2784);
nand U6716 (N_6716,N_1472,N_1354);
or U6717 (N_6717,N_3649,N_3682);
or U6718 (N_6718,N_627,N_2314);
nor U6719 (N_6719,N_3062,N_3621);
nor U6720 (N_6720,N_2435,N_2357);
xor U6721 (N_6721,N_1230,N_1511);
nand U6722 (N_6722,N_464,N_690);
or U6723 (N_6723,N_726,N_2969);
and U6724 (N_6724,N_3159,N_686);
or U6725 (N_6725,N_3419,N_567);
and U6726 (N_6726,N_572,N_1076);
or U6727 (N_6727,N_3948,N_3117);
or U6728 (N_6728,N_1288,N_245);
nor U6729 (N_6729,N_2009,N_1698);
nor U6730 (N_6730,N_2576,N_1446);
nor U6731 (N_6731,N_3800,N_936);
or U6732 (N_6732,N_1007,N_3140);
nand U6733 (N_6733,N_2659,N_251);
xnor U6734 (N_6734,N_2232,N_2463);
nand U6735 (N_6735,N_2230,N_1608);
nand U6736 (N_6736,N_559,N_1662);
xor U6737 (N_6737,N_188,N_759);
nor U6738 (N_6738,N_3132,N_511);
and U6739 (N_6739,N_3410,N_722);
or U6740 (N_6740,N_783,N_931);
and U6741 (N_6741,N_2677,N_1038);
nand U6742 (N_6742,N_2140,N_3980);
nand U6743 (N_6743,N_1434,N_1265);
and U6744 (N_6744,N_3803,N_1928);
nand U6745 (N_6745,N_2077,N_888);
xnor U6746 (N_6746,N_2532,N_3844);
nand U6747 (N_6747,N_2704,N_1300);
and U6748 (N_6748,N_2557,N_333);
and U6749 (N_6749,N_71,N_2199);
nand U6750 (N_6750,N_765,N_1826);
nand U6751 (N_6751,N_252,N_1555);
or U6752 (N_6752,N_625,N_3466);
nor U6753 (N_6753,N_1869,N_2669);
nand U6754 (N_6754,N_1776,N_2647);
or U6755 (N_6755,N_3370,N_3594);
or U6756 (N_6756,N_500,N_1018);
or U6757 (N_6757,N_3500,N_1007);
nor U6758 (N_6758,N_2997,N_2795);
nor U6759 (N_6759,N_3988,N_2122);
nor U6760 (N_6760,N_3750,N_3913);
nand U6761 (N_6761,N_3725,N_1649);
and U6762 (N_6762,N_3546,N_2324);
and U6763 (N_6763,N_2956,N_2905);
nand U6764 (N_6764,N_3906,N_3372);
and U6765 (N_6765,N_2375,N_291);
or U6766 (N_6766,N_846,N_3117);
nand U6767 (N_6767,N_527,N_715);
xor U6768 (N_6768,N_1531,N_254);
or U6769 (N_6769,N_736,N_1112);
nand U6770 (N_6770,N_2890,N_2976);
xnor U6771 (N_6771,N_2567,N_3031);
nor U6772 (N_6772,N_117,N_1167);
nand U6773 (N_6773,N_1002,N_3474);
or U6774 (N_6774,N_478,N_3127);
nor U6775 (N_6775,N_1352,N_2993);
or U6776 (N_6776,N_3041,N_3662);
or U6777 (N_6777,N_1158,N_857);
or U6778 (N_6778,N_2251,N_1117);
nand U6779 (N_6779,N_498,N_1076);
and U6780 (N_6780,N_452,N_1028);
or U6781 (N_6781,N_1663,N_1928);
nor U6782 (N_6782,N_1211,N_1208);
or U6783 (N_6783,N_38,N_1397);
nor U6784 (N_6784,N_1491,N_1720);
nor U6785 (N_6785,N_3727,N_818);
nor U6786 (N_6786,N_1747,N_299);
or U6787 (N_6787,N_1884,N_1958);
and U6788 (N_6788,N_1957,N_837);
and U6789 (N_6789,N_1059,N_2941);
xor U6790 (N_6790,N_3278,N_1234);
and U6791 (N_6791,N_1281,N_136);
nor U6792 (N_6792,N_3496,N_2048);
and U6793 (N_6793,N_2880,N_2592);
or U6794 (N_6794,N_120,N_1767);
xor U6795 (N_6795,N_3402,N_66);
nor U6796 (N_6796,N_959,N_533);
nor U6797 (N_6797,N_1976,N_3566);
and U6798 (N_6798,N_2454,N_186);
nor U6799 (N_6799,N_1849,N_213);
nand U6800 (N_6800,N_1893,N_238);
and U6801 (N_6801,N_999,N_369);
xnor U6802 (N_6802,N_3919,N_3421);
nor U6803 (N_6803,N_2204,N_2525);
and U6804 (N_6804,N_3866,N_3821);
or U6805 (N_6805,N_542,N_1465);
and U6806 (N_6806,N_2205,N_1610);
nor U6807 (N_6807,N_1893,N_1927);
and U6808 (N_6808,N_2241,N_640);
and U6809 (N_6809,N_3053,N_1123);
or U6810 (N_6810,N_2442,N_812);
nor U6811 (N_6811,N_2670,N_2189);
xor U6812 (N_6812,N_3665,N_3722);
and U6813 (N_6813,N_559,N_3318);
or U6814 (N_6814,N_841,N_828);
and U6815 (N_6815,N_819,N_1489);
or U6816 (N_6816,N_3355,N_474);
nor U6817 (N_6817,N_867,N_579);
nor U6818 (N_6818,N_3553,N_424);
nor U6819 (N_6819,N_3832,N_3532);
nand U6820 (N_6820,N_1843,N_726);
nand U6821 (N_6821,N_1138,N_124);
or U6822 (N_6822,N_853,N_2630);
nand U6823 (N_6823,N_1499,N_444);
nor U6824 (N_6824,N_1585,N_3562);
or U6825 (N_6825,N_1169,N_3368);
and U6826 (N_6826,N_3122,N_3484);
nand U6827 (N_6827,N_1375,N_2528);
and U6828 (N_6828,N_2526,N_2931);
nand U6829 (N_6829,N_1341,N_2658);
nand U6830 (N_6830,N_47,N_400);
nor U6831 (N_6831,N_2935,N_1676);
or U6832 (N_6832,N_2330,N_1994);
or U6833 (N_6833,N_3406,N_3667);
nor U6834 (N_6834,N_142,N_1290);
or U6835 (N_6835,N_3894,N_1059);
or U6836 (N_6836,N_2125,N_1841);
or U6837 (N_6837,N_3644,N_167);
and U6838 (N_6838,N_1918,N_3341);
nor U6839 (N_6839,N_2419,N_1048);
and U6840 (N_6840,N_50,N_3014);
and U6841 (N_6841,N_1957,N_1733);
or U6842 (N_6842,N_2847,N_3040);
and U6843 (N_6843,N_2671,N_1514);
nand U6844 (N_6844,N_1958,N_715);
xnor U6845 (N_6845,N_1456,N_1557);
nor U6846 (N_6846,N_1000,N_283);
or U6847 (N_6847,N_681,N_2578);
nor U6848 (N_6848,N_2884,N_615);
and U6849 (N_6849,N_1608,N_2297);
or U6850 (N_6850,N_3665,N_1007);
nor U6851 (N_6851,N_2516,N_3092);
nand U6852 (N_6852,N_539,N_2932);
nand U6853 (N_6853,N_3457,N_1855);
or U6854 (N_6854,N_3664,N_2208);
nor U6855 (N_6855,N_467,N_1248);
nand U6856 (N_6856,N_387,N_3710);
nor U6857 (N_6857,N_3846,N_22);
and U6858 (N_6858,N_1821,N_433);
nor U6859 (N_6859,N_935,N_1624);
nand U6860 (N_6860,N_80,N_1194);
nor U6861 (N_6861,N_369,N_311);
nand U6862 (N_6862,N_1094,N_2825);
nand U6863 (N_6863,N_2456,N_1565);
or U6864 (N_6864,N_348,N_1436);
xor U6865 (N_6865,N_840,N_3372);
nand U6866 (N_6866,N_1247,N_3940);
or U6867 (N_6867,N_3850,N_3969);
xnor U6868 (N_6868,N_1889,N_3956);
nor U6869 (N_6869,N_3813,N_11);
nand U6870 (N_6870,N_2432,N_1614);
nand U6871 (N_6871,N_1330,N_3020);
xor U6872 (N_6872,N_3279,N_3192);
and U6873 (N_6873,N_3948,N_786);
nand U6874 (N_6874,N_3498,N_1398);
nand U6875 (N_6875,N_3642,N_3554);
or U6876 (N_6876,N_279,N_3757);
and U6877 (N_6877,N_3960,N_2474);
or U6878 (N_6878,N_2154,N_1790);
xnor U6879 (N_6879,N_496,N_384);
nand U6880 (N_6880,N_1824,N_174);
and U6881 (N_6881,N_2871,N_3385);
and U6882 (N_6882,N_3147,N_3081);
and U6883 (N_6883,N_751,N_181);
nand U6884 (N_6884,N_17,N_3418);
nand U6885 (N_6885,N_1454,N_2013);
and U6886 (N_6886,N_1604,N_2042);
nor U6887 (N_6887,N_3597,N_3275);
xor U6888 (N_6888,N_1889,N_1194);
xnor U6889 (N_6889,N_1432,N_2081);
or U6890 (N_6890,N_1511,N_3902);
nand U6891 (N_6891,N_1504,N_3121);
nand U6892 (N_6892,N_3838,N_1833);
nand U6893 (N_6893,N_2460,N_3940);
nor U6894 (N_6894,N_3778,N_3138);
nor U6895 (N_6895,N_1773,N_2976);
nor U6896 (N_6896,N_1280,N_1418);
or U6897 (N_6897,N_53,N_2876);
nor U6898 (N_6898,N_3646,N_585);
or U6899 (N_6899,N_1291,N_3705);
nor U6900 (N_6900,N_3355,N_2592);
or U6901 (N_6901,N_3494,N_3867);
nor U6902 (N_6902,N_975,N_2954);
or U6903 (N_6903,N_741,N_231);
nor U6904 (N_6904,N_3675,N_223);
and U6905 (N_6905,N_3656,N_2965);
nor U6906 (N_6906,N_802,N_1197);
nor U6907 (N_6907,N_3379,N_3046);
nor U6908 (N_6908,N_3176,N_1440);
nand U6909 (N_6909,N_3124,N_3891);
nand U6910 (N_6910,N_2750,N_3080);
or U6911 (N_6911,N_2862,N_2880);
nand U6912 (N_6912,N_3708,N_508);
and U6913 (N_6913,N_2574,N_2007);
xnor U6914 (N_6914,N_231,N_2797);
nand U6915 (N_6915,N_3759,N_3645);
and U6916 (N_6916,N_367,N_294);
nor U6917 (N_6917,N_2518,N_1665);
nand U6918 (N_6918,N_2818,N_3019);
or U6919 (N_6919,N_857,N_1617);
and U6920 (N_6920,N_2469,N_896);
nand U6921 (N_6921,N_304,N_3759);
nand U6922 (N_6922,N_2842,N_3381);
nand U6923 (N_6923,N_1224,N_1384);
nand U6924 (N_6924,N_2707,N_3678);
or U6925 (N_6925,N_422,N_3921);
nand U6926 (N_6926,N_2812,N_985);
nand U6927 (N_6927,N_3935,N_447);
nor U6928 (N_6928,N_2006,N_112);
nand U6929 (N_6929,N_2667,N_1925);
xnor U6930 (N_6930,N_129,N_3575);
and U6931 (N_6931,N_1386,N_2502);
nor U6932 (N_6932,N_471,N_395);
nand U6933 (N_6933,N_3540,N_3530);
nand U6934 (N_6934,N_267,N_3053);
nand U6935 (N_6935,N_823,N_2227);
and U6936 (N_6936,N_3451,N_3475);
nand U6937 (N_6937,N_651,N_3732);
and U6938 (N_6938,N_2155,N_1776);
nor U6939 (N_6939,N_2669,N_3800);
and U6940 (N_6940,N_3425,N_519);
nor U6941 (N_6941,N_638,N_1590);
or U6942 (N_6942,N_3005,N_3308);
nor U6943 (N_6943,N_641,N_3578);
and U6944 (N_6944,N_2800,N_3356);
and U6945 (N_6945,N_204,N_2027);
nor U6946 (N_6946,N_1482,N_3973);
xnor U6947 (N_6947,N_2258,N_518);
xor U6948 (N_6948,N_3821,N_583);
nor U6949 (N_6949,N_106,N_1977);
and U6950 (N_6950,N_434,N_2345);
or U6951 (N_6951,N_1580,N_523);
or U6952 (N_6952,N_2815,N_3453);
xnor U6953 (N_6953,N_1705,N_1310);
and U6954 (N_6954,N_1256,N_3947);
nand U6955 (N_6955,N_325,N_1692);
nor U6956 (N_6956,N_2052,N_898);
nand U6957 (N_6957,N_587,N_2424);
nand U6958 (N_6958,N_182,N_1870);
and U6959 (N_6959,N_3650,N_2000);
or U6960 (N_6960,N_3822,N_706);
or U6961 (N_6961,N_3140,N_2202);
nor U6962 (N_6962,N_3812,N_3114);
xor U6963 (N_6963,N_1956,N_659);
nor U6964 (N_6964,N_3034,N_1983);
or U6965 (N_6965,N_721,N_3745);
nor U6966 (N_6966,N_1302,N_657);
and U6967 (N_6967,N_2438,N_2777);
and U6968 (N_6968,N_212,N_752);
nor U6969 (N_6969,N_1057,N_2287);
nand U6970 (N_6970,N_1583,N_3739);
xnor U6971 (N_6971,N_2913,N_255);
and U6972 (N_6972,N_2214,N_846);
nor U6973 (N_6973,N_3794,N_2775);
and U6974 (N_6974,N_3469,N_1830);
xnor U6975 (N_6975,N_1360,N_692);
nand U6976 (N_6976,N_1237,N_2438);
and U6977 (N_6977,N_3663,N_3440);
nand U6978 (N_6978,N_2228,N_1022);
or U6979 (N_6979,N_3758,N_3994);
xnor U6980 (N_6980,N_1561,N_3328);
and U6981 (N_6981,N_792,N_1638);
and U6982 (N_6982,N_1059,N_538);
xor U6983 (N_6983,N_336,N_2632);
and U6984 (N_6984,N_2425,N_984);
or U6985 (N_6985,N_3946,N_1769);
or U6986 (N_6986,N_1996,N_25);
and U6987 (N_6987,N_1395,N_3454);
or U6988 (N_6988,N_1296,N_3729);
nand U6989 (N_6989,N_3290,N_3722);
nor U6990 (N_6990,N_3358,N_681);
or U6991 (N_6991,N_58,N_665);
or U6992 (N_6992,N_3156,N_2321);
and U6993 (N_6993,N_3968,N_470);
nand U6994 (N_6994,N_3876,N_2129);
and U6995 (N_6995,N_3815,N_1817);
nor U6996 (N_6996,N_2241,N_438);
nand U6997 (N_6997,N_2432,N_1763);
nor U6998 (N_6998,N_334,N_1912);
nand U6999 (N_6999,N_2193,N_290);
or U7000 (N_7000,N_1758,N_3887);
nor U7001 (N_7001,N_711,N_430);
and U7002 (N_7002,N_86,N_578);
or U7003 (N_7003,N_684,N_3231);
nand U7004 (N_7004,N_2353,N_275);
nor U7005 (N_7005,N_3408,N_1811);
and U7006 (N_7006,N_2790,N_710);
nor U7007 (N_7007,N_2291,N_2133);
or U7008 (N_7008,N_2897,N_2169);
nor U7009 (N_7009,N_861,N_2439);
nor U7010 (N_7010,N_2839,N_653);
nor U7011 (N_7011,N_3196,N_1651);
xor U7012 (N_7012,N_1290,N_1640);
xnor U7013 (N_7013,N_3427,N_3079);
nand U7014 (N_7014,N_688,N_2026);
or U7015 (N_7015,N_1118,N_2909);
or U7016 (N_7016,N_1329,N_1540);
and U7017 (N_7017,N_1749,N_3902);
nor U7018 (N_7018,N_3154,N_3139);
or U7019 (N_7019,N_2085,N_3199);
xor U7020 (N_7020,N_347,N_124);
xnor U7021 (N_7021,N_3492,N_3209);
nor U7022 (N_7022,N_3710,N_1687);
or U7023 (N_7023,N_3707,N_729);
nand U7024 (N_7024,N_299,N_3751);
nand U7025 (N_7025,N_3423,N_2407);
nor U7026 (N_7026,N_2562,N_2343);
xor U7027 (N_7027,N_569,N_1805);
nand U7028 (N_7028,N_1478,N_1176);
or U7029 (N_7029,N_647,N_3877);
nor U7030 (N_7030,N_3759,N_1521);
nand U7031 (N_7031,N_3644,N_3700);
and U7032 (N_7032,N_1927,N_2521);
or U7033 (N_7033,N_1205,N_3106);
and U7034 (N_7034,N_2363,N_855);
or U7035 (N_7035,N_795,N_3838);
nor U7036 (N_7036,N_3893,N_238);
nand U7037 (N_7037,N_3673,N_41);
nand U7038 (N_7038,N_463,N_617);
or U7039 (N_7039,N_2338,N_305);
nand U7040 (N_7040,N_1639,N_813);
nand U7041 (N_7041,N_2521,N_15);
nand U7042 (N_7042,N_522,N_3788);
and U7043 (N_7043,N_97,N_978);
nor U7044 (N_7044,N_2124,N_3990);
nor U7045 (N_7045,N_301,N_2770);
or U7046 (N_7046,N_2622,N_1851);
nand U7047 (N_7047,N_90,N_89);
xor U7048 (N_7048,N_2566,N_3963);
nor U7049 (N_7049,N_2912,N_441);
nand U7050 (N_7050,N_2532,N_2773);
nand U7051 (N_7051,N_2986,N_711);
or U7052 (N_7052,N_3264,N_138);
xor U7053 (N_7053,N_400,N_2250);
nand U7054 (N_7054,N_2940,N_2651);
nand U7055 (N_7055,N_1051,N_773);
xor U7056 (N_7056,N_1243,N_2973);
or U7057 (N_7057,N_1187,N_708);
and U7058 (N_7058,N_1946,N_1251);
xnor U7059 (N_7059,N_1906,N_3721);
or U7060 (N_7060,N_1170,N_2291);
nand U7061 (N_7061,N_2346,N_1893);
nand U7062 (N_7062,N_3092,N_3192);
and U7063 (N_7063,N_2632,N_2141);
xor U7064 (N_7064,N_2393,N_311);
or U7065 (N_7065,N_139,N_702);
nand U7066 (N_7066,N_181,N_881);
or U7067 (N_7067,N_1359,N_3156);
or U7068 (N_7068,N_747,N_3027);
nand U7069 (N_7069,N_3593,N_1987);
nand U7070 (N_7070,N_135,N_1775);
or U7071 (N_7071,N_3152,N_1822);
nor U7072 (N_7072,N_3340,N_2635);
nand U7073 (N_7073,N_3238,N_2817);
nand U7074 (N_7074,N_3603,N_158);
or U7075 (N_7075,N_360,N_978);
nor U7076 (N_7076,N_3393,N_3726);
xnor U7077 (N_7077,N_10,N_702);
nor U7078 (N_7078,N_1874,N_2982);
nand U7079 (N_7079,N_389,N_1075);
and U7080 (N_7080,N_3014,N_2336);
xnor U7081 (N_7081,N_2384,N_3792);
and U7082 (N_7082,N_3965,N_431);
or U7083 (N_7083,N_274,N_488);
or U7084 (N_7084,N_3551,N_1092);
nor U7085 (N_7085,N_2579,N_423);
nand U7086 (N_7086,N_3415,N_1688);
xor U7087 (N_7087,N_845,N_2739);
and U7088 (N_7088,N_938,N_779);
and U7089 (N_7089,N_3618,N_2222);
nand U7090 (N_7090,N_3443,N_2126);
nor U7091 (N_7091,N_456,N_2492);
and U7092 (N_7092,N_3129,N_1751);
nor U7093 (N_7093,N_3747,N_440);
xnor U7094 (N_7094,N_3897,N_2422);
and U7095 (N_7095,N_93,N_1039);
or U7096 (N_7096,N_3184,N_2081);
nor U7097 (N_7097,N_652,N_1004);
nand U7098 (N_7098,N_3260,N_1323);
or U7099 (N_7099,N_3510,N_3671);
and U7100 (N_7100,N_2554,N_1369);
nor U7101 (N_7101,N_581,N_2988);
nor U7102 (N_7102,N_3466,N_3682);
nor U7103 (N_7103,N_1630,N_3162);
or U7104 (N_7104,N_647,N_344);
or U7105 (N_7105,N_1390,N_425);
nand U7106 (N_7106,N_867,N_1784);
and U7107 (N_7107,N_2379,N_2324);
nor U7108 (N_7108,N_1986,N_329);
xnor U7109 (N_7109,N_519,N_436);
and U7110 (N_7110,N_1144,N_536);
and U7111 (N_7111,N_2390,N_676);
xnor U7112 (N_7112,N_542,N_2361);
nor U7113 (N_7113,N_215,N_1078);
and U7114 (N_7114,N_16,N_3170);
and U7115 (N_7115,N_703,N_2821);
nor U7116 (N_7116,N_1625,N_2556);
nand U7117 (N_7117,N_788,N_1249);
or U7118 (N_7118,N_1562,N_3592);
or U7119 (N_7119,N_2728,N_872);
and U7120 (N_7120,N_2972,N_3458);
or U7121 (N_7121,N_2098,N_2211);
xor U7122 (N_7122,N_3740,N_1262);
nor U7123 (N_7123,N_3632,N_3354);
and U7124 (N_7124,N_1915,N_740);
xor U7125 (N_7125,N_2567,N_3002);
xor U7126 (N_7126,N_1950,N_3540);
or U7127 (N_7127,N_1612,N_1308);
nand U7128 (N_7128,N_547,N_3053);
xnor U7129 (N_7129,N_507,N_1781);
nor U7130 (N_7130,N_3759,N_389);
and U7131 (N_7131,N_751,N_3249);
or U7132 (N_7132,N_1363,N_1276);
nand U7133 (N_7133,N_1925,N_3230);
and U7134 (N_7134,N_3174,N_2538);
xnor U7135 (N_7135,N_518,N_3780);
or U7136 (N_7136,N_880,N_522);
and U7137 (N_7137,N_3387,N_1593);
nor U7138 (N_7138,N_2013,N_3567);
nor U7139 (N_7139,N_1246,N_3133);
and U7140 (N_7140,N_2110,N_628);
and U7141 (N_7141,N_1013,N_2482);
nor U7142 (N_7142,N_90,N_2419);
nor U7143 (N_7143,N_106,N_3676);
nand U7144 (N_7144,N_2923,N_2485);
nand U7145 (N_7145,N_1976,N_3820);
and U7146 (N_7146,N_1935,N_475);
and U7147 (N_7147,N_2422,N_3099);
or U7148 (N_7148,N_3101,N_1053);
or U7149 (N_7149,N_3192,N_3443);
nand U7150 (N_7150,N_1112,N_1429);
and U7151 (N_7151,N_3380,N_1918);
nor U7152 (N_7152,N_3964,N_949);
nor U7153 (N_7153,N_3090,N_1571);
nand U7154 (N_7154,N_2214,N_3860);
nand U7155 (N_7155,N_1627,N_3923);
or U7156 (N_7156,N_235,N_640);
nor U7157 (N_7157,N_3059,N_2589);
nand U7158 (N_7158,N_3067,N_3799);
nor U7159 (N_7159,N_3529,N_1190);
nor U7160 (N_7160,N_533,N_1207);
or U7161 (N_7161,N_2831,N_995);
and U7162 (N_7162,N_1992,N_3918);
nand U7163 (N_7163,N_3052,N_561);
nand U7164 (N_7164,N_822,N_3529);
nor U7165 (N_7165,N_2466,N_902);
xnor U7166 (N_7166,N_3934,N_3694);
or U7167 (N_7167,N_3588,N_3787);
or U7168 (N_7168,N_1576,N_2712);
nand U7169 (N_7169,N_2667,N_1232);
and U7170 (N_7170,N_2953,N_2442);
nor U7171 (N_7171,N_1200,N_668);
nor U7172 (N_7172,N_1573,N_3299);
nor U7173 (N_7173,N_3349,N_288);
and U7174 (N_7174,N_1650,N_1018);
nand U7175 (N_7175,N_1150,N_210);
or U7176 (N_7176,N_3920,N_2339);
or U7177 (N_7177,N_2604,N_2065);
nand U7178 (N_7178,N_1563,N_2892);
and U7179 (N_7179,N_2854,N_3943);
nand U7180 (N_7180,N_2595,N_572);
nand U7181 (N_7181,N_2223,N_2582);
and U7182 (N_7182,N_3999,N_3257);
xnor U7183 (N_7183,N_1504,N_26);
and U7184 (N_7184,N_3482,N_1645);
and U7185 (N_7185,N_2737,N_3630);
or U7186 (N_7186,N_3321,N_2882);
or U7187 (N_7187,N_3534,N_970);
nand U7188 (N_7188,N_3995,N_913);
nor U7189 (N_7189,N_2988,N_652);
nand U7190 (N_7190,N_1350,N_3557);
or U7191 (N_7191,N_1238,N_2791);
nor U7192 (N_7192,N_1024,N_41);
nor U7193 (N_7193,N_826,N_466);
xnor U7194 (N_7194,N_2716,N_158);
nand U7195 (N_7195,N_3199,N_3253);
xnor U7196 (N_7196,N_2033,N_1121);
and U7197 (N_7197,N_2755,N_81);
or U7198 (N_7198,N_1669,N_295);
or U7199 (N_7199,N_1570,N_689);
nand U7200 (N_7200,N_581,N_2411);
and U7201 (N_7201,N_1872,N_2084);
and U7202 (N_7202,N_3247,N_856);
nand U7203 (N_7203,N_1259,N_1601);
nand U7204 (N_7204,N_2324,N_314);
and U7205 (N_7205,N_2092,N_1169);
and U7206 (N_7206,N_188,N_236);
nand U7207 (N_7207,N_1539,N_849);
xnor U7208 (N_7208,N_754,N_1688);
xor U7209 (N_7209,N_664,N_298);
nor U7210 (N_7210,N_297,N_3489);
nand U7211 (N_7211,N_2767,N_2306);
nor U7212 (N_7212,N_1354,N_2478);
or U7213 (N_7213,N_1680,N_3215);
xor U7214 (N_7214,N_180,N_1230);
nand U7215 (N_7215,N_2924,N_1020);
and U7216 (N_7216,N_2319,N_1466);
nand U7217 (N_7217,N_1078,N_968);
nor U7218 (N_7218,N_3574,N_2015);
or U7219 (N_7219,N_2032,N_1041);
and U7220 (N_7220,N_2343,N_3840);
or U7221 (N_7221,N_3577,N_1091);
nand U7222 (N_7222,N_3177,N_1086);
or U7223 (N_7223,N_801,N_2456);
nand U7224 (N_7224,N_3253,N_2090);
nand U7225 (N_7225,N_10,N_3108);
nand U7226 (N_7226,N_3084,N_1483);
xor U7227 (N_7227,N_1455,N_782);
nand U7228 (N_7228,N_2246,N_1696);
and U7229 (N_7229,N_826,N_948);
xor U7230 (N_7230,N_1531,N_626);
and U7231 (N_7231,N_2673,N_189);
nand U7232 (N_7232,N_692,N_178);
nor U7233 (N_7233,N_2566,N_3378);
and U7234 (N_7234,N_1927,N_3028);
and U7235 (N_7235,N_108,N_2893);
nor U7236 (N_7236,N_1837,N_2004);
nor U7237 (N_7237,N_3941,N_1664);
xor U7238 (N_7238,N_2002,N_987);
and U7239 (N_7239,N_2578,N_2329);
xor U7240 (N_7240,N_462,N_221);
and U7241 (N_7241,N_134,N_1867);
or U7242 (N_7242,N_3933,N_3546);
nor U7243 (N_7243,N_3774,N_3522);
or U7244 (N_7244,N_1924,N_2626);
or U7245 (N_7245,N_596,N_74);
and U7246 (N_7246,N_67,N_1808);
and U7247 (N_7247,N_2361,N_1742);
or U7248 (N_7248,N_2461,N_2143);
and U7249 (N_7249,N_1117,N_2245);
nor U7250 (N_7250,N_1563,N_2080);
nand U7251 (N_7251,N_438,N_1727);
or U7252 (N_7252,N_2680,N_2442);
nor U7253 (N_7253,N_3261,N_3264);
nor U7254 (N_7254,N_3541,N_1344);
nor U7255 (N_7255,N_1453,N_2003);
nor U7256 (N_7256,N_321,N_2035);
or U7257 (N_7257,N_891,N_2680);
nor U7258 (N_7258,N_1520,N_608);
nand U7259 (N_7259,N_1087,N_2953);
xnor U7260 (N_7260,N_2374,N_1467);
nor U7261 (N_7261,N_3515,N_2898);
or U7262 (N_7262,N_3635,N_2740);
xor U7263 (N_7263,N_561,N_144);
or U7264 (N_7264,N_913,N_2046);
nand U7265 (N_7265,N_3101,N_1793);
and U7266 (N_7266,N_0,N_3126);
or U7267 (N_7267,N_2471,N_2434);
and U7268 (N_7268,N_3360,N_2874);
nand U7269 (N_7269,N_303,N_3376);
nor U7270 (N_7270,N_3613,N_957);
nand U7271 (N_7271,N_3320,N_2279);
or U7272 (N_7272,N_2550,N_2199);
nor U7273 (N_7273,N_3804,N_261);
or U7274 (N_7274,N_1183,N_2216);
and U7275 (N_7275,N_3622,N_453);
and U7276 (N_7276,N_1360,N_3206);
nand U7277 (N_7277,N_3605,N_3862);
nor U7278 (N_7278,N_1415,N_2281);
nor U7279 (N_7279,N_3216,N_1961);
xor U7280 (N_7280,N_3655,N_1618);
or U7281 (N_7281,N_3119,N_1530);
xnor U7282 (N_7282,N_831,N_3874);
and U7283 (N_7283,N_1715,N_2171);
nor U7284 (N_7284,N_3587,N_3121);
nor U7285 (N_7285,N_265,N_1118);
and U7286 (N_7286,N_1979,N_730);
nor U7287 (N_7287,N_1106,N_3188);
and U7288 (N_7288,N_3560,N_1798);
nor U7289 (N_7289,N_1902,N_1610);
and U7290 (N_7290,N_634,N_1790);
and U7291 (N_7291,N_1683,N_3658);
nand U7292 (N_7292,N_3235,N_3210);
nand U7293 (N_7293,N_3430,N_3103);
or U7294 (N_7294,N_252,N_1649);
nand U7295 (N_7295,N_1751,N_3070);
and U7296 (N_7296,N_1013,N_443);
or U7297 (N_7297,N_1876,N_451);
or U7298 (N_7298,N_3869,N_1240);
and U7299 (N_7299,N_1925,N_2415);
and U7300 (N_7300,N_1238,N_2971);
or U7301 (N_7301,N_1201,N_2320);
nand U7302 (N_7302,N_1131,N_3596);
or U7303 (N_7303,N_59,N_896);
nand U7304 (N_7304,N_130,N_3627);
and U7305 (N_7305,N_3681,N_3255);
and U7306 (N_7306,N_987,N_729);
xnor U7307 (N_7307,N_854,N_1722);
nor U7308 (N_7308,N_573,N_736);
and U7309 (N_7309,N_2478,N_508);
nand U7310 (N_7310,N_912,N_3392);
or U7311 (N_7311,N_3113,N_3352);
nor U7312 (N_7312,N_829,N_644);
xor U7313 (N_7313,N_1350,N_3221);
or U7314 (N_7314,N_2170,N_3266);
nor U7315 (N_7315,N_3152,N_1485);
nand U7316 (N_7316,N_2828,N_3923);
xnor U7317 (N_7317,N_477,N_299);
nand U7318 (N_7318,N_2495,N_3834);
nor U7319 (N_7319,N_1882,N_450);
xnor U7320 (N_7320,N_3912,N_2864);
nand U7321 (N_7321,N_1720,N_890);
and U7322 (N_7322,N_3839,N_1554);
nor U7323 (N_7323,N_2163,N_1773);
or U7324 (N_7324,N_1176,N_3779);
and U7325 (N_7325,N_760,N_5);
or U7326 (N_7326,N_1354,N_2723);
or U7327 (N_7327,N_2756,N_2892);
xor U7328 (N_7328,N_2845,N_1884);
nand U7329 (N_7329,N_2107,N_3465);
or U7330 (N_7330,N_791,N_1113);
or U7331 (N_7331,N_2676,N_3293);
or U7332 (N_7332,N_2168,N_1138);
nor U7333 (N_7333,N_2679,N_2241);
nand U7334 (N_7334,N_2472,N_3318);
and U7335 (N_7335,N_3852,N_1230);
nand U7336 (N_7336,N_2178,N_3951);
nand U7337 (N_7337,N_1708,N_1270);
and U7338 (N_7338,N_3260,N_3385);
nor U7339 (N_7339,N_301,N_3211);
nand U7340 (N_7340,N_146,N_3706);
and U7341 (N_7341,N_1951,N_3611);
nand U7342 (N_7342,N_527,N_2870);
nor U7343 (N_7343,N_3664,N_3349);
or U7344 (N_7344,N_3194,N_3054);
nor U7345 (N_7345,N_1627,N_3024);
and U7346 (N_7346,N_2382,N_559);
nor U7347 (N_7347,N_1891,N_1837);
nor U7348 (N_7348,N_3859,N_3945);
nand U7349 (N_7349,N_1678,N_875);
xor U7350 (N_7350,N_3329,N_3085);
and U7351 (N_7351,N_139,N_2217);
nand U7352 (N_7352,N_2993,N_1986);
or U7353 (N_7353,N_722,N_415);
or U7354 (N_7354,N_951,N_516);
xnor U7355 (N_7355,N_1402,N_2308);
or U7356 (N_7356,N_2275,N_1926);
and U7357 (N_7357,N_2828,N_3972);
or U7358 (N_7358,N_276,N_3401);
nor U7359 (N_7359,N_1290,N_3875);
xor U7360 (N_7360,N_2183,N_2431);
or U7361 (N_7361,N_1876,N_623);
nor U7362 (N_7362,N_1963,N_1892);
or U7363 (N_7363,N_328,N_3030);
nor U7364 (N_7364,N_1480,N_1337);
nand U7365 (N_7365,N_1983,N_1008);
and U7366 (N_7366,N_2724,N_1637);
nor U7367 (N_7367,N_3434,N_3355);
and U7368 (N_7368,N_1657,N_2850);
and U7369 (N_7369,N_2452,N_3266);
xnor U7370 (N_7370,N_1978,N_3857);
and U7371 (N_7371,N_1068,N_2978);
or U7372 (N_7372,N_2987,N_1351);
or U7373 (N_7373,N_792,N_3849);
xnor U7374 (N_7374,N_28,N_368);
or U7375 (N_7375,N_881,N_386);
or U7376 (N_7376,N_496,N_1198);
or U7377 (N_7377,N_1425,N_3056);
nor U7378 (N_7378,N_1192,N_3916);
nand U7379 (N_7379,N_2986,N_2475);
nand U7380 (N_7380,N_3195,N_534);
nand U7381 (N_7381,N_2069,N_3316);
nor U7382 (N_7382,N_2020,N_2312);
nand U7383 (N_7383,N_2720,N_3120);
and U7384 (N_7384,N_3091,N_359);
nor U7385 (N_7385,N_399,N_1045);
and U7386 (N_7386,N_1146,N_3253);
or U7387 (N_7387,N_3785,N_3129);
and U7388 (N_7388,N_2584,N_1900);
nor U7389 (N_7389,N_1412,N_3755);
or U7390 (N_7390,N_3383,N_3741);
nand U7391 (N_7391,N_3965,N_152);
and U7392 (N_7392,N_930,N_259);
nor U7393 (N_7393,N_3572,N_3515);
or U7394 (N_7394,N_3552,N_1171);
nor U7395 (N_7395,N_3137,N_107);
and U7396 (N_7396,N_3062,N_3837);
nor U7397 (N_7397,N_2802,N_1937);
nand U7398 (N_7398,N_561,N_2635);
and U7399 (N_7399,N_3871,N_2536);
nand U7400 (N_7400,N_1755,N_406);
and U7401 (N_7401,N_1687,N_647);
or U7402 (N_7402,N_3391,N_3153);
or U7403 (N_7403,N_1894,N_1048);
or U7404 (N_7404,N_2257,N_568);
and U7405 (N_7405,N_3231,N_3268);
xnor U7406 (N_7406,N_3680,N_1590);
nor U7407 (N_7407,N_816,N_1318);
and U7408 (N_7408,N_2202,N_1636);
nor U7409 (N_7409,N_2272,N_2486);
or U7410 (N_7410,N_1810,N_1881);
and U7411 (N_7411,N_3245,N_827);
and U7412 (N_7412,N_2922,N_1094);
nand U7413 (N_7413,N_163,N_987);
nor U7414 (N_7414,N_3769,N_2060);
nand U7415 (N_7415,N_2189,N_1667);
or U7416 (N_7416,N_3477,N_3234);
and U7417 (N_7417,N_3305,N_2146);
nand U7418 (N_7418,N_1753,N_3268);
nand U7419 (N_7419,N_1686,N_3763);
or U7420 (N_7420,N_487,N_2211);
nor U7421 (N_7421,N_179,N_2945);
nor U7422 (N_7422,N_3008,N_2997);
or U7423 (N_7423,N_1847,N_329);
nor U7424 (N_7424,N_1765,N_1759);
xnor U7425 (N_7425,N_2545,N_152);
nor U7426 (N_7426,N_2342,N_2410);
nor U7427 (N_7427,N_490,N_806);
or U7428 (N_7428,N_2123,N_738);
nand U7429 (N_7429,N_2160,N_1279);
or U7430 (N_7430,N_1691,N_531);
nand U7431 (N_7431,N_3749,N_1287);
and U7432 (N_7432,N_2623,N_953);
or U7433 (N_7433,N_3839,N_484);
and U7434 (N_7434,N_3028,N_1720);
xnor U7435 (N_7435,N_1520,N_3841);
nor U7436 (N_7436,N_3853,N_3891);
xor U7437 (N_7437,N_3707,N_2333);
nor U7438 (N_7438,N_515,N_1414);
or U7439 (N_7439,N_1907,N_3920);
or U7440 (N_7440,N_3950,N_2011);
or U7441 (N_7441,N_1644,N_1818);
nor U7442 (N_7442,N_3428,N_1944);
nor U7443 (N_7443,N_574,N_3361);
xor U7444 (N_7444,N_84,N_402);
nand U7445 (N_7445,N_2784,N_1093);
nor U7446 (N_7446,N_1990,N_3692);
or U7447 (N_7447,N_3541,N_1066);
nor U7448 (N_7448,N_710,N_825);
nand U7449 (N_7449,N_1871,N_2287);
or U7450 (N_7450,N_507,N_3405);
nor U7451 (N_7451,N_2874,N_3791);
and U7452 (N_7452,N_2722,N_450);
nor U7453 (N_7453,N_2173,N_234);
and U7454 (N_7454,N_1825,N_3263);
xnor U7455 (N_7455,N_3097,N_1188);
nor U7456 (N_7456,N_3523,N_3010);
or U7457 (N_7457,N_457,N_2280);
nand U7458 (N_7458,N_496,N_1930);
or U7459 (N_7459,N_3737,N_1217);
and U7460 (N_7460,N_834,N_717);
nor U7461 (N_7461,N_2995,N_1817);
xor U7462 (N_7462,N_3915,N_1779);
and U7463 (N_7463,N_3177,N_3058);
xnor U7464 (N_7464,N_1777,N_2835);
nor U7465 (N_7465,N_2979,N_3776);
and U7466 (N_7466,N_211,N_624);
and U7467 (N_7467,N_698,N_3532);
or U7468 (N_7468,N_1076,N_2219);
and U7469 (N_7469,N_2301,N_773);
or U7470 (N_7470,N_2143,N_1225);
nor U7471 (N_7471,N_3379,N_1201);
and U7472 (N_7472,N_3016,N_1171);
nand U7473 (N_7473,N_1136,N_2051);
nor U7474 (N_7474,N_1987,N_218);
and U7475 (N_7475,N_61,N_387);
or U7476 (N_7476,N_3710,N_1515);
nor U7477 (N_7477,N_257,N_3958);
nand U7478 (N_7478,N_2925,N_2291);
nor U7479 (N_7479,N_1077,N_3165);
nor U7480 (N_7480,N_1000,N_3697);
or U7481 (N_7481,N_2038,N_2760);
nor U7482 (N_7482,N_1109,N_2615);
nor U7483 (N_7483,N_2907,N_1844);
nand U7484 (N_7484,N_2671,N_2605);
or U7485 (N_7485,N_1282,N_3277);
nor U7486 (N_7486,N_3064,N_2173);
and U7487 (N_7487,N_2779,N_3541);
nand U7488 (N_7488,N_2833,N_3273);
nand U7489 (N_7489,N_3957,N_1750);
and U7490 (N_7490,N_2827,N_3812);
nand U7491 (N_7491,N_2828,N_3673);
and U7492 (N_7492,N_2039,N_1044);
or U7493 (N_7493,N_3206,N_683);
nor U7494 (N_7494,N_650,N_1005);
nand U7495 (N_7495,N_3093,N_3755);
and U7496 (N_7496,N_2329,N_3838);
xnor U7497 (N_7497,N_1647,N_3978);
and U7498 (N_7498,N_1037,N_1980);
and U7499 (N_7499,N_2746,N_3303);
nor U7500 (N_7500,N_543,N_62);
and U7501 (N_7501,N_2328,N_729);
or U7502 (N_7502,N_1659,N_2384);
or U7503 (N_7503,N_1110,N_3653);
nor U7504 (N_7504,N_2523,N_1658);
nor U7505 (N_7505,N_1840,N_3888);
nand U7506 (N_7506,N_1459,N_93);
xnor U7507 (N_7507,N_1484,N_1754);
nor U7508 (N_7508,N_688,N_2894);
and U7509 (N_7509,N_3880,N_514);
nand U7510 (N_7510,N_3200,N_2326);
nand U7511 (N_7511,N_257,N_261);
nor U7512 (N_7512,N_1980,N_3617);
nand U7513 (N_7513,N_757,N_3874);
or U7514 (N_7514,N_3541,N_3477);
nand U7515 (N_7515,N_2614,N_431);
or U7516 (N_7516,N_1518,N_2968);
nor U7517 (N_7517,N_388,N_2608);
and U7518 (N_7518,N_3357,N_2492);
or U7519 (N_7519,N_3540,N_1583);
nand U7520 (N_7520,N_1880,N_301);
and U7521 (N_7521,N_1060,N_1232);
nand U7522 (N_7522,N_2082,N_1618);
and U7523 (N_7523,N_1908,N_441);
and U7524 (N_7524,N_542,N_936);
nand U7525 (N_7525,N_1381,N_836);
and U7526 (N_7526,N_2048,N_2371);
nand U7527 (N_7527,N_1485,N_3254);
nand U7528 (N_7528,N_2975,N_312);
or U7529 (N_7529,N_415,N_3210);
xor U7530 (N_7530,N_1244,N_1002);
nor U7531 (N_7531,N_2097,N_2285);
nor U7532 (N_7532,N_819,N_734);
nand U7533 (N_7533,N_3123,N_2579);
nand U7534 (N_7534,N_46,N_795);
nor U7535 (N_7535,N_194,N_112);
nor U7536 (N_7536,N_1867,N_3561);
or U7537 (N_7537,N_248,N_2081);
nand U7538 (N_7538,N_1504,N_1684);
nor U7539 (N_7539,N_129,N_3301);
nor U7540 (N_7540,N_3179,N_2803);
nor U7541 (N_7541,N_2489,N_2447);
and U7542 (N_7542,N_2701,N_1092);
nand U7543 (N_7543,N_3331,N_1828);
or U7544 (N_7544,N_1553,N_44);
and U7545 (N_7545,N_149,N_60);
or U7546 (N_7546,N_219,N_1729);
nand U7547 (N_7547,N_2924,N_2252);
nand U7548 (N_7548,N_1701,N_3935);
nor U7549 (N_7549,N_49,N_2975);
or U7550 (N_7550,N_1027,N_1410);
nand U7551 (N_7551,N_1951,N_701);
nor U7552 (N_7552,N_708,N_2619);
and U7553 (N_7553,N_862,N_311);
xnor U7554 (N_7554,N_2300,N_3988);
and U7555 (N_7555,N_2229,N_890);
nand U7556 (N_7556,N_3551,N_2163);
and U7557 (N_7557,N_3971,N_1807);
or U7558 (N_7558,N_1119,N_3688);
and U7559 (N_7559,N_3656,N_3158);
nand U7560 (N_7560,N_1932,N_2449);
or U7561 (N_7561,N_1096,N_3609);
nor U7562 (N_7562,N_3974,N_270);
nand U7563 (N_7563,N_1933,N_495);
nand U7564 (N_7564,N_399,N_3915);
or U7565 (N_7565,N_196,N_1983);
and U7566 (N_7566,N_1882,N_2052);
or U7567 (N_7567,N_1445,N_3274);
or U7568 (N_7568,N_1558,N_1000);
or U7569 (N_7569,N_3959,N_3621);
and U7570 (N_7570,N_2391,N_2675);
and U7571 (N_7571,N_746,N_1932);
nor U7572 (N_7572,N_3339,N_2502);
nand U7573 (N_7573,N_2452,N_1567);
nand U7574 (N_7574,N_3944,N_3814);
nand U7575 (N_7575,N_1247,N_2016);
xnor U7576 (N_7576,N_2955,N_595);
or U7577 (N_7577,N_2562,N_780);
or U7578 (N_7578,N_3246,N_3578);
nand U7579 (N_7579,N_927,N_1564);
or U7580 (N_7580,N_1780,N_44);
or U7581 (N_7581,N_1491,N_804);
and U7582 (N_7582,N_2316,N_3176);
nand U7583 (N_7583,N_3823,N_3321);
xnor U7584 (N_7584,N_1223,N_1963);
xnor U7585 (N_7585,N_3548,N_3119);
nor U7586 (N_7586,N_495,N_2066);
nand U7587 (N_7587,N_2279,N_3184);
and U7588 (N_7588,N_138,N_2960);
nor U7589 (N_7589,N_3979,N_683);
and U7590 (N_7590,N_2921,N_1569);
nor U7591 (N_7591,N_3994,N_3246);
xor U7592 (N_7592,N_407,N_1752);
and U7593 (N_7593,N_3686,N_3359);
or U7594 (N_7594,N_638,N_2378);
and U7595 (N_7595,N_525,N_2788);
nand U7596 (N_7596,N_1065,N_1083);
or U7597 (N_7597,N_2802,N_1169);
nor U7598 (N_7598,N_1188,N_2634);
nor U7599 (N_7599,N_2098,N_2735);
and U7600 (N_7600,N_3885,N_2662);
nand U7601 (N_7601,N_1758,N_1500);
nand U7602 (N_7602,N_673,N_941);
nor U7603 (N_7603,N_1574,N_1357);
or U7604 (N_7604,N_1645,N_3186);
and U7605 (N_7605,N_965,N_1288);
nand U7606 (N_7606,N_3931,N_1326);
nand U7607 (N_7607,N_2497,N_2673);
nand U7608 (N_7608,N_117,N_3419);
nor U7609 (N_7609,N_2619,N_2883);
and U7610 (N_7610,N_1987,N_3318);
and U7611 (N_7611,N_3786,N_197);
nor U7612 (N_7612,N_3068,N_616);
nor U7613 (N_7613,N_1536,N_1327);
nor U7614 (N_7614,N_2256,N_740);
and U7615 (N_7615,N_2447,N_3813);
nor U7616 (N_7616,N_1588,N_3384);
nand U7617 (N_7617,N_1833,N_2778);
and U7618 (N_7618,N_3843,N_1947);
nor U7619 (N_7619,N_1341,N_2553);
xor U7620 (N_7620,N_3050,N_1527);
xor U7621 (N_7621,N_3094,N_1630);
and U7622 (N_7622,N_3094,N_3670);
nor U7623 (N_7623,N_548,N_256);
nand U7624 (N_7624,N_2202,N_1650);
and U7625 (N_7625,N_3038,N_1209);
xnor U7626 (N_7626,N_3547,N_2503);
xnor U7627 (N_7627,N_653,N_1981);
nand U7628 (N_7628,N_2294,N_770);
or U7629 (N_7629,N_2665,N_708);
and U7630 (N_7630,N_1527,N_1463);
or U7631 (N_7631,N_225,N_476);
and U7632 (N_7632,N_3646,N_3325);
xnor U7633 (N_7633,N_278,N_2987);
nor U7634 (N_7634,N_81,N_3315);
nand U7635 (N_7635,N_1257,N_3762);
xor U7636 (N_7636,N_2228,N_1819);
or U7637 (N_7637,N_3639,N_1584);
and U7638 (N_7638,N_2860,N_1638);
nor U7639 (N_7639,N_554,N_1071);
or U7640 (N_7640,N_2876,N_3949);
nand U7641 (N_7641,N_2592,N_2531);
nand U7642 (N_7642,N_2146,N_673);
and U7643 (N_7643,N_259,N_3637);
nand U7644 (N_7644,N_1800,N_2686);
or U7645 (N_7645,N_3897,N_1590);
nand U7646 (N_7646,N_1808,N_301);
and U7647 (N_7647,N_1151,N_1454);
and U7648 (N_7648,N_547,N_2233);
and U7649 (N_7649,N_1143,N_2571);
xor U7650 (N_7650,N_3534,N_2011);
and U7651 (N_7651,N_399,N_601);
nor U7652 (N_7652,N_3568,N_206);
and U7653 (N_7653,N_1815,N_1763);
nor U7654 (N_7654,N_3773,N_214);
nor U7655 (N_7655,N_3252,N_3395);
nor U7656 (N_7656,N_2781,N_1384);
nand U7657 (N_7657,N_1625,N_2945);
nor U7658 (N_7658,N_3363,N_843);
or U7659 (N_7659,N_2256,N_352);
and U7660 (N_7660,N_1935,N_79);
nor U7661 (N_7661,N_223,N_650);
nor U7662 (N_7662,N_3817,N_597);
nor U7663 (N_7663,N_3051,N_1940);
or U7664 (N_7664,N_3743,N_1237);
or U7665 (N_7665,N_2082,N_3700);
and U7666 (N_7666,N_1185,N_1663);
nor U7667 (N_7667,N_3189,N_1623);
or U7668 (N_7668,N_3072,N_2138);
or U7669 (N_7669,N_2129,N_1559);
nor U7670 (N_7670,N_369,N_753);
nor U7671 (N_7671,N_1819,N_2840);
and U7672 (N_7672,N_109,N_1902);
nor U7673 (N_7673,N_962,N_143);
nand U7674 (N_7674,N_435,N_386);
xor U7675 (N_7675,N_2074,N_1212);
or U7676 (N_7676,N_2264,N_2473);
nand U7677 (N_7677,N_184,N_77);
and U7678 (N_7678,N_3309,N_2018);
nand U7679 (N_7679,N_2187,N_3093);
or U7680 (N_7680,N_3207,N_1745);
and U7681 (N_7681,N_2254,N_2228);
or U7682 (N_7682,N_903,N_1963);
nor U7683 (N_7683,N_3942,N_586);
nor U7684 (N_7684,N_2286,N_3446);
or U7685 (N_7685,N_166,N_1071);
xnor U7686 (N_7686,N_1640,N_3392);
or U7687 (N_7687,N_1919,N_3285);
nand U7688 (N_7688,N_1687,N_3308);
nor U7689 (N_7689,N_2316,N_544);
nor U7690 (N_7690,N_1906,N_2512);
nor U7691 (N_7691,N_3934,N_3929);
nand U7692 (N_7692,N_3780,N_3996);
nand U7693 (N_7693,N_1162,N_1365);
and U7694 (N_7694,N_1939,N_3174);
nand U7695 (N_7695,N_2555,N_3594);
nor U7696 (N_7696,N_1420,N_1118);
and U7697 (N_7697,N_1275,N_3903);
nor U7698 (N_7698,N_1784,N_3367);
nand U7699 (N_7699,N_220,N_2788);
nor U7700 (N_7700,N_657,N_1004);
nand U7701 (N_7701,N_3072,N_1069);
nand U7702 (N_7702,N_1193,N_132);
xnor U7703 (N_7703,N_3152,N_3056);
nand U7704 (N_7704,N_1301,N_2830);
and U7705 (N_7705,N_3785,N_2010);
or U7706 (N_7706,N_1714,N_681);
nand U7707 (N_7707,N_3180,N_919);
or U7708 (N_7708,N_3616,N_158);
or U7709 (N_7709,N_3958,N_1728);
xnor U7710 (N_7710,N_1741,N_1175);
nand U7711 (N_7711,N_3255,N_3052);
nor U7712 (N_7712,N_3254,N_3936);
nor U7713 (N_7713,N_3538,N_2994);
nor U7714 (N_7714,N_656,N_2935);
xnor U7715 (N_7715,N_3098,N_3148);
nor U7716 (N_7716,N_2620,N_3527);
or U7717 (N_7717,N_1928,N_508);
nand U7718 (N_7718,N_1725,N_3417);
and U7719 (N_7719,N_668,N_682);
or U7720 (N_7720,N_113,N_359);
nand U7721 (N_7721,N_1308,N_1925);
nor U7722 (N_7722,N_2131,N_2436);
and U7723 (N_7723,N_3590,N_2089);
nand U7724 (N_7724,N_1184,N_2810);
and U7725 (N_7725,N_1480,N_3323);
or U7726 (N_7726,N_2174,N_3603);
or U7727 (N_7727,N_3902,N_1539);
or U7728 (N_7728,N_1434,N_2445);
or U7729 (N_7729,N_1504,N_3927);
or U7730 (N_7730,N_27,N_3058);
nor U7731 (N_7731,N_3189,N_3137);
and U7732 (N_7732,N_992,N_3550);
xnor U7733 (N_7733,N_2243,N_1216);
nand U7734 (N_7734,N_1871,N_3709);
nor U7735 (N_7735,N_229,N_1406);
or U7736 (N_7736,N_2993,N_2098);
nor U7737 (N_7737,N_3464,N_3527);
or U7738 (N_7738,N_1817,N_3010);
and U7739 (N_7739,N_1665,N_3394);
nor U7740 (N_7740,N_3681,N_943);
or U7741 (N_7741,N_1436,N_3413);
or U7742 (N_7742,N_3504,N_609);
or U7743 (N_7743,N_1750,N_1833);
nand U7744 (N_7744,N_2707,N_582);
and U7745 (N_7745,N_1356,N_3033);
and U7746 (N_7746,N_2955,N_1492);
nor U7747 (N_7747,N_825,N_3399);
nand U7748 (N_7748,N_268,N_3707);
or U7749 (N_7749,N_727,N_2995);
and U7750 (N_7750,N_1935,N_1463);
and U7751 (N_7751,N_3574,N_2551);
nor U7752 (N_7752,N_3747,N_464);
nor U7753 (N_7753,N_1008,N_3174);
or U7754 (N_7754,N_317,N_568);
nor U7755 (N_7755,N_1976,N_79);
nor U7756 (N_7756,N_3647,N_3643);
and U7757 (N_7757,N_3438,N_2100);
nor U7758 (N_7758,N_23,N_2872);
and U7759 (N_7759,N_3222,N_517);
nand U7760 (N_7760,N_102,N_2785);
nand U7761 (N_7761,N_3814,N_207);
nand U7762 (N_7762,N_2515,N_108);
xor U7763 (N_7763,N_1798,N_611);
nand U7764 (N_7764,N_1880,N_0);
nor U7765 (N_7765,N_3844,N_701);
and U7766 (N_7766,N_343,N_3284);
or U7767 (N_7767,N_1621,N_2816);
and U7768 (N_7768,N_3500,N_2188);
nor U7769 (N_7769,N_3867,N_3014);
and U7770 (N_7770,N_1823,N_2211);
xnor U7771 (N_7771,N_3183,N_88);
nand U7772 (N_7772,N_2676,N_2336);
and U7773 (N_7773,N_3365,N_1261);
and U7774 (N_7774,N_1100,N_3548);
nor U7775 (N_7775,N_1099,N_366);
and U7776 (N_7776,N_2231,N_527);
or U7777 (N_7777,N_2205,N_2801);
xor U7778 (N_7778,N_912,N_3102);
and U7779 (N_7779,N_525,N_3443);
and U7780 (N_7780,N_3272,N_3167);
and U7781 (N_7781,N_117,N_705);
and U7782 (N_7782,N_3830,N_2894);
or U7783 (N_7783,N_1461,N_3593);
xor U7784 (N_7784,N_822,N_3566);
nand U7785 (N_7785,N_2278,N_3848);
and U7786 (N_7786,N_3543,N_988);
nand U7787 (N_7787,N_124,N_1149);
or U7788 (N_7788,N_1557,N_3605);
or U7789 (N_7789,N_1894,N_760);
nand U7790 (N_7790,N_698,N_3683);
or U7791 (N_7791,N_1595,N_3958);
and U7792 (N_7792,N_2466,N_385);
and U7793 (N_7793,N_2392,N_847);
xor U7794 (N_7794,N_1391,N_88);
or U7795 (N_7795,N_1650,N_2945);
or U7796 (N_7796,N_745,N_1445);
or U7797 (N_7797,N_3793,N_1223);
xor U7798 (N_7798,N_2740,N_2280);
nor U7799 (N_7799,N_2692,N_538);
nor U7800 (N_7800,N_2477,N_2121);
and U7801 (N_7801,N_2355,N_2530);
and U7802 (N_7802,N_774,N_2998);
and U7803 (N_7803,N_3661,N_3529);
nor U7804 (N_7804,N_634,N_1018);
and U7805 (N_7805,N_2940,N_2583);
and U7806 (N_7806,N_786,N_862);
and U7807 (N_7807,N_851,N_1486);
and U7808 (N_7808,N_2114,N_2928);
or U7809 (N_7809,N_2962,N_718);
and U7810 (N_7810,N_740,N_169);
xnor U7811 (N_7811,N_2243,N_2791);
xor U7812 (N_7812,N_2,N_363);
or U7813 (N_7813,N_1820,N_2124);
nor U7814 (N_7814,N_415,N_1531);
or U7815 (N_7815,N_930,N_452);
nand U7816 (N_7816,N_1999,N_3174);
and U7817 (N_7817,N_1993,N_3134);
nand U7818 (N_7818,N_1660,N_3571);
or U7819 (N_7819,N_1739,N_2529);
or U7820 (N_7820,N_1375,N_2971);
and U7821 (N_7821,N_661,N_2807);
nor U7822 (N_7822,N_650,N_648);
nor U7823 (N_7823,N_1058,N_2605);
nand U7824 (N_7824,N_3632,N_3081);
or U7825 (N_7825,N_3320,N_3973);
or U7826 (N_7826,N_1009,N_2046);
nand U7827 (N_7827,N_3614,N_1295);
xor U7828 (N_7828,N_2936,N_942);
nor U7829 (N_7829,N_135,N_1789);
nand U7830 (N_7830,N_2538,N_1882);
nor U7831 (N_7831,N_2497,N_2709);
or U7832 (N_7832,N_1311,N_833);
xnor U7833 (N_7833,N_2622,N_3600);
or U7834 (N_7834,N_1024,N_3299);
nand U7835 (N_7835,N_3410,N_59);
or U7836 (N_7836,N_2617,N_850);
and U7837 (N_7837,N_990,N_311);
and U7838 (N_7838,N_3512,N_2063);
nand U7839 (N_7839,N_2444,N_3552);
xor U7840 (N_7840,N_1759,N_1293);
and U7841 (N_7841,N_3603,N_3352);
nor U7842 (N_7842,N_3523,N_1518);
and U7843 (N_7843,N_1377,N_2667);
nand U7844 (N_7844,N_2657,N_373);
and U7845 (N_7845,N_1935,N_3177);
or U7846 (N_7846,N_2294,N_162);
and U7847 (N_7847,N_528,N_33);
nor U7848 (N_7848,N_810,N_845);
and U7849 (N_7849,N_1154,N_3619);
nand U7850 (N_7850,N_2993,N_2377);
and U7851 (N_7851,N_2600,N_2590);
or U7852 (N_7852,N_632,N_2849);
and U7853 (N_7853,N_2462,N_1712);
xor U7854 (N_7854,N_1122,N_640);
xnor U7855 (N_7855,N_222,N_475);
nand U7856 (N_7856,N_3087,N_2193);
nand U7857 (N_7857,N_596,N_2472);
nor U7858 (N_7858,N_827,N_3113);
nand U7859 (N_7859,N_3739,N_720);
and U7860 (N_7860,N_1679,N_3771);
or U7861 (N_7861,N_301,N_1026);
and U7862 (N_7862,N_3471,N_3636);
nand U7863 (N_7863,N_2339,N_2780);
nand U7864 (N_7864,N_1631,N_875);
nor U7865 (N_7865,N_1869,N_2608);
or U7866 (N_7866,N_814,N_388);
and U7867 (N_7867,N_492,N_2215);
or U7868 (N_7868,N_2694,N_3175);
or U7869 (N_7869,N_823,N_1904);
nor U7870 (N_7870,N_2222,N_998);
nor U7871 (N_7871,N_3594,N_262);
nor U7872 (N_7872,N_1197,N_3795);
and U7873 (N_7873,N_3840,N_2009);
nor U7874 (N_7874,N_1561,N_2469);
nor U7875 (N_7875,N_3740,N_1528);
and U7876 (N_7876,N_1970,N_1187);
or U7877 (N_7877,N_692,N_288);
or U7878 (N_7878,N_2281,N_2908);
nor U7879 (N_7879,N_1016,N_80);
nor U7880 (N_7880,N_2939,N_2415);
nand U7881 (N_7881,N_3878,N_2552);
and U7882 (N_7882,N_3067,N_3014);
nor U7883 (N_7883,N_3055,N_1528);
and U7884 (N_7884,N_2661,N_152);
nor U7885 (N_7885,N_51,N_1620);
nor U7886 (N_7886,N_2580,N_2550);
nand U7887 (N_7887,N_3643,N_415);
or U7888 (N_7888,N_300,N_921);
xor U7889 (N_7889,N_3147,N_543);
or U7890 (N_7890,N_268,N_1954);
nand U7891 (N_7891,N_1097,N_810);
or U7892 (N_7892,N_1711,N_495);
nor U7893 (N_7893,N_1923,N_2661);
and U7894 (N_7894,N_338,N_1215);
or U7895 (N_7895,N_2006,N_1406);
xnor U7896 (N_7896,N_1729,N_2946);
xnor U7897 (N_7897,N_441,N_3150);
xnor U7898 (N_7898,N_958,N_228);
nand U7899 (N_7899,N_532,N_2420);
and U7900 (N_7900,N_3773,N_3187);
nor U7901 (N_7901,N_2399,N_3244);
nor U7902 (N_7902,N_2078,N_1616);
and U7903 (N_7903,N_1073,N_580);
or U7904 (N_7904,N_1910,N_24);
or U7905 (N_7905,N_945,N_518);
and U7906 (N_7906,N_2311,N_2383);
nand U7907 (N_7907,N_2345,N_1830);
nand U7908 (N_7908,N_3720,N_2064);
and U7909 (N_7909,N_3065,N_770);
nor U7910 (N_7910,N_1606,N_1136);
xor U7911 (N_7911,N_719,N_717);
or U7912 (N_7912,N_3837,N_3537);
or U7913 (N_7913,N_56,N_2806);
nor U7914 (N_7914,N_3623,N_399);
nor U7915 (N_7915,N_1810,N_2646);
and U7916 (N_7916,N_1341,N_2608);
nor U7917 (N_7917,N_1667,N_976);
or U7918 (N_7918,N_3229,N_71);
nand U7919 (N_7919,N_3227,N_240);
or U7920 (N_7920,N_2933,N_379);
or U7921 (N_7921,N_969,N_2390);
nor U7922 (N_7922,N_3709,N_1348);
and U7923 (N_7923,N_2967,N_3992);
and U7924 (N_7924,N_2691,N_1369);
nor U7925 (N_7925,N_2105,N_3446);
or U7926 (N_7926,N_843,N_982);
nand U7927 (N_7927,N_1715,N_2289);
nand U7928 (N_7928,N_3024,N_640);
or U7929 (N_7929,N_1451,N_2427);
nand U7930 (N_7930,N_516,N_2681);
and U7931 (N_7931,N_1414,N_2800);
or U7932 (N_7932,N_2779,N_2679);
nor U7933 (N_7933,N_3668,N_2347);
nand U7934 (N_7934,N_2944,N_3091);
nand U7935 (N_7935,N_3285,N_1084);
nand U7936 (N_7936,N_3225,N_1541);
or U7937 (N_7937,N_620,N_2766);
xnor U7938 (N_7938,N_517,N_1667);
nor U7939 (N_7939,N_695,N_4);
xnor U7940 (N_7940,N_863,N_3642);
or U7941 (N_7941,N_2952,N_1328);
or U7942 (N_7942,N_132,N_3587);
nand U7943 (N_7943,N_3157,N_961);
nor U7944 (N_7944,N_2211,N_852);
xor U7945 (N_7945,N_3025,N_3071);
nor U7946 (N_7946,N_2002,N_2083);
or U7947 (N_7947,N_1767,N_610);
or U7948 (N_7948,N_149,N_3809);
nand U7949 (N_7949,N_1119,N_2379);
and U7950 (N_7950,N_787,N_3028);
nor U7951 (N_7951,N_3834,N_135);
and U7952 (N_7952,N_3286,N_102);
nand U7953 (N_7953,N_779,N_254);
or U7954 (N_7954,N_3354,N_557);
nand U7955 (N_7955,N_2363,N_877);
or U7956 (N_7956,N_980,N_2173);
and U7957 (N_7957,N_1159,N_1201);
and U7958 (N_7958,N_3372,N_1488);
nor U7959 (N_7959,N_1043,N_1046);
nor U7960 (N_7960,N_1663,N_2828);
xor U7961 (N_7961,N_28,N_2817);
nor U7962 (N_7962,N_1504,N_1110);
or U7963 (N_7963,N_1813,N_1463);
nand U7964 (N_7964,N_3327,N_2779);
or U7965 (N_7965,N_2302,N_2910);
nor U7966 (N_7966,N_1569,N_1715);
nor U7967 (N_7967,N_1182,N_1642);
nand U7968 (N_7968,N_3538,N_1947);
xnor U7969 (N_7969,N_2992,N_3457);
nor U7970 (N_7970,N_2475,N_2890);
and U7971 (N_7971,N_0,N_3143);
nand U7972 (N_7972,N_3492,N_1446);
nor U7973 (N_7973,N_1037,N_3592);
nor U7974 (N_7974,N_2539,N_652);
or U7975 (N_7975,N_1987,N_558);
and U7976 (N_7976,N_3244,N_988);
or U7977 (N_7977,N_1751,N_2034);
xor U7978 (N_7978,N_2668,N_3423);
or U7979 (N_7979,N_2157,N_3158);
nor U7980 (N_7980,N_1289,N_1482);
or U7981 (N_7981,N_132,N_833);
and U7982 (N_7982,N_1406,N_2197);
nor U7983 (N_7983,N_751,N_3141);
nand U7984 (N_7984,N_3883,N_1462);
and U7985 (N_7985,N_1470,N_1591);
nand U7986 (N_7986,N_3249,N_3296);
or U7987 (N_7987,N_1156,N_1744);
xor U7988 (N_7988,N_3312,N_978);
nand U7989 (N_7989,N_1536,N_3728);
or U7990 (N_7990,N_2679,N_3204);
xor U7991 (N_7991,N_858,N_442);
nor U7992 (N_7992,N_2845,N_1075);
and U7993 (N_7993,N_1887,N_3567);
or U7994 (N_7994,N_2300,N_2728);
nor U7995 (N_7995,N_625,N_147);
nand U7996 (N_7996,N_1692,N_806);
and U7997 (N_7997,N_3148,N_296);
and U7998 (N_7998,N_116,N_1295);
nand U7999 (N_7999,N_3996,N_1655);
or U8000 (N_8000,N_6234,N_6021);
nor U8001 (N_8001,N_6174,N_5335);
xnor U8002 (N_8002,N_7393,N_6548);
nand U8003 (N_8003,N_5851,N_5937);
and U8004 (N_8004,N_5381,N_6982);
and U8005 (N_8005,N_5104,N_6339);
or U8006 (N_8006,N_4905,N_7784);
or U8007 (N_8007,N_7668,N_4643);
or U8008 (N_8008,N_7652,N_5622);
nand U8009 (N_8009,N_4511,N_7759);
and U8010 (N_8010,N_5441,N_5052);
nand U8011 (N_8011,N_5110,N_6360);
nand U8012 (N_8012,N_6652,N_6611);
or U8013 (N_8013,N_6004,N_5339);
nand U8014 (N_8014,N_5760,N_7565);
or U8015 (N_8015,N_4428,N_7206);
nor U8016 (N_8016,N_7514,N_4683);
and U8017 (N_8017,N_4531,N_4030);
and U8018 (N_8018,N_7821,N_5037);
nand U8019 (N_8019,N_7405,N_5227);
xnor U8020 (N_8020,N_7458,N_6162);
nand U8021 (N_8021,N_4677,N_4150);
xnor U8022 (N_8022,N_5428,N_6210);
nand U8023 (N_8023,N_5567,N_6328);
and U8024 (N_8024,N_6878,N_4353);
and U8025 (N_8025,N_5089,N_4293);
xnor U8026 (N_8026,N_7991,N_5855);
nor U8027 (N_8027,N_5954,N_4480);
or U8028 (N_8028,N_6736,N_4751);
or U8029 (N_8029,N_6421,N_5880);
nand U8030 (N_8030,N_5312,N_7208);
nand U8031 (N_8031,N_4957,N_5891);
nor U8032 (N_8032,N_5776,N_5009);
and U8033 (N_8033,N_4354,N_6791);
nand U8034 (N_8034,N_7920,N_6465);
nor U8035 (N_8035,N_4307,N_7533);
and U8036 (N_8036,N_4926,N_6017);
nand U8037 (N_8037,N_5158,N_4109);
nand U8038 (N_8038,N_7748,N_7572);
or U8039 (N_8039,N_7142,N_6294);
or U8040 (N_8040,N_6940,N_5848);
or U8041 (N_8041,N_4686,N_5644);
and U8042 (N_8042,N_5006,N_4372);
nand U8043 (N_8043,N_7765,N_5296);
or U8044 (N_8044,N_4871,N_5723);
or U8045 (N_8045,N_6515,N_6894);
nor U8046 (N_8046,N_6077,N_4043);
xor U8047 (N_8047,N_7425,N_7223);
or U8048 (N_8048,N_5191,N_5958);
and U8049 (N_8049,N_6400,N_4908);
nor U8050 (N_8050,N_5002,N_6965);
nand U8051 (N_8051,N_4029,N_6680);
xor U8052 (N_8052,N_4430,N_4093);
and U8053 (N_8053,N_4964,N_5933);
nor U8054 (N_8054,N_6132,N_5968);
nor U8055 (N_8055,N_4861,N_6527);
or U8056 (N_8056,N_7104,N_6186);
nand U8057 (N_8057,N_5430,N_6641);
and U8058 (N_8058,N_4987,N_6441);
or U8059 (N_8059,N_7253,N_6484);
and U8060 (N_8060,N_5143,N_5361);
and U8061 (N_8061,N_4989,N_6771);
nor U8062 (N_8062,N_4786,N_7723);
xor U8063 (N_8063,N_5539,N_4244);
and U8064 (N_8064,N_6322,N_6623);
nand U8065 (N_8065,N_5198,N_6840);
nand U8066 (N_8066,N_6414,N_7460);
or U8067 (N_8067,N_7640,N_6737);
nor U8068 (N_8068,N_5627,N_6738);
nand U8069 (N_8069,N_5400,N_6825);
and U8070 (N_8070,N_6806,N_4838);
nand U8071 (N_8071,N_6459,N_6601);
nor U8072 (N_8072,N_7065,N_5168);
nand U8073 (N_8073,N_5688,N_7793);
nor U8074 (N_8074,N_5226,N_6659);
and U8075 (N_8075,N_5549,N_6143);
and U8076 (N_8076,N_5307,N_7710);
nor U8077 (N_8077,N_5086,N_4586);
or U8078 (N_8078,N_5444,N_7694);
xor U8079 (N_8079,N_4077,N_4363);
nor U8080 (N_8080,N_4993,N_5249);
nor U8081 (N_8081,N_7676,N_4384);
or U8082 (N_8082,N_4065,N_5738);
and U8083 (N_8083,N_7165,N_4489);
and U8084 (N_8084,N_7919,N_5016);
xor U8085 (N_8085,N_4562,N_5453);
xor U8086 (N_8086,N_4919,N_5893);
or U8087 (N_8087,N_6585,N_6408);
and U8088 (N_8088,N_4950,N_4979);
and U8089 (N_8089,N_5969,N_6745);
or U8090 (N_8090,N_5011,N_6325);
nand U8091 (N_8091,N_4546,N_6110);
nand U8092 (N_8092,N_7121,N_4529);
nand U8093 (N_8093,N_5753,N_7896);
or U8094 (N_8094,N_7207,N_4212);
nand U8095 (N_8095,N_7977,N_4120);
nand U8096 (N_8096,N_7270,N_6241);
or U8097 (N_8097,N_7578,N_5140);
nand U8098 (N_8098,N_6751,N_6502);
or U8099 (N_8099,N_4581,N_6253);
nand U8100 (N_8100,N_7587,N_7147);
xor U8101 (N_8101,N_5984,N_7268);
or U8102 (N_8102,N_4717,N_5945);
nand U8103 (N_8103,N_7833,N_7297);
or U8104 (N_8104,N_4321,N_6897);
nor U8105 (N_8105,N_5693,N_4361);
and U8106 (N_8106,N_5625,N_4323);
nand U8107 (N_8107,N_5565,N_6196);
nor U8108 (N_8108,N_7382,N_4854);
and U8109 (N_8109,N_6813,N_5548);
and U8110 (N_8110,N_6910,N_7352);
xor U8111 (N_8111,N_4659,N_4375);
or U8112 (N_8112,N_7626,N_4213);
nand U8113 (N_8113,N_4742,N_6353);
and U8114 (N_8114,N_5390,N_6563);
nand U8115 (N_8115,N_5422,N_6352);
and U8116 (N_8116,N_7842,N_7944);
and U8117 (N_8117,N_5317,N_6921);
nor U8118 (N_8118,N_6090,N_5239);
xor U8119 (N_8119,N_4167,N_6428);
nor U8120 (N_8120,N_4526,N_4470);
nand U8121 (N_8121,N_7687,N_6372);
and U8122 (N_8122,N_5481,N_4154);
xnor U8123 (N_8123,N_7952,N_7247);
or U8124 (N_8124,N_6158,N_6541);
or U8125 (N_8125,N_7851,N_7138);
nor U8126 (N_8126,N_6349,N_5582);
nor U8127 (N_8127,N_5202,N_4235);
xnor U8128 (N_8128,N_5150,N_5781);
nand U8129 (N_8129,N_5777,N_6514);
xor U8130 (N_8130,N_7998,N_7588);
or U8131 (N_8131,N_4798,N_5613);
nand U8132 (N_8132,N_5094,N_6833);
and U8133 (N_8133,N_5939,N_7342);
nand U8134 (N_8134,N_6284,N_4118);
and U8135 (N_8135,N_5664,N_5176);
xor U8136 (N_8136,N_5656,N_7251);
and U8137 (N_8137,N_6307,N_6521);
nand U8138 (N_8138,N_5008,N_7701);
nand U8139 (N_8139,N_6775,N_4910);
or U8140 (N_8140,N_6370,N_5208);
and U8141 (N_8141,N_7126,N_5899);
or U8142 (N_8142,N_5780,N_4945);
nor U8143 (N_8143,N_4924,N_6547);
or U8144 (N_8144,N_5145,N_5064);
and U8145 (N_8145,N_7880,N_7642);
nor U8146 (N_8146,N_7924,N_5683);
or U8147 (N_8147,N_6655,N_5185);
and U8148 (N_8148,N_6823,N_7937);
and U8149 (N_8149,N_5531,N_4792);
xor U8150 (N_8150,N_4911,N_4644);
nand U8151 (N_8151,N_7261,N_6313);
or U8152 (N_8152,N_6262,N_6803);
and U8153 (N_8153,N_7431,N_6707);
nor U8154 (N_8154,N_4149,N_6092);
nand U8155 (N_8155,N_6069,N_7331);
nor U8156 (N_8156,N_5618,N_6340);
xnor U8157 (N_8157,N_4498,N_6014);
xnor U8158 (N_8158,N_5343,N_5655);
nand U8159 (N_8159,N_7507,N_7579);
nand U8160 (N_8160,N_4007,N_6801);
xor U8161 (N_8161,N_6213,N_7461);
nand U8162 (N_8162,N_4523,N_5234);
and U8163 (N_8163,N_4638,N_6617);
nor U8164 (N_8164,N_6175,N_4815);
nor U8165 (N_8165,N_4730,N_6012);
xor U8166 (N_8166,N_6198,N_6734);
nor U8167 (N_8167,N_4210,N_5579);
xnor U8168 (N_8168,N_7362,N_6148);
xor U8169 (N_8169,N_7894,N_5333);
nor U8170 (N_8170,N_6804,N_6867);
or U8171 (N_8171,N_4600,N_6396);
and U8172 (N_8172,N_4934,N_7738);
or U8173 (N_8173,N_4432,N_7190);
or U8174 (N_8174,N_5213,N_6634);
and U8175 (N_8175,N_7446,N_7941);
and U8176 (N_8176,N_5915,N_7289);
nor U8177 (N_8177,N_6391,N_5261);
and U8178 (N_8178,N_6251,N_4483);
and U8179 (N_8179,N_6819,N_4646);
or U8180 (N_8180,N_6487,N_6651);
or U8181 (N_8181,N_5587,N_7319);
xnor U8182 (N_8182,N_6821,N_7503);
or U8183 (N_8183,N_4334,N_4294);
and U8184 (N_8184,N_5259,N_5906);
or U8185 (N_8185,N_5812,N_5236);
nor U8186 (N_8186,N_7046,N_6298);
or U8187 (N_8187,N_7561,N_7210);
xnor U8188 (N_8188,N_4814,N_6336);
or U8189 (N_8189,N_5133,N_6233);
nor U8190 (N_8190,N_7231,N_4999);
or U8191 (N_8191,N_6893,N_6619);
nor U8192 (N_8192,N_5815,N_4982);
nor U8193 (N_8193,N_6691,N_5269);
nor U8194 (N_8194,N_7810,N_6777);
and U8195 (N_8195,N_7275,N_7848);
nand U8196 (N_8196,N_7856,N_7013);
nor U8197 (N_8197,N_5147,N_7334);
nor U8198 (N_8198,N_4469,N_6979);
nand U8199 (N_8199,N_7504,N_4147);
nand U8200 (N_8200,N_6928,N_6224);
and U8201 (N_8201,N_4055,N_4909);
and U8202 (N_8202,N_7288,N_5817);
and U8203 (N_8203,N_4699,N_4128);
or U8204 (N_8204,N_7908,N_7695);
nand U8205 (N_8205,N_4094,N_5602);
or U8206 (N_8206,N_4124,N_7513);
nor U8207 (N_8207,N_4368,N_5106);
nor U8208 (N_8208,N_6333,N_4448);
nor U8209 (N_8209,N_5454,N_6693);
and U8210 (N_8210,N_6113,N_7990);
nand U8211 (N_8211,N_7538,N_5493);
nand U8212 (N_8212,N_7753,N_6495);
xnor U8213 (N_8213,N_6503,N_7160);
and U8214 (N_8214,N_6104,N_7867);
and U8215 (N_8215,N_6057,N_7246);
and U8216 (N_8216,N_6816,N_4169);
or U8217 (N_8217,N_6705,N_4411);
and U8218 (N_8218,N_4605,N_7512);
nand U8219 (N_8219,N_7408,N_7492);
or U8220 (N_8220,N_4178,N_5300);
and U8221 (N_8221,N_6319,N_7844);
xnor U8222 (N_8222,N_4484,N_5540);
and U8223 (N_8223,N_6448,N_6572);
nor U8224 (N_8224,N_6443,N_4870);
nand U8225 (N_8225,N_4920,N_4975);
or U8226 (N_8226,N_4338,N_7674);
and U8227 (N_8227,N_7024,N_5669);
nor U8228 (N_8228,N_6781,N_4679);
or U8229 (N_8229,N_7644,N_7700);
nand U8230 (N_8230,N_6366,N_6130);
or U8231 (N_8231,N_6712,N_4016);
nand U8232 (N_8232,N_4512,N_7549);
or U8233 (N_8233,N_6907,N_4245);
xnor U8234 (N_8234,N_6157,N_4085);
and U8235 (N_8235,N_4041,N_4276);
nand U8236 (N_8236,N_7789,N_4104);
nand U8237 (N_8237,N_6163,N_4764);
or U8238 (N_8238,N_7974,N_5763);
nor U8239 (N_8239,N_5134,N_5291);
xor U8240 (N_8240,N_7455,N_5347);
nor U8241 (N_8241,N_6031,N_6598);
nor U8242 (N_8242,N_7375,N_4239);
nand U8243 (N_8243,N_7332,N_5120);
or U8244 (N_8244,N_5866,N_4032);
nand U8245 (N_8245,N_5066,N_5792);
and U8246 (N_8246,N_6675,N_6365);
nor U8247 (N_8247,N_4892,N_5524);
nor U8248 (N_8248,N_7711,N_7778);
nor U8249 (N_8249,N_5964,N_5243);
and U8250 (N_8250,N_4602,N_4330);
xor U8251 (N_8251,N_4986,N_5476);
nor U8252 (N_8252,N_7258,N_5165);
or U8253 (N_8253,N_6433,N_5405);
nand U8254 (N_8254,N_4702,N_4025);
or U8255 (N_8255,N_5636,N_4896);
xor U8256 (N_8256,N_4132,N_7547);
or U8257 (N_8257,N_4027,N_6106);
or U8258 (N_8258,N_5729,N_5330);
nor U8259 (N_8259,N_4355,N_4127);
nor U8260 (N_8260,N_7448,N_6604);
or U8261 (N_8261,N_4860,N_7073);
xor U8262 (N_8262,N_4535,N_5180);
or U8263 (N_8263,N_7038,N_7598);
xnor U8264 (N_8264,N_7757,N_6694);
and U8265 (N_8265,N_6373,N_6794);
xnor U8266 (N_8266,N_5502,N_7806);
or U8267 (N_8267,N_5975,N_4876);
nor U8268 (N_8268,N_7645,N_7389);
or U8269 (N_8269,N_5003,N_7916);
xnor U8270 (N_8270,N_7675,N_6729);
nand U8271 (N_8271,N_4705,N_4386);
or U8272 (N_8272,N_4096,N_7020);
nor U8273 (N_8273,N_5124,N_5705);
nor U8274 (N_8274,N_5038,N_4273);
xnor U8275 (N_8275,N_7797,N_5256);
xor U8276 (N_8276,N_4655,N_5995);
or U8277 (N_8277,N_5513,N_7294);
nor U8278 (N_8278,N_6037,N_6599);
nand U8279 (N_8279,N_6149,N_7387);
and U8280 (N_8280,N_4112,N_4229);
or U8281 (N_8281,N_7752,N_4394);
nor U8282 (N_8282,N_5398,N_6131);
nand U8283 (N_8283,N_7545,N_6756);
and U8284 (N_8284,N_5316,N_4853);
nand U8285 (N_8285,N_4847,N_7080);
nor U8286 (N_8286,N_4929,N_6039);
nor U8287 (N_8287,N_5241,N_4116);
nor U8288 (N_8288,N_6159,N_6024);
nand U8289 (N_8289,N_5341,N_6197);
xor U8290 (N_8290,N_4520,N_5950);
nor U8291 (N_8291,N_4339,N_6882);
and U8292 (N_8292,N_5963,N_6595);
nand U8293 (N_8293,N_6466,N_7730);
or U8294 (N_8294,N_4665,N_5161);
nand U8295 (N_8295,N_7282,N_7067);
nor U8296 (N_8296,N_4505,N_4251);
or U8297 (N_8297,N_7917,N_6123);
nand U8298 (N_8298,N_6948,N_6941);
nand U8299 (N_8299,N_4305,N_6918);
and U8300 (N_8300,N_7438,N_5581);
and U8301 (N_8301,N_6172,N_6864);
or U8302 (N_8302,N_5834,N_5114);
nand U8303 (N_8303,N_7415,N_7279);
nand U8304 (N_8304,N_4687,N_5860);
or U8305 (N_8305,N_6915,N_6597);
nand U8306 (N_8306,N_7592,N_4227);
nand U8307 (N_8307,N_4021,N_4201);
and U8308 (N_8308,N_6925,N_7324);
or U8309 (N_8309,N_5634,N_7427);
xor U8310 (N_8310,N_5835,N_6114);
nand U8311 (N_8311,N_4832,N_7875);
nor U8312 (N_8312,N_7301,N_6676);
and U8313 (N_8313,N_7418,N_7604);
nor U8314 (N_8314,N_5624,N_6117);
nand U8315 (N_8315,N_4688,N_4509);
nor U8316 (N_8316,N_5357,N_6030);
nand U8317 (N_8317,N_5856,N_6025);
nand U8318 (N_8318,N_4954,N_5650);
and U8319 (N_8319,N_7744,N_5026);
or U8320 (N_8320,N_5647,N_5642);
or U8321 (N_8321,N_4789,N_6557);
nand U8322 (N_8322,N_7594,N_7731);
nor U8323 (N_8323,N_4740,N_4566);
xor U8324 (N_8324,N_4139,N_7566);
or U8325 (N_8325,N_5036,N_5745);
nand U8326 (N_8326,N_5414,N_7337);
or U8327 (N_8327,N_6829,N_4095);
or U8328 (N_8328,N_7457,N_7997);
or U8329 (N_8329,N_7761,N_4062);
or U8330 (N_8330,N_4736,N_7262);
or U8331 (N_8331,N_7182,N_4491);
and U8332 (N_8332,N_5402,N_6455);
and U8333 (N_8333,N_5324,N_6103);
or U8334 (N_8334,N_6086,N_6740);
nand U8335 (N_8335,N_5854,N_4599);
and U8336 (N_8336,N_4774,N_4866);
nand U8337 (N_8337,N_5747,N_4099);
and U8338 (N_8338,N_4081,N_6364);
or U8339 (N_8339,N_5336,N_4915);
nor U8340 (N_8340,N_6817,N_5649);
xnor U8341 (N_8341,N_6629,N_7060);
nor U8342 (N_8342,N_7157,N_5040);
or U8343 (N_8343,N_5048,N_4195);
nor U8344 (N_8344,N_4947,N_4186);
or U8345 (N_8345,N_7094,N_5248);
xor U8346 (N_8346,N_7395,N_6297);
and U8347 (N_8347,N_7167,N_7827);
and U8348 (N_8348,N_4111,N_7176);
and U8349 (N_8349,N_4466,N_5735);
xor U8350 (N_8350,N_4435,N_7417);
or U8351 (N_8351,N_6683,N_4996);
nor U8352 (N_8352,N_5551,N_6420);
and U8353 (N_8353,N_4881,N_7322);
nand U8354 (N_8354,N_7713,N_4517);
nand U8355 (N_8355,N_5974,N_5626);
xor U8356 (N_8356,N_5832,N_4477);
and U8357 (N_8357,N_4883,N_7361);
nor U8358 (N_8358,N_5271,N_5668);
and U8359 (N_8359,N_5557,N_7568);
and U8360 (N_8360,N_6964,N_4170);
xnor U8361 (N_8361,N_5018,N_5097);
or U8362 (N_8362,N_5603,N_6167);
or U8363 (N_8363,N_7107,N_7150);
nor U8364 (N_8364,N_7226,N_4174);
and U8365 (N_8365,N_5759,N_4628);
or U8366 (N_8366,N_7882,N_5352);
nor U8367 (N_8367,N_4233,N_5506);
nand U8368 (N_8368,N_6977,N_7906);
nor U8369 (N_8369,N_4749,N_6207);
nand U8370 (N_8370,N_5087,N_4904);
or U8371 (N_8371,N_6885,N_7825);
or U8372 (N_8372,N_6033,N_6717);
nor U8373 (N_8373,N_6192,N_6891);
or U8374 (N_8374,N_4652,N_6437);
or U8375 (N_8375,N_6750,N_7168);
xor U8376 (N_8376,N_6082,N_4966);
and U8377 (N_8377,N_6008,N_5842);
xor U8378 (N_8378,N_5919,N_6140);
nor U8379 (N_8379,N_4221,N_5462);
and U8380 (N_8380,N_7025,N_7993);
nand U8381 (N_8381,N_6768,N_6263);
or U8382 (N_8382,N_6247,N_4759);
or U8383 (N_8383,N_4582,N_5314);
nor U8384 (N_8384,N_6108,N_4344);
xnor U8385 (N_8385,N_4826,N_7328);
or U8386 (N_8386,N_5309,N_4779);
nor U8387 (N_8387,N_6758,N_6903);
or U8388 (N_8388,N_7873,N_6002);
nand U8389 (N_8389,N_6956,N_6718);
and U8390 (N_8390,N_5806,N_6960);
nand U8391 (N_8391,N_4342,N_7029);
and U8392 (N_8392,N_4575,N_6274);
nand U8393 (N_8393,N_6304,N_6227);
nand U8394 (N_8394,N_5042,N_6136);
and U8395 (N_8395,N_5305,N_6554);
or U8396 (N_8396,N_6824,N_6722);
or U8397 (N_8397,N_5553,N_7441);
xor U8398 (N_8398,N_5878,N_6181);
xnor U8399 (N_8399,N_7493,N_4921);
or U8400 (N_8400,N_4907,N_5519);
nand U8401 (N_8401,N_5894,N_6456);
or U8402 (N_8402,N_4366,N_4260);
and U8403 (N_8403,N_4583,N_7829);
xnor U8404 (N_8404,N_7527,N_6790);
nor U8405 (N_8405,N_7381,N_4230);
nor U8406 (N_8406,N_4555,N_7307);
nand U8407 (N_8407,N_4267,N_7741);
xnor U8408 (N_8408,N_4851,N_6630);
nor U8409 (N_8409,N_5631,N_7973);
nand U8410 (N_8410,N_7085,N_7661);
nand U8411 (N_8411,N_6011,N_7905);
and U8412 (N_8412,N_7763,N_4616);
nand U8413 (N_8413,N_6594,N_7428);
or U8414 (N_8414,N_6375,N_6506);
and U8415 (N_8415,N_5284,N_4691);
or U8416 (N_8416,N_6731,N_6013);
or U8417 (N_8417,N_7312,N_5537);
xor U8418 (N_8418,N_6249,N_4387);
nand U8419 (N_8419,N_4048,N_6116);
and U8420 (N_8420,N_6682,N_6637);
nand U8421 (N_8421,N_4978,N_7726);
nor U8422 (N_8422,N_6861,N_7648);
and U8423 (N_8423,N_5512,N_7816);
nor U8424 (N_8424,N_6426,N_6331);
nand U8425 (N_8425,N_4817,N_6055);
or U8426 (N_8426,N_4984,N_7003);
xnor U8427 (N_8427,N_4923,N_6997);
nor U8428 (N_8428,N_6709,N_7161);
nor U8429 (N_8429,N_4540,N_4316);
nor U8430 (N_8430,N_6590,N_5113);
and U8431 (N_8431,N_7992,N_6673);
and U8432 (N_8432,N_7414,N_6963);
nand U8433 (N_8433,N_4673,N_6688);
and U8434 (N_8434,N_5646,N_4959);
or U8435 (N_8435,N_5670,N_6388);
nand U8436 (N_8436,N_6020,N_7740);
and U8437 (N_8437,N_7177,N_7144);
xor U8438 (N_8438,N_7634,N_6529);
nor U8439 (N_8439,N_7883,N_6808);
or U8440 (N_8440,N_7623,N_7651);
xor U8441 (N_8441,N_7179,N_4087);
or U8442 (N_8442,N_7296,N_6684);
or U8443 (N_8443,N_4503,N_5332);
or U8444 (N_8444,N_6983,N_6762);
or U8445 (N_8445,N_7988,N_4585);
nor U8446 (N_8446,N_4356,N_5700);
nand U8447 (N_8447,N_7786,N_4894);
nor U8448 (N_8448,N_7666,N_6505);
nor U8449 (N_8449,N_7911,N_5550);
xnor U8450 (N_8450,N_5900,N_4823);
nand U8451 (N_8451,N_7704,N_5578);
nor U8452 (N_8452,N_4684,N_7249);
nand U8453 (N_8453,N_5074,N_5073);
nor U8454 (N_8454,N_5844,N_5961);
nand U8455 (N_8455,N_6577,N_7123);
and U8456 (N_8456,N_7450,N_5767);
nand U8457 (N_8457,N_7658,N_7811);
and U8458 (N_8458,N_5100,N_4849);
nor U8459 (N_8459,N_7985,N_6458);
and U8460 (N_8460,N_4977,N_6812);
nor U8461 (N_8461,N_5645,N_7028);
nand U8462 (N_8462,N_7734,N_4023);
and U8463 (N_8463,N_4393,N_7398);
xor U8464 (N_8464,N_5769,N_5667);
nor U8465 (N_8465,N_5193,N_7865);
nand U8466 (N_8466,N_5132,N_5566);
nor U8467 (N_8467,N_4278,N_5711);
nor U8468 (N_8468,N_7617,N_4492);
nand U8469 (N_8469,N_4468,N_4024);
nor U8470 (N_8470,N_5943,N_4295);
nor U8471 (N_8471,N_5913,N_6341);
or U8472 (N_8472,N_5751,N_4258);
and U8473 (N_8473,N_5156,N_4946);
or U8474 (N_8474,N_5103,N_5809);
and U8475 (N_8475,N_4941,N_5993);
and U8476 (N_8476,N_6147,N_4001);
or U8477 (N_8477,N_4047,N_6853);
or U8478 (N_8478,N_6656,N_4998);
nand U8479 (N_8479,N_5515,N_6876);
and U8480 (N_8480,N_6238,N_5277);
and U8481 (N_8481,N_4460,N_7198);
nor U8482 (N_8482,N_6063,N_6786);
nand U8483 (N_8483,N_5730,N_4649);
and U8484 (N_8484,N_5302,N_6672);
nand U8485 (N_8485,N_7615,N_4359);
and U8486 (N_8486,N_5205,N_4775);
nor U8487 (N_8487,N_5850,N_6991);
nor U8488 (N_8488,N_4114,N_6283);
nand U8489 (N_8489,N_6497,N_5580);
nand U8490 (N_8490,N_7534,N_5959);
nand U8491 (N_8491,N_4385,N_5482);
xor U8492 (N_8492,N_7532,N_7649);
xnor U8493 (N_8493,N_7099,N_7197);
xnor U8494 (N_8494,N_4414,N_7915);
xnor U8495 (N_8495,N_4869,N_5863);
and U8496 (N_8496,N_7963,N_7773);
and U8497 (N_8497,N_6368,N_4565);
nand U8498 (N_8498,N_6767,N_5301);
or U8499 (N_8499,N_4548,N_5793);
and U8500 (N_8500,N_6468,N_5740);
or U8501 (N_8501,N_5199,N_5450);
nand U8502 (N_8502,N_5484,N_7386);
and U8503 (N_8503,N_5214,N_7475);
nor U8504 (N_8504,N_5872,N_6990);
nand U8505 (N_8505,N_5167,N_6003);
or U8506 (N_8506,N_4637,N_5687);
xor U8507 (N_8507,N_5823,N_7805);
nand U8508 (N_8508,N_5836,N_7113);
xor U8509 (N_8509,N_4804,N_5859);
and U8510 (N_8510,N_7895,N_6695);
nand U8511 (N_8511,N_5956,N_6865);
nor U8512 (N_8512,N_5908,N_6430);
or U8513 (N_8513,N_6052,N_7042);
and U8514 (N_8514,N_6687,N_5356);
and U8515 (N_8515,N_7931,N_7057);
or U8516 (N_8516,N_5350,N_7472);
nor U8517 (N_8517,N_5216,N_6785);
nor U8518 (N_8518,N_4141,N_6256);
or U8519 (N_8519,N_5788,N_7378);
or U8520 (N_8520,N_5845,N_6308);
and U8521 (N_8521,N_7897,N_7228);
nand U8522 (N_8522,N_5574,N_5365);
nor U8523 (N_8523,N_6254,N_7585);
or U8524 (N_8524,N_6721,N_7435);
or U8525 (N_8525,N_6509,N_5395);
or U8526 (N_8526,N_4828,N_5413);
nand U8527 (N_8527,N_7553,N_6671);
nand U8528 (N_8528,N_6996,N_6409);
and U8529 (N_8529,N_4310,N_5472);
nand U8530 (N_8530,N_6133,N_6464);
xnor U8531 (N_8531,N_6007,N_5883);
nor U8532 (N_8532,N_5604,N_6129);
nor U8533 (N_8533,N_5612,N_7982);
or U8534 (N_8534,N_6995,N_7618);
and U8535 (N_8535,N_4791,N_6438);
or U8536 (N_8536,N_5709,N_6935);
nor U8537 (N_8537,N_7217,N_6899);
nor U8538 (N_8538,N_4445,N_6839);
nor U8539 (N_8539,N_7235,N_5265);
nand U8540 (N_8540,N_6223,N_7664);
nand U8541 (N_8541,N_7551,N_7501);
nor U8542 (N_8542,N_7403,N_4564);
or U8543 (N_8543,N_5072,N_7166);
or U8544 (N_8544,N_6334,N_4550);
xnor U8545 (N_8545,N_4058,N_6265);
and U8546 (N_8546,N_6470,N_5327);
nand U8547 (N_8547,N_6036,N_6627);
and U8548 (N_8548,N_7277,N_7540);
nor U8549 (N_8549,N_7374,N_6874);
xnor U8550 (N_8550,N_5386,N_6987);
or U8551 (N_8551,N_4442,N_4389);
or U8552 (N_8552,N_6854,N_7716);
nor U8553 (N_8553,N_6067,N_7358);
and U8554 (N_8554,N_7336,N_6203);
and U8555 (N_8555,N_5951,N_7141);
and U8556 (N_8556,N_4242,N_7520);
or U8557 (N_8557,N_4951,N_6795);
nand U8558 (N_8558,N_5192,N_7058);
nand U8559 (N_8559,N_4315,N_6994);
and U8560 (N_8560,N_4639,N_4724);
nand U8561 (N_8561,N_4259,N_4171);
nand U8562 (N_8562,N_7923,N_5771);
nor U8563 (N_8563,N_6884,N_7788);
and U8564 (N_8564,N_7023,N_7900);
nor U8565 (N_8565,N_6746,N_6875);
and U8566 (N_8566,N_4119,N_5861);
or U8567 (N_8567,N_4396,N_6632);
or U8568 (N_8568,N_5989,N_6164);
xnor U8569 (N_8569,N_4961,N_4318);
or U8570 (N_8570,N_4379,N_4204);
nor U8571 (N_8571,N_5654,N_5242);
xnor U8572 (N_8572,N_5293,N_6508);
nor U8573 (N_8573,N_6872,N_5764);
nor U8574 (N_8574,N_7066,N_6958);
or U8575 (N_8575,N_7665,N_7346);
nand U8576 (N_8576,N_7241,N_5204);
nor U8577 (N_8577,N_7498,N_7078);
xnor U8578 (N_8578,N_4203,N_4610);
nand U8579 (N_8579,N_7442,N_6317);
nor U8580 (N_8580,N_5534,N_7864);
xor U8581 (N_8581,N_5490,N_5977);
or U8582 (N_8582,N_6385,N_4657);
and U8583 (N_8583,N_5283,N_4937);
xor U8584 (N_8584,N_7563,N_6139);
nand U8585 (N_8585,N_6968,N_6985);
or U8586 (N_8586,N_7950,N_7015);
nor U8587 (N_8587,N_6073,N_7948);
xor U8588 (N_8588,N_5325,N_4199);
or U8589 (N_8589,N_6533,N_6526);
nor U8590 (N_8590,N_4082,N_6165);
nand U8591 (N_8591,N_5452,N_4624);
nand U8592 (N_8592,N_4835,N_7380);
nor U8593 (N_8593,N_4232,N_6060);
and U8594 (N_8594,N_5971,N_7869);
xnor U8595 (N_8595,N_6664,N_5039);
or U8596 (N_8596,N_7353,N_6525);
nand U8597 (N_8597,N_4594,N_4514);
and U8598 (N_8598,N_4080,N_5116);
or U8599 (N_8599,N_5371,N_7285);
and U8600 (N_8600,N_4668,N_7215);
and U8601 (N_8601,N_5427,N_6102);
nor U8602 (N_8602,N_7134,N_7088);
nand U8603 (N_8603,N_6828,N_4026);
nand U8604 (N_8604,N_7027,N_7096);
nor U8605 (N_8605,N_5783,N_4568);
and U8606 (N_8606,N_4733,N_5230);
nand U8607 (N_8607,N_7620,N_6271);
and U8608 (N_8608,N_5019,N_7707);
or U8609 (N_8609,N_7794,N_5569);
or U8610 (N_8610,N_4144,N_4187);
nor U8611 (N_8611,N_7278,N_6942);
nor U8612 (N_8612,N_4709,N_4272);
nor U8613 (N_8613,N_7295,N_5838);
nor U8614 (N_8614,N_4965,N_7887);
nor U8615 (N_8615,N_5732,N_5633);
and U8616 (N_8616,N_4884,N_4824);
or U8617 (N_8617,N_7556,N_6299);
nand U8618 (N_8618,N_5762,N_6988);
and U8619 (N_8619,N_5013,N_7383);
nand U8620 (N_8620,N_5629,N_6491);
nor U8621 (N_8621,N_7304,N_7767);
xnor U8622 (N_8622,N_5354,N_6678);
or U8623 (N_8623,N_6887,N_7127);
nand U8624 (N_8624,N_5211,N_7084);
nand U8625 (N_8625,N_6488,N_4038);
or U8626 (N_8626,N_7964,N_6326);
or U8627 (N_8627,N_4214,N_4788);
or U8628 (N_8628,N_4443,N_6501);
nor U8629 (N_8629,N_4401,N_5677);
nand U8630 (N_8630,N_7684,N_5885);
nand U8631 (N_8631,N_7120,N_7571);
nor U8632 (N_8632,N_5281,N_7530);
and U8633 (N_8633,N_4157,N_7886);
and U8634 (N_8634,N_5443,N_7031);
and U8635 (N_8635,N_7227,N_4075);
and U8636 (N_8636,N_7774,N_4612);
and U8637 (N_8637,N_6926,N_7591);
and U8638 (N_8638,N_5601,N_6973);
and U8639 (N_8639,N_5153,N_5572);
and U8640 (N_8640,N_4635,N_7879);
or U8641 (N_8641,N_4893,N_6635);
nand U8642 (N_8642,N_7517,N_4015);
nand U8643 (N_8643,N_5870,N_5507);
and U8644 (N_8644,N_4900,N_5879);
and U8645 (N_8645,N_6216,N_4224);
nand U8646 (N_8646,N_4208,N_5366);
xnor U8647 (N_8647,N_5810,N_7302);
or U8648 (N_8648,N_6761,N_6573);
or U8649 (N_8649,N_6765,N_4617);
nand U8650 (N_8650,N_5896,N_5118);
nand U8651 (N_8651,N_7691,N_7156);
nand U8652 (N_8652,N_7807,N_7601);
nor U8653 (N_8653,N_6681,N_4350);
nor U8654 (N_8654,N_4899,N_5235);
nor U8655 (N_8655,N_7030,N_7100);
or U8656 (N_8656,N_7835,N_5303);
or U8657 (N_8657,N_6065,N_5232);
nand U8658 (N_8658,N_7017,N_7610);
nand U8659 (N_8659,N_7609,N_6259);
or U8660 (N_8660,N_6564,N_7595);
nor U8661 (N_8661,N_5178,N_6028);
xor U8662 (N_8662,N_6107,N_6517);
nand U8663 (N_8663,N_4341,N_5628);
and U8664 (N_8664,N_7893,N_6933);
or U8665 (N_8665,N_6834,N_4059);
xnor U8666 (N_8666,N_4013,N_5004);
nor U8667 (N_8667,N_7852,N_5275);
nand U8668 (N_8668,N_6261,N_4345);
nor U8669 (N_8669,N_5682,N_5270);
or U8670 (N_8670,N_5496,N_7343);
nand U8671 (N_8671,N_6109,N_4005);
nand U8672 (N_8672,N_5614,N_7779);
nor U8673 (N_8673,N_5384,N_4142);
nand U8674 (N_8674,N_6846,N_4268);
and U8675 (N_8675,N_6361,N_7070);
or U8676 (N_8676,N_4179,N_5716);
or U8677 (N_8677,N_4949,N_6383);
nor U8678 (N_8678,N_5163,N_4358);
nor U8679 (N_8679,N_6555,N_6321);
nand U8680 (N_8680,N_4536,N_5611);
xor U8681 (N_8681,N_6749,N_4061);
xor U8682 (N_8682,N_7429,N_7298);
and U8683 (N_8683,N_5585,N_7470);
nor U8684 (N_8684,N_5938,N_6536);
nor U8685 (N_8685,N_4177,N_7091);
or U8686 (N_8686,N_6362,N_4846);
nand U8687 (N_8687,N_7290,N_5934);
nand U8688 (N_8688,N_6301,N_5698);
or U8689 (N_8689,N_6217,N_6125);
xor U8690 (N_8690,N_7432,N_4761);
nand U8691 (N_8691,N_6574,N_4615);
nand U8692 (N_8692,N_4773,N_4611);
nand U8693 (N_8693,N_4842,N_4819);
or U8694 (N_8694,N_6074,N_5456);
or U8695 (N_8695,N_6371,N_6625);
or U8696 (N_8696,N_4642,N_4083);
or U8697 (N_8697,N_6607,N_6088);
xor U8698 (N_8698,N_5697,N_5536);
nor U8699 (N_8699,N_6551,N_5596);
and U8700 (N_8700,N_6993,N_7466);
and U8701 (N_8701,N_6405,N_6920);
and U8702 (N_8702,N_5756,N_5573);
or U8703 (N_8703,N_5505,N_7801);
or U8704 (N_8704,N_6293,N_6787);
nor U8705 (N_8705,N_4902,N_6931);
nand U8706 (N_8706,N_5015,N_5535);
xnor U8707 (N_8707,N_5805,N_5115);
or U8708 (N_8708,N_6592,N_4584);
or U8709 (N_8709,N_4400,N_5822);
xnor U8710 (N_8710,N_6855,N_6231);
nor U8711 (N_8711,N_7483,N_6415);
or U8712 (N_8712,N_7885,N_4559);
nor U8713 (N_8713,N_6399,N_5912);
or U8714 (N_8714,N_5720,N_4682);
and U8715 (N_8715,N_4158,N_6744);
and U8716 (N_8716,N_7281,N_5690);
xnor U8717 (N_8717,N_5149,N_7519);
xor U8718 (N_8718,N_4288,N_4429);
and U8719 (N_8719,N_7394,N_7681);
or U8720 (N_8720,N_5396,N_4754);
or U8721 (N_8721,N_7818,N_5606);
or U8722 (N_8722,N_4173,N_7196);
nand U8723 (N_8723,N_6534,N_6119);
nand U8724 (N_8724,N_4457,N_6984);
or U8725 (N_8725,N_5387,N_7377);
or U8726 (N_8726,N_4306,N_5186);
nor U8727 (N_8727,N_7980,N_5797);
nand U8728 (N_8728,N_4552,N_6300);
nor U8729 (N_8729,N_6402,N_7663);
nor U8730 (N_8730,N_4397,N_6431);
and U8731 (N_8731,N_5731,N_5742);
or U8732 (N_8732,N_7087,N_7682);
nand U8733 (N_8733,N_4827,N_6302);
or U8734 (N_8734,N_6559,N_6270);
nor U8735 (N_8735,N_4044,N_6739);
and U8736 (N_8736,N_4390,N_5882);
and U8737 (N_8737,N_5674,N_4728);
or U8738 (N_8738,N_6292,N_4403);
and U8739 (N_8739,N_4108,N_7308);
nand U8740 (N_8740,N_6650,N_6474);
nor U8741 (N_8741,N_4454,N_6706);
and U8742 (N_8742,N_6809,N_6538);
xor U8743 (N_8743,N_6257,N_5096);
and U8744 (N_8744,N_7211,N_4940);
or U8745 (N_8745,N_5045,N_6240);
nand U8746 (N_8746,N_5895,N_6613);
and U8747 (N_8747,N_7531,N_5007);
or U8748 (N_8748,N_4631,N_7611);
nand U8749 (N_8749,N_4383,N_6826);
or U8750 (N_8750,N_5022,N_7272);
and U8751 (N_8751,N_4347,N_6154);
and U8752 (N_8752,N_6134,N_4440);
nor U8753 (N_8753,N_4834,N_4282);
nand U8754 (N_8754,N_4068,N_7573);
nor U8755 (N_8755,N_4322,N_5821);
nor U8756 (N_8756,N_4971,N_7696);
nor U8757 (N_8757,N_7650,N_6460);
or U8758 (N_8758,N_6005,N_4402);
or U8759 (N_8759,N_5408,N_4329);
and U8760 (N_8760,N_4314,N_5378);
nand U8761 (N_8761,N_6580,N_7116);
nor U8762 (N_8762,N_4348,N_5916);
and U8763 (N_8763,N_6168,N_5542);
nand U8764 (N_8764,N_6626,N_6215);
nor U8765 (N_8765,N_6498,N_7291);
nor U8766 (N_8766,N_4346,N_7673);
or U8767 (N_8767,N_7978,N_4455);
xnor U8768 (N_8768,N_5552,N_7702);
nand U8769 (N_8769,N_7449,N_6602);
and U8770 (N_8770,N_7400,N_4580);
nand U8771 (N_8771,N_4560,N_6911);
or U8772 (N_8772,N_7348,N_7005);
nand U8773 (N_8773,N_6946,N_7715);
or U8774 (N_8774,N_4264,N_5445);
nand U8775 (N_8775,N_7929,N_7558);
or U8776 (N_8776,N_7956,N_5813);
nand U8777 (N_8777,N_4981,N_6085);
nor U8778 (N_8778,N_4822,N_5533);
and U8779 (N_8779,N_6622,N_4569);
nand U8780 (N_8780,N_6155,N_6273);
nand U8781 (N_8781,N_7233,N_7054);
nand U8782 (N_8782,N_5902,N_4879);
or U8783 (N_8783,N_4012,N_6230);
or U8784 (N_8784,N_5928,N_6959);
or U8785 (N_8785,N_4859,N_7180);
or U8786 (N_8786,N_4134,N_5442);
or U8787 (N_8787,N_6079,N_6584);
xor U8788 (N_8788,N_7209,N_7315);
nand U8789 (N_8789,N_7175,N_4931);
xnor U8790 (N_8790,N_6183,N_6348);
nor U8791 (N_8791,N_5245,N_4707);
nor U8792 (N_8792,N_5044,N_6900);
nand U8793 (N_8793,N_7284,N_4714);
nor U8794 (N_8794,N_6204,N_5520);
nand U8795 (N_8795,N_6612,N_7152);
nand U8796 (N_8796,N_5532,N_7575);
nand U8797 (N_8797,N_4507,N_4217);
or U8798 (N_8798,N_7213,N_4839);
or U8799 (N_8799,N_4422,N_7853);
nor U8800 (N_8800,N_7056,N_6716);
nand U8801 (N_8801,N_4739,N_5197);
nand U8802 (N_8802,N_5075,N_5014);
xnor U8803 (N_8803,N_5229,N_5841);
nor U8804 (N_8804,N_4241,N_4302);
nor U8805 (N_8805,N_4256,N_4106);
xnor U8806 (N_8806,N_4496,N_7544);
nand U8807 (N_8807,N_4499,N_6725);
and U8808 (N_8808,N_5394,N_5554);
nand U8809 (N_8809,N_4388,N_6056);
or U8810 (N_8810,N_6500,N_6582);
nand U8811 (N_8811,N_4837,N_6001);
or U8812 (N_8812,N_5803,N_5607);
and U8813 (N_8813,N_5867,N_4486);
nand U8814 (N_8814,N_4645,N_7918);
or U8815 (N_8815,N_7654,N_7724);
nor U8816 (N_8816,N_4250,N_5374);
and U8817 (N_8817,N_5789,N_6544);
or U8818 (N_8818,N_6608,N_7254);
nor U8819 (N_8819,N_7889,N_4613);
or U8820 (N_8820,N_4577,N_4122);
or U8821 (N_8821,N_4183,N_7717);
nor U8822 (N_8822,N_6191,N_6764);
or U8823 (N_8823,N_7014,N_5795);
and U8824 (N_8824,N_4760,N_4793);
nor U8825 (N_8825,N_4727,N_5960);
and U8826 (N_8826,N_4189,N_4045);
nand U8827 (N_8827,N_5109,N_7739);
and U8828 (N_8828,N_6218,N_7638);
nand U8829 (N_8829,N_4587,N_5501);
and U8830 (N_8830,N_4299,N_6176);
and U8831 (N_8831,N_6232,N_6735);
and U8832 (N_8832,N_7259,N_7232);
nor U8833 (N_8833,N_4084,N_7491);
or U8834 (N_8834,N_7936,N_5021);
and U8835 (N_8835,N_5148,N_4159);
and U8836 (N_8836,N_4017,N_4010);
nor U8837 (N_8837,N_6609,N_5779);
xor U8838 (N_8838,N_6837,N_7722);
or U8839 (N_8839,N_5084,N_4796);
and U8840 (N_8840,N_6708,N_4482);
and U8841 (N_8841,N_4225,N_7489);
nand U8842 (N_8842,N_7939,N_5262);
nand U8843 (N_8843,N_4475,N_6969);
and U8844 (N_8844,N_5558,N_6413);
and U8845 (N_8845,N_6763,N_7373);
or U8846 (N_8846,N_7815,N_7347);
nand U8847 (N_8847,N_7721,N_6344);
nor U8848 (N_8848,N_5266,N_6710);
nand U8849 (N_8849,N_7946,N_7699);
or U8850 (N_8850,N_4967,N_5831);
nor U8851 (N_8851,N_5639,N_4236);
xor U8852 (N_8852,N_4105,N_7055);
xnor U8853 (N_8853,N_5661,N_7101);
nor U8854 (N_8854,N_7181,N_6374);
nor U8855 (N_8855,N_6145,N_4970);
nand U8856 (N_8856,N_5733,N_5376);
and U8857 (N_8857,N_7872,N_5397);
nand U8858 (N_8858,N_6188,N_7705);
nand U8859 (N_8859,N_4436,N_5985);
nand U8860 (N_8860,N_6645,N_7131);
nand U8861 (N_8861,N_5328,N_6856);
or U8862 (N_8862,N_5923,N_7145);
nand U8863 (N_8863,N_7357,N_5367);
nor U8864 (N_8864,N_7468,N_6668);
nand U8865 (N_8865,N_6295,N_7218);
nand U8866 (N_8866,N_6211,N_6866);
and U8867 (N_8867,N_7185,N_7567);
and U8868 (N_8868,N_7521,N_7975);
and U8869 (N_8869,N_7524,N_4309);
and U8870 (N_8870,N_6567,N_5479);
and U8871 (N_8871,N_6700,N_4129);
and U8872 (N_8872,N_6404,N_6075);
and U8873 (N_8873,N_6260,N_6045);
nand U8874 (N_8874,N_5342,N_5942);
nor U8875 (N_8875,N_7849,N_5840);
or U8876 (N_8876,N_6472,N_5485);
nand U8877 (N_8877,N_7820,N_5085);
xnor U8878 (N_8878,N_7795,N_6290);
nor U8879 (N_8879,N_5282,N_5033);
or U8880 (N_8880,N_5320,N_4513);
or U8881 (N_8881,N_5154,N_4462);
and U8882 (N_8882,N_4632,N_7471);
nor U8883 (N_8883,N_5594,N_6141);
and U8884 (N_8884,N_5362,N_5173);
or U8885 (N_8885,N_6811,N_6583);
or U8886 (N_8886,N_7619,N_4110);
and U8887 (N_8887,N_6061,N_6160);
and U8888 (N_8888,N_4176,N_5406);
and U8889 (N_8889,N_7355,N_4231);
or U8890 (N_8890,N_4502,N_5299);
or U8891 (N_8891,N_7733,N_7436);
and U8892 (N_8892,N_6436,N_4901);
or U8893 (N_8893,N_5728,N_6954);
nor U8894 (N_8894,N_4604,N_6904);
and U8895 (N_8895,N_6394,N_5869);
or U8896 (N_8896,N_4420,N_6118);
nor U8897 (N_8897,N_5058,N_7996);
nand U8898 (N_8898,N_4184,N_4678);
nand U8899 (N_8899,N_5724,N_4234);
or U8900 (N_8900,N_6704,N_5068);
and U8901 (N_8901,N_4916,N_5446);
and U8902 (N_8902,N_5112,N_6229);
and U8903 (N_8903,N_6442,N_5240);
nor U8904 (N_8904,N_5544,N_4618);
and U8905 (N_8905,N_6105,N_7095);
nor U8906 (N_8906,N_7495,N_4766);
and U8907 (N_8907,N_4464,N_6796);
xor U8908 (N_8908,N_4524,N_4776);
nand U8909 (N_8909,N_6901,N_7581);
and U8910 (N_8910,N_5179,N_6345);
nand U8911 (N_8911,N_7679,N_6511);
nor U8912 (N_8912,N_7560,N_4497);
or U8913 (N_8913,N_5621,N_4228);
and U8914 (N_8914,N_6357,N_7612);
and U8915 (N_8915,N_6315,N_6342);
xor U8916 (N_8916,N_5164,N_6078);
nor U8917 (N_8917,N_6111,N_4731);
nand U8918 (N_8918,N_7995,N_4528);
nor U8919 (N_8919,N_4681,N_6552);
nor U8920 (N_8920,N_6169,N_5139);
or U8921 (N_8921,N_7041,N_7224);
nor U8922 (N_8922,N_4320,N_7469);
or U8923 (N_8923,N_4438,N_5696);
or U8924 (N_8924,N_5752,N_4249);
and U8925 (N_8925,N_7102,N_5217);
nand U8926 (N_8926,N_6714,N_7760);
or U8927 (N_8927,N_4248,N_4533);
nor U8928 (N_8928,N_6628,N_5136);
and U8929 (N_8929,N_6089,N_4541);
and U8930 (N_8930,N_6759,N_7413);
nand U8931 (N_8931,N_6220,N_5431);
nand U8932 (N_8932,N_7635,N_6966);
or U8933 (N_8933,N_6091,N_4423);
and U8934 (N_8934,N_5653,N_6836);
xnor U8935 (N_8935,N_5591,N_5455);
and U8936 (N_8936,N_4539,N_7356);
and U8937 (N_8937,N_7874,N_5471);
nand U8938 (N_8938,N_6944,N_5510);
and U8939 (N_8939,N_7130,N_4734);
and U8940 (N_8940,N_6906,N_5129);
nand U8941 (N_8941,N_7799,N_5331);
nor U8942 (N_8942,N_6152,N_4983);
and U8943 (N_8943,N_7089,N_5804);
nand U8944 (N_8944,N_7111,N_7426);
xor U8945 (N_8945,N_5458,N_7824);
and U8946 (N_8946,N_5685,N_7940);
and U8947 (N_8947,N_4629,N_6462);
nor U8948 (N_8948,N_7437,N_5409);
and U8949 (N_8949,N_7022,N_7756);
nand U8950 (N_8950,N_6266,N_5279);
or U8951 (N_8951,N_5105,N_6296);
nand U8952 (N_8952,N_7871,N_6276);
nor U8953 (N_8953,N_6499,N_5119);
nand U8954 (N_8954,N_7582,N_6049);
and U8955 (N_8955,N_4805,N_6614);
nor U8956 (N_8956,N_4404,N_7957);
nor U8957 (N_8957,N_4270,N_5734);
xnor U8958 (N_8958,N_6182,N_4406);
or U8959 (N_8959,N_4781,N_7770);
or U8960 (N_8960,N_7399,N_6967);
and U8961 (N_8961,N_7597,N_5255);
nor U8962 (N_8962,N_4121,N_4078);
and U8963 (N_8963,N_6101,N_7792);
nor U8964 (N_8964,N_6449,N_7892);
nor U8965 (N_8965,N_4266,N_5024);
xor U8966 (N_8966,N_4399,N_5772);
xnor U8967 (N_8967,N_4777,N_7079);
or U8968 (N_8968,N_6034,N_7629);
nand U8969 (N_8969,N_6312,N_7237);
or U8970 (N_8970,N_7103,N_5448);
nand U8971 (N_8971,N_5610,N_6543);
nand U8972 (N_8972,N_4530,N_7550);
and U8973 (N_8973,N_7271,N_5061);
and U8974 (N_8974,N_6644,N_4922);
or U8975 (N_8975,N_4680,N_7628);
nand U8976 (N_8976,N_7943,N_5794);
or U8977 (N_8977,N_5691,N_6081);
nor U8978 (N_8978,N_4857,N_6728);
nor U8979 (N_8979,N_5658,N_7169);
nand U8980 (N_8980,N_4461,N_6489);
or U8981 (N_8981,N_5076,N_6354);
and U8982 (N_8982,N_6252,N_4867);
nand U8983 (N_8983,N_7942,N_7032);
xor U8984 (N_8984,N_6621,N_6978);
nor U8985 (N_8985,N_5798,N_5111);
or U8986 (N_8986,N_6772,N_5528);
nand U8987 (N_8987,N_5791,N_7776);
nor U8988 (N_8988,N_6843,N_4473);
xnor U8989 (N_8989,N_6044,N_4803);
nor U8990 (N_8990,N_7542,N_5041);
and U8991 (N_8991,N_4747,N_5056);
nor U8992 (N_8992,N_6913,N_5714);
and U8993 (N_8993,N_7240,N_5032);
nor U8994 (N_8994,N_5839,N_4146);
or U8995 (N_8995,N_6367,N_7034);
nor U8996 (N_8996,N_7049,N_5598);
and U8997 (N_8997,N_7407,N_5684);
nand U8998 (N_8998,N_4033,N_7934);
and U8999 (N_8999,N_5874,N_4597);
and U9000 (N_9000,N_4696,N_6976);
nand U9001 (N_9001,N_4693,N_4138);
or U9002 (N_9002,N_7214,N_4419);
nor U9003 (N_9003,N_7006,N_6027);
or U9004 (N_9004,N_6050,N_7194);
or U9005 (N_9005,N_4718,N_4625);
or U9006 (N_9006,N_7846,N_7945);
nor U9007 (N_9007,N_7048,N_6883);
and U9008 (N_9008,N_7683,N_5207);
xor U9009 (N_9009,N_6323,N_5982);
nor U9010 (N_9010,N_5525,N_5280);
xor U9011 (N_9011,N_4778,N_4052);
nor U9012 (N_9012,N_6318,N_4218);
nand U9013 (N_9013,N_7912,N_4765);
nor U9014 (N_9014,N_7506,N_7999);
and U9015 (N_9015,N_5922,N_7845);
nor U9016 (N_9016,N_4521,N_6860);
and U9017 (N_9017,N_7329,N_5348);
or U9018 (N_9018,N_5313,N_4744);
nand U9019 (N_9019,N_5393,N_6048);
or U9020 (N_9020,N_7010,N_6146);
or U9021 (N_9021,N_6532,N_6537);
or U9022 (N_9022,N_6847,N_4863);
or U9023 (N_9023,N_7970,N_7011);
xor U9024 (N_9024,N_5932,N_5035);
or U9025 (N_9025,N_4992,N_4813);
nor U9026 (N_9026,N_4133,N_4726);
or U9027 (N_9027,N_7230,N_6427);
nor U9028 (N_9028,N_4936,N_5141);
nor U9029 (N_9029,N_6094,N_6006);
and U9030 (N_9030,N_7891,N_4113);
and U9031 (N_9031,N_7708,N_4175);
nand U9032 (N_9032,N_4948,N_7245);
nand U9033 (N_9033,N_7557,N_7802);
or U9034 (N_9034,N_4117,N_4913);
nand U9035 (N_9035,N_5051,N_7093);
or U9036 (N_9036,N_7725,N_7053);
or U9037 (N_9037,N_4928,N_5345);
nand U9038 (N_9038,N_5464,N_7888);
and U9039 (N_9039,N_4831,N_4903);
or U9040 (N_9040,N_5377,N_7430);
nand U9041 (N_9041,N_7117,N_6406);
xor U9042 (N_9042,N_5754,N_6112);
nor U9043 (N_9043,N_7019,N_4490);
nand U9044 (N_9044,N_6369,N_4534);
nor U9045 (N_9045,N_7984,N_6235);
or U9046 (N_9046,N_7782,N_4525);
and U9047 (N_9047,N_5412,N_5643);
and U9048 (N_9048,N_6000,N_6397);
nor U9049 (N_9049,N_4333,N_6766);
and U9050 (N_9050,N_7423,N_7959);
nand U9051 (N_9051,N_7881,N_4072);
nand U9052 (N_9052,N_7884,N_7204);
and U9053 (N_9053,N_5483,N_4226);
xor U9054 (N_9054,N_5518,N_5128);
or U9055 (N_9055,N_5273,N_6279);
nor U9056 (N_9056,N_7485,N_4421);
or U9057 (N_9057,N_6510,N_5092);
or U9058 (N_9058,N_4785,N_5251);
nor U9059 (N_9059,N_7486,N_6774);
nor U9060 (N_9060,N_5010,N_4880);
nand U9061 (N_9061,N_7497,N_7222);
and U9062 (N_9062,N_5595,N_7406);
or U9063 (N_9063,N_7636,N_7769);
and U9064 (N_9064,N_4073,N_4279);
or U9065 (N_9065,N_6454,N_6138);
or U9066 (N_9066,N_4974,N_4969);
nor U9067 (N_9067,N_6713,N_4051);
nor U9068 (N_9068,N_4285,N_6351);
nor U9069 (N_9069,N_4162,N_6411);
nand U9070 (N_9070,N_7735,N_5088);
and U9071 (N_9071,N_7340,N_5410);
or U9072 (N_9072,N_4769,N_5561);
nor U9073 (N_9073,N_4271,N_4938);
and U9074 (N_9074,N_7480,N_4829);
nand U9075 (N_9075,N_5920,N_7135);
nand U9076 (N_9076,N_6486,N_6938);
xor U9077 (N_9077,N_4060,N_7273);
or U9078 (N_9078,N_7928,N_6376);
or U9079 (N_9079,N_4097,N_5722);
xnor U9080 (N_9080,N_4064,N_5503);
and U9081 (N_9081,N_4886,N_6435);
or U9082 (N_9082,N_5295,N_6588);
nand U9083 (N_9083,N_6949,N_5868);
nor U9084 (N_9084,N_6802,N_6358);
or U9085 (N_9085,N_7481,N_6912);
nand U9086 (N_9086,N_4153,N_5799);
nand U9087 (N_9087,N_6962,N_6851);
xor U9088 (N_9088,N_7391,N_5030);
or U9089 (N_9089,N_4927,N_5433);
and U9090 (N_9090,N_5474,N_7798);
and U9091 (N_9091,N_4544,N_4197);
nor U9092 (N_9092,N_4427,N_5460);
or U9093 (N_9093,N_5166,N_5368);
or U9094 (N_9094,N_5766,N_4850);
nor U9095 (N_9095,N_4522,N_7330);
nand U9096 (N_9096,N_6264,N_4092);
nand U9097 (N_9097,N_7286,N_7602);
or U9098 (N_9098,N_4891,N_5253);
xor U9099 (N_9099,N_4806,N_6403);
and U9100 (N_9100,N_5375,N_5319);
xnor U9101 (N_9101,N_7979,N_4958);
or U9102 (N_9102,N_5593,N_7459);
nor U9103 (N_9103,N_7372,N_7749);
and U9104 (N_9104,N_4200,N_7541);
and U9105 (N_9105,N_4692,N_5672);
or U9106 (N_9106,N_5623,N_7154);
nand U9107 (N_9107,N_6047,N_7743);
xnor U9108 (N_9108,N_5886,N_4160);
nor U9109 (N_9109,N_5162,N_7689);
nor U9110 (N_9110,N_6952,N_7641);
nor U9111 (N_9111,N_5308,N_7719);
or U9112 (N_9112,N_7163,N_6303);
nor U9113 (N_9113,N_6953,N_5135);
nor U9114 (N_9114,N_4296,N_5926);
xor U9115 (N_9115,N_4885,N_7878);
nand U9116 (N_9116,N_5310,N_6778);
or U9117 (N_9117,N_4008,N_6267);
nor U9118 (N_9118,N_4518,N_7510);
nand U9119 (N_9119,N_6546,N_7518);
nor U9120 (N_9120,N_4382,N_5903);
xnor U9121 (N_9121,N_5787,N_5563);
or U9122 (N_9122,N_7657,N_6482);
nand U9123 (N_9123,N_7004,N_4066);
or U9124 (N_9124,N_7149,N_5005);
and U9125 (N_9125,N_6869,N_7397);
or U9126 (N_9126,N_6504,N_4161);
and U9127 (N_9127,N_6616,N_7826);
or U9128 (N_9128,N_4551,N_6310);
nand U9129 (N_9129,N_7174,N_5818);
nor U9130 (N_9130,N_7633,N_4750);
and U9131 (N_9131,N_7434,N_7098);
nand U9132 (N_9132,N_4795,N_4968);
and U9133 (N_9133,N_5715,N_7606);
nor U9134 (N_9134,N_6793,N_6723);
nand U9135 (N_9135,N_4243,N_6359);
nor U9136 (N_9136,N_5706,N_7953);
nor U9137 (N_9137,N_7775,N_5898);
xor U9138 (N_9138,N_5917,N_4515);
nor U9139 (N_9139,N_5616,N_7090);
or U9140 (N_9140,N_4800,N_6040);
xnor U9141 (N_9141,N_4408,N_4166);
nor U9142 (N_9142,N_7947,N_4493);
xnor U9143 (N_9143,N_4810,N_6066);
nand U9144 (N_9144,N_6269,N_5304);
or U9145 (N_9145,N_6919,N_5337);
and U9146 (N_9146,N_4247,N_7363);
xor U9147 (N_9147,N_5749,N_4205);
and U9148 (N_9148,N_5498,N_7855);
and U9149 (N_9149,N_4667,N_7630);
nand U9150 (N_9150,N_6540,N_4855);
nand U9151 (N_9151,N_5244,N_4447);
nor U9152 (N_9152,N_7236,N_6769);
nor U9153 (N_9153,N_4312,N_5849);
nor U9154 (N_9154,N_6309,N_7967);
nor U9155 (N_9155,N_6142,N_4723);
or U9156 (N_9156,N_5415,N_4988);
and U9157 (N_9157,N_5218,N_5702);
or U9158 (N_9158,N_5775,N_4504);
and U9159 (N_9159,N_7445,N_7718);
or U9160 (N_9160,N_6226,N_7300);
nor U9161 (N_9161,N_4756,N_7043);
and U9162 (N_9162,N_6820,N_4215);
and U9163 (N_9163,N_6490,N_5449);
nand U9164 (N_9164,N_7496,N_4508);
and U9165 (N_9165,N_4418,N_5065);
and U9166 (N_9166,N_5527,N_7574);
xnor U9167 (N_9167,N_7248,N_7239);
or U9168 (N_9168,N_5228,N_6788);
xnor U9169 (N_9169,N_4069,N_5108);
and U9170 (N_9170,N_5892,N_5487);
or U9171 (N_9171,N_4889,N_4656);
nand U9172 (N_9172,N_7861,N_4131);
nor U9173 (N_9173,N_4182,N_5082);
nor U9174 (N_9174,N_7452,N_4767);
nor U9175 (N_9175,N_6667,N_7781);
and U9176 (N_9176,N_4287,N_5272);
nor U9177 (N_9177,N_7608,N_6518);
nand U9178 (N_9178,N_4194,N_4596);
nor U9179 (N_9179,N_4269,N_7907);
and U9180 (N_9180,N_6305,N_6446);
nor U9181 (N_9181,N_5543,N_7171);
xnor U9182 (N_9182,N_7727,N_7001);
nor U9183 (N_9183,N_5718,N_5770);
xor U9184 (N_9184,N_7754,N_4762);
and U9185 (N_9185,N_4689,N_7863);
or U9186 (N_9186,N_7583,N_4672);
nand U9187 (N_9187,N_7909,N_7814);
and U9188 (N_9188,N_6387,N_4453);
or U9189 (N_9189,N_7838,N_6471);
and U9190 (N_9190,N_6732,N_7220);
or U9191 (N_9191,N_6880,N_7670);
and U9192 (N_9192,N_7539,N_7350);
and U9193 (N_9193,N_4698,N_6807);
nor U9194 (N_9194,N_4809,N_5358);
and U9195 (N_9195,N_5517,N_5034);
and U9196 (N_9196,N_5080,N_6565);
nor U9197 (N_9197,N_4840,N_6620);
nor U9198 (N_9198,N_4476,N_5833);
nand U9199 (N_9199,N_5736,N_6035);
nor U9200 (N_9200,N_6193,N_5978);
and U9201 (N_9201,N_5758,N_6019);
nand U9202 (N_9202,N_7146,N_4784);
nand U9203 (N_9203,N_4895,N_5853);
and U9204 (N_9204,N_6600,N_4223);
nand U9205 (N_9205,N_6476,N_4216);
and U9206 (N_9206,N_7772,N_6393);
or U9207 (N_9207,N_4002,N_7201);
and U9208 (N_9208,N_7837,N_7371);
nand U9209 (N_9209,N_4451,N_5784);
nand U9210 (N_9210,N_4963,N_6898);
nor U9211 (N_9211,N_7026,N_6566);
nand U9212 (N_9212,N_5757,N_7463);
nand U9213 (N_9213,N_7122,N_5881);
nor U9214 (N_9214,N_4003,N_6291);
or U9215 (N_9215,N_6120,N_5142);
nand U9216 (N_9216,N_7836,N_7009);
and U9217 (N_9217,N_5953,N_5028);
or U9218 (N_9218,N_5160,N_7522);
nor U9219 (N_9219,N_4735,N_4100);
nand U9220 (N_9220,N_4812,N_7075);
nand U9221 (N_9221,N_4014,N_4664);
nor U9222 (N_9222,N_5382,N_4042);
nand U9223 (N_9223,N_5288,N_6558);
nand U9224 (N_9224,N_7274,N_5619);
nand U9225 (N_9225,N_6477,N_6010);
nand U9226 (N_9226,N_7925,N_7841);
or U9227 (N_9227,N_6576,N_5555);
or U9228 (N_9228,N_4953,N_4722);
and U9229 (N_9229,N_6083,N_4089);
nand U9230 (N_9230,N_6023,N_7421);
and U9231 (N_9231,N_5876,N_7791);
and U9232 (N_9232,N_7128,N_7453);
and U9233 (N_9233,N_4039,N_7712);
nand U9234 (N_9234,N_5509,N_5260);
nor U9235 (N_9235,N_4841,N_7570);
nand U9236 (N_9236,N_4875,N_6126);
xnor U9237 (N_9237,N_6715,N_7830);
nand U9238 (N_9238,N_4771,N_6153);
or U9239 (N_9239,N_6852,N_6275);
or U9240 (N_9240,N_5290,N_7316);
nand U9241 (N_9241,N_5617,N_4820);
nand U9242 (N_9242,N_7118,N_7968);
xor U9243 (N_9243,N_5523,N_5023);
xnor U9244 (N_9244,N_4426,N_6742);
or U9245 (N_9245,N_7616,N_7809);
and U9246 (N_9246,N_4136,N_5182);
xnor U9247 (N_9247,N_7800,N_6748);
xnor U9248 (N_9248,N_7045,N_7543);
or U9249 (N_9249,N_5289,N_5746);
or U9250 (N_9250,N_5605,N_4034);
and U9251 (N_9251,N_6784,N_4906);
nand U9252 (N_9252,N_6698,N_6311);
nand U9253 (N_9253,N_7420,N_4398);
nand U9254 (N_9254,N_5095,N_7823);
or U9255 (N_9255,N_4662,N_7370);
nor U9256 (N_9256,N_5755,N_7904);
nor U9257 (N_9257,N_6610,N_5516);
nand U9258 (N_9258,N_6239,N_6289);
nor U9259 (N_9259,N_4211,N_4107);
nor U9260 (N_9260,N_7859,N_5344);
nand U9261 (N_9261,N_4209,N_4130);
and U9262 (N_9262,N_5632,N_5996);
or U9263 (N_9263,N_7972,N_7276);
nand U9264 (N_9264,N_5530,N_5846);
and U9265 (N_9265,N_5159,N_6989);
and U9266 (N_9266,N_4782,N_5914);
or U9267 (N_9267,N_5057,N_4685);
nand U9268 (N_9268,N_4960,N_6479);
or U9269 (N_9269,N_7762,N_7751);
nor U9270 (N_9270,N_6757,N_7857);
xnor U9271 (N_9271,N_7926,N_6480);
and U9272 (N_9272,N_5500,N_4088);
or U9273 (N_9273,N_6439,N_4621);
nor U9274 (N_9274,N_4864,N_6422);
nor U9275 (N_9275,N_5692,N_4407);
and U9276 (N_9276,N_5363,N_6492);
and U9277 (N_9277,N_6281,N_6699);
xor U9278 (N_9278,N_6842,N_4821);
and U9279 (N_9279,N_7746,N_6857);
or U9280 (N_9280,N_6752,N_5562);
nor U9281 (N_9281,N_5589,N_4145);
nor U9282 (N_9282,N_4070,N_7188);
xnor U9283 (N_9283,N_6288,N_6467);
xor U9284 (N_9284,N_5488,N_4343);
and U9285 (N_9285,N_6171,N_4364);
nor U9286 (N_9286,N_5435,N_7477);
nand U9287 (N_9287,N_7083,N_5999);
or U9288 (N_9288,N_5246,N_5404);
nor U9289 (N_9289,N_6199,N_4619);
or U9290 (N_9290,N_4874,N_5373);
and U9291 (N_9291,N_4590,N_5665);
nor U9292 (N_9292,N_4768,N_6377);
nor U9293 (N_9293,N_4163,N_4036);
or U9294 (N_9294,N_6070,N_5138);
and U9295 (N_9295,N_6905,N_6212);
or U9296 (N_9296,N_5322,N_6818);
or U9297 (N_9297,N_5494,N_5949);
or U9298 (N_9298,N_6879,N_4446);
nor U9299 (N_9299,N_4465,N_4729);
nand U9300 (N_9300,N_6286,N_7500);
and U9301 (N_9301,N_4381,N_4606);
nor U9302 (N_9302,N_7139,N_6797);
or U9303 (N_9303,N_4543,N_4298);
and U9304 (N_9304,N_4360,N_7287);
nand U9305 (N_9305,N_6282,N_5379);
nand U9306 (N_9306,N_7847,N_7265);
nor U9307 (N_9307,N_6658,N_7624);
xor U9308 (N_9308,N_4277,N_5825);
and U9309 (N_9309,N_5568,N_4955);
nor U9310 (N_9310,N_6320,N_5340);
and U9311 (N_9311,N_7505,N_4836);
and U9312 (N_9312,N_7068,N_6280);
and U9313 (N_9313,N_7335,N_6225);
and U9314 (N_9314,N_4391,N_4395);
or U9315 (N_9315,N_5315,N_7808);
and U9316 (N_9316,N_5905,N_7580);
nand U9317 (N_9317,N_6058,N_5117);
nor U9318 (N_9318,N_4634,N_6568);
and U9319 (N_9319,N_7728,N_7590);
or U9320 (N_9320,N_6690,N_7199);
and U9321 (N_9321,N_5391,N_4697);
and U9322 (N_9322,N_4660,N_5401);
or U9323 (N_9323,N_5183,N_7921);
nor U9324 (N_9324,N_5708,N_7678);
xnor U9325 (N_9325,N_4463,N_7018);
and U9326 (N_9326,N_5773,N_7106);
nand U9327 (N_9327,N_7320,N_5190);
nor U9328 (N_9328,N_5238,N_7832);
nand U9329 (N_9329,N_4102,N_5712);
xnor U9330 (N_9330,N_7193,N_4439);
and U9331 (N_9331,N_7467,N_7317);
and U9332 (N_9332,N_4488,N_7155);
nor U9333 (N_9333,N_5220,N_5440);
or U9334 (N_9334,N_7764,N_4006);
and U9335 (N_9335,N_4519,N_4057);
or U9336 (N_9336,N_6009,N_6927);
or U9337 (N_9337,N_5447,N_7935);
nand U9338 (N_9338,N_4994,N_6792);
nor U9339 (N_9339,N_6578,N_4495);
nor U9340 (N_9340,N_4332,N_5970);
and U9341 (N_9341,N_4897,N_6194);
or U9342 (N_9342,N_5053,N_6561);
and U9343 (N_9343,N_7195,N_6800);
nand U9344 (N_9344,N_7360,N_6200);
nor U9345 (N_9345,N_7706,N_7354);
or U9346 (N_9346,N_4825,N_5695);
nor U9347 (N_9347,N_4752,N_5748);
nand U9348 (N_9348,N_7600,N_4076);
and U9349 (N_9349,N_4701,N_5966);
and U9350 (N_9350,N_5830,N_5575);
nand U9351 (N_9351,N_5750,N_7388);
and U9352 (N_9352,N_5062,N_7960);
nand U9353 (N_9353,N_4297,N_5267);
and U9354 (N_9354,N_4053,N_6896);
nand U9355 (N_9355,N_4074,N_5025);
and U9356 (N_9356,N_5206,N_7192);
or U9357 (N_9357,N_7164,N_4661);
and U9358 (N_9358,N_4011,N_6624);
nor U9359 (N_9359,N_5877,N_6412);
nand U9360 (N_9360,N_5992,N_4031);
or U9361 (N_9361,N_5820,N_4720);
nand U9362 (N_9362,N_6398,N_4086);
nand U9363 (N_9363,N_5615,N_4608);
xnor U9364 (N_9364,N_7244,N_4261);
nor U9365 (N_9365,N_7012,N_4252);
and U9366 (N_9366,N_4755,N_6647);
nand U9367 (N_9367,N_6407,N_6440);
xnor U9368 (N_9368,N_7392,N_7323);
nor U9369 (N_9369,N_4254,N_6950);
nand U9370 (N_9370,N_7771,N_6779);
and U9371 (N_9371,N_7951,N_5761);
nor U9372 (N_9372,N_7184,N_5434);
xor U9373 (N_9373,N_5864,N_6447);
and U9374 (N_9374,N_6782,N_6338);
or U9375 (N_9375,N_4369,N_6244);
nor U9376 (N_9376,N_7516,N_4168);
or U9377 (N_9377,N_5419,N_5233);
and U9378 (N_9378,N_5790,N_4845);
nand U9379 (N_9379,N_5499,N_4811);
nand U9380 (N_9380,N_6914,N_4352);
and U9381 (N_9381,N_7697,N_4050);
nor U9382 (N_9382,N_4746,N_6755);
nand U9383 (N_9383,N_5194,N_4286);
or U9384 (N_9384,N_6100,N_4155);
and U9385 (N_9385,N_4573,N_6053);
nor U9386 (N_9386,N_7325,N_4022);
or U9387 (N_9387,N_6258,N_6587);
nand U9388 (N_9388,N_6423,N_5063);
or U9389 (N_9389,N_5436,N_7750);
nor U9390 (N_9390,N_5099,N_7639);
and U9391 (N_9391,N_7433,N_6332);
xnor U9392 (N_9392,N_5466,N_5884);
or U9393 (N_9393,N_4725,N_5807);
and U9394 (N_9394,N_6184,N_4325);
or U9395 (N_9395,N_5678,N_7368);
and U9396 (N_9396,N_6679,N_6640);
and U9397 (N_9397,N_5407,N_7525);
nand U9398 (N_9398,N_4362,N_4004);
nand U9399 (N_9399,N_6350,N_4485);
nor U9400 (N_9400,N_5676,N_4135);
xnor U9401 (N_9401,N_7243,N_7369);
or U9402 (N_9402,N_6892,N_7714);
nand U9403 (N_9403,N_4220,N_7690);
and U9404 (N_9404,N_7523,N_6179);
nand U9405 (N_9405,N_5768,N_6099);
nand U9406 (N_9406,N_7384,N_7187);
xnor U9407 (N_9407,N_5495,N_4487);
nand U9408 (N_9408,N_6805,N_4450);
or U9409 (N_9409,N_6916,N_5209);
nor U9410 (N_9410,N_5254,N_6195);
and U9411 (N_9411,N_6209,N_5931);
nor U9412 (N_9412,N_6062,N_4787);
nand U9413 (N_9413,N_7021,N_4695);
nor U9414 (N_9414,N_6228,N_5321);
and U9415 (N_9415,N_5429,N_7971);
nor U9416 (N_9416,N_6696,N_5480);
nor U9417 (N_9417,N_7819,N_5721);
xor U9418 (N_9418,N_7444,N_6666);
nor U9419 (N_9419,N_5837,N_4592);
nor U9420 (N_9420,N_4674,N_6242);
nor U9421 (N_9421,N_7509,N_4991);
nor U9422 (N_9422,N_5887,N_7831);
nand U9423 (N_9423,N_4237,N_7170);
or U9424 (N_9424,N_6523,N_4956);
nor U9425 (N_9425,N_7178,N_4882);
nand U9426 (N_9426,N_4802,N_6337);
or U9427 (N_9427,N_6095,N_6863);
and U9428 (N_9428,N_5980,N_7659);
nor U9429 (N_9429,N_7854,N_4620);
nor U9430 (N_9430,N_7462,N_6593);
or U9431 (N_9431,N_4651,N_4308);
or U9432 (N_9432,N_4844,N_5388);
and U9433 (N_9433,N_7484,N_4758);
nand U9434 (N_9434,N_5570,N_4020);
and U9435 (N_9435,N_7114,N_6827);
and U9436 (N_9436,N_7655,N_5189);
and U9437 (N_9437,N_7482,N_4636);
nand U9438 (N_9438,N_7877,N_6417);
and U9439 (N_9439,N_6512,N_4340);
and U9440 (N_9440,N_4995,N_4563);
nor U9441 (N_9441,N_6562,N_7016);
nor U9442 (N_9442,N_6161,N_7698);
and U9443 (N_9443,N_5276,N_7173);
nor U9444 (N_9444,N_5071,N_4547);
xnor U9445 (N_9445,N_4872,N_5323);
or U9446 (N_9446,N_5098,N_4570);
nor U9447 (N_9447,N_5719,N_5294);
and U9448 (N_9448,N_6643,N_4997);
and U9449 (N_9449,N_5703,N_7110);
xor U9450 (N_9450,N_5292,N_7860);
and U9451 (N_9451,N_7868,N_6124);
and U9452 (N_9452,N_6378,N_6848);
or U9453 (N_9453,N_6306,N_7737);
or U9454 (N_9454,N_6754,N_5990);
xor U9455 (N_9455,N_5416,N_4797);
or U9456 (N_9456,N_4700,N_4090);
and U9457 (N_9457,N_5564,N_5935);
and U9458 (N_9458,N_7411,N_5017);
and U9459 (N_9459,N_6733,N_4188);
and U9460 (N_9460,N_4327,N_6937);
nand U9461 (N_9461,N_6381,N_4510);
xor U9462 (N_9462,N_4932,N_4289);
xnor U9463 (N_9463,N_4663,N_7309);
or U9464 (N_9464,N_5862,N_5609);
nand U9465 (N_9465,N_7535,N_4222);
or U9466 (N_9466,N_5987,N_6205);
or U9467 (N_9467,N_4887,N_6434);
and U9468 (N_9468,N_4783,N_5967);
xnor U9469 (N_9469,N_4925,N_6579);
xor U9470 (N_9470,N_7577,N_4799);
or U9471 (N_9471,N_4640,N_4943);
or U9472 (N_9472,N_7949,N_5468);
or U9473 (N_9473,N_5944,N_7416);
nand U9474 (N_9474,N_4745,N_5608);
nor U9475 (N_9475,N_5946,N_4262);
nor U9476 (N_9476,N_7914,N_6316);
nor U9477 (N_9477,N_7007,N_7796);
or U9478 (N_9478,N_6961,N_6268);
nor U9479 (N_9479,N_5852,N_5546);
xor U9480 (N_9480,N_7508,N_5187);
or U9481 (N_9481,N_4858,N_6444);
nor U9482 (N_9482,N_4115,N_7787);
nor U9483 (N_9483,N_5637,N_4848);
nand U9484 (N_9484,N_5389,N_7292);
xor U9485 (N_9485,N_6743,N_6097);
or U9486 (N_9486,N_5223,N_6815);
and U9487 (N_9487,N_7082,N_5306);
or U9488 (N_9488,N_6185,N_5910);
and U9489 (N_9489,N_7647,N_5597);
nor U9490 (N_9490,N_6222,N_5181);
and U9491 (N_9491,N_7047,N_5201);
or U9492 (N_9492,N_6451,N_4737);
xor U9493 (N_9493,N_6703,N_7376);
or U9494 (N_9494,N_6343,N_5050);
nand U9495 (N_9495,N_5998,N_7822);
nand U9496 (N_9496,N_4598,N_4148);
or U9497 (N_9497,N_6445,N_5778);
nand U9498 (N_9498,N_7955,N_5785);
and U9499 (N_9499,N_7858,N_6390);
nand U9500 (N_9500,N_6701,N_7747);
nand U9501 (N_9501,N_5224,N_5083);
nor U9502 (N_9502,N_7603,N_6636);
nand U9503 (N_9503,N_7562,N_7410);
xor U9504 (N_9504,N_7396,N_7511);
nor U9505 (N_9505,N_7321,N_6830);
xnor U9506 (N_9506,N_4648,N_7367);
nor U9507 (N_9507,N_5972,N_4578);
nor U9508 (N_9508,N_7593,N_6355);
or U9509 (N_9509,N_7729,N_7269);
nor U9510 (N_9510,N_6741,N_4479);
nand U9511 (N_9511,N_4675,N_7962);
nand U9512 (N_9512,N_6943,N_6018);
and U9513 (N_9513,N_6702,N_5237);
nand U9514 (N_9514,N_4807,N_4202);
xnor U9515 (N_9515,N_4313,N_5620);
nor U9516 (N_9516,N_6889,N_6909);
nor U9517 (N_9517,N_7385,N_6418);
and U9518 (N_9518,N_6457,N_7488);
and U9519 (N_9519,N_6450,N_4472);
nand U9520 (N_9520,N_4962,N_6980);
nor U9521 (N_9521,N_6151,N_7870);
or U9522 (N_9522,N_7693,N_5929);
or U9523 (N_9523,N_7586,N_6190);
and U9524 (N_9524,N_7076,N_4413);
nand U9525 (N_9525,N_6022,N_5508);
and U9526 (N_9526,N_5069,N_7439);
and U9527 (N_9527,N_7260,N_5941);
and U9528 (N_9528,N_6507,N_6064);
nand U9529 (N_9529,N_4035,N_6255);
nor U9530 (N_9530,N_7086,N_5081);
nor U9531 (N_9531,N_6776,N_7680);
nor U9532 (N_9532,N_5212,N_5121);
nand U9533 (N_9533,N_5713,N_7526);
and U9534 (N_9534,N_6934,N_4888);
and U9535 (N_9535,N_4527,N_7621);
xor U9536 (N_9536,N_5774,N_6386);
nand U9537 (N_9537,N_6026,N_4371);
and U9538 (N_9538,N_6493,N_7404);
nor U9539 (N_9539,N_4772,N_5997);
nor U9540 (N_9540,N_6016,N_7234);
and U9541 (N_9541,N_5666,N_4719);
nand U9542 (N_9542,N_4567,N_4558);
nand U9543 (N_9543,N_6890,N_5177);
nor U9544 (N_9544,N_6038,N_5264);
nor U9545 (N_9545,N_6144,N_5828);
nor U9546 (N_9546,N_5829,N_5737);
nand U9547 (N_9547,N_5635,N_5802);
and U9548 (N_9548,N_6380,N_6711);
nor U9549 (N_9549,N_6873,N_7584);
or U9550 (N_9550,N_6697,N_4019);
and U9551 (N_9551,N_6475,N_6041);
and U9552 (N_9552,N_7703,N_7736);
nand U9553 (N_9553,N_6389,N_6043);
and U9554 (N_9554,N_7862,N_4410);
nor U9555 (N_9555,N_6661,N_6662);
or U9556 (N_9556,N_5219,N_4738);
and U9557 (N_9557,N_5599,N_5976);
or U9558 (N_9558,N_4576,N_4704);
nor U9559 (N_9559,N_4654,N_7327);
or U9560 (N_9560,N_4156,N_4458);
and U9561 (N_9561,N_4603,N_5093);
or U9562 (N_9562,N_5584,N_6363);
nor U9563 (N_9563,N_5640,N_4942);
nand U9564 (N_9564,N_6663,N_7876);
and U9565 (N_9565,N_6556,N_6452);
nor U9566 (N_9566,N_6871,N_6947);
nor U9567 (N_9567,N_5907,N_4079);
or U9568 (N_9568,N_4324,N_6615);
and U9569 (N_9569,N_5067,N_5699);
xnor U9570 (N_9570,N_4808,N_6485);
nor U9571 (N_9571,N_7364,N_4650);
nor U9572 (N_9572,N_7063,N_5986);
and U9573 (N_9573,N_6189,N_6329);
nand U9574 (N_9574,N_6686,N_6084);
nand U9575 (N_9575,N_4589,N_7052);
nor U9576 (N_9576,N_4973,N_4280);
nor U9577 (N_9577,N_5175,N_5965);
nand U9578 (N_9578,N_6560,N_7465);
and U9579 (N_9579,N_6524,N_5203);
xor U9580 (N_9580,N_4357,N_4532);
or U9581 (N_9581,N_4622,N_7528);
and U9582 (N_9582,N_6481,N_6059);
or U9583 (N_9583,N_4716,N_4985);
nand U9584 (N_9584,N_6780,N_6724);
or U9585 (N_9585,N_4918,N_6822);
xnor U9586 (N_9586,N_5125,N_6076);
or U9587 (N_9587,N_6221,N_5369);
nand U9588 (N_9588,N_7183,N_7390);
nor U9589 (N_9589,N_7479,N_7050);
and U9590 (N_9590,N_6424,N_5743);
nor U9591 (N_9591,N_5808,N_5155);
and U9592 (N_9592,N_4538,N_7256);
or U9593 (N_9593,N_5560,N_4877);
xnor U9594 (N_9594,N_4290,N_7158);
or U9595 (N_9595,N_5888,N_5816);
nand U9596 (N_9596,N_7109,N_4506);
xor U9597 (N_9597,N_5586,N_7631);
nor U9598 (N_9598,N_6888,N_4151);
nor U9599 (N_9599,N_6844,N_7564);
or U9600 (N_9600,N_7293,N_6528);
nand U9601 (N_9601,N_7464,N_5152);
or U9602 (N_9602,N_7033,N_5169);
and U9603 (N_9603,N_6093,N_5648);
nor U9604 (N_9604,N_7529,N_5927);
xnor U9605 (N_9605,N_6314,N_4326);
or U9606 (N_9606,N_5819,N_6981);
xor U9607 (N_9607,N_7219,N_5486);
and U9608 (N_9608,N_6957,N_7143);
nor U9609 (N_9609,N_5059,N_4292);
xnor U9610 (N_9610,N_4207,N_5504);
or U9611 (N_9611,N_7172,N_6535);
nand U9612 (N_9612,N_5727,N_4191);
nor U9613 (N_9613,N_4780,N_6649);
and U9614 (N_9614,N_4046,N_4481);
nand U9615 (N_9615,N_4253,N_7685);
nand U9616 (N_9616,N_7305,N_6870);
and U9617 (N_9617,N_7456,N_5020);
xnor U9618 (N_9618,N_5268,N_4049);
nor U9619 (N_9619,N_5590,N_7344);
nand U9620 (N_9620,N_7189,N_4370);
and U9621 (N_9621,N_5355,N_6214);
xor U9622 (N_9622,N_4304,N_6726);
nor U9623 (N_9623,N_4818,N_5298);
nand U9624 (N_9624,N_6285,N_7338);
nand U9625 (N_9625,N_5871,N_7229);
nor U9626 (N_9626,N_5897,N_4437);
nand U9627 (N_9627,N_6924,N_7989);
nand U9628 (N_9628,N_7040,N_7151);
and U9629 (N_9629,N_5399,N_6121);
nor U9630 (N_9630,N_7692,N_6902);
nor U9631 (N_9631,N_6881,N_7933);
nor U9632 (N_9632,N_6974,N_6054);
and U9633 (N_9633,N_6335,N_7137);
nand U9634 (N_9634,N_5188,N_5046);
nor U9635 (N_9635,N_6838,N_7899);
or U9636 (N_9636,N_4912,N_5744);
nor U9637 (N_9637,N_4416,N_4670);
and U9638 (N_9638,N_5475,N_6877);
nand U9639 (N_9639,N_7646,N_6219);
xor U9640 (N_9640,N_7954,N_5469);
or U9641 (N_9641,N_7159,N_7412);
nand U9642 (N_9642,N_7069,N_4303);
or U9643 (N_9643,N_4054,N_5130);
nand U9644 (N_9644,N_6930,N_6677);
or U9645 (N_9645,N_7777,N_6530);
nand U9646 (N_9646,N_6799,N_6542);
or U9647 (N_9647,N_5824,N_5681);
nor U9648 (N_9648,N_5925,N_5385);
nand U9649 (N_9649,N_5936,N_5278);
or U9650 (N_9650,N_7643,N_5814);
nor U9651 (N_9651,N_4865,N_6685);
or U9652 (N_9652,N_7359,N_5329);
and U9653 (N_9653,N_4703,N_7780);
nor U9654 (N_9654,N_5911,N_6581);
nor U9655 (N_9655,N_7133,N_6596);
nor U9656 (N_9656,N_5423,N_5497);
nor U9657 (N_9657,N_4862,N_6760);
and U9658 (N_9658,N_4623,N_6071);
nand U9659 (N_9659,N_5890,N_4690);
nand U9660 (N_9660,N_5184,N_7902);
nor U9661 (N_9661,N_7671,N_5027);
xnor U9662 (N_9662,N_5652,N_7419);
xnor U9663 (N_9663,N_4647,N_7938);
nor U9664 (N_9664,N_5421,N_5710);
xor U9665 (N_9665,N_4633,N_7732);
nor U9666 (N_9666,N_5137,N_4378);
nor U9667 (N_9667,N_7494,N_4009);
nand U9668 (N_9668,N_6248,N_4641);
and U9669 (N_9669,N_7124,N_4708);
nand U9670 (N_9670,N_4238,N_6945);
nor U9671 (N_9671,N_7366,N_7930);
xnor U9672 (N_9672,N_4856,N_6999);
or U9673 (N_9673,N_7981,N_6015);
or U9674 (N_9674,N_5078,N_5146);
nand U9675 (N_9675,N_5847,N_4367);
and U9676 (N_9676,N_5461,N_4337);
xnor U9677 (N_9677,N_5600,N_6180);
nand U9678 (N_9678,N_5043,N_4449);
and U9679 (N_9679,N_4944,N_7422);
or U9680 (N_9680,N_6657,N_5221);
xor U9681 (N_9681,N_4627,N_6747);
nand U9682 (N_9682,N_6633,N_6122);
or U9683 (N_9683,N_7785,N_5511);
or U9684 (N_9684,N_6494,N_5439);
nor U9685 (N_9685,N_6473,N_7454);
nor U9686 (N_9686,N_4609,N_7447);
and U9687 (N_9687,N_7039,N_4424);
xnor U9688 (N_9688,N_4409,N_5286);
and U9689 (N_9689,N_6478,N_7927);
or U9690 (N_9690,N_4561,N_7129);
xor U9691 (N_9691,N_6545,N_5514);
nand U9692 (N_9692,N_4801,N_5196);
nand U9693 (N_9693,N_4794,N_6720);
nor U9694 (N_9694,N_7890,N_7036);
nor U9695 (N_9695,N_4474,N_5360);
and U9696 (N_9696,N_7969,N_5123);
nor U9697 (N_9697,N_4917,N_5492);
xnor U9698 (N_9698,N_7499,N_5477);
and U9699 (N_9699,N_7349,N_5489);
or U9700 (N_9700,N_6886,N_4757);
and U9701 (N_9701,N_4328,N_5538);
nor U9702 (N_9702,N_5437,N_7476);
or U9703 (N_9703,N_7783,N_4542);
or U9704 (N_9704,N_5875,N_7490);
nand U9705 (N_9705,N_5662,N_5418);
nand U9706 (N_9706,N_5991,N_5463);
or U9707 (N_9707,N_5459,N_7072);
or U9708 (N_9708,N_5909,N_6177);
and U9709 (N_9709,N_5547,N_5403);
xnor U9710 (N_9710,N_6798,N_6638);
nor U9711 (N_9711,N_4056,N_6137);
nand U9712 (N_9712,N_4467,N_5131);
nand U9713 (N_9713,N_4349,N_4152);
nor U9714 (N_9714,N_6922,N_4588);
nand U9715 (N_9715,N_5983,N_6654);
nand U9716 (N_9716,N_6278,N_6277);
xor U9717 (N_9717,N_7768,N_6042);
and U9718 (N_9718,N_6955,N_4494);
or U9719 (N_9719,N_5857,N_6096);
or U9720 (N_9720,N_7898,N_7614);
and U9721 (N_9721,N_4101,N_5311);
and U9722 (N_9722,N_7424,N_5172);
xnor U9723 (N_9723,N_6206,N_7720);
nor U9724 (N_9724,N_6970,N_7667);
nand U9725 (N_9725,N_7632,N_4190);
and U9726 (N_9726,N_7669,N_5955);
nor U9727 (N_9727,N_5924,N_4549);
nand U9728 (N_9728,N_7653,N_5694);
nand U9729 (N_9729,N_5988,N_4240);
nor U9730 (N_9730,N_6324,N_5470);
or U9731 (N_9731,N_7686,N_6150);
and U9732 (N_9732,N_6516,N_7987);
xnor U9733 (N_9733,N_6068,N_5210);
nand U9734 (N_9734,N_5424,N_4990);
or U9735 (N_9735,N_4425,N_5047);
nand U9736 (N_9736,N_4816,N_7555);
nor U9737 (N_9737,N_4571,N_6591);
and U9738 (N_9738,N_6783,N_5811);
nand U9739 (N_9739,N_4198,N_5679);
nor U9740 (N_9740,N_5901,N_5588);
xor U9741 (N_9741,N_6859,N_4471);
nand U9742 (N_9742,N_5556,N_5800);
or U9743 (N_9743,N_4376,N_7804);
nand U9744 (N_9744,N_5000,N_4028);
nand U9745 (N_9745,N_5370,N_6522);
or U9746 (N_9746,N_7333,N_4284);
or U9747 (N_9747,N_5349,N_5680);
and U9748 (N_9748,N_5739,N_4263);
nand U9749 (N_9749,N_5630,N_5478);
and U9750 (N_9750,N_4180,N_5170);
and U9751 (N_9751,N_7576,N_5451);
and U9752 (N_9752,N_6170,N_7966);
nor U9753 (N_9753,N_6575,N_5122);
nor U9754 (N_9754,N_5420,N_7828);
and U9755 (N_9755,N_5571,N_5529);
or U9756 (N_9756,N_5287,N_4255);
nor U9757 (N_9757,N_5250,N_7035);
xnor U9758 (N_9758,N_7002,N_7790);
xnor U9759 (N_9759,N_5889,N_4172);
or U9760 (N_9760,N_4669,N_7162);
nor U9761 (N_9761,N_5491,N_6939);
xnor U9762 (N_9762,N_5559,N_4000);
nor U9763 (N_9763,N_5704,N_6550);
nor U9764 (N_9764,N_7637,N_6929);
and U9765 (N_9765,N_7548,N_5380);
nor U9766 (N_9766,N_6236,N_7817);
or U9767 (N_9767,N_7221,N_7607);
and U9768 (N_9768,N_7379,N_4098);
nor U9769 (N_9769,N_6356,N_6603);
or U9770 (N_9770,N_5338,N_5673);
or U9771 (N_9771,N_7077,N_5247);
xor U9772 (N_9772,N_6841,N_6187);
nand U9773 (N_9773,N_7688,N_7559);
xnor U9774 (N_9774,N_5843,N_4452);
nand U9775 (N_9775,N_6051,N_5707);
or U9776 (N_9776,N_7840,N_5994);
and U9777 (N_9777,N_6932,N_5231);
xnor U9778 (N_9778,N_7283,N_6917);
and U9779 (N_9779,N_5962,N_6972);
nor U9780 (N_9780,N_5263,N_7339);
nand U9781 (N_9781,N_5411,N_4501);
or U9782 (N_9782,N_5521,N_7994);
xor U9783 (N_9783,N_7345,N_7202);
nand U9784 (N_9784,N_7250,N_6519);
nor U9785 (N_9785,N_4614,N_4091);
or U9786 (N_9786,N_6327,N_7473);
or U9787 (N_9787,N_4412,N_4317);
nor U9788 (N_9788,N_6586,N_6166);
nand U9789 (N_9789,N_6202,N_6401);
or U9790 (N_9790,N_7613,N_7554);
and U9791 (N_9791,N_6029,N_4830);
nand U9792 (N_9792,N_5663,N_4335);
or U9793 (N_9793,N_4275,N_7242);
nand U9794 (N_9794,N_4868,N_6895);
and U9795 (N_9795,N_4557,N_5726);
nand U9796 (N_9796,N_6639,N_7487);
xor U9797 (N_9797,N_6862,N_7965);
nand U9798 (N_9798,N_6730,N_5865);
and U9799 (N_9799,N_5425,N_6631);
and U9800 (N_9800,N_5334,N_7766);
nor U9801 (N_9801,N_7061,N_6936);
nand U9802 (N_9802,N_5049,N_6483);
xnor U9803 (N_9803,N_6072,N_6346);
xor U9804 (N_9804,N_7742,N_5473);
or U9805 (N_9805,N_4843,N_5318);
nor U9806 (N_9806,N_7901,N_4300);
nand U9807 (N_9807,N_4713,N_7148);
nor U9808 (N_9808,N_7451,N_5873);
or U9809 (N_9809,N_6115,N_6461);
nand U9810 (N_9810,N_6098,N_7267);
or U9811 (N_9811,N_4852,N_6156);
nand U9812 (N_9812,N_7515,N_4192);
nor U9813 (N_9813,N_6287,N_4374);
nor U9814 (N_9814,N_5921,N_7812);
or U9815 (N_9815,N_5126,N_5741);
and U9816 (N_9816,N_6513,N_6080);
nor U9817 (N_9817,N_4898,N_6463);
and U9818 (N_9818,N_4377,N_5102);
nor U9819 (N_9819,N_6810,N_5297);
nor U9820 (N_9820,N_4444,N_7225);
xnor U9821 (N_9821,N_5671,N_5252);
or U9822 (N_9822,N_5957,N_6727);
nor U9823 (N_9823,N_4392,N_5465);
or U9824 (N_9824,N_7910,N_7443);
or U9825 (N_9825,N_5796,N_7071);
nor U9826 (N_9826,N_7081,N_5070);
nor U9827 (N_9827,N_5522,N_4595);
nor U9828 (N_9828,N_6849,N_6272);
and U9829 (N_9829,N_7203,N_7662);
and U9830 (N_9830,N_6653,N_5725);
nand U9831 (N_9831,N_5657,N_6520);
or U9832 (N_9832,N_4478,N_7409);
nor U9833 (N_9833,N_5801,N_7709);
and U9834 (N_9834,N_4500,N_5858);
nor U9835 (N_9835,N_7119,N_7008);
or U9836 (N_9836,N_6835,N_4040);
nand U9837 (N_9837,N_5686,N_6858);
or U9838 (N_9838,N_6453,N_6606);
xnor U9839 (N_9839,N_5782,N_7000);
and U9840 (N_9840,N_7299,N_5952);
and U9841 (N_9841,N_7112,N_5918);
or U9842 (N_9842,N_4554,N_7961);
or U9843 (N_9843,N_7059,N_7976);
nand U9844 (N_9844,N_7745,N_4833);
nand U9845 (N_9845,N_7105,N_7672);
nand U9846 (N_9846,N_6689,N_4914);
or U9847 (N_9847,N_6178,N_4431);
or U9848 (N_9848,N_7755,N_4063);
nor U9849 (N_9849,N_6832,N_5079);
or U9850 (N_9850,N_4143,N_4671);
nor U9851 (N_9851,N_4164,N_5258);
nand U9852 (N_9852,N_6665,N_6128);
and U9853 (N_9853,N_5689,N_4319);
nand U9854 (N_9854,N_6660,N_7037);
nor U9855 (N_9855,N_4939,N_5577);
and U9856 (N_9856,N_6087,N_5215);
nor U9857 (N_9857,N_4415,N_6379);
nor U9858 (N_9858,N_5930,N_4545);
or U9859 (N_9859,N_5031,N_4732);
nor U9860 (N_9860,N_6646,N_7252);
nand U9861 (N_9861,N_7986,N_4721);
or U9862 (N_9862,N_7958,N_5101);
nand U9863 (N_9863,N_7264,N_7625);
and U9864 (N_9864,N_7813,N_4630);
and U9865 (N_9865,N_4456,N_4283);
nand U9866 (N_9866,N_6469,N_6243);
nor U9867 (N_9867,N_4441,N_4591);
nor U9868 (N_9868,N_6669,N_4553);
and U9869 (N_9869,N_7136,N_6923);
nor U9870 (N_9870,N_6589,N_5225);
and U9871 (N_9871,N_5765,N_6951);
xnor U9872 (N_9872,N_7440,N_7903);
and U9873 (N_9873,N_7097,N_5174);
nor U9874 (N_9874,N_5346,N_5940);
or U9875 (N_9875,N_4331,N_7044);
xnor U9876 (N_9876,N_4067,N_6719);
nor U9877 (N_9877,N_7108,N_4257);
and U9878 (N_9878,N_7062,N_7306);
nand U9879 (N_9879,N_6046,N_4980);
and U9880 (N_9880,N_6814,N_7474);
and U9881 (N_9881,N_6330,N_4516);
or U9882 (N_9882,N_5054,N_6908);
and U9883 (N_9883,N_7478,N_4715);
nand U9884 (N_9884,N_7153,N_7552);
nand U9885 (N_9885,N_4607,N_4935);
nand U9886 (N_9886,N_7311,N_4181);
nor U9887 (N_9887,N_5638,N_4741);
or U9888 (N_9888,N_5351,N_7064);
nand U9889 (N_9889,N_5285,N_4137);
nor U9890 (N_9890,N_5973,N_7212);
and U9891 (N_9891,N_6250,N_5171);
and U9892 (N_9892,N_7280,N_5222);
nand U9893 (N_9893,N_6382,N_5660);
nand U9894 (N_9894,N_6642,N_7132);
and U9895 (N_9895,N_7266,N_4206);
and U9896 (N_9896,N_5127,N_7092);
or U9897 (N_9897,N_4694,N_4311);
and U9898 (N_9898,N_7932,N_5392);
nor U9899 (N_9899,N_4601,N_5467);
or U9900 (N_9900,N_4336,N_4976);
or U9901 (N_9901,N_6246,N_6789);
nand U9902 (N_9902,N_4301,N_7310);
nand U9903 (N_9903,N_4712,N_6432);
nand U9904 (N_9904,N_7303,N_5432);
or U9905 (N_9905,N_4743,N_6395);
nor U9906 (N_9906,N_4572,N_5274);
nor U9907 (N_9907,N_4653,N_6392);
or U9908 (N_9908,N_4434,N_7589);
or U9909 (N_9909,N_7839,N_6539);
or U9910 (N_9910,N_4574,N_7596);
nor U9911 (N_9911,N_5353,N_4658);
or U9912 (N_9912,N_5545,N_6245);
nand U9913 (N_9913,N_7186,N_4666);
or U9914 (N_9914,N_5077,N_6571);
nor U9915 (N_9915,N_5948,N_6831);
xor U9916 (N_9916,N_7536,N_4930);
xor U9917 (N_9917,N_5090,N_6975);
and U9918 (N_9918,N_5659,N_5786);
or U9919 (N_9919,N_7263,N_4890);
or U9920 (N_9920,N_7866,N_5372);
nand U9921 (N_9921,N_4373,N_7051);
and U9922 (N_9922,N_7314,N_6570);
or U9923 (N_9923,N_5526,N_4933);
and U9924 (N_9924,N_6992,N_7922);
and U9925 (N_9925,N_7191,N_7502);
and U9926 (N_9926,N_7834,N_7758);
nand U9927 (N_9927,N_5364,N_4265);
xor U9928 (N_9928,N_4676,N_5541);
nor U9929 (N_9929,N_4748,N_5904);
nand U9930 (N_9930,N_5717,N_7627);
xor U9931 (N_9931,N_5947,N_6429);
nor U9932 (N_9932,N_7351,N_6173);
nand U9933 (N_9933,N_4037,N_6998);
and U9934 (N_9934,N_7850,N_5592);
or U9935 (N_9935,N_5417,N_4140);
xor U9936 (N_9936,N_4126,N_4459);
or U9937 (N_9937,N_4952,N_7660);
xnor U9938 (N_9938,N_6850,N_7200);
and U9939 (N_9939,N_5151,N_5060);
nor U9940 (N_9940,N_4185,N_6237);
nand U9941 (N_9941,N_7205,N_6127);
nor U9942 (N_9942,N_7622,N_5107);
and U9943 (N_9943,N_4537,N_7074);
and U9944 (N_9944,N_4365,N_7326);
nand U9945 (N_9945,N_4770,N_4706);
nor U9946 (N_9946,N_6496,N_4125);
nand U9947 (N_9947,N_7546,N_6845);
xnor U9948 (N_9948,N_5001,N_7140);
and U9949 (N_9949,N_7216,N_7677);
or U9950 (N_9950,N_7313,N_4763);
nand U9951 (N_9951,N_6618,N_5583);
and U9952 (N_9952,N_5827,N_4405);
nand U9953 (N_9953,N_5326,N_4878);
or U9954 (N_9954,N_6549,N_6753);
nor U9955 (N_9955,N_4196,N_5257);
or U9956 (N_9956,N_7803,N_6032);
nand U9957 (N_9957,N_7605,N_7913);
nand U9958 (N_9958,N_4579,N_7983);
nor U9959 (N_9959,N_7569,N_6773);
nor U9960 (N_9960,N_5979,N_4433);
nor U9961 (N_9961,N_6553,N_7656);
or U9962 (N_9962,N_4219,N_5012);
nor U9963 (N_9963,N_6648,N_4018);
or U9964 (N_9964,N_7402,N_4281);
nor U9965 (N_9965,N_4291,N_6135);
nor U9966 (N_9966,N_4103,N_5651);
nor U9967 (N_9967,N_4123,N_6425);
or U9968 (N_9968,N_6971,N_4274);
xor U9969 (N_9969,N_6770,N_5438);
or U9970 (N_9970,N_5576,N_6670);
or U9971 (N_9971,N_7318,N_5359);
nand U9972 (N_9972,N_4873,N_6201);
nor U9973 (N_9973,N_5195,N_5157);
nand U9974 (N_9974,N_4593,N_6531);
or U9975 (N_9975,N_5641,N_4711);
xor U9976 (N_9976,N_7599,N_5055);
or U9977 (N_9977,N_6868,N_6674);
nor U9978 (N_9978,N_4556,N_4972);
nor U9979 (N_9979,N_4071,N_6384);
and U9980 (N_9980,N_7238,N_7537);
nand U9981 (N_9981,N_4626,N_6208);
nand U9982 (N_9982,N_7257,N_6986);
nor U9983 (N_9983,N_4417,N_5701);
nand U9984 (N_9984,N_5457,N_6569);
nand U9985 (N_9985,N_4790,N_5383);
nand U9986 (N_9986,N_4351,N_6692);
nor U9987 (N_9987,N_7341,N_5826);
nand U9988 (N_9988,N_5029,N_7843);
nor U9989 (N_9989,N_5200,N_7255);
or U9990 (N_9990,N_6605,N_5144);
nor U9991 (N_9991,N_6410,N_4710);
nand U9992 (N_9992,N_6419,N_7401);
nor U9993 (N_9993,N_7365,N_4193);
nor U9994 (N_9994,N_7125,N_4165);
and U9995 (N_9995,N_5675,N_7115);
nand U9996 (N_9996,N_6416,N_5981);
nor U9997 (N_9997,N_5426,N_6347);
nor U9998 (N_9998,N_4246,N_4753);
nor U9999 (N_9999,N_4380,N_5091);
and U10000 (N_10000,N_6456,N_5151);
and U10001 (N_10001,N_5481,N_4673);
and U10002 (N_10002,N_4291,N_6634);
or U10003 (N_10003,N_4141,N_7979);
or U10004 (N_10004,N_6391,N_4645);
nor U10005 (N_10005,N_6677,N_5556);
and U10006 (N_10006,N_6069,N_7447);
or U10007 (N_10007,N_4881,N_7146);
nor U10008 (N_10008,N_5501,N_7739);
and U10009 (N_10009,N_4316,N_4114);
or U10010 (N_10010,N_6201,N_4292);
nor U10011 (N_10011,N_6786,N_6859);
xnor U10012 (N_10012,N_6553,N_7842);
or U10013 (N_10013,N_6352,N_7109);
or U10014 (N_10014,N_5785,N_4086);
nor U10015 (N_10015,N_7592,N_4147);
xnor U10016 (N_10016,N_5993,N_4077);
nand U10017 (N_10017,N_6685,N_6165);
and U10018 (N_10018,N_5450,N_7756);
and U10019 (N_10019,N_7437,N_5197);
and U10020 (N_10020,N_5940,N_4612);
nand U10021 (N_10021,N_5535,N_4420);
nor U10022 (N_10022,N_5578,N_7390);
nand U10023 (N_10023,N_5046,N_4589);
or U10024 (N_10024,N_5041,N_7028);
xnor U10025 (N_10025,N_7528,N_6976);
or U10026 (N_10026,N_7704,N_4071);
nor U10027 (N_10027,N_4322,N_4284);
nor U10028 (N_10028,N_6930,N_4777);
or U10029 (N_10029,N_5224,N_6168);
or U10030 (N_10030,N_5989,N_5374);
and U10031 (N_10031,N_5131,N_5490);
or U10032 (N_10032,N_5047,N_6554);
nand U10033 (N_10033,N_5914,N_5927);
nand U10034 (N_10034,N_5298,N_6183);
and U10035 (N_10035,N_5848,N_4340);
nor U10036 (N_10036,N_4835,N_7768);
nand U10037 (N_10037,N_4383,N_5684);
nand U10038 (N_10038,N_5606,N_4860);
and U10039 (N_10039,N_6375,N_7082);
nor U10040 (N_10040,N_5795,N_4759);
xnor U10041 (N_10041,N_5649,N_5719);
nand U10042 (N_10042,N_6264,N_5229);
or U10043 (N_10043,N_5688,N_6541);
nand U10044 (N_10044,N_5416,N_6836);
and U10045 (N_10045,N_6054,N_5967);
or U10046 (N_10046,N_5238,N_6072);
nor U10047 (N_10047,N_6016,N_4235);
nor U10048 (N_10048,N_6400,N_5030);
xor U10049 (N_10049,N_4789,N_5428);
and U10050 (N_10050,N_6674,N_4697);
nor U10051 (N_10051,N_5673,N_7876);
and U10052 (N_10052,N_5334,N_4775);
nor U10053 (N_10053,N_5303,N_6394);
nand U10054 (N_10054,N_4215,N_5312);
nand U10055 (N_10055,N_5743,N_6202);
or U10056 (N_10056,N_5800,N_4460);
or U10057 (N_10057,N_7295,N_7368);
nand U10058 (N_10058,N_6664,N_7929);
and U10059 (N_10059,N_6860,N_7116);
xnor U10060 (N_10060,N_7932,N_5346);
nor U10061 (N_10061,N_5480,N_5909);
nand U10062 (N_10062,N_4100,N_6216);
and U10063 (N_10063,N_7478,N_7066);
nor U10064 (N_10064,N_7384,N_4821);
xor U10065 (N_10065,N_4226,N_5800);
or U10066 (N_10066,N_6865,N_5963);
and U10067 (N_10067,N_5353,N_7313);
nand U10068 (N_10068,N_6848,N_7468);
and U10069 (N_10069,N_7105,N_4296);
or U10070 (N_10070,N_6303,N_4174);
and U10071 (N_10071,N_5382,N_4899);
nor U10072 (N_10072,N_6706,N_4014);
and U10073 (N_10073,N_5311,N_5206);
or U10074 (N_10074,N_5997,N_4044);
nand U10075 (N_10075,N_5186,N_5860);
nand U10076 (N_10076,N_6785,N_5115);
or U10077 (N_10077,N_6925,N_7846);
nor U10078 (N_10078,N_5224,N_6338);
nand U10079 (N_10079,N_6548,N_4570);
xnor U10080 (N_10080,N_5785,N_5906);
or U10081 (N_10081,N_5711,N_7573);
and U10082 (N_10082,N_6730,N_4766);
and U10083 (N_10083,N_6945,N_4393);
and U10084 (N_10084,N_6020,N_4644);
nand U10085 (N_10085,N_6679,N_7090);
nor U10086 (N_10086,N_6173,N_7069);
nand U10087 (N_10087,N_4549,N_5228);
nand U10088 (N_10088,N_6400,N_7912);
and U10089 (N_10089,N_4264,N_7614);
nor U10090 (N_10090,N_7338,N_6372);
and U10091 (N_10091,N_5827,N_7993);
and U10092 (N_10092,N_4231,N_6681);
nor U10093 (N_10093,N_4596,N_5018);
or U10094 (N_10094,N_4480,N_6462);
or U10095 (N_10095,N_5424,N_6743);
or U10096 (N_10096,N_4458,N_4021);
and U10097 (N_10097,N_7407,N_5276);
or U10098 (N_10098,N_4320,N_4424);
nand U10099 (N_10099,N_4243,N_4196);
nor U10100 (N_10100,N_5918,N_4384);
or U10101 (N_10101,N_4878,N_7558);
and U10102 (N_10102,N_6134,N_6991);
and U10103 (N_10103,N_7222,N_5922);
and U10104 (N_10104,N_4149,N_4883);
or U10105 (N_10105,N_6959,N_5960);
or U10106 (N_10106,N_4473,N_7426);
and U10107 (N_10107,N_5161,N_4806);
or U10108 (N_10108,N_4437,N_6276);
and U10109 (N_10109,N_5556,N_6696);
nor U10110 (N_10110,N_4953,N_7162);
xnor U10111 (N_10111,N_4905,N_5692);
nor U10112 (N_10112,N_6714,N_4947);
and U10113 (N_10113,N_5285,N_4340);
xnor U10114 (N_10114,N_7405,N_7980);
and U10115 (N_10115,N_4336,N_6408);
and U10116 (N_10116,N_5542,N_7088);
nor U10117 (N_10117,N_6885,N_6185);
xor U10118 (N_10118,N_7960,N_6297);
or U10119 (N_10119,N_5688,N_7181);
xor U10120 (N_10120,N_5787,N_5545);
nor U10121 (N_10121,N_4767,N_5093);
nand U10122 (N_10122,N_6315,N_5451);
nand U10123 (N_10123,N_6009,N_4004);
and U10124 (N_10124,N_6254,N_5181);
and U10125 (N_10125,N_7348,N_7197);
and U10126 (N_10126,N_5488,N_4699);
or U10127 (N_10127,N_5738,N_7047);
and U10128 (N_10128,N_7528,N_4434);
nor U10129 (N_10129,N_5131,N_6076);
nor U10130 (N_10130,N_6350,N_5178);
nand U10131 (N_10131,N_7965,N_6622);
nand U10132 (N_10132,N_5082,N_7589);
or U10133 (N_10133,N_5553,N_6065);
nor U10134 (N_10134,N_5838,N_4403);
or U10135 (N_10135,N_6189,N_4102);
nand U10136 (N_10136,N_4342,N_5319);
or U10137 (N_10137,N_7500,N_5965);
and U10138 (N_10138,N_7166,N_6790);
nand U10139 (N_10139,N_5657,N_5452);
nand U10140 (N_10140,N_5923,N_7765);
and U10141 (N_10141,N_5607,N_4436);
nand U10142 (N_10142,N_7111,N_7339);
nor U10143 (N_10143,N_7627,N_6365);
and U10144 (N_10144,N_5182,N_7649);
nor U10145 (N_10145,N_6075,N_5555);
xor U10146 (N_10146,N_5945,N_5039);
nor U10147 (N_10147,N_4027,N_4433);
nor U10148 (N_10148,N_6581,N_4473);
nand U10149 (N_10149,N_6146,N_6885);
or U10150 (N_10150,N_6279,N_5661);
and U10151 (N_10151,N_5365,N_5042);
or U10152 (N_10152,N_5450,N_6393);
nor U10153 (N_10153,N_6626,N_6897);
and U10154 (N_10154,N_4099,N_7489);
nand U10155 (N_10155,N_6712,N_5735);
or U10156 (N_10156,N_7939,N_4805);
and U10157 (N_10157,N_6743,N_7826);
nand U10158 (N_10158,N_4848,N_5209);
or U10159 (N_10159,N_5978,N_7506);
or U10160 (N_10160,N_4876,N_5137);
and U10161 (N_10161,N_4311,N_7166);
nand U10162 (N_10162,N_7049,N_6979);
and U10163 (N_10163,N_7346,N_4458);
and U10164 (N_10164,N_4205,N_5124);
nor U10165 (N_10165,N_6065,N_6791);
nor U10166 (N_10166,N_7795,N_4089);
nor U10167 (N_10167,N_7353,N_5262);
and U10168 (N_10168,N_6674,N_6474);
and U10169 (N_10169,N_6084,N_6181);
or U10170 (N_10170,N_6851,N_4978);
and U10171 (N_10171,N_7034,N_6127);
or U10172 (N_10172,N_4704,N_6150);
xor U10173 (N_10173,N_5612,N_5185);
or U10174 (N_10174,N_5189,N_4482);
nand U10175 (N_10175,N_5557,N_6578);
or U10176 (N_10176,N_4892,N_4475);
nand U10177 (N_10177,N_6476,N_4939);
and U10178 (N_10178,N_5996,N_6866);
or U10179 (N_10179,N_5881,N_7219);
and U10180 (N_10180,N_4826,N_7686);
xor U10181 (N_10181,N_7680,N_4840);
nand U10182 (N_10182,N_4227,N_4091);
or U10183 (N_10183,N_5322,N_4098);
or U10184 (N_10184,N_5492,N_5238);
nor U10185 (N_10185,N_6631,N_7116);
nor U10186 (N_10186,N_5231,N_6294);
nor U10187 (N_10187,N_6954,N_5249);
nor U10188 (N_10188,N_7311,N_5164);
xnor U10189 (N_10189,N_7407,N_4068);
and U10190 (N_10190,N_6752,N_7039);
and U10191 (N_10191,N_5062,N_5727);
and U10192 (N_10192,N_5124,N_7096);
and U10193 (N_10193,N_5436,N_6667);
nand U10194 (N_10194,N_5660,N_5189);
nor U10195 (N_10195,N_4700,N_5279);
or U10196 (N_10196,N_4479,N_6512);
or U10197 (N_10197,N_7084,N_6696);
nand U10198 (N_10198,N_5200,N_5965);
nand U10199 (N_10199,N_4670,N_4611);
nor U10200 (N_10200,N_7056,N_6315);
nor U10201 (N_10201,N_4323,N_6267);
nand U10202 (N_10202,N_6251,N_6615);
nor U10203 (N_10203,N_7821,N_4052);
nand U10204 (N_10204,N_7219,N_4409);
or U10205 (N_10205,N_5653,N_4432);
nand U10206 (N_10206,N_7547,N_5806);
nor U10207 (N_10207,N_7122,N_7529);
xnor U10208 (N_10208,N_4375,N_5461);
nor U10209 (N_10209,N_4550,N_5707);
or U10210 (N_10210,N_7322,N_7062);
and U10211 (N_10211,N_5691,N_4693);
nor U10212 (N_10212,N_7424,N_7197);
nand U10213 (N_10213,N_4286,N_5589);
or U10214 (N_10214,N_7772,N_7078);
nand U10215 (N_10215,N_4099,N_5387);
and U10216 (N_10216,N_4054,N_5389);
nor U10217 (N_10217,N_7874,N_7763);
or U10218 (N_10218,N_4242,N_5802);
and U10219 (N_10219,N_4762,N_6007);
nor U10220 (N_10220,N_6327,N_5499);
nor U10221 (N_10221,N_4156,N_4301);
and U10222 (N_10222,N_5594,N_5072);
nor U10223 (N_10223,N_7931,N_5336);
nand U10224 (N_10224,N_5733,N_6085);
nor U10225 (N_10225,N_7331,N_5755);
or U10226 (N_10226,N_5586,N_5212);
nor U10227 (N_10227,N_4975,N_6224);
and U10228 (N_10228,N_6456,N_4099);
nand U10229 (N_10229,N_6128,N_6895);
nand U10230 (N_10230,N_6823,N_6649);
nor U10231 (N_10231,N_6755,N_5428);
or U10232 (N_10232,N_7918,N_7072);
xor U10233 (N_10233,N_6743,N_7303);
nor U10234 (N_10234,N_4965,N_7827);
nand U10235 (N_10235,N_5237,N_4853);
and U10236 (N_10236,N_6723,N_6179);
nand U10237 (N_10237,N_7615,N_4153);
nor U10238 (N_10238,N_7383,N_5107);
or U10239 (N_10239,N_5900,N_7598);
xor U10240 (N_10240,N_4709,N_7318);
nand U10241 (N_10241,N_5243,N_7743);
nor U10242 (N_10242,N_5380,N_5350);
or U10243 (N_10243,N_6942,N_5221);
nand U10244 (N_10244,N_5706,N_7994);
xor U10245 (N_10245,N_4432,N_5381);
xnor U10246 (N_10246,N_4185,N_4609);
or U10247 (N_10247,N_5900,N_6759);
or U10248 (N_10248,N_6563,N_6670);
and U10249 (N_10249,N_6824,N_6476);
xor U10250 (N_10250,N_7869,N_6224);
nand U10251 (N_10251,N_4793,N_4927);
and U10252 (N_10252,N_7031,N_7166);
and U10253 (N_10253,N_4745,N_6654);
or U10254 (N_10254,N_5716,N_5503);
nand U10255 (N_10255,N_4800,N_7634);
or U10256 (N_10256,N_5581,N_4076);
xor U10257 (N_10257,N_5395,N_4398);
and U10258 (N_10258,N_7435,N_5170);
and U10259 (N_10259,N_4377,N_7683);
xnor U10260 (N_10260,N_6221,N_7145);
nand U10261 (N_10261,N_5311,N_7330);
nand U10262 (N_10262,N_4160,N_5766);
and U10263 (N_10263,N_4436,N_4117);
nor U10264 (N_10264,N_4547,N_6974);
and U10265 (N_10265,N_7290,N_4896);
nor U10266 (N_10266,N_7943,N_5324);
nor U10267 (N_10267,N_6463,N_6940);
and U10268 (N_10268,N_6875,N_4215);
and U10269 (N_10269,N_6215,N_7062);
or U10270 (N_10270,N_6033,N_4130);
nor U10271 (N_10271,N_7861,N_5314);
xor U10272 (N_10272,N_6751,N_7274);
or U10273 (N_10273,N_4543,N_5949);
nand U10274 (N_10274,N_5301,N_5091);
nor U10275 (N_10275,N_6710,N_5228);
or U10276 (N_10276,N_4455,N_4046);
nor U10277 (N_10277,N_6564,N_7389);
nor U10278 (N_10278,N_6106,N_6486);
or U10279 (N_10279,N_7022,N_5946);
nor U10280 (N_10280,N_7484,N_5880);
or U10281 (N_10281,N_5346,N_5744);
or U10282 (N_10282,N_4283,N_4750);
nand U10283 (N_10283,N_5865,N_6219);
nor U10284 (N_10284,N_6858,N_7275);
nor U10285 (N_10285,N_6129,N_5800);
and U10286 (N_10286,N_6684,N_6687);
and U10287 (N_10287,N_5190,N_4912);
or U10288 (N_10288,N_5998,N_6587);
nand U10289 (N_10289,N_4355,N_7579);
or U10290 (N_10290,N_7403,N_5241);
or U10291 (N_10291,N_7317,N_7508);
or U10292 (N_10292,N_5053,N_6587);
and U10293 (N_10293,N_6539,N_5179);
and U10294 (N_10294,N_5256,N_4033);
or U10295 (N_10295,N_7976,N_5709);
nand U10296 (N_10296,N_5114,N_4715);
or U10297 (N_10297,N_6574,N_7180);
nand U10298 (N_10298,N_7729,N_7956);
and U10299 (N_10299,N_6575,N_4341);
or U10300 (N_10300,N_4174,N_7159);
and U10301 (N_10301,N_7251,N_7680);
nor U10302 (N_10302,N_4877,N_4611);
or U10303 (N_10303,N_7517,N_4667);
or U10304 (N_10304,N_4172,N_5408);
xor U10305 (N_10305,N_7177,N_5894);
or U10306 (N_10306,N_5458,N_5794);
or U10307 (N_10307,N_7079,N_5401);
nor U10308 (N_10308,N_7085,N_4579);
nand U10309 (N_10309,N_7801,N_6349);
or U10310 (N_10310,N_6030,N_6088);
nand U10311 (N_10311,N_6224,N_7090);
nor U10312 (N_10312,N_5355,N_4870);
and U10313 (N_10313,N_5634,N_4587);
or U10314 (N_10314,N_5194,N_4564);
nor U10315 (N_10315,N_6920,N_7209);
xor U10316 (N_10316,N_5095,N_6626);
or U10317 (N_10317,N_7749,N_4557);
nor U10318 (N_10318,N_4094,N_6306);
and U10319 (N_10319,N_4125,N_5312);
nand U10320 (N_10320,N_6810,N_4007);
and U10321 (N_10321,N_6243,N_5449);
and U10322 (N_10322,N_7304,N_5464);
or U10323 (N_10323,N_7785,N_5810);
and U10324 (N_10324,N_4484,N_7440);
or U10325 (N_10325,N_5012,N_7090);
nand U10326 (N_10326,N_4442,N_7762);
and U10327 (N_10327,N_5687,N_5140);
nor U10328 (N_10328,N_5974,N_6532);
nor U10329 (N_10329,N_5088,N_7615);
nand U10330 (N_10330,N_5826,N_5776);
nand U10331 (N_10331,N_5396,N_5273);
or U10332 (N_10332,N_5427,N_5719);
nand U10333 (N_10333,N_7684,N_7144);
xor U10334 (N_10334,N_7431,N_5860);
nand U10335 (N_10335,N_6065,N_4064);
nor U10336 (N_10336,N_6477,N_7258);
or U10337 (N_10337,N_5467,N_6686);
nor U10338 (N_10338,N_6003,N_6045);
and U10339 (N_10339,N_5788,N_7672);
and U10340 (N_10340,N_5175,N_6599);
nor U10341 (N_10341,N_7634,N_7359);
nand U10342 (N_10342,N_4208,N_6188);
or U10343 (N_10343,N_7049,N_7361);
nor U10344 (N_10344,N_4151,N_4992);
and U10345 (N_10345,N_5247,N_7459);
nor U10346 (N_10346,N_6464,N_5511);
nor U10347 (N_10347,N_6163,N_7410);
nand U10348 (N_10348,N_5801,N_7449);
or U10349 (N_10349,N_7494,N_4467);
or U10350 (N_10350,N_5217,N_7609);
nand U10351 (N_10351,N_7319,N_7826);
nand U10352 (N_10352,N_6856,N_4430);
nand U10353 (N_10353,N_7986,N_4476);
nand U10354 (N_10354,N_7757,N_5998);
nor U10355 (N_10355,N_5475,N_5006);
or U10356 (N_10356,N_6839,N_6576);
or U10357 (N_10357,N_6311,N_4811);
and U10358 (N_10358,N_6634,N_4857);
nor U10359 (N_10359,N_6108,N_6530);
and U10360 (N_10360,N_4222,N_6098);
nor U10361 (N_10361,N_5449,N_7904);
nor U10362 (N_10362,N_4533,N_6113);
or U10363 (N_10363,N_5251,N_6878);
and U10364 (N_10364,N_6777,N_5363);
and U10365 (N_10365,N_6078,N_4082);
and U10366 (N_10366,N_4313,N_7659);
nor U10367 (N_10367,N_4984,N_5042);
nand U10368 (N_10368,N_5074,N_5987);
xnor U10369 (N_10369,N_4151,N_6237);
nand U10370 (N_10370,N_7203,N_4249);
or U10371 (N_10371,N_6529,N_7281);
or U10372 (N_10372,N_6445,N_4430);
and U10373 (N_10373,N_7165,N_5354);
nor U10374 (N_10374,N_6142,N_6813);
nor U10375 (N_10375,N_6574,N_6406);
nor U10376 (N_10376,N_6775,N_6661);
and U10377 (N_10377,N_6988,N_5674);
or U10378 (N_10378,N_6427,N_7893);
and U10379 (N_10379,N_4450,N_4580);
nand U10380 (N_10380,N_5176,N_6624);
and U10381 (N_10381,N_6911,N_7725);
nand U10382 (N_10382,N_5818,N_4097);
nand U10383 (N_10383,N_5794,N_6331);
xnor U10384 (N_10384,N_7041,N_4863);
or U10385 (N_10385,N_4539,N_7237);
nor U10386 (N_10386,N_5656,N_7722);
and U10387 (N_10387,N_5390,N_7367);
and U10388 (N_10388,N_4674,N_4691);
and U10389 (N_10389,N_5369,N_4457);
nand U10390 (N_10390,N_6864,N_6656);
or U10391 (N_10391,N_4839,N_5515);
or U10392 (N_10392,N_7551,N_5882);
nor U10393 (N_10393,N_6739,N_6752);
nor U10394 (N_10394,N_7463,N_7783);
nor U10395 (N_10395,N_4133,N_6972);
and U10396 (N_10396,N_4306,N_7010);
or U10397 (N_10397,N_6255,N_6079);
or U10398 (N_10398,N_6653,N_4310);
or U10399 (N_10399,N_7043,N_4045);
and U10400 (N_10400,N_5794,N_4521);
nand U10401 (N_10401,N_7394,N_7780);
nor U10402 (N_10402,N_7559,N_7780);
and U10403 (N_10403,N_6919,N_5984);
nand U10404 (N_10404,N_4336,N_6569);
or U10405 (N_10405,N_7915,N_7993);
or U10406 (N_10406,N_5316,N_4726);
nor U10407 (N_10407,N_5701,N_5201);
nand U10408 (N_10408,N_4062,N_7950);
and U10409 (N_10409,N_7456,N_6483);
nand U10410 (N_10410,N_4077,N_4267);
or U10411 (N_10411,N_7143,N_5175);
and U10412 (N_10412,N_6779,N_5082);
nand U10413 (N_10413,N_4887,N_5292);
nor U10414 (N_10414,N_4593,N_5021);
nand U10415 (N_10415,N_4414,N_4731);
and U10416 (N_10416,N_4218,N_7225);
or U10417 (N_10417,N_4125,N_4106);
and U10418 (N_10418,N_7461,N_7516);
nand U10419 (N_10419,N_4704,N_6464);
nand U10420 (N_10420,N_6488,N_5499);
and U10421 (N_10421,N_6211,N_6628);
and U10422 (N_10422,N_4916,N_7575);
nor U10423 (N_10423,N_5916,N_6654);
nand U10424 (N_10424,N_4054,N_5656);
xor U10425 (N_10425,N_6092,N_5624);
nand U10426 (N_10426,N_4623,N_4585);
nor U10427 (N_10427,N_7560,N_7380);
and U10428 (N_10428,N_6862,N_4265);
nor U10429 (N_10429,N_7498,N_4191);
and U10430 (N_10430,N_4964,N_4833);
or U10431 (N_10431,N_4720,N_5239);
or U10432 (N_10432,N_5766,N_7684);
nand U10433 (N_10433,N_6074,N_4476);
xnor U10434 (N_10434,N_4017,N_7803);
and U10435 (N_10435,N_6089,N_6189);
nor U10436 (N_10436,N_7995,N_4530);
or U10437 (N_10437,N_7225,N_7554);
and U10438 (N_10438,N_6277,N_5987);
or U10439 (N_10439,N_6238,N_7477);
and U10440 (N_10440,N_4842,N_6081);
and U10441 (N_10441,N_4210,N_7613);
and U10442 (N_10442,N_5196,N_5866);
and U10443 (N_10443,N_4958,N_7143);
xnor U10444 (N_10444,N_4830,N_7635);
and U10445 (N_10445,N_5954,N_5347);
or U10446 (N_10446,N_7434,N_6219);
nand U10447 (N_10447,N_4258,N_5285);
nor U10448 (N_10448,N_6839,N_7937);
nor U10449 (N_10449,N_5836,N_4859);
or U10450 (N_10450,N_4544,N_6932);
xor U10451 (N_10451,N_5763,N_4080);
or U10452 (N_10452,N_7617,N_5254);
or U10453 (N_10453,N_4422,N_7339);
or U10454 (N_10454,N_7093,N_5978);
or U10455 (N_10455,N_7196,N_4683);
xnor U10456 (N_10456,N_6557,N_5425);
xor U10457 (N_10457,N_7135,N_6362);
nand U10458 (N_10458,N_7493,N_4110);
nand U10459 (N_10459,N_5109,N_6011);
nand U10460 (N_10460,N_5321,N_7478);
nor U10461 (N_10461,N_7043,N_6853);
or U10462 (N_10462,N_5116,N_7641);
or U10463 (N_10463,N_6358,N_4025);
nor U10464 (N_10464,N_5828,N_6493);
nor U10465 (N_10465,N_6845,N_4619);
or U10466 (N_10466,N_5609,N_5506);
nor U10467 (N_10467,N_6330,N_5642);
nand U10468 (N_10468,N_5586,N_6954);
and U10469 (N_10469,N_5733,N_6778);
nor U10470 (N_10470,N_6026,N_4656);
nand U10471 (N_10471,N_6699,N_7749);
or U10472 (N_10472,N_7084,N_5137);
and U10473 (N_10473,N_5315,N_7563);
and U10474 (N_10474,N_5990,N_7676);
and U10475 (N_10475,N_7897,N_7724);
nor U10476 (N_10476,N_6036,N_5292);
or U10477 (N_10477,N_7928,N_7895);
nor U10478 (N_10478,N_4082,N_7306);
nor U10479 (N_10479,N_7237,N_4650);
nand U10480 (N_10480,N_5213,N_5115);
xnor U10481 (N_10481,N_5548,N_7138);
xnor U10482 (N_10482,N_6566,N_5301);
xor U10483 (N_10483,N_4033,N_6711);
or U10484 (N_10484,N_6602,N_4200);
nand U10485 (N_10485,N_7828,N_5025);
or U10486 (N_10486,N_5770,N_5959);
or U10487 (N_10487,N_5204,N_4648);
and U10488 (N_10488,N_4556,N_7551);
and U10489 (N_10489,N_7789,N_7884);
or U10490 (N_10490,N_6918,N_7510);
nand U10491 (N_10491,N_7859,N_6843);
xnor U10492 (N_10492,N_6855,N_6010);
nand U10493 (N_10493,N_5424,N_7878);
and U10494 (N_10494,N_6472,N_5303);
xor U10495 (N_10495,N_6471,N_6868);
nor U10496 (N_10496,N_6545,N_6995);
and U10497 (N_10497,N_5233,N_6873);
or U10498 (N_10498,N_7582,N_7193);
nor U10499 (N_10499,N_6723,N_5105);
nor U10500 (N_10500,N_6562,N_4807);
nand U10501 (N_10501,N_6842,N_6978);
nand U10502 (N_10502,N_7389,N_5287);
and U10503 (N_10503,N_5777,N_6341);
nand U10504 (N_10504,N_4748,N_5827);
and U10505 (N_10505,N_5269,N_4850);
nor U10506 (N_10506,N_7252,N_7998);
or U10507 (N_10507,N_6161,N_5168);
xor U10508 (N_10508,N_5255,N_5025);
nor U10509 (N_10509,N_4007,N_5204);
and U10510 (N_10510,N_4732,N_4016);
nor U10511 (N_10511,N_7330,N_4969);
and U10512 (N_10512,N_6047,N_7518);
nand U10513 (N_10513,N_5669,N_7740);
or U10514 (N_10514,N_6567,N_7298);
nand U10515 (N_10515,N_6558,N_5085);
nand U10516 (N_10516,N_7125,N_4951);
and U10517 (N_10517,N_7399,N_7296);
and U10518 (N_10518,N_4281,N_6539);
nor U10519 (N_10519,N_4557,N_5763);
nand U10520 (N_10520,N_4409,N_5553);
or U10521 (N_10521,N_7784,N_5893);
nor U10522 (N_10522,N_5811,N_4559);
or U10523 (N_10523,N_4361,N_7714);
or U10524 (N_10524,N_5084,N_6529);
or U10525 (N_10525,N_6225,N_5563);
nor U10526 (N_10526,N_7285,N_6901);
nand U10527 (N_10527,N_4164,N_6981);
nor U10528 (N_10528,N_6483,N_6150);
and U10529 (N_10529,N_4244,N_4153);
nor U10530 (N_10530,N_4723,N_7186);
nor U10531 (N_10531,N_7846,N_7440);
or U10532 (N_10532,N_5500,N_5123);
or U10533 (N_10533,N_7944,N_5285);
nor U10534 (N_10534,N_5427,N_7498);
and U10535 (N_10535,N_7727,N_6638);
or U10536 (N_10536,N_7640,N_6871);
nand U10537 (N_10537,N_7075,N_5240);
and U10538 (N_10538,N_5518,N_5782);
nand U10539 (N_10539,N_6325,N_4582);
nand U10540 (N_10540,N_6152,N_6162);
nor U10541 (N_10541,N_4401,N_7249);
nand U10542 (N_10542,N_5719,N_4999);
or U10543 (N_10543,N_4355,N_5748);
or U10544 (N_10544,N_5036,N_6639);
nor U10545 (N_10545,N_6065,N_6372);
nand U10546 (N_10546,N_4475,N_6290);
nand U10547 (N_10547,N_7547,N_6586);
or U10548 (N_10548,N_4694,N_6188);
xnor U10549 (N_10549,N_5833,N_7444);
and U10550 (N_10550,N_7997,N_7873);
or U10551 (N_10551,N_6777,N_5453);
and U10552 (N_10552,N_5107,N_5754);
nor U10553 (N_10553,N_6949,N_6836);
or U10554 (N_10554,N_4018,N_4224);
or U10555 (N_10555,N_6502,N_7657);
nor U10556 (N_10556,N_4884,N_7348);
nand U10557 (N_10557,N_4974,N_6533);
and U10558 (N_10558,N_5548,N_4090);
or U10559 (N_10559,N_5192,N_7768);
or U10560 (N_10560,N_6243,N_4469);
nand U10561 (N_10561,N_7150,N_5926);
nor U10562 (N_10562,N_6463,N_6962);
nor U10563 (N_10563,N_7646,N_7909);
or U10564 (N_10564,N_4838,N_7427);
and U10565 (N_10565,N_4728,N_7471);
or U10566 (N_10566,N_6421,N_4452);
nor U10567 (N_10567,N_4356,N_5890);
nor U10568 (N_10568,N_6618,N_7893);
nand U10569 (N_10569,N_7632,N_4955);
nand U10570 (N_10570,N_7808,N_4818);
or U10571 (N_10571,N_6063,N_5344);
and U10572 (N_10572,N_4506,N_6755);
and U10573 (N_10573,N_6056,N_4707);
xnor U10574 (N_10574,N_7351,N_5821);
nor U10575 (N_10575,N_5332,N_5714);
xnor U10576 (N_10576,N_4586,N_5947);
nand U10577 (N_10577,N_7897,N_4794);
nand U10578 (N_10578,N_7539,N_5134);
nor U10579 (N_10579,N_5063,N_4690);
nor U10580 (N_10580,N_4218,N_6099);
or U10581 (N_10581,N_4461,N_4785);
xor U10582 (N_10582,N_5488,N_5094);
xnor U10583 (N_10583,N_4889,N_6238);
and U10584 (N_10584,N_6863,N_5533);
or U10585 (N_10585,N_7131,N_5939);
and U10586 (N_10586,N_5891,N_5239);
nand U10587 (N_10587,N_6909,N_4558);
nand U10588 (N_10588,N_6306,N_7532);
or U10589 (N_10589,N_4285,N_7699);
and U10590 (N_10590,N_4730,N_5010);
nor U10591 (N_10591,N_5923,N_7264);
xnor U10592 (N_10592,N_5621,N_7671);
nand U10593 (N_10593,N_4232,N_5256);
xor U10594 (N_10594,N_4755,N_5632);
xor U10595 (N_10595,N_6012,N_5774);
nor U10596 (N_10596,N_4325,N_7473);
and U10597 (N_10597,N_5659,N_5459);
and U10598 (N_10598,N_7873,N_4714);
and U10599 (N_10599,N_7351,N_7623);
nor U10600 (N_10600,N_7719,N_7876);
nor U10601 (N_10601,N_6718,N_5280);
and U10602 (N_10602,N_6980,N_7521);
and U10603 (N_10603,N_7746,N_4916);
nand U10604 (N_10604,N_7542,N_4112);
or U10605 (N_10605,N_4397,N_5588);
xnor U10606 (N_10606,N_4910,N_6234);
nor U10607 (N_10607,N_7914,N_6550);
nor U10608 (N_10608,N_6583,N_6200);
nand U10609 (N_10609,N_7003,N_6899);
nor U10610 (N_10610,N_5007,N_6554);
nand U10611 (N_10611,N_7762,N_5534);
nand U10612 (N_10612,N_7160,N_4766);
or U10613 (N_10613,N_6698,N_7728);
nor U10614 (N_10614,N_4093,N_5783);
or U10615 (N_10615,N_4746,N_6092);
nand U10616 (N_10616,N_4394,N_5948);
nand U10617 (N_10617,N_6369,N_6746);
nor U10618 (N_10618,N_7279,N_6927);
nor U10619 (N_10619,N_4344,N_4320);
nor U10620 (N_10620,N_5612,N_7146);
and U10621 (N_10621,N_6424,N_5292);
and U10622 (N_10622,N_7364,N_6672);
or U10623 (N_10623,N_6251,N_5983);
nand U10624 (N_10624,N_7306,N_6492);
nor U10625 (N_10625,N_7544,N_7651);
or U10626 (N_10626,N_6999,N_4164);
nor U10627 (N_10627,N_6549,N_7441);
and U10628 (N_10628,N_5022,N_5161);
and U10629 (N_10629,N_6977,N_6001);
nor U10630 (N_10630,N_4374,N_5392);
xnor U10631 (N_10631,N_6394,N_6567);
nor U10632 (N_10632,N_5442,N_7742);
nand U10633 (N_10633,N_7496,N_6688);
nor U10634 (N_10634,N_6818,N_6859);
or U10635 (N_10635,N_4736,N_6594);
nor U10636 (N_10636,N_5223,N_6365);
nor U10637 (N_10637,N_6720,N_6529);
and U10638 (N_10638,N_4237,N_4089);
nor U10639 (N_10639,N_5140,N_5807);
and U10640 (N_10640,N_5985,N_6990);
or U10641 (N_10641,N_5122,N_7832);
nor U10642 (N_10642,N_4229,N_4570);
xnor U10643 (N_10643,N_6008,N_6200);
nor U10644 (N_10644,N_7886,N_7613);
nand U10645 (N_10645,N_4079,N_6611);
and U10646 (N_10646,N_4778,N_6185);
nand U10647 (N_10647,N_4999,N_5619);
or U10648 (N_10648,N_4941,N_4945);
and U10649 (N_10649,N_6055,N_7465);
nand U10650 (N_10650,N_4453,N_5310);
nor U10651 (N_10651,N_6957,N_6154);
xnor U10652 (N_10652,N_4357,N_4976);
nor U10653 (N_10653,N_7986,N_6881);
nor U10654 (N_10654,N_4759,N_6968);
xor U10655 (N_10655,N_7034,N_4002);
nand U10656 (N_10656,N_5374,N_7102);
nor U10657 (N_10657,N_6430,N_5061);
nor U10658 (N_10658,N_6703,N_6181);
nor U10659 (N_10659,N_7330,N_4975);
nor U10660 (N_10660,N_4442,N_4665);
nor U10661 (N_10661,N_6150,N_4774);
or U10662 (N_10662,N_5154,N_6353);
nand U10663 (N_10663,N_4906,N_6236);
and U10664 (N_10664,N_5944,N_6416);
and U10665 (N_10665,N_5532,N_7516);
xor U10666 (N_10666,N_7130,N_6168);
xor U10667 (N_10667,N_4818,N_7252);
or U10668 (N_10668,N_7370,N_5436);
nand U10669 (N_10669,N_6101,N_7487);
nand U10670 (N_10670,N_6340,N_6823);
xor U10671 (N_10671,N_7994,N_7209);
or U10672 (N_10672,N_4110,N_5421);
and U10673 (N_10673,N_4339,N_5505);
and U10674 (N_10674,N_5855,N_6263);
nand U10675 (N_10675,N_7684,N_6448);
nand U10676 (N_10676,N_7303,N_5178);
nor U10677 (N_10677,N_4056,N_7721);
xor U10678 (N_10678,N_5189,N_6226);
nor U10679 (N_10679,N_5091,N_5701);
xor U10680 (N_10680,N_6478,N_7404);
and U10681 (N_10681,N_7413,N_7187);
nor U10682 (N_10682,N_4160,N_6384);
nand U10683 (N_10683,N_4758,N_7584);
nor U10684 (N_10684,N_4053,N_4605);
or U10685 (N_10685,N_7720,N_6667);
xor U10686 (N_10686,N_5010,N_6893);
nor U10687 (N_10687,N_4825,N_5136);
and U10688 (N_10688,N_7101,N_5854);
nor U10689 (N_10689,N_4193,N_7929);
nor U10690 (N_10690,N_6866,N_6039);
nand U10691 (N_10691,N_6871,N_7944);
xor U10692 (N_10692,N_6446,N_7817);
and U10693 (N_10693,N_6286,N_6093);
xor U10694 (N_10694,N_5923,N_4088);
nand U10695 (N_10695,N_5454,N_6665);
nor U10696 (N_10696,N_6040,N_6259);
or U10697 (N_10697,N_4366,N_7101);
nand U10698 (N_10698,N_6547,N_5802);
and U10699 (N_10699,N_6340,N_4533);
and U10700 (N_10700,N_5777,N_4158);
xnor U10701 (N_10701,N_4013,N_4730);
and U10702 (N_10702,N_6328,N_4703);
nor U10703 (N_10703,N_5800,N_5363);
nor U10704 (N_10704,N_6693,N_6628);
nand U10705 (N_10705,N_6744,N_5631);
or U10706 (N_10706,N_4253,N_5125);
or U10707 (N_10707,N_7720,N_5606);
nor U10708 (N_10708,N_4500,N_7389);
or U10709 (N_10709,N_4823,N_6173);
or U10710 (N_10710,N_7369,N_6835);
or U10711 (N_10711,N_5629,N_7597);
nand U10712 (N_10712,N_5581,N_7921);
xor U10713 (N_10713,N_5490,N_7833);
nand U10714 (N_10714,N_5296,N_6868);
or U10715 (N_10715,N_4507,N_6691);
nor U10716 (N_10716,N_5143,N_7896);
nand U10717 (N_10717,N_4365,N_4529);
xnor U10718 (N_10718,N_4465,N_5672);
xor U10719 (N_10719,N_6185,N_6796);
and U10720 (N_10720,N_4469,N_4889);
nor U10721 (N_10721,N_7199,N_7893);
and U10722 (N_10722,N_4539,N_7064);
or U10723 (N_10723,N_7293,N_4735);
xor U10724 (N_10724,N_6367,N_5889);
nor U10725 (N_10725,N_7017,N_4319);
nand U10726 (N_10726,N_5973,N_4309);
and U10727 (N_10727,N_4331,N_6765);
or U10728 (N_10728,N_7749,N_5241);
and U10729 (N_10729,N_7887,N_6740);
or U10730 (N_10730,N_6730,N_5048);
xor U10731 (N_10731,N_6302,N_6970);
or U10732 (N_10732,N_5959,N_6368);
nor U10733 (N_10733,N_5217,N_4085);
and U10734 (N_10734,N_4828,N_6576);
nand U10735 (N_10735,N_4643,N_6325);
or U10736 (N_10736,N_5553,N_6984);
nand U10737 (N_10737,N_5834,N_5423);
nand U10738 (N_10738,N_4904,N_7023);
xnor U10739 (N_10739,N_5757,N_6154);
or U10740 (N_10740,N_6120,N_6707);
nor U10741 (N_10741,N_4658,N_4470);
nand U10742 (N_10742,N_6835,N_4138);
nand U10743 (N_10743,N_7757,N_7565);
xnor U10744 (N_10744,N_5113,N_6860);
and U10745 (N_10745,N_7296,N_4328);
xnor U10746 (N_10746,N_4850,N_5955);
nand U10747 (N_10747,N_5254,N_5942);
and U10748 (N_10748,N_4455,N_4622);
nand U10749 (N_10749,N_6171,N_6814);
nor U10750 (N_10750,N_5716,N_6388);
nor U10751 (N_10751,N_5275,N_7026);
nor U10752 (N_10752,N_5146,N_6052);
and U10753 (N_10753,N_5820,N_5150);
and U10754 (N_10754,N_6021,N_7165);
and U10755 (N_10755,N_5202,N_6305);
nor U10756 (N_10756,N_5432,N_6073);
and U10757 (N_10757,N_5960,N_4116);
or U10758 (N_10758,N_4435,N_7807);
xor U10759 (N_10759,N_6807,N_5130);
nand U10760 (N_10760,N_7242,N_4439);
xor U10761 (N_10761,N_5455,N_7775);
nor U10762 (N_10762,N_5744,N_5419);
nor U10763 (N_10763,N_5738,N_4456);
nand U10764 (N_10764,N_5196,N_5091);
nand U10765 (N_10765,N_7417,N_4289);
or U10766 (N_10766,N_7199,N_7065);
or U10767 (N_10767,N_7421,N_6578);
nand U10768 (N_10768,N_4479,N_7510);
or U10769 (N_10769,N_6063,N_6381);
nand U10770 (N_10770,N_5150,N_4105);
nand U10771 (N_10771,N_7258,N_6043);
and U10772 (N_10772,N_7424,N_6753);
nor U10773 (N_10773,N_4225,N_4707);
and U10774 (N_10774,N_6969,N_5171);
or U10775 (N_10775,N_6962,N_7891);
nand U10776 (N_10776,N_4776,N_5838);
nand U10777 (N_10777,N_4850,N_6054);
or U10778 (N_10778,N_4763,N_4854);
and U10779 (N_10779,N_6541,N_5363);
and U10780 (N_10780,N_6320,N_6486);
xor U10781 (N_10781,N_7885,N_6642);
nand U10782 (N_10782,N_4993,N_6493);
or U10783 (N_10783,N_7913,N_6701);
nand U10784 (N_10784,N_7935,N_4032);
and U10785 (N_10785,N_7409,N_5578);
nand U10786 (N_10786,N_7680,N_5126);
nor U10787 (N_10787,N_5826,N_5569);
or U10788 (N_10788,N_7431,N_7460);
and U10789 (N_10789,N_6605,N_7055);
nor U10790 (N_10790,N_7924,N_5904);
xor U10791 (N_10791,N_7423,N_7347);
nor U10792 (N_10792,N_7147,N_7510);
or U10793 (N_10793,N_4780,N_7212);
nand U10794 (N_10794,N_7024,N_7954);
nand U10795 (N_10795,N_4121,N_4284);
nor U10796 (N_10796,N_5705,N_5502);
and U10797 (N_10797,N_7661,N_6530);
nand U10798 (N_10798,N_6498,N_4623);
nor U10799 (N_10799,N_6765,N_6783);
nand U10800 (N_10800,N_6854,N_7215);
nor U10801 (N_10801,N_6881,N_7613);
and U10802 (N_10802,N_6937,N_6354);
or U10803 (N_10803,N_5127,N_7523);
nand U10804 (N_10804,N_5677,N_6417);
and U10805 (N_10805,N_7364,N_4339);
and U10806 (N_10806,N_6024,N_4260);
nor U10807 (N_10807,N_6830,N_5492);
nor U10808 (N_10808,N_7885,N_4244);
nand U10809 (N_10809,N_6927,N_5727);
nor U10810 (N_10810,N_4248,N_6722);
nand U10811 (N_10811,N_5720,N_5690);
nand U10812 (N_10812,N_4999,N_6870);
nand U10813 (N_10813,N_5885,N_6248);
and U10814 (N_10814,N_6882,N_7919);
xnor U10815 (N_10815,N_5409,N_6108);
or U10816 (N_10816,N_7363,N_5274);
nor U10817 (N_10817,N_4343,N_6167);
or U10818 (N_10818,N_7403,N_6814);
nand U10819 (N_10819,N_6499,N_6040);
or U10820 (N_10820,N_4481,N_7301);
or U10821 (N_10821,N_6550,N_7100);
or U10822 (N_10822,N_5790,N_7624);
or U10823 (N_10823,N_7102,N_5527);
or U10824 (N_10824,N_7849,N_4632);
or U10825 (N_10825,N_6332,N_7049);
and U10826 (N_10826,N_4784,N_7913);
nor U10827 (N_10827,N_6716,N_5914);
nand U10828 (N_10828,N_5343,N_5756);
nor U10829 (N_10829,N_5758,N_5025);
nand U10830 (N_10830,N_7735,N_6131);
and U10831 (N_10831,N_6256,N_4492);
nand U10832 (N_10832,N_5138,N_4554);
nor U10833 (N_10833,N_6539,N_6689);
or U10834 (N_10834,N_5157,N_4194);
xor U10835 (N_10835,N_7452,N_7059);
or U10836 (N_10836,N_6282,N_4826);
nand U10837 (N_10837,N_5902,N_4317);
and U10838 (N_10838,N_6815,N_6510);
nand U10839 (N_10839,N_4131,N_7399);
xnor U10840 (N_10840,N_4253,N_7977);
xnor U10841 (N_10841,N_4118,N_4554);
nor U10842 (N_10842,N_4018,N_4598);
nand U10843 (N_10843,N_6702,N_6826);
xor U10844 (N_10844,N_4553,N_6454);
and U10845 (N_10845,N_5797,N_6881);
nor U10846 (N_10846,N_5659,N_7482);
nor U10847 (N_10847,N_6636,N_7705);
or U10848 (N_10848,N_5593,N_5146);
nor U10849 (N_10849,N_4185,N_6157);
xor U10850 (N_10850,N_4206,N_5359);
nor U10851 (N_10851,N_6187,N_6078);
nor U10852 (N_10852,N_4438,N_7210);
nand U10853 (N_10853,N_6012,N_7495);
and U10854 (N_10854,N_7968,N_5828);
nor U10855 (N_10855,N_4273,N_4601);
nor U10856 (N_10856,N_7347,N_6488);
nor U10857 (N_10857,N_4369,N_7467);
nor U10858 (N_10858,N_7916,N_6196);
nor U10859 (N_10859,N_7374,N_6489);
and U10860 (N_10860,N_6496,N_4795);
and U10861 (N_10861,N_7652,N_4911);
and U10862 (N_10862,N_4594,N_5131);
or U10863 (N_10863,N_6938,N_5813);
nor U10864 (N_10864,N_5698,N_7772);
nand U10865 (N_10865,N_5536,N_4986);
or U10866 (N_10866,N_5071,N_7402);
xor U10867 (N_10867,N_5592,N_5347);
and U10868 (N_10868,N_6342,N_5866);
nor U10869 (N_10869,N_4043,N_6590);
or U10870 (N_10870,N_5559,N_5252);
xnor U10871 (N_10871,N_6456,N_5915);
or U10872 (N_10872,N_4846,N_6805);
and U10873 (N_10873,N_5753,N_4891);
xor U10874 (N_10874,N_4799,N_6632);
and U10875 (N_10875,N_6185,N_5816);
and U10876 (N_10876,N_7596,N_7377);
xnor U10877 (N_10877,N_5212,N_4580);
or U10878 (N_10878,N_7927,N_5948);
nand U10879 (N_10879,N_6410,N_6252);
xor U10880 (N_10880,N_5145,N_5341);
nor U10881 (N_10881,N_7979,N_7451);
nor U10882 (N_10882,N_7397,N_4174);
xnor U10883 (N_10883,N_5546,N_6191);
xnor U10884 (N_10884,N_4806,N_7416);
nand U10885 (N_10885,N_6831,N_6124);
nand U10886 (N_10886,N_4923,N_7231);
or U10887 (N_10887,N_6999,N_6359);
and U10888 (N_10888,N_7863,N_6124);
and U10889 (N_10889,N_6831,N_4818);
nand U10890 (N_10890,N_4300,N_7206);
nor U10891 (N_10891,N_7239,N_6439);
nor U10892 (N_10892,N_5298,N_4409);
nor U10893 (N_10893,N_7748,N_5867);
or U10894 (N_10894,N_4846,N_7789);
or U10895 (N_10895,N_7305,N_5681);
or U10896 (N_10896,N_6097,N_5151);
nor U10897 (N_10897,N_6786,N_6383);
xor U10898 (N_10898,N_4463,N_7135);
nand U10899 (N_10899,N_6641,N_6267);
and U10900 (N_10900,N_7385,N_6303);
xor U10901 (N_10901,N_6318,N_7473);
and U10902 (N_10902,N_7876,N_5626);
and U10903 (N_10903,N_6014,N_4002);
nand U10904 (N_10904,N_4702,N_7491);
nor U10905 (N_10905,N_7924,N_6362);
nor U10906 (N_10906,N_7507,N_7020);
and U10907 (N_10907,N_4102,N_5872);
nor U10908 (N_10908,N_7419,N_4065);
nor U10909 (N_10909,N_6752,N_4039);
nand U10910 (N_10910,N_4244,N_5962);
and U10911 (N_10911,N_4045,N_6326);
nor U10912 (N_10912,N_4727,N_7689);
nand U10913 (N_10913,N_7343,N_6280);
xnor U10914 (N_10914,N_6076,N_4762);
and U10915 (N_10915,N_6772,N_4219);
or U10916 (N_10916,N_4371,N_6727);
nor U10917 (N_10917,N_7027,N_7682);
nor U10918 (N_10918,N_4338,N_5086);
nand U10919 (N_10919,N_6634,N_5377);
xnor U10920 (N_10920,N_6313,N_6497);
or U10921 (N_10921,N_6045,N_6573);
and U10922 (N_10922,N_4241,N_5543);
nand U10923 (N_10923,N_5758,N_6023);
nand U10924 (N_10924,N_5385,N_7307);
or U10925 (N_10925,N_5809,N_4095);
or U10926 (N_10926,N_7407,N_6397);
nand U10927 (N_10927,N_4744,N_7663);
and U10928 (N_10928,N_6345,N_7242);
nor U10929 (N_10929,N_6063,N_7673);
nor U10930 (N_10930,N_6143,N_7674);
or U10931 (N_10931,N_6850,N_6168);
or U10932 (N_10932,N_7522,N_5180);
nand U10933 (N_10933,N_4071,N_7465);
nand U10934 (N_10934,N_5105,N_6260);
nand U10935 (N_10935,N_6863,N_7721);
xnor U10936 (N_10936,N_5022,N_6509);
xnor U10937 (N_10937,N_4969,N_4557);
and U10938 (N_10938,N_5117,N_5309);
or U10939 (N_10939,N_7947,N_4676);
or U10940 (N_10940,N_5630,N_6283);
and U10941 (N_10941,N_5270,N_6477);
nor U10942 (N_10942,N_7848,N_4955);
or U10943 (N_10943,N_5880,N_5070);
nor U10944 (N_10944,N_4009,N_4524);
nor U10945 (N_10945,N_5909,N_4243);
xor U10946 (N_10946,N_5995,N_5399);
and U10947 (N_10947,N_7583,N_6239);
and U10948 (N_10948,N_6660,N_6890);
xor U10949 (N_10949,N_4705,N_4245);
or U10950 (N_10950,N_4863,N_5182);
and U10951 (N_10951,N_6316,N_6488);
and U10952 (N_10952,N_6914,N_4507);
nand U10953 (N_10953,N_6928,N_5054);
nor U10954 (N_10954,N_4451,N_4646);
and U10955 (N_10955,N_5821,N_6002);
xor U10956 (N_10956,N_6137,N_5282);
and U10957 (N_10957,N_4871,N_7591);
nor U10958 (N_10958,N_6986,N_6329);
nor U10959 (N_10959,N_7260,N_6634);
and U10960 (N_10960,N_6616,N_5134);
xnor U10961 (N_10961,N_6286,N_5505);
nand U10962 (N_10962,N_6180,N_4184);
nor U10963 (N_10963,N_4780,N_7102);
nand U10964 (N_10964,N_7372,N_6754);
nor U10965 (N_10965,N_4833,N_7666);
or U10966 (N_10966,N_4152,N_7560);
nor U10967 (N_10967,N_7132,N_5975);
nand U10968 (N_10968,N_6079,N_6626);
and U10969 (N_10969,N_5251,N_6589);
or U10970 (N_10970,N_6933,N_6289);
or U10971 (N_10971,N_6179,N_4030);
nor U10972 (N_10972,N_5471,N_6007);
xnor U10973 (N_10973,N_4745,N_5891);
nand U10974 (N_10974,N_6817,N_6336);
nor U10975 (N_10975,N_7770,N_7891);
and U10976 (N_10976,N_6269,N_6048);
or U10977 (N_10977,N_4677,N_6044);
xor U10978 (N_10978,N_7337,N_7795);
and U10979 (N_10979,N_6044,N_7486);
or U10980 (N_10980,N_6061,N_7321);
xnor U10981 (N_10981,N_6379,N_4776);
and U10982 (N_10982,N_5700,N_7786);
nor U10983 (N_10983,N_7378,N_4011);
nand U10984 (N_10984,N_6419,N_6700);
xor U10985 (N_10985,N_7248,N_6762);
and U10986 (N_10986,N_6697,N_7334);
xor U10987 (N_10987,N_7233,N_6443);
nand U10988 (N_10988,N_5656,N_7201);
or U10989 (N_10989,N_4140,N_6074);
or U10990 (N_10990,N_7458,N_6318);
or U10991 (N_10991,N_6757,N_7703);
or U10992 (N_10992,N_4223,N_6294);
and U10993 (N_10993,N_6308,N_6711);
nand U10994 (N_10994,N_5302,N_7109);
nand U10995 (N_10995,N_4928,N_5806);
or U10996 (N_10996,N_6825,N_7789);
nor U10997 (N_10997,N_4092,N_7709);
nor U10998 (N_10998,N_7386,N_6570);
or U10999 (N_10999,N_7964,N_7439);
nand U11000 (N_11000,N_5816,N_6423);
and U11001 (N_11001,N_7924,N_4984);
nor U11002 (N_11002,N_7800,N_7564);
nor U11003 (N_11003,N_5690,N_4708);
xor U11004 (N_11004,N_7346,N_5694);
nand U11005 (N_11005,N_6245,N_5396);
xnor U11006 (N_11006,N_4463,N_6471);
and U11007 (N_11007,N_4820,N_5984);
nor U11008 (N_11008,N_5221,N_6517);
nand U11009 (N_11009,N_7972,N_7071);
nor U11010 (N_11010,N_5280,N_4761);
and U11011 (N_11011,N_5228,N_7816);
or U11012 (N_11012,N_7152,N_5259);
and U11013 (N_11013,N_6140,N_5957);
and U11014 (N_11014,N_5629,N_6605);
or U11015 (N_11015,N_5494,N_6857);
nand U11016 (N_11016,N_6685,N_4003);
nand U11017 (N_11017,N_6237,N_4243);
nor U11018 (N_11018,N_7243,N_6848);
or U11019 (N_11019,N_5031,N_4167);
nand U11020 (N_11020,N_6122,N_5367);
and U11021 (N_11021,N_6521,N_4363);
nor U11022 (N_11022,N_5860,N_7635);
nor U11023 (N_11023,N_7374,N_5793);
and U11024 (N_11024,N_7180,N_7539);
and U11025 (N_11025,N_7831,N_6579);
and U11026 (N_11026,N_7532,N_4196);
nand U11027 (N_11027,N_6149,N_7605);
nor U11028 (N_11028,N_5961,N_6262);
or U11029 (N_11029,N_7780,N_7249);
xor U11030 (N_11030,N_7708,N_6448);
or U11031 (N_11031,N_7326,N_4109);
and U11032 (N_11032,N_5199,N_4048);
xnor U11033 (N_11033,N_7938,N_6368);
and U11034 (N_11034,N_6177,N_5991);
nor U11035 (N_11035,N_4095,N_6492);
xnor U11036 (N_11036,N_7184,N_4544);
or U11037 (N_11037,N_4831,N_6568);
nor U11038 (N_11038,N_7560,N_5998);
nor U11039 (N_11039,N_6381,N_6961);
nor U11040 (N_11040,N_5139,N_7346);
nor U11041 (N_11041,N_4707,N_7464);
and U11042 (N_11042,N_4557,N_5703);
nor U11043 (N_11043,N_6381,N_5731);
nand U11044 (N_11044,N_6603,N_6522);
and U11045 (N_11045,N_4312,N_5890);
xor U11046 (N_11046,N_4902,N_7677);
nand U11047 (N_11047,N_5172,N_5012);
nand U11048 (N_11048,N_7636,N_7585);
and U11049 (N_11049,N_6947,N_4627);
xor U11050 (N_11050,N_6038,N_6216);
xnor U11051 (N_11051,N_6953,N_7446);
or U11052 (N_11052,N_7012,N_4095);
or U11053 (N_11053,N_5689,N_7073);
and U11054 (N_11054,N_6721,N_5626);
xor U11055 (N_11055,N_6059,N_4458);
nor U11056 (N_11056,N_6666,N_4750);
nor U11057 (N_11057,N_4587,N_5587);
nor U11058 (N_11058,N_7688,N_7487);
xnor U11059 (N_11059,N_7486,N_4590);
and U11060 (N_11060,N_6951,N_4299);
and U11061 (N_11061,N_6079,N_6309);
and U11062 (N_11062,N_5259,N_4056);
nor U11063 (N_11063,N_7808,N_5745);
xnor U11064 (N_11064,N_7239,N_6116);
or U11065 (N_11065,N_4637,N_4738);
xor U11066 (N_11066,N_4444,N_4617);
or U11067 (N_11067,N_5436,N_4196);
nand U11068 (N_11068,N_7776,N_6985);
and U11069 (N_11069,N_5037,N_6530);
nand U11070 (N_11070,N_6174,N_4888);
nor U11071 (N_11071,N_5789,N_6344);
nand U11072 (N_11072,N_5595,N_7609);
xor U11073 (N_11073,N_4742,N_6640);
nand U11074 (N_11074,N_4737,N_6353);
and U11075 (N_11075,N_5874,N_6189);
nor U11076 (N_11076,N_4475,N_6722);
nor U11077 (N_11077,N_6315,N_4845);
nand U11078 (N_11078,N_7895,N_7507);
nand U11079 (N_11079,N_4718,N_4563);
and U11080 (N_11080,N_7184,N_5923);
nor U11081 (N_11081,N_7764,N_4056);
or U11082 (N_11082,N_5470,N_5395);
and U11083 (N_11083,N_7865,N_5959);
nand U11084 (N_11084,N_7923,N_5675);
or U11085 (N_11085,N_5657,N_7400);
or U11086 (N_11086,N_6666,N_5788);
nand U11087 (N_11087,N_4588,N_5950);
and U11088 (N_11088,N_4723,N_7077);
or U11089 (N_11089,N_4607,N_4522);
or U11090 (N_11090,N_6565,N_4021);
and U11091 (N_11091,N_5712,N_6377);
xnor U11092 (N_11092,N_7661,N_7537);
xor U11093 (N_11093,N_6246,N_7861);
and U11094 (N_11094,N_7502,N_4832);
and U11095 (N_11095,N_4641,N_5517);
or U11096 (N_11096,N_6005,N_6128);
or U11097 (N_11097,N_7882,N_4197);
nand U11098 (N_11098,N_5822,N_7397);
nand U11099 (N_11099,N_4686,N_5811);
or U11100 (N_11100,N_6224,N_5500);
nand U11101 (N_11101,N_5080,N_5085);
nor U11102 (N_11102,N_4518,N_5666);
xnor U11103 (N_11103,N_4054,N_6542);
or U11104 (N_11104,N_5038,N_5061);
or U11105 (N_11105,N_5512,N_6768);
and U11106 (N_11106,N_7588,N_4311);
or U11107 (N_11107,N_5363,N_4847);
and U11108 (N_11108,N_4314,N_7874);
nand U11109 (N_11109,N_4808,N_7476);
or U11110 (N_11110,N_7861,N_4099);
nor U11111 (N_11111,N_7766,N_6740);
nor U11112 (N_11112,N_7342,N_6049);
nand U11113 (N_11113,N_5918,N_6387);
nor U11114 (N_11114,N_7779,N_6219);
and U11115 (N_11115,N_4730,N_4564);
nor U11116 (N_11116,N_4525,N_4969);
nand U11117 (N_11117,N_4182,N_5058);
or U11118 (N_11118,N_7497,N_4498);
nand U11119 (N_11119,N_7890,N_6018);
and U11120 (N_11120,N_6744,N_6774);
nand U11121 (N_11121,N_6899,N_5783);
and U11122 (N_11122,N_5778,N_6866);
xor U11123 (N_11123,N_5618,N_4006);
and U11124 (N_11124,N_4862,N_6087);
nand U11125 (N_11125,N_4364,N_6867);
and U11126 (N_11126,N_6698,N_5020);
and U11127 (N_11127,N_5685,N_5255);
nand U11128 (N_11128,N_4759,N_6528);
nor U11129 (N_11129,N_7467,N_4304);
nor U11130 (N_11130,N_4167,N_4972);
nor U11131 (N_11131,N_5609,N_7187);
xnor U11132 (N_11132,N_4517,N_6360);
nand U11133 (N_11133,N_6550,N_5254);
nor U11134 (N_11134,N_7230,N_4990);
nor U11135 (N_11135,N_5059,N_4955);
nor U11136 (N_11136,N_7033,N_6874);
xor U11137 (N_11137,N_7260,N_6646);
xnor U11138 (N_11138,N_6978,N_4502);
nor U11139 (N_11139,N_7105,N_7594);
or U11140 (N_11140,N_7699,N_5317);
nor U11141 (N_11141,N_4125,N_5434);
or U11142 (N_11142,N_4823,N_6911);
xor U11143 (N_11143,N_5895,N_5494);
nor U11144 (N_11144,N_6102,N_6014);
nand U11145 (N_11145,N_4628,N_6627);
xnor U11146 (N_11146,N_4969,N_7169);
or U11147 (N_11147,N_4113,N_7532);
nor U11148 (N_11148,N_7240,N_7619);
nand U11149 (N_11149,N_7926,N_5535);
nor U11150 (N_11150,N_6597,N_6475);
nor U11151 (N_11151,N_6767,N_4276);
nand U11152 (N_11152,N_6324,N_7853);
or U11153 (N_11153,N_6140,N_6415);
or U11154 (N_11154,N_4009,N_6606);
nand U11155 (N_11155,N_5763,N_7855);
or U11156 (N_11156,N_6758,N_4545);
nand U11157 (N_11157,N_6420,N_7090);
or U11158 (N_11158,N_6386,N_5502);
or U11159 (N_11159,N_7434,N_5902);
nor U11160 (N_11160,N_5504,N_6069);
and U11161 (N_11161,N_7805,N_6181);
or U11162 (N_11162,N_6957,N_4158);
nand U11163 (N_11163,N_7736,N_7015);
and U11164 (N_11164,N_6995,N_6741);
or U11165 (N_11165,N_6279,N_4305);
or U11166 (N_11166,N_7027,N_7842);
nand U11167 (N_11167,N_4014,N_7270);
and U11168 (N_11168,N_7357,N_5216);
xor U11169 (N_11169,N_5421,N_4315);
and U11170 (N_11170,N_7621,N_6984);
nand U11171 (N_11171,N_5505,N_4806);
nor U11172 (N_11172,N_4108,N_6267);
xor U11173 (N_11173,N_4725,N_4326);
and U11174 (N_11174,N_6796,N_4923);
xnor U11175 (N_11175,N_7089,N_5510);
and U11176 (N_11176,N_5445,N_5319);
nand U11177 (N_11177,N_6314,N_6725);
and U11178 (N_11178,N_7198,N_5959);
nand U11179 (N_11179,N_4081,N_4227);
or U11180 (N_11180,N_4754,N_6587);
nor U11181 (N_11181,N_4134,N_6586);
xnor U11182 (N_11182,N_5190,N_7993);
and U11183 (N_11183,N_4543,N_4701);
nand U11184 (N_11184,N_5680,N_4639);
xor U11185 (N_11185,N_7872,N_5745);
nor U11186 (N_11186,N_7174,N_4734);
and U11187 (N_11187,N_6223,N_6425);
xor U11188 (N_11188,N_7241,N_7604);
nor U11189 (N_11189,N_4201,N_7662);
and U11190 (N_11190,N_4745,N_4121);
xor U11191 (N_11191,N_7695,N_4602);
and U11192 (N_11192,N_6227,N_5127);
or U11193 (N_11193,N_4246,N_4104);
xor U11194 (N_11194,N_6111,N_7116);
xnor U11195 (N_11195,N_6186,N_6763);
nand U11196 (N_11196,N_7166,N_5273);
xnor U11197 (N_11197,N_6556,N_5151);
or U11198 (N_11198,N_7015,N_7232);
or U11199 (N_11199,N_4905,N_5230);
and U11200 (N_11200,N_6009,N_4800);
nand U11201 (N_11201,N_7005,N_6837);
nor U11202 (N_11202,N_5680,N_5780);
or U11203 (N_11203,N_5365,N_4539);
or U11204 (N_11204,N_4011,N_7954);
or U11205 (N_11205,N_7341,N_6874);
nor U11206 (N_11206,N_7742,N_7696);
nand U11207 (N_11207,N_6226,N_7109);
or U11208 (N_11208,N_6942,N_6045);
nand U11209 (N_11209,N_7036,N_6064);
or U11210 (N_11210,N_4281,N_7996);
nor U11211 (N_11211,N_4835,N_7062);
and U11212 (N_11212,N_7446,N_5857);
xor U11213 (N_11213,N_4682,N_4733);
or U11214 (N_11214,N_4085,N_5196);
xnor U11215 (N_11215,N_7272,N_6263);
nor U11216 (N_11216,N_6753,N_7292);
nand U11217 (N_11217,N_4048,N_4696);
and U11218 (N_11218,N_5487,N_4984);
and U11219 (N_11219,N_7280,N_5993);
or U11220 (N_11220,N_5917,N_6712);
nand U11221 (N_11221,N_7895,N_4521);
nor U11222 (N_11222,N_4424,N_5186);
nor U11223 (N_11223,N_5774,N_7871);
or U11224 (N_11224,N_4088,N_6647);
nand U11225 (N_11225,N_6971,N_6275);
nand U11226 (N_11226,N_4327,N_6901);
xnor U11227 (N_11227,N_5464,N_6968);
and U11228 (N_11228,N_6022,N_6770);
nor U11229 (N_11229,N_6305,N_5166);
xor U11230 (N_11230,N_5238,N_6948);
and U11231 (N_11231,N_5691,N_7174);
nand U11232 (N_11232,N_4801,N_7062);
or U11233 (N_11233,N_5253,N_5273);
xor U11234 (N_11234,N_6643,N_4118);
nor U11235 (N_11235,N_5556,N_7320);
xnor U11236 (N_11236,N_4917,N_6491);
and U11237 (N_11237,N_7337,N_4031);
or U11238 (N_11238,N_5055,N_4645);
nand U11239 (N_11239,N_5609,N_7640);
xor U11240 (N_11240,N_6450,N_7226);
nand U11241 (N_11241,N_7795,N_6889);
xnor U11242 (N_11242,N_7028,N_6188);
xnor U11243 (N_11243,N_7042,N_5560);
and U11244 (N_11244,N_6842,N_7899);
or U11245 (N_11245,N_5032,N_4503);
nor U11246 (N_11246,N_7587,N_4017);
and U11247 (N_11247,N_7162,N_5647);
or U11248 (N_11248,N_5045,N_6981);
nor U11249 (N_11249,N_4122,N_4213);
nor U11250 (N_11250,N_5038,N_6801);
nand U11251 (N_11251,N_5722,N_6636);
nand U11252 (N_11252,N_6521,N_5999);
xnor U11253 (N_11253,N_4397,N_4266);
nand U11254 (N_11254,N_7380,N_7314);
nor U11255 (N_11255,N_7993,N_6418);
and U11256 (N_11256,N_5063,N_4185);
nor U11257 (N_11257,N_6060,N_5354);
or U11258 (N_11258,N_7379,N_5590);
xnor U11259 (N_11259,N_6288,N_6661);
nand U11260 (N_11260,N_5015,N_6220);
nor U11261 (N_11261,N_4327,N_5107);
or U11262 (N_11262,N_6130,N_5155);
and U11263 (N_11263,N_6318,N_4881);
or U11264 (N_11264,N_7349,N_7623);
nor U11265 (N_11265,N_7145,N_4546);
xnor U11266 (N_11266,N_4297,N_7516);
or U11267 (N_11267,N_4861,N_5231);
xor U11268 (N_11268,N_5302,N_6020);
xnor U11269 (N_11269,N_6057,N_6759);
or U11270 (N_11270,N_4996,N_5479);
nand U11271 (N_11271,N_6826,N_7158);
xor U11272 (N_11272,N_7751,N_5392);
nand U11273 (N_11273,N_6369,N_6038);
xor U11274 (N_11274,N_4488,N_7323);
and U11275 (N_11275,N_5151,N_5942);
or U11276 (N_11276,N_7896,N_4291);
or U11277 (N_11277,N_6306,N_5770);
nor U11278 (N_11278,N_4427,N_6840);
xnor U11279 (N_11279,N_7485,N_7023);
and U11280 (N_11280,N_6139,N_4018);
or U11281 (N_11281,N_7090,N_7471);
or U11282 (N_11282,N_4795,N_5195);
nor U11283 (N_11283,N_5424,N_7489);
and U11284 (N_11284,N_6075,N_4476);
or U11285 (N_11285,N_4958,N_5092);
or U11286 (N_11286,N_7571,N_6480);
nor U11287 (N_11287,N_5724,N_5596);
or U11288 (N_11288,N_7752,N_7256);
xnor U11289 (N_11289,N_5701,N_5676);
nor U11290 (N_11290,N_6300,N_4797);
nor U11291 (N_11291,N_4592,N_4463);
nor U11292 (N_11292,N_7644,N_4112);
nor U11293 (N_11293,N_6682,N_4026);
xor U11294 (N_11294,N_6645,N_6973);
or U11295 (N_11295,N_4874,N_4182);
nand U11296 (N_11296,N_4124,N_6573);
and U11297 (N_11297,N_4294,N_6897);
and U11298 (N_11298,N_4326,N_4809);
and U11299 (N_11299,N_5650,N_4745);
nor U11300 (N_11300,N_7767,N_6911);
xnor U11301 (N_11301,N_5957,N_5413);
and U11302 (N_11302,N_7643,N_6785);
nor U11303 (N_11303,N_6859,N_7575);
nand U11304 (N_11304,N_7837,N_7387);
nor U11305 (N_11305,N_7880,N_7590);
or U11306 (N_11306,N_5494,N_7672);
and U11307 (N_11307,N_4572,N_5932);
nor U11308 (N_11308,N_7456,N_4038);
or U11309 (N_11309,N_4423,N_5763);
nor U11310 (N_11310,N_5413,N_6527);
or U11311 (N_11311,N_4189,N_7589);
nand U11312 (N_11312,N_6467,N_7157);
nor U11313 (N_11313,N_4189,N_5860);
nand U11314 (N_11314,N_7123,N_4089);
or U11315 (N_11315,N_7884,N_5749);
nor U11316 (N_11316,N_4100,N_4434);
nor U11317 (N_11317,N_4334,N_6536);
and U11318 (N_11318,N_4820,N_7016);
nand U11319 (N_11319,N_6782,N_5313);
or U11320 (N_11320,N_7450,N_6985);
or U11321 (N_11321,N_5951,N_5975);
xnor U11322 (N_11322,N_4781,N_4960);
xnor U11323 (N_11323,N_4536,N_6910);
nor U11324 (N_11324,N_4627,N_6635);
and U11325 (N_11325,N_5024,N_5809);
nand U11326 (N_11326,N_6413,N_5117);
and U11327 (N_11327,N_6419,N_6437);
or U11328 (N_11328,N_7364,N_6323);
and U11329 (N_11329,N_5249,N_7655);
nor U11330 (N_11330,N_4041,N_5613);
and U11331 (N_11331,N_5272,N_7876);
nor U11332 (N_11332,N_4929,N_5357);
nor U11333 (N_11333,N_7223,N_5373);
nand U11334 (N_11334,N_4507,N_7401);
and U11335 (N_11335,N_5965,N_5674);
or U11336 (N_11336,N_6892,N_6449);
or U11337 (N_11337,N_6368,N_4393);
and U11338 (N_11338,N_7191,N_4148);
nor U11339 (N_11339,N_7688,N_7308);
nor U11340 (N_11340,N_4322,N_5054);
nor U11341 (N_11341,N_5967,N_6236);
nand U11342 (N_11342,N_4330,N_6620);
or U11343 (N_11343,N_6762,N_6315);
nand U11344 (N_11344,N_7628,N_5352);
nand U11345 (N_11345,N_4861,N_4144);
or U11346 (N_11346,N_6459,N_5552);
or U11347 (N_11347,N_5269,N_7125);
and U11348 (N_11348,N_6993,N_7109);
xnor U11349 (N_11349,N_7902,N_5531);
xor U11350 (N_11350,N_4015,N_7849);
and U11351 (N_11351,N_7717,N_5439);
nand U11352 (N_11352,N_5797,N_6179);
or U11353 (N_11353,N_4956,N_4096);
or U11354 (N_11354,N_7805,N_4740);
and U11355 (N_11355,N_6149,N_7422);
or U11356 (N_11356,N_4948,N_5633);
nand U11357 (N_11357,N_5668,N_5758);
or U11358 (N_11358,N_7039,N_7563);
and U11359 (N_11359,N_6272,N_4946);
nand U11360 (N_11360,N_4399,N_4410);
and U11361 (N_11361,N_7002,N_5909);
and U11362 (N_11362,N_5204,N_4265);
nand U11363 (N_11363,N_5042,N_5648);
xor U11364 (N_11364,N_5025,N_4544);
nor U11365 (N_11365,N_5265,N_4073);
xnor U11366 (N_11366,N_4584,N_7455);
nand U11367 (N_11367,N_4325,N_4296);
or U11368 (N_11368,N_4737,N_4725);
nand U11369 (N_11369,N_7971,N_6128);
and U11370 (N_11370,N_5366,N_6049);
nand U11371 (N_11371,N_7600,N_4787);
xor U11372 (N_11372,N_4826,N_5168);
nand U11373 (N_11373,N_7470,N_5081);
nor U11374 (N_11374,N_7485,N_5782);
nor U11375 (N_11375,N_7566,N_6890);
nand U11376 (N_11376,N_5283,N_6059);
nand U11377 (N_11377,N_4146,N_7959);
and U11378 (N_11378,N_7561,N_5465);
and U11379 (N_11379,N_7708,N_4194);
or U11380 (N_11380,N_7606,N_5400);
xor U11381 (N_11381,N_5258,N_5175);
nor U11382 (N_11382,N_4339,N_5889);
xor U11383 (N_11383,N_4767,N_6285);
or U11384 (N_11384,N_7045,N_5333);
nor U11385 (N_11385,N_7317,N_7366);
nor U11386 (N_11386,N_7771,N_7953);
xnor U11387 (N_11387,N_7722,N_4889);
or U11388 (N_11388,N_5936,N_4877);
and U11389 (N_11389,N_6541,N_4566);
nor U11390 (N_11390,N_6494,N_6270);
and U11391 (N_11391,N_6536,N_4040);
nor U11392 (N_11392,N_6906,N_5068);
nand U11393 (N_11393,N_4689,N_4738);
and U11394 (N_11394,N_4900,N_7399);
or U11395 (N_11395,N_7739,N_6703);
or U11396 (N_11396,N_7471,N_4740);
and U11397 (N_11397,N_6805,N_7290);
or U11398 (N_11398,N_5910,N_6195);
xor U11399 (N_11399,N_7387,N_5705);
and U11400 (N_11400,N_7131,N_5719);
xnor U11401 (N_11401,N_4216,N_7168);
nand U11402 (N_11402,N_4043,N_4370);
or U11403 (N_11403,N_7388,N_5402);
or U11404 (N_11404,N_6942,N_6436);
or U11405 (N_11405,N_5160,N_7030);
nand U11406 (N_11406,N_4481,N_4590);
nand U11407 (N_11407,N_7245,N_6215);
and U11408 (N_11408,N_6562,N_5163);
nor U11409 (N_11409,N_7855,N_6946);
nand U11410 (N_11410,N_5561,N_6655);
and U11411 (N_11411,N_4649,N_5651);
and U11412 (N_11412,N_7647,N_7610);
and U11413 (N_11413,N_5387,N_6094);
nand U11414 (N_11414,N_6625,N_6833);
nand U11415 (N_11415,N_5580,N_6874);
nor U11416 (N_11416,N_5085,N_6164);
nor U11417 (N_11417,N_5087,N_7746);
and U11418 (N_11418,N_6336,N_7920);
and U11419 (N_11419,N_6658,N_7230);
nand U11420 (N_11420,N_6288,N_7427);
or U11421 (N_11421,N_7794,N_6942);
xor U11422 (N_11422,N_5514,N_4423);
nand U11423 (N_11423,N_5119,N_7323);
nor U11424 (N_11424,N_5668,N_6247);
nor U11425 (N_11425,N_7387,N_7126);
and U11426 (N_11426,N_5628,N_7677);
nand U11427 (N_11427,N_7530,N_6019);
or U11428 (N_11428,N_6296,N_7002);
nand U11429 (N_11429,N_7683,N_4560);
nand U11430 (N_11430,N_7385,N_4166);
nand U11431 (N_11431,N_5671,N_6061);
or U11432 (N_11432,N_6752,N_5390);
or U11433 (N_11433,N_4973,N_5522);
nor U11434 (N_11434,N_7805,N_7752);
and U11435 (N_11435,N_4728,N_5023);
and U11436 (N_11436,N_5112,N_6301);
nand U11437 (N_11437,N_5691,N_4863);
nand U11438 (N_11438,N_4776,N_4463);
or U11439 (N_11439,N_4001,N_6983);
nor U11440 (N_11440,N_7126,N_4047);
and U11441 (N_11441,N_4313,N_5749);
nand U11442 (N_11442,N_4786,N_4561);
nor U11443 (N_11443,N_7970,N_4453);
and U11444 (N_11444,N_5761,N_5213);
and U11445 (N_11445,N_6946,N_5995);
nor U11446 (N_11446,N_5722,N_7709);
nor U11447 (N_11447,N_6523,N_4056);
nand U11448 (N_11448,N_4942,N_5807);
xnor U11449 (N_11449,N_4178,N_5050);
nand U11450 (N_11450,N_4175,N_6845);
and U11451 (N_11451,N_4494,N_6399);
nand U11452 (N_11452,N_5086,N_6357);
nand U11453 (N_11453,N_5189,N_4924);
or U11454 (N_11454,N_6467,N_4835);
or U11455 (N_11455,N_7744,N_6339);
and U11456 (N_11456,N_5729,N_7448);
nand U11457 (N_11457,N_5706,N_4111);
nor U11458 (N_11458,N_4704,N_7654);
or U11459 (N_11459,N_5372,N_5811);
nand U11460 (N_11460,N_7878,N_7144);
nand U11461 (N_11461,N_7905,N_7780);
and U11462 (N_11462,N_7651,N_7715);
or U11463 (N_11463,N_5729,N_4270);
or U11464 (N_11464,N_6284,N_4081);
xnor U11465 (N_11465,N_7837,N_6932);
and U11466 (N_11466,N_6657,N_7429);
nor U11467 (N_11467,N_5802,N_6944);
nand U11468 (N_11468,N_5606,N_7784);
and U11469 (N_11469,N_5944,N_7031);
nor U11470 (N_11470,N_7232,N_4113);
and U11471 (N_11471,N_5734,N_6319);
nand U11472 (N_11472,N_5661,N_5358);
xor U11473 (N_11473,N_4427,N_7120);
nand U11474 (N_11474,N_6472,N_6156);
and U11475 (N_11475,N_5482,N_7177);
and U11476 (N_11476,N_7560,N_7842);
or U11477 (N_11477,N_6188,N_5984);
nand U11478 (N_11478,N_7589,N_7454);
nor U11479 (N_11479,N_5624,N_6328);
or U11480 (N_11480,N_6363,N_7834);
or U11481 (N_11481,N_5382,N_5561);
and U11482 (N_11482,N_5918,N_4321);
nand U11483 (N_11483,N_7009,N_7735);
nor U11484 (N_11484,N_6398,N_5889);
nand U11485 (N_11485,N_5813,N_5301);
or U11486 (N_11486,N_6508,N_7397);
nand U11487 (N_11487,N_6279,N_5181);
or U11488 (N_11488,N_7518,N_7692);
nand U11489 (N_11489,N_6789,N_6264);
xnor U11490 (N_11490,N_7830,N_4827);
or U11491 (N_11491,N_7884,N_7477);
or U11492 (N_11492,N_4537,N_7731);
and U11493 (N_11493,N_7988,N_6957);
and U11494 (N_11494,N_4980,N_6931);
nor U11495 (N_11495,N_4155,N_4035);
and U11496 (N_11496,N_7611,N_5730);
nand U11497 (N_11497,N_6730,N_5842);
and U11498 (N_11498,N_4930,N_4397);
or U11499 (N_11499,N_6383,N_6623);
and U11500 (N_11500,N_4493,N_4748);
nor U11501 (N_11501,N_5439,N_6160);
xnor U11502 (N_11502,N_6346,N_6391);
and U11503 (N_11503,N_6583,N_6912);
nor U11504 (N_11504,N_5991,N_7128);
xnor U11505 (N_11505,N_7778,N_7594);
or U11506 (N_11506,N_6641,N_4163);
nor U11507 (N_11507,N_5933,N_7986);
and U11508 (N_11508,N_5690,N_7155);
and U11509 (N_11509,N_7644,N_5992);
or U11510 (N_11510,N_5845,N_7083);
or U11511 (N_11511,N_7543,N_4093);
nand U11512 (N_11512,N_4210,N_7842);
or U11513 (N_11513,N_7497,N_5840);
nand U11514 (N_11514,N_4249,N_5267);
or U11515 (N_11515,N_5405,N_6165);
and U11516 (N_11516,N_4847,N_4554);
nor U11517 (N_11517,N_7850,N_4492);
nand U11518 (N_11518,N_7494,N_4275);
or U11519 (N_11519,N_4387,N_7803);
and U11520 (N_11520,N_4710,N_6053);
nor U11521 (N_11521,N_4363,N_5924);
nor U11522 (N_11522,N_6696,N_7767);
nand U11523 (N_11523,N_7854,N_6429);
and U11524 (N_11524,N_6558,N_6551);
nor U11525 (N_11525,N_7763,N_6761);
nor U11526 (N_11526,N_7621,N_4676);
or U11527 (N_11527,N_4022,N_7803);
and U11528 (N_11528,N_7225,N_4142);
nor U11529 (N_11529,N_6504,N_7135);
xnor U11530 (N_11530,N_7435,N_5260);
and U11531 (N_11531,N_6846,N_7868);
or U11532 (N_11532,N_5474,N_4618);
or U11533 (N_11533,N_7427,N_7252);
nor U11534 (N_11534,N_4909,N_7270);
or U11535 (N_11535,N_4578,N_7719);
and U11536 (N_11536,N_6269,N_5098);
and U11537 (N_11537,N_4318,N_5758);
or U11538 (N_11538,N_5575,N_6827);
and U11539 (N_11539,N_7436,N_6739);
and U11540 (N_11540,N_4183,N_7790);
xnor U11541 (N_11541,N_6905,N_4644);
xnor U11542 (N_11542,N_4955,N_4065);
nor U11543 (N_11543,N_7683,N_5143);
nand U11544 (N_11544,N_4914,N_5029);
and U11545 (N_11545,N_4990,N_6348);
and U11546 (N_11546,N_7680,N_6383);
nor U11547 (N_11547,N_5177,N_6978);
nor U11548 (N_11548,N_5958,N_5918);
xor U11549 (N_11549,N_4998,N_6059);
nor U11550 (N_11550,N_6427,N_4081);
and U11551 (N_11551,N_7775,N_6386);
xnor U11552 (N_11552,N_4760,N_6604);
nand U11553 (N_11553,N_4415,N_5927);
nor U11554 (N_11554,N_7959,N_4944);
xor U11555 (N_11555,N_4821,N_6394);
and U11556 (N_11556,N_5378,N_4507);
and U11557 (N_11557,N_6120,N_7301);
or U11558 (N_11558,N_6971,N_4398);
nor U11559 (N_11559,N_6308,N_6785);
xnor U11560 (N_11560,N_7941,N_6572);
nand U11561 (N_11561,N_7668,N_5440);
or U11562 (N_11562,N_6902,N_7550);
or U11563 (N_11563,N_5341,N_6497);
nor U11564 (N_11564,N_6265,N_7309);
nor U11565 (N_11565,N_4459,N_6638);
nand U11566 (N_11566,N_5594,N_4036);
nand U11567 (N_11567,N_5150,N_5159);
nand U11568 (N_11568,N_7847,N_5747);
and U11569 (N_11569,N_7538,N_7686);
and U11570 (N_11570,N_5148,N_5957);
xnor U11571 (N_11571,N_4027,N_6038);
or U11572 (N_11572,N_4333,N_4575);
or U11573 (N_11573,N_7706,N_6216);
and U11574 (N_11574,N_6695,N_4597);
or U11575 (N_11575,N_4348,N_5304);
and U11576 (N_11576,N_5998,N_6000);
or U11577 (N_11577,N_4461,N_5896);
nor U11578 (N_11578,N_6942,N_7914);
nor U11579 (N_11579,N_4125,N_6601);
or U11580 (N_11580,N_6916,N_7988);
nand U11581 (N_11581,N_5214,N_6452);
or U11582 (N_11582,N_4134,N_4535);
nand U11583 (N_11583,N_6112,N_6281);
or U11584 (N_11584,N_7199,N_5779);
xor U11585 (N_11585,N_7458,N_4887);
nor U11586 (N_11586,N_6856,N_5258);
nor U11587 (N_11587,N_4396,N_6077);
and U11588 (N_11588,N_6623,N_7650);
nand U11589 (N_11589,N_5246,N_7790);
nor U11590 (N_11590,N_6354,N_7965);
nand U11591 (N_11591,N_7869,N_6111);
and U11592 (N_11592,N_7357,N_5803);
or U11593 (N_11593,N_6308,N_7560);
or U11594 (N_11594,N_5011,N_5199);
nand U11595 (N_11595,N_7871,N_5036);
or U11596 (N_11596,N_5111,N_5368);
or U11597 (N_11597,N_7740,N_5580);
nor U11598 (N_11598,N_5334,N_4741);
or U11599 (N_11599,N_6558,N_6689);
nor U11600 (N_11600,N_7840,N_5461);
nor U11601 (N_11601,N_6189,N_4185);
nand U11602 (N_11602,N_6984,N_7162);
or U11603 (N_11603,N_5923,N_6486);
xnor U11604 (N_11604,N_4922,N_7948);
nand U11605 (N_11605,N_7288,N_4594);
nand U11606 (N_11606,N_5362,N_6257);
nor U11607 (N_11607,N_4093,N_4276);
or U11608 (N_11608,N_6710,N_5537);
and U11609 (N_11609,N_6835,N_6778);
nor U11610 (N_11610,N_5441,N_4812);
and U11611 (N_11611,N_7438,N_5459);
or U11612 (N_11612,N_7415,N_6329);
nand U11613 (N_11613,N_7218,N_4759);
and U11614 (N_11614,N_6892,N_5360);
and U11615 (N_11615,N_4946,N_4192);
and U11616 (N_11616,N_6049,N_5326);
or U11617 (N_11617,N_4922,N_6451);
nor U11618 (N_11618,N_5733,N_7036);
nand U11619 (N_11619,N_6885,N_7274);
and U11620 (N_11620,N_6153,N_4385);
or U11621 (N_11621,N_6061,N_6237);
nand U11622 (N_11622,N_6325,N_5832);
nor U11623 (N_11623,N_6194,N_6228);
xor U11624 (N_11624,N_6238,N_6845);
or U11625 (N_11625,N_6635,N_6149);
and U11626 (N_11626,N_4316,N_4098);
nand U11627 (N_11627,N_5755,N_4290);
or U11628 (N_11628,N_5140,N_4408);
xnor U11629 (N_11629,N_5229,N_7143);
nand U11630 (N_11630,N_4496,N_5657);
nor U11631 (N_11631,N_7461,N_5420);
and U11632 (N_11632,N_7168,N_6296);
or U11633 (N_11633,N_6067,N_4357);
and U11634 (N_11634,N_7374,N_6333);
and U11635 (N_11635,N_6540,N_4275);
or U11636 (N_11636,N_4567,N_4307);
or U11637 (N_11637,N_6312,N_4113);
or U11638 (N_11638,N_7569,N_7705);
nand U11639 (N_11639,N_4235,N_5471);
and U11640 (N_11640,N_5234,N_7393);
nor U11641 (N_11641,N_7144,N_5385);
and U11642 (N_11642,N_6151,N_6601);
nor U11643 (N_11643,N_7986,N_7282);
or U11644 (N_11644,N_5864,N_6670);
xor U11645 (N_11645,N_6058,N_6188);
and U11646 (N_11646,N_5408,N_4409);
nand U11647 (N_11647,N_5179,N_7447);
xnor U11648 (N_11648,N_4335,N_7302);
and U11649 (N_11649,N_4394,N_6087);
or U11650 (N_11650,N_6441,N_6256);
and U11651 (N_11651,N_4427,N_7153);
nor U11652 (N_11652,N_7857,N_7740);
nor U11653 (N_11653,N_6137,N_4499);
and U11654 (N_11654,N_5585,N_5354);
and U11655 (N_11655,N_5181,N_7443);
xor U11656 (N_11656,N_6711,N_4965);
nor U11657 (N_11657,N_6186,N_7699);
xnor U11658 (N_11658,N_5255,N_6700);
nor U11659 (N_11659,N_7307,N_4425);
nand U11660 (N_11660,N_7248,N_6643);
nor U11661 (N_11661,N_4410,N_4113);
and U11662 (N_11662,N_4710,N_6860);
nand U11663 (N_11663,N_4664,N_6041);
nor U11664 (N_11664,N_6890,N_7199);
or U11665 (N_11665,N_7619,N_6676);
nor U11666 (N_11666,N_4514,N_6256);
or U11667 (N_11667,N_7949,N_5041);
nand U11668 (N_11668,N_4232,N_6844);
xnor U11669 (N_11669,N_5389,N_7034);
nor U11670 (N_11670,N_4947,N_6677);
and U11671 (N_11671,N_5349,N_7644);
nand U11672 (N_11672,N_6666,N_7441);
nand U11673 (N_11673,N_6693,N_5742);
nor U11674 (N_11674,N_5095,N_6907);
nor U11675 (N_11675,N_5181,N_6303);
and U11676 (N_11676,N_4259,N_7942);
and U11677 (N_11677,N_7808,N_4964);
and U11678 (N_11678,N_7393,N_4474);
nor U11679 (N_11679,N_4833,N_6315);
nand U11680 (N_11680,N_7168,N_6478);
nor U11681 (N_11681,N_6559,N_6006);
nand U11682 (N_11682,N_7109,N_6983);
and U11683 (N_11683,N_7229,N_6342);
nor U11684 (N_11684,N_4808,N_5348);
xnor U11685 (N_11685,N_5078,N_4097);
nand U11686 (N_11686,N_6654,N_4450);
nand U11687 (N_11687,N_7627,N_5007);
and U11688 (N_11688,N_6043,N_5459);
and U11689 (N_11689,N_6248,N_4988);
and U11690 (N_11690,N_5898,N_4886);
nor U11691 (N_11691,N_5237,N_5526);
nor U11692 (N_11692,N_7840,N_6454);
nor U11693 (N_11693,N_7472,N_6538);
xor U11694 (N_11694,N_6930,N_4268);
or U11695 (N_11695,N_5495,N_5350);
nand U11696 (N_11696,N_6381,N_5194);
xnor U11697 (N_11697,N_4397,N_5026);
or U11698 (N_11698,N_6926,N_7937);
or U11699 (N_11699,N_4329,N_6550);
nor U11700 (N_11700,N_6283,N_4838);
and U11701 (N_11701,N_4837,N_7290);
or U11702 (N_11702,N_7912,N_4075);
nor U11703 (N_11703,N_6454,N_7416);
and U11704 (N_11704,N_6137,N_6662);
nand U11705 (N_11705,N_6962,N_7311);
or U11706 (N_11706,N_6343,N_7364);
nor U11707 (N_11707,N_6990,N_4571);
xor U11708 (N_11708,N_7817,N_4836);
xnor U11709 (N_11709,N_4019,N_4560);
xnor U11710 (N_11710,N_6511,N_5074);
or U11711 (N_11711,N_6286,N_6283);
xnor U11712 (N_11712,N_7846,N_5252);
nand U11713 (N_11713,N_6992,N_7370);
or U11714 (N_11714,N_7914,N_5647);
or U11715 (N_11715,N_5841,N_7242);
or U11716 (N_11716,N_5669,N_7303);
and U11717 (N_11717,N_5782,N_7462);
and U11718 (N_11718,N_7578,N_4413);
and U11719 (N_11719,N_5225,N_5228);
nand U11720 (N_11720,N_6664,N_6452);
nand U11721 (N_11721,N_5195,N_5546);
nand U11722 (N_11722,N_4820,N_6180);
nor U11723 (N_11723,N_4485,N_5907);
or U11724 (N_11724,N_6677,N_5471);
and U11725 (N_11725,N_5485,N_7690);
xor U11726 (N_11726,N_6276,N_5777);
or U11727 (N_11727,N_5299,N_5051);
and U11728 (N_11728,N_5835,N_6666);
or U11729 (N_11729,N_7615,N_5274);
nand U11730 (N_11730,N_7739,N_6006);
nor U11731 (N_11731,N_6538,N_4972);
xnor U11732 (N_11732,N_4623,N_6270);
nor U11733 (N_11733,N_6411,N_4874);
or U11734 (N_11734,N_7515,N_6220);
or U11735 (N_11735,N_4595,N_7218);
nor U11736 (N_11736,N_4063,N_6996);
xnor U11737 (N_11737,N_7793,N_5631);
nand U11738 (N_11738,N_6505,N_6069);
nor U11739 (N_11739,N_6994,N_7200);
or U11740 (N_11740,N_5143,N_5419);
nand U11741 (N_11741,N_6646,N_6857);
or U11742 (N_11742,N_5300,N_4862);
and U11743 (N_11743,N_7805,N_5119);
nand U11744 (N_11744,N_6290,N_7037);
and U11745 (N_11745,N_6558,N_6670);
and U11746 (N_11746,N_5740,N_5288);
nor U11747 (N_11747,N_7942,N_4472);
nor U11748 (N_11748,N_6996,N_5387);
nand U11749 (N_11749,N_5629,N_6712);
xor U11750 (N_11750,N_6400,N_7151);
nor U11751 (N_11751,N_6496,N_4958);
or U11752 (N_11752,N_5452,N_4978);
nand U11753 (N_11753,N_4611,N_5533);
nor U11754 (N_11754,N_4991,N_6604);
nand U11755 (N_11755,N_4718,N_4862);
nor U11756 (N_11756,N_6930,N_4094);
or U11757 (N_11757,N_5500,N_6570);
nor U11758 (N_11758,N_7405,N_5209);
and U11759 (N_11759,N_6211,N_6928);
nor U11760 (N_11760,N_4172,N_5877);
xnor U11761 (N_11761,N_4905,N_5936);
or U11762 (N_11762,N_6060,N_4367);
nor U11763 (N_11763,N_5256,N_7916);
xnor U11764 (N_11764,N_7711,N_7997);
or U11765 (N_11765,N_4386,N_7607);
and U11766 (N_11766,N_7290,N_4904);
xor U11767 (N_11767,N_4722,N_7134);
nor U11768 (N_11768,N_5414,N_4079);
or U11769 (N_11769,N_6941,N_4080);
nor U11770 (N_11770,N_6113,N_4132);
or U11771 (N_11771,N_5060,N_4389);
xor U11772 (N_11772,N_7471,N_6329);
nand U11773 (N_11773,N_7309,N_7879);
nor U11774 (N_11774,N_7585,N_6419);
nand U11775 (N_11775,N_6129,N_5076);
or U11776 (N_11776,N_6360,N_5619);
nor U11777 (N_11777,N_5162,N_5104);
or U11778 (N_11778,N_7367,N_6981);
nand U11779 (N_11779,N_6883,N_5625);
nor U11780 (N_11780,N_5606,N_6606);
or U11781 (N_11781,N_4565,N_4726);
nand U11782 (N_11782,N_7967,N_6342);
and U11783 (N_11783,N_7294,N_6507);
nor U11784 (N_11784,N_6307,N_4044);
or U11785 (N_11785,N_6631,N_5828);
nor U11786 (N_11786,N_4195,N_6057);
and U11787 (N_11787,N_6677,N_7539);
nor U11788 (N_11788,N_4586,N_7667);
or U11789 (N_11789,N_6453,N_6127);
nand U11790 (N_11790,N_7352,N_5758);
nand U11791 (N_11791,N_6312,N_7539);
nor U11792 (N_11792,N_6925,N_5631);
xor U11793 (N_11793,N_5179,N_4449);
or U11794 (N_11794,N_4515,N_7394);
nor U11795 (N_11795,N_6985,N_5416);
xor U11796 (N_11796,N_7648,N_6082);
and U11797 (N_11797,N_5941,N_6930);
or U11798 (N_11798,N_6468,N_4353);
nor U11799 (N_11799,N_7410,N_4830);
and U11800 (N_11800,N_7375,N_6974);
or U11801 (N_11801,N_5044,N_4663);
nor U11802 (N_11802,N_7747,N_4049);
nor U11803 (N_11803,N_4181,N_6409);
and U11804 (N_11804,N_6312,N_6863);
nand U11805 (N_11805,N_5271,N_7009);
nor U11806 (N_11806,N_5736,N_4308);
and U11807 (N_11807,N_7720,N_6590);
and U11808 (N_11808,N_4126,N_6771);
or U11809 (N_11809,N_5354,N_5932);
nor U11810 (N_11810,N_4300,N_5864);
nor U11811 (N_11811,N_4256,N_7904);
nand U11812 (N_11812,N_6980,N_5121);
xor U11813 (N_11813,N_7782,N_7817);
and U11814 (N_11814,N_4706,N_4119);
nor U11815 (N_11815,N_5230,N_7956);
xor U11816 (N_11816,N_7526,N_4444);
xnor U11817 (N_11817,N_6097,N_5772);
or U11818 (N_11818,N_4077,N_4350);
and U11819 (N_11819,N_4209,N_4854);
or U11820 (N_11820,N_5235,N_7863);
nor U11821 (N_11821,N_4911,N_6676);
xor U11822 (N_11822,N_6083,N_6597);
nand U11823 (N_11823,N_5621,N_4479);
nand U11824 (N_11824,N_5794,N_4248);
or U11825 (N_11825,N_6373,N_7909);
xor U11826 (N_11826,N_5629,N_7656);
or U11827 (N_11827,N_4662,N_4398);
nand U11828 (N_11828,N_7510,N_7149);
and U11829 (N_11829,N_7628,N_4459);
nand U11830 (N_11830,N_4809,N_5643);
nor U11831 (N_11831,N_7741,N_5426);
nor U11832 (N_11832,N_7629,N_4806);
or U11833 (N_11833,N_6026,N_4735);
nand U11834 (N_11834,N_7441,N_4660);
and U11835 (N_11835,N_7127,N_4698);
or U11836 (N_11836,N_7432,N_4361);
nand U11837 (N_11837,N_5456,N_6289);
nand U11838 (N_11838,N_6197,N_6122);
and U11839 (N_11839,N_7646,N_4034);
nand U11840 (N_11840,N_5710,N_4451);
or U11841 (N_11841,N_5272,N_4001);
or U11842 (N_11842,N_5861,N_7793);
and U11843 (N_11843,N_7730,N_7100);
xnor U11844 (N_11844,N_7516,N_4037);
nor U11845 (N_11845,N_5112,N_7258);
nand U11846 (N_11846,N_6702,N_6242);
or U11847 (N_11847,N_5105,N_6075);
nand U11848 (N_11848,N_5668,N_4582);
and U11849 (N_11849,N_5455,N_6719);
nor U11850 (N_11850,N_4165,N_6956);
nor U11851 (N_11851,N_6962,N_7573);
xor U11852 (N_11852,N_5187,N_7155);
or U11853 (N_11853,N_7778,N_5391);
and U11854 (N_11854,N_5799,N_6506);
and U11855 (N_11855,N_7639,N_7880);
nand U11856 (N_11856,N_7210,N_5875);
nor U11857 (N_11857,N_7530,N_6902);
or U11858 (N_11858,N_4203,N_4692);
nand U11859 (N_11859,N_7240,N_5504);
nor U11860 (N_11860,N_5081,N_7812);
nand U11861 (N_11861,N_4477,N_5578);
and U11862 (N_11862,N_6313,N_5576);
nand U11863 (N_11863,N_5034,N_7826);
nor U11864 (N_11864,N_4092,N_5832);
or U11865 (N_11865,N_4581,N_4605);
and U11866 (N_11866,N_7697,N_6159);
nor U11867 (N_11867,N_6442,N_7136);
or U11868 (N_11868,N_5539,N_4484);
or U11869 (N_11869,N_4029,N_6809);
and U11870 (N_11870,N_6815,N_6073);
nor U11871 (N_11871,N_5448,N_7790);
nor U11872 (N_11872,N_4636,N_6391);
nor U11873 (N_11873,N_7145,N_6826);
or U11874 (N_11874,N_4569,N_4219);
nand U11875 (N_11875,N_6328,N_5309);
and U11876 (N_11876,N_6143,N_7937);
xor U11877 (N_11877,N_4202,N_5047);
nand U11878 (N_11878,N_6517,N_4640);
nor U11879 (N_11879,N_5162,N_5270);
nand U11880 (N_11880,N_7924,N_7248);
or U11881 (N_11881,N_4187,N_6900);
nor U11882 (N_11882,N_5928,N_7454);
or U11883 (N_11883,N_4508,N_6416);
xnor U11884 (N_11884,N_7551,N_4686);
or U11885 (N_11885,N_6620,N_4060);
nand U11886 (N_11886,N_6702,N_7525);
and U11887 (N_11887,N_6245,N_7145);
nor U11888 (N_11888,N_5820,N_6583);
or U11889 (N_11889,N_5541,N_6209);
nand U11890 (N_11890,N_6046,N_7656);
and U11891 (N_11891,N_4989,N_4998);
and U11892 (N_11892,N_4915,N_7732);
nor U11893 (N_11893,N_4372,N_7033);
and U11894 (N_11894,N_7680,N_6661);
or U11895 (N_11895,N_4512,N_5214);
or U11896 (N_11896,N_7540,N_6982);
or U11897 (N_11897,N_6326,N_7150);
nand U11898 (N_11898,N_4187,N_5947);
or U11899 (N_11899,N_5323,N_4514);
nand U11900 (N_11900,N_6390,N_6930);
and U11901 (N_11901,N_4014,N_7607);
nor U11902 (N_11902,N_6091,N_7107);
and U11903 (N_11903,N_7294,N_5821);
or U11904 (N_11904,N_7567,N_5394);
nand U11905 (N_11905,N_7774,N_7619);
and U11906 (N_11906,N_6935,N_5591);
nand U11907 (N_11907,N_6968,N_6474);
nand U11908 (N_11908,N_5114,N_6591);
and U11909 (N_11909,N_7969,N_7985);
nand U11910 (N_11910,N_6327,N_6192);
nand U11911 (N_11911,N_4107,N_7284);
nor U11912 (N_11912,N_7597,N_4786);
and U11913 (N_11913,N_5245,N_5906);
nand U11914 (N_11914,N_7532,N_5899);
nand U11915 (N_11915,N_4880,N_5761);
nor U11916 (N_11916,N_4557,N_4611);
nor U11917 (N_11917,N_7349,N_4237);
xor U11918 (N_11918,N_5161,N_7064);
nand U11919 (N_11919,N_6283,N_4349);
and U11920 (N_11920,N_4524,N_7074);
and U11921 (N_11921,N_4979,N_7973);
and U11922 (N_11922,N_5063,N_6776);
nand U11923 (N_11923,N_6131,N_4622);
nor U11924 (N_11924,N_4729,N_6776);
nand U11925 (N_11925,N_7238,N_6820);
nor U11926 (N_11926,N_6362,N_7097);
or U11927 (N_11927,N_5781,N_7659);
and U11928 (N_11928,N_4803,N_5377);
nand U11929 (N_11929,N_5956,N_7396);
nand U11930 (N_11930,N_4251,N_4628);
and U11931 (N_11931,N_4252,N_6612);
and U11932 (N_11932,N_7609,N_5984);
or U11933 (N_11933,N_4153,N_7291);
nand U11934 (N_11934,N_4387,N_6221);
and U11935 (N_11935,N_5565,N_6172);
nand U11936 (N_11936,N_4891,N_5872);
and U11937 (N_11937,N_4421,N_5310);
and U11938 (N_11938,N_5182,N_5652);
or U11939 (N_11939,N_7339,N_5366);
nor U11940 (N_11940,N_4573,N_5387);
and U11941 (N_11941,N_4333,N_6092);
or U11942 (N_11942,N_6284,N_4595);
and U11943 (N_11943,N_6448,N_4685);
or U11944 (N_11944,N_5646,N_7862);
nor U11945 (N_11945,N_4953,N_4387);
xnor U11946 (N_11946,N_6284,N_4820);
nor U11947 (N_11947,N_6656,N_6231);
or U11948 (N_11948,N_6855,N_4135);
xor U11949 (N_11949,N_4206,N_7497);
nor U11950 (N_11950,N_6579,N_7078);
nor U11951 (N_11951,N_6677,N_6808);
nand U11952 (N_11952,N_4240,N_6353);
xor U11953 (N_11953,N_5286,N_6675);
or U11954 (N_11954,N_7181,N_7510);
nor U11955 (N_11955,N_7554,N_6164);
or U11956 (N_11956,N_7094,N_5653);
or U11957 (N_11957,N_4561,N_4159);
nor U11958 (N_11958,N_4508,N_6663);
nor U11959 (N_11959,N_6157,N_7256);
or U11960 (N_11960,N_5706,N_7999);
nor U11961 (N_11961,N_4006,N_6178);
nor U11962 (N_11962,N_6059,N_5385);
nand U11963 (N_11963,N_7364,N_6803);
nand U11964 (N_11964,N_5903,N_6716);
nand U11965 (N_11965,N_6017,N_5482);
or U11966 (N_11966,N_7035,N_6112);
or U11967 (N_11967,N_7402,N_4429);
and U11968 (N_11968,N_4158,N_4992);
nor U11969 (N_11969,N_7992,N_5954);
or U11970 (N_11970,N_6196,N_7404);
or U11971 (N_11971,N_5131,N_7062);
nand U11972 (N_11972,N_7130,N_6754);
and U11973 (N_11973,N_5712,N_7946);
nor U11974 (N_11974,N_4881,N_4707);
and U11975 (N_11975,N_5310,N_6092);
nand U11976 (N_11976,N_4250,N_5460);
xor U11977 (N_11977,N_6094,N_5736);
nand U11978 (N_11978,N_4167,N_5497);
nand U11979 (N_11979,N_5185,N_6806);
nand U11980 (N_11980,N_6294,N_7273);
nand U11981 (N_11981,N_4383,N_4443);
nor U11982 (N_11982,N_6924,N_6149);
and U11983 (N_11983,N_6481,N_7685);
nor U11984 (N_11984,N_7356,N_5321);
nor U11985 (N_11985,N_4891,N_7218);
and U11986 (N_11986,N_5335,N_5179);
or U11987 (N_11987,N_7460,N_4382);
nor U11988 (N_11988,N_7169,N_6172);
and U11989 (N_11989,N_4712,N_5660);
nand U11990 (N_11990,N_6510,N_7075);
xnor U11991 (N_11991,N_5062,N_6659);
nand U11992 (N_11992,N_5054,N_6680);
nor U11993 (N_11993,N_7187,N_7112);
and U11994 (N_11994,N_5547,N_6816);
nor U11995 (N_11995,N_6360,N_7345);
nand U11996 (N_11996,N_4549,N_7597);
nand U11997 (N_11997,N_6833,N_6696);
and U11998 (N_11998,N_7776,N_4541);
nor U11999 (N_11999,N_6535,N_4392);
nor U12000 (N_12000,N_10740,N_8952);
or U12001 (N_12001,N_10393,N_8850);
nand U12002 (N_12002,N_9351,N_9222);
and U12003 (N_12003,N_8150,N_11101);
or U12004 (N_12004,N_9100,N_8123);
nand U12005 (N_12005,N_11942,N_8064);
nand U12006 (N_12006,N_9725,N_10857);
nand U12007 (N_12007,N_10410,N_8414);
nand U12008 (N_12008,N_10426,N_11756);
nor U12009 (N_12009,N_11172,N_9070);
or U12010 (N_12010,N_11194,N_8199);
nor U12011 (N_12011,N_10450,N_9611);
nor U12012 (N_12012,N_10596,N_8392);
or U12013 (N_12013,N_10974,N_11411);
nand U12014 (N_12014,N_9096,N_11285);
and U12015 (N_12015,N_11896,N_10792);
nor U12016 (N_12016,N_11080,N_9650);
nand U12017 (N_12017,N_10047,N_8760);
nand U12018 (N_12018,N_8041,N_9921);
nand U12019 (N_12019,N_10335,N_8457);
nand U12020 (N_12020,N_8489,N_10808);
nor U12021 (N_12021,N_11118,N_8055);
nand U12022 (N_12022,N_11076,N_10522);
nor U12023 (N_12023,N_11195,N_10790);
nor U12024 (N_12024,N_10435,N_10349);
nand U12025 (N_12025,N_9486,N_10846);
nand U12026 (N_12026,N_9082,N_9771);
nand U12027 (N_12027,N_10397,N_10971);
nand U12028 (N_12028,N_11584,N_10782);
nand U12029 (N_12029,N_10563,N_10616);
nor U12030 (N_12030,N_11311,N_8344);
nor U12031 (N_12031,N_11250,N_10549);
nand U12032 (N_12032,N_10281,N_9064);
nand U12033 (N_12033,N_9261,N_9020);
nand U12034 (N_12034,N_9001,N_11854);
xor U12035 (N_12035,N_10487,N_10609);
and U12036 (N_12036,N_9561,N_11853);
and U12037 (N_12037,N_11647,N_8535);
nor U12038 (N_12038,N_9981,N_9189);
nor U12039 (N_12039,N_9792,N_11639);
and U12040 (N_12040,N_10245,N_11028);
nor U12041 (N_12041,N_8555,N_11634);
and U12042 (N_12042,N_8407,N_9498);
or U12043 (N_12043,N_11061,N_11970);
xnor U12044 (N_12044,N_11774,N_11981);
and U12045 (N_12045,N_8839,N_9854);
or U12046 (N_12046,N_8808,N_8718);
nor U12047 (N_12047,N_10650,N_9426);
xor U12048 (N_12048,N_8805,N_10139);
nor U12049 (N_12049,N_9699,N_10479);
nor U12050 (N_12050,N_10380,N_9566);
nor U12051 (N_12051,N_11660,N_9316);
nor U12052 (N_12052,N_8128,N_9573);
nand U12053 (N_12053,N_9761,N_11966);
nor U12054 (N_12054,N_9909,N_9060);
and U12055 (N_12055,N_8737,N_10020);
or U12056 (N_12056,N_9799,N_8696);
nor U12057 (N_12057,N_8670,N_8481);
and U12058 (N_12058,N_8245,N_8885);
or U12059 (N_12059,N_11887,N_9801);
nor U12060 (N_12060,N_10986,N_8447);
or U12061 (N_12061,N_8558,N_11099);
nor U12062 (N_12062,N_11553,N_9037);
or U12063 (N_12063,N_8834,N_9267);
or U12064 (N_12064,N_9820,N_11054);
and U12065 (N_12065,N_9968,N_11425);
and U12066 (N_12066,N_10724,N_11294);
nor U12067 (N_12067,N_11699,N_9103);
or U12068 (N_12068,N_11763,N_9508);
or U12069 (N_12069,N_10779,N_8940);
nor U12070 (N_12070,N_11108,N_11560);
nor U12071 (N_12071,N_8334,N_9401);
and U12072 (N_12072,N_9819,N_11807);
nor U12073 (N_12073,N_11885,N_9900);
and U12074 (N_12074,N_9623,N_10990);
nand U12075 (N_12075,N_8568,N_8847);
xor U12076 (N_12076,N_9376,N_8620);
nand U12077 (N_12077,N_11579,N_9235);
or U12078 (N_12078,N_9569,N_11592);
or U12079 (N_12079,N_11295,N_11969);
nand U12080 (N_12080,N_9260,N_11765);
nand U12081 (N_12081,N_11809,N_9529);
or U12082 (N_12082,N_8849,N_11288);
nor U12083 (N_12083,N_8543,N_10844);
and U12084 (N_12084,N_10743,N_9974);
nand U12085 (N_12085,N_9145,N_9838);
and U12086 (N_12086,N_8008,N_11671);
nor U12087 (N_12087,N_10082,N_9523);
and U12088 (N_12088,N_10728,N_8956);
nand U12089 (N_12089,N_11606,N_9582);
nor U12090 (N_12090,N_8417,N_8591);
nand U12091 (N_12091,N_8275,N_11545);
nor U12092 (N_12092,N_9580,N_11060);
xor U12093 (N_12093,N_8350,N_9507);
nand U12094 (N_12094,N_10817,N_11741);
or U12095 (N_12095,N_10710,N_9294);
and U12096 (N_12096,N_10278,N_11367);
nand U12097 (N_12097,N_10761,N_9217);
or U12098 (N_12098,N_11052,N_9411);
or U12099 (N_12099,N_9285,N_11502);
nor U12100 (N_12100,N_11074,N_9199);
nor U12101 (N_12101,N_8538,N_8108);
or U12102 (N_12102,N_10361,N_9911);
and U12103 (N_12103,N_10698,N_8587);
nand U12104 (N_12104,N_8460,N_10482);
or U12105 (N_12105,N_10658,N_8459);
nand U12106 (N_12106,N_8342,N_10336);
or U12107 (N_12107,N_10227,N_11486);
nand U12108 (N_12108,N_11494,N_11743);
and U12109 (N_12109,N_11730,N_9884);
nand U12110 (N_12110,N_8794,N_10804);
nand U12111 (N_12111,N_8063,N_9436);
and U12112 (N_12112,N_8540,N_10136);
nand U12113 (N_12113,N_9214,N_9723);
nand U12114 (N_12114,N_9534,N_10237);
or U12115 (N_12115,N_10063,N_11707);
or U12116 (N_12116,N_9485,N_10443);
or U12117 (N_12117,N_11575,N_11622);
and U12118 (N_12118,N_10205,N_11492);
nand U12119 (N_12119,N_8755,N_11668);
xor U12120 (N_12120,N_9333,N_9961);
or U12121 (N_12121,N_11040,N_10294);
or U12122 (N_12122,N_11376,N_10832);
nor U12123 (N_12123,N_8405,N_10198);
and U12124 (N_12124,N_10555,N_11605);
or U12125 (N_12125,N_8118,N_9137);
nor U12126 (N_12126,N_11064,N_8933);
nand U12127 (N_12127,N_11534,N_11443);
nor U12128 (N_12128,N_9581,N_10216);
nor U12129 (N_12129,N_9949,N_11006);
and U12130 (N_12130,N_11163,N_9129);
or U12131 (N_12131,N_11362,N_8689);
xnor U12132 (N_12132,N_8131,N_8375);
nand U12133 (N_12133,N_8018,N_9750);
nand U12134 (N_12134,N_8564,N_8364);
or U12135 (N_12135,N_9034,N_10599);
xor U12136 (N_12136,N_10718,N_10920);
nand U12137 (N_12137,N_9047,N_8906);
or U12138 (N_12138,N_8341,N_10876);
nor U12139 (N_12139,N_9039,N_11428);
nand U12140 (N_12140,N_11351,N_8362);
or U12141 (N_12141,N_11547,N_9991);
or U12142 (N_12142,N_8652,N_10392);
or U12143 (N_12143,N_10271,N_8817);
and U12144 (N_12144,N_11232,N_11812);
or U12145 (N_12145,N_8778,N_8090);
and U12146 (N_12146,N_10352,N_11273);
nand U12147 (N_12147,N_9857,N_9067);
or U12148 (N_12148,N_11281,N_8410);
xor U12149 (N_12149,N_9334,N_8099);
or U12150 (N_12150,N_8918,N_10636);
and U12151 (N_12151,N_9906,N_10733);
nand U12152 (N_12152,N_9538,N_11350);
or U12153 (N_12153,N_10663,N_9410);
or U12154 (N_12154,N_8235,N_8458);
nor U12155 (N_12155,N_9239,N_11435);
or U12156 (N_12156,N_9065,N_11434);
xor U12157 (N_12157,N_8867,N_8901);
nand U12158 (N_12158,N_11858,N_9447);
or U12159 (N_12159,N_11037,N_9172);
and U12160 (N_12160,N_10333,N_10454);
or U12161 (N_12161,N_10535,N_8265);
nor U12162 (N_12162,N_8989,N_11272);
or U12163 (N_12163,N_9694,N_9841);
xnor U12164 (N_12164,N_10356,N_10096);
or U12165 (N_12165,N_9689,N_9099);
nor U12166 (N_12166,N_11026,N_9632);
nor U12167 (N_12167,N_9703,N_9338);
nand U12168 (N_12168,N_11215,N_8355);
nand U12169 (N_12169,N_9955,N_10912);
nor U12170 (N_12170,N_8452,N_9008);
nand U12171 (N_12171,N_9437,N_9228);
nor U12172 (N_12172,N_10843,N_9717);
and U12173 (N_12173,N_9640,N_9871);
nor U12174 (N_12174,N_8425,N_8957);
or U12175 (N_12175,N_10554,N_10418);
xor U12176 (N_12176,N_10931,N_9361);
xnor U12177 (N_12177,N_8946,N_10727);
nand U12178 (N_12178,N_11017,N_10452);
nand U12179 (N_12179,N_10326,N_10993);
nor U12180 (N_12180,N_10131,N_8557);
or U12181 (N_12181,N_11649,N_8043);
xnor U12182 (N_12182,N_8647,N_8511);
nor U12183 (N_12183,N_10010,N_11354);
nand U12184 (N_12184,N_10716,N_8667);
nor U12185 (N_12185,N_9688,N_8263);
or U12186 (N_12186,N_10623,N_9933);
nor U12187 (N_12187,N_9598,N_9300);
or U12188 (N_12188,N_11828,N_11466);
xnor U12189 (N_12189,N_8403,N_10648);
xnor U12190 (N_12190,N_10826,N_11246);
or U12191 (N_12191,N_9387,N_10343);
nor U12192 (N_12192,N_8967,N_11818);
and U12193 (N_12193,N_11777,N_8610);
nor U12194 (N_12194,N_8488,N_8152);
and U12195 (N_12195,N_9083,N_10477);
or U12196 (N_12196,N_9992,N_11531);
nand U12197 (N_12197,N_10107,N_9501);
nand U12198 (N_12198,N_9506,N_10634);
nor U12199 (N_12199,N_9557,N_9310);
xor U12200 (N_12200,N_9004,N_10962);
nand U12201 (N_12201,N_10066,N_11972);
or U12202 (N_12202,N_11721,N_9674);
nor U12203 (N_12203,N_8175,N_8005);
nand U12204 (N_12204,N_9031,N_9389);
and U12205 (N_12205,N_8714,N_8735);
or U12206 (N_12206,N_8859,N_9420);
and U12207 (N_12207,N_9280,N_9676);
or U12208 (N_12208,N_10958,N_8366);
nand U12209 (N_12209,N_11100,N_9385);
and U12210 (N_12210,N_8765,N_10263);
nand U12211 (N_12211,N_8868,N_10647);
and U12212 (N_12212,N_10488,N_10945);
and U12213 (N_12213,N_11779,N_9864);
and U12214 (N_12214,N_9328,N_10592);
or U12215 (N_12215,N_8923,N_9291);
nor U12216 (N_12216,N_9954,N_10468);
nor U12217 (N_12217,N_8462,N_8177);
or U12218 (N_12218,N_8479,N_8533);
and U12219 (N_12219,N_9363,N_8571);
xor U12220 (N_12220,N_8603,N_8130);
and U12221 (N_12221,N_11033,N_10436);
nor U12222 (N_12222,N_9358,N_8013);
or U12223 (N_12223,N_9038,N_10784);
xnor U12224 (N_12224,N_11306,N_9619);
and U12225 (N_12225,N_8575,N_9883);
nand U12226 (N_12226,N_8451,N_11129);
and U12227 (N_12227,N_11365,N_11451);
and U12228 (N_12228,N_8276,N_11624);
nand U12229 (N_12229,N_10508,N_9695);
or U12230 (N_12230,N_10369,N_8733);
nand U12231 (N_12231,N_8328,N_9434);
or U12232 (N_12232,N_9600,N_10785);
nor U12233 (N_12233,N_8665,N_9033);
nor U12234 (N_12234,N_10607,N_9938);
nand U12235 (N_12235,N_11136,N_10730);
and U12236 (N_12236,N_9740,N_9169);
nand U12237 (N_12237,N_8640,N_8633);
and U12238 (N_12238,N_8030,N_8544);
or U12239 (N_12239,N_11906,N_11817);
or U12240 (N_12240,N_11319,N_9517);
and U12241 (N_12241,N_9692,N_11926);
nand U12242 (N_12242,N_8779,N_11923);
nor U12243 (N_12243,N_10988,N_11918);
nand U12244 (N_12244,N_11197,N_10519);
nor U12245 (N_12245,N_8856,N_11968);
and U12246 (N_12246,N_9299,N_10935);
and U12247 (N_12247,N_9945,N_11401);
or U12248 (N_12248,N_11039,N_11702);
and U12249 (N_12249,N_11866,N_10168);
or U12250 (N_12250,N_8329,N_11338);
and U12251 (N_12251,N_8047,N_9835);
nand U12252 (N_12252,N_10654,N_8502);
or U12253 (N_12253,N_10871,N_10032);
or U12254 (N_12254,N_8581,N_8877);
xor U12255 (N_12255,N_10880,N_9112);
nand U12256 (N_12256,N_10702,N_10191);
and U12257 (N_12257,N_8282,N_9629);
xor U12258 (N_12258,N_10328,N_11089);
and U12259 (N_12259,N_8307,N_8529);
or U12260 (N_12260,N_11192,N_11835);
or U12261 (N_12261,N_9605,N_10464);
and U12262 (N_12262,N_9175,N_9312);
nor U12263 (N_12263,N_10241,N_11978);
or U12264 (N_12264,N_11045,N_8438);
and U12265 (N_12265,N_8035,N_9532);
nand U12266 (N_12266,N_11175,N_11432);
nor U12267 (N_12267,N_8060,N_9014);
or U12268 (N_12268,N_8306,N_10850);
or U12269 (N_12269,N_10415,N_9638);
nand U12270 (N_12270,N_9758,N_9276);
nor U12271 (N_12271,N_8728,N_8873);
and U12272 (N_12272,N_9832,N_8322);
nand U12273 (N_12273,N_8872,N_8209);
and U12274 (N_12274,N_11751,N_10174);
nand U12275 (N_12275,N_11188,N_9610);
nor U12276 (N_12276,N_8052,N_8139);
or U12277 (N_12277,N_9324,N_8632);
and U12278 (N_12278,N_8394,N_11859);
and U12279 (N_12279,N_8297,N_9726);
nor U12280 (N_12280,N_11395,N_11985);
nor U12281 (N_12281,N_10902,N_11317);
or U12282 (N_12282,N_10422,N_8596);
nor U12283 (N_12283,N_9322,N_9466);
xnor U12284 (N_12284,N_11568,N_10573);
nand U12285 (N_12285,N_11944,N_10089);
and U12286 (N_12286,N_8019,N_8819);
nand U12287 (N_12287,N_8323,N_11482);
or U12288 (N_12288,N_10048,N_10715);
nor U12289 (N_12289,N_9062,N_11307);
and U12290 (N_12290,N_8113,N_11726);
nand U12291 (N_12291,N_9348,N_8220);
nand U12292 (N_12292,N_8091,N_11417);
nand U12293 (N_12293,N_10805,N_11599);
nor U12294 (N_12294,N_8774,N_11056);
and U12295 (N_12295,N_10806,N_9525);
nor U12296 (N_12296,N_11361,N_11766);
or U12297 (N_12297,N_8864,N_9236);
xor U12298 (N_12298,N_11352,N_10219);
and U12299 (N_12299,N_11007,N_11030);
nor U12300 (N_12300,N_11947,N_10346);
nor U12301 (N_12301,N_8356,N_10540);
nor U12302 (N_12302,N_10949,N_8697);
nor U12303 (N_12303,N_11032,N_9547);
xor U12304 (N_12304,N_9412,N_11051);
or U12305 (N_12305,N_10695,N_11416);
and U12306 (N_12306,N_11328,N_11041);
nand U12307 (N_12307,N_9647,N_11924);
or U12308 (N_12308,N_8663,N_9986);
and U12309 (N_12309,N_8908,N_9318);
xor U12310 (N_12310,N_10025,N_11528);
and U12311 (N_12311,N_8509,N_9844);
or U12312 (N_12312,N_11468,N_10802);
nand U12313 (N_12313,N_11050,N_11607);
and U12314 (N_12314,N_11834,N_8699);
or U12315 (N_12315,N_10652,N_10918);
nand U12316 (N_12316,N_9077,N_11196);
nor U12317 (N_12317,N_11655,N_8734);
nand U12318 (N_12318,N_9029,N_11217);
nor U12319 (N_12319,N_8766,N_11864);
and U12320 (N_12320,N_9427,N_9802);
and U12321 (N_12321,N_8319,N_8507);
nor U12322 (N_12322,N_11683,N_10156);
xnor U12323 (N_12323,N_10167,N_10079);
xnor U12324 (N_12324,N_9521,N_8333);
nand U12325 (N_12325,N_8752,N_11912);
nand U12326 (N_12326,N_11474,N_9452);
nor U12327 (N_12327,N_10366,N_10123);
and U12328 (N_12328,N_9831,N_8751);
xor U12329 (N_12329,N_9862,N_9646);
nand U12330 (N_12330,N_10858,N_11692);
or U12331 (N_12331,N_9621,N_8324);
xor U12332 (N_12332,N_8384,N_8268);
nand U12333 (N_12333,N_9978,N_8609);
nand U12334 (N_12334,N_8241,N_9293);
and U12335 (N_12335,N_8830,N_11857);
nor U12336 (N_12336,N_11018,N_10372);
nand U12337 (N_12337,N_11375,N_11705);
nand U12338 (N_12338,N_9548,N_10385);
nor U12339 (N_12339,N_9362,N_8916);
and U12340 (N_12340,N_8659,N_9115);
or U12341 (N_12341,N_10196,N_8694);
or U12342 (N_12342,N_11934,N_10713);
and U12343 (N_12343,N_10105,N_8926);
nor U12344 (N_12344,N_9317,N_9249);
nand U12345 (N_12345,N_10316,N_11020);
nor U12346 (N_12346,N_10524,N_9359);
or U12347 (N_12347,N_8441,N_8695);
or U12348 (N_12348,N_9141,N_8784);
nand U12349 (N_12349,N_11404,N_9118);
and U12350 (N_12350,N_11300,N_8812);
nor U12351 (N_12351,N_8327,N_11764);
and U12352 (N_12352,N_9794,N_8953);
and U12353 (N_12353,N_9846,N_9965);
or U12354 (N_12354,N_10255,N_10407);
or U12355 (N_12355,N_11685,N_10905);
and U12356 (N_12356,N_9630,N_10217);
nor U12357 (N_12357,N_10491,N_8829);
xor U12358 (N_12358,N_11405,N_10190);
nand U12359 (N_12359,N_8683,N_8016);
xnor U12360 (N_12360,N_11590,N_10224);
nand U12361 (N_12361,N_11327,N_9618);
nand U12362 (N_12362,N_8339,N_10117);
nor U12363 (N_12363,N_8146,N_9715);
or U12364 (N_12364,N_11057,N_9952);
or U12365 (N_12365,N_8051,N_11048);
or U12366 (N_12366,N_10019,N_10666);
nand U12367 (N_12367,N_10906,N_11304);
and U12368 (N_12368,N_8790,N_8869);
or U12369 (N_12369,N_10788,N_9360);
nor U12370 (N_12370,N_11641,N_11626);
nand U12371 (N_12371,N_9275,N_9057);
nor U12372 (N_12372,N_9539,N_10406);
nand U12373 (N_12373,N_11868,N_9815);
or U12374 (N_12374,N_9413,N_9421);
nand U12375 (N_12375,N_10513,N_9795);
and U12376 (N_12376,N_9927,N_8803);
xnor U12377 (N_12377,N_8379,N_10864);
or U12378 (N_12378,N_9603,N_11455);
or U12379 (N_12379,N_9576,N_9828);
nor U12380 (N_12380,N_11359,N_11990);
nor U12381 (N_12381,N_8731,N_10100);
or U12382 (N_12382,N_11959,N_10431);
or U12383 (N_12383,N_10753,N_11261);
or U12384 (N_12384,N_11380,N_8296);
nand U12385 (N_12385,N_9350,N_8523);
or U12386 (N_12386,N_11625,N_11044);
nand U12387 (N_12387,N_8022,N_11187);
or U12388 (N_12388,N_8082,N_9139);
nor U12389 (N_12389,N_8622,N_10894);
nor U12390 (N_12390,N_11090,N_11378);
or U12391 (N_12391,N_9661,N_10417);
or U12392 (N_12392,N_8257,N_9036);
nand U12393 (N_12393,N_9469,N_8625);
nand U12394 (N_12394,N_10615,N_10296);
or U12395 (N_12395,N_9549,N_10595);
nand U12396 (N_12396,N_8684,N_8227);
nor U12397 (N_12397,N_10106,N_9399);
or U12398 (N_12398,N_10757,N_9306);
nand U12399 (N_12399,N_11177,N_9069);
nor U12400 (N_12400,N_11711,N_9969);
nand U12401 (N_12401,N_9806,N_10505);
and U12402 (N_12402,N_8531,N_8589);
and U12403 (N_12403,N_11648,N_9853);
nand U12404 (N_12404,N_8127,N_10489);
nand U12405 (N_12405,N_11189,N_9781);
nor U12406 (N_12406,N_11672,N_9474);
or U12407 (N_12407,N_10357,N_8888);
nor U12408 (N_12408,N_10474,N_11900);
nor U12409 (N_12409,N_10341,N_10548);
nand U12410 (N_12410,N_8773,N_9205);
or U12411 (N_12411,N_9196,N_8896);
nand U12412 (N_12412,N_9754,N_11308);
or U12413 (N_12413,N_10176,N_10527);
nand U12414 (N_12414,N_11004,N_8229);
nand U12415 (N_12415,N_11022,N_10500);
or U12416 (N_12416,N_10583,N_10432);
nor U12417 (N_12417,N_9425,N_8965);
and U12418 (N_12418,N_10360,N_11305);
and U12419 (N_12419,N_8092,N_9970);
nor U12420 (N_12420,N_8308,N_11496);
nand U12421 (N_12421,N_8086,N_11752);
or U12422 (N_12422,N_8722,N_11754);
and U12423 (N_12423,N_10498,N_8184);
nand U12424 (N_12424,N_10109,N_8865);
or U12425 (N_12425,N_8250,N_10321);
nand U12426 (N_12426,N_8806,N_9929);
nand U12427 (N_12427,N_11550,N_10381);
nand U12428 (N_12428,N_10893,N_11334);
and U12429 (N_12429,N_8505,N_8929);
or U12430 (N_12430,N_11077,N_10083);
nor U12431 (N_12431,N_11190,N_9868);
nand U12432 (N_12432,N_8206,N_11469);
nand U12433 (N_12433,N_11513,N_8706);
nor U12434 (N_12434,N_10310,N_9114);
nor U12435 (N_12435,N_9564,N_9010);
nor U12436 (N_12436,N_8182,N_8491);
nand U12437 (N_12437,N_9084,N_9966);
nand U12438 (N_12438,N_8170,N_11613);
and U12439 (N_12439,N_8454,N_10175);
xnor U12440 (N_12440,N_11512,N_10374);
or U12441 (N_12441,N_10531,N_8948);
nand U12442 (N_12442,N_8517,N_9049);
nor U12443 (N_12443,N_9246,N_8247);
nor U12444 (N_12444,N_11214,N_9651);
nand U12445 (N_12445,N_10424,N_11949);
nand U12446 (N_12446,N_9476,N_9032);
or U12447 (N_12447,N_11204,N_11587);
and U12448 (N_12448,N_10445,N_8133);
nand U12449 (N_12449,N_10632,N_11916);
nor U12450 (N_12450,N_9918,N_8293);
or U12451 (N_12451,N_9023,N_11663);
nor U12452 (N_12452,N_8653,N_8391);
or U12453 (N_12453,N_10157,N_9989);
xor U12454 (N_12454,N_9304,N_11958);
or U12455 (N_12455,N_9928,N_9659);
nand U12456 (N_12456,N_10585,N_8312);
or U12457 (N_12457,N_11563,N_9415);
or U12458 (N_12458,N_8053,N_9985);
nor U12459 (N_12459,N_8661,N_8370);
nor U12460 (N_12460,N_8676,N_11497);
xnor U12461 (N_12461,N_8708,N_8823);
nand U12462 (N_12462,N_8927,N_8471);
nand U12463 (N_12463,N_11637,N_11446);
nand U12464 (N_12464,N_9731,N_9719);
nor U12465 (N_12465,N_10171,N_10597);
nor U12466 (N_12466,N_10758,N_9074);
nand U12467 (N_12467,N_8105,N_11744);
or U12468 (N_12468,N_11248,N_11687);
nand U12469 (N_12469,N_11166,N_8122);
or U12470 (N_12470,N_11005,N_11874);
or U12471 (N_12471,N_11369,N_10539);
and U12472 (N_12472,N_8725,N_9151);
nor U12473 (N_12473,N_10518,N_11768);
nand U12474 (N_12474,N_11238,N_9814);
nor U12475 (N_12475,N_8607,N_9546);
or U12476 (N_12476,N_8613,N_8892);
and U12477 (N_12477,N_9833,N_11453);
and U12478 (N_12478,N_10103,N_9156);
nor U12479 (N_12479,N_11340,N_11666);
or U12480 (N_12480,N_11010,N_10095);
nand U12481 (N_12481,N_9988,N_10701);
and U12482 (N_12482,N_9994,N_10319);
and U12483 (N_12483,N_8239,N_10226);
or U12484 (N_12484,N_9336,N_9011);
nand U12485 (N_12485,N_9655,N_9824);
nor U12486 (N_12486,N_10252,N_9493);
xnor U12487 (N_12487,N_8255,N_11895);
or U12488 (N_12488,N_11123,N_11385);
nand U12489 (N_12489,N_9256,N_8443);
nor U12490 (N_12490,N_8693,N_10969);
or U12491 (N_12491,N_8782,N_8000);
nand U12492 (N_12492,N_10645,N_11806);
or U12493 (N_12493,N_9191,N_10127);
and U12494 (N_12494,N_10760,N_10188);
nand U12495 (N_12495,N_9673,N_9471);
nand U12496 (N_12496,N_10789,N_11292);
nor U12497 (N_12497,N_10831,N_10441);
or U12498 (N_12498,N_9686,N_8945);
or U12499 (N_12499,N_10193,N_10416);
nor U12500 (N_12500,N_9181,N_9553);
and U12501 (N_12501,N_9459,N_9662);
xor U12502 (N_12502,N_9917,N_11597);
nand U12503 (N_12503,N_11794,N_11391);
or U12504 (N_12504,N_8467,N_9908);
or U12505 (N_12505,N_11387,N_10960);
or U12506 (N_12506,N_8813,N_8848);
or U12507 (N_12507,N_11266,N_8506);
and U12508 (N_12508,N_11329,N_10017);
or U12509 (N_12509,N_8814,N_9912);
nor U12510 (N_12510,N_8033,N_9109);
nand U12511 (N_12511,N_10249,N_8903);
nand U12512 (N_12512,N_8756,N_8820);
nand U12513 (N_12513,N_10903,N_8213);
and U12514 (N_12514,N_8497,N_8567);
nor U12515 (N_12515,N_8550,N_10447);
nand U12516 (N_12516,N_11619,N_10244);
and U12517 (N_12517,N_10633,N_10794);
nand U12518 (N_12518,N_9024,N_10504);
xor U12519 (N_12519,N_11820,N_11580);
or U12520 (N_12520,N_10959,N_11221);
nand U12521 (N_12521,N_10126,N_9608);
nand U12522 (N_12522,N_9948,N_11669);
or U12523 (N_12523,N_8899,N_9266);
and U12524 (N_12524,N_10869,N_9448);
and U12525 (N_12525,N_10957,N_11686);
or U12526 (N_12526,N_9158,N_8202);
and U12527 (N_12527,N_8346,N_8729);
nand U12528 (N_12528,N_10815,N_10150);
or U12529 (N_12529,N_11952,N_10622);
nand U12530 (N_12530,N_10394,N_9536);
or U12531 (N_12531,N_10284,N_11254);
or U12532 (N_12532,N_10460,N_9424);
xor U12533 (N_12533,N_11249,N_8576);
or U12534 (N_12534,N_9737,N_8891);
nor U12535 (N_12535,N_10617,N_8741);
nand U12536 (N_12536,N_10384,N_10642);
or U12537 (N_12537,N_11802,N_9735);
nand U12538 (N_12538,N_9394,N_10863);
nor U12539 (N_12539,N_9690,N_9777);
nor U12540 (N_12540,N_9542,N_8107);
or U12541 (N_12541,N_11742,N_11128);
xor U12542 (N_12542,N_10301,N_9110);
or U12543 (N_12543,N_9105,N_10342);
or U12544 (N_12544,N_10532,N_10865);
or U12545 (N_12545,N_9453,N_11991);
nand U12546 (N_12546,N_9013,N_8993);
xnor U12547 (N_12547,N_8310,N_8191);
nor U12548 (N_12548,N_11415,N_10625);
nor U12549 (N_12549,N_8709,N_10981);
or U12550 (N_12550,N_11816,N_9850);
and U12551 (N_12551,N_10911,N_9937);
or U12552 (N_12552,N_10183,N_11903);
xnor U12553 (N_12553,N_10391,N_8915);
and U12554 (N_12554,N_11481,N_11680);
nand U12555 (N_12555,N_11551,N_10218);
xnor U12556 (N_12556,N_9007,N_11348);
xor U12557 (N_12557,N_10013,N_11739);
nor U12558 (N_12558,N_11475,N_8330);
and U12559 (N_12559,N_10472,N_10781);
and U12560 (N_12560,N_10449,N_10292);
nand U12561 (N_12561,N_9873,N_11602);
or U12562 (N_12562,N_8998,N_8588);
or U12563 (N_12563,N_9418,N_8500);
nor U12564 (N_12564,N_9840,N_11325);
xnor U12565 (N_12565,N_8583,N_11141);
nor U12566 (N_12566,N_8846,N_9441);
or U12567 (N_12567,N_8955,N_9356);
or U12568 (N_12568,N_11398,N_9681);
xnor U12569 (N_12569,N_11784,N_10890);
and U12570 (N_12570,N_9787,N_11220);
nor U12571 (N_12571,N_9229,N_9620);
or U12572 (N_12572,N_10386,N_11091);
or U12573 (N_12573,N_9430,N_9417);
and U12574 (N_12574,N_11986,N_11654);
xor U12575 (N_12575,N_9073,N_9046);
nand U12576 (N_12576,N_11257,N_10809);
nor U12577 (N_12577,N_9575,N_8148);
nor U12578 (N_12578,N_9821,N_11289);
or U12579 (N_12579,N_9003,N_11526);
nor U12580 (N_12580,N_9583,N_11268);
nor U12581 (N_12581,N_8793,N_8377);
and U12582 (N_12582,N_9219,N_10128);
nor U12583 (N_12583,N_10068,N_9633);
xor U12584 (N_12584,N_8802,N_11333);
and U12585 (N_12585,N_9307,N_10348);
or U12586 (N_12586,N_11012,N_9563);
nor U12587 (N_12587,N_11132,N_8142);
or U12588 (N_12588,N_9930,N_11047);
nand U12589 (N_12589,N_9785,N_9473);
or U12590 (N_12590,N_10172,N_10603);
nand U12591 (N_12591,N_10347,N_10521);
nand U12592 (N_12592,N_10051,N_11775);
nor U12593 (N_12593,N_9058,N_8553);
or U12594 (N_12594,N_8014,N_8058);
and U12595 (N_12595,N_8103,N_9371);
nor U12596 (N_12596,N_9179,N_10315);
and U12597 (N_12597,N_11945,N_10529);
nand U12598 (N_12598,N_11447,N_10938);
nor U12599 (N_12599,N_8548,N_10242);
and U12600 (N_12600,N_10201,N_9272);
or U12601 (N_12601,N_8599,N_8186);
or U12602 (N_12602,N_9535,N_11689);
nand U12603 (N_12603,N_8851,N_8389);
and U12604 (N_12604,N_9054,N_8455);
nand U12605 (N_12605,N_11559,N_10236);
xnor U12606 (N_12606,N_9130,N_8298);
nand U12607 (N_12607,N_11558,N_8449);
xor U12608 (N_12608,N_11245,N_8145);
nand U12609 (N_12609,N_8961,N_11718);
or U12610 (N_12610,N_9388,N_8114);
and U12611 (N_12611,N_10985,N_8338);
and U12612 (N_12612,N_8563,N_11140);
nor U12613 (N_12613,N_10009,N_10362);
nor U12614 (N_12614,N_9419,N_10414);
nand U12615 (N_12615,N_11600,N_11879);
nand U12616 (N_12616,N_8619,N_10552);
nor U12617 (N_12617,N_11727,N_10024);
or U12618 (N_12618,N_11734,N_11500);
and U12619 (N_12619,N_8870,N_8763);
nand U12620 (N_12620,N_8972,N_11384);
and U12621 (N_12621,N_8036,N_8566);
xor U12622 (N_12622,N_11423,N_10948);
and U12623 (N_12623,N_10163,N_11235);
nor U12624 (N_12624,N_9045,N_8413);
and U12625 (N_12625,N_11510,N_11104);
and U12626 (N_12626,N_9072,N_8504);
nor U12627 (N_12627,N_8277,N_10114);
nand U12628 (N_12628,N_10575,N_8866);
or U12629 (N_12629,N_9198,N_8963);
or U12630 (N_12630,N_10057,N_10641);
nor U12631 (N_12631,N_11429,N_9248);
nand U12632 (N_12632,N_9939,N_10104);
or U12633 (N_12633,N_8821,N_11612);
nand U12634 (N_12634,N_10638,N_8197);
or U12635 (N_12635,N_9170,N_10533);
or U12636 (N_12636,N_9377,N_9347);
nand U12637 (N_12637,N_9422,N_10134);
and U12638 (N_12638,N_10312,N_8478);
nor U12639 (N_12639,N_10485,N_10991);
and U12640 (N_12640,N_11899,N_11865);
or U12641 (N_12641,N_11658,N_9936);
nand U12642 (N_12642,N_8490,N_11997);
and U12643 (N_12643,N_8210,N_9984);
nand U12644 (N_12644,N_8875,N_8421);
or U12645 (N_12645,N_9019,N_10769);
nand U12646 (N_12646,N_8801,N_9606);
or U12647 (N_12647,N_9216,N_11603);
and U12648 (N_12648,N_8260,N_10928);
nor U12649 (N_12649,N_11083,N_8840);
nor U12650 (N_12650,N_10665,N_11346);
nand U12651 (N_12651,N_9764,N_10182);
nand U12652 (N_12652,N_11407,N_11016);
or U12653 (N_12653,N_10455,N_10584);
nand U12654 (N_12654,N_8109,N_11540);
nor U12655 (N_12655,N_8201,N_9382);
nand U12656 (N_12656,N_10137,N_9218);
and U12657 (N_12657,N_8404,N_8302);
nor U12658 (N_12658,N_10084,N_9998);
and U12659 (N_12659,N_11335,N_11539);
or U12660 (N_12660,N_11856,N_11713);
nand U12661 (N_12661,N_9055,N_11463);
and U12662 (N_12662,N_11495,N_8954);
and U12663 (N_12663,N_9977,N_11125);
and U12664 (N_12664,N_9732,N_11904);
and U12665 (N_12665,N_8669,N_10277);
nand U12666 (N_12666,N_10119,N_8195);
or U12667 (N_12667,N_8180,N_10900);
or U12668 (N_12668,N_9593,N_10933);
xnor U12669 (N_12669,N_8468,N_9500);
nand U12670 (N_12670,N_8273,N_9488);
or U12671 (N_12671,N_8015,N_9378);
or U12672 (N_12672,N_9631,N_10243);
and U12673 (N_12673,N_10087,N_8519);
nor U12674 (N_12674,N_8761,N_10562);
nand U12675 (N_12675,N_10678,N_10503);
xor U12676 (N_12676,N_11167,N_9636);
or U12677 (N_12677,N_8434,N_11542);
xor U12678 (N_12678,N_8349,N_11460);
or U12679 (N_12679,N_11509,N_9742);
nor U12680 (N_12680,N_11871,N_8208);
nand U12681 (N_12681,N_8396,N_10274);
and U12682 (N_12682,N_11749,N_8069);
xor U12683 (N_12683,N_9194,N_11957);
and U12684 (N_12684,N_9596,N_10699);
nand U12685 (N_12685,N_10866,N_8982);
or U12686 (N_12686,N_8534,N_9006);
and U12687 (N_12687,N_9559,N_10746);
and U12688 (N_12688,N_9515,N_9622);
and U12689 (N_12689,N_11491,N_11159);
xnor U12690 (N_12690,N_10069,N_8898);
nor U12691 (N_12691,N_11691,N_11811);
or U12692 (N_12692,N_11343,N_11964);
or U12693 (N_12693,N_9530,N_10670);
nor U12694 (N_12694,N_10883,N_10687);
nand U12695 (N_12695,N_9423,N_11615);
nor U12696 (N_12696,N_8037,N_11265);
nor U12697 (N_12697,N_8173,N_8828);
nand U12698 (N_12698,N_9327,N_10398);
nand U12699 (N_12699,N_10996,N_10588);
or U12700 (N_12700,N_10194,N_9472);
nor U12701 (N_12701,N_10542,N_8552);
nor U12702 (N_12702,N_8401,N_11943);
nor U12703 (N_12703,N_10983,N_9745);
or U12704 (N_12704,N_8088,N_10140);
nor U12705 (N_12705,N_11312,N_10772);
or U12706 (N_12706,N_11913,N_10547);
nor U12707 (N_12707,N_9392,N_11795);
xnor U12708 (N_12708,N_11260,N_11069);
nor U12709 (N_12709,N_11965,N_11860);
or U12710 (N_12710,N_11392,N_10400);
xnor U12711 (N_12711,N_9133,N_10011);
nand U12712 (N_12712,N_8775,N_11808);
nor U12713 (N_12713,N_9238,N_11670);
xor U12714 (N_12714,N_8083,N_10141);
xnor U12715 (N_12715,N_8657,N_11869);
xnor U12716 (N_12716,N_8730,N_11498);
and U12717 (N_12717,N_10054,N_8499);
nor U12718 (N_12718,N_10965,N_11601);
nand U12719 (N_12719,N_10517,N_9709);
and U12720 (N_12720,N_11151,N_8155);
nand U12721 (N_12721,N_10803,N_11881);
xor U12722 (N_12722,N_10978,N_9081);
nand U12723 (N_12723,N_10085,N_8279);
nand U12724 (N_12724,N_8097,N_11242);
or U12725 (N_12725,N_9223,N_11501);
nor U12726 (N_12726,N_10834,N_10124);
nand U12727 (N_12727,N_10737,N_10731);
and U12728 (N_12728,N_8135,N_8554);
nor U12729 (N_12729,N_9779,N_11948);
or U12730 (N_12730,N_9449,N_11158);
and U12731 (N_12731,N_11788,N_11829);
or U12732 (N_12732,N_8162,N_11722);
and U12733 (N_12733,N_10481,N_9499);
nor U12734 (N_12734,N_11459,N_10387);
nor U12735 (N_12735,N_9321,N_9672);
nor U12736 (N_12736,N_8369,N_8393);
or U12737 (N_12737,N_8666,N_9812);
xnor U12738 (N_12738,N_8440,N_10053);
nand U12739 (N_12739,N_10036,N_11695);
and U12740 (N_12740,N_10530,N_9749);
nand U12741 (N_12741,N_9960,N_8378);
or U12742 (N_12742,N_10816,N_8980);
nand U12743 (N_12743,N_9591,N_11803);
and U12744 (N_12744,N_9904,N_11422);
nand U12745 (N_12745,N_8674,N_9247);
nand U12746 (N_12746,N_8721,N_8634);
nor U12747 (N_12747,N_9439,N_9519);
nand U12748 (N_12748,N_10742,N_9634);
and U12749 (N_12749,N_11426,N_9892);
or U12750 (N_12750,N_8672,N_8501);
nand U12751 (N_12751,N_11518,N_10502);
nor U12752 (N_12752,N_11419,N_9455);
and U12753 (N_12753,N_11753,N_9706);
xor U12754 (N_12754,N_9168,N_8029);
xnor U12755 (N_12755,N_9428,N_9309);
nor U12756 (N_12756,N_8542,N_9784);
and U12757 (N_12757,N_10169,N_8626);
and U12758 (N_12758,N_8541,N_10311);
and U12759 (N_12759,N_9215,N_8390);
xor U12760 (N_12760,N_9085,N_10688);
xor U12761 (N_12761,N_10228,N_8577);
nor U12762 (N_12762,N_10231,N_8742);
nand U12763 (N_12763,N_10872,N_10257);
xor U12764 (N_12764,N_10473,N_9117);
or U12765 (N_12765,N_11731,N_10692);
and U12766 (N_12766,N_8461,N_10951);
and U12767 (N_12767,N_8132,N_11183);
nand U12768 (N_12768,N_11458,N_10515);
or U12769 (N_12769,N_11522,N_10693);
nand U12770 (N_12770,N_9278,N_9343);
nand U12771 (N_12771,N_11356,N_9180);
or U12772 (N_12772,N_11480,N_11845);
or U12773 (N_12773,N_9721,N_8335);
nor U12774 (N_12774,N_11656,N_9762);
xnor U12775 (N_12775,N_11374,N_9477);
or U12776 (N_12776,N_11746,N_9658);
nand U12777 (N_12777,N_10922,N_10113);
nor U12778 (N_12778,N_10484,N_9541);
and U12779 (N_12779,N_11149,N_10877);
and U12780 (N_12780,N_11431,N_11013);
nand U12781 (N_12781,N_10302,N_8266);
and U12782 (N_12782,N_10253,N_10736);
nor U12783 (N_12783,N_10553,N_8791);
and U12784 (N_12784,N_9956,N_10664);
or U12785 (N_12785,N_9987,N_10039);
nor U12786 (N_12786,N_11569,N_10637);
or U12787 (N_12787,N_9352,N_10179);
nor U12788 (N_12788,N_11921,N_8288);
nor U12789 (N_12789,N_11867,N_9693);
and U12790 (N_12790,N_10215,N_8748);
nand U12791 (N_12791,N_11031,N_10898);
nor U12792 (N_12792,N_11313,N_10571);
and U12793 (N_12793,N_9545,N_11441);
nand U12794 (N_12794,N_9080,N_8757);
and U12795 (N_12795,N_10574,N_8237);
nand U12796 (N_12796,N_8050,N_11116);
or U12797 (N_12797,N_9178,N_11855);
and U12798 (N_12798,N_8682,N_8004);
nand U12799 (N_12799,N_10110,N_8522);
nor U12800 (N_12800,N_11152,N_10478);
nand U12801 (N_12801,N_11745,N_10158);
nand U12802 (N_12802,N_10076,N_10028);
nand U12803 (N_12803,N_10287,N_9830);
or U12804 (N_12804,N_9971,N_8456);
nand U12805 (N_12805,N_8853,N_9107);
or U12806 (N_12806,N_11473,N_8977);
nand U12807 (N_12807,N_10101,N_11210);
xor U12808 (N_12808,N_10889,N_10186);
and U12809 (N_12809,N_9098,N_10512);
nand U12810 (N_12810,N_8267,N_8190);
nand U12811 (N_12811,N_11200,N_8188);
nor U12812 (N_12812,N_9091,N_8236);
and U12813 (N_12813,N_10735,N_9319);
or U12814 (N_12814,N_8442,N_10081);
or U12815 (N_12815,N_9044,N_10722);
nor U12816 (N_12816,N_11520,N_10836);
or U12817 (N_12817,N_9270,N_11577);
and U12818 (N_12818,N_9005,N_8171);
or U12819 (N_12819,N_10199,N_9757);
and U12820 (N_12820,N_11892,N_9882);
nor U12821 (N_12821,N_8432,N_8428);
xnor U12822 (N_12822,N_11493,N_9886);
xor U12823 (N_12823,N_8565,N_9607);
and U12824 (N_12824,N_10332,N_9221);
nor U12825 (N_12825,N_11478,N_11049);
and U12826 (N_12826,N_9116,N_11135);
and U12827 (N_12827,N_8975,N_10247);
and U12828 (N_12828,N_8824,N_9274);
and U12829 (N_12829,N_10014,N_8238);
nand U12830 (N_12830,N_11082,N_11393);
or U12831 (N_12831,N_10550,N_11345);
nand U12832 (N_12832,N_8970,N_11841);
xnor U12833 (N_12833,N_9612,N_9140);
or U12834 (N_12834,N_9405,N_10330);
xor U12835 (N_12835,N_11236,N_10470);
or U12836 (N_12836,N_11693,N_8416);
or U12837 (N_12837,N_8352,N_10061);
nand U12838 (N_12838,N_11562,N_8299);
or U12839 (N_12839,N_10304,N_10860);
or U12840 (N_12840,N_10538,N_10752);
and U12841 (N_12841,N_9305,N_10222);
nand U12842 (N_12842,N_9301,N_10306);
or U12843 (N_12843,N_11593,N_11604);
or U12844 (N_12844,N_8524,N_9017);
nand U12845 (N_12845,N_11170,N_11696);
nand U12846 (N_12846,N_10590,N_11103);
nand U12847 (N_12847,N_11025,N_11259);
nand U12848 (N_12848,N_9433,N_11735);
and U12849 (N_12849,N_10520,N_8463);
nor U12850 (N_12850,N_11003,N_11063);
xor U12851 (N_12851,N_8810,N_10345);
nand U12852 (N_12852,N_11409,N_8886);
nor U12853 (N_12853,N_11684,N_10344);
or U12854 (N_12854,N_9143,N_11544);
and U12855 (N_12855,N_10855,N_8526);
or U12856 (N_12856,N_11661,N_8023);
and U12857 (N_12857,N_11276,N_9531);
nand U12858 (N_12858,N_10845,N_8687);
nand U12859 (N_12859,N_11623,N_9146);
nor U12860 (N_12860,N_9713,N_8746);
nor U12861 (N_12861,N_11038,N_10285);
and U12862 (N_12862,N_10501,N_8010);
or U12863 (N_12863,N_9190,N_10425);
nor U12864 (N_12864,N_11954,N_11382);
nand U12865 (N_12865,N_8612,N_10262);
nand U12866 (N_12866,N_10998,N_11977);
or U12867 (N_12867,N_11092,N_11863);
and U12868 (N_12868,N_8189,N_8753);
nor U12869 (N_12869,N_9863,N_9752);
or U12870 (N_12870,N_10496,N_9252);
xnor U12871 (N_12871,N_9789,N_11000);
nand U12872 (N_12872,N_8313,N_11179);
nand U12873 (N_12873,N_10463,N_11830);
nand U12874 (N_12874,N_8860,N_10408);
nand U12875 (N_12875,N_9147,N_9481);
and U12876 (N_12876,N_9357,N_11323);
nor U12877 (N_12877,N_8650,N_8638);
and U12878 (N_12878,N_10919,N_8978);
nor U12879 (N_12879,N_11667,N_10796);
nor U12880 (N_12880,N_11543,N_8979);
nand U12881 (N_12881,N_8644,N_10099);
and U12882 (N_12882,N_10497,N_9839);
and U12883 (N_12883,N_11219,N_8020);
nor U12884 (N_12884,N_8645,N_9193);
nor U12885 (N_12885,N_11571,N_11055);
nor U12886 (N_12886,N_11836,N_9041);
nor U12887 (N_12887,N_9056,N_11798);
and U12888 (N_12888,N_10887,N_9429);
nand U12889 (N_12889,N_8002,N_10712);
nor U12890 (N_12890,N_9335,N_10956);
and U12891 (N_12891,N_10810,N_8116);
nor U12892 (N_12892,N_11678,N_8862);
xnor U12893 (N_12893,N_9670,N_9490);
or U12894 (N_12894,N_9920,N_10091);
and U12895 (N_12895,N_10955,N_8584);
or U12896 (N_12896,N_11224,N_8818);
or U12897 (N_12897,N_10494,N_9220);
xor U12898 (N_12898,N_10776,N_11898);
nor U12899 (N_12899,N_11872,N_8469);
or U12900 (N_12900,N_10823,N_11636);
or U12901 (N_12901,N_9957,N_10050);
nor U12902 (N_12902,N_11299,N_9101);
nand U12903 (N_12903,N_11143,N_9484);
or U12904 (N_12904,N_11824,N_11488);
nor U12905 (N_12905,N_11535,N_8147);
and U12906 (N_12906,N_10674,N_8153);
and U12907 (N_12907,N_8656,N_9462);
and U12908 (N_12908,N_8129,N_8586);
xnor U12909 (N_12909,N_11596,N_10777);
and U12910 (N_12910,N_9132,N_10453);
or U12911 (N_12911,N_10111,N_8272);
and U12912 (N_12912,N_10358,N_11213);
or U12913 (N_12913,N_9432,N_9946);
and U12914 (N_12914,N_11632,N_8453);
nor U12915 (N_12915,N_8724,N_11504);
nor U12916 (N_12916,N_9369,N_9915);
or U12917 (N_12917,N_9078,N_11377);
and U12918 (N_12918,N_10608,N_8999);
xnor U12919 (N_12919,N_10173,N_11878);
nor U12920 (N_12920,N_9811,N_10992);
or U12921 (N_12921,N_11755,N_8590);
and U12922 (N_12922,N_10382,N_10937);
nand U12923 (N_12923,N_11093,N_8960);
and U12924 (N_12924,N_8783,N_8253);
nand U12925 (N_12925,N_10525,N_10423);
and U12926 (N_12926,N_11538,N_9154);
nand U12927 (N_12927,N_10878,N_11673);
or U12928 (N_12928,N_11034,N_11530);
xor U12929 (N_12929,N_10421,N_9710);
or U12930 (N_12930,N_11507,N_8681);
or U12931 (N_12931,N_9770,N_8795);
nand U12932 (N_12932,N_10272,N_11759);
or U12933 (N_12933,N_10486,N_10879);
nor U12934 (N_12934,N_11216,N_9584);
nand U12935 (N_12935,N_8894,N_8061);
nor U12936 (N_12936,N_10528,N_10213);
or U12937 (N_12937,N_11347,N_11643);
xor U12938 (N_12938,N_8910,N_11758);
or U12939 (N_12939,N_11888,N_11231);
and U12940 (N_12940,N_8017,N_10646);
or U12941 (N_12941,N_9931,N_8580);
and U12942 (N_12942,N_9373,N_9540);
xnor U12943 (N_12943,N_11573,N_11708);
nand U12944 (N_12944,N_11111,N_9393);
nor U12945 (N_12945,N_11247,N_9503);
xor U12946 (N_12946,N_10669,N_8578);
nor U12947 (N_12947,N_10275,N_10283);
nor U12948 (N_12948,N_11582,N_8762);
nor U12949 (N_12949,N_8311,N_10064);
and U12950 (N_12950,N_10145,N_8628);
and U12951 (N_12951,N_11440,N_9128);
nand U12952 (N_12952,N_8079,N_8922);
or U12953 (N_12953,N_9468,N_10404);
or U12954 (N_12954,N_11980,N_11086);
and U12955 (N_12955,N_10567,N_8855);
and U12956 (N_12956,N_11652,N_11107);
or U12957 (N_12957,N_10711,N_10927);
nor U12958 (N_12958,N_8920,N_9730);
or U12959 (N_12959,N_11609,N_10839);
and U12960 (N_12960,N_9842,N_10560);
or U12961 (N_12961,N_10129,N_8605);
nand U12962 (N_12962,N_11982,N_9865);
nand U12963 (N_12963,N_8232,N_9457);
xor U12964 (N_12964,N_8592,N_11438);
nand U12965 (N_12965,N_9768,N_9798);
or U12966 (N_12966,N_10545,N_10685);
xor U12967 (N_12967,N_11662,N_10675);
nor U12968 (N_12968,N_11701,N_11164);
nor U12969 (N_12969,N_8711,N_10807);
and U12970 (N_12970,N_11072,N_10078);
and U12971 (N_12971,N_9166,N_11344);
and U12972 (N_12972,N_10763,N_11229);
nand U12973 (N_12973,N_10605,N_9443);
and U12974 (N_12974,N_11396,N_10246);
nor U12975 (N_12975,N_11406,N_8001);
and U12976 (N_12976,N_9973,N_8138);
nor U12977 (N_12977,N_10072,N_11618);
and U12978 (N_12978,N_11046,N_10197);
or U12979 (N_12979,N_11804,N_10412);
and U12980 (N_12980,N_9135,N_9679);
or U12981 (N_12981,N_10943,N_11971);
nand U12982 (N_12982,N_11113,N_11773);
nor U12983 (N_12983,N_9570,N_11688);
or U12984 (N_12984,N_10726,N_8712);
and U12985 (N_12985,N_9409,N_8743);
or U12986 (N_12986,N_8412,N_9183);
nand U12987 (N_12987,N_10142,N_11174);
and U12988 (N_12988,N_8318,N_9283);
or U12989 (N_12989,N_9403,N_9910);
nor U12990 (N_12990,N_9344,N_10006);
nand U12991 (N_12991,N_10577,N_9097);
and U12992 (N_12992,N_10780,N_8991);
nor U12993 (N_12993,N_8483,N_11861);
nor U12994 (N_12994,N_10493,N_9654);
xnor U12995 (N_12995,N_10413,N_10033);
and U12996 (N_12996,N_8951,N_9197);
and U12997 (N_12997,N_11171,N_11014);
nand U12998 (N_12998,N_10696,N_8515);
xor U12999 (N_12999,N_10671,N_11767);
and U13000 (N_13000,N_8046,N_9494);
nand U13001 (N_13001,N_10828,N_11457);
and U13002 (N_13002,N_8120,N_9944);
or U13003 (N_13003,N_8719,N_11243);
nand U13004 (N_13004,N_10997,N_8985);
nor U13005 (N_13005,N_11994,N_11800);
nand U13006 (N_13006,N_8947,N_8262);
and U13007 (N_13007,N_11732,N_9173);
nand U13008 (N_13008,N_11631,N_10686);
nor U13009 (N_13009,N_10604,N_10747);
and U13010 (N_13010,N_10537,N_8874);
and U13011 (N_13011,N_11436,N_11421);
nand U13012 (N_13012,N_9543,N_11984);
nor U13013 (N_13013,N_10120,N_10041);
and U13014 (N_13014,N_8498,N_8376);
and U13015 (N_13015,N_10684,N_10368);
nor U13016 (N_13016,N_9996,N_8942);
xor U13017 (N_13017,N_11097,N_9053);
nand U13018 (N_13018,N_11059,N_9625);
or U13019 (N_13019,N_9880,N_11925);
and U13020 (N_13020,N_10558,N_10787);
nor U13021 (N_13021,N_8251,N_10212);
and U13022 (N_13022,N_10427,N_8797);
nor U13023 (N_13023,N_8158,N_9174);
nor U13024 (N_13024,N_8281,N_10184);
nor U13025 (N_13025,N_9776,N_11931);
nand U13026 (N_13026,N_10353,N_8003);
and U13027 (N_13027,N_10018,N_10700);
nor U13028 (N_13028,N_10543,N_8546);
nor U13029 (N_13029,N_9874,N_9465);
or U13030 (N_13030,N_8075,N_10783);
or U13031 (N_13031,N_11646,N_9513);
nor U13032 (N_13032,N_10075,N_8905);
nand U13033 (N_13033,N_9760,N_11258);
or U13034 (N_13034,N_9680,N_10614);
and U13035 (N_13035,N_9279,N_9263);
and U13036 (N_13036,N_10620,N_11805);
nor U13037 (N_13037,N_8863,N_9187);
or U13038 (N_13038,N_8007,N_8673);
nand U13039 (N_13039,N_10220,N_8031);
nor U13040 (N_13040,N_11902,N_8925);
nand U13041 (N_13041,N_11357,N_9337);
xor U13042 (N_13042,N_9953,N_9311);
or U13043 (N_13043,N_9496,N_9066);
nor U13044 (N_13044,N_10004,N_10483);
or U13045 (N_13045,N_8121,N_9404);
nor U13046 (N_13046,N_9208,N_9495);
nand U13047 (N_13047,N_10395,N_11282);
and U13048 (N_13048,N_8549,N_11134);
nor U13049 (N_13049,N_10885,N_11102);
or U13050 (N_13050,N_10339,N_10000);
nor U13051 (N_13051,N_8032,N_8068);
and U13052 (N_13052,N_11303,N_10621);
or U13053 (N_13053,N_10324,N_11389);
and U13054 (N_13054,N_8934,N_11420);
nand U13055 (N_13055,N_10759,N_9786);
nand U13056 (N_13056,N_9914,N_8513);
nand U13057 (N_13057,N_9879,N_9366);
or U13058 (N_13058,N_10932,N_9959);
nand U13059 (N_13059,N_10260,N_11442);
and U13060 (N_13060,N_9381,N_8889);
or U13061 (N_13061,N_9711,N_8648);
xor U13062 (N_13062,N_11209,N_10058);
and U13063 (N_13063,N_9516,N_9691);
or U13064 (N_13064,N_11847,N_11366);
nor U13065 (N_13065,N_11585,N_11043);
and U13066 (N_13066,N_9159,N_11848);
nor U13067 (N_13067,N_8228,N_8705);
and U13068 (N_13068,N_11379,N_10739);
or U13069 (N_13069,N_9251,N_10649);
xor U13070 (N_13070,N_8739,N_11998);
or U13071 (N_13071,N_8572,N_9822);
nor U13072 (N_13072,N_10299,N_8562);
nand U13073 (N_13073,N_11208,N_8635);
and U13074 (N_13074,N_8642,N_8686);
nand U13075 (N_13075,N_11035,N_11075);
nand U13076 (N_13076,N_11412,N_8510);
and U13077 (N_13077,N_10429,N_10995);
and U13078 (N_13078,N_10704,N_10052);
and U13079 (N_13079,N_11703,N_11070);
nand U13080 (N_13080,N_10975,N_8537);
nand U13081 (N_13081,N_9601,N_10254);
nor U13082 (N_13082,N_10030,N_10067);
xor U13083 (N_13083,N_8493,N_11517);
nand U13084 (N_13084,N_9755,N_10576);
nor U13085 (N_13085,N_9847,N_9237);
xnor U13086 (N_13086,N_10853,N_9059);
and U13087 (N_13087,N_9766,N_9675);
or U13088 (N_13088,N_10941,N_11021);
nor U13089 (N_13089,N_10465,N_11207);
nand U13090 (N_13090,N_8192,N_9325);
xor U13091 (N_13091,N_8781,N_11677);
nor U13092 (N_13092,N_9514,N_11789);
or U13093 (N_13093,N_11024,N_8959);
or U13094 (N_13094,N_11318,N_8315);
xor U13095 (N_13095,N_11290,N_9667);
nor U13096 (N_13096,N_9780,N_10775);
nor U13097 (N_13097,N_9823,N_8560);
and U13098 (N_13098,N_9308,N_9111);
nand U13099 (N_13099,N_10177,N_10327);
nand U13100 (N_13100,N_9527,N_8136);
nand U13101 (N_13101,N_10371,N_10559);
nor U13102 (N_13102,N_8309,N_8215);
nor U13103 (N_13103,N_11911,N_11381);
xor U13104 (N_13104,N_10390,N_10824);
or U13105 (N_13105,N_8574,N_10942);
and U13106 (N_13106,N_10035,N_9253);
or U13107 (N_13107,N_10192,N_11198);
nand U13108 (N_13108,N_9995,N_8777);
or U13109 (N_13109,N_11564,N_9804);
nand U13110 (N_13110,N_9224,N_8382);
nand U13111 (N_13111,N_9354,N_8363);
and U13112 (N_13112,N_9809,N_9271);
or U13113 (N_13113,N_8119,N_9592);
and U13114 (N_13114,N_11716,N_10896);
and U13115 (N_13115,N_11565,N_10659);
nor U13116 (N_13116,N_10690,N_11418);
xnor U13117 (N_13117,N_10766,N_11645);
nor U13118 (N_13118,N_11138,N_9520);
xnor U13119 (N_13119,N_11770,N_9803);
and U13120 (N_13120,N_10833,N_9233);
nand U13121 (N_13121,N_10279,N_10325);
and U13122 (N_13122,N_10027,N_8843);
or U13123 (N_13123,N_9296,N_9763);
nor U13124 (N_13124,N_11001,N_8680);
and U13125 (N_13125,N_8284,N_9230);
and U13126 (N_13126,N_10135,N_9051);
nand U13127 (N_13127,N_8570,N_10162);
nand U13128 (N_13128,N_9790,N_10467);
nand U13129 (N_13129,N_11489,N_9510);
nor U13130 (N_13130,N_11084,N_11877);
nand U13131 (N_13131,N_11355,N_9483);
or U13132 (N_13132,N_9808,N_9165);
nor U13133 (N_13133,N_10492,N_11621);
nand U13134 (N_13134,N_10899,N_8117);
or U13135 (N_13135,N_8966,N_10351);
or U13136 (N_13136,N_10738,N_9845);
nor U13137 (N_13137,N_8402,N_11448);
and U13138 (N_13138,N_9119,N_8286);
nand U13139 (N_13139,N_8780,N_11169);
nand U13140 (N_13140,N_9087,N_9590);
and U13141 (N_13141,N_11586,N_8044);
or U13142 (N_13142,N_11704,N_10206);
and U13143 (N_13143,N_8038,N_9398);
or U13144 (N_13144,N_9551,N_8617);
nand U13145 (N_13145,N_8240,N_10401);
nor U13146 (N_13146,N_9200,N_11719);
nor U13147 (N_13147,N_8494,N_10181);
nor U13148 (N_13148,N_10544,N_10466);
nor U13149 (N_13149,N_8137,N_9624);
nand U13150 (N_13150,N_10661,N_11205);
nand U13151 (N_13151,N_11728,N_9772);
nand U13152 (N_13152,N_11961,N_10754);
nand U13153 (N_13153,N_9281,N_9120);
and U13154 (N_13154,N_8597,N_8800);
xnor U13155 (N_13155,N_8340,N_10055);
nand U13156 (N_13156,N_9153,N_9626);
nor U13157 (N_13157,N_8539,N_10925);
nor U13158 (N_13158,N_8295,N_10225);
xor U13159 (N_13159,N_8100,N_9518);
nand U13160 (N_13160,N_9163,N_9018);
nand U13161 (N_13161,N_9810,N_8231);
nand U13162 (N_13162,N_9615,N_11154);
xnor U13163 (N_13163,N_11371,N_11567);
and U13164 (N_13164,N_11144,N_9050);
or U13165 (N_13165,N_8651,N_8163);
and U13166 (N_13166,N_11747,N_8649);
nand U13167 (N_13167,N_9152,N_11675);
nor U13168 (N_13168,N_9284,N_8437);
and U13169 (N_13169,N_11252,N_10093);
and U13170 (N_13170,N_10534,N_9454);
or U13171 (N_13171,N_10709,N_8556);
nand U13172 (N_13172,N_11640,N_11160);
xnor U13173 (N_13173,N_9913,N_9289);
and U13174 (N_13174,N_11527,N_10298);
nor U13175 (N_13175,N_11561,N_10966);
nor U13176 (N_13176,N_10264,N_10021);
and U13177 (N_13177,N_10202,N_11218);
nor U13178 (N_13178,N_9562,N_10060);
and U13179 (N_13179,N_8630,N_8786);
or U13180 (N_13180,N_11157,N_11724);
nand U13181 (N_13181,N_8579,N_9903);
nor U13182 (N_13182,N_10723,N_9142);
nand U13183 (N_13183,N_8770,N_10631);
nand U13184 (N_13184,N_10837,N_11087);
and U13185 (N_13185,N_8688,N_10375);
or U13186 (N_13186,N_9512,N_8677);
nor U13187 (N_13187,N_10313,N_9446);
and U13188 (N_13188,N_8200,N_11121);
nand U13189 (N_13189,N_10112,N_10926);
xor U13190 (N_13190,N_8895,N_10676);
xnor U13191 (N_13191,N_8641,N_9161);
nor U13192 (N_13192,N_9767,N_10768);
nor U13193 (N_13193,N_11065,N_11124);
nor U13194 (N_13194,N_8071,N_10600);
or U13195 (N_13195,N_8842,N_8917);
nand U13196 (N_13196,N_8124,N_8902);
nand U13197 (N_13197,N_10673,N_9315);
and U13198 (N_13198,N_10229,N_11314);
nand U13199 (N_13199,N_10448,N_8604);
nor U13200 (N_13200,N_9297,N_9791);
nand U13201 (N_13201,N_8359,N_8387);
xor U13202 (N_13202,N_11349,N_10305);
and U13203 (N_13203,N_9286,N_9722);
nand U13204 (N_13204,N_8040,N_9788);
and U13205 (N_13205,N_8503,N_10268);
or U13206 (N_13206,N_11414,N_10821);
and U13207 (N_13207,N_8527,N_11095);
and U13208 (N_13208,N_9855,N_9924);
nand U13209 (N_13209,N_8418,N_8154);
nor U13210 (N_13210,N_11712,N_10459);
nand U13211 (N_13211,N_10115,N_9326);
nor U13212 (N_13212,N_8446,N_9579);
nand U13213 (N_13213,N_8283,N_11941);
xor U13214 (N_13214,N_8248,N_9148);
nor U13215 (N_13215,N_11748,N_8703);
and U13216 (N_13216,N_9475,N_9144);
nor U13217 (N_13217,N_8157,N_11165);
and U13218 (N_13218,N_8941,N_9858);
nand U13219 (N_13219,N_11725,N_10037);
nand U13220 (N_13220,N_10046,N_11106);
nand U13221 (N_13221,N_10256,N_11541);
and U13222 (N_13222,N_8547,N_8858);
or U13223 (N_13223,N_11909,N_9028);
xnor U13224 (N_13224,N_11574,N_8702);
or U13225 (N_13225,N_10689,N_9277);
nor U13226 (N_13226,N_11993,N_11275);
and U13227 (N_13227,N_8048,N_10133);
nor U13228 (N_13228,N_8011,N_11115);
and U13229 (N_13229,N_11516,N_11723);
xnor U13230 (N_13230,N_9890,N_9391);
nor U13231 (N_13231,N_8049,N_10118);
and U13232 (N_13232,N_11147,N_11914);
and U13233 (N_13233,N_9554,N_9980);
xor U13234 (N_13234,N_11917,N_10745);
and U13235 (N_13235,N_9982,N_10044);
or U13236 (N_13236,N_8512,N_8054);
xnor U13237 (N_13237,N_11114,N_11778);
and U13238 (N_13238,N_9492,N_9355);
and U13239 (N_13239,N_10144,N_10835);
nor U13240 (N_13240,N_11119,N_8345);
nor U13241 (N_13241,N_8883,N_9756);
nand U13242 (N_13242,N_8179,N_10830);
or U13243 (N_13243,N_11515,N_11360);
or U13244 (N_13244,N_9577,N_10239);
nor U13245 (N_13245,N_8006,N_11552);
and U13246 (N_13246,N_9435,N_11485);
or U13247 (N_13247,N_8931,N_11595);
nor U13248 (N_13248,N_9902,N_8487);
nand U13249 (N_13249,N_9979,N_10750);
and U13250 (N_13250,N_8039,N_8316);
or U13251 (N_13251,N_9704,N_11142);
nor U13252 (N_13252,N_9827,N_11821);
nand U13253 (N_13253,N_11437,N_9964);
and U13254 (N_13254,N_9875,N_11470);
nand U13255 (N_13255,N_8087,N_11400);
or U13256 (N_13256,N_9185,N_11233);
and U13257 (N_13257,N_9323,N_8292);
or U13258 (N_13258,N_11882,N_11301);
nor U13259 (N_13259,N_11955,N_8374);
nor U13260 (N_13260,N_8076,N_8698);
xor U13261 (N_13261,N_8618,N_9881);
xor U13262 (N_13262,N_9314,N_8747);
nand U13263 (N_13263,N_11709,N_10340);
and U13264 (N_13264,N_10934,N_9628);
nor U13265 (N_13265,N_10303,N_9926);
nor U13266 (N_13266,N_8585,N_10691);
nor U13267 (N_13267,N_10221,N_8836);
and U13268 (N_13268,N_8983,N_9048);
nand U13269 (N_13269,N_11697,N_9491);
nor U13270 (N_13270,N_8700,N_8772);
nor U13271 (N_13271,N_9250,N_11987);
and U13272 (N_13272,N_10627,N_8582);
nand U13273 (N_13273,N_9245,N_11109);
or U13274 (N_13274,N_10286,N_11588);
or U13275 (N_13275,N_9702,N_10355);
xnor U13276 (N_13276,N_9195,N_9227);
or U13277 (N_13277,N_10628,N_8198);
nand U13278 (N_13278,N_11461,N_11094);
nor U13279 (N_13279,N_9016,N_10038);
and U13280 (N_13280,N_9657,N_10770);
and U13281 (N_13281,N_10875,N_8360);
nor U13282 (N_13282,N_10697,N_10334);
or U13283 (N_13283,N_10097,N_10043);
and U13284 (N_13284,N_11309,N_11810);
or U13285 (N_13285,N_8816,N_10705);
xor U13286 (N_13286,N_9782,N_8713);
or U13287 (N_13287,N_8831,N_9950);
nand U13288 (N_13288,N_11608,N_10437);
and U13289 (N_13289,N_9257,N_8988);
or U13290 (N_13290,N_8477,N_9442);
nand U13291 (N_13291,N_11068,N_9861);
and U13292 (N_13292,N_10778,N_10572);
nor U13293 (N_13293,N_11053,N_8832);
nand U13294 (N_13294,N_10976,N_11837);
nor U13295 (N_13295,N_10913,N_9565);
and U13296 (N_13296,N_9734,N_8600);
or U13297 (N_13297,N_8476,N_11342);
or U13298 (N_13298,N_10917,N_8854);
and U13299 (N_13299,N_9700,N_11320);
and U13300 (N_13300,N_11390,N_11832);
nand U13301 (N_13301,N_9102,N_10601);
nand U13302 (N_13302,N_8383,N_10012);
and U13303 (N_13303,N_8878,N_9589);
and U13304 (N_13304,N_9340,N_10428);
or U13305 (N_13305,N_9747,N_11353);
nand U13306 (N_13306,N_11995,N_9456);
and U13307 (N_13307,N_8371,N_8287);
or U13308 (N_13308,N_8907,N_10874);
or U13309 (N_13309,N_8833,N_11737);
and U13310 (N_13310,N_9438,N_9859);
xor U13311 (N_13311,N_9445,N_8857);
or U13312 (N_13312,N_8367,N_10377);
xor U13313 (N_13313,N_9716,N_8258);
nor U13314 (N_13314,N_9877,N_10557);
nor U13315 (N_13315,N_11402,N_11536);
nor U13316 (N_13316,N_10270,N_10897);
nand U13317 (N_13317,N_10153,N_8769);
and U13318 (N_13318,N_8172,N_9895);
xor U13319 (N_13319,N_11614,N_8072);
nor U13320 (N_13320,N_11729,N_9396);
xor U13321 (N_13321,N_10619,N_11270);
nor U13322 (N_13322,N_10291,N_9669);
or U13323 (N_13323,N_11454,N_9365);
xnor U13324 (N_13324,N_10568,N_11846);
or U13325 (N_13325,N_11694,N_11757);
and U13326 (N_13326,N_9364,N_11525);
xor U13327 (N_13327,N_8508,N_11071);
nor U13328 (N_13328,N_10266,N_10007);
xor U13329 (N_13329,N_9648,N_9851);
and U13330 (N_13330,N_9951,N_10098);
or U13331 (N_13331,N_11424,N_9131);
and U13332 (N_13332,N_10160,N_9602);
or U13333 (N_13333,N_8045,N_8009);
or U13334 (N_13334,N_8156,N_9617);
nor U13335 (N_13335,N_9643,N_11844);
or U13336 (N_13336,N_11733,N_9265);
nor U13337 (N_13337,N_11332,N_10211);
or U13338 (N_13338,N_10786,N_11554);
nor U13339 (N_13339,N_9123,N_9431);
or U13340 (N_13340,N_8411,N_11505);
and U13341 (N_13341,N_9022,N_8472);
and U13342 (N_13342,N_10829,N_9320);
nor U13343 (N_13343,N_10267,N_11211);
or U13344 (N_13344,N_8559,N_10510);
and U13345 (N_13345,N_9150,N_10977);
nor U13346 (N_13346,N_11815,N_9552);
and U13347 (N_13347,N_10884,N_10598);
or U13348 (N_13348,N_10606,N_9402);
or U13349 (N_13349,N_9368,N_9160);
and U13350 (N_13350,N_8841,N_11397);
nand U13351 (N_13351,N_11813,N_8811);
or U13352 (N_13352,N_11081,N_10861);
nand U13353 (N_13353,N_11532,N_10578);
or U13354 (N_13354,N_11799,N_9907);
nor U13355 (N_13355,N_11548,N_11664);
nand U13356 (N_13356,N_11506,N_11326);
xor U13357 (N_13357,N_10660,N_8495);
nor U13358 (N_13358,N_10847,N_8744);
and U13359 (N_13359,N_10984,N_9497);
nor U13360 (N_13360,N_10813,N_11228);
nor U13361 (N_13361,N_10471,N_11962);
and U13362 (N_13362,N_10307,N_11950);
nand U13363 (N_13363,N_10506,N_10462);
xnor U13364 (N_13364,N_9653,N_10442);
and U13365 (N_13365,N_10411,N_8149);
nand U13366 (N_13366,N_11126,N_8073);
xor U13367 (N_13367,N_10954,N_9997);
and U13368 (N_13368,N_10989,N_10376);
and U13369 (N_13369,N_11791,N_10851);
nor U13370 (N_13370,N_8219,N_8385);
xnor U13371 (N_13371,N_10914,N_8520);
nand U13372 (N_13372,N_9652,N_10148);
nand U13373 (N_13373,N_9818,N_10579);
nor U13374 (N_13374,N_9867,N_10002);
nand U13375 (N_13375,N_11831,N_8289);
or U13376 (N_13376,N_10008,N_11876);
and U13377 (N_13377,N_9061,N_8303);
nand U13378 (N_13378,N_9395,N_9225);
nor U13379 (N_13379,N_8317,N_8938);
or U13380 (N_13380,N_8799,N_8904);
nor U13381 (N_13381,N_11681,N_8594);
nand U13382 (N_13382,N_8326,N_10630);
and U13383 (N_13383,N_11015,N_8337);
nand U13384 (N_13384,N_11938,N_8636);
and U13385 (N_13385,N_8595,N_8225);
and U13386 (N_13386,N_9406,N_11893);
and U13387 (N_13387,N_9942,N_10122);
nand U13388 (N_13388,N_9574,N_8353);
nand U13389 (N_13389,N_11283,N_9793);
and U13390 (N_13390,N_10819,N_11939);
and U13391 (N_13391,N_11156,N_11117);
or U13392 (N_13392,N_8754,N_10827);
and U13393 (N_13393,N_11822,N_8406);
nand U13394 (N_13394,N_11112,N_8400);
nor U13395 (N_13395,N_11907,N_11316);
nor U13396 (N_13396,N_11331,N_8193);
nand U13397 (N_13397,N_8962,N_10365);
or U13398 (N_13398,N_10741,N_8637);
nand U13399 (N_13399,N_11533,N_8325);
and U13400 (N_13400,N_8042,N_9932);
nor U13401 (N_13401,N_9571,N_10767);
nor U13402 (N_13402,N_8936,N_10797);
or U13403 (N_13403,N_8809,N_10982);
nand U13404 (N_13404,N_11296,N_10765);
xnor U13405 (N_13405,N_9089,N_10929);
and U13406 (N_13406,N_10308,N_9186);
nand U13407 (N_13407,N_8627,N_10591);
xor U13408 (N_13408,N_8624,N_10910);
and U13409 (N_13409,N_11992,N_10240);
nand U13410 (N_13410,N_10908,N_10364);
nor U13411 (N_13411,N_10526,N_9330);
nand U13412 (N_13412,N_8932,N_10507);
nand U13413 (N_13413,N_11960,N_10108);
nor U13414 (N_13414,N_11814,N_9511);
or U13415 (N_13415,N_8361,N_8408);
nand U13416 (N_13416,N_11849,N_8611);
and U13417 (N_13417,N_8827,N_10439);
nor U13418 (N_13418,N_8057,N_9919);
nor U13419 (N_13419,N_8835,N_9604);
xnor U13420 (N_13420,N_10551,N_11974);
nand U13421 (N_13421,N_11738,N_8395);
and U13422 (N_13422,N_9687,N_10403);
nor U13423 (N_13423,N_9482,N_8196);
nand U13424 (N_13424,N_9012,N_8140);
or U13425 (N_13425,N_11139,N_8964);
nand U13426 (N_13426,N_11787,N_9544);
nand U13427 (N_13427,N_10744,N_8643);
or U13428 (N_13428,N_10026,N_8473);
or U13429 (N_13429,N_10430,N_11058);
xnor U13430 (N_13430,N_10812,N_9727);
nand U13431 (N_13431,N_9176,N_11324);
and U13432 (N_13432,N_9800,N_10944);
and U13433 (N_13433,N_9204,N_8357);
nand U13434 (N_13434,N_10062,N_10402);
and U13435 (N_13435,N_8399,N_10195);
nor U13436 (N_13436,N_10056,N_9751);
xnor U13437 (N_13437,N_9467,N_11452);
or U13438 (N_13438,N_10717,N_8028);
nand U13439 (N_13439,N_10729,N_9502);
nand U13440 (N_13440,N_10329,N_10164);
and U13441 (N_13441,N_10248,N_8516);
nand U13442 (N_13442,N_9231,N_10801);
nor U13443 (N_13443,N_8768,N_9095);
xor U13444 (N_13444,N_11598,N_8879);
and U13445 (N_13445,N_10300,N_10862);
nand U13446 (N_13446,N_10882,N_10771);
or U13447 (N_13447,N_8897,N_11408);
nor U13448 (N_13448,N_8716,N_10921);
and U13449 (N_13449,N_11537,N_8758);
and U13450 (N_13450,N_9922,N_8185);
xnor U13451 (N_13451,N_9295,N_11740);
nand U13452 (N_13452,N_8243,N_10322);
or U13453 (N_13453,N_9030,N_10610);
nor U13454 (N_13454,N_10092,N_8314);
xor U13455 (N_13455,N_8089,N_10679);
and U13456 (N_13456,N_11937,N_10189);
and U13457 (N_13457,N_8269,N_9901);
and U13458 (N_13458,N_9678,N_10818);
and U13459 (N_13459,N_9860,N_10420);
and U13460 (N_13460,N_10848,N_9071);
nor U13461 (N_13461,N_8930,N_10476);
and U13462 (N_13462,N_11193,N_11433);
or U13463 (N_13463,N_9843,N_8601);
or U13464 (N_13464,N_8436,N_9461);
nand U13465 (N_13465,N_10151,N_10331);
nand U13466 (N_13466,N_9641,N_11137);
or U13467 (N_13467,N_10359,N_11130);
or U13468 (N_13468,N_11449,N_9616);
and U13469 (N_13469,N_10611,N_9287);
or U13470 (N_13470,N_11503,N_10276);
or U13471 (N_13471,N_8561,N_9935);
or U13472 (N_13472,N_9748,N_11122);
and U13473 (N_13473,N_10842,N_9290);
nand U13474 (N_13474,N_10901,N_9113);
or U13475 (N_13475,N_8776,N_11524);
or U13476 (N_13476,N_8996,N_8427);
nor U13477 (N_13477,N_8671,N_8826);
and U13478 (N_13478,N_10457,N_11383);
nor U13479 (N_13479,N_9480,N_11783);
or U13480 (N_13480,N_11322,N_9627);
nor U13481 (N_13481,N_9234,N_11477);
and U13482 (N_13482,N_9349,N_8615);
nand U13483 (N_13483,N_8373,N_11241);
or U13484 (N_13484,N_8950,N_10892);
and U13485 (N_13485,N_11920,N_9025);
nand U13486 (N_13486,N_11935,N_8913);
nor U13487 (N_13487,N_10444,N_9665);
nand U13488 (N_13488,N_8532,N_10999);
or U13489 (N_13489,N_10373,N_9783);
or U13490 (N_13490,N_10720,N_11922);
or U13491 (N_13491,N_9572,N_10644);
xnor U13492 (N_13492,N_10323,N_8887);
and U13493 (N_13493,N_10963,N_10822);
or U13494 (N_13494,N_8159,N_9866);
or U13495 (N_13495,N_10475,N_9940);
or U13496 (N_13496,N_11027,N_11201);
and U13497 (N_13497,N_10250,N_11953);
nor U13498 (N_13498,N_10180,N_9136);
nand U13499 (N_13499,N_9273,N_11467);
nand U13500 (N_13500,N_10451,N_11576);
nand U13501 (N_13501,N_10370,N_9164);
nand U13502 (N_13502,N_10405,N_11042);
or U13503 (N_13503,N_10461,N_9644);
or U13504 (N_13504,N_8151,N_8723);
or U13505 (N_13505,N_8211,N_8274);
nor U13506 (N_13506,N_11717,N_8736);
and U13507 (N_13507,N_11199,N_8997);
and U13508 (N_13508,N_11008,N_8518);
and U13509 (N_13509,N_11989,N_9241);
or U13510 (N_13510,N_9108,N_8409);
nand U13511 (N_13511,N_9660,N_9458);
or U13512 (N_13512,N_8085,N_9797);
or U13513 (N_13513,N_8852,N_11287);
nand U13514 (N_13514,N_8678,N_11976);
nor U13515 (N_13515,N_9255,N_9015);
or U13516 (N_13516,N_10672,N_8837);
nor U13517 (N_13517,N_9226,N_10706);
nor U13518 (N_13518,N_10626,N_8429);
and U13519 (N_13519,N_9796,N_10994);
and U13520 (N_13520,N_9134,N_10102);
and U13521 (N_13521,N_8181,N_9505);
xor U13522 (N_13522,N_11430,N_9121);
or U13523 (N_13523,N_10261,N_11088);
and U13524 (N_13524,N_8990,N_8106);
or U13525 (N_13525,N_8707,N_11127);
nor U13526 (N_13526,N_10755,N_8912);
and U13527 (N_13527,N_10320,N_8065);
nor U13528 (N_13528,N_8514,N_10338);
nor U13529 (N_13529,N_10795,N_9390);
nor U13530 (N_13530,N_11826,N_11244);
xor U13531 (N_13531,N_9383,N_10946);
and U13532 (N_13532,N_11616,N_9887);
and U13533 (N_13533,N_9202,N_10756);
nand U13534 (N_13534,N_10970,N_10154);
xnor U13535 (N_13535,N_11635,N_8025);
nand U13536 (N_13536,N_9370,N_9367);
or U13537 (N_13537,N_9962,N_9211);
nand U13538 (N_13538,N_10049,N_11776);
or U13539 (N_13539,N_8838,N_10121);
nand U13540 (N_13540,N_11523,N_9262);
or U13541 (N_13541,N_10419,N_8928);
and U13542 (N_13542,N_11657,N_8919);
or U13543 (N_13543,N_8261,N_10034);
and U13544 (N_13544,N_10947,N_11659);
and U13545 (N_13545,N_10071,N_8176);
xor U13546 (N_13546,N_11886,N_11761);
nand U13547 (N_13547,N_8264,N_8161);
nor U13548 (N_13548,N_10282,N_8221);
or U13549 (N_13549,N_9254,N_9375);
and U13550 (N_13550,N_9259,N_10396);
or U13551 (N_13551,N_11336,N_10799);
nand U13552 (N_13552,N_10235,N_10125);
nand U13553 (N_13553,N_8861,N_9162);
or U13554 (N_13554,N_8290,N_10029);
or U13555 (N_13555,N_8167,N_10318);
or U13556 (N_13556,N_10258,N_11894);
or U13557 (N_13557,N_9171,N_10556);
and U13558 (N_13558,N_11302,N_8807);
nor U13559 (N_13559,N_10210,N_8614);
and U13560 (N_13560,N_8166,N_11581);
nor U13561 (N_13561,N_9656,N_10094);
nor U13562 (N_13562,N_10383,N_8679);
or U13563 (N_13563,N_8924,N_9963);
or U13564 (N_13564,N_9509,N_8254);
nor U13565 (N_13565,N_8435,N_10639);
xor U13566 (N_13566,N_11780,N_9303);
nand U13567 (N_13567,N_10023,N_10791);
xnor U13568 (N_13568,N_9878,N_9155);
or U13569 (N_13569,N_8710,N_10059);
and U13570 (N_13570,N_10146,N_10138);
nand U13571 (N_13571,N_9897,N_8125);
and U13572 (N_13572,N_10165,N_8986);
and U13573 (N_13573,N_10438,N_9759);
nor U13574 (N_13574,N_8530,N_9487);
or U13575 (N_13575,N_11842,N_10972);
and U13576 (N_13576,N_9192,N_8545);
nor U13577 (N_13577,N_11665,N_9341);
nand U13578 (N_13578,N_9585,N_8331);
nor U13579 (N_13579,N_9052,N_8111);
nand U13580 (N_13580,N_8415,N_10238);
and U13581 (N_13581,N_10725,N_8433);
nand U13582 (N_13582,N_8602,N_9177);
xnor U13583 (N_13583,N_10870,N_9264);
and U13584 (N_13584,N_9210,N_11620);
nor U13585 (N_13585,N_9397,N_11444);
and U13586 (N_13586,N_10314,N_8727);
or U13587 (N_13587,N_11131,N_10495);
and U13588 (N_13588,N_9104,N_11462);
and U13589 (N_13589,N_9898,N_11594);
xnor U13590 (N_13590,N_9242,N_9068);
and U13591 (N_13591,N_8492,N_9313);
xor U13592 (N_13592,N_11801,N_8764);
nor U13593 (N_13593,N_9414,N_9852);
or U13594 (N_13594,N_10016,N_11339);
nor U13595 (N_13595,N_9872,N_9743);
nor U13596 (N_13596,N_11206,N_10683);
and U13597 (N_13597,N_10088,N_11897);
or U13598 (N_13598,N_9407,N_9739);
nand U13599 (N_13599,N_11439,N_11096);
nor U13600 (N_13600,N_8321,N_11951);
nand U13601 (N_13601,N_9834,N_8658);
nor U13602 (N_13602,N_11085,N_9244);
and U13603 (N_13603,N_8212,N_11870);
nand U13604 (N_13604,N_11905,N_10793);
nand U13605 (N_13605,N_8450,N_10570);
and U13606 (N_13606,N_11264,N_8165);
nand U13607 (N_13607,N_8691,N_11628);
nand U13608 (N_13608,N_10207,N_9240);
nand U13609 (N_13609,N_9464,N_8976);
or U13610 (N_13610,N_9374,N_10940);
or U13611 (N_13611,N_9586,N_11079);
and U13612 (N_13612,N_8305,N_10677);
xnor U13613 (N_13613,N_11173,N_9684);
or U13614 (N_13614,N_8168,N_11120);
xnor U13615 (N_13615,N_8160,N_8692);
xor U13616 (N_13616,N_8621,N_8280);
nor U13617 (N_13617,N_10541,N_9870);
or U13618 (N_13618,N_11009,N_8388);
or U13619 (N_13619,N_10159,N_11291);
and U13620 (N_13620,N_9002,N_9958);
nand U13621 (N_13621,N_10968,N_10873);
or U13622 (N_13622,N_10045,N_11203);
or U13623 (N_13623,N_9092,N_8397);
and U13624 (N_13624,N_10309,N_8465);
or U13625 (N_13625,N_11557,N_8654);
nand U13626 (N_13626,N_8573,N_9905);
or U13627 (N_13627,N_11862,N_10297);
nor U13628 (N_13628,N_10764,N_10867);
nor U13629 (N_13629,N_11690,N_11521);
nand U13630 (N_13630,N_8448,N_9157);
xnor U13631 (N_13631,N_10881,N_9088);
nor U13632 (N_13632,N_10602,N_11760);
and U13633 (N_13633,N_9094,N_8771);
and U13634 (N_13634,N_11150,N_10800);
nor U13635 (N_13635,N_10856,N_10820);
nand U13636 (N_13636,N_8224,N_9460);
and U13637 (N_13637,N_11067,N_10209);
or U13638 (N_13638,N_11279,N_10409);
nand U13639 (N_13639,N_9504,N_11337);
nor U13640 (N_13640,N_11280,N_9869);
or U13641 (N_13641,N_10070,N_11427);
or U13642 (N_13642,N_11153,N_11471);
or U13643 (N_13643,N_10909,N_9975);
nor U13644 (N_13644,N_8419,N_9213);
and U13645 (N_13645,N_9635,N_8598);
nor U13646 (N_13646,N_8398,N_8223);
or U13647 (N_13647,N_11750,N_10773);
nor U13648 (N_13648,N_10681,N_11610);
nand U13649 (N_13649,N_9666,N_10166);
xor U13650 (N_13650,N_9560,N_8104);
nand U13651 (N_13651,N_8464,N_10594);
nor U13652 (N_13652,N_9894,N_11251);
or U13653 (N_13653,N_9329,N_10682);
or U13654 (N_13654,N_11110,N_11715);
nand U13655 (N_13655,N_11476,N_9288);
nand U13656 (N_13656,N_10214,N_11908);
or U13657 (N_13657,N_10987,N_8732);
nor U13658 (N_13658,N_9738,N_11933);
nand U13659 (N_13659,N_8871,N_10748);
nand U13660 (N_13660,N_8380,N_11988);
nand U13661 (N_13661,N_9876,N_11963);
or U13662 (N_13662,N_11679,N_10536);
or U13663 (N_13663,N_10916,N_9258);
and U13664 (N_13664,N_10155,N_9698);
and U13665 (N_13665,N_10259,N_9597);
and U13666 (N_13666,N_8278,N_9416);
nor U13667 (N_13667,N_11880,N_10868);
and U13668 (N_13668,N_11823,N_9947);
or U13669 (N_13669,N_9817,N_11373);
and U13670 (N_13670,N_9268,N_8704);
nand U13671 (N_13671,N_11212,N_10293);
nor U13672 (N_13672,N_8143,N_11890);
nand U13673 (N_13673,N_11825,N_9207);
nand U13674 (N_13674,N_8246,N_8690);
nand U13675 (N_13675,N_10446,N_8203);
nor U13676 (N_13676,N_11321,N_10511);
and U13677 (N_13677,N_11237,N_10273);
nand U13678 (N_13678,N_8884,N_8662);
or U13679 (N_13679,N_10895,N_11178);
nand U13680 (N_13680,N_9063,N_11286);
nor U13681 (N_13681,N_10350,N_8062);
or U13682 (N_13682,N_11184,N_8881);
nand U13683 (N_13683,N_10456,N_8971);
and U13684 (N_13684,N_9943,N_8095);
xnor U13685 (N_13685,N_10317,N_10643);
xor U13686 (N_13686,N_9026,N_10516);
and U13687 (N_13687,N_9556,N_8059);
nor U13688 (N_13688,N_11792,N_10653);
or U13689 (N_13689,N_10161,N_10031);
nor U13690 (N_13690,N_9773,N_10208);
nor U13691 (N_13691,N_11566,N_9816);
and U13692 (N_13692,N_8244,N_10289);
nand U13693 (N_13693,N_9201,N_8348);
or U13694 (N_13694,N_10849,N_11146);
or U13695 (N_13695,N_9345,N_8992);
nand U13696 (N_13696,N_8876,N_9353);
or U13697 (N_13697,N_8164,N_11884);
or U13698 (N_13698,N_10200,N_8968);
or U13699 (N_13699,N_9899,N_11256);
and U13700 (N_13700,N_8995,N_10586);
and U13701 (N_13701,N_9891,N_9339);
xor U13702 (N_13702,N_11979,N_11036);
or U13703 (N_13703,N_10838,N_8074);
xor U13704 (N_13704,N_9744,N_9384);
nor U13705 (N_13705,N_9837,N_8304);
nand U13706 (N_13706,N_9848,N_10953);
nand U13707 (N_13707,N_11168,N_9451);
nor U13708 (N_13708,N_8921,N_8720);
nand U13709 (N_13709,N_10523,N_9741);
nor U13710 (N_13710,N_11180,N_9400);
xor U13711 (N_13711,N_10612,N_9934);
xnor U13712 (N_13712,N_11967,N_10022);
nor U13713 (N_13713,N_11511,N_8759);
xor U13714 (N_13714,N_11284,N_9668);
or U13715 (N_13715,N_8242,N_11182);
nor U13716 (N_13716,N_8070,N_9885);
xor U13717 (N_13717,N_8271,N_8974);
or U13718 (N_13718,N_10185,N_11358);
and U13719 (N_13719,N_9167,N_9076);
and U13720 (N_13720,N_10703,N_11840);
and U13721 (N_13721,N_9753,N_10458);
and U13722 (N_13722,N_11793,N_11202);
nand U13723 (N_13723,N_10566,N_11297);
or U13724 (N_13724,N_9849,N_8749);
and U13725 (N_13725,N_11514,N_9009);
nor U13726 (N_13726,N_10509,N_9043);
or U13727 (N_13727,N_11239,N_11873);
nand U13728 (N_13728,N_9203,N_8593);
xor U13729 (N_13729,N_11267,N_11394);
xnor U13730 (N_13730,N_11983,N_10367);
and U13731 (N_13731,N_10841,N_9106);
or U13732 (N_13732,N_8067,N_8880);
or U13733 (N_13733,N_8126,N_10924);
nor U13734 (N_13734,N_9035,N_11936);
or U13735 (N_13735,N_10811,N_11771);
or U13736 (N_13736,N_9138,N_9040);
and U13737 (N_13737,N_10152,N_9122);
nand U13738 (N_13738,N_11274,N_8381);
and U13739 (N_13739,N_9983,N_9685);
or U13740 (N_13740,N_8664,N_11833);
xnor U13741 (N_13741,N_10979,N_11364);
and U13742 (N_13742,N_10721,N_10074);
nand U13743 (N_13743,N_11073,N_10589);
and U13744 (N_13744,N_11932,N_10147);
nor U13745 (N_13745,N_10232,N_9813);
and U13746 (N_13746,N_11255,N_10132);
nor U13747 (N_13747,N_10073,N_11368);
nand U13748 (N_13748,N_8233,N_8174);
nor U13749 (N_13749,N_9683,N_8021);
or U13750 (N_13750,N_11066,N_11710);
xor U13751 (N_13751,N_10561,N_8300);
nand U13752 (N_13752,N_9470,N_9682);
and U13753 (N_13753,N_8285,N_11827);
nand U13754 (N_13754,N_9778,N_11410);
nand U13755 (N_13755,N_10581,N_9728);
or U13756 (N_13756,N_9993,N_11627);
xnor U13757 (N_13757,N_8420,N_8616);
and U13758 (N_13758,N_8026,N_11450);
nand U13759 (N_13759,N_10593,N_10090);
nor U13760 (N_13760,N_8115,N_9386);
and U13761 (N_13761,N_10116,N_8701);
nor U13762 (N_13762,N_11472,N_10774);
nand U13763 (N_13763,N_8973,N_9000);
or U13764 (N_13764,N_9916,N_11956);
nand U13765 (N_13765,N_8141,N_10565);
nor U13766 (N_13766,N_8882,N_10749);
or U13767 (N_13767,N_11226,N_10042);
nor U13768 (N_13768,N_9379,N_8482);
nand U13769 (N_13769,N_9550,N_11519);
nor U13770 (N_13770,N_9126,N_9479);
nand U13771 (N_13771,N_8740,N_11078);
or U13772 (N_13772,N_8914,N_11133);
nand U13773 (N_13773,N_8386,N_9707);
and U13774 (N_13774,N_9774,N_8094);
nor U13775 (N_13775,N_11222,N_10433);
nor U13776 (N_13776,N_8102,N_11002);
nand U13777 (N_13777,N_8911,N_11162);
nor U13778 (N_13778,N_8372,N_8738);
nand U13779 (N_13779,N_10204,N_8909);
nor U13780 (N_13780,N_8569,N_11310);
nand U13781 (N_13781,N_9302,N_10223);
nor U13782 (N_13782,N_9528,N_8715);
nand U13783 (N_13783,N_9967,N_8256);
nand U13784 (N_13784,N_8484,N_11875);
and U13785 (N_13785,N_9888,N_9149);
or U13786 (N_13786,N_10499,N_11278);
nand U13787 (N_13787,N_9663,N_11011);
and U13788 (N_13788,N_8466,N_11263);
xor U13789 (N_13789,N_8027,N_9637);
nor U13790 (N_13790,N_8475,N_10337);
or U13791 (N_13791,N_11819,N_10854);
nand U13792 (N_13792,N_11591,N_8426);
nor U13793 (N_13793,N_11464,N_11891);
nand U13794 (N_13794,N_10613,N_8034);
and U13795 (N_13795,N_11487,N_10680);
and U13796 (N_13796,N_8660,N_9440);
and U13797 (N_13797,N_8796,N_8066);
and U13798 (N_13798,N_8056,N_11633);
or U13799 (N_13799,N_9578,N_8084);
nand U13800 (N_13800,N_9588,N_11901);
or U13801 (N_13801,N_11910,N_11445);
and U13802 (N_13802,N_8606,N_10640);
nor U13803 (N_13803,N_11674,N_11617);
or U13804 (N_13804,N_9696,N_8798);
nand U13805 (N_13805,N_8944,N_9079);
and U13806 (N_13806,N_9372,N_8187);
or U13807 (N_13807,N_10825,N_9332);
and U13808 (N_13808,N_9594,N_11700);
xnor U13809 (N_13809,N_10546,N_11578);
nor U13810 (N_13810,N_9042,N_11186);
nor U13811 (N_13811,N_11889,N_11234);
nor U13812 (N_13812,N_10656,N_10149);
or U13813 (N_13813,N_11650,N_8994);
and U13814 (N_13814,N_11413,N_9613);
nand U13815 (N_13815,N_8785,N_8207);
or U13816 (N_13816,N_8336,N_8726);
nand U13817 (N_13817,N_10708,N_9522);
nor U13818 (N_13818,N_8234,N_10939);
xnor U13819 (N_13819,N_9720,N_8424);
nand U13820 (N_13820,N_9836,N_8012);
and U13821 (N_13821,N_9733,N_11927);
xor U13822 (N_13822,N_8204,N_8981);
and U13823 (N_13823,N_9609,N_11388);
or U13824 (N_13824,N_8745,N_11029);
and U13825 (N_13825,N_11223,N_11181);
and U13826 (N_13826,N_8987,N_10354);
nor U13827 (N_13827,N_10269,N_9444);
nand U13828 (N_13828,N_8470,N_9489);
nand U13829 (N_13829,N_9718,N_8216);
and U13830 (N_13830,N_8984,N_9708);
and U13831 (N_13831,N_10732,N_11946);
nand U13832 (N_13832,N_11456,N_11399);
xnor U13833 (N_13833,N_11781,N_9941);
or U13834 (N_13834,N_10065,N_9649);
xor U13835 (N_13835,N_9775,N_8675);
and U13836 (N_13836,N_8365,N_8080);
nor U13837 (N_13837,N_9243,N_10434);
nor U13838 (N_13838,N_9212,N_10569);
nor U13839 (N_13839,N_11642,N_9595);
nand U13840 (N_13840,N_11839,N_9724);
nor U13841 (N_13841,N_11583,N_11638);
or U13842 (N_13842,N_10265,N_8767);
or U13843 (N_13843,N_9765,N_11796);
nor U13844 (N_13844,N_10936,N_11883);
xor U13845 (N_13845,N_10514,N_11370);
nor U13846 (N_13846,N_10230,N_11372);
and U13847 (N_13847,N_9807,N_10288);
xnor U13848 (N_13848,N_11363,N_9587);
or U13849 (N_13849,N_10280,N_10170);
and U13850 (N_13850,N_10582,N_9027);
nor U13851 (N_13851,N_11644,N_8226);
and U13852 (N_13852,N_8935,N_9697);
nand U13853 (N_13853,N_8815,N_11240);
and U13854 (N_13854,N_10080,N_10798);
or U13855 (N_13855,N_8217,N_9298);
xor U13856 (N_13856,N_10490,N_10657);
nand U13857 (N_13857,N_11611,N_10852);
or U13858 (N_13858,N_10399,N_8358);
and U13859 (N_13859,N_8958,N_11225);
nor U13860 (N_13860,N_10077,N_9826);
nor U13861 (N_13861,N_8024,N_10930);
or U13862 (N_13862,N_10587,N_11589);
nand U13863 (N_13863,N_8845,N_10130);
and U13864 (N_13864,N_8252,N_10086);
nand U13865 (N_13865,N_10950,N_9292);
or U13866 (N_13866,N_10668,N_8623);
and U13867 (N_13867,N_9463,N_9021);
or U13868 (N_13868,N_11529,N_8893);
nand U13869 (N_13869,N_11023,N_11930);
nand U13870 (N_13870,N_10840,N_11262);
and U13871 (N_13871,N_11928,N_8343);
nor U13872 (N_13872,N_8939,N_10480);
nor U13873 (N_13873,N_8528,N_11570);
nand U13874 (N_13874,N_11484,N_11555);
or U13875 (N_13875,N_9209,N_9182);
nand U13876 (N_13876,N_11940,N_10379);
nor U13877 (N_13877,N_11277,N_10964);
or U13878 (N_13878,N_9555,N_10290);
xor U13879 (N_13879,N_8183,N_11851);
and U13880 (N_13880,N_8900,N_11785);
nand U13881 (N_13881,N_10859,N_9526);
or U13882 (N_13882,N_11148,N_10005);
nor U13883 (N_13883,N_10003,N_11720);
xor U13884 (N_13884,N_8789,N_10363);
or U13885 (N_13885,N_8249,N_9184);
or U13886 (N_13886,N_9825,N_11185);
nor U13887 (N_13887,N_9829,N_10886);
or U13888 (N_13888,N_8685,N_11508);
nand U13889 (N_13889,N_8525,N_9736);
or U13890 (N_13890,N_8949,N_9639);
and U13891 (N_13891,N_9701,N_11838);
nand U13892 (N_13892,N_11556,N_9342);
and U13893 (N_13893,N_10719,N_8486);
nor U13894 (N_13894,N_11145,N_8368);
or U13895 (N_13895,N_9124,N_10967);
or U13896 (N_13896,N_8178,N_11629);
or U13897 (N_13897,N_8134,N_8825);
or U13898 (N_13898,N_9714,N_11714);
nor U13899 (N_13899,N_11341,N_10904);
and U13900 (N_13900,N_9524,N_8214);
nor U13901 (N_13901,N_11386,N_8485);
or U13902 (N_13902,N_10203,N_10714);
or U13903 (N_13903,N_10251,N_10891);
or U13904 (N_13904,N_9533,N_8081);
and U13905 (N_13905,N_8890,N_11996);
nor U13906 (N_13906,N_8077,N_10389);
or U13907 (N_13907,N_11403,N_11546);
xor U13908 (N_13908,N_10564,N_10233);
or U13909 (N_13909,N_9677,N_8354);
and U13910 (N_13910,N_10178,N_9712);
nor U13911 (N_13911,N_8301,N_9075);
nor U13912 (N_13912,N_9925,N_8422);
nand U13913 (N_13913,N_8112,N_10469);
or U13914 (N_13914,N_9642,N_10961);
nand U13915 (N_13915,N_9537,N_8474);
nand U13916 (N_13916,N_9990,N_11191);
or U13917 (N_13917,N_11852,N_8218);
nand U13918 (N_13918,N_10440,N_8101);
nor U13919 (N_13919,N_10187,N_8750);
or U13920 (N_13920,N_8969,N_10923);
or U13921 (N_13921,N_10040,N_8551);
nand U13922 (N_13922,N_10015,N_11330);
nor U13923 (N_13923,N_11572,N_9729);
or U13924 (N_13924,N_10624,N_10655);
or U13925 (N_13925,N_10907,N_9450);
and U13926 (N_13926,N_11490,N_11769);
or U13927 (N_13927,N_11019,N_9380);
or U13928 (N_13928,N_8347,N_11230);
xnor U13929 (N_13929,N_11479,N_8480);
or U13930 (N_13930,N_11843,N_11155);
nand U13931 (N_13931,N_10973,N_8943);
and U13932 (N_13932,N_11253,N_11062);
nor U13933 (N_13933,N_11736,N_11293);
or U13934 (N_13934,N_8423,N_8291);
or U13935 (N_13935,N_9893,N_9568);
and U13936 (N_13936,N_9346,N_10814);
or U13937 (N_13937,N_8222,N_9188);
nand U13938 (N_13938,N_9232,N_11929);
nand U13939 (N_13939,N_11999,N_11797);
or U13940 (N_13940,N_9206,N_11499);
xnor U13941 (N_13941,N_9127,N_8169);
xor U13942 (N_13942,N_10751,N_8521);
nand U13943 (N_13943,N_10980,N_8844);
nor U13944 (N_13944,N_10952,N_9671);
nor U13945 (N_13945,N_11915,N_9558);
nand U13946 (N_13946,N_8194,N_11630);
nor U13947 (N_13947,N_10888,N_8444);
and U13948 (N_13948,N_11786,N_9125);
and U13949 (N_13949,N_9282,N_8717);
nand U13950 (N_13950,N_8078,N_11973);
nor U13951 (N_13951,N_11161,N_8631);
nor U13952 (N_13952,N_11975,N_9093);
nand U13953 (N_13953,N_9976,N_11269);
nand U13954 (N_13954,N_8629,N_10001);
nor U13955 (N_13955,N_9645,N_9769);
or U13956 (N_13956,N_10618,N_8259);
and U13957 (N_13957,N_11176,N_8792);
or U13958 (N_13958,N_11271,N_8668);
nor U13959 (N_13959,N_10234,N_8093);
nor U13960 (N_13960,N_9664,N_8646);
xor U13961 (N_13961,N_8496,N_9614);
nand U13962 (N_13962,N_8608,N_11227);
nor U13963 (N_13963,N_9705,N_11682);
nor U13964 (N_13964,N_11465,N_10707);
and U13965 (N_13965,N_9408,N_9269);
or U13966 (N_13966,N_10662,N_9896);
xor U13967 (N_13967,N_8439,N_11772);
xnor U13968 (N_13968,N_8096,N_11782);
xor U13969 (N_13969,N_10378,N_8294);
nor U13970 (N_13970,N_9331,N_9478);
and U13971 (N_13971,N_8430,N_8655);
xor U13972 (N_13972,N_10762,N_11483);
nand U13973 (N_13973,N_9567,N_11790);
nand U13974 (N_13974,N_10667,N_11298);
nor U13975 (N_13975,N_9599,N_11651);
xor U13976 (N_13976,N_8098,N_10915);
nor U13977 (N_13977,N_8205,N_8536);
nand U13978 (N_13978,N_8230,N_11919);
and U13979 (N_13979,N_9090,N_10295);
nand U13980 (N_13980,N_11676,N_9805);
xnor U13981 (N_13981,N_8351,N_8639);
nor U13982 (N_13982,N_11850,N_8144);
nand U13983 (N_13983,N_9972,N_10694);
xnor U13984 (N_13984,N_8445,N_11698);
nand U13985 (N_13985,N_8270,N_9999);
nand U13986 (N_13986,N_8804,N_11706);
xnor U13987 (N_13987,N_10143,N_10388);
or U13988 (N_13988,N_8788,N_11762);
nor U13989 (N_13989,N_9086,N_11105);
nand U13990 (N_13990,N_10629,N_9856);
and U13991 (N_13991,N_10734,N_10580);
nor U13992 (N_13992,N_9923,N_11653);
nand U13993 (N_13993,N_11549,N_8110);
or U13994 (N_13994,N_9746,N_10635);
nand U13995 (N_13995,N_8787,N_8937);
nor U13996 (N_13996,N_11098,N_8332);
nand U13997 (N_13997,N_10651,N_8431);
xnor U13998 (N_13998,N_11315,N_8320);
or U13999 (N_13999,N_9889,N_8822);
or U14000 (N_14000,N_8401,N_11103);
nand U14001 (N_14001,N_8348,N_10231);
and U14002 (N_14002,N_11437,N_10279);
and U14003 (N_14003,N_11498,N_9272);
and U14004 (N_14004,N_10681,N_8610);
nand U14005 (N_14005,N_10138,N_10487);
or U14006 (N_14006,N_8282,N_10125);
nand U14007 (N_14007,N_8918,N_11275);
or U14008 (N_14008,N_8308,N_11196);
or U14009 (N_14009,N_11503,N_11773);
nand U14010 (N_14010,N_9907,N_10894);
or U14011 (N_14011,N_9383,N_9185);
or U14012 (N_14012,N_10741,N_8570);
xor U14013 (N_14013,N_8986,N_9424);
nor U14014 (N_14014,N_11997,N_9278);
or U14015 (N_14015,N_9305,N_9533);
nor U14016 (N_14016,N_9566,N_11998);
and U14017 (N_14017,N_10902,N_10945);
nor U14018 (N_14018,N_10647,N_8168);
or U14019 (N_14019,N_11242,N_9377);
nor U14020 (N_14020,N_11399,N_8884);
nand U14021 (N_14021,N_8833,N_10133);
nand U14022 (N_14022,N_10217,N_8350);
or U14023 (N_14023,N_9207,N_9942);
xnor U14024 (N_14024,N_8460,N_10435);
and U14025 (N_14025,N_8970,N_9202);
or U14026 (N_14026,N_11653,N_8530);
or U14027 (N_14027,N_8852,N_11144);
and U14028 (N_14028,N_8517,N_10904);
nand U14029 (N_14029,N_8304,N_9692);
and U14030 (N_14030,N_8100,N_11051);
and U14031 (N_14031,N_9186,N_9028);
nor U14032 (N_14032,N_9133,N_10593);
nor U14033 (N_14033,N_9372,N_9538);
or U14034 (N_14034,N_10931,N_9406);
nor U14035 (N_14035,N_10594,N_8752);
or U14036 (N_14036,N_9905,N_8034);
nor U14037 (N_14037,N_8665,N_10829);
nor U14038 (N_14038,N_9025,N_9868);
and U14039 (N_14039,N_11430,N_10087);
nand U14040 (N_14040,N_10372,N_10026);
nand U14041 (N_14041,N_9499,N_8183);
or U14042 (N_14042,N_10090,N_8211);
or U14043 (N_14043,N_9641,N_11518);
or U14044 (N_14044,N_11064,N_8387);
and U14045 (N_14045,N_10666,N_9428);
nor U14046 (N_14046,N_8822,N_11375);
and U14047 (N_14047,N_9292,N_9044);
or U14048 (N_14048,N_9971,N_9466);
and U14049 (N_14049,N_8373,N_9660);
or U14050 (N_14050,N_9496,N_9800);
and U14051 (N_14051,N_11561,N_8181);
nor U14052 (N_14052,N_8912,N_8141);
and U14053 (N_14053,N_9436,N_11518);
nor U14054 (N_14054,N_10811,N_11296);
and U14055 (N_14055,N_11610,N_8987);
and U14056 (N_14056,N_10013,N_11541);
nand U14057 (N_14057,N_8146,N_8036);
nor U14058 (N_14058,N_8962,N_11169);
or U14059 (N_14059,N_9322,N_8432);
or U14060 (N_14060,N_9425,N_8739);
and U14061 (N_14061,N_10049,N_11597);
nand U14062 (N_14062,N_9697,N_9879);
xnor U14063 (N_14063,N_10682,N_8115);
and U14064 (N_14064,N_8184,N_8872);
and U14065 (N_14065,N_10730,N_10289);
or U14066 (N_14066,N_11003,N_11146);
xor U14067 (N_14067,N_8175,N_9580);
or U14068 (N_14068,N_10804,N_8490);
or U14069 (N_14069,N_11724,N_11530);
and U14070 (N_14070,N_11555,N_8590);
xnor U14071 (N_14071,N_10878,N_10276);
nor U14072 (N_14072,N_8175,N_10705);
nor U14073 (N_14073,N_11348,N_9313);
nand U14074 (N_14074,N_11950,N_9513);
and U14075 (N_14075,N_10785,N_11910);
nor U14076 (N_14076,N_10308,N_11938);
nor U14077 (N_14077,N_9983,N_9296);
nand U14078 (N_14078,N_10906,N_11518);
and U14079 (N_14079,N_9673,N_9520);
nand U14080 (N_14080,N_11617,N_8252);
and U14081 (N_14081,N_10255,N_9646);
or U14082 (N_14082,N_11496,N_10072);
nand U14083 (N_14083,N_10569,N_8851);
nand U14084 (N_14084,N_11917,N_9308);
and U14085 (N_14085,N_10181,N_8316);
nand U14086 (N_14086,N_10632,N_8003);
nor U14087 (N_14087,N_10162,N_8683);
or U14088 (N_14088,N_9546,N_10203);
nor U14089 (N_14089,N_8162,N_10479);
and U14090 (N_14090,N_11427,N_8283);
and U14091 (N_14091,N_10157,N_11340);
or U14092 (N_14092,N_8989,N_11372);
or U14093 (N_14093,N_8811,N_10790);
nand U14094 (N_14094,N_10011,N_10017);
nand U14095 (N_14095,N_9730,N_8931);
nand U14096 (N_14096,N_11114,N_8465);
and U14097 (N_14097,N_9444,N_11184);
xor U14098 (N_14098,N_9028,N_10467);
nand U14099 (N_14099,N_10200,N_9914);
nand U14100 (N_14100,N_11496,N_8620);
or U14101 (N_14101,N_11973,N_11115);
and U14102 (N_14102,N_9421,N_11869);
and U14103 (N_14103,N_10153,N_8976);
xnor U14104 (N_14104,N_11870,N_10362);
nor U14105 (N_14105,N_8009,N_9532);
nand U14106 (N_14106,N_8143,N_8412);
nor U14107 (N_14107,N_10358,N_8736);
nor U14108 (N_14108,N_11308,N_10308);
nand U14109 (N_14109,N_9923,N_9882);
and U14110 (N_14110,N_9226,N_8749);
or U14111 (N_14111,N_11949,N_8269);
nor U14112 (N_14112,N_9567,N_8368);
or U14113 (N_14113,N_10635,N_9482);
nand U14114 (N_14114,N_10430,N_9495);
or U14115 (N_14115,N_9071,N_10240);
xor U14116 (N_14116,N_11872,N_10515);
and U14117 (N_14117,N_11409,N_8587);
or U14118 (N_14118,N_10144,N_10409);
nand U14119 (N_14119,N_9408,N_8255);
and U14120 (N_14120,N_11142,N_9284);
or U14121 (N_14121,N_9203,N_10456);
nand U14122 (N_14122,N_11163,N_10756);
and U14123 (N_14123,N_8630,N_9926);
nand U14124 (N_14124,N_8245,N_8875);
and U14125 (N_14125,N_8441,N_10642);
or U14126 (N_14126,N_8559,N_10239);
nand U14127 (N_14127,N_8008,N_9813);
and U14128 (N_14128,N_10781,N_8654);
nor U14129 (N_14129,N_11010,N_11236);
and U14130 (N_14130,N_11827,N_11130);
and U14131 (N_14131,N_9395,N_9630);
and U14132 (N_14132,N_11928,N_8866);
or U14133 (N_14133,N_10501,N_10648);
nor U14134 (N_14134,N_11345,N_11491);
xor U14135 (N_14135,N_8415,N_8723);
nand U14136 (N_14136,N_11902,N_8044);
nand U14137 (N_14137,N_9938,N_9214);
and U14138 (N_14138,N_8120,N_9772);
xnor U14139 (N_14139,N_11732,N_11345);
nand U14140 (N_14140,N_9819,N_11835);
nor U14141 (N_14141,N_9345,N_10297);
nand U14142 (N_14142,N_10137,N_8647);
xor U14143 (N_14143,N_11883,N_10338);
and U14144 (N_14144,N_10015,N_8432);
nor U14145 (N_14145,N_8437,N_9038);
nor U14146 (N_14146,N_8229,N_9666);
or U14147 (N_14147,N_10045,N_8706);
nand U14148 (N_14148,N_9881,N_11184);
nand U14149 (N_14149,N_8529,N_9060);
nand U14150 (N_14150,N_10152,N_11353);
and U14151 (N_14151,N_11030,N_11373);
or U14152 (N_14152,N_8944,N_9805);
nand U14153 (N_14153,N_8398,N_10232);
nor U14154 (N_14154,N_9103,N_11703);
and U14155 (N_14155,N_8911,N_11354);
or U14156 (N_14156,N_11151,N_11430);
and U14157 (N_14157,N_9738,N_9602);
and U14158 (N_14158,N_10839,N_10687);
or U14159 (N_14159,N_10353,N_8420);
xnor U14160 (N_14160,N_9703,N_8221);
and U14161 (N_14161,N_8831,N_8562);
and U14162 (N_14162,N_10637,N_9349);
or U14163 (N_14163,N_10373,N_10102);
nand U14164 (N_14164,N_8809,N_9393);
or U14165 (N_14165,N_10373,N_9790);
nor U14166 (N_14166,N_11563,N_10192);
nand U14167 (N_14167,N_9561,N_9861);
or U14168 (N_14168,N_8343,N_8044);
or U14169 (N_14169,N_11858,N_10809);
xor U14170 (N_14170,N_11712,N_10708);
or U14171 (N_14171,N_9804,N_11213);
and U14172 (N_14172,N_8664,N_8782);
nand U14173 (N_14173,N_8105,N_11155);
nand U14174 (N_14174,N_8300,N_11763);
xnor U14175 (N_14175,N_8717,N_8926);
nand U14176 (N_14176,N_10143,N_9712);
nand U14177 (N_14177,N_9095,N_8377);
nand U14178 (N_14178,N_9077,N_9765);
nor U14179 (N_14179,N_8190,N_9461);
xnor U14180 (N_14180,N_10215,N_11267);
and U14181 (N_14181,N_11665,N_10812);
xnor U14182 (N_14182,N_8180,N_8836);
nand U14183 (N_14183,N_8474,N_11163);
nor U14184 (N_14184,N_9111,N_11850);
and U14185 (N_14185,N_9891,N_8959);
or U14186 (N_14186,N_9436,N_10912);
nand U14187 (N_14187,N_9329,N_11186);
and U14188 (N_14188,N_11402,N_9874);
or U14189 (N_14189,N_10177,N_8261);
nor U14190 (N_14190,N_10698,N_11101);
nor U14191 (N_14191,N_10388,N_8379);
and U14192 (N_14192,N_11299,N_10781);
or U14193 (N_14193,N_8199,N_9245);
xnor U14194 (N_14194,N_10544,N_11327);
or U14195 (N_14195,N_10694,N_9120);
xor U14196 (N_14196,N_10264,N_9306);
nand U14197 (N_14197,N_9737,N_11049);
and U14198 (N_14198,N_10295,N_9629);
or U14199 (N_14199,N_10430,N_9137);
or U14200 (N_14200,N_10350,N_10431);
or U14201 (N_14201,N_9134,N_9820);
xnor U14202 (N_14202,N_11631,N_11194);
nand U14203 (N_14203,N_8137,N_8378);
xnor U14204 (N_14204,N_9486,N_9398);
and U14205 (N_14205,N_11031,N_10798);
or U14206 (N_14206,N_10529,N_8150);
nand U14207 (N_14207,N_10137,N_8871);
and U14208 (N_14208,N_10454,N_10208);
nand U14209 (N_14209,N_9552,N_8589);
and U14210 (N_14210,N_10615,N_10486);
nor U14211 (N_14211,N_8768,N_11062);
nand U14212 (N_14212,N_11638,N_10292);
xnor U14213 (N_14213,N_10232,N_11139);
nor U14214 (N_14214,N_9344,N_9359);
or U14215 (N_14215,N_11042,N_10293);
xor U14216 (N_14216,N_8110,N_9299);
xnor U14217 (N_14217,N_9748,N_11593);
and U14218 (N_14218,N_11794,N_8724);
or U14219 (N_14219,N_8238,N_10393);
nand U14220 (N_14220,N_9728,N_9011);
and U14221 (N_14221,N_10282,N_11708);
or U14222 (N_14222,N_11649,N_9758);
nor U14223 (N_14223,N_10266,N_8351);
and U14224 (N_14224,N_8738,N_9356);
xor U14225 (N_14225,N_8939,N_9458);
and U14226 (N_14226,N_8894,N_9212);
xor U14227 (N_14227,N_9416,N_10746);
and U14228 (N_14228,N_9466,N_9579);
and U14229 (N_14229,N_10817,N_9218);
nor U14230 (N_14230,N_8473,N_8631);
or U14231 (N_14231,N_10216,N_10117);
xnor U14232 (N_14232,N_9439,N_11026);
nor U14233 (N_14233,N_11259,N_8273);
nor U14234 (N_14234,N_9408,N_11208);
or U14235 (N_14235,N_11769,N_9665);
or U14236 (N_14236,N_8127,N_10826);
or U14237 (N_14237,N_10982,N_10665);
nand U14238 (N_14238,N_8346,N_10847);
nor U14239 (N_14239,N_11982,N_10048);
nor U14240 (N_14240,N_10375,N_10676);
nand U14241 (N_14241,N_8390,N_10154);
or U14242 (N_14242,N_9975,N_11139);
nand U14243 (N_14243,N_11696,N_8385);
nor U14244 (N_14244,N_11164,N_11892);
nor U14245 (N_14245,N_8298,N_10901);
or U14246 (N_14246,N_8693,N_9709);
nand U14247 (N_14247,N_11936,N_8848);
and U14248 (N_14248,N_9458,N_11835);
nor U14249 (N_14249,N_11169,N_9565);
xor U14250 (N_14250,N_9175,N_10034);
nor U14251 (N_14251,N_11743,N_8984);
nor U14252 (N_14252,N_8269,N_10557);
nor U14253 (N_14253,N_8190,N_8532);
or U14254 (N_14254,N_8216,N_8167);
nor U14255 (N_14255,N_9451,N_11155);
nor U14256 (N_14256,N_8241,N_10200);
or U14257 (N_14257,N_8997,N_9125);
and U14258 (N_14258,N_11331,N_10390);
nor U14259 (N_14259,N_9565,N_11807);
and U14260 (N_14260,N_9149,N_11491);
or U14261 (N_14261,N_11021,N_11151);
and U14262 (N_14262,N_10866,N_11694);
nor U14263 (N_14263,N_10165,N_11046);
nor U14264 (N_14264,N_10129,N_9544);
and U14265 (N_14265,N_11823,N_8040);
nand U14266 (N_14266,N_8788,N_11994);
xnor U14267 (N_14267,N_9114,N_8793);
nor U14268 (N_14268,N_9917,N_8141);
and U14269 (N_14269,N_11913,N_8128);
nor U14270 (N_14270,N_8459,N_9451);
nand U14271 (N_14271,N_8585,N_8811);
or U14272 (N_14272,N_11144,N_11058);
xor U14273 (N_14273,N_9933,N_10495);
nand U14274 (N_14274,N_11792,N_9188);
or U14275 (N_14275,N_11901,N_10002);
xnor U14276 (N_14276,N_10507,N_9112);
or U14277 (N_14277,N_9149,N_10177);
or U14278 (N_14278,N_9545,N_9641);
nand U14279 (N_14279,N_8688,N_11001);
and U14280 (N_14280,N_8539,N_8289);
or U14281 (N_14281,N_8644,N_10551);
nor U14282 (N_14282,N_10002,N_8730);
xor U14283 (N_14283,N_8565,N_8804);
nand U14284 (N_14284,N_10911,N_8356);
nor U14285 (N_14285,N_11718,N_9078);
nand U14286 (N_14286,N_10974,N_9399);
or U14287 (N_14287,N_8129,N_10480);
nand U14288 (N_14288,N_8018,N_11790);
nand U14289 (N_14289,N_9425,N_11414);
nand U14290 (N_14290,N_11596,N_10781);
nor U14291 (N_14291,N_11428,N_10617);
or U14292 (N_14292,N_11539,N_11534);
and U14293 (N_14293,N_11650,N_11603);
nor U14294 (N_14294,N_8855,N_8708);
nand U14295 (N_14295,N_9921,N_8371);
or U14296 (N_14296,N_11281,N_8513);
and U14297 (N_14297,N_10884,N_10483);
or U14298 (N_14298,N_8164,N_9903);
and U14299 (N_14299,N_8405,N_8503);
or U14300 (N_14300,N_11396,N_11899);
nor U14301 (N_14301,N_11793,N_9606);
nand U14302 (N_14302,N_8751,N_10577);
and U14303 (N_14303,N_10529,N_11290);
nand U14304 (N_14304,N_11919,N_9929);
nand U14305 (N_14305,N_8123,N_10562);
and U14306 (N_14306,N_11876,N_9105);
xor U14307 (N_14307,N_8938,N_9719);
nor U14308 (N_14308,N_10579,N_8644);
and U14309 (N_14309,N_8840,N_8406);
or U14310 (N_14310,N_8442,N_10573);
and U14311 (N_14311,N_11963,N_8196);
or U14312 (N_14312,N_11109,N_8878);
and U14313 (N_14313,N_11713,N_10415);
and U14314 (N_14314,N_9637,N_11802);
or U14315 (N_14315,N_8665,N_9747);
nand U14316 (N_14316,N_11867,N_9808);
nand U14317 (N_14317,N_9295,N_9864);
and U14318 (N_14318,N_10494,N_8112);
xnor U14319 (N_14319,N_8877,N_9117);
nor U14320 (N_14320,N_11941,N_10206);
nor U14321 (N_14321,N_9790,N_8729);
nor U14322 (N_14322,N_8691,N_9932);
nand U14323 (N_14323,N_8694,N_10542);
nor U14324 (N_14324,N_9045,N_11330);
nor U14325 (N_14325,N_11147,N_10086);
or U14326 (N_14326,N_11700,N_10251);
nand U14327 (N_14327,N_8322,N_10967);
and U14328 (N_14328,N_10924,N_9513);
nand U14329 (N_14329,N_10258,N_10137);
nand U14330 (N_14330,N_11215,N_9388);
and U14331 (N_14331,N_10775,N_11066);
nand U14332 (N_14332,N_8711,N_11607);
nor U14333 (N_14333,N_11898,N_9845);
and U14334 (N_14334,N_10968,N_11048);
nor U14335 (N_14335,N_9784,N_8628);
nor U14336 (N_14336,N_8356,N_9785);
or U14337 (N_14337,N_10379,N_9838);
and U14338 (N_14338,N_10898,N_9455);
nand U14339 (N_14339,N_8869,N_8439);
nor U14340 (N_14340,N_9273,N_10902);
nand U14341 (N_14341,N_8498,N_11499);
or U14342 (N_14342,N_11705,N_11267);
nand U14343 (N_14343,N_10588,N_11650);
nor U14344 (N_14344,N_10293,N_11146);
and U14345 (N_14345,N_11937,N_10326);
nand U14346 (N_14346,N_11702,N_9927);
nand U14347 (N_14347,N_8469,N_10064);
nor U14348 (N_14348,N_11165,N_8413);
nor U14349 (N_14349,N_11429,N_8025);
or U14350 (N_14350,N_8324,N_8757);
nand U14351 (N_14351,N_11974,N_9299);
nand U14352 (N_14352,N_9001,N_9918);
nor U14353 (N_14353,N_9036,N_8613);
and U14354 (N_14354,N_8193,N_10642);
and U14355 (N_14355,N_8458,N_8566);
and U14356 (N_14356,N_8364,N_8087);
or U14357 (N_14357,N_8172,N_11618);
nor U14358 (N_14358,N_8008,N_8350);
nor U14359 (N_14359,N_8967,N_9140);
nor U14360 (N_14360,N_8410,N_11449);
and U14361 (N_14361,N_11092,N_10403);
nor U14362 (N_14362,N_9409,N_8154);
xnor U14363 (N_14363,N_11190,N_8869);
nand U14364 (N_14364,N_9442,N_8304);
or U14365 (N_14365,N_10105,N_8805);
nand U14366 (N_14366,N_9738,N_9866);
or U14367 (N_14367,N_10807,N_11561);
nor U14368 (N_14368,N_8712,N_10410);
nor U14369 (N_14369,N_10940,N_9884);
or U14370 (N_14370,N_8226,N_8611);
and U14371 (N_14371,N_10643,N_8567);
nand U14372 (N_14372,N_10912,N_8008);
and U14373 (N_14373,N_8833,N_11558);
or U14374 (N_14374,N_11705,N_11246);
and U14375 (N_14375,N_9035,N_10228);
and U14376 (N_14376,N_9505,N_8395);
xnor U14377 (N_14377,N_11089,N_11833);
nand U14378 (N_14378,N_9778,N_10846);
or U14379 (N_14379,N_9661,N_11144);
and U14380 (N_14380,N_11841,N_10647);
nor U14381 (N_14381,N_8251,N_11802);
nor U14382 (N_14382,N_10105,N_8372);
and U14383 (N_14383,N_8242,N_10877);
nor U14384 (N_14384,N_8843,N_11071);
nand U14385 (N_14385,N_9516,N_8627);
nor U14386 (N_14386,N_11111,N_9285);
nor U14387 (N_14387,N_10451,N_9286);
nand U14388 (N_14388,N_8692,N_8307);
or U14389 (N_14389,N_11025,N_10527);
nor U14390 (N_14390,N_10714,N_11498);
nand U14391 (N_14391,N_10382,N_9769);
nand U14392 (N_14392,N_10635,N_9446);
nor U14393 (N_14393,N_9948,N_10749);
and U14394 (N_14394,N_11039,N_10683);
and U14395 (N_14395,N_10895,N_11298);
nand U14396 (N_14396,N_9412,N_10612);
nor U14397 (N_14397,N_9631,N_8244);
nand U14398 (N_14398,N_8242,N_11151);
or U14399 (N_14399,N_9321,N_10665);
and U14400 (N_14400,N_9310,N_8843);
or U14401 (N_14401,N_11116,N_9933);
nand U14402 (N_14402,N_9335,N_11628);
nor U14403 (N_14403,N_11918,N_9474);
nor U14404 (N_14404,N_8743,N_8759);
nor U14405 (N_14405,N_9548,N_10232);
or U14406 (N_14406,N_9896,N_11597);
nand U14407 (N_14407,N_8908,N_8900);
xor U14408 (N_14408,N_9903,N_11894);
or U14409 (N_14409,N_11444,N_10824);
and U14410 (N_14410,N_8396,N_8523);
xor U14411 (N_14411,N_9845,N_11755);
and U14412 (N_14412,N_10701,N_10492);
nand U14413 (N_14413,N_11573,N_11967);
nor U14414 (N_14414,N_8360,N_11099);
xor U14415 (N_14415,N_11105,N_10475);
nor U14416 (N_14416,N_11079,N_9785);
and U14417 (N_14417,N_11006,N_11595);
nor U14418 (N_14418,N_9230,N_8153);
nor U14419 (N_14419,N_11261,N_8173);
xor U14420 (N_14420,N_10405,N_10896);
nor U14421 (N_14421,N_11126,N_10097);
nor U14422 (N_14422,N_11364,N_8355);
or U14423 (N_14423,N_9719,N_8960);
and U14424 (N_14424,N_10550,N_10177);
nand U14425 (N_14425,N_10766,N_11720);
nand U14426 (N_14426,N_11507,N_8614);
nor U14427 (N_14427,N_8987,N_9506);
or U14428 (N_14428,N_11749,N_9514);
and U14429 (N_14429,N_10278,N_11999);
or U14430 (N_14430,N_11345,N_9342);
and U14431 (N_14431,N_9273,N_10929);
and U14432 (N_14432,N_8116,N_8894);
or U14433 (N_14433,N_8357,N_10831);
xor U14434 (N_14434,N_11090,N_10439);
and U14435 (N_14435,N_10885,N_10992);
or U14436 (N_14436,N_8741,N_9567);
and U14437 (N_14437,N_10985,N_8471);
nand U14438 (N_14438,N_9930,N_8107);
or U14439 (N_14439,N_10627,N_10801);
nor U14440 (N_14440,N_8100,N_10306);
nor U14441 (N_14441,N_8957,N_8357);
or U14442 (N_14442,N_11636,N_9694);
xor U14443 (N_14443,N_8581,N_8975);
and U14444 (N_14444,N_11952,N_10593);
nand U14445 (N_14445,N_9074,N_8423);
xor U14446 (N_14446,N_8682,N_11847);
nor U14447 (N_14447,N_11315,N_10508);
nand U14448 (N_14448,N_10432,N_8647);
or U14449 (N_14449,N_11724,N_10320);
nand U14450 (N_14450,N_8393,N_11599);
nor U14451 (N_14451,N_9980,N_11852);
and U14452 (N_14452,N_11000,N_9913);
nor U14453 (N_14453,N_8440,N_10246);
or U14454 (N_14454,N_8483,N_11177);
and U14455 (N_14455,N_10308,N_8087);
xnor U14456 (N_14456,N_11129,N_9842);
or U14457 (N_14457,N_11374,N_10991);
nand U14458 (N_14458,N_10509,N_9478);
nor U14459 (N_14459,N_10998,N_9370);
and U14460 (N_14460,N_11824,N_8289);
nand U14461 (N_14461,N_11947,N_9952);
xnor U14462 (N_14462,N_8602,N_8497);
nand U14463 (N_14463,N_11185,N_8119);
or U14464 (N_14464,N_8768,N_11553);
or U14465 (N_14465,N_11002,N_8244);
nand U14466 (N_14466,N_11523,N_8613);
or U14467 (N_14467,N_10553,N_11843);
nor U14468 (N_14468,N_9239,N_11097);
nand U14469 (N_14469,N_11399,N_10141);
or U14470 (N_14470,N_8231,N_10564);
or U14471 (N_14471,N_9485,N_10805);
or U14472 (N_14472,N_10878,N_10801);
and U14473 (N_14473,N_11991,N_9368);
nor U14474 (N_14474,N_9785,N_11130);
or U14475 (N_14475,N_9373,N_10598);
or U14476 (N_14476,N_8495,N_8917);
or U14477 (N_14477,N_8996,N_9842);
nor U14478 (N_14478,N_11169,N_9789);
nand U14479 (N_14479,N_11605,N_11826);
and U14480 (N_14480,N_10516,N_11383);
nand U14481 (N_14481,N_10211,N_8903);
nor U14482 (N_14482,N_8031,N_10532);
or U14483 (N_14483,N_8228,N_9221);
or U14484 (N_14484,N_10827,N_8141);
nand U14485 (N_14485,N_11652,N_10078);
xor U14486 (N_14486,N_9877,N_9227);
nand U14487 (N_14487,N_11758,N_9411);
or U14488 (N_14488,N_9010,N_11989);
nor U14489 (N_14489,N_9145,N_9239);
xor U14490 (N_14490,N_11777,N_10455);
nor U14491 (N_14491,N_11028,N_8083);
and U14492 (N_14492,N_11113,N_10635);
and U14493 (N_14493,N_9046,N_9602);
nor U14494 (N_14494,N_8336,N_10302);
and U14495 (N_14495,N_9227,N_10265);
nor U14496 (N_14496,N_10858,N_10939);
nand U14497 (N_14497,N_11976,N_8516);
or U14498 (N_14498,N_8481,N_9423);
xor U14499 (N_14499,N_8105,N_10169);
or U14500 (N_14500,N_8205,N_8998);
nor U14501 (N_14501,N_9761,N_10697);
or U14502 (N_14502,N_9718,N_11299);
xnor U14503 (N_14503,N_11968,N_9261);
nand U14504 (N_14504,N_9758,N_11245);
nand U14505 (N_14505,N_9796,N_11212);
and U14506 (N_14506,N_9861,N_8502);
nand U14507 (N_14507,N_11425,N_10173);
nor U14508 (N_14508,N_9675,N_8495);
or U14509 (N_14509,N_8977,N_10278);
xnor U14510 (N_14510,N_11148,N_9038);
xnor U14511 (N_14511,N_8817,N_10943);
or U14512 (N_14512,N_10950,N_8659);
or U14513 (N_14513,N_10330,N_10094);
nor U14514 (N_14514,N_11641,N_8518);
and U14515 (N_14515,N_11552,N_9660);
nand U14516 (N_14516,N_11688,N_10433);
nand U14517 (N_14517,N_10490,N_10236);
nor U14518 (N_14518,N_10265,N_8534);
nand U14519 (N_14519,N_11624,N_9426);
nor U14520 (N_14520,N_11451,N_8535);
or U14521 (N_14521,N_8106,N_11116);
and U14522 (N_14522,N_9307,N_8851);
and U14523 (N_14523,N_11272,N_8765);
and U14524 (N_14524,N_10378,N_10863);
nor U14525 (N_14525,N_11155,N_9936);
and U14526 (N_14526,N_11980,N_11234);
nand U14527 (N_14527,N_8053,N_8805);
nor U14528 (N_14528,N_11449,N_11567);
or U14529 (N_14529,N_11767,N_8223);
and U14530 (N_14530,N_8152,N_9871);
or U14531 (N_14531,N_8989,N_10883);
nand U14532 (N_14532,N_10665,N_11984);
nor U14533 (N_14533,N_10904,N_8221);
nor U14534 (N_14534,N_8211,N_10132);
and U14535 (N_14535,N_11349,N_11523);
or U14536 (N_14536,N_8212,N_10947);
xor U14537 (N_14537,N_8647,N_10045);
or U14538 (N_14538,N_8952,N_8452);
and U14539 (N_14539,N_11978,N_8246);
or U14540 (N_14540,N_11648,N_8945);
and U14541 (N_14541,N_10527,N_9793);
and U14542 (N_14542,N_8711,N_9302);
or U14543 (N_14543,N_11880,N_9243);
nand U14544 (N_14544,N_10619,N_11388);
or U14545 (N_14545,N_8677,N_8203);
nand U14546 (N_14546,N_11368,N_11321);
nor U14547 (N_14547,N_11088,N_10926);
or U14548 (N_14548,N_10606,N_8593);
nor U14549 (N_14549,N_8623,N_8334);
or U14550 (N_14550,N_8713,N_8946);
or U14551 (N_14551,N_10192,N_8359);
nor U14552 (N_14552,N_8090,N_8469);
xnor U14553 (N_14553,N_8342,N_9806);
or U14554 (N_14554,N_8023,N_9896);
and U14555 (N_14555,N_11185,N_11613);
and U14556 (N_14556,N_9670,N_11217);
or U14557 (N_14557,N_8578,N_11988);
and U14558 (N_14558,N_10791,N_8491);
xor U14559 (N_14559,N_10562,N_9759);
nor U14560 (N_14560,N_8296,N_11415);
nor U14561 (N_14561,N_10327,N_9191);
or U14562 (N_14562,N_10165,N_11839);
and U14563 (N_14563,N_8577,N_11990);
nor U14564 (N_14564,N_11660,N_8509);
xor U14565 (N_14565,N_10150,N_8465);
and U14566 (N_14566,N_8447,N_9007);
nor U14567 (N_14567,N_11585,N_9826);
nor U14568 (N_14568,N_10259,N_8912);
or U14569 (N_14569,N_11101,N_9558);
and U14570 (N_14570,N_9850,N_8254);
and U14571 (N_14571,N_11831,N_11868);
and U14572 (N_14572,N_11929,N_9443);
xor U14573 (N_14573,N_10236,N_9032);
nand U14574 (N_14574,N_11969,N_11490);
nor U14575 (N_14575,N_9325,N_8059);
or U14576 (N_14576,N_9008,N_10330);
nand U14577 (N_14577,N_11340,N_8709);
or U14578 (N_14578,N_9145,N_10771);
nor U14579 (N_14579,N_8394,N_9780);
xnor U14580 (N_14580,N_8274,N_8153);
nand U14581 (N_14581,N_10168,N_11452);
and U14582 (N_14582,N_11801,N_8785);
and U14583 (N_14583,N_10253,N_9856);
nand U14584 (N_14584,N_9375,N_9629);
nand U14585 (N_14585,N_8352,N_9918);
xor U14586 (N_14586,N_10149,N_10132);
and U14587 (N_14587,N_8399,N_11849);
or U14588 (N_14588,N_8281,N_11611);
nor U14589 (N_14589,N_10047,N_11364);
or U14590 (N_14590,N_8339,N_8649);
nor U14591 (N_14591,N_9607,N_11112);
and U14592 (N_14592,N_10574,N_9864);
xnor U14593 (N_14593,N_9874,N_8385);
nor U14594 (N_14594,N_9173,N_11239);
and U14595 (N_14595,N_9511,N_11471);
nor U14596 (N_14596,N_9796,N_11790);
or U14597 (N_14597,N_11595,N_10568);
and U14598 (N_14598,N_10842,N_10571);
and U14599 (N_14599,N_8221,N_9140);
and U14600 (N_14600,N_11945,N_11161);
nand U14601 (N_14601,N_8881,N_11707);
or U14602 (N_14602,N_9368,N_10064);
nand U14603 (N_14603,N_8606,N_10444);
nand U14604 (N_14604,N_11507,N_10217);
and U14605 (N_14605,N_11175,N_8582);
nand U14606 (N_14606,N_9061,N_10789);
or U14607 (N_14607,N_10343,N_9560);
or U14608 (N_14608,N_8369,N_8712);
and U14609 (N_14609,N_9444,N_8097);
nand U14610 (N_14610,N_11360,N_11041);
or U14611 (N_14611,N_10321,N_9031);
and U14612 (N_14612,N_9617,N_8782);
nor U14613 (N_14613,N_11427,N_9289);
xor U14614 (N_14614,N_8528,N_8654);
or U14615 (N_14615,N_10540,N_11860);
nand U14616 (N_14616,N_11443,N_9285);
or U14617 (N_14617,N_8977,N_11638);
and U14618 (N_14618,N_10131,N_8187);
or U14619 (N_14619,N_11175,N_10709);
nor U14620 (N_14620,N_11927,N_8790);
xor U14621 (N_14621,N_11321,N_10758);
xor U14622 (N_14622,N_10933,N_10687);
and U14623 (N_14623,N_10640,N_9033);
xnor U14624 (N_14624,N_10057,N_8396);
or U14625 (N_14625,N_9485,N_9351);
nand U14626 (N_14626,N_8507,N_8949);
or U14627 (N_14627,N_9759,N_10669);
and U14628 (N_14628,N_8677,N_8273);
nand U14629 (N_14629,N_8685,N_9258);
nor U14630 (N_14630,N_9809,N_9177);
nor U14631 (N_14631,N_9179,N_11702);
nor U14632 (N_14632,N_10327,N_8239);
xor U14633 (N_14633,N_8056,N_9686);
or U14634 (N_14634,N_10972,N_10515);
or U14635 (N_14635,N_8528,N_11811);
or U14636 (N_14636,N_11362,N_11054);
or U14637 (N_14637,N_10816,N_9038);
nor U14638 (N_14638,N_10716,N_9538);
or U14639 (N_14639,N_11187,N_10960);
or U14640 (N_14640,N_8072,N_8112);
nand U14641 (N_14641,N_10731,N_11841);
nand U14642 (N_14642,N_11483,N_9423);
and U14643 (N_14643,N_9115,N_8943);
nand U14644 (N_14644,N_10051,N_9264);
nand U14645 (N_14645,N_8411,N_8125);
and U14646 (N_14646,N_9478,N_10529);
or U14647 (N_14647,N_8474,N_9620);
and U14648 (N_14648,N_8242,N_10272);
nand U14649 (N_14649,N_9947,N_8223);
nor U14650 (N_14650,N_8239,N_10633);
and U14651 (N_14651,N_8247,N_8630);
and U14652 (N_14652,N_9083,N_10498);
nand U14653 (N_14653,N_10774,N_10866);
nand U14654 (N_14654,N_9746,N_9620);
and U14655 (N_14655,N_9436,N_11765);
and U14656 (N_14656,N_11439,N_9207);
xor U14657 (N_14657,N_11619,N_8680);
nand U14658 (N_14658,N_8490,N_11843);
and U14659 (N_14659,N_10930,N_9302);
nor U14660 (N_14660,N_9341,N_10066);
nand U14661 (N_14661,N_9438,N_11385);
or U14662 (N_14662,N_10223,N_8810);
and U14663 (N_14663,N_9561,N_9699);
nor U14664 (N_14664,N_10494,N_8796);
nor U14665 (N_14665,N_11965,N_8181);
or U14666 (N_14666,N_11580,N_10999);
nand U14667 (N_14667,N_10458,N_10766);
or U14668 (N_14668,N_8909,N_11587);
nor U14669 (N_14669,N_11872,N_9853);
or U14670 (N_14670,N_10653,N_9450);
xor U14671 (N_14671,N_11256,N_8619);
nand U14672 (N_14672,N_11973,N_10142);
and U14673 (N_14673,N_11106,N_10680);
xor U14674 (N_14674,N_8828,N_11779);
nor U14675 (N_14675,N_9263,N_11220);
or U14676 (N_14676,N_9443,N_10396);
or U14677 (N_14677,N_11672,N_9136);
or U14678 (N_14678,N_10918,N_11829);
or U14679 (N_14679,N_8036,N_9906);
or U14680 (N_14680,N_11152,N_10142);
or U14681 (N_14681,N_11534,N_9320);
nor U14682 (N_14682,N_11017,N_11352);
nand U14683 (N_14683,N_10183,N_8912);
nor U14684 (N_14684,N_8342,N_8161);
nand U14685 (N_14685,N_8033,N_9438);
xor U14686 (N_14686,N_10979,N_11677);
nand U14687 (N_14687,N_10530,N_9151);
or U14688 (N_14688,N_8173,N_9992);
and U14689 (N_14689,N_11593,N_9638);
and U14690 (N_14690,N_10753,N_8205);
or U14691 (N_14691,N_8354,N_10332);
and U14692 (N_14692,N_8144,N_9842);
nor U14693 (N_14693,N_10543,N_11307);
and U14694 (N_14694,N_11121,N_11135);
nor U14695 (N_14695,N_10478,N_10421);
nand U14696 (N_14696,N_9323,N_8161);
nor U14697 (N_14697,N_11967,N_8009);
nand U14698 (N_14698,N_9465,N_9505);
or U14699 (N_14699,N_8449,N_10556);
nor U14700 (N_14700,N_8232,N_10847);
nor U14701 (N_14701,N_8480,N_8826);
or U14702 (N_14702,N_10132,N_10024);
nand U14703 (N_14703,N_9250,N_11446);
or U14704 (N_14704,N_8651,N_11461);
or U14705 (N_14705,N_10850,N_8795);
nor U14706 (N_14706,N_9913,N_11764);
nand U14707 (N_14707,N_9932,N_9382);
or U14708 (N_14708,N_9056,N_8863);
xnor U14709 (N_14709,N_9443,N_11451);
nor U14710 (N_14710,N_10199,N_11897);
nand U14711 (N_14711,N_9147,N_8610);
and U14712 (N_14712,N_11799,N_8258);
and U14713 (N_14713,N_9681,N_10864);
or U14714 (N_14714,N_8103,N_10820);
nor U14715 (N_14715,N_9302,N_11120);
nor U14716 (N_14716,N_8514,N_8759);
nand U14717 (N_14717,N_9156,N_9973);
nand U14718 (N_14718,N_11729,N_9802);
nand U14719 (N_14719,N_8980,N_10152);
or U14720 (N_14720,N_9311,N_9415);
and U14721 (N_14721,N_10852,N_9991);
or U14722 (N_14722,N_10197,N_9397);
and U14723 (N_14723,N_10748,N_9985);
nor U14724 (N_14724,N_9902,N_8828);
or U14725 (N_14725,N_11347,N_8209);
nor U14726 (N_14726,N_8177,N_8738);
and U14727 (N_14727,N_8080,N_10863);
nand U14728 (N_14728,N_11799,N_8427);
and U14729 (N_14729,N_10373,N_8308);
nor U14730 (N_14730,N_11380,N_8103);
xor U14731 (N_14731,N_10270,N_8095);
or U14732 (N_14732,N_9081,N_9355);
nor U14733 (N_14733,N_9154,N_8882);
or U14734 (N_14734,N_10520,N_10644);
or U14735 (N_14735,N_11318,N_10309);
and U14736 (N_14736,N_9027,N_9570);
nand U14737 (N_14737,N_8110,N_8156);
nor U14738 (N_14738,N_9492,N_10083);
or U14739 (N_14739,N_8033,N_10361);
or U14740 (N_14740,N_9349,N_8089);
and U14741 (N_14741,N_9534,N_11189);
nor U14742 (N_14742,N_9771,N_11138);
xor U14743 (N_14743,N_9146,N_8471);
or U14744 (N_14744,N_8323,N_8201);
nand U14745 (N_14745,N_10070,N_8477);
or U14746 (N_14746,N_8665,N_10972);
nor U14747 (N_14747,N_8860,N_8226);
nor U14748 (N_14748,N_11543,N_11593);
or U14749 (N_14749,N_8047,N_11092);
and U14750 (N_14750,N_11817,N_8266);
nor U14751 (N_14751,N_10489,N_11250);
or U14752 (N_14752,N_8669,N_11815);
and U14753 (N_14753,N_9808,N_8077);
xnor U14754 (N_14754,N_11354,N_10381);
or U14755 (N_14755,N_8378,N_8359);
and U14756 (N_14756,N_9693,N_10493);
and U14757 (N_14757,N_9422,N_8295);
and U14758 (N_14758,N_9694,N_11421);
or U14759 (N_14759,N_10497,N_8852);
or U14760 (N_14760,N_8512,N_8577);
and U14761 (N_14761,N_11020,N_9234);
or U14762 (N_14762,N_8411,N_8934);
nand U14763 (N_14763,N_9749,N_8355);
nand U14764 (N_14764,N_10764,N_10579);
nand U14765 (N_14765,N_9604,N_10209);
or U14766 (N_14766,N_10677,N_10514);
and U14767 (N_14767,N_8472,N_9073);
xor U14768 (N_14768,N_8454,N_9224);
nor U14769 (N_14769,N_8763,N_10200);
and U14770 (N_14770,N_9292,N_9587);
and U14771 (N_14771,N_9310,N_11695);
or U14772 (N_14772,N_8402,N_8134);
or U14773 (N_14773,N_10505,N_8628);
nor U14774 (N_14774,N_9627,N_10263);
nand U14775 (N_14775,N_8387,N_11217);
or U14776 (N_14776,N_8531,N_10299);
and U14777 (N_14777,N_8589,N_10874);
or U14778 (N_14778,N_8186,N_9002);
nand U14779 (N_14779,N_10664,N_10819);
nor U14780 (N_14780,N_10084,N_9477);
or U14781 (N_14781,N_10292,N_8139);
and U14782 (N_14782,N_10725,N_9678);
nor U14783 (N_14783,N_11778,N_10510);
or U14784 (N_14784,N_10292,N_9446);
xnor U14785 (N_14785,N_9704,N_11867);
nand U14786 (N_14786,N_10476,N_9585);
and U14787 (N_14787,N_10070,N_11371);
or U14788 (N_14788,N_8869,N_8349);
or U14789 (N_14789,N_9639,N_11509);
nand U14790 (N_14790,N_8539,N_10350);
nor U14791 (N_14791,N_9340,N_10930);
nor U14792 (N_14792,N_9975,N_11085);
nand U14793 (N_14793,N_8987,N_9530);
nor U14794 (N_14794,N_10517,N_10754);
nand U14795 (N_14795,N_11759,N_10991);
nor U14796 (N_14796,N_11360,N_9370);
or U14797 (N_14797,N_10807,N_8016);
or U14798 (N_14798,N_9728,N_11278);
or U14799 (N_14799,N_11229,N_9779);
nand U14800 (N_14800,N_8576,N_8992);
nand U14801 (N_14801,N_9174,N_9786);
nor U14802 (N_14802,N_8582,N_8713);
nand U14803 (N_14803,N_9418,N_10855);
nor U14804 (N_14804,N_9803,N_11577);
nand U14805 (N_14805,N_8963,N_10542);
nand U14806 (N_14806,N_8921,N_10132);
and U14807 (N_14807,N_9876,N_11590);
nand U14808 (N_14808,N_11277,N_9235);
nor U14809 (N_14809,N_10965,N_10191);
nand U14810 (N_14810,N_9762,N_9740);
nor U14811 (N_14811,N_10689,N_8735);
or U14812 (N_14812,N_11702,N_8148);
xor U14813 (N_14813,N_8249,N_10445);
nor U14814 (N_14814,N_10075,N_11809);
or U14815 (N_14815,N_11996,N_9558);
and U14816 (N_14816,N_10228,N_9775);
nand U14817 (N_14817,N_10840,N_11678);
nand U14818 (N_14818,N_11291,N_8541);
and U14819 (N_14819,N_11368,N_8278);
and U14820 (N_14820,N_8303,N_8212);
and U14821 (N_14821,N_9021,N_11133);
or U14822 (N_14822,N_8008,N_8171);
nor U14823 (N_14823,N_8997,N_11834);
and U14824 (N_14824,N_10303,N_11183);
nor U14825 (N_14825,N_8181,N_8695);
nand U14826 (N_14826,N_10761,N_10934);
xnor U14827 (N_14827,N_10485,N_10462);
nand U14828 (N_14828,N_11929,N_8705);
nor U14829 (N_14829,N_10756,N_9109);
xnor U14830 (N_14830,N_10165,N_9010);
nand U14831 (N_14831,N_8858,N_10234);
nor U14832 (N_14832,N_8167,N_8571);
and U14833 (N_14833,N_8278,N_10948);
nand U14834 (N_14834,N_9478,N_11911);
nand U14835 (N_14835,N_8193,N_11335);
nor U14836 (N_14836,N_9386,N_11849);
and U14837 (N_14837,N_9291,N_9729);
and U14838 (N_14838,N_8223,N_11164);
or U14839 (N_14839,N_8683,N_11370);
nor U14840 (N_14840,N_10576,N_10170);
nand U14841 (N_14841,N_10635,N_11918);
nand U14842 (N_14842,N_10777,N_8318);
nor U14843 (N_14843,N_10250,N_11698);
or U14844 (N_14844,N_8730,N_9047);
or U14845 (N_14845,N_10362,N_11498);
xnor U14846 (N_14846,N_11959,N_8811);
nor U14847 (N_14847,N_9693,N_10518);
nor U14848 (N_14848,N_8659,N_10167);
nor U14849 (N_14849,N_8070,N_10181);
or U14850 (N_14850,N_8161,N_11519);
or U14851 (N_14851,N_11564,N_10638);
nor U14852 (N_14852,N_8427,N_11152);
xor U14853 (N_14853,N_11745,N_10765);
nand U14854 (N_14854,N_11639,N_11090);
nand U14855 (N_14855,N_11446,N_8229);
xnor U14856 (N_14856,N_9106,N_10285);
or U14857 (N_14857,N_11991,N_9054);
nand U14858 (N_14858,N_9221,N_11501);
nor U14859 (N_14859,N_11293,N_9181);
or U14860 (N_14860,N_8200,N_8992);
nand U14861 (N_14861,N_10233,N_10604);
and U14862 (N_14862,N_10983,N_8935);
nor U14863 (N_14863,N_10543,N_8638);
and U14864 (N_14864,N_10204,N_8630);
and U14865 (N_14865,N_11696,N_11185);
xor U14866 (N_14866,N_9045,N_11363);
nor U14867 (N_14867,N_9601,N_9579);
nand U14868 (N_14868,N_9492,N_8311);
and U14869 (N_14869,N_8161,N_9435);
xnor U14870 (N_14870,N_10974,N_10999);
nor U14871 (N_14871,N_10044,N_10880);
or U14872 (N_14872,N_10235,N_10230);
and U14873 (N_14873,N_10081,N_9616);
nor U14874 (N_14874,N_9785,N_9873);
nand U14875 (N_14875,N_9367,N_8416);
or U14876 (N_14876,N_8327,N_9010);
or U14877 (N_14877,N_8929,N_9208);
nand U14878 (N_14878,N_9868,N_11449);
or U14879 (N_14879,N_11220,N_11839);
nand U14880 (N_14880,N_10212,N_11885);
or U14881 (N_14881,N_9987,N_11650);
nor U14882 (N_14882,N_10823,N_9294);
and U14883 (N_14883,N_8068,N_8387);
and U14884 (N_14884,N_9725,N_11895);
nand U14885 (N_14885,N_10267,N_8934);
xor U14886 (N_14886,N_8700,N_9357);
nor U14887 (N_14887,N_8590,N_8836);
nor U14888 (N_14888,N_8322,N_10602);
nor U14889 (N_14889,N_8442,N_10750);
or U14890 (N_14890,N_11052,N_10802);
nand U14891 (N_14891,N_8915,N_9665);
nand U14892 (N_14892,N_9192,N_11634);
or U14893 (N_14893,N_11940,N_9982);
nand U14894 (N_14894,N_10900,N_9650);
nor U14895 (N_14895,N_8290,N_10796);
nand U14896 (N_14896,N_10117,N_11525);
xnor U14897 (N_14897,N_8222,N_10944);
nor U14898 (N_14898,N_11545,N_10990);
xnor U14899 (N_14899,N_9056,N_11313);
and U14900 (N_14900,N_8132,N_8952);
nor U14901 (N_14901,N_8665,N_8255);
nor U14902 (N_14902,N_8245,N_9099);
nand U14903 (N_14903,N_9577,N_11355);
or U14904 (N_14904,N_8156,N_10171);
nor U14905 (N_14905,N_9733,N_11135);
nor U14906 (N_14906,N_9739,N_8875);
nand U14907 (N_14907,N_8883,N_11206);
nand U14908 (N_14908,N_9059,N_10849);
nor U14909 (N_14909,N_10324,N_8323);
nand U14910 (N_14910,N_10293,N_9065);
nand U14911 (N_14911,N_11503,N_9691);
or U14912 (N_14912,N_8699,N_11144);
nand U14913 (N_14913,N_9904,N_9869);
nand U14914 (N_14914,N_10990,N_10724);
or U14915 (N_14915,N_10412,N_10633);
and U14916 (N_14916,N_11569,N_8953);
nand U14917 (N_14917,N_11805,N_11161);
nor U14918 (N_14918,N_11130,N_8025);
nor U14919 (N_14919,N_10339,N_8640);
and U14920 (N_14920,N_9841,N_9923);
or U14921 (N_14921,N_9272,N_9485);
xor U14922 (N_14922,N_9357,N_9577);
and U14923 (N_14923,N_10755,N_9374);
xnor U14924 (N_14924,N_8062,N_11581);
nand U14925 (N_14925,N_10553,N_9274);
xor U14926 (N_14926,N_10681,N_9650);
nor U14927 (N_14927,N_10326,N_10047);
nand U14928 (N_14928,N_9293,N_11640);
nand U14929 (N_14929,N_9119,N_8596);
xnor U14930 (N_14930,N_11899,N_9779);
nand U14931 (N_14931,N_8318,N_11496);
nor U14932 (N_14932,N_10154,N_9446);
or U14933 (N_14933,N_11475,N_8530);
xnor U14934 (N_14934,N_11800,N_8556);
and U14935 (N_14935,N_10352,N_8330);
xnor U14936 (N_14936,N_8791,N_10041);
nand U14937 (N_14937,N_11758,N_10542);
nor U14938 (N_14938,N_10956,N_10628);
and U14939 (N_14939,N_8940,N_11387);
or U14940 (N_14940,N_10930,N_11862);
and U14941 (N_14941,N_10770,N_10372);
nand U14942 (N_14942,N_9341,N_11031);
nor U14943 (N_14943,N_8091,N_11517);
or U14944 (N_14944,N_10087,N_9798);
or U14945 (N_14945,N_9968,N_9583);
or U14946 (N_14946,N_8865,N_10096);
nand U14947 (N_14947,N_8392,N_9778);
or U14948 (N_14948,N_11936,N_10890);
xor U14949 (N_14949,N_9175,N_10141);
nand U14950 (N_14950,N_8938,N_8433);
and U14951 (N_14951,N_11010,N_8365);
nor U14952 (N_14952,N_11255,N_8972);
nor U14953 (N_14953,N_11138,N_10584);
nor U14954 (N_14954,N_11729,N_10812);
and U14955 (N_14955,N_9397,N_8159);
nor U14956 (N_14956,N_8809,N_10667);
xor U14957 (N_14957,N_9674,N_10222);
and U14958 (N_14958,N_8103,N_8255);
and U14959 (N_14959,N_10324,N_11352);
or U14960 (N_14960,N_10664,N_10568);
nor U14961 (N_14961,N_9740,N_9027);
or U14962 (N_14962,N_11137,N_10685);
and U14963 (N_14963,N_10580,N_9471);
or U14964 (N_14964,N_8041,N_10890);
nor U14965 (N_14965,N_9939,N_10267);
nand U14966 (N_14966,N_8972,N_11857);
nand U14967 (N_14967,N_9612,N_8124);
xnor U14968 (N_14968,N_9336,N_10292);
nor U14969 (N_14969,N_8231,N_10499);
nor U14970 (N_14970,N_10318,N_10899);
or U14971 (N_14971,N_9434,N_8694);
and U14972 (N_14972,N_11129,N_11317);
nand U14973 (N_14973,N_10872,N_8444);
nor U14974 (N_14974,N_11920,N_9322);
and U14975 (N_14975,N_9405,N_11507);
nor U14976 (N_14976,N_11972,N_8375);
nor U14977 (N_14977,N_9667,N_9755);
nor U14978 (N_14978,N_9733,N_10668);
or U14979 (N_14979,N_9035,N_9062);
or U14980 (N_14980,N_11255,N_11567);
nor U14981 (N_14981,N_9826,N_9818);
xor U14982 (N_14982,N_11709,N_10414);
or U14983 (N_14983,N_10079,N_8168);
nor U14984 (N_14984,N_9995,N_10248);
nor U14985 (N_14985,N_8508,N_9596);
nand U14986 (N_14986,N_9102,N_10713);
nor U14987 (N_14987,N_11153,N_10086);
or U14988 (N_14988,N_11115,N_8337);
nor U14989 (N_14989,N_9292,N_10363);
and U14990 (N_14990,N_10158,N_10867);
nor U14991 (N_14991,N_9583,N_10285);
nor U14992 (N_14992,N_8973,N_9063);
and U14993 (N_14993,N_11589,N_10054);
nor U14994 (N_14994,N_10213,N_8739);
xnor U14995 (N_14995,N_8450,N_9199);
and U14996 (N_14996,N_8727,N_10264);
nor U14997 (N_14997,N_8299,N_8398);
nor U14998 (N_14998,N_8923,N_11139);
nand U14999 (N_14999,N_11365,N_11930);
and U15000 (N_15000,N_9341,N_8905);
or U15001 (N_15001,N_9422,N_8806);
xor U15002 (N_15002,N_11124,N_11773);
nor U15003 (N_15003,N_9224,N_10949);
or U15004 (N_15004,N_9784,N_9160);
nor U15005 (N_15005,N_8145,N_9347);
or U15006 (N_15006,N_8633,N_8339);
and U15007 (N_15007,N_9152,N_11239);
nor U15008 (N_15008,N_8220,N_11527);
and U15009 (N_15009,N_8326,N_11464);
xnor U15010 (N_15010,N_11007,N_10050);
nand U15011 (N_15011,N_10379,N_9921);
nand U15012 (N_15012,N_11191,N_8469);
nand U15013 (N_15013,N_8505,N_11480);
or U15014 (N_15014,N_8822,N_10283);
and U15015 (N_15015,N_8115,N_10036);
xnor U15016 (N_15016,N_9999,N_8618);
or U15017 (N_15017,N_9367,N_9238);
nor U15018 (N_15018,N_8637,N_11936);
and U15019 (N_15019,N_11908,N_8855);
nand U15020 (N_15020,N_11776,N_10230);
and U15021 (N_15021,N_8115,N_10232);
xnor U15022 (N_15022,N_9551,N_9165);
or U15023 (N_15023,N_10064,N_8087);
nand U15024 (N_15024,N_10457,N_8239);
nand U15025 (N_15025,N_10506,N_8945);
xnor U15026 (N_15026,N_9221,N_11206);
nand U15027 (N_15027,N_8929,N_8752);
nand U15028 (N_15028,N_9307,N_8087);
nand U15029 (N_15029,N_8334,N_9132);
xor U15030 (N_15030,N_10913,N_8363);
or U15031 (N_15031,N_11194,N_8448);
nand U15032 (N_15032,N_10223,N_11645);
or U15033 (N_15033,N_11681,N_9377);
nor U15034 (N_15034,N_10572,N_8933);
nand U15035 (N_15035,N_8174,N_10319);
and U15036 (N_15036,N_8605,N_8880);
xor U15037 (N_15037,N_11501,N_11123);
and U15038 (N_15038,N_11884,N_10579);
and U15039 (N_15039,N_11055,N_10059);
nor U15040 (N_15040,N_9102,N_8070);
and U15041 (N_15041,N_9854,N_10708);
and U15042 (N_15042,N_11072,N_9420);
xor U15043 (N_15043,N_8046,N_9139);
or U15044 (N_15044,N_10369,N_9264);
nor U15045 (N_15045,N_10681,N_10989);
or U15046 (N_15046,N_8949,N_11645);
and U15047 (N_15047,N_8089,N_9485);
and U15048 (N_15048,N_9171,N_10055);
and U15049 (N_15049,N_10997,N_11880);
or U15050 (N_15050,N_8603,N_11284);
and U15051 (N_15051,N_8496,N_9704);
or U15052 (N_15052,N_11933,N_10174);
nand U15053 (N_15053,N_11163,N_9084);
and U15054 (N_15054,N_11934,N_8848);
and U15055 (N_15055,N_10524,N_9020);
and U15056 (N_15056,N_10396,N_9068);
or U15057 (N_15057,N_9724,N_10323);
or U15058 (N_15058,N_11880,N_9294);
or U15059 (N_15059,N_10514,N_9676);
or U15060 (N_15060,N_9434,N_10940);
or U15061 (N_15061,N_10339,N_8587);
nor U15062 (N_15062,N_11353,N_11940);
nand U15063 (N_15063,N_11376,N_8496);
xnor U15064 (N_15064,N_11463,N_9557);
nand U15065 (N_15065,N_10322,N_11443);
nor U15066 (N_15066,N_9089,N_11937);
nand U15067 (N_15067,N_11310,N_10316);
or U15068 (N_15068,N_10442,N_9797);
nand U15069 (N_15069,N_8280,N_9712);
nor U15070 (N_15070,N_9504,N_9624);
nand U15071 (N_15071,N_9748,N_8679);
nand U15072 (N_15072,N_11862,N_9989);
or U15073 (N_15073,N_11870,N_10122);
nand U15074 (N_15074,N_11280,N_8413);
nand U15075 (N_15075,N_10854,N_10245);
or U15076 (N_15076,N_10508,N_11928);
and U15077 (N_15077,N_11688,N_11205);
nor U15078 (N_15078,N_10331,N_10672);
xnor U15079 (N_15079,N_9180,N_11756);
and U15080 (N_15080,N_8008,N_10495);
nor U15081 (N_15081,N_8158,N_9252);
nand U15082 (N_15082,N_8518,N_9958);
xnor U15083 (N_15083,N_10605,N_11593);
or U15084 (N_15084,N_9363,N_8076);
nor U15085 (N_15085,N_11193,N_11039);
nand U15086 (N_15086,N_10250,N_8077);
xor U15087 (N_15087,N_9828,N_9778);
and U15088 (N_15088,N_11819,N_9120);
nand U15089 (N_15089,N_11784,N_10654);
nand U15090 (N_15090,N_11644,N_8687);
nand U15091 (N_15091,N_9312,N_9859);
nor U15092 (N_15092,N_11010,N_9543);
nor U15093 (N_15093,N_9800,N_11525);
and U15094 (N_15094,N_10886,N_9071);
xnor U15095 (N_15095,N_8527,N_11753);
or U15096 (N_15096,N_11639,N_10801);
or U15097 (N_15097,N_11938,N_10995);
or U15098 (N_15098,N_8140,N_8083);
nor U15099 (N_15099,N_8879,N_8433);
or U15100 (N_15100,N_11112,N_10361);
or U15101 (N_15101,N_9114,N_11943);
nand U15102 (N_15102,N_9089,N_11688);
nand U15103 (N_15103,N_9486,N_11458);
and U15104 (N_15104,N_8519,N_11404);
or U15105 (N_15105,N_8676,N_9169);
and U15106 (N_15106,N_9611,N_9016);
and U15107 (N_15107,N_8524,N_9903);
xnor U15108 (N_15108,N_11270,N_8596);
and U15109 (N_15109,N_8519,N_11311);
and U15110 (N_15110,N_8216,N_11871);
nand U15111 (N_15111,N_8005,N_10150);
or U15112 (N_15112,N_9064,N_9444);
nor U15113 (N_15113,N_10536,N_10736);
or U15114 (N_15114,N_10809,N_9370);
xor U15115 (N_15115,N_8440,N_8890);
nor U15116 (N_15116,N_9540,N_10693);
or U15117 (N_15117,N_11495,N_10829);
nand U15118 (N_15118,N_8602,N_10037);
nor U15119 (N_15119,N_10203,N_11844);
and U15120 (N_15120,N_11303,N_9594);
or U15121 (N_15121,N_9496,N_10222);
nor U15122 (N_15122,N_10556,N_11662);
and U15123 (N_15123,N_9310,N_9900);
or U15124 (N_15124,N_11333,N_10418);
nand U15125 (N_15125,N_9458,N_10317);
xnor U15126 (N_15126,N_9062,N_10518);
xnor U15127 (N_15127,N_8648,N_8302);
or U15128 (N_15128,N_9829,N_8994);
and U15129 (N_15129,N_10549,N_9134);
nand U15130 (N_15130,N_8129,N_9557);
nor U15131 (N_15131,N_9482,N_8199);
and U15132 (N_15132,N_10723,N_11314);
or U15133 (N_15133,N_11571,N_10456);
nor U15134 (N_15134,N_10164,N_10534);
nand U15135 (N_15135,N_11866,N_11849);
and U15136 (N_15136,N_11378,N_8964);
and U15137 (N_15137,N_11777,N_9144);
or U15138 (N_15138,N_11606,N_9258);
nand U15139 (N_15139,N_9503,N_8031);
nor U15140 (N_15140,N_9228,N_11701);
and U15141 (N_15141,N_9194,N_8387);
nor U15142 (N_15142,N_9203,N_8265);
or U15143 (N_15143,N_8611,N_8520);
xnor U15144 (N_15144,N_10905,N_11735);
xor U15145 (N_15145,N_11883,N_8027);
nand U15146 (N_15146,N_9504,N_9662);
nor U15147 (N_15147,N_8736,N_11173);
and U15148 (N_15148,N_11438,N_8808);
and U15149 (N_15149,N_8571,N_8649);
nor U15150 (N_15150,N_10722,N_8933);
and U15151 (N_15151,N_10068,N_11872);
and U15152 (N_15152,N_11984,N_10896);
nor U15153 (N_15153,N_9377,N_11115);
nor U15154 (N_15154,N_9010,N_11478);
nor U15155 (N_15155,N_10915,N_9757);
or U15156 (N_15156,N_8312,N_8135);
xnor U15157 (N_15157,N_8091,N_9641);
nand U15158 (N_15158,N_11766,N_11197);
nand U15159 (N_15159,N_11440,N_8057);
nor U15160 (N_15160,N_10549,N_11422);
nand U15161 (N_15161,N_9646,N_8610);
or U15162 (N_15162,N_9551,N_9322);
nand U15163 (N_15163,N_9228,N_10456);
xor U15164 (N_15164,N_11504,N_8553);
nand U15165 (N_15165,N_9261,N_11662);
and U15166 (N_15166,N_10272,N_11681);
nand U15167 (N_15167,N_10770,N_8158);
nand U15168 (N_15168,N_10074,N_9275);
nand U15169 (N_15169,N_10262,N_10067);
and U15170 (N_15170,N_10088,N_9729);
nor U15171 (N_15171,N_8816,N_9954);
or U15172 (N_15172,N_8783,N_8672);
and U15173 (N_15173,N_8440,N_11022);
or U15174 (N_15174,N_8349,N_11612);
nor U15175 (N_15175,N_8004,N_11846);
and U15176 (N_15176,N_10799,N_10312);
and U15177 (N_15177,N_9486,N_11538);
and U15178 (N_15178,N_8734,N_9505);
nor U15179 (N_15179,N_10891,N_11562);
xnor U15180 (N_15180,N_9936,N_8096);
or U15181 (N_15181,N_10212,N_10883);
or U15182 (N_15182,N_11146,N_9416);
nand U15183 (N_15183,N_11792,N_9312);
nor U15184 (N_15184,N_8381,N_10227);
and U15185 (N_15185,N_9596,N_9266);
nor U15186 (N_15186,N_10011,N_11674);
nor U15187 (N_15187,N_8530,N_10474);
nand U15188 (N_15188,N_8123,N_10996);
nor U15189 (N_15189,N_10710,N_11113);
nand U15190 (N_15190,N_10490,N_10405);
nand U15191 (N_15191,N_10902,N_8973);
or U15192 (N_15192,N_10648,N_10779);
and U15193 (N_15193,N_11446,N_9593);
and U15194 (N_15194,N_11050,N_10387);
or U15195 (N_15195,N_8177,N_10064);
xnor U15196 (N_15196,N_10827,N_11902);
nor U15197 (N_15197,N_11596,N_11713);
nand U15198 (N_15198,N_10908,N_8158);
xor U15199 (N_15199,N_9297,N_9020);
nor U15200 (N_15200,N_8988,N_9460);
nor U15201 (N_15201,N_10046,N_9927);
nand U15202 (N_15202,N_9770,N_11119);
or U15203 (N_15203,N_9300,N_11755);
and U15204 (N_15204,N_9417,N_9486);
nor U15205 (N_15205,N_9529,N_9894);
nor U15206 (N_15206,N_10965,N_9664);
nor U15207 (N_15207,N_8652,N_11441);
or U15208 (N_15208,N_10816,N_10697);
nand U15209 (N_15209,N_11303,N_10580);
and U15210 (N_15210,N_11198,N_8639);
or U15211 (N_15211,N_9024,N_10710);
xor U15212 (N_15212,N_9945,N_9468);
nand U15213 (N_15213,N_8529,N_11370);
nand U15214 (N_15214,N_8452,N_8665);
nor U15215 (N_15215,N_8325,N_10654);
nor U15216 (N_15216,N_11518,N_10228);
nor U15217 (N_15217,N_11188,N_10596);
or U15218 (N_15218,N_10205,N_10422);
nand U15219 (N_15219,N_8642,N_11300);
nor U15220 (N_15220,N_8101,N_9481);
or U15221 (N_15221,N_8138,N_9020);
nand U15222 (N_15222,N_8064,N_11113);
and U15223 (N_15223,N_11011,N_11187);
and U15224 (N_15224,N_9769,N_10415);
nor U15225 (N_15225,N_8999,N_10162);
and U15226 (N_15226,N_8315,N_9061);
and U15227 (N_15227,N_11331,N_10040);
nor U15228 (N_15228,N_10630,N_9147);
nor U15229 (N_15229,N_9366,N_11197);
nor U15230 (N_15230,N_9327,N_11299);
and U15231 (N_15231,N_9537,N_9810);
nand U15232 (N_15232,N_9531,N_11614);
nor U15233 (N_15233,N_11666,N_10250);
nor U15234 (N_15234,N_8667,N_10352);
and U15235 (N_15235,N_11405,N_8327);
or U15236 (N_15236,N_9328,N_8484);
nand U15237 (N_15237,N_8766,N_11053);
nand U15238 (N_15238,N_10194,N_8842);
or U15239 (N_15239,N_11895,N_11880);
nand U15240 (N_15240,N_9963,N_10038);
and U15241 (N_15241,N_11759,N_8194);
nor U15242 (N_15242,N_11169,N_10502);
nor U15243 (N_15243,N_9237,N_8895);
nand U15244 (N_15244,N_9466,N_9983);
nor U15245 (N_15245,N_8482,N_8909);
nor U15246 (N_15246,N_10562,N_9761);
nor U15247 (N_15247,N_10183,N_10444);
nand U15248 (N_15248,N_9851,N_10742);
or U15249 (N_15249,N_11631,N_9786);
and U15250 (N_15250,N_11486,N_10585);
xnor U15251 (N_15251,N_11921,N_9023);
and U15252 (N_15252,N_9379,N_8357);
or U15253 (N_15253,N_8377,N_8689);
nand U15254 (N_15254,N_11845,N_10764);
and U15255 (N_15255,N_10337,N_11439);
and U15256 (N_15256,N_10876,N_9703);
and U15257 (N_15257,N_8305,N_9070);
xnor U15258 (N_15258,N_9464,N_8522);
or U15259 (N_15259,N_9643,N_10346);
or U15260 (N_15260,N_8947,N_10346);
and U15261 (N_15261,N_8549,N_8258);
nor U15262 (N_15262,N_10366,N_9437);
nor U15263 (N_15263,N_10508,N_11591);
or U15264 (N_15264,N_11627,N_8349);
xnor U15265 (N_15265,N_10633,N_8572);
or U15266 (N_15266,N_8197,N_11753);
nand U15267 (N_15267,N_9152,N_8924);
or U15268 (N_15268,N_10189,N_8432);
xor U15269 (N_15269,N_11936,N_10673);
nor U15270 (N_15270,N_9734,N_9604);
or U15271 (N_15271,N_8300,N_10451);
nand U15272 (N_15272,N_11249,N_8760);
nor U15273 (N_15273,N_9604,N_10855);
or U15274 (N_15274,N_8689,N_9289);
or U15275 (N_15275,N_11487,N_9968);
nor U15276 (N_15276,N_8903,N_8082);
xnor U15277 (N_15277,N_10572,N_11886);
and U15278 (N_15278,N_9129,N_11876);
nand U15279 (N_15279,N_9478,N_11393);
nand U15280 (N_15280,N_8342,N_10568);
or U15281 (N_15281,N_11404,N_9600);
nand U15282 (N_15282,N_10896,N_9095);
and U15283 (N_15283,N_10339,N_11574);
nor U15284 (N_15284,N_11553,N_11888);
nor U15285 (N_15285,N_10161,N_10693);
or U15286 (N_15286,N_10183,N_9502);
nor U15287 (N_15287,N_8658,N_10367);
and U15288 (N_15288,N_8558,N_11629);
and U15289 (N_15289,N_10585,N_11596);
or U15290 (N_15290,N_10599,N_11302);
and U15291 (N_15291,N_9662,N_10374);
and U15292 (N_15292,N_8641,N_10319);
nand U15293 (N_15293,N_11919,N_10588);
nor U15294 (N_15294,N_10096,N_10712);
or U15295 (N_15295,N_11321,N_10799);
nor U15296 (N_15296,N_9791,N_9584);
and U15297 (N_15297,N_11480,N_11496);
nor U15298 (N_15298,N_9486,N_9992);
xnor U15299 (N_15299,N_9099,N_9521);
or U15300 (N_15300,N_11694,N_8577);
nor U15301 (N_15301,N_10635,N_10515);
or U15302 (N_15302,N_9812,N_9920);
and U15303 (N_15303,N_11983,N_8522);
xnor U15304 (N_15304,N_10394,N_9596);
or U15305 (N_15305,N_8932,N_10226);
nor U15306 (N_15306,N_11198,N_9220);
xor U15307 (N_15307,N_11022,N_11039);
and U15308 (N_15308,N_10790,N_9785);
and U15309 (N_15309,N_8457,N_11828);
nand U15310 (N_15310,N_9294,N_9326);
nor U15311 (N_15311,N_11911,N_11306);
nand U15312 (N_15312,N_11155,N_11555);
and U15313 (N_15313,N_11260,N_8839);
nand U15314 (N_15314,N_10396,N_11137);
nor U15315 (N_15315,N_11133,N_8658);
or U15316 (N_15316,N_11173,N_11976);
or U15317 (N_15317,N_11039,N_11937);
and U15318 (N_15318,N_10238,N_9637);
xor U15319 (N_15319,N_10454,N_10585);
or U15320 (N_15320,N_8468,N_10109);
or U15321 (N_15321,N_10009,N_11585);
nand U15322 (N_15322,N_11274,N_9695);
or U15323 (N_15323,N_10986,N_8641);
nor U15324 (N_15324,N_10567,N_10056);
xnor U15325 (N_15325,N_11634,N_10300);
nor U15326 (N_15326,N_9008,N_8043);
and U15327 (N_15327,N_9639,N_9943);
or U15328 (N_15328,N_9199,N_11199);
nand U15329 (N_15329,N_11383,N_9682);
or U15330 (N_15330,N_11445,N_9286);
nand U15331 (N_15331,N_9714,N_11989);
nand U15332 (N_15332,N_9930,N_10783);
nand U15333 (N_15333,N_10747,N_8076);
and U15334 (N_15334,N_11028,N_9054);
and U15335 (N_15335,N_11564,N_11932);
or U15336 (N_15336,N_10216,N_9578);
and U15337 (N_15337,N_8184,N_11194);
and U15338 (N_15338,N_8358,N_8322);
nor U15339 (N_15339,N_9911,N_10980);
nand U15340 (N_15340,N_8583,N_8453);
nor U15341 (N_15341,N_11426,N_11392);
nor U15342 (N_15342,N_10995,N_9660);
or U15343 (N_15343,N_9701,N_8982);
and U15344 (N_15344,N_8574,N_8490);
and U15345 (N_15345,N_10129,N_11927);
nor U15346 (N_15346,N_10367,N_9191);
or U15347 (N_15347,N_9466,N_8297);
nor U15348 (N_15348,N_9060,N_9570);
xor U15349 (N_15349,N_11563,N_11632);
xnor U15350 (N_15350,N_10888,N_10117);
xor U15351 (N_15351,N_9168,N_8592);
and U15352 (N_15352,N_8852,N_8549);
nor U15353 (N_15353,N_10217,N_9355);
nor U15354 (N_15354,N_9015,N_9461);
nor U15355 (N_15355,N_11878,N_9993);
or U15356 (N_15356,N_10541,N_11800);
nor U15357 (N_15357,N_10353,N_10689);
nor U15358 (N_15358,N_10499,N_10613);
nor U15359 (N_15359,N_10954,N_11537);
nand U15360 (N_15360,N_8985,N_11364);
or U15361 (N_15361,N_10765,N_9314);
nor U15362 (N_15362,N_11231,N_11843);
nor U15363 (N_15363,N_9350,N_9974);
nor U15364 (N_15364,N_10384,N_10557);
nand U15365 (N_15365,N_11007,N_9111);
nor U15366 (N_15366,N_10018,N_10338);
xor U15367 (N_15367,N_9900,N_9133);
nor U15368 (N_15368,N_8261,N_8096);
nor U15369 (N_15369,N_10846,N_9698);
or U15370 (N_15370,N_9520,N_11032);
and U15371 (N_15371,N_9082,N_8394);
xnor U15372 (N_15372,N_8382,N_9024);
or U15373 (N_15373,N_10392,N_9793);
nand U15374 (N_15374,N_10586,N_9842);
nand U15375 (N_15375,N_10078,N_11246);
nand U15376 (N_15376,N_10423,N_9972);
nand U15377 (N_15377,N_10984,N_11761);
nor U15378 (N_15378,N_8912,N_8222);
nand U15379 (N_15379,N_8328,N_8059);
or U15380 (N_15380,N_10126,N_11043);
nor U15381 (N_15381,N_9696,N_11071);
nor U15382 (N_15382,N_8139,N_9032);
nand U15383 (N_15383,N_11881,N_8818);
nor U15384 (N_15384,N_9198,N_11684);
nor U15385 (N_15385,N_9508,N_11348);
and U15386 (N_15386,N_9258,N_10273);
or U15387 (N_15387,N_9129,N_11854);
nor U15388 (N_15388,N_11137,N_9558);
nor U15389 (N_15389,N_9545,N_9247);
xor U15390 (N_15390,N_9740,N_9524);
and U15391 (N_15391,N_9826,N_11698);
and U15392 (N_15392,N_11689,N_9057);
nor U15393 (N_15393,N_9016,N_8276);
nand U15394 (N_15394,N_9017,N_11901);
nor U15395 (N_15395,N_10072,N_11284);
or U15396 (N_15396,N_10321,N_11351);
nor U15397 (N_15397,N_8157,N_9072);
nand U15398 (N_15398,N_9452,N_9532);
nand U15399 (N_15399,N_11138,N_8016);
nor U15400 (N_15400,N_10700,N_8482);
and U15401 (N_15401,N_9433,N_10125);
and U15402 (N_15402,N_11838,N_10949);
and U15403 (N_15403,N_9781,N_11593);
and U15404 (N_15404,N_8771,N_8054);
nand U15405 (N_15405,N_10819,N_10323);
or U15406 (N_15406,N_9160,N_10616);
nand U15407 (N_15407,N_10582,N_9988);
nand U15408 (N_15408,N_10989,N_10151);
nor U15409 (N_15409,N_8113,N_8859);
nand U15410 (N_15410,N_8840,N_9903);
nor U15411 (N_15411,N_11423,N_11766);
or U15412 (N_15412,N_11759,N_10631);
nand U15413 (N_15413,N_10084,N_10180);
and U15414 (N_15414,N_11392,N_11644);
or U15415 (N_15415,N_8826,N_10147);
nand U15416 (N_15416,N_11674,N_9422);
xor U15417 (N_15417,N_8737,N_8692);
and U15418 (N_15418,N_8481,N_8966);
nand U15419 (N_15419,N_8342,N_11689);
or U15420 (N_15420,N_8006,N_8269);
nor U15421 (N_15421,N_10810,N_8874);
and U15422 (N_15422,N_9923,N_8812);
and U15423 (N_15423,N_10289,N_9850);
or U15424 (N_15424,N_8450,N_9967);
or U15425 (N_15425,N_8209,N_8387);
and U15426 (N_15426,N_8833,N_11571);
or U15427 (N_15427,N_9524,N_11479);
or U15428 (N_15428,N_11231,N_9975);
nand U15429 (N_15429,N_8403,N_8081);
or U15430 (N_15430,N_10894,N_11120);
or U15431 (N_15431,N_10560,N_9967);
nor U15432 (N_15432,N_8556,N_8443);
nand U15433 (N_15433,N_11625,N_11496);
xor U15434 (N_15434,N_11238,N_9356);
or U15435 (N_15435,N_9799,N_8594);
and U15436 (N_15436,N_10791,N_8705);
or U15437 (N_15437,N_11902,N_11483);
and U15438 (N_15438,N_8639,N_8437);
and U15439 (N_15439,N_10453,N_8125);
xnor U15440 (N_15440,N_8345,N_8177);
nand U15441 (N_15441,N_10657,N_10924);
or U15442 (N_15442,N_11535,N_9618);
nand U15443 (N_15443,N_8332,N_8362);
nor U15444 (N_15444,N_8526,N_9635);
or U15445 (N_15445,N_11053,N_11525);
nor U15446 (N_15446,N_10156,N_10821);
and U15447 (N_15447,N_9806,N_10022);
or U15448 (N_15448,N_8181,N_10127);
xor U15449 (N_15449,N_9425,N_9164);
and U15450 (N_15450,N_11080,N_10651);
xnor U15451 (N_15451,N_11179,N_8088);
or U15452 (N_15452,N_8293,N_8951);
and U15453 (N_15453,N_11209,N_8172);
nand U15454 (N_15454,N_10894,N_8188);
or U15455 (N_15455,N_9066,N_9727);
nand U15456 (N_15456,N_8246,N_11170);
or U15457 (N_15457,N_9453,N_9140);
or U15458 (N_15458,N_8245,N_10164);
and U15459 (N_15459,N_11133,N_10200);
xnor U15460 (N_15460,N_8518,N_8800);
nor U15461 (N_15461,N_10238,N_8828);
and U15462 (N_15462,N_10527,N_8906);
nand U15463 (N_15463,N_10283,N_9756);
nor U15464 (N_15464,N_8701,N_10441);
or U15465 (N_15465,N_8594,N_8971);
nor U15466 (N_15466,N_11867,N_8256);
nand U15467 (N_15467,N_10397,N_11240);
and U15468 (N_15468,N_10153,N_10452);
or U15469 (N_15469,N_11213,N_9857);
nor U15470 (N_15470,N_8302,N_10454);
and U15471 (N_15471,N_8036,N_9085);
nor U15472 (N_15472,N_9783,N_8358);
nand U15473 (N_15473,N_8689,N_11183);
nand U15474 (N_15474,N_10622,N_8460);
or U15475 (N_15475,N_11241,N_9331);
nand U15476 (N_15476,N_10387,N_10453);
and U15477 (N_15477,N_9983,N_8439);
and U15478 (N_15478,N_9810,N_8083);
or U15479 (N_15479,N_8973,N_10482);
nand U15480 (N_15480,N_9950,N_8012);
or U15481 (N_15481,N_11709,N_9863);
and U15482 (N_15482,N_11182,N_9617);
and U15483 (N_15483,N_9238,N_11970);
nor U15484 (N_15484,N_8975,N_10104);
and U15485 (N_15485,N_9476,N_10430);
nor U15486 (N_15486,N_11003,N_10031);
nand U15487 (N_15487,N_9507,N_8083);
nor U15488 (N_15488,N_8791,N_10541);
nor U15489 (N_15489,N_8760,N_10899);
or U15490 (N_15490,N_10168,N_11332);
nand U15491 (N_15491,N_9278,N_10332);
nor U15492 (N_15492,N_11256,N_8031);
nand U15493 (N_15493,N_9587,N_9338);
or U15494 (N_15494,N_8483,N_10618);
nor U15495 (N_15495,N_11180,N_9501);
nor U15496 (N_15496,N_10964,N_9428);
or U15497 (N_15497,N_8143,N_8809);
or U15498 (N_15498,N_8145,N_10560);
nor U15499 (N_15499,N_11903,N_11735);
and U15500 (N_15500,N_8521,N_8703);
nor U15501 (N_15501,N_10912,N_10063);
xor U15502 (N_15502,N_9212,N_9487);
xor U15503 (N_15503,N_8908,N_9100);
xnor U15504 (N_15504,N_9319,N_9509);
xnor U15505 (N_15505,N_10471,N_9154);
or U15506 (N_15506,N_11416,N_8334);
nor U15507 (N_15507,N_9367,N_8230);
or U15508 (N_15508,N_10915,N_11698);
nand U15509 (N_15509,N_8246,N_9854);
and U15510 (N_15510,N_11070,N_9276);
nand U15511 (N_15511,N_8310,N_9320);
nor U15512 (N_15512,N_9969,N_9625);
nand U15513 (N_15513,N_10200,N_8808);
or U15514 (N_15514,N_9151,N_8693);
nor U15515 (N_15515,N_10800,N_10154);
or U15516 (N_15516,N_10894,N_8868);
nand U15517 (N_15517,N_10796,N_9585);
and U15518 (N_15518,N_8364,N_10760);
and U15519 (N_15519,N_9379,N_9745);
xor U15520 (N_15520,N_8956,N_9587);
or U15521 (N_15521,N_10649,N_8459);
nand U15522 (N_15522,N_8067,N_9389);
and U15523 (N_15523,N_11379,N_9852);
and U15524 (N_15524,N_9781,N_11933);
nand U15525 (N_15525,N_9950,N_8871);
and U15526 (N_15526,N_10776,N_11932);
nand U15527 (N_15527,N_8666,N_8504);
nand U15528 (N_15528,N_11376,N_11172);
or U15529 (N_15529,N_9544,N_9356);
nor U15530 (N_15530,N_11516,N_11242);
and U15531 (N_15531,N_9134,N_8234);
nand U15532 (N_15532,N_8565,N_10985);
xnor U15533 (N_15533,N_10730,N_8628);
and U15534 (N_15534,N_11740,N_9525);
or U15535 (N_15535,N_9693,N_9381);
and U15536 (N_15536,N_8770,N_10064);
or U15537 (N_15537,N_8388,N_11832);
and U15538 (N_15538,N_9457,N_9257);
nor U15539 (N_15539,N_8272,N_10908);
and U15540 (N_15540,N_8378,N_10935);
and U15541 (N_15541,N_11003,N_10967);
nand U15542 (N_15542,N_8120,N_8184);
nor U15543 (N_15543,N_8067,N_10992);
nand U15544 (N_15544,N_10352,N_9293);
or U15545 (N_15545,N_9721,N_11985);
nor U15546 (N_15546,N_11452,N_8115);
and U15547 (N_15547,N_8448,N_11636);
and U15548 (N_15548,N_8164,N_9049);
nand U15549 (N_15549,N_9766,N_11465);
nand U15550 (N_15550,N_11778,N_10640);
xor U15551 (N_15551,N_10848,N_9718);
nor U15552 (N_15552,N_11571,N_8949);
nand U15553 (N_15553,N_9910,N_9560);
and U15554 (N_15554,N_8522,N_9012);
or U15555 (N_15555,N_9115,N_10260);
nor U15556 (N_15556,N_10581,N_11123);
nor U15557 (N_15557,N_9510,N_11328);
and U15558 (N_15558,N_11768,N_11808);
and U15559 (N_15559,N_11919,N_8632);
nand U15560 (N_15560,N_9129,N_10369);
or U15561 (N_15561,N_9938,N_11556);
nand U15562 (N_15562,N_10776,N_10380);
nor U15563 (N_15563,N_10491,N_10933);
xor U15564 (N_15564,N_10633,N_11276);
xor U15565 (N_15565,N_9251,N_9186);
and U15566 (N_15566,N_10226,N_10063);
nand U15567 (N_15567,N_9215,N_8123);
or U15568 (N_15568,N_9110,N_11239);
nand U15569 (N_15569,N_8392,N_9456);
nand U15570 (N_15570,N_11466,N_10774);
xnor U15571 (N_15571,N_9951,N_8819);
nor U15572 (N_15572,N_11480,N_10423);
or U15573 (N_15573,N_11469,N_10081);
and U15574 (N_15574,N_10135,N_11701);
or U15575 (N_15575,N_10055,N_9174);
nor U15576 (N_15576,N_8056,N_10381);
and U15577 (N_15577,N_8146,N_9062);
nor U15578 (N_15578,N_9278,N_8128);
nor U15579 (N_15579,N_9020,N_11506);
nand U15580 (N_15580,N_8206,N_10303);
and U15581 (N_15581,N_8996,N_11645);
and U15582 (N_15582,N_8717,N_8028);
xnor U15583 (N_15583,N_10087,N_8336);
or U15584 (N_15584,N_10464,N_8219);
or U15585 (N_15585,N_11496,N_11914);
nor U15586 (N_15586,N_8998,N_8876);
and U15587 (N_15587,N_8436,N_9368);
xor U15588 (N_15588,N_9297,N_10978);
nor U15589 (N_15589,N_8422,N_11784);
and U15590 (N_15590,N_8971,N_8473);
nor U15591 (N_15591,N_8884,N_9436);
or U15592 (N_15592,N_11270,N_10816);
xnor U15593 (N_15593,N_8792,N_10465);
nor U15594 (N_15594,N_11960,N_11414);
xor U15595 (N_15595,N_11648,N_9067);
nor U15596 (N_15596,N_8354,N_8468);
and U15597 (N_15597,N_10428,N_10443);
or U15598 (N_15598,N_11679,N_10289);
or U15599 (N_15599,N_8755,N_9356);
nor U15600 (N_15600,N_10897,N_10744);
or U15601 (N_15601,N_11747,N_9885);
and U15602 (N_15602,N_10658,N_11567);
nor U15603 (N_15603,N_8448,N_10172);
and U15604 (N_15604,N_9105,N_11680);
nand U15605 (N_15605,N_11101,N_8352);
and U15606 (N_15606,N_10226,N_8961);
nand U15607 (N_15607,N_9594,N_11722);
nand U15608 (N_15608,N_10505,N_8995);
nand U15609 (N_15609,N_10156,N_10779);
nand U15610 (N_15610,N_8708,N_10564);
and U15611 (N_15611,N_10609,N_11928);
nor U15612 (N_15612,N_9705,N_8348);
nand U15613 (N_15613,N_11387,N_8303);
nand U15614 (N_15614,N_10409,N_9315);
nand U15615 (N_15615,N_9425,N_10747);
nor U15616 (N_15616,N_11646,N_8103);
or U15617 (N_15617,N_9781,N_11735);
nor U15618 (N_15618,N_9183,N_10132);
nand U15619 (N_15619,N_10508,N_10416);
and U15620 (N_15620,N_11011,N_10914);
xnor U15621 (N_15621,N_8702,N_10124);
nor U15622 (N_15622,N_8169,N_9649);
xor U15623 (N_15623,N_11293,N_8748);
or U15624 (N_15624,N_9524,N_9319);
and U15625 (N_15625,N_8427,N_8688);
or U15626 (N_15626,N_11900,N_9907);
and U15627 (N_15627,N_9764,N_9332);
or U15628 (N_15628,N_10751,N_11395);
xor U15629 (N_15629,N_8260,N_9937);
nand U15630 (N_15630,N_8592,N_8079);
and U15631 (N_15631,N_10639,N_8022);
nand U15632 (N_15632,N_10463,N_8480);
nand U15633 (N_15633,N_8593,N_10912);
nand U15634 (N_15634,N_9958,N_8297);
nor U15635 (N_15635,N_8877,N_10355);
nand U15636 (N_15636,N_9251,N_11061);
and U15637 (N_15637,N_9966,N_8804);
and U15638 (N_15638,N_10694,N_11338);
or U15639 (N_15639,N_8131,N_9527);
nor U15640 (N_15640,N_10200,N_9665);
nand U15641 (N_15641,N_10309,N_8315);
nor U15642 (N_15642,N_10204,N_9762);
and U15643 (N_15643,N_10594,N_8577);
and U15644 (N_15644,N_11941,N_9952);
and U15645 (N_15645,N_11448,N_11520);
nor U15646 (N_15646,N_8687,N_9475);
and U15647 (N_15647,N_8012,N_8104);
nand U15648 (N_15648,N_10489,N_11337);
and U15649 (N_15649,N_10050,N_10095);
and U15650 (N_15650,N_9110,N_8134);
nand U15651 (N_15651,N_11152,N_11018);
nand U15652 (N_15652,N_10909,N_8726);
xor U15653 (N_15653,N_9431,N_11368);
or U15654 (N_15654,N_10402,N_8543);
and U15655 (N_15655,N_10583,N_10586);
or U15656 (N_15656,N_8322,N_10939);
nor U15657 (N_15657,N_11558,N_9852);
nand U15658 (N_15658,N_8660,N_11180);
nor U15659 (N_15659,N_11847,N_10698);
and U15660 (N_15660,N_10519,N_11579);
nor U15661 (N_15661,N_9054,N_10711);
or U15662 (N_15662,N_10854,N_9961);
or U15663 (N_15663,N_11988,N_8168);
and U15664 (N_15664,N_10971,N_9896);
nor U15665 (N_15665,N_8039,N_11768);
nand U15666 (N_15666,N_8669,N_8710);
xnor U15667 (N_15667,N_8598,N_8740);
and U15668 (N_15668,N_8684,N_8911);
nand U15669 (N_15669,N_10640,N_11864);
and U15670 (N_15670,N_8992,N_8215);
nor U15671 (N_15671,N_8158,N_11796);
and U15672 (N_15672,N_8820,N_11439);
xor U15673 (N_15673,N_11154,N_9007);
and U15674 (N_15674,N_8136,N_9791);
and U15675 (N_15675,N_11941,N_10174);
xor U15676 (N_15676,N_9638,N_11509);
and U15677 (N_15677,N_8132,N_8491);
or U15678 (N_15678,N_9687,N_10522);
nand U15679 (N_15679,N_9774,N_11489);
nand U15680 (N_15680,N_10976,N_8698);
nor U15681 (N_15681,N_9911,N_9786);
nor U15682 (N_15682,N_11754,N_11631);
nand U15683 (N_15683,N_11013,N_9380);
or U15684 (N_15684,N_9450,N_8187);
or U15685 (N_15685,N_11205,N_8533);
or U15686 (N_15686,N_8741,N_10546);
nand U15687 (N_15687,N_10658,N_9473);
nand U15688 (N_15688,N_8809,N_10232);
or U15689 (N_15689,N_10166,N_10519);
xor U15690 (N_15690,N_8161,N_9858);
nor U15691 (N_15691,N_11132,N_9964);
and U15692 (N_15692,N_8527,N_11428);
nor U15693 (N_15693,N_10614,N_11052);
or U15694 (N_15694,N_11589,N_11300);
or U15695 (N_15695,N_11941,N_9671);
or U15696 (N_15696,N_11856,N_11644);
nor U15697 (N_15697,N_9697,N_11825);
xnor U15698 (N_15698,N_9403,N_10219);
nand U15699 (N_15699,N_8171,N_10863);
or U15700 (N_15700,N_11591,N_9639);
nand U15701 (N_15701,N_8876,N_11546);
xnor U15702 (N_15702,N_9253,N_9551);
nand U15703 (N_15703,N_10868,N_8746);
nor U15704 (N_15704,N_9477,N_10427);
or U15705 (N_15705,N_11516,N_11477);
nand U15706 (N_15706,N_9581,N_11042);
and U15707 (N_15707,N_9634,N_11422);
or U15708 (N_15708,N_8444,N_8738);
nand U15709 (N_15709,N_9947,N_8938);
and U15710 (N_15710,N_8548,N_8000);
nor U15711 (N_15711,N_11105,N_9059);
and U15712 (N_15712,N_11913,N_9175);
and U15713 (N_15713,N_9329,N_8769);
and U15714 (N_15714,N_8842,N_11180);
nand U15715 (N_15715,N_9331,N_11392);
nor U15716 (N_15716,N_10342,N_10762);
xnor U15717 (N_15717,N_11712,N_11297);
or U15718 (N_15718,N_8982,N_10025);
nor U15719 (N_15719,N_8071,N_11199);
nor U15720 (N_15720,N_11886,N_11275);
and U15721 (N_15721,N_10097,N_9238);
and U15722 (N_15722,N_11964,N_10460);
nor U15723 (N_15723,N_10391,N_11949);
nor U15724 (N_15724,N_9452,N_11734);
nand U15725 (N_15725,N_8810,N_10515);
or U15726 (N_15726,N_11258,N_8835);
or U15727 (N_15727,N_9696,N_8195);
or U15728 (N_15728,N_8450,N_8756);
or U15729 (N_15729,N_8770,N_11929);
or U15730 (N_15730,N_9458,N_8152);
and U15731 (N_15731,N_8504,N_9847);
and U15732 (N_15732,N_11918,N_11068);
and U15733 (N_15733,N_10022,N_11107);
nand U15734 (N_15734,N_8306,N_11725);
nor U15735 (N_15735,N_8894,N_9633);
nor U15736 (N_15736,N_10800,N_11883);
or U15737 (N_15737,N_9172,N_11896);
or U15738 (N_15738,N_9363,N_11295);
nor U15739 (N_15739,N_8145,N_11158);
nand U15740 (N_15740,N_10066,N_10007);
and U15741 (N_15741,N_9793,N_10444);
and U15742 (N_15742,N_8901,N_11104);
xor U15743 (N_15743,N_10777,N_11129);
and U15744 (N_15744,N_10166,N_11566);
xor U15745 (N_15745,N_10027,N_9876);
and U15746 (N_15746,N_8124,N_9031);
or U15747 (N_15747,N_9871,N_11843);
nand U15748 (N_15748,N_11392,N_11871);
xnor U15749 (N_15749,N_10557,N_8073);
and U15750 (N_15750,N_10662,N_11472);
and U15751 (N_15751,N_11092,N_9312);
nand U15752 (N_15752,N_10792,N_10278);
or U15753 (N_15753,N_10856,N_8225);
nand U15754 (N_15754,N_8055,N_9600);
nor U15755 (N_15755,N_9516,N_10882);
and U15756 (N_15756,N_11366,N_8018);
nand U15757 (N_15757,N_9568,N_11779);
or U15758 (N_15758,N_11541,N_9711);
or U15759 (N_15759,N_10115,N_11599);
nor U15760 (N_15760,N_9859,N_9730);
nor U15761 (N_15761,N_11628,N_8875);
nand U15762 (N_15762,N_11459,N_9036);
nor U15763 (N_15763,N_10517,N_8744);
and U15764 (N_15764,N_8834,N_10012);
and U15765 (N_15765,N_11738,N_8417);
nand U15766 (N_15766,N_11149,N_10330);
or U15767 (N_15767,N_10176,N_9269);
nor U15768 (N_15768,N_10603,N_11066);
xor U15769 (N_15769,N_8628,N_9567);
xnor U15770 (N_15770,N_10407,N_9295);
and U15771 (N_15771,N_8559,N_10022);
nand U15772 (N_15772,N_8026,N_11590);
or U15773 (N_15773,N_9573,N_11975);
nand U15774 (N_15774,N_8915,N_9327);
nand U15775 (N_15775,N_9503,N_11310);
or U15776 (N_15776,N_9836,N_8982);
or U15777 (N_15777,N_9519,N_10683);
or U15778 (N_15778,N_10412,N_11117);
or U15779 (N_15779,N_9037,N_9927);
or U15780 (N_15780,N_11017,N_10836);
or U15781 (N_15781,N_10088,N_9959);
nand U15782 (N_15782,N_10850,N_11568);
nor U15783 (N_15783,N_8472,N_11857);
xor U15784 (N_15784,N_11062,N_11223);
nor U15785 (N_15785,N_11374,N_9356);
nand U15786 (N_15786,N_11564,N_8518);
xnor U15787 (N_15787,N_11568,N_10256);
nand U15788 (N_15788,N_8958,N_11029);
and U15789 (N_15789,N_11831,N_9023);
nand U15790 (N_15790,N_8876,N_8507);
xnor U15791 (N_15791,N_8719,N_10704);
nand U15792 (N_15792,N_9848,N_8325);
or U15793 (N_15793,N_11394,N_8282);
nor U15794 (N_15794,N_8086,N_8522);
nand U15795 (N_15795,N_10594,N_10079);
nand U15796 (N_15796,N_11734,N_9189);
or U15797 (N_15797,N_9460,N_10740);
nor U15798 (N_15798,N_9750,N_10172);
nor U15799 (N_15799,N_10141,N_8978);
and U15800 (N_15800,N_10467,N_11597);
nor U15801 (N_15801,N_11440,N_11239);
and U15802 (N_15802,N_8596,N_9668);
and U15803 (N_15803,N_9403,N_11280);
and U15804 (N_15804,N_10816,N_10376);
xnor U15805 (N_15805,N_11406,N_9065);
nor U15806 (N_15806,N_10459,N_11755);
and U15807 (N_15807,N_10864,N_10668);
xor U15808 (N_15808,N_8858,N_11343);
and U15809 (N_15809,N_10329,N_9769);
nand U15810 (N_15810,N_9934,N_8771);
or U15811 (N_15811,N_11662,N_9595);
and U15812 (N_15812,N_11357,N_9864);
nor U15813 (N_15813,N_11731,N_10836);
nor U15814 (N_15814,N_11495,N_8287);
or U15815 (N_15815,N_10507,N_9023);
and U15816 (N_15816,N_10885,N_8833);
nor U15817 (N_15817,N_8562,N_10343);
nand U15818 (N_15818,N_11917,N_10600);
nand U15819 (N_15819,N_11423,N_8469);
nand U15820 (N_15820,N_9390,N_10267);
nand U15821 (N_15821,N_10069,N_8549);
or U15822 (N_15822,N_9591,N_10083);
or U15823 (N_15823,N_8725,N_10159);
nand U15824 (N_15824,N_10732,N_10436);
nand U15825 (N_15825,N_10618,N_11832);
and U15826 (N_15826,N_9794,N_10594);
or U15827 (N_15827,N_8932,N_11124);
xor U15828 (N_15828,N_11247,N_9909);
nand U15829 (N_15829,N_8233,N_11545);
and U15830 (N_15830,N_9385,N_9894);
nand U15831 (N_15831,N_10647,N_9161);
xor U15832 (N_15832,N_9688,N_11092);
and U15833 (N_15833,N_11753,N_9015);
nand U15834 (N_15834,N_11654,N_8503);
and U15835 (N_15835,N_9880,N_9376);
and U15836 (N_15836,N_9028,N_8348);
or U15837 (N_15837,N_8399,N_11214);
nand U15838 (N_15838,N_8256,N_11833);
nor U15839 (N_15839,N_9990,N_10385);
nand U15840 (N_15840,N_8796,N_11455);
nor U15841 (N_15841,N_8391,N_11352);
nor U15842 (N_15842,N_8653,N_11050);
or U15843 (N_15843,N_9987,N_10374);
and U15844 (N_15844,N_9821,N_8276);
nor U15845 (N_15845,N_11258,N_11565);
and U15846 (N_15846,N_8816,N_11385);
and U15847 (N_15847,N_8375,N_9185);
and U15848 (N_15848,N_8062,N_9297);
and U15849 (N_15849,N_8874,N_10924);
or U15850 (N_15850,N_10447,N_11155);
and U15851 (N_15851,N_11699,N_10100);
nor U15852 (N_15852,N_11335,N_8771);
xor U15853 (N_15853,N_11259,N_11820);
xnor U15854 (N_15854,N_9874,N_8665);
nor U15855 (N_15855,N_8798,N_11558);
nor U15856 (N_15856,N_9936,N_11715);
nand U15857 (N_15857,N_10644,N_9414);
nor U15858 (N_15858,N_9393,N_8008);
and U15859 (N_15859,N_8152,N_10866);
or U15860 (N_15860,N_10712,N_8757);
nand U15861 (N_15861,N_11878,N_8950);
and U15862 (N_15862,N_9449,N_9887);
or U15863 (N_15863,N_11911,N_11594);
nand U15864 (N_15864,N_8858,N_11667);
nor U15865 (N_15865,N_10756,N_8607);
xnor U15866 (N_15866,N_11313,N_10441);
nor U15867 (N_15867,N_11954,N_9078);
and U15868 (N_15868,N_9193,N_10646);
nor U15869 (N_15869,N_10487,N_11765);
nor U15870 (N_15870,N_10758,N_10644);
nand U15871 (N_15871,N_10764,N_11783);
nor U15872 (N_15872,N_11142,N_10017);
xnor U15873 (N_15873,N_8249,N_11472);
or U15874 (N_15874,N_10821,N_11716);
nor U15875 (N_15875,N_9581,N_11905);
or U15876 (N_15876,N_10030,N_8864);
nand U15877 (N_15877,N_10231,N_11173);
and U15878 (N_15878,N_10009,N_8857);
or U15879 (N_15879,N_8041,N_8510);
and U15880 (N_15880,N_8694,N_9723);
xnor U15881 (N_15881,N_8422,N_10557);
nand U15882 (N_15882,N_10047,N_8324);
and U15883 (N_15883,N_9324,N_8694);
xor U15884 (N_15884,N_9477,N_8146);
nand U15885 (N_15885,N_10472,N_9869);
nand U15886 (N_15886,N_11629,N_10583);
or U15887 (N_15887,N_8022,N_11444);
and U15888 (N_15888,N_9713,N_10488);
or U15889 (N_15889,N_9766,N_9525);
nor U15890 (N_15890,N_8193,N_11969);
or U15891 (N_15891,N_8305,N_8240);
and U15892 (N_15892,N_8911,N_9507);
and U15893 (N_15893,N_8818,N_9486);
xnor U15894 (N_15894,N_9022,N_11359);
or U15895 (N_15895,N_8670,N_11594);
nand U15896 (N_15896,N_8349,N_8989);
and U15897 (N_15897,N_11044,N_9446);
nor U15898 (N_15898,N_10045,N_11381);
or U15899 (N_15899,N_8638,N_10481);
nand U15900 (N_15900,N_9000,N_11815);
xnor U15901 (N_15901,N_8841,N_8312);
nand U15902 (N_15902,N_8171,N_11917);
xnor U15903 (N_15903,N_10695,N_9611);
nor U15904 (N_15904,N_10911,N_11236);
nand U15905 (N_15905,N_10834,N_9370);
nor U15906 (N_15906,N_9875,N_10890);
or U15907 (N_15907,N_9552,N_11270);
xnor U15908 (N_15908,N_11500,N_9723);
or U15909 (N_15909,N_8870,N_11586);
nand U15910 (N_15910,N_11303,N_11858);
nor U15911 (N_15911,N_8098,N_10696);
or U15912 (N_15912,N_9816,N_8814);
nor U15913 (N_15913,N_10286,N_10530);
nand U15914 (N_15914,N_9913,N_8869);
nand U15915 (N_15915,N_11010,N_9844);
nor U15916 (N_15916,N_8860,N_8017);
nor U15917 (N_15917,N_10785,N_10142);
xor U15918 (N_15918,N_8884,N_9993);
or U15919 (N_15919,N_10019,N_11630);
nand U15920 (N_15920,N_11446,N_11610);
and U15921 (N_15921,N_9698,N_11822);
nor U15922 (N_15922,N_11884,N_11365);
nand U15923 (N_15923,N_10135,N_8635);
and U15924 (N_15924,N_10525,N_11229);
xor U15925 (N_15925,N_10656,N_10500);
nand U15926 (N_15926,N_11008,N_11346);
nor U15927 (N_15927,N_10806,N_9587);
nor U15928 (N_15928,N_8640,N_9173);
or U15929 (N_15929,N_10342,N_9187);
and U15930 (N_15930,N_8850,N_8407);
and U15931 (N_15931,N_11018,N_11673);
and U15932 (N_15932,N_9869,N_8930);
or U15933 (N_15933,N_11952,N_10210);
and U15934 (N_15934,N_10311,N_8224);
and U15935 (N_15935,N_8618,N_8534);
xnor U15936 (N_15936,N_9601,N_9708);
nand U15937 (N_15937,N_9414,N_9885);
nor U15938 (N_15938,N_9713,N_9409);
nor U15939 (N_15939,N_9646,N_9733);
or U15940 (N_15940,N_9850,N_10394);
nor U15941 (N_15941,N_9824,N_9042);
nor U15942 (N_15942,N_8480,N_9864);
and U15943 (N_15943,N_10975,N_9600);
and U15944 (N_15944,N_9577,N_10850);
or U15945 (N_15945,N_8347,N_8848);
and U15946 (N_15946,N_9092,N_11307);
and U15947 (N_15947,N_8735,N_10422);
nand U15948 (N_15948,N_9027,N_8890);
and U15949 (N_15949,N_9403,N_9382);
nand U15950 (N_15950,N_10474,N_11582);
nand U15951 (N_15951,N_9382,N_9444);
and U15952 (N_15952,N_8541,N_11372);
and U15953 (N_15953,N_11798,N_8432);
and U15954 (N_15954,N_11489,N_8636);
or U15955 (N_15955,N_8982,N_8639);
and U15956 (N_15956,N_9145,N_9063);
nor U15957 (N_15957,N_11346,N_9270);
xnor U15958 (N_15958,N_9257,N_9022);
or U15959 (N_15959,N_8193,N_10704);
and U15960 (N_15960,N_11272,N_10684);
xor U15961 (N_15961,N_9825,N_8322);
and U15962 (N_15962,N_8682,N_9542);
nor U15963 (N_15963,N_10276,N_11504);
nor U15964 (N_15964,N_9066,N_8803);
and U15965 (N_15965,N_8361,N_10730);
or U15966 (N_15966,N_8494,N_11320);
nand U15967 (N_15967,N_10211,N_9368);
or U15968 (N_15968,N_9857,N_8883);
xnor U15969 (N_15969,N_9585,N_10217);
and U15970 (N_15970,N_9294,N_9559);
nor U15971 (N_15971,N_9609,N_10450);
or U15972 (N_15972,N_8371,N_10503);
nand U15973 (N_15973,N_11232,N_10170);
or U15974 (N_15974,N_10863,N_8181);
nor U15975 (N_15975,N_8602,N_9413);
or U15976 (N_15976,N_11330,N_11033);
nand U15977 (N_15977,N_8438,N_9493);
nand U15978 (N_15978,N_9889,N_9211);
nand U15979 (N_15979,N_11028,N_10382);
nor U15980 (N_15980,N_11121,N_10831);
nand U15981 (N_15981,N_9870,N_11668);
nor U15982 (N_15982,N_10152,N_10621);
xnor U15983 (N_15983,N_8550,N_10468);
and U15984 (N_15984,N_8493,N_11333);
xor U15985 (N_15985,N_8506,N_10009);
nor U15986 (N_15986,N_8195,N_8627);
nor U15987 (N_15987,N_10085,N_8356);
nor U15988 (N_15988,N_9402,N_11606);
or U15989 (N_15989,N_10749,N_10659);
and U15990 (N_15990,N_11836,N_11886);
and U15991 (N_15991,N_9972,N_9786);
nor U15992 (N_15992,N_9295,N_9354);
nor U15993 (N_15993,N_9396,N_11796);
xor U15994 (N_15994,N_8265,N_9868);
and U15995 (N_15995,N_8531,N_9153);
and U15996 (N_15996,N_11259,N_10003);
or U15997 (N_15997,N_8081,N_11399);
nand U15998 (N_15998,N_8507,N_9294);
nor U15999 (N_15999,N_11825,N_10316);
and U16000 (N_16000,N_15827,N_12627);
or U16001 (N_16001,N_12776,N_13830);
xor U16002 (N_16002,N_12743,N_14820);
and U16003 (N_16003,N_15120,N_12405);
and U16004 (N_16004,N_14228,N_12634);
and U16005 (N_16005,N_14427,N_12865);
nor U16006 (N_16006,N_12086,N_13143);
and U16007 (N_16007,N_15984,N_13123);
nand U16008 (N_16008,N_13663,N_13646);
nand U16009 (N_16009,N_13145,N_13415);
or U16010 (N_16010,N_13723,N_15973);
or U16011 (N_16011,N_14026,N_15908);
and U16012 (N_16012,N_15452,N_12957);
and U16013 (N_16013,N_15166,N_13768);
nand U16014 (N_16014,N_12510,N_13613);
and U16015 (N_16015,N_14307,N_14382);
and U16016 (N_16016,N_12829,N_15619);
or U16017 (N_16017,N_12479,N_14889);
nor U16018 (N_16018,N_14533,N_12664);
and U16019 (N_16019,N_15212,N_14224);
xor U16020 (N_16020,N_15253,N_12099);
xnor U16021 (N_16021,N_15260,N_15726);
nor U16022 (N_16022,N_15170,N_15457);
nor U16023 (N_16023,N_12144,N_15962);
nand U16024 (N_16024,N_15405,N_13810);
or U16025 (N_16025,N_14740,N_15736);
and U16026 (N_16026,N_14407,N_14952);
nor U16027 (N_16027,N_14730,N_15073);
nand U16028 (N_16028,N_15278,N_14115);
nand U16029 (N_16029,N_13995,N_14032);
nand U16030 (N_16030,N_13465,N_14636);
nor U16031 (N_16031,N_12445,N_14966);
nor U16032 (N_16032,N_12301,N_12791);
and U16033 (N_16033,N_13999,N_13552);
nand U16034 (N_16034,N_14790,N_13784);
xor U16035 (N_16035,N_13837,N_13140);
nand U16036 (N_16036,N_12140,N_14592);
and U16037 (N_16037,N_13960,N_13326);
or U16038 (N_16038,N_15413,N_14666);
nor U16039 (N_16039,N_13059,N_13407);
nand U16040 (N_16040,N_14805,N_15256);
nor U16041 (N_16041,N_13794,N_15410);
and U16042 (N_16042,N_15434,N_12695);
and U16043 (N_16043,N_14799,N_12775);
nor U16044 (N_16044,N_12989,N_15785);
nor U16045 (N_16045,N_13321,N_13472);
or U16046 (N_16046,N_13406,N_13139);
and U16047 (N_16047,N_12545,N_14641);
and U16048 (N_16048,N_15177,N_15066);
xnor U16049 (N_16049,N_12593,N_13453);
and U16050 (N_16050,N_14368,N_14974);
nor U16051 (N_16051,N_15014,N_15733);
or U16052 (N_16052,N_15495,N_12732);
xnor U16053 (N_16053,N_13260,N_15527);
nor U16054 (N_16054,N_14051,N_14833);
or U16055 (N_16055,N_12252,N_12498);
nor U16056 (N_16056,N_12841,N_12191);
nand U16057 (N_16057,N_14242,N_13316);
or U16058 (N_16058,N_14342,N_13628);
nand U16059 (N_16059,N_14275,N_15969);
xnor U16060 (N_16060,N_15860,N_15341);
nor U16061 (N_16061,N_15850,N_15661);
or U16062 (N_16062,N_15490,N_15044);
or U16063 (N_16063,N_13207,N_14306);
or U16064 (N_16064,N_13939,N_13184);
or U16065 (N_16065,N_15872,N_15467);
or U16066 (N_16066,N_13413,N_13197);
nand U16067 (N_16067,N_12685,N_13542);
nand U16068 (N_16068,N_15417,N_14718);
nor U16069 (N_16069,N_12423,N_13745);
xnor U16070 (N_16070,N_14043,N_15725);
or U16071 (N_16071,N_14300,N_13958);
nor U16072 (N_16072,N_13392,N_12183);
nor U16073 (N_16073,N_12861,N_15288);
nor U16074 (N_16074,N_15760,N_15659);
xnor U16075 (N_16075,N_15091,N_15141);
nor U16076 (N_16076,N_15747,N_15812);
nand U16077 (N_16077,N_12234,N_15754);
nor U16078 (N_16078,N_15772,N_12605);
nor U16079 (N_16079,N_13269,N_13511);
or U16080 (N_16080,N_14020,N_14894);
nor U16081 (N_16081,N_15562,N_15198);
nor U16082 (N_16082,N_14377,N_12657);
and U16083 (N_16083,N_14262,N_14201);
nor U16084 (N_16084,N_12859,N_14548);
nor U16085 (N_16085,N_14083,N_12670);
nor U16086 (N_16086,N_14831,N_13899);
nand U16087 (N_16087,N_14128,N_13494);
or U16088 (N_16088,N_15636,N_12203);
and U16089 (N_16089,N_13291,N_13838);
nand U16090 (N_16090,N_14074,N_14953);
or U16091 (N_16091,N_14492,N_12933);
and U16092 (N_16092,N_14880,N_13711);
nand U16093 (N_16093,N_14322,N_15142);
nand U16094 (N_16094,N_15420,N_14346);
and U16095 (N_16095,N_13584,N_15590);
or U16096 (N_16096,N_15670,N_15397);
or U16097 (N_16097,N_13560,N_15102);
nand U16098 (N_16098,N_12900,N_13875);
and U16099 (N_16099,N_14650,N_12230);
and U16100 (N_16100,N_13074,N_12754);
and U16101 (N_16101,N_12669,N_15823);
nor U16102 (N_16102,N_12796,N_13105);
nor U16103 (N_16103,N_15498,N_13485);
or U16104 (N_16104,N_15153,N_15067);
or U16105 (N_16105,N_14119,N_13893);
nor U16106 (N_16106,N_14168,N_15508);
or U16107 (N_16107,N_15666,N_12644);
or U16108 (N_16108,N_15920,N_13595);
nand U16109 (N_16109,N_12066,N_12939);
xor U16110 (N_16110,N_15199,N_12977);
nor U16111 (N_16111,N_12388,N_13342);
and U16112 (N_16112,N_12986,N_12390);
nand U16113 (N_16113,N_15591,N_14775);
or U16114 (N_16114,N_12538,N_14496);
or U16115 (N_16115,N_14612,N_14056);
and U16116 (N_16116,N_12629,N_14808);
or U16117 (N_16117,N_15978,N_15429);
nand U16118 (N_16118,N_12557,N_13573);
nor U16119 (N_16119,N_15228,N_12168);
or U16120 (N_16120,N_14215,N_13057);
or U16121 (N_16121,N_13660,N_13644);
or U16122 (N_16122,N_12642,N_15727);
or U16123 (N_16123,N_14369,N_15791);
nor U16124 (N_16124,N_14018,N_15547);
and U16125 (N_16125,N_13871,N_13412);
and U16126 (N_16126,N_13183,N_12693);
or U16127 (N_16127,N_15255,N_12408);
and U16128 (N_16128,N_15479,N_13509);
nor U16129 (N_16129,N_12744,N_14418);
nand U16130 (N_16130,N_14095,N_13028);
nor U16131 (N_16131,N_12990,N_14449);
nor U16132 (N_16132,N_12023,N_15686);
xor U16133 (N_16133,N_13164,N_15456);
nand U16134 (N_16134,N_14747,N_12561);
or U16135 (N_16135,N_15721,N_13303);
xor U16136 (N_16136,N_14383,N_15939);
or U16137 (N_16137,N_15882,N_13525);
xor U16138 (N_16138,N_13047,N_14338);
nand U16139 (N_16139,N_12962,N_13213);
or U16140 (N_16140,N_13701,N_14127);
and U16141 (N_16141,N_12482,N_14025);
nand U16142 (N_16142,N_15330,N_12332);
nand U16143 (N_16143,N_13440,N_12209);
and U16144 (N_16144,N_12480,N_13668);
nand U16145 (N_16145,N_12508,N_14815);
nand U16146 (N_16146,N_14595,N_13118);
or U16147 (N_16147,N_13828,N_13530);
nor U16148 (N_16148,N_12417,N_15319);
and U16149 (N_16149,N_15524,N_15543);
or U16150 (N_16150,N_14345,N_14375);
xnor U16151 (N_16151,N_12727,N_13795);
and U16152 (N_16152,N_13270,N_15271);
nor U16153 (N_16153,N_12152,N_12467);
xor U16154 (N_16154,N_14862,N_14395);
xnor U16155 (N_16155,N_15502,N_14325);
nand U16156 (N_16156,N_12300,N_12849);
nand U16157 (N_16157,N_14603,N_13892);
nor U16158 (N_16158,N_13228,N_14936);
and U16159 (N_16159,N_12293,N_12952);
xor U16160 (N_16160,N_12572,N_12641);
nand U16161 (N_16161,N_12495,N_14513);
or U16162 (N_16162,N_12832,N_13603);
and U16163 (N_16163,N_14009,N_12029);
or U16164 (N_16164,N_12391,N_15618);
and U16165 (N_16165,N_13776,N_13961);
nand U16166 (N_16166,N_15575,N_15099);
xnor U16167 (N_16167,N_12863,N_14841);
nor U16168 (N_16168,N_15767,N_12027);
nor U16169 (N_16169,N_13385,N_13643);
xor U16170 (N_16170,N_12367,N_12430);
xor U16171 (N_16171,N_12675,N_15796);
nand U16172 (N_16172,N_13704,N_13083);
or U16173 (N_16173,N_15399,N_13821);
xnor U16174 (N_16174,N_15633,N_12689);
and U16175 (N_16175,N_12236,N_13223);
or U16176 (N_16176,N_14002,N_13313);
or U16177 (N_16177,N_13879,N_14263);
nor U16178 (N_16178,N_15235,N_13447);
or U16179 (N_16179,N_15678,N_15477);
and U16180 (N_16180,N_15337,N_13499);
and U16181 (N_16181,N_15246,N_14870);
or U16182 (N_16182,N_14622,N_13675);
nor U16183 (N_16183,N_15862,N_15101);
and U16184 (N_16184,N_12412,N_14273);
or U16185 (N_16185,N_13426,N_13731);
or U16186 (N_16186,N_13421,N_14472);
nand U16187 (N_16187,N_12292,N_14837);
nand U16188 (N_16188,N_13559,N_14205);
nand U16189 (N_16189,N_14042,N_12741);
or U16190 (N_16190,N_14583,N_12456);
nor U16191 (N_16191,N_15665,N_14951);
and U16192 (N_16192,N_13881,N_15061);
nor U16193 (N_16193,N_12840,N_13479);
nor U16194 (N_16194,N_14264,N_14071);
nand U16195 (N_16195,N_14473,N_14426);
nand U16196 (N_16196,N_14839,N_13227);
xor U16197 (N_16197,N_13247,N_15040);
nand U16198 (N_16198,N_15994,N_15647);
or U16199 (N_16199,N_14725,N_15879);
and U16200 (N_16200,N_14296,N_14531);
and U16201 (N_16201,N_15864,N_14336);
nand U16202 (N_16202,N_13092,N_14102);
nor U16203 (N_16203,N_12531,N_12478);
xor U16204 (N_16204,N_14406,N_13214);
and U16205 (N_16205,N_13687,N_14447);
and U16206 (N_16206,N_12081,N_13898);
and U16207 (N_16207,N_12768,N_14064);
or U16208 (N_16208,N_15422,N_13642);
or U16209 (N_16209,N_15890,N_13135);
nand U16210 (N_16210,N_15194,N_14291);
nand U16211 (N_16211,N_13921,N_13980);
nand U16212 (N_16212,N_13306,N_13416);
and U16213 (N_16213,N_15913,N_12416);
and U16214 (N_16214,N_12373,N_12360);
and U16215 (N_16215,N_15111,N_15139);
xnor U16216 (N_16216,N_14590,N_15289);
or U16217 (N_16217,N_12368,N_14853);
nor U16218 (N_16218,N_13659,N_14192);
nand U16219 (N_16219,N_13751,N_13331);
nand U16220 (N_16220,N_13176,N_12746);
nand U16221 (N_16221,N_13201,N_12453);
or U16222 (N_16222,N_12909,N_13901);
nand U16223 (N_16223,N_15145,N_12337);
or U16224 (N_16224,N_12378,N_13318);
nor U16225 (N_16225,N_15026,N_14647);
nor U16226 (N_16226,N_12331,N_12087);
nor U16227 (N_16227,N_12343,N_15027);
nand U16228 (N_16228,N_14453,N_13437);
nand U16229 (N_16229,N_12160,N_14527);
nand U16230 (N_16230,N_13622,N_14804);
and U16231 (N_16231,N_14663,N_13855);
nand U16232 (N_16232,N_14742,N_14659);
and U16233 (N_16233,N_15828,N_13244);
nor U16234 (N_16234,N_13815,N_12499);
or U16235 (N_16235,N_12774,N_14667);
and U16236 (N_16236,N_15005,N_14525);
nor U16237 (N_16237,N_15564,N_13593);
nor U16238 (N_16238,N_14764,N_15906);
and U16239 (N_16239,N_14357,N_13051);
nor U16240 (N_16240,N_14037,N_15209);
nor U16241 (N_16241,N_15266,N_13189);
nand U16242 (N_16242,N_14225,N_12477);
xor U16243 (N_16243,N_15262,N_15176);
nor U16244 (N_16244,N_13035,N_15086);
or U16245 (N_16245,N_15902,N_14186);
and U16246 (N_16246,N_12162,N_12616);
and U16247 (N_16247,N_12275,N_13488);
and U16248 (N_16248,N_13112,N_15787);
or U16249 (N_16249,N_14339,N_14293);
nand U16250 (N_16250,N_13826,N_14122);
xnor U16251 (N_16251,N_14784,N_14567);
xor U16252 (N_16252,N_12836,N_15391);
nor U16253 (N_16253,N_14564,N_15105);
or U16254 (N_16254,N_12874,N_15757);
xnor U16255 (N_16255,N_12917,N_13279);
xor U16256 (N_16256,N_14237,N_15651);
xnor U16257 (N_16257,N_13082,N_15560);
or U16258 (N_16258,N_15691,N_12712);
nand U16259 (N_16259,N_15357,N_14487);
or U16260 (N_16260,N_13931,N_13376);
or U16261 (N_16261,N_15991,N_15358);
and U16262 (N_16262,N_15197,N_12635);
or U16263 (N_16263,N_14930,N_13919);
and U16264 (N_16264,N_13635,N_14643);
nand U16265 (N_16265,N_13816,N_13590);
nor U16266 (N_16266,N_15933,N_15745);
or U16267 (N_16267,N_14173,N_13229);
nand U16268 (N_16268,N_15532,N_12937);
or U16269 (N_16269,N_15512,N_14090);
or U16270 (N_16270,N_15234,N_12154);
or U16271 (N_16271,N_14781,N_13271);
or U16272 (N_16272,N_12138,N_15660);
or U16273 (N_16273,N_13597,N_12680);
and U16274 (N_16274,N_13913,N_15576);
and U16275 (N_16275,N_14142,N_15655);
or U16276 (N_16276,N_12097,N_14485);
and U16277 (N_16277,N_15259,N_12399);
xnor U16278 (N_16278,N_13363,N_13411);
nor U16279 (N_16279,N_15949,N_14290);
or U16280 (N_16280,N_13422,N_15640);
nor U16281 (N_16281,N_14459,N_15641);
xnor U16282 (N_16282,N_14304,N_12497);
nand U16283 (N_16283,N_13558,N_14464);
nand U16284 (N_16284,N_14579,N_13948);
and U16285 (N_16285,N_14668,N_15401);
or U16286 (N_16286,N_14305,N_14744);
nor U16287 (N_16287,N_12913,N_12061);
and U16288 (N_16288,N_12911,N_13505);
xor U16289 (N_16289,N_12830,N_13872);
and U16290 (N_16290,N_12339,N_15443);
or U16291 (N_16291,N_15738,N_15814);
and U16292 (N_16292,N_15281,N_14027);
xnor U16293 (N_16293,N_14356,N_15742);
nor U16294 (N_16294,N_14999,N_15542);
and U16295 (N_16295,N_13529,N_13918);
nand U16296 (N_16296,N_15961,N_15634);
xnor U16297 (N_16297,N_15096,N_15138);
and U16298 (N_16298,N_15342,N_13191);
or U16299 (N_16299,N_15517,N_14926);
xor U16300 (N_16300,N_14566,N_12556);
or U16301 (N_16301,N_12181,N_14467);
or U16302 (N_16302,N_12994,N_14905);
and U16303 (N_16303,N_15593,N_14259);
or U16304 (N_16304,N_14249,N_13832);
and U16305 (N_16305,N_12036,N_12812);
nand U16306 (N_16306,N_15200,N_14415);
or U16307 (N_16307,N_14363,N_14422);
nand U16308 (N_16308,N_15987,N_13110);
and U16309 (N_16309,N_15333,N_14469);
and U16310 (N_16310,N_13026,N_14500);
or U16311 (N_16311,N_14493,N_13365);
nand U16312 (N_16312,N_14807,N_15471);
or U16313 (N_16313,N_12244,N_14114);
nand U16314 (N_16314,N_15607,N_13592);
nand U16315 (N_16315,N_13434,N_13717);
nand U16316 (N_16316,N_12566,N_14945);
nor U16317 (N_16317,N_15140,N_13172);
or U16318 (N_16318,N_13766,N_12170);
or U16319 (N_16319,N_13755,N_14252);
and U16320 (N_16320,N_12505,N_15841);
or U16321 (N_16321,N_15613,N_12839);
nor U16322 (N_16322,N_13483,N_15930);
or U16323 (N_16323,N_12764,N_12038);
nor U16324 (N_16324,N_14780,N_12838);
or U16325 (N_16325,N_12098,N_14108);
and U16326 (N_16326,N_12030,N_12021);
nand U16327 (N_16327,N_12983,N_14298);
or U16328 (N_16328,N_14787,N_13924);
nor U16329 (N_16329,N_15798,N_12858);
and U16330 (N_16330,N_12193,N_12686);
nand U16331 (N_16331,N_14964,N_15071);
and U16332 (N_16332,N_13375,N_12080);
nand U16333 (N_16333,N_13027,N_13095);
and U16334 (N_16334,N_13917,N_15004);
nor U16335 (N_16335,N_13612,N_12147);
nor U16336 (N_16336,N_15440,N_12060);
nor U16337 (N_16337,N_14700,N_13393);
nor U16338 (N_16338,N_12327,N_13004);
or U16339 (N_16339,N_13161,N_15956);
and U16340 (N_16340,N_12222,N_14859);
or U16341 (N_16341,N_15497,N_14771);
nand U16342 (N_16342,N_14028,N_13192);
nand U16343 (N_16343,N_12235,N_12366);
nor U16344 (N_16344,N_12625,N_12772);
nand U16345 (N_16345,N_14125,N_13408);
and U16346 (N_16346,N_13536,N_15076);
nand U16347 (N_16347,N_14928,N_14637);
or U16348 (N_16348,N_15597,N_12512);
or U16349 (N_16349,N_14190,N_15941);
nor U16350 (N_16350,N_13144,N_12617);
nor U16351 (N_16351,N_15531,N_13076);
nand U16352 (N_16352,N_14661,N_12554);
or U16353 (N_16353,N_15699,N_13930);
nor U16354 (N_16354,N_12600,N_13521);
and U16355 (N_16355,N_15904,N_15696);
nand U16356 (N_16356,N_15032,N_13840);
nand U16357 (N_16357,N_13891,N_12521);
and U16358 (N_16358,N_12012,N_13429);
nand U16359 (N_16359,N_14266,N_15919);
or U16360 (N_16360,N_13741,N_14856);
or U16361 (N_16361,N_13812,N_12525);
or U16362 (N_16362,N_15290,N_14792);
nand U16363 (N_16363,N_13134,N_12398);
and U16364 (N_16364,N_12458,N_13932);
nor U16365 (N_16365,N_12185,N_13596);
nand U16366 (N_16366,N_13927,N_13014);
nor U16367 (N_16367,N_15998,N_15816);
nor U16368 (N_16368,N_14904,N_15297);
or U16369 (N_16369,N_12259,N_13341);
nor U16370 (N_16370,N_14310,N_15586);
and U16371 (N_16371,N_15608,N_12780);
nor U16372 (N_16372,N_15786,N_14331);
or U16373 (N_16373,N_15390,N_13371);
nor U16374 (N_16374,N_15205,N_13276);
and U16375 (N_16375,N_15276,N_13733);
nor U16376 (N_16376,N_12349,N_13506);
nor U16377 (N_16377,N_13888,N_15668);
and U16378 (N_16378,N_14677,N_15845);
xor U16379 (N_16379,N_14942,N_15104);
nor U16380 (N_16380,N_13272,N_12713);
nand U16381 (N_16381,N_15624,N_15267);
and U16382 (N_16382,N_15094,N_15866);
and U16383 (N_16383,N_15952,N_12017);
or U16384 (N_16384,N_15954,N_15081);
nor U16385 (N_16385,N_12363,N_12663);
nand U16386 (N_16386,N_13116,N_13650);
and U16387 (N_16387,N_12431,N_12033);
or U16388 (N_16388,N_15803,N_15018);
nor U16389 (N_16389,N_14269,N_13364);
and U16390 (N_16390,N_12661,N_14658);
nand U16391 (N_16391,N_15598,N_12553);
nand U16392 (N_16392,N_15716,N_13743);
nand U16393 (N_16393,N_15677,N_12681);
xnor U16394 (N_16394,N_12148,N_15982);
nor U16395 (N_16395,N_13078,N_12878);
xor U16396 (N_16396,N_13137,N_15368);
or U16397 (N_16397,N_15874,N_14549);
xnor U16398 (N_16398,N_12006,N_12919);
nor U16399 (N_16399,N_13010,N_14465);
and U16400 (N_16400,N_15213,N_14099);
or U16401 (N_16401,N_15243,N_15628);
and U16402 (N_16402,N_12647,N_14711);
or U16403 (N_16403,N_14302,N_14408);
nand U16404 (N_16404,N_15192,N_14483);
xnor U16405 (N_16405,N_13327,N_15327);
or U16406 (N_16406,N_15306,N_14717);
nand U16407 (N_16407,N_14550,N_13162);
nor U16408 (N_16408,N_14208,N_13423);
nor U16409 (N_16409,N_15447,N_12935);
nand U16410 (N_16410,N_13524,N_13772);
and U16411 (N_16411,N_12044,N_13289);
and U16412 (N_16412,N_14748,N_13261);
or U16413 (N_16413,N_13902,N_15367);
and U16414 (N_16414,N_13389,N_15692);
xor U16415 (N_16415,N_15189,N_14359);
nor U16416 (N_16416,N_12393,N_14005);
nand U16417 (N_16417,N_15848,N_15284);
and U16418 (N_16418,N_12402,N_15568);
and U16419 (N_16419,N_13791,N_13890);
nand U16420 (N_16420,N_14340,N_14210);
and U16421 (N_16421,N_15662,N_13975);
or U16422 (N_16422,N_13096,N_15445);
xnor U16423 (N_16423,N_14022,N_12317);
or U16424 (N_16424,N_14983,N_14349);
or U16425 (N_16425,N_12837,N_12206);
nand U16426 (N_16426,N_14970,N_13240);
or U16427 (N_16427,N_12090,N_15748);
nand U16428 (N_16428,N_15623,N_13574);
and U16429 (N_16429,N_15753,N_12464);
nor U16430 (N_16430,N_14137,N_14975);
nand U16431 (N_16431,N_15286,N_12314);
or U16432 (N_16432,N_14482,N_14000);
and U16433 (N_16433,N_13006,N_15298);
or U16434 (N_16434,N_13972,N_15698);
or U16435 (N_16435,N_14016,N_15448);
nor U16436 (N_16436,N_14844,N_14720);
or U16437 (N_16437,N_13950,N_13532);
and U16438 (N_16438,N_12740,N_15300);
nand U16439 (N_16439,N_13058,N_14414);
and U16440 (N_16440,N_12062,N_13388);
or U16441 (N_16441,N_12125,N_14167);
and U16442 (N_16442,N_12396,N_14706);
nor U16443 (N_16443,N_13575,N_15707);
nand U16444 (N_16444,N_12192,N_14536);
and U16445 (N_16445,N_15047,N_12873);
and U16446 (N_16446,N_15480,N_12719);
xor U16447 (N_16447,N_12823,N_12034);
and U16448 (N_16448,N_13209,N_12050);
or U16449 (N_16449,N_13955,N_15492);
and U16450 (N_16450,N_14917,N_13462);
and U16451 (N_16451,N_12221,N_15540);
nor U16452 (N_16452,N_12626,N_13049);
nor U16453 (N_16453,N_13109,N_15779);
and U16454 (N_16454,N_12658,N_12526);
and U16455 (N_16455,N_15997,N_15574);
nand U16456 (N_16456,N_12586,N_12386);
and U16457 (N_16457,N_15824,N_12834);
nor U16458 (N_16458,N_14958,N_13707);
nor U16459 (N_16459,N_15155,N_13545);
nand U16460 (N_16460,N_14052,N_13199);
and U16461 (N_16461,N_14374,N_14959);
nand U16462 (N_16462,N_12753,N_15468);
nor U16463 (N_16463,N_15844,N_15051);
nor U16464 (N_16464,N_13284,N_14347);
and U16465 (N_16465,N_15936,N_15349);
nor U16466 (N_16466,N_15674,N_14861);
nor U16467 (N_16467,N_15788,N_13749);
xor U16468 (N_16468,N_15122,N_14789);
and U16469 (N_16469,N_14625,N_15559);
or U16470 (N_16470,N_12371,N_15159);
xor U16471 (N_16471,N_13645,N_15755);
nor U16472 (N_16472,N_15895,N_13971);
xnor U16473 (N_16473,N_14685,N_14295);
nor U16474 (N_16474,N_13758,N_13329);
and U16475 (N_16475,N_13103,N_15307);
and U16476 (N_16476,N_12734,N_12345);
and U16477 (N_16477,N_14933,N_15264);
nand U16478 (N_16478,N_13068,N_15441);
nand U16479 (N_16479,N_15567,N_14814);
nand U16480 (N_16480,N_15513,N_12319);
and U16481 (N_16481,N_14088,N_14708);
and U16482 (N_16482,N_13583,N_13850);
nor U16483 (N_16483,N_15996,N_13322);
or U16484 (N_16484,N_15315,N_12220);
and U16485 (N_16485,N_13834,N_15589);
or U16486 (N_16486,N_12418,N_13661);
nor U16487 (N_16487,N_13259,N_12156);
or U16488 (N_16488,N_15020,N_15351);
or U16489 (N_16489,N_14559,N_14682);
and U16490 (N_16490,N_14222,N_15972);
nor U16491 (N_16491,N_12042,N_13173);
nand U16492 (N_16492,N_12093,N_13195);
nand U16493 (N_16493,N_15380,N_14479);
or U16494 (N_16494,N_14539,N_12843);
nand U16495 (N_16495,N_13349,N_14523);
nor U16496 (N_16496,N_14152,N_14394);
or U16497 (N_16497,N_13237,N_12427);
and U16498 (N_16498,N_15112,N_12524);
xor U16499 (N_16499,N_13773,N_13805);
nand U16500 (N_16500,N_14204,N_15818);
or U16501 (N_16501,N_14593,N_13267);
nor U16502 (N_16502,N_15424,N_13641);
nand U16503 (N_16503,N_14420,N_12736);
nor U16504 (N_16504,N_12999,N_14334);
and U16505 (N_16505,N_14553,N_13021);
nor U16506 (N_16506,N_13252,N_15732);
and U16507 (N_16507,N_14121,N_14562);
nand U16508 (N_16508,N_14628,N_12804);
nand U16509 (N_16509,N_12987,N_13730);
and U16510 (N_16510,N_15326,N_13507);
or U16511 (N_16511,N_12903,N_14697);
nand U16512 (N_16512,N_14207,N_12720);
nor U16513 (N_16513,N_12618,N_14961);
nor U16514 (N_16514,N_12981,N_12892);
nor U16515 (N_16515,N_12808,N_15435);
or U16516 (N_16516,N_12888,N_14801);
nor U16517 (N_16517,N_12132,N_13020);
xor U16518 (N_16518,N_14376,N_13860);
xor U16519 (N_16519,N_12920,N_14842);
nor U16520 (N_16520,N_14796,N_14312);
or U16521 (N_16521,N_12142,N_13557);
nor U16522 (N_16522,N_15187,N_13884);
nor U16523 (N_16523,N_13204,N_15510);
nand U16524 (N_16524,N_14149,N_15293);
and U16525 (N_16525,N_15250,N_14779);
or U16526 (N_16526,N_12494,N_15064);
xor U16527 (N_16527,N_13219,N_14316);
and U16528 (N_16528,N_12546,N_13679);
nor U16529 (N_16529,N_13620,N_14572);
or U16530 (N_16530,N_13174,N_15491);
nor U16531 (N_16531,N_13377,N_13211);
nor U16532 (N_16532,N_12704,N_13464);
nand U16533 (N_16533,N_12569,N_15815);
nand U16534 (N_16534,N_15313,N_15861);
and U16535 (N_16535,N_13196,N_12509);
nor U16536 (N_16536,N_12815,N_15609);
and U16537 (N_16537,N_14956,N_14529);
nand U16538 (N_16538,N_13383,N_14921);
nand U16539 (N_16539,N_12382,N_14630);
and U16540 (N_16540,N_12186,N_15374);
xor U16541 (N_16541,N_15310,N_14367);
xnor U16542 (N_16542,N_12974,N_12630);
nand U16543 (N_16543,N_12005,N_14797);
or U16544 (N_16544,N_13066,N_13782);
xnor U16545 (N_16545,N_15778,N_14895);
or U16546 (N_16546,N_13097,N_13009);
and U16547 (N_16547,N_12071,N_14508);
nor U16548 (N_16548,N_13065,N_14721);
or U16549 (N_16549,N_15868,N_15888);
nor U16550 (N_16550,N_13222,N_13340);
xnor U16551 (N_16551,N_14001,N_13430);
and U16552 (N_16552,N_12971,N_13001);
nand U16553 (N_16553,N_13293,N_14082);
nand U16554 (N_16554,N_13215,N_12507);
nand U16555 (N_16555,N_15588,N_14411);
nand U16556 (N_16556,N_13579,N_14869);
and U16557 (N_16557,N_14087,N_12930);
nor U16558 (N_16558,N_12846,N_13477);
and U16559 (N_16559,N_15127,N_14848);
nand U16560 (N_16560,N_12700,N_13869);
nand U16561 (N_16561,N_13452,N_12921);
and U16562 (N_16562,N_15834,N_12536);
and U16563 (N_16563,N_12073,N_15438);
nand U16564 (N_16564,N_15119,N_15007);
and U16565 (N_16565,N_14934,N_12130);
and U16566 (N_16566,N_13916,N_15777);
and U16567 (N_16567,N_15953,N_12204);
nor U16568 (N_16568,N_14410,N_13601);
nand U16569 (N_16569,N_15592,N_15928);
or U16570 (N_16570,N_14507,N_15070);
nand U16571 (N_16571,N_15820,N_12585);
or U16572 (N_16572,N_13651,N_13496);
xor U16573 (N_16573,N_15396,N_12486);
or U16574 (N_16574,N_13455,N_14845);
and U16575 (N_16575,N_13040,N_15911);
and U16576 (N_16576,N_13205,N_14218);
nor U16577 (N_16577,N_13716,N_13640);
nor U16578 (N_16578,N_12898,N_14750);
or U16579 (N_16579,N_15923,N_15799);
nor U16580 (N_16580,N_12790,N_15218);
nor U16581 (N_16581,N_12157,N_13807);
nor U16582 (N_16582,N_13978,N_13315);
or U16583 (N_16583,N_12710,N_14800);
or U16584 (N_16584,N_13578,N_12574);
nor U16585 (N_16585,N_13937,N_14832);
nor U16586 (N_16586,N_14745,N_12271);
nand U16587 (N_16587,N_15995,N_13604);
or U16588 (N_16588,N_13188,N_15751);
and U16589 (N_16589,N_12184,N_14280);
and U16590 (N_16590,N_12350,N_13077);
or U16591 (N_16591,N_12308,N_14574);
or U16592 (N_16592,N_14519,N_12628);
and U16593 (N_16593,N_13417,N_13347);
or U16594 (N_16594,N_12852,N_14286);
or U16595 (N_16595,N_13617,N_14971);
nor U16596 (N_16596,N_15340,N_13726);
and U16597 (N_16597,N_14955,N_14358);
and U16598 (N_16598,N_13526,N_15783);
nand U16599 (N_16599,N_14417,N_13992);
nor U16600 (N_16600,N_13450,N_12963);
and U16601 (N_16601,N_13556,N_12896);
nand U16602 (N_16602,N_15428,N_15049);
nand U16603 (N_16603,N_12523,N_15817);
xnor U16604 (N_16604,N_13940,N_13101);
xnor U16605 (N_16605,N_13637,N_12562);
xnor U16606 (N_16606,N_14413,N_15360);
nand U16607 (N_16607,N_13963,N_13959);
nor U16608 (N_16608,N_14752,N_12868);
or U16609 (N_16609,N_15299,N_12076);
nand U16610 (N_16610,N_13121,N_13263);
xnor U16611 (N_16611,N_12894,N_12650);
or U16612 (N_16612,N_13115,N_15355);
nor U16613 (N_16613,N_13522,N_13862);
or U16614 (N_16614,N_14757,N_15700);
and U16615 (N_16615,N_13718,N_15263);
nor U16616 (N_16616,N_14915,N_15606);
nor U16617 (N_16617,N_13216,N_14591);
and U16618 (N_16618,N_13833,N_12998);
or U16619 (N_16619,N_15173,N_13801);
nand U16620 (N_16620,N_12760,N_15673);
xor U16621 (N_16621,N_14033,N_13305);
xnor U16622 (N_16622,N_14435,N_15643);
nor U16623 (N_16623,N_12440,N_15937);
nor U16624 (N_16624,N_13348,N_12276);
xor U16625 (N_16625,N_12907,N_13569);
or U16626 (N_16626,N_15175,N_15129);
nor U16627 (N_16627,N_15762,N_14003);
and U16628 (N_16628,N_12065,N_12159);
nand U16629 (N_16629,N_14791,N_14758);
nand U16630 (N_16630,N_12232,N_15690);
xnor U16631 (N_16631,N_14440,N_14147);
nor U16632 (N_16632,N_12908,N_14132);
and U16633 (N_16633,N_14284,N_14055);
and U16634 (N_16634,N_15831,N_15764);
nand U16635 (N_16635,N_14399,N_12122);
nand U16636 (N_16636,N_15539,N_13132);
nor U16637 (N_16637,N_15537,N_13907);
nor U16638 (N_16638,N_13533,N_12844);
and U16639 (N_16639,N_14437,N_12651);
and U16640 (N_16640,N_15217,N_13947);
or U16641 (N_16641,N_15781,N_12737);
and U16642 (N_16642,N_15459,N_13359);
or U16643 (N_16643,N_12988,N_13674);
nor U16644 (N_16644,N_12241,N_15292);
nor U16645 (N_16645,N_14209,N_12289);
nor U16646 (N_16646,N_15769,N_12517);
or U16647 (N_16647,N_13548,N_12264);
or U16648 (N_16648,N_13056,N_15320);
or U16649 (N_16649,N_12053,N_14546);
nor U16650 (N_16650,N_15811,N_15885);
or U16651 (N_16651,N_12596,N_12528);
nor U16652 (N_16652,N_13742,N_13594);
and U16653 (N_16653,N_13131,N_14092);
nand U16654 (N_16654,N_14881,N_15638);
xnor U16655 (N_16655,N_13988,N_15265);
nand U16656 (N_16656,N_12288,N_13920);
nand U16657 (N_16657,N_14515,N_13451);
or U16658 (N_16658,N_15648,N_13649);
xnor U16659 (N_16659,N_12799,N_14066);
nand U16660 (N_16660,N_15680,N_14526);
and U16661 (N_16661,N_12118,N_13029);
or U16662 (N_16662,N_13541,N_15534);
xor U16663 (N_16663,N_12601,N_14978);
nor U16664 (N_16664,N_14013,N_14520);
and U16665 (N_16665,N_12749,N_14069);
nand U16666 (N_16666,N_13344,N_13476);
xnor U16667 (N_16667,N_12000,N_13190);
or U16668 (N_16668,N_14893,N_15083);
or U16669 (N_16669,N_15309,N_15756);
nor U16670 (N_16670,N_12707,N_14922);
xnor U16671 (N_16671,N_15909,N_12568);
xnor U16672 (N_16672,N_13676,N_13954);
and U16673 (N_16673,N_13069,N_13256);
or U16674 (N_16674,N_12520,N_15379);
nand U16675 (N_16675,N_13946,N_15172);
nand U16676 (N_16676,N_14672,N_12096);
nand U16677 (N_16677,N_15203,N_13953);
and U16678 (N_16678,N_12255,N_13433);
xnor U16679 (N_16679,N_12009,N_14456);
nor U16680 (N_16680,N_15054,N_15897);
and U16681 (N_16681,N_15347,N_14746);
xor U16682 (N_16682,N_14193,N_14557);
nor U16683 (N_16683,N_14932,N_12443);
or U16684 (N_16684,N_14409,N_14048);
nor U16685 (N_16685,N_14913,N_15917);
nand U16686 (N_16686,N_15202,N_12679);
and U16687 (N_16687,N_15179,N_14008);
nor U16688 (N_16688,N_12225,N_13126);
or U16689 (N_16689,N_12436,N_12800);
and U16690 (N_16690,N_12294,N_12672);
and U16691 (N_16691,N_14311,N_13949);
xnor U16692 (N_16692,N_15971,N_13255);
or U16693 (N_16693,N_14158,N_13692);
xnor U16694 (N_16694,N_13550,N_13079);
or U16695 (N_16695,N_14196,N_12759);
xor U16696 (N_16696,N_14163,N_12954);
or U16697 (N_16697,N_14714,N_15905);
and U16698 (N_16698,N_13665,N_14140);
or U16699 (N_16699,N_13230,N_13372);
xnor U16700 (N_16700,N_13241,N_13586);
nand U16701 (N_16701,N_14044,N_15947);
nand U16702 (N_16702,N_13866,N_14332);
nor U16703 (N_16703,N_14432,N_13817);
and U16704 (N_16704,N_14235,N_15211);
nand U16705 (N_16705,N_13979,N_14843);
or U16706 (N_16706,N_14530,N_14247);
and U16707 (N_16707,N_14772,N_13814);
xor U16708 (N_16708,N_15999,N_13588);
nor U16709 (N_16709,N_12716,N_12136);
and U16710 (N_16710,N_14704,N_12662);
or U16711 (N_16711,N_14034,N_15436);
or U16712 (N_16712,N_12581,N_12794);
and U16713 (N_16713,N_13467,N_13387);
and U16714 (N_16714,N_14433,N_14610);
and U16715 (N_16715,N_15439,N_13328);
or U16716 (N_16716,N_13369,N_14702);
nand U16717 (N_16717,N_14824,N_13740);
nand U16718 (N_16718,N_15344,N_14812);
and U16719 (N_16719,N_15561,N_15106);
or U16720 (N_16720,N_12706,N_13852);
nor U16721 (N_16721,N_12442,N_12872);
nand U16722 (N_16722,N_13038,N_13352);
and U16723 (N_16723,N_12660,N_12454);
and U16724 (N_16724,N_14642,N_15002);
or U16725 (N_16725,N_14555,N_15146);
and U16726 (N_16726,N_14818,N_15729);
or U16727 (N_16727,N_14317,N_12290);
and U16728 (N_16728,N_14371,N_13159);
nand U16729 (N_16729,N_15100,N_15273);
nor U16730 (N_16730,N_14233,N_12471);
and U16731 (N_16731,N_15715,N_13886);
and U16732 (N_16732,N_14486,N_12483);
nor U16733 (N_16733,N_12539,N_15871);
nor U16734 (N_16734,N_14608,N_12978);
and U16735 (N_16735,N_12195,N_15376);
xnor U16736 (N_16736,N_13474,N_15516);
nand U16737 (N_16737,N_12711,N_15653);
or U16738 (N_16738,N_12251,N_15829);
nand U16739 (N_16739,N_13091,N_13634);
or U16740 (N_16740,N_15622,N_13966);
and U16741 (N_16741,N_12697,N_12281);
nor U16742 (N_16742,N_12291,N_14067);
nor U16743 (N_16743,N_14098,N_15843);
nand U16744 (N_16744,N_13580,N_15835);
or U16745 (N_16745,N_12424,N_14060);
and U16746 (N_16746,N_15979,N_12637);
and U16747 (N_16747,N_13775,N_13928);
nor U16748 (N_16748,N_12778,N_12652);
or U16749 (N_16749,N_12484,N_14751);
nand U16750 (N_16750,N_15530,N_14144);
and U16751 (N_16751,N_14762,N_15556);
or U16752 (N_16752,N_12380,N_13370);
or U16753 (N_16753,N_14920,N_14944);
and U16754 (N_16754,N_12214,N_14785);
nand U16755 (N_16755,N_15421,N_12698);
nand U16756 (N_16756,N_14189,N_15414);
xnor U16757 (N_16757,N_12135,N_13878);
xnor U16758 (N_16758,N_12109,N_14480);
nand U16759 (N_16759,N_13242,N_12648);
or U16760 (N_16760,N_13626,N_12847);
nor U16761 (N_16761,N_13338,N_13576);
nand U16762 (N_16762,N_13425,N_14116);
or U16763 (N_16763,N_13623,N_12432);
nor U16764 (N_16764,N_13625,N_12102);
nand U16765 (N_16765,N_13905,N_14656);
nand U16766 (N_16766,N_12419,N_15077);
and U16767 (N_16767,N_15740,N_14911);
nand U16768 (N_16768,N_14887,N_15889);
xnor U16769 (N_16769,N_14646,N_15958);
nand U16770 (N_16770,N_12299,N_15001);
nand U16771 (N_16771,N_15110,N_12756);
or U16772 (N_16772,N_14191,N_12083);
xor U16773 (N_16773,N_14111,N_15565);
nor U16774 (N_16774,N_13378,N_14397);
or U16775 (N_16775,N_14716,N_15022);
nor U16776 (N_16776,N_14973,N_15719);
nor U16777 (N_16777,N_14231,N_13041);
nand U16778 (N_16778,N_15305,N_12855);
nand U16779 (N_16779,N_15734,N_15507);
nor U16780 (N_16780,N_14906,N_12826);
nor U16781 (N_16781,N_14653,N_15134);
and U16782 (N_16782,N_12735,N_15169);
or U16783 (N_16783,N_14888,N_12682);
xor U16784 (N_16784,N_14826,N_13249);
nor U16785 (N_16785,N_15730,N_13486);
nor U16786 (N_16786,N_12422,N_12819);
and U16787 (N_16787,N_12046,N_15950);
nand U16788 (N_16788,N_12752,N_13599);
nand U16789 (N_16789,N_14011,N_13317);
nor U16790 (N_16790,N_13350,N_15035);
nand U16791 (N_16791,N_15806,N_12223);
nand U16792 (N_16792,N_14691,N_14385);
nor U16793 (N_16793,N_14314,N_13165);
xor U16794 (N_16794,N_14260,N_14372);
or U16795 (N_16795,N_14118,N_15394);
nand U16796 (N_16796,N_14126,N_15989);
and U16797 (N_16797,N_14162,N_15015);
or U16798 (N_16798,N_14524,N_14100);
and U16799 (N_16799,N_14159,N_14161);
nor U16800 (N_16800,N_12260,N_14876);
nor U16801 (N_16801,N_13809,N_14997);
or U16802 (N_16802,N_15934,N_13771);
nand U16803 (N_16803,N_12365,N_15993);
xnor U16804 (N_16804,N_12429,N_14819);
and U16805 (N_16805,N_13563,N_13128);
and U16806 (N_16806,N_12024,N_14244);
or U16807 (N_16807,N_13210,N_13459);
nor U16808 (N_16808,N_12848,N_14091);
or U16809 (N_16809,N_15282,N_14400);
nor U16810 (N_16810,N_13678,N_12179);
and U16811 (N_16811,N_13098,N_13909);
nand U16812 (N_16812,N_13608,N_15722);
or U16813 (N_16813,N_13294,N_12853);
nand U16814 (N_16814,N_14875,N_14501);
or U16815 (N_16815,N_15682,N_12325);
and U16816 (N_16816,N_12375,N_14169);
or U16817 (N_16817,N_15450,N_15222);
nand U16818 (N_16818,N_14200,N_12226);
nor U16819 (N_16819,N_13774,N_12943);
nor U16820 (N_16820,N_13770,N_15365);
nand U16821 (N_16821,N_15251,N_15453);
nor U16822 (N_16822,N_15478,N_13484);
nor U16823 (N_16823,N_15158,N_14767);
nand U16824 (N_16824,N_12013,N_15663);
xnor U16825 (N_16825,N_13081,N_13591);
nor U16826 (N_16826,N_14139,N_14141);
xnor U16827 (N_16827,N_13292,N_13813);
or U16828 (N_16828,N_13245,N_13070);
and U16829 (N_16829,N_15345,N_15887);
nor U16830 (N_16830,N_12321,N_13444);
nand U16831 (N_16831,N_12668,N_14885);
and U16832 (N_16832,N_13234,N_15204);
nor U16833 (N_16833,N_12474,N_12315);
nor U16834 (N_16834,N_15210,N_13796);
and U16835 (N_16835,N_14613,N_15963);
nand U16836 (N_16836,N_15269,N_15915);
or U16837 (N_16837,N_15667,N_15085);
and U16838 (N_16838,N_14094,N_14522);
nand U16839 (N_16839,N_13523,N_14600);
nand U16840 (N_16840,N_12945,N_12374);
nand U16841 (N_16841,N_14425,N_13861);
or U16842 (N_16842,N_13842,N_13053);
nor U16843 (N_16843,N_12708,N_14599);
nand U16844 (N_16844,N_13468,N_12678);
or U16845 (N_16845,N_12488,N_12056);
nor U16846 (N_16846,N_12973,N_14722);
or U16847 (N_16847,N_13225,N_13657);
nor U16848 (N_16848,N_12493,N_13647);
nor U16849 (N_16849,N_15759,N_15676);
nor U16850 (N_16850,N_15582,N_13273);
nor U16851 (N_16851,N_12246,N_14084);
nor U16852 (N_16852,N_13120,N_15886);
nor U16853 (N_16853,N_14840,N_15840);
or U16854 (N_16854,N_12072,N_12979);
nand U16855 (N_16855,N_13735,N_13712);
and U16856 (N_16856,N_15308,N_13539);
and U16857 (N_16857,N_12805,N_13848);
or U16858 (N_16858,N_15744,N_13705);
or U16859 (N_16859,N_12057,N_13089);
xor U16860 (N_16860,N_15021,N_12854);
nor U16861 (N_16861,N_15415,N_15792);
and U16862 (N_16862,N_14670,N_13926);
or U16863 (N_16863,N_13857,N_14217);
nand U16864 (N_16864,N_12460,N_14988);
nor U16865 (N_16865,N_15821,N_14874);
or U16866 (N_16866,N_15519,N_14391);
nand U16867 (N_16867,N_15511,N_13685);
nand U16868 (N_16868,N_14146,N_14621);
nand U16869 (N_16869,N_13697,N_14669);
or U16870 (N_16870,N_12955,N_13581);
or U16871 (N_16871,N_13469,N_15241);
nor U16872 (N_16872,N_15809,N_15124);
or U16873 (N_16873,N_14614,N_15180);
and U16874 (N_16874,N_15095,N_13302);
or U16875 (N_16875,N_13985,N_12323);
or U16876 (N_16876,N_15881,N_13461);
and U16877 (N_16877,N_14827,N_15472);
or U16878 (N_16878,N_15437,N_13602);
and U16879 (N_16879,N_12793,N_14778);
and U16880 (N_16880,N_13759,N_12451);
xnor U16881 (N_16881,N_12699,N_14015);
or U16882 (N_16882,N_12129,N_12304);
nor U16883 (N_16883,N_15851,N_12379);
or U16884 (N_16884,N_12901,N_13831);
nand U16885 (N_16885,N_14665,N_13689);
nor U16886 (N_16886,N_15901,N_12439);
or U16887 (N_16887,N_14444,N_14255);
nand U16888 (N_16888,N_14138,N_15940);
nand U16889 (N_16889,N_13667,N_15951);
nand U16890 (N_16890,N_13146,N_13516);
or U16891 (N_16891,N_12054,N_13800);
nand U16892 (N_16892,N_12638,N_15830);
and U16893 (N_16893,N_15125,N_14925);
nand U16894 (N_16894,N_14364,N_14929);
nand U16895 (N_16895,N_14532,N_14330);
nor U16896 (N_16896,N_14017,N_12797);
or U16897 (N_16897,N_15587,N_15794);
and U16898 (N_16898,N_14578,N_13714);
and U16899 (N_16899,N_13080,N_13309);
or U16900 (N_16900,N_14980,N_14381);
and U16901 (N_16901,N_12624,N_13033);
nand U16902 (N_16902,N_13157,N_14806);
or U16903 (N_16903,N_12673,N_13510);
nor U16904 (N_16904,N_13339,N_15318);
or U16905 (N_16905,N_12243,N_15503);
xor U16906 (N_16906,N_14581,N_12895);
nor U16907 (N_16907,N_12659,N_13233);
nand U16908 (N_16908,N_14388,N_14327);
or U16909 (N_16909,N_12516,N_14662);
nor U16910 (N_16910,N_13155,N_14402);
or U16911 (N_16911,N_15109,N_14534);
nand U16912 (N_16912,N_15287,N_12178);
or U16913 (N_16913,N_14313,N_12404);
nor U16914 (N_16914,N_12103,N_14967);
nor U16915 (N_16915,N_15059,N_13356);
and U16916 (N_16916,N_13152,N_15386);
and U16917 (N_16917,N_13565,N_12941);
or U16918 (N_16918,N_13000,N_14143);
nand U16919 (N_16919,N_15079,N_12692);
nand U16920 (N_16920,N_14477,N_14279);
nand U16921 (N_16921,N_15028,N_12766);
nor U16922 (N_16922,N_14821,N_12492);
or U16923 (N_16923,N_13738,N_12862);
nand U16924 (N_16924,N_12284,N_14494);
and U16925 (N_16925,N_15208,N_15361);
and U16926 (N_16926,N_15965,N_15375);
nand U16927 (N_16927,N_13262,N_15646);
nand U16928 (N_16928,N_12723,N_13653);
nand U16929 (N_16929,N_15912,N_13537);
nor U16930 (N_16930,N_14096,N_15240);
or U16931 (N_16931,N_15338,N_12296);
xor U16932 (N_16932,N_15922,N_14439);
or U16933 (N_16933,N_13606,N_12400);
and U16934 (N_16934,N_13265,N_15323);
nor U16935 (N_16935,N_14816,N_13060);
nor U16936 (N_16936,N_12182,N_15750);
nand U16937 (N_16937,N_14871,N_15985);
or U16938 (N_16938,N_12446,N_13067);
and U16939 (N_16939,N_14366,N_13354);
xnor U16940 (N_16940,N_14019,N_14318);
or U16941 (N_16941,N_12959,N_13401);
or U16942 (N_16942,N_12248,N_12002);
nor U16943 (N_16943,N_14671,N_14731);
or U16944 (N_16944,N_15910,N_12763);
and U16945 (N_16945,N_15839,N_15041);
and U16946 (N_16946,N_12543,N_12807);
xnor U16947 (N_16947,N_13605,N_15884);
and U16948 (N_16948,N_13686,N_14351);
and U16949 (N_16949,N_15117,N_12351);
nand U16950 (N_16950,N_15136,N_13652);
nand U16951 (N_16951,N_12155,N_12588);
nand U16952 (N_16952,N_13418,N_15003);
xor U16953 (N_16953,N_15481,N_12785);
and U16954 (N_16954,N_14573,N_15065);
nor U16955 (N_16955,N_15462,N_13935);
xor U16956 (N_16956,N_12387,N_13278);
nor U16957 (N_16957,N_13936,N_14623);
or U16958 (N_16958,N_12519,N_12355);
nand U16959 (N_16959,N_13231,N_13783);
or U16960 (N_16960,N_12964,N_12397);
nor U16961 (N_16961,N_14065,N_14221);
nor U16962 (N_16962,N_13384,N_13275);
nor U16963 (N_16963,N_12210,N_13843);
nor U16964 (N_16964,N_14616,N_13064);
and U16965 (N_16965,N_12997,N_14179);
nor U16966 (N_16966,N_13615,N_13436);
nor U16967 (N_16967,N_15423,N_13224);
xor U16968 (N_16968,N_14655,N_15148);
or U16969 (N_16969,N_15533,N_14113);
and U16970 (N_16970,N_13386,N_15030);
and U16971 (N_16971,N_12890,N_12114);
xor U16972 (N_16972,N_12407,N_15242);
or U16973 (N_16973,N_15832,N_12032);
or U16974 (N_16974,N_15163,N_14057);
nand U16975 (N_16975,N_14112,N_13264);
nand U16976 (N_16976,N_15637,N_15419);
xnor U16977 (N_16977,N_12489,N_12333);
nor U16978 (N_16978,N_15938,N_14634);
nand U16979 (N_16979,N_14836,N_12750);
or U16980 (N_16980,N_12224,N_13691);
nor U16981 (N_16981,N_12984,N_14430);
or U16982 (N_16982,N_13122,N_12729);
or U16983 (N_16983,N_14651,N_15957);
nor U16984 (N_16984,N_15621,N_14503);
nand U16985 (N_16985,N_14618,N_12877);
nor U16986 (N_16986,N_13896,N_12468);
nor U16987 (N_16987,N_12268,N_12547);
and U16988 (N_16988,N_15042,N_15880);
nor U16989 (N_16989,N_13108,N_15093);
and U16990 (N_16990,N_13206,N_14851);
and U16991 (N_16991,N_12576,N_13631);
xor U16992 (N_16992,N_14786,N_12469);
xnor U16993 (N_16993,N_15190,N_14038);
nor U16994 (N_16994,N_14398,N_15891);
nand U16995 (N_16995,N_13471,N_15706);
nand U16996 (N_16996,N_12298,N_15201);
nand U16997 (N_16997,N_14596,N_14211);
nor U16998 (N_16998,N_12950,N_12335);
and U16999 (N_16999,N_14177,N_13996);
or U17000 (N_17000,N_13658,N_15869);
or U17001 (N_17001,N_12665,N_12879);
nand U17002 (N_17002,N_15206,N_15196);
nor U17003 (N_17003,N_14151,N_13478);
or U17004 (N_17004,N_14949,N_15088);
nand U17005 (N_17005,N_12761,N_12143);
nand U17006 (N_17006,N_14914,N_12573);
and U17007 (N_17007,N_15916,N_14441);
and U17008 (N_17008,N_14106,N_13504);
or U17009 (N_17009,N_12751,N_14517);
nand U17010 (N_17010,N_12947,N_13806);
nand U17011 (N_17011,N_13203,N_13760);
and U17012 (N_17012,N_13251,N_13087);
or U17013 (N_17013,N_13002,N_15826);
nor U17014 (N_17014,N_12411,N_13218);
and U17015 (N_17015,N_14976,N_12100);
nor U17016 (N_17016,N_13473,N_13693);
nor U17017 (N_17017,N_12219,N_13688);
nand U17018 (N_17018,N_13253,N_14431);
nand U17019 (N_17019,N_15541,N_12421);
nor U17020 (N_17020,N_15011,N_15494);
or U17021 (N_17021,N_15808,N_14696);
or U17022 (N_17022,N_14145,N_12864);
and U17023 (N_17023,N_12960,N_15232);
and U17024 (N_17024,N_13282,N_14587);
and U17025 (N_17025,N_14605,N_12124);
xor U17026 (N_17026,N_12216,N_14769);
nand U17027 (N_17027,N_14461,N_12555);
nor U17028 (N_17028,N_15544,N_12891);
nor U17029 (N_17029,N_15400,N_12876);
and U17030 (N_17030,N_12043,N_12534);
nor U17031 (N_17031,N_14278,N_13792);
and U17032 (N_17032,N_12063,N_13779);
nand U17033 (N_17033,N_13019,N_15151);
nand U17034 (N_17034,N_14903,N_12612);
and U17035 (N_17035,N_15723,N_15274);
and U17036 (N_17036,N_15062,N_14101);
or U17037 (N_17037,N_12589,N_13296);
or U17038 (N_17038,N_14240,N_15705);
or U17039 (N_17039,N_14457,N_12809);
xnor U17040 (N_17040,N_14878,N_15741);
or U17041 (N_17041,N_13915,N_13099);
and U17042 (N_17042,N_14699,N_14521);
or U17043 (N_17043,N_14979,N_14156);
nand U17044 (N_17044,N_12915,N_13609);
or U17045 (N_17045,N_14868,N_15161);
xor U17046 (N_17046,N_12410,N_15056);
or U17047 (N_17047,N_14884,N_14136);
or U17048 (N_17048,N_14575,N_12857);
and U17049 (N_17049,N_12201,N_13319);
nand U17050 (N_17050,N_15031,N_15892);
and U17051 (N_17051,N_13343,N_14261);
or U17052 (N_17052,N_13320,N_13818);
nand U17053 (N_17053,N_13368,N_12649);
nand U17054 (N_17054,N_13513,N_13765);
or U17055 (N_17055,N_14315,N_14203);
or U17056 (N_17056,N_13822,N_15853);
nor U17057 (N_17057,N_15107,N_12123);
and U17058 (N_17058,N_12948,N_12615);
or U17059 (N_17059,N_12028,N_12560);
nor U17060 (N_17060,N_12549,N_12646);
or U17061 (N_17061,N_15893,N_13824);
nor U17062 (N_17062,N_12067,N_12916);
or U17063 (N_17063,N_14384,N_12420);
and U17064 (N_17064,N_15496,N_13086);
nand U17065 (N_17065,N_12787,N_12015);
nand U17066 (N_17066,N_13419,N_15486);
nor U17067 (N_17067,N_13208,N_15239);
nor U17068 (N_17068,N_12297,N_15546);
or U17069 (N_17069,N_15797,N_13846);
or U17070 (N_17070,N_15285,N_15029);
nand U17071 (N_17071,N_14489,N_15025);
nor U17072 (N_17072,N_13402,N_15316);
nor U17073 (N_17073,N_15296,N_14213);
nor U17074 (N_17074,N_12084,N_15554);
nor U17075 (N_17075,N_15353,N_13424);
xnor U17076 (N_17076,N_15378,N_12413);
nor U17077 (N_17077,N_14230,N_14729);
nor U17078 (N_17078,N_15894,N_12272);
or U17079 (N_17079,N_14470,N_14673);
and U17080 (N_17080,N_13063,N_14380);
nor U17081 (N_17081,N_12187,N_13045);
nand U17082 (N_17082,N_12091,N_12684);
and U17083 (N_17083,N_12982,N_14632);
nor U17084 (N_17084,N_14040,N_15143);
nand U17085 (N_17085,N_15877,N_12329);
or U17086 (N_17086,N_15214,N_15430);
nand U17087 (N_17087,N_12048,N_13298);
or U17088 (N_17088,N_12738,N_14741);
xnor U17089 (N_17089,N_12172,N_15499);
nor U17090 (N_17090,N_12266,N_12835);
nand U17091 (N_17091,N_13104,N_15149);
and U17092 (N_17092,N_12166,N_12258);
xnor U17093 (N_17093,N_14897,N_12312);
xor U17094 (N_17094,N_14847,N_15529);
nor U17095 (N_17095,N_15515,N_13458);
and U17096 (N_17096,N_13706,N_13181);
and U17097 (N_17097,N_15489,N_13720);
or U17098 (N_17098,N_15182,N_13793);
nor U17099 (N_17099,N_12558,N_12904);
or U17100 (N_17100,N_14991,N_12806);
or U17101 (N_17101,N_15152,N_14423);
nor U17102 (N_17102,N_13867,N_15019);
and U17103 (N_17103,N_13904,N_12095);
and U17104 (N_17104,N_15370,N_12929);
nor U17105 (N_17105,N_15601,N_14353);
and U17106 (N_17106,N_13553,N_12934);
or U17107 (N_17107,N_12883,N_12595);
or U17108 (N_17108,N_14899,N_13125);
nor U17109 (N_17109,N_13034,N_15525);
and U17110 (N_17110,N_12666,N_14962);
or U17111 (N_17111,N_13744,N_12640);
and U17112 (N_17112,N_14462,N_14756);
or U17113 (N_17113,N_12770,N_14130);
nand U17114 (N_17114,N_15859,N_15944);
nor U17115 (N_17115,N_13508,N_13797);
and U17116 (N_17116,N_15975,N_14320);
and U17117 (N_17117,N_13970,N_12850);
xnor U17118 (N_17118,N_14188,N_12383);
nand U17119 (N_17119,N_14765,N_14551);
and U17120 (N_17120,N_12818,N_12535);
xor U17121 (N_17121,N_15878,N_14822);
and U17122 (N_17122,N_13672,N_14390);
nor U17123 (N_17123,N_13943,N_12307);
nor U17124 (N_17124,N_12671,N_14838);
nor U17125 (N_17125,N_15116,N_12435);
and U17126 (N_17126,N_12961,N_13016);
nand U17127 (N_17127,N_14947,N_14782);
and U17128 (N_17128,N_14157,N_12798);
nor U17129 (N_17129,N_15039,N_12762);
and U17130 (N_17130,N_13062,N_15131);
and U17131 (N_17131,N_12972,N_13334);
nor U17132 (N_17132,N_12016,N_14195);
or U17133 (N_17133,N_12886,N_15932);
or U17134 (N_17134,N_12326,N_13906);
and U17135 (N_17135,N_15168,N_15484);
xnor U17136 (N_17136,N_15959,N_15033);
nand U17137 (N_17137,N_13517,N_15123);
nand U17138 (N_17138,N_13951,N_12470);
nand U17139 (N_17139,N_12717,N_12801);
or U17140 (N_17140,N_12906,N_12542);
or U17141 (N_17141,N_15332,N_14760);
or U17142 (N_17142,N_12197,N_13399);
and U17143 (N_17143,N_13169,N_13106);
nor U17144 (N_17144,N_14588,N_14793);
nor U17145 (N_17145,N_14712,N_15291);
and U17146 (N_17146,N_12511,N_13600);
and U17147 (N_17147,N_13397,N_13737);
or U17148 (N_17148,N_14582,N_14448);
or U17149 (N_17149,N_15509,N_15627);
and U17150 (N_17150,N_14246,N_13702);
nor U17151 (N_17151,N_14241,N_15771);
nand U17152 (N_17152,N_15283,N_15113);
nor U17153 (N_17153,N_14689,N_13864);
or U17154 (N_17154,N_12384,N_13610);
and U17155 (N_17155,N_13236,N_14164);
nand U17156 (N_17156,N_12490,N_12991);
nand U17157 (N_17157,N_12218,N_15279);
xor U17158 (N_17158,N_15685,N_12926);
nor U17159 (N_17159,N_12824,N_12564);
or U17160 (N_17160,N_14495,N_15577);
nand U17161 (N_17161,N_12247,N_15470);
nor U17162 (N_17162,N_12270,N_15579);
or U17163 (N_17163,N_13427,N_15475);
or U17164 (N_17164,N_12395,N_15602);
nand U17165 (N_17165,N_15693,N_15382);
nand U17166 (N_17166,N_15825,N_15346);
xnor U17167 (N_17167,N_13487,N_13257);
or U17168 (N_17168,N_14963,N_12233);
nand U17169 (N_17169,N_13239,N_14864);
and U17170 (N_17170,N_14541,N_12466);
nand U17171 (N_17171,N_13194,N_12212);
or U17172 (N_17172,N_12827,N_15328);
nor U17173 (N_17173,N_13587,N_15082);
nand U17174 (N_17174,N_14504,N_13254);
nor U17175 (N_17175,N_15090,N_15907);
or U17176 (N_17176,N_15165,N_15063);
nor U17177 (N_17177,N_14686,N_12342);
nand U17178 (N_17178,N_14811,N_14684);
nor U17179 (N_17179,N_13011,N_12932);
and U17180 (N_17180,N_13102,N_14968);
or U17181 (N_17181,N_12506,N_14226);
nand U17182 (N_17182,N_15458,N_15523);
nor U17183 (N_17183,N_14570,N_14558);
xnor U17184 (N_17184,N_14029,N_15801);
xnor U17185 (N_17185,N_13185,N_15258);
nor U17186 (N_17186,N_13789,N_15611);
nor U17187 (N_17187,N_15074,N_14265);
nor U17188 (N_17188,N_15247,N_13147);
nor U17189 (N_17189,N_15528,N_14267);
nand U17190 (N_17190,N_12931,N_12502);
and U17191 (N_17191,N_12320,N_14535);
nand U17192 (N_17192,N_14537,N_15504);
nor U17193 (N_17193,N_15449,N_13624);
and U17194 (N_17194,N_15404,N_15272);
and U17195 (N_17195,N_14282,N_12340);
and U17196 (N_17196,N_14737,N_14270);
nand U17197 (N_17197,N_13700,N_12131);
and U17198 (N_17198,N_13976,N_15461);
and U17199 (N_17199,N_12828,N_14181);
or U17200 (N_17200,N_15046,N_15118);
nand U17201 (N_17201,N_13198,N_14627);
xnor U17202 (N_17202,N_14446,N_13819);
nor U17203 (N_17203,N_13052,N_12444);
nand U17204 (N_17204,N_12346,N_14850);
and U17205 (N_17205,N_12426,N_12249);
nor U17206 (N_17206,N_12026,N_14089);
nor U17207 (N_17207,N_12047,N_15977);
and U17208 (N_17208,N_12820,N_12104);
or U17209 (N_17209,N_14059,N_15605);
and U17210 (N_17210,N_14910,N_14611);
nand U17211 (N_17211,N_15870,N_12636);
nand U17212 (N_17212,N_13345,N_14041);
and U17213 (N_17213,N_14301,N_13571);
xnor U17214 (N_17214,N_15359,N_14251);
nand U17215 (N_17215,N_13380,N_12579);
nand U17216 (N_17216,N_15233,N_15964);
nand U17217 (N_17217,N_12070,N_12369);
or U17218 (N_17218,N_13682,N_14931);
or U17219 (N_17219,N_12747,N_15207);
nand U17220 (N_17220,N_12923,N_12361);
nand U17221 (N_17221,N_14938,N_14354);
and U17222 (N_17222,N_15615,N_12639);
nand U17223 (N_17223,N_14344,N_14788);
and U17224 (N_17224,N_15992,N_12606);
nor U17225 (N_17225,N_14097,N_14458);
and U17226 (N_17226,N_13756,N_14941);
and U17227 (N_17227,N_13911,N_14617);
and U17228 (N_17228,N_13332,N_13638);
or U17229 (N_17229,N_12110,N_14010);
nand U17230 (N_17230,N_13498,N_12116);
xnor U17231 (N_17231,N_14937,N_15520);
or U17232 (N_17232,N_13502,N_15658);
and U17233 (N_17233,N_15455,N_14277);
nand U17234 (N_17234,N_13088,N_13090);
nand U17235 (N_17235,N_12465,N_14987);
xor U17236 (N_17236,N_13175,N_12302);
nand U17237 (N_17237,N_15223,N_15968);
nand U17238 (N_17238,N_14852,N_14776);
and U17239 (N_17239,N_12487,N_14992);
and U17240 (N_17240,N_12295,N_12604);
nand U17241 (N_17241,N_14424,N_14585);
nor U17242 (N_17242,N_14036,N_15584);
nor U17243 (N_17243,N_13870,N_13877);
nor U17244 (N_17244,N_15810,N_15768);
or U17245 (N_17245,N_15720,N_14103);
nand U17246 (N_17246,N_15572,N_15573);
nand U17247 (N_17247,N_12020,N_13301);
and U17248 (N_17248,N_15108,N_14421);
xnor U17249 (N_17249,N_13897,N_13750);
and U17250 (N_17250,N_13858,N_13420);
nand U17251 (N_17251,N_12088,N_12733);
and U17252 (N_17252,N_12583,N_14223);
nand U17253 (N_17253,N_13835,N_12578);
or U17254 (N_17254,N_15935,N_15270);
and U17255 (N_17255,N_14370,N_13013);
xor U17256 (N_17256,N_14081,N_15697);
and U17257 (N_17257,N_13983,N_14511);
and U17258 (N_17258,N_12385,N_15229);
or U17259 (N_17259,N_14276,N_15926);
nor U17260 (N_17260,N_14995,N_12310);
xnor U17261 (N_17261,N_12153,N_13017);
and U17262 (N_17262,N_15115,N_14185);
or U17263 (N_17263,N_14045,N_15038);
nand U17264 (N_17264,N_15863,N_12643);
nand U17265 (N_17265,N_12039,N_12587);
or U17266 (N_17266,N_14990,N_15013);
nand U17267 (N_17267,N_15238,N_13585);
nand U17268 (N_17268,N_15596,N_12591);
xnor U17269 (N_17269,N_14309,N_15334);
nor U17270 (N_17270,N_14386,N_13490);
and U17271 (N_17271,N_14077,N_12055);
and U17272 (N_17272,N_15652,N_12563);
nor U17273 (N_17273,N_13409,N_14021);
nand U17274 (N_17274,N_13616,N_15681);
nand U17275 (N_17275,N_13863,N_13967);
or U17276 (N_17276,N_15854,N_13777);
nand U17277 (N_17277,N_13681,N_14227);
nand U17278 (N_17278,N_13154,N_15144);
and U17279 (N_17279,N_12316,N_15714);
xnor U17280 (N_17280,N_15231,N_14918);
or U17281 (N_17281,N_14619,N_14078);
nand U17282 (N_17282,N_12529,N_13696);
nor U17283 (N_17283,N_14660,N_12966);
nor U17284 (N_17284,N_13023,N_13956);
nor U17285 (N_17285,N_12171,N_13727);
nor U17286 (N_17286,N_15746,N_15103);
or U17287 (N_17287,N_14093,N_12107);
nand U17288 (N_17288,N_12918,N_14180);
nor U17289 (N_17289,N_12771,N_13394);
nand U17290 (N_17290,N_13690,N_13500);
nand U17291 (N_17291,N_13540,N_12352);
xor U17292 (N_17292,N_15060,N_14626);
or U17293 (N_17293,N_13280,N_13482);
xnor U17294 (N_17294,N_15896,N_15372);
and U17295 (N_17295,N_13859,N_14160);
and U17296 (N_17296,N_14679,N_15147);
or U17297 (N_17297,N_13868,N_14236);
or U17298 (N_17298,N_12094,N_14728);
nor U17299 (N_17299,N_14117,N_15545);
nand U17300 (N_17300,N_12748,N_12603);
nor U17301 (N_17301,N_14175,N_15689);
nand U17302 (N_17302,N_14924,N_13621);
xnor U17303 (N_17303,N_14872,N_14328);
nand U17304 (N_17304,N_14996,N_12261);
nor U17305 (N_17305,N_12860,N_14373);
nand U17306 (N_17306,N_14597,N_14960);
nor U17307 (N_17307,N_15743,N_13018);
nand U17308 (N_17308,N_12359,N_13876);
nor U17309 (N_17309,N_13561,N_14676);
and U17310 (N_17310,N_15336,N_15650);
xor U17311 (N_17311,N_15215,N_14698);
and U17312 (N_17312,N_15538,N_12765);
or U17313 (N_17313,N_13178,N_15629);
nor U17314 (N_17314,N_13820,N_12303);
nand U17315 (N_17315,N_12120,N_15034);
nor U17316 (N_17316,N_15943,N_14429);
nand U17317 (N_17317,N_12105,N_13170);
and U17318 (N_17318,N_13614,N_14258);
nand U17319 (N_17319,N_13664,N_12782);
nor U17320 (N_17320,N_12211,N_14710);
or U17321 (N_17321,N_13829,N_12240);
and U17322 (N_17322,N_14569,N_14909);
nand U17323 (N_17323,N_14707,N_12082);
and U17324 (N_17324,N_15931,N_15639);
and U17325 (N_17325,N_13232,N_15505);
or U17326 (N_17326,N_14049,N_14484);
or U17327 (N_17327,N_15098,N_14912);
or U17328 (N_17328,N_13404,N_13324);
xor U17329 (N_17329,N_12889,N_14648);
and U17330 (N_17330,N_15569,N_12822);
or U17331 (N_17331,N_13084,N_15694);
nor U17332 (N_17332,N_13544,N_13994);
nand U17333 (N_17333,N_15802,N_12189);
nand U17334 (N_17334,N_12633,N_15550);
nor U17335 (N_17335,N_12540,N_13311);
or U17336 (N_17336,N_13355,N_12949);
or U17337 (N_17337,N_12274,N_13491);
nand U17338 (N_17338,N_12473,N_12683);
and U17339 (N_17339,N_12530,N_14989);
and U17340 (N_17340,N_14633,N_12548);
nor U17341 (N_17341,N_13514,N_13435);
or U17342 (N_17342,N_13977,N_13046);
and U17343 (N_17343,N_14981,N_13577);
or U17344 (N_17344,N_13598,N_14681);
nor U17345 (N_17345,N_13535,N_15701);
nor U17346 (N_17346,N_14723,N_13684);
and U17347 (N_17347,N_14738,N_12825);
nor U17348 (N_17348,N_14499,N_12217);
and U17349 (N_17349,N_12938,N_13666);
nand U17350 (N_17350,N_13130,N_14846);
or U17351 (N_17351,N_12513,N_14849);
and U17352 (N_17352,N_12336,N_13748);
and U17353 (N_17353,N_13780,N_15536);
xnor U17354 (N_17354,N_15500,N_15483);
and U17355 (N_17355,N_12199,N_14753);
and U17356 (N_17356,N_13151,N_13333);
xnor U17357 (N_17357,N_15664,N_15416);
nand U17358 (N_17358,N_13297,N_13851);
nand U17359 (N_17359,N_15227,N_13729);
or U17360 (N_17360,N_14879,N_15858);
or U17361 (N_17361,N_12565,N_15553);
nand U17362 (N_17362,N_12282,N_12654);
and U17363 (N_17363,N_15133,N_15925);
nor U17364 (N_17364,N_13695,N_15427);
nand U17365 (N_17365,N_13193,N_14104);
nand U17366 (N_17366,N_14571,N_13671);
nor U17367 (N_17367,N_13441,N_14468);
nor U17368 (N_17368,N_13398,N_13050);
nor U17369 (N_17369,N_12126,N_15010);
nand U17370 (N_17370,N_12967,N_15366);
or U17371 (N_17371,N_15248,N_12213);
nand U17372 (N_17372,N_13456,N_12040);
or U17373 (N_17373,N_13220,N_15321);
nor U17374 (N_17374,N_14148,N_15451);
nand U17375 (N_17375,N_12256,N_15710);
and U17376 (N_17376,N_15581,N_15875);
nand U17377 (N_17377,N_12953,N_13968);
nor U17378 (N_17378,N_14900,N_15645);
nor U17379 (N_17379,N_12503,N_13432);
and U17380 (N_17380,N_12976,N_14594);
and U17381 (N_17381,N_14281,N_15224);
or U17382 (N_17382,N_15914,N_13632);
or U17383 (N_17383,N_13325,N_12724);
or U17384 (N_17384,N_14075,N_14568);
xnor U17385 (N_17385,N_13788,N_12866);
nand U17386 (N_17386,N_14726,N_12035);
xor U17387 (N_17387,N_12392,N_14560);
nor U17388 (N_17388,N_15617,N_12344);
nor U17389 (N_17389,N_14073,N_14491);
xor U17390 (N_17390,N_14561,N_12975);
nor U17391 (N_17391,N_13790,N_15657);
and U17392 (N_17392,N_13785,N_14584);
nand U17393 (N_17393,N_15431,N_12993);
xor U17394 (N_17394,N_12514,N_14257);
nand U17395 (N_17395,N_15128,N_12687);
xor U17396 (N_17396,N_14030,N_14749);
nor U17397 (N_17397,N_13856,N_15948);
nor U17398 (N_17398,N_13713,N_15687);
or U17399 (N_17399,N_14321,N_15731);
nand U17400 (N_17400,N_14946,N_12433);
xnor U17401 (N_17401,N_15012,N_15776);
and U17402 (N_17402,N_14194,N_12059);
nor U17403 (N_17403,N_12205,N_15135);
or U17404 (N_17404,N_13519,N_12377);
nand U17405 (N_17405,N_12176,N_15594);
nor U17406 (N_17406,N_14552,N_15236);
nor U17407 (N_17407,N_14743,N_12899);
or U17408 (N_17408,N_12810,N_15114);
or U17409 (N_17409,N_12541,N_13295);
nand U17410 (N_17410,N_13179,N_12910);
nor U17411 (N_17411,N_12169,N_12265);
nand U17412 (N_17412,N_14927,N_14733);
nand U17413 (N_17413,N_14350,N_15045);
or U17414 (N_17414,N_13366,N_15711);
nand U17415 (N_17415,N_13543,N_12146);
nand U17416 (N_17416,N_12278,N_13562);
or U17417 (N_17417,N_14490,N_13929);
nand U17418 (N_17418,N_12415,N_14454);
and U17419 (N_17419,N_13582,N_12582);
nor U17420 (N_17420,N_14855,N_12757);
nand U17421 (N_17421,N_13781,N_12049);
nor U17422 (N_17422,N_12777,N_12037);
nor U17423 (N_17423,N_12324,N_13266);
xnor U17424 (N_17424,N_12215,N_13732);
and U17425 (N_17425,N_14238,N_12347);
nand U17426 (N_17426,N_12239,N_15383);
nor U17427 (N_17427,N_13942,N_14690);
xnor U17428 (N_17428,N_14629,N_12190);
nand U17429 (N_17429,N_14923,N_14220);
nor U17430 (N_17430,N_14129,N_14631);
and U17431 (N_17431,N_15718,N_13177);
nand U17432 (N_17432,N_13235,N_13914);
nand U17433 (N_17433,N_13414,N_13475);
nand U17434 (N_17434,N_15728,N_14086);
nand U17435 (N_17435,N_12238,N_13258);
or U17436 (N_17436,N_13629,N_12968);
nor U17437 (N_17437,N_13989,N_14892);
or U17438 (N_17438,N_13808,N_14948);
or U17439 (N_17439,N_15800,N_14516);
or U17440 (N_17440,N_14652,N_15856);
and U17441 (N_17441,N_12677,N_12940);
nand U17442 (N_17442,N_15600,N_15252);
or U17443 (N_17443,N_14705,N_12739);
xnor U17444 (N_17444,N_13895,N_12257);
xnor U17445 (N_17445,N_14727,N_14512);
or U17446 (N_17446,N_15735,N_12106);
nand U17447 (N_17447,N_13073,N_13677);
and U17448 (N_17448,N_13287,N_14058);
nor U17449 (N_17449,N_13885,N_13991);
and U17450 (N_17450,N_12928,N_12196);
or U17451 (N_17451,N_14287,N_15501);
nor U17452 (N_17452,N_12718,N_13619);
or U17453 (N_17453,N_13555,N_14640);
or U17454 (N_17454,N_13438,N_12607);
nor U17455 (N_17455,N_12077,N_13823);
nor U17456 (N_17456,N_14253,N_14014);
nand U17457 (N_17457,N_13802,N_15631);
or U17458 (N_17458,N_14908,N_12089);
and U17459 (N_17459,N_15412,N_13811);
and U17460 (N_17460,N_14907,N_13156);
nand U17461 (N_17461,N_14556,N_15183);
xor U17462 (N_17462,N_12773,N_15960);
xor U17463 (N_17463,N_15043,N_14187);
and U17464 (N_17464,N_15301,N_14502);
and U17465 (N_17465,N_15758,N_14972);
nand U17466 (N_17466,N_14362,N_15585);
nand U17467 (N_17467,N_12694,N_15521);
or U17468 (N_17468,N_13182,N_14813);
nor U17469 (N_17469,N_13217,N_13721);
or U17470 (N_17470,N_13136,N_14678);
nor U17471 (N_17471,N_13202,N_15990);
and U17472 (N_17472,N_13528,N_14694);
nand U17473 (N_17473,N_15876,N_15675);
and U17474 (N_17474,N_13168,N_15058);
nor U17475 (N_17475,N_15981,N_13998);
nand U17476 (N_17476,N_13403,N_14214);
or U17477 (N_17477,N_12884,N_13374);
nor U17478 (N_17478,N_13880,N_13518);
nand U17479 (N_17479,N_12875,N_14124);
nand U17480 (N_17480,N_13003,N_14835);
or U17481 (N_17481,N_12608,N_13075);
and U17482 (N_17482,N_12758,N_14609);
nand U17483 (N_17483,N_15277,N_14063);
nand U17484 (N_17484,N_12362,N_13844);
and U17485 (N_17485,N_14935,N_13221);
and U17486 (N_17486,N_14445,N_15181);
nor U17487 (N_17487,N_12623,N_14443);
or U17488 (N_17488,N_15280,N_15976);
or U17489 (N_17489,N_13250,N_12551);
nand U17490 (N_17490,N_12245,N_15364);
or U17491 (N_17491,N_12722,N_14540);
and U17492 (N_17492,N_13281,N_15092);
and U17493 (N_17493,N_13445,N_14735);
and U17494 (N_17494,N_12370,N_15857);
and U17495 (N_17495,N_15927,N_15406);
and U17496 (N_17496,N_14047,N_13274);
nor U17497 (N_17497,N_13361,N_15805);
nand U17498 (N_17498,N_12121,N_12286);
nor U17499 (N_17499,N_13448,N_15630);
nor U17500 (N_17500,N_14455,N_12406);
and U17501 (N_17501,N_14954,N_13728);
or U17502 (N_17502,N_15036,N_15626);
nand U17503 (N_17503,N_14182,N_13457);
xor U17504 (N_17504,N_13973,N_12428);
or U17505 (N_17505,N_14734,N_14254);
nor U17506 (N_17506,N_15766,N_12119);
nand U17507 (N_17507,N_14183,N_13934);
or U17508 (N_17508,N_12078,N_15403);
xor U17509 (N_17509,N_13285,N_15080);
nor U17510 (N_17510,N_13962,N_13912);
or U17511 (N_17511,N_12194,N_12726);
nand U17512 (N_17512,N_13428,N_15518);
and U17513 (N_17513,N_13031,N_12691);
nand U17514 (N_17514,N_13515,N_14860);
nor U17515 (N_17515,N_14248,N_15552);
nor U17516 (N_17516,N_12676,N_12742);
nor U17517 (N_17517,N_13158,N_12598);
xor U17518 (N_17518,N_14466,N_13618);
and U17519 (N_17519,N_15048,N_14939);
and U17520 (N_17520,N_12011,N_15237);
and U17521 (N_17521,N_13656,N_15986);
nor U17522 (N_17522,N_13764,N_13889);
and U17523 (N_17523,N_12019,N_15220);
nor U17524 (N_17524,N_15425,N_12452);
or U17525 (N_17525,N_15244,N_12594);
nand U17526 (N_17526,N_15988,N_14024);
nor U17527 (N_17527,N_12912,N_13804);
nand U17528 (N_17528,N_13527,N_15918);
xor U17529 (N_17529,N_15684,N_15571);
nor U17530 (N_17530,N_13323,N_13757);
or U17531 (N_17531,N_13248,N_13719);
nor U17532 (N_17532,N_14715,N_12527);
nor U17533 (N_17533,N_13836,N_14150);
and U17534 (N_17534,N_15089,N_13042);
and U17535 (N_17535,N_15132,N_14054);
or U17536 (N_17536,N_12242,N_12714);
nand U17537 (N_17537,N_14198,N_14604);
and U17538 (N_17538,N_15493,N_14285);
nor U17539 (N_17539,N_13048,N_14703);
and U17540 (N_17540,N_12645,N_14460);
nor U17541 (N_17541,N_14817,N_14283);
nor U17542 (N_17542,N_15446,N_14109);
or U17543 (N_17543,N_12845,N_14858);
nor U17544 (N_17544,N_12051,N_12688);
and U17545 (N_17545,N_13736,N_15130);
and U17546 (N_17546,N_13570,N_15656);
nand U17547 (N_17547,N_13630,N_12725);
nand U17548 (N_17548,N_15749,N_12614);
and U17549 (N_17549,N_15195,N_14229);
nand U17550 (N_17550,N_15226,N_15709);
nand U17551 (N_17551,N_14664,N_12620);
nand U17552 (N_17552,N_13734,N_14863);
and U17553 (N_17553,N_12448,N_15191);
nor U17554 (N_17554,N_13534,N_14405);
xnor U17555 (N_17555,N_14620,N_13008);
nand U17556 (N_17556,N_15072,N_12792);
nand U17557 (N_17557,N_14768,N_15466);
nor U17558 (N_17558,N_12784,N_12522);
and U17559 (N_17559,N_12833,N_13987);
or U17560 (N_17560,N_12064,N_14607);
nor U17561 (N_17561,N_13910,N_12437);
nand U17562 (N_17562,N_15087,N_13246);
nor U17563 (N_17563,N_12577,N_12111);
or U17564 (N_17564,N_12537,N_14154);
nor U17565 (N_17565,N_12389,N_12052);
or U17566 (N_17566,N_13798,N_15185);
and U17567 (N_17567,N_12409,N_12198);
nor U17568 (N_17568,N_12177,N_12701);
nor U17569 (N_17569,N_13061,N_15335);
nor U17570 (N_17570,N_15514,N_13431);
xnor U17571 (N_17571,N_14403,N_15852);
or U17572 (N_17572,N_14341,N_14481);
or U17573 (N_17573,N_15257,N_13094);
nor U17574 (N_17574,N_15604,N_12273);
and U17575 (N_17575,N_13133,N_15903);
nand U17576 (N_17576,N_13984,N_15314);
nor U17577 (N_17577,N_14436,N_12150);
nor U17578 (N_17578,N_13107,N_12202);
or U17579 (N_17579,N_13243,N_12831);
and U17580 (N_17580,N_13974,N_15804);
nor U17581 (N_17581,N_13314,N_13803);
nor U17582 (N_17582,N_13346,N_14866);
nor U17583 (N_17583,N_15426,N_12269);
nor U17584 (N_17584,N_14873,N_14308);
or U17585 (N_17585,N_13071,N_13149);
or U17586 (N_17586,N_12280,N_14323);
nor U17587 (N_17587,N_14412,N_13787);
nor U17588 (N_17588,N_12814,N_13360);
or U17589 (N_17589,N_15371,N_12767);
or U17590 (N_17590,N_15275,N_14378);
or U17591 (N_17591,N_15487,N_12461);
and U17592 (N_17592,N_15649,N_12069);
nand U17593 (N_17593,N_13015,N_12075);
nand U17594 (N_17594,N_14239,N_12958);
xor U17595 (N_17595,N_13400,N_14709);
or U17596 (N_17596,N_14547,N_13752);
or U17597 (N_17597,N_14695,N_12022);
nor U17598 (N_17598,N_12394,N_15712);
nand U17599 (N_17599,N_14896,N_13883);
or U17600 (N_17600,N_13300,N_14166);
and U17601 (N_17601,N_14898,N_14606);
and U17602 (N_17602,N_13611,N_14172);
and U17603 (N_17603,N_14802,N_14982);
and U17604 (N_17604,N_12079,N_12515);
nand U17605 (N_17605,N_14206,N_14212);
nor U17606 (N_17606,N_12995,N_12425);
nand U17607 (N_17607,N_12161,N_15819);
and U17608 (N_17608,N_12112,N_12141);
nand U17609 (N_17609,N_14739,N_14289);
and U17610 (N_17610,N_15078,N_15473);
and U17611 (N_17611,N_14834,N_12158);
nand U17612 (N_17612,N_13503,N_15654);
nand U17613 (N_17613,N_13148,N_14586);
xor U17614 (N_17614,N_13495,N_13922);
and U17615 (N_17615,N_14463,N_13673);
or U17616 (N_17616,N_14984,N_12897);
nor U17617 (N_17617,N_14050,N_13538);
nor U17618 (N_17618,N_12167,N_14759);
xor U17619 (N_17619,N_12322,N_13925);
and U17620 (N_17620,N_14105,N_13531);
xor U17621 (N_17621,N_15765,N_15294);
or U17622 (N_17622,N_12882,N_12354);
nor U17623 (N_17623,N_12414,N_14969);
nor U17624 (N_17624,N_12944,N_13054);
and U17625 (N_17625,N_12602,N_12263);
nor U17626 (N_17626,N_14680,N_12481);
or U17627 (N_17627,N_15679,N_15052);
nor U17628 (N_17628,N_14348,N_12992);
nor U17629 (N_17629,N_12552,N_13933);
or U17630 (N_17630,N_13725,N_15775);
nor U17631 (N_17631,N_12802,N_14763);
and U17632 (N_17632,N_13166,N_14361);
nand U17633 (N_17633,N_15488,N_12500);
nand U17634 (N_17634,N_14563,N_13268);
or U17635 (N_17635,N_15037,N_15460);
nand U17636 (N_17636,N_15595,N_14755);
or U17637 (N_17637,N_13362,N_12250);
or U17638 (N_17638,N_15160,N_12496);
nor U17639 (N_17639,N_12237,N_14580);
or U17640 (N_17640,N_15268,N_15849);
nor U17641 (N_17641,N_12330,N_15583);
nor U17642 (N_17642,N_15465,N_12004);
and U17643 (N_17643,N_14649,N_13708);
and U17644 (N_17644,N_12705,N_13390);
or U17645 (N_17645,N_14657,N_12173);
xnor U17646 (N_17646,N_13564,N_15409);
or U17647 (N_17647,N_14538,N_15482);
or U17648 (N_17648,N_12789,N_15924);
or U17649 (N_17649,N_15384,N_13030);
or U17650 (N_17650,N_13489,N_14509);
or U17651 (N_17651,N_15773,N_13908);
and U17652 (N_17652,N_12134,N_15945);
nand U17653 (N_17653,N_15899,N_14761);
nor U17654 (N_17654,N_15000,N_15713);
or U17655 (N_17655,N_12485,N_14478);
and U17656 (N_17656,N_13036,N_14061);
nand U17657 (N_17657,N_13330,N_12151);
and U17658 (N_17658,N_12631,N_14986);
and U17659 (N_17659,N_12267,N_14624);
nand U17660 (N_17660,N_12985,N_15167);
and U17661 (N_17661,N_12491,N_14170);
or U17662 (N_17662,N_13497,N_12356);
or U17663 (N_17663,N_12597,N_15898);
or U17664 (N_17664,N_13454,N_14438);
nand U17665 (N_17665,N_12008,N_12450);
and U17666 (N_17666,N_14877,N_14965);
nand U17667 (N_17667,N_14303,N_12285);
nand U17668 (N_17668,N_13938,N_12372);
nand U17669 (N_17669,N_13044,N_12501);
xor U17670 (N_17670,N_12936,N_14865);
xor U17671 (N_17671,N_15373,N_12867);
and U17672 (N_17672,N_14635,N_15855);
xor U17673 (N_17673,N_13446,N_12745);
or U17674 (N_17674,N_15156,N_12970);
nor U17675 (N_17675,N_12376,N_13114);
or U17676 (N_17676,N_14589,N_13039);
nor U17677 (N_17677,N_15395,N_15254);
nor U17678 (N_17678,N_13853,N_15703);
or U17679 (N_17679,N_15761,N_13470);
xor U17680 (N_17680,N_14615,N_15343);
or U17681 (N_17681,N_12455,N_14396);
nand U17682 (N_17682,N_13007,N_12730);
or U17683 (N_17683,N_12786,N_15955);
and U17684 (N_17684,N_14754,N_15126);
nor U17685 (N_17685,N_13357,N_14977);
or U17686 (N_17686,N_14271,N_14891);
and U17687 (N_17687,N_13288,N_15846);
nand U17688 (N_17688,N_14645,N_12441);
xor U17689 (N_17689,N_15865,N_15929);
or U17690 (N_17690,N_15317,N_13382);
xnor U17691 (N_17691,N_13944,N_12813);
and U17692 (N_17692,N_15388,N_12358);
and U17693 (N_17693,N_14393,N_15946);
nor U17694 (N_17694,N_13290,N_14451);
nor U17695 (N_17695,N_13952,N_13986);
nand U17696 (N_17696,N_13379,N_15219);
or U17697 (N_17697,N_13981,N_15770);
or U17698 (N_17698,N_15752,N_13969);
xor U17699 (N_17699,N_14039,N_15717);
xor U17700 (N_17700,N_14692,N_15407);
and U17701 (N_17701,N_14601,N_13589);
or U17702 (N_17702,N_14404,N_13113);
nor U17703 (N_17703,N_14940,N_14272);
or U17704 (N_17704,N_13724,N_14135);
nor U17705 (N_17705,N_12925,N_13845);
nor U17706 (N_17706,N_15097,N_15245);
nand U17707 (N_17707,N_12127,N_14133);
or U17708 (N_17708,N_15708,N_15522);
and U17709 (N_17709,N_14333,N_12821);
nor U17710 (N_17710,N_15836,N_15053);
or U17711 (N_17711,N_14216,N_13160);
and U17712 (N_17712,N_14544,N_15137);
nand U17713 (N_17713,N_14639,N_15967);
nor U17714 (N_17714,N_12622,N_15164);
or U17715 (N_17715,N_14199,N_15789);
and U17716 (N_17716,N_12592,N_14202);
nand U17717 (N_17717,N_15057,N_12003);
and U17718 (N_17718,N_12287,N_15311);
nor U17719 (N_17719,N_12674,N_14957);
nand U17720 (N_17720,N_12715,N_12728);
and U17721 (N_17721,N_15837,N_15303);
nor U17722 (N_17722,N_12703,N_12655);
and U17723 (N_17723,N_14072,N_13990);
nand U17724 (N_17724,N_15312,N_12007);
and U17725 (N_17725,N_15432,N_15121);
nor U17726 (N_17726,N_13551,N_12180);
nor U17727 (N_17727,N_15642,N_12045);
and U17728 (N_17728,N_15980,N_15578);
nor U17729 (N_17729,N_14329,N_15671);
nor U17730 (N_17730,N_15162,N_13100);
nor U17731 (N_17731,N_14777,N_12313);
nand U17732 (N_17732,N_13849,N_12068);
nand U17733 (N_17733,N_13786,N_13754);
xnor U17734 (N_17734,N_12885,N_15339);
or U17735 (N_17735,N_15974,N_12667);
or U17736 (N_17736,N_14107,N_12309);
nand U17737 (N_17737,N_15331,N_12783);
nand U17738 (N_17738,N_12208,N_15669);
and U17739 (N_17739,N_13709,N_15724);
nor U17740 (N_17740,N_14719,N_13648);
nand U17741 (N_17741,N_14598,N_12200);
and U17742 (N_17742,N_13167,N_14577);
nand U17743 (N_17743,N_15790,N_15171);
nand U17744 (N_17744,N_13763,N_15506);
and U17745 (N_17745,N_15178,N_13882);
xnor U17746 (N_17746,N_14576,N_15150);
nand U17747 (N_17747,N_14062,N_14299);
or U17748 (N_17748,N_14416,N_14774);
and U17749 (N_17749,N_14476,N_12025);
nand U17750 (N_17750,N_13187,N_12924);
nor U17751 (N_17751,N_14518,N_14335);
or U17752 (N_17752,N_14766,N_12584);
xnor U17753 (N_17753,N_13546,N_12946);
or U17754 (N_17754,N_12690,N_14825);
nand U17755 (N_17755,N_12956,N_13554);
nor U17756 (N_17756,N_13900,N_15672);
nand U17757 (N_17757,N_12449,N_15566);
nand U17758 (N_17758,N_14219,N_12653);
nand U17759 (N_17759,N_14890,N_12092);
and U17760 (N_17760,N_12613,N_13769);
and U17761 (N_17761,N_14387,N_13442);
or U17762 (N_17762,N_13982,N_14554);
nor U17763 (N_17763,N_13746,N_15249);
nor U17764 (N_17764,N_13654,N_14545);
nand U17765 (N_17765,N_12348,N_14498);
xor U17766 (N_17766,N_14798,N_15464);
and U17767 (N_17767,N_14184,N_15381);
or U17768 (N_17768,N_14256,N_14497);
nand U17769 (N_17769,N_14007,N_15354);
nor U17770 (N_17770,N_14474,N_14809);
or U17771 (N_17771,N_13335,N_15763);
or U17772 (N_17772,N_12856,N_12980);
xnor U17773 (N_17773,N_12575,N_15942);
or U17774 (N_17774,N_13286,N_13694);
or U17775 (N_17775,N_14352,N_15557);
nand U17776 (N_17776,N_14171,N_12128);
nand U17777 (N_17777,N_15068,N_14046);
or U17778 (N_17778,N_15433,N_13141);
xnor U17779 (N_17779,N_12842,N_12108);
nand U17780 (N_17780,N_12518,N_15635);
and U17781 (N_17781,N_14450,N_12811);
nand U17782 (N_17782,N_12781,N_13410);
nand U17783 (N_17783,N_14803,N_13117);
and U17784 (N_17784,N_13391,N_15369);
nand U17785 (N_17785,N_13670,N_14023);
or U17786 (N_17786,N_13480,N_14292);
or U17787 (N_17787,N_12207,N_14070);
or U17788 (N_17788,N_15008,N_13439);
nand U17789 (N_17789,N_12570,N_14857);
or U17790 (N_17790,N_12476,N_13367);
nor U17791 (N_17791,N_14176,N_15356);
nor U17792 (N_17792,N_14943,N_14178);
nor U17793 (N_17793,N_14031,N_12031);
nor U17794 (N_17794,N_12851,N_14379);
nor U17795 (N_17795,N_13481,N_12696);
nand U17796 (N_17796,N_14120,N_15216);
xnor U17797 (N_17797,N_12632,N_15739);
nor U17798 (N_17798,N_12475,N_15408);
nand U17799 (N_17799,N_15580,N_13358);
nor U17800 (N_17800,N_13683,N_12334);
or U17801 (N_17801,N_13093,N_13022);
nand U17802 (N_17802,N_15230,N_14542);
xor U17803 (N_17803,N_15186,N_12457);
nand U17804 (N_17804,N_14337,N_14452);
nand U17805 (N_17805,N_13568,N_14006);
xor U17806 (N_17806,N_12311,N_15023);
or U17807 (N_17807,N_15632,N_14076);
and U17808 (N_17808,N_15016,N_14823);
or U17809 (N_17809,N_13312,N_12599);
and U17810 (N_17810,N_13032,N_12228);
nand U17811 (N_17811,N_12927,N_13024);
and U17812 (N_17812,N_15966,N_12544);
xor U17813 (N_17813,N_15983,N_13874);
xnor U17814 (N_17814,N_14654,N_15193);
or U17815 (N_17815,N_14510,N_13993);
nand U17816 (N_17816,N_15325,N_15603);
or U17817 (N_17817,N_12779,N_14392);
or U17818 (N_17818,N_12580,N_12621);
or U17819 (N_17819,N_12550,N_13903);
xnor U17820 (N_17820,N_12619,N_14882);
nor U17821 (N_17821,N_13111,N_13337);
and U17822 (N_17822,N_13520,N_14197);
and U17823 (N_17823,N_12769,N_15352);
or U17824 (N_17824,N_13127,N_15006);
or U17825 (N_17825,N_15225,N_14174);
or U17826 (N_17826,N_14528,N_12969);
nor U17827 (N_17827,N_15704,N_12942);
or U17828 (N_17828,N_13072,N_14505);
xnor U17829 (N_17829,N_14080,N_14488);
nand U17830 (N_17830,N_14675,N_13762);
nor U17831 (N_17831,N_15551,N_13778);
nor U17832 (N_17832,N_12788,N_13722);
nand U17833 (N_17833,N_15570,N_13085);
nor U17834 (N_17834,N_13680,N_14916);
nand U17835 (N_17835,N_14245,N_14355);
or U17836 (N_17836,N_12145,N_12709);
nand U17837 (N_17837,N_15463,N_13138);
nor U17838 (N_17838,N_13655,N_12462);
nand U17839 (N_17839,N_15221,N_13396);
nand U17840 (N_17840,N_14736,N_14419);
nand U17841 (N_17841,N_15454,N_14810);
nand U17842 (N_17842,N_14998,N_15174);
nor U17843 (N_17843,N_12229,N_13633);
nand U17844 (N_17844,N_14773,N_15558);
nor U17845 (N_17845,N_13299,N_12283);
and U17846 (N_17846,N_12965,N_13761);
nor U17847 (N_17847,N_15599,N_15418);
nor U17848 (N_17848,N_12459,N_15795);
xnor U17849 (N_17849,N_14401,N_14674);
nor U17850 (N_17850,N_13572,N_12231);
nand U17851 (N_17851,N_14428,N_12188);
nand U17852 (N_17852,N_12357,N_13037);
nor U17853 (N_17853,N_13012,N_12803);
and U17854 (N_17854,N_14155,N_15184);
xnor U17855 (N_17855,N_14294,N_12164);
xnor U17856 (N_17856,N_15695,N_13200);
nand U17857 (N_17857,N_13767,N_12905);
xor U17858 (N_17858,N_12341,N_13180);
nor U17859 (N_17859,N_14012,N_13827);
nor U17860 (N_17860,N_14274,N_12338);
nor U17861 (N_17861,N_13753,N_14319);
nor U17862 (N_17862,N_13997,N_15610);
nand U17863 (N_17863,N_12504,N_14360);
xnor U17864 (N_17864,N_14829,N_15474);
nor U17865 (N_17865,N_15883,N_14794);
nand U17866 (N_17866,N_15620,N_14442);
nand U17867 (N_17867,N_13839,N_13566);
or U17868 (N_17868,N_13739,N_13150);
nor U17869 (N_17869,N_13841,N_12434);
nand U17870 (N_17870,N_12279,N_13825);
nor U17871 (N_17871,N_12922,N_14471);
xor U17872 (N_17872,N_14902,N_15050);
nand U17873 (N_17873,N_15348,N_15625);
nand U17874 (N_17874,N_15387,N_14867);
and U17875 (N_17875,N_12795,N_12149);
and U17876 (N_17876,N_15612,N_15683);
and U17877 (N_17877,N_15780,N_13129);
nor U17878 (N_17878,N_12731,N_13865);
and U17879 (N_17879,N_13124,N_15389);
or U17880 (N_17880,N_15476,N_12702);
xnor U17881 (N_17881,N_12305,N_15873);
xor U17882 (N_17882,N_14783,N_13715);
nor U17883 (N_17883,N_14883,N_15411);
and U17884 (N_17884,N_12328,N_13636);
nor U17885 (N_17885,N_12277,N_14232);
xor U17886 (N_17886,N_15350,N_12609);
or U17887 (N_17887,N_13307,N_14565);
nor U17888 (N_17888,N_12438,N_13153);
nand U17889 (N_17889,N_15324,N_14830);
nor U17890 (N_17890,N_14506,N_12996);
and U17891 (N_17891,N_13923,N_12447);
or U17892 (N_17892,N_15702,N_14324);
or U17893 (N_17893,N_15304,N_12165);
nor U17894 (N_17894,N_13607,N_15549);
or U17895 (N_17895,N_13873,N_13945);
nand U17896 (N_17896,N_15084,N_15838);
nor U17897 (N_17897,N_14297,N_13847);
xor U17898 (N_17898,N_12253,N_14389);
nor U17899 (N_17899,N_13512,N_14644);
and U17900 (N_17900,N_12115,N_15402);
and U17901 (N_17901,N_13171,N_12532);
or U17902 (N_17902,N_14110,N_12163);
nand U17903 (N_17903,N_15363,N_12656);
or U17904 (N_17904,N_14134,N_14250);
or U17905 (N_17905,N_13493,N_12817);
nand U17906 (N_17906,N_13055,N_14828);
xor U17907 (N_17907,N_15017,N_12318);
nand U17908 (N_17908,N_14234,N_15469);
nand U17909 (N_17909,N_14732,N_13238);
and U17910 (N_17910,N_14079,N_14153);
and U17911 (N_17911,N_13547,N_14701);
nor U17912 (N_17912,N_13163,N_12869);
or U17913 (N_17913,N_15261,N_13142);
nor U17914 (N_17914,N_14434,N_14053);
and U17915 (N_17915,N_14638,N_14994);
and U17916 (N_17916,N_13639,N_13353);
xor U17917 (N_17917,N_12871,N_14165);
or U17918 (N_17918,N_15188,N_15614);
and U17919 (N_17919,N_12085,N_12816);
nor U17920 (N_17920,N_15157,N_13887);
nor U17921 (N_17921,N_13662,N_13395);
or U17922 (N_17922,N_13381,N_12893);
nand U17923 (N_17923,N_13710,N_13310);
and U17924 (N_17924,N_13336,N_15822);
nor U17925 (N_17925,N_15295,N_12101);
nand U17926 (N_17926,N_12381,N_12881);
and U17927 (N_17927,N_14683,N_14365);
nor U17928 (N_17928,N_13025,N_15009);
or U17929 (N_17929,N_12074,N_13460);
and U17930 (N_17930,N_15392,N_15563);
or U17931 (N_17931,N_14004,N_15807);
nand U17932 (N_17932,N_15362,N_12117);
nor U17933 (N_17933,N_12364,N_14693);
xor U17934 (N_17934,N_12755,N_15774);
nor U17935 (N_17935,N_15377,N_13703);
or U17936 (N_17936,N_15385,N_15069);
nand U17937 (N_17937,N_12887,N_13351);
nand U17938 (N_17938,N_14886,N_14901);
nand U17939 (N_17939,N_14688,N_12403);
xor U17940 (N_17940,N_13226,N_15784);
nand U17941 (N_17941,N_15055,N_12175);
nand U17942 (N_17942,N_12174,N_14343);
and U17943 (N_17943,N_15833,N_15555);
xor U17944 (N_17944,N_15444,N_14985);
and U17945 (N_17945,N_15024,N_12721);
xor U17946 (N_17946,N_12010,N_15644);
and U17947 (N_17947,N_15842,N_15813);
or U17948 (N_17948,N_14326,N_15154);
xor U17949 (N_17949,N_12018,N_13941);
and U17950 (N_17950,N_13043,N_12902);
nor U17951 (N_17951,N_13501,N_14243);
and U17952 (N_17952,N_13405,N_13304);
nand U17953 (N_17953,N_12139,N_14035);
xor U17954 (N_17954,N_15793,N_12133);
and U17955 (N_17955,N_13669,N_12058);
nand U17956 (N_17956,N_12262,N_12401);
and U17957 (N_17957,N_12353,N_14085);
or U17958 (N_17958,N_15322,N_14543);
and U17959 (N_17959,N_15847,N_15485);
nor U17960 (N_17960,N_15616,N_15867);
nand U17961 (N_17961,N_15526,N_12870);
nand U17962 (N_17962,N_13894,N_12611);
and U17963 (N_17963,N_14268,N_15329);
or U17964 (N_17964,N_12880,N_13698);
or U17965 (N_17965,N_13747,N_13186);
xor U17966 (N_17966,N_13549,N_14713);
or U17967 (N_17967,N_12113,N_14770);
and U17968 (N_17968,N_13463,N_12610);
xnor U17969 (N_17969,N_15921,N_13699);
xor U17970 (N_17970,N_14854,N_14514);
and U17971 (N_17971,N_14602,N_15302);
nor U17972 (N_17972,N_13212,N_12590);
or U17973 (N_17973,N_15970,N_15548);
or U17974 (N_17974,N_12571,N_12472);
or U17975 (N_17975,N_14950,N_15393);
nor U17976 (N_17976,N_15535,N_13308);
nor U17977 (N_17977,N_13005,N_15737);
nor U17978 (N_17978,N_13466,N_12137);
nor U17979 (N_17979,N_13283,N_13627);
nor U17980 (N_17980,N_12914,N_15398);
nand U17981 (N_17981,N_14068,N_13492);
and U17982 (N_17982,N_14475,N_12001);
nor U17983 (N_17983,N_13373,N_12463);
nor U17984 (N_17984,N_13957,N_13277);
nand U17985 (N_17985,N_15688,N_12014);
nor U17986 (N_17986,N_14919,N_14795);
nand U17987 (N_17987,N_13854,N_12567);
nand U17988 (N_17988,N_15075,N_13567);
nand U17989 (N_17989,N_15442,N_12559);
or U17990 (N_17990,N_13449,N_12306);
xnor U17991 (N_17991,N_12041,N_12227);
and U17992 (N_17992,N_13965,N_14131);
or U17993 (N_17993,N_13964,N_12254);
or U17994 (N_17994,N_12533,N_14123);
nor U17995 (N_17995,N_14724,N_14687);
nand U17996 (N_17996,N_15900,N_14288);
nand U17997 (N_17997,N_13119,N_15782);
nor U17998 (N_17998,N_13443,N_13799);
xor U17999 (N_17999,N_12951,N_14993);
nand U18000 (N_18000,N_15301,N_15970);
nand U18001 (N_18001,N_15707,N_14605);
nor U18002 (N_18002,N_15195,N_12928);
xor U18003 (N_18003,N_14514,N_14342);
and U18004 (N_18004,N_14480,N_14201);
xor U18005 (N_18005,N_14482,N_12228);
or U18006 (N_18006,N_12946,N_13928);
or U18007 (N_18007,N_14767,N_14280);
nor U18008 (N_18008,N_14675,N_12956);
nor U18009 (N_18009,N_15000,N_12183);
or U18010 (N_18010,N_13494,N_12247);
nand U18011 (N_18011,N_12168,N_15319);
and U18012 (N_18012,N_14566,N_12030);
nor U18013 (N_18013,N_12025,N_13217);
nand U18014 (N_18014,N_15896,N_12657);
or U18015 (N_18015,N_15519,N_13344);
nand U18016 (N_18016,N_14911,N_12448);
or U18017 (N_18017,N_15356,N_15701);
xor U18018 (N_18018,N_15214,N_15245);
nor U18019 (N_18019,N_14657,N_13473);
and U18020 (N_18020,N_14337,N_13329);
and U18021 (N_18021,N_12235,N_13629);
or U18022 (N_18022,N_13497,N_13412);
or U18023 (N_18023,N_14315,N_14779);
xor U18024 (N_18024,N_14864,N_14167);
nand U18025 (N_18025,N_13850,N_15825);
or U18026 (N_18026,N_12517,N_13243);
nor U18027 (N_18027,N_15545,N_13762);
nor U18028 (N_18028,N_14523,N_15665);
nand U18029 (N_18029,N_15242,N_15183);
and U18030 (N_18030,N_15449,N_13455);
nor U18031 (N_18031,N_12279,N_12670);
and U18032 (N_18032,N_12431,N_13033);
or U18033 (N_18033,N_12149,N_15741);
nor U18034 (N_18034,N_14187,N_15740);
nor U18035 (N_18035,N_13000,N_12445);
or U18036 (N_18036,N_14632,N_12362);
and U18037 (N_18037,N_14827,N_12630);
and U18038 (N_18038,N_14780,N_14023);
or U18039 (N_18039,N_14359,N_15890);
or U18040 (N_18040,N_12665,N_15990);
or U18041 (N_18041,N_13916,N_12308);
and U18042 (N_18042,N_13576,N_15195);
and U18043 (N_18043,N_13018,N_12900);
nor U18044 (N_18044,N_13945,N_13688);
nand U18045 (N_18045,N_15561,N_13596);
or U18046 (N_18046,N_14340,N_14654);
or U18047 (N_18047,N_14916,N_15711);
and U18048 (N_18048,N_14979,N_13211);
or U18049 (N_18049,N_14327,N_12487);
nor U18050 (N_18050,N_14576,N_12218);
and U18051 (N_18051,N_14554,N_13846);
nor U18052 (N_18052,N_13158,N_14201);
or U18053 (N_18053,N_14632,N_13921);
and U18054 (N_18054,N_15648,N_15108);
xor U18055 (N_18055,N_12360,N_15573);
or U18056 (N_18056,N_13992,N_12551);
and U18057 (N_18057,N_13865,N_12151);
nor U18058 (N_18058,N_12703,N_13616);
xnor U18059 (N_18059,N_15531,N_14810);
and U18060 (N_18060,N_12527,N_12437);
nor U18061 (N_18061,N_15475,N_13390);
nor U18062 (N_18062,N_12489,N_12296);
nand U18063 (N_18063,N_12118,N_15347);
nand U18064 (N_18064,N_13902,N_12155);
and U18065 (N_18065,N_13740,N_14195);
xor U18066 (N_18066,N_15627,N_14747);
nor U18067 (N_18067,N_13765,N_13588);
nor U18068 (N_18068,N_14661,N_14067);
xnor U18069 (N_18069,N_12617,N_14977);
nor U18070 (N_18070,N_15785,N_14049);
nand U18071 (N_18071,N_12092,N_14127);
and U18072 (N_18072,N_15206,N_13151);
or U18073 (N_18073,N_14317,N_15765);
nor U18074 (N_18074,N_12747,N_12109);
or U18075 (N_18075,N_14373,N_13735);
nor U18076 (N_18076,N_12509,N_13180);
and U18077 (N_18077,N_12754,N_13455);
nand U18078 (N_18078,N_13853,N_12016);
xnor U18079 (N_18079,N_14463,N_15836);
nand U18080 (N_18080,N_15193,N_13267);
nor U18081 (N_18081,N_12111,N_14140);
and U18082 (N_18082,N_13546,N_14611);
xnor U18083 (N_18083,N_15879,N_14315);
or U18084 (N_18084,N_15855,N_12623);
nor U18085 (N_18085,N_15703,N_12148);
xnor U18086 (N_18086,N_14808,N_12770);
and U18087 (N_18087,N_12736,N_14196);
nor U18088 (N_18088,N_15931,N_12498);
nand U18089 (N_18089,N_13429,N_14411);
nor U18090 (N_18090,N_14756,N_15811);
nand U18091 (N_18091,N_15760,N_13443);
and U18092 (N_18092,N_13299,N_15460);
and U18093 (N_18093,N_15294,N_12828);
nand U18094 (N_18094,N_13621,N_12529);
nand U18095 (N_18095,N_14138,N_13768);
nand U18096 (N_18096,N_12903,N_13639);
nor U18097 (N_18097,N_15069,N_12825);
xnor U18098 (N_18098,N_13489,N_14590);
xnor U18099 (N_18099,N_14813,N_13990);
or U18100 (N_18100,N_13977,N_15424);
nand U18101 (N_18101,N_13647,N_15839);
nor U18102 (N_18102,N_12883,N_13366);
nand U18103 (N_18103,N_13914,N_13617);
or U18104 (N_18104,N_14309,N_15975);
nor U18105 (N_18105,N_15228,N_12963);
nand U18106 (N_18106,N_15194,N_14528);
or U18107 (N_18107,N_13690,N_14764);
xnor U18108 (N_18108,N_13368,N_13741);
or U18109 (N_18109,N_12020,N_14603);
and U18110 (N_18110,N_12903,N_12220);
nand U18111 (N_18111,N_12822,N_12686);
and U18112 (N_18112,N_14157,N_13584);
and U18113 (N_18113,N_13025,N_13287);
and U18114 (N_18114,N_14802,N_14525);
nor U18115 (N_18115,N_13832,N_14982);
nor U18116 (N_18116,N_14344,N_12495);
or U18117 (N_18117,N_14294,N_15130);
or U18118 (N_18118,N_14103,N_12627);
and U18119 (N_18119,N_14854,N_13183);
or U18120 (N_18120,N_12918,N_12907);
or U18121 (N_18121,N_13217,N_14801);
xnor U18122 (N_18122,N_14514,N_12333);
or U18123 (N_18123,N_15470,N_12642);
nor U18124 (N_18124,N_15442,N_13487);
or U18125 (N_18125,N_14527,N_13108);
and U18126 (N_18126,N_12719,N_15294);
or U18127 (N_18127,N_12959,N_13769);
nand U18128 (N_18128,N_14165,N_13387);
nand U18129 (N_18129,N_12984,N_13957);
xnor U18130 (N_18130,N_13775,N_15226);
xor U18131 (N_18131,N_14137,N_13681);
or U18132 (N_18132,N_13896,N_15164);
and U18133 (N_18133,N_13343,N_12020);
nand U18134 (N_18134,N_14327,N_12146);
nor U18135 (N_18135,N_13250,N_12229);
xnor U18136 (N_18136,N_14020,N_15126);
nand U18137 (N_18137,N_14807,N_15591);
xor U18138 (N_18138,N_14395,N_13709);
and U18139 (N_18139,N_13597,N_12691);
nand U18140 (N_18140,N_14516,N_12643);
nand U18141 (N_18141,N_13673,N_13236);
or U18142 (N_18142,N_12782,N_12964);
or U18143 (N_18143,N_15850,N_13630);
or U18144 (N_18144,N_14659,N_13388);
nand U18145 (N_18145,N_12425,N_14225);
nor U18146 (N_18146,N_12347,N_14654);
nand U18147 (N_18147,N_14993,N_13761);
nand U18148 (N_18148,N_13049,N_12315);
or U18149 (N_18149,N_13712,N_15472);
nand U18150 (N_18150,N_13473,N_12590);
xor U18151 (N_18151,N_14855,N_12031);
nor U18152 (N_18152,N_13768,N_13113);
xnor U18153 (N_18153,N_14454,N_14986);
nor U18154 (N_18154,N_12060,N_13308);
or U18155 (N_18155,N_12634,N_15870);
nor U18156 (N_18156,N_12110,N_14016);
nor U18157 (N_18157,N_13045,N_13900);
xor U18158 (N_18158,N_12111,N_13229);
nor U18159 (N_18159,N_12127,N_13067);
or U18160 (N_18160,N_15585,N_13412);
or U18161 (N_18161,N_13185,N_12298);
and U18162 (N_18162,N_14021,N_14974);
and U18163 (N_18163,N_13277,N_13206);
nand U18164 (N_18164,N_15717,N_15450);
xnor U18165 (N_18165,N_12808,N_14519);
nor U18166 (N_18166,N_12038,N_13952);
and U18167 (N_18167,N_14446,N_15092);
nand U18168 (N_18168,N_12549,N_15588);
nand U18169 (N_18169,N_15873,N_14094);
nand U18170 (N_18170,N_15740,N_12402);
or U18171 (N_18171,N_14206,N_13734);
nor U18172 (N_18172,N_15463,N_13408);
and U18173 (N_18173,N_13921,N_14990);
nand U18174 (N_18174,N_15312,N_14224);
nor U18175 (N_18175,N_15632,N_13957);
xnor U18176 (N_18176,N_13954,N_14897);
and U18177 (N_18177,N_14116,N_12368);
nor U18178 (N_18178,N_13596,N_14355);
or U18179 (N_18179,N_13659,N_12340);
and U18180 (N_18180,N_12153,N_15051);
nand U18181 (N_18181,N_14535,N_14569);
and U18182 (N_18182,N_13215,N_12114);
and U18183 (N_18183,N_13016,N_13941);
nand U18184 (N_18184,N_12545,N_14442);
and U18185 (N_18185,N_15688,N_12186);
and U18186 (N_18186,N_13243,N_13964);
or U18187 (N_18187,N_13938,N_13033);
or U18188 (N_18188,N_12355,N_15847);
nand U18189 (N_18189,N_14289,N_14029);
or U18190 (N_18190,N_13646,N_13944);
and U18191 (N_18191,N_12586,N_15458);
and U18192 (N_18192,N_15835,N_14988);
or U18193 (N_18193,N_12766,N_12812);
or U18194 (N_18194,N_13842,N_15683);
or U18195 (N_18195,N_14928,N_15667);
or U18196 (N_18196,N_13109,N_12366);
xor U18197 (N_18197,N_12378,N_12221);
xnor U18198 (N_18198,N_14631,N_12307);
nand U18199 (N_18199,N_12519,N_15206);
nand U18200 (N_18200,N_13083,N_14501);
and U18201 (N_18201,N_12742,N_12947);
or U18202 (N_18202,N_12393,N_15903);
nand U18203 (N_18203,N_14907,N_13450);
nor U18204 (N_18204,N_15959,N_12139);
xor U18205 (N_18205,N_13453,N_12104);
or U18206 (N_18206,N_13366,N_13402);
or U18207 (N_18207,N_14958,N_14185);
or U18208 (N_18208,N_15013,N_15131);
or U18209 (N_18209,N_14179,N_12791);
or U18210 (N_18210,N_13460,N_13894);
and U18211 (N_18211,N_15115,N_12620);
nor U18212 (N_18212,N_15336,N_12959);
nor U18213 (N_18213,N_13832,N_12309);
and U18214 (N_18214,N_12360,N_15082);
and U18215 (N_18215,N_13634,N_13893);
nor U18216 (N_18216,N_12781,N_12260);
nand U18217 (N_18217,N_15895,N_13992);
nor U18218 (N_18218,N_12206,N_12910);
nor U18219 (N_18219,N_13950,N_15126);
and U18220 (N_18220,N_13159,N_14847);
nand U18221 (N_18221,N_12209,N_12472);
and U18222 (N_18222,N_14614,N_12765);
or U18223 (N_18223,N_12409,N_12149);
nand U18224 (N_18224,N_15770,N_15449);
nand U18225 (N_18225,N_12697,N_15232);
nor U18226 (N_18226,N_13160,N_14557);
xnor U18227 (N_18227,N_14277,N_12674);
nor U18228 (N_18228,N_12173,N_12582);
nand U18229 (N_18229,N_15917,N_13513);
xnor U18230 (N_18230,N_14585,N_15309);
nand U18231 (N_18231,N_12652,N_15355);
nor U18232 (N_18232,N_14294,N_15726);
and U18233 (N_18233,N_13726,N_13497);
or U18234 (N_18234,N_15892,N_14319);
or U18235 (N_18235,N_12824,N_15380);
nand U18236 (N_18236,N_13756,N_12401);
or U18237 (N_18237,N_14787,N_12830);
xnor U18238 (N_18238,N_15926,N_13823);
or U18239 (N_18239,N_15751,N_12019);
and U18240 (N_18240,N_14903,N_12203);
and U18241 (N_18241,N_13149,N_14443);
nand U18242 (N_18242,N_12443,N_15975);
and U18243 (N_18243,N_15489,N_14626);
xor U18244 (N_18244,N_15705,N_12245);
nor U18245 (N_18245,N_14404,N_12272);
nor U18246 (N_18246,N_13217,N_12556);
xor U18247 (N_18247,N_15792,N_14670);
nor U18248 (N_18248,N_14455,N_13010);
and U18249 (N_18249,N_12215,N_15783);
or U18250 (N_18250,N_14184,N_12438);
nand U18251 (N_18251,N_15528,N_13941);
nand U18252 (N_18252,N_15368,N_13470);
and U18253 (N_18253,N_12300,N_14021);
nand U18254 (N_18254,N_12681,N_13410);
or U18255 (N_18255,N_12460,N_14186);
or U18256 (N_18256,N_13437,N_12872);
xor U18257 (N_18257,N_13255,N_15273);
or U18258 (N_18258,N_12623,N_13323);
xnor U18259 (N_18259,N_14544,N_15953);
nor U18260 (N_18260,N_12302,N_15172);
nand U18261 (N_18261,N_14079,N_14726);
nand U18262 (N_18262,N_15751,N_14967);
nand U18263 (N_18263,N_12231,N_12302);
nand U18264 (N_18264,N_14214,N_15774);
nand U18265 (N_18265,N_13916,N_14553);
nor U18266 (N_18266,N_13837,N_15369);
nor U18267 (N_18267,N_12118,N_12781);
nand U18268 (N_18268,N_12807,N_13435);
nor U18269 (N_18269,N_12472,N_13008);
nor U18270 (N_18270,N_14552,N_12842);
or U18271 (N_18271,N_13749,N_14284);
xnor U18272 (N_18272,N_14197,N_12953);
or U18273 (N_18273,N_12672,N_15710);
or U18274 (N_18274,N_15481,N_15647);
nor U18275 (N_18275,N_13684,N_13600);
nor U18276 (N_18276,N_15122,N_15688);
or U18277 (N_18277,N_13117,N_15169);
nor U18278 (N_18278,N_12555,N_15178);
nor U18279 (N_18279,N_15290,N_13141);
nand U18280 (N_18280,N_14569,N_12744);
xnor U18281 (N_18281,N_13243,N_14343);
xor U18282 (N_18282,N_13543,N_13077);
nor U18283 (N_18283,N_14559,N_13490);
nor U18284 (N_18284,N_13007,N_12757);
nand U18285 (N_18285,N_13866,N_13517);
nand U18286 (N_18286,N_14487,N_12643);
and U18287 (N_18287,N_12253,N_12916);
nor U18288 (N_18288,N_12512,N_14779);
and U18289 (N_18289,N_15604,N_12720);
nor U18290 (N_18290,N_12164,N_13208);
nand U18291 (N_18291,N_15158,N_15925);
and U18292 (N_18292,N_12680,N_13019);
or U18293 (N_18293,N_15994,N_12960);
nor U18294 (N_18294,N_13816,N_13850);
nor U18295 (N_18295,N_15530,N_12891);
nor U18296 (N_18296,N_13227,N_13657);
nand U18297 (N_18297,N_13551,N_14165);
nor U18298 (N_18298,N_15274,N_12508);
nor U18299 (N_18299,N_12142,N_13099);
nor U18300 (N_18300,N_14197,N_13362);
nor U18301 (N_18301,N_12377,N_15787);
nand U18302 (N_18302,N_12275,N_15526);
nand U18303 (N_18303,N_13475,N_13861);
nand U18304 (N_18304,N_12240,N_12008);
or U18305 (N_18305,N_14501,N_14918);
nor U18306 (N_18306,N_12720,N_13587);
or U18307 (N_18307,N_12079,N_14096);
nand U18308 (N_18308,N_15202,N_13658);
and U18309 (N_18309,N_12926,N_14925);
and U18310 (N_18310,N_15261,N_13069);
or U18311 (N_18311,N_13091,N_12689);
and U18312 (N_18312,N_15054,N_13403);
xnor U18313 (N_18313,N_14774,N_15172);
xor U18314 (N_18314,N_15645,N_15179);
or U18315 (N_18315,N_12069,N_14933);
and U18316 (N_18316,N_15565,N_15679);
nand U18317 (N_18317,N_15006,N_13283);
or U18318 (N_18318,N_15171,N_15667);
or U18319 (N_18319,N_15287,N_15568);
or U18320 (N_18320,N_12935,N_14893);
and U18321 (N_18321,N_13467,N_13965);
nor U18322 (N_18322,N_15041,N_15907);
or U18323 (N_18323,N_12659,N_12417);
nand U18324 (N_18324,N_13427,N_15576);
and U18325 (N_18325,N_15940,N_15372);
nor U18326 (N_18326,N_12071,N_14211);
nor U18327 (N_18327,N_12957,N_14488);
or U18328 (N_18328,N_15787,N_14834);
nand U18329 (N_18329,N_14924,N_15199);
or U18330 (N_18330,N_15510,N_12232);
nor U18331 (N_18331,N_15898,N_12698);
nand U18332 (N_18332,N_12408,N_15763);
nand U18333 (N_18333,N_14949,N_12531);
nand U18334 (N_18334,N_13900,N_13366);
nand U18335 (N_18335,N_13387,N_15334);
nor U18336 (N_18336,N_12931,N_13343);
nand U18337 (N_18337,N_13933,N_13366);
and U18338 (N_18338,N_15645,N_13946);
and U18339 (N_18339,N_14285,N_15191);
nor U18340 (N_18340,N_15955,N_13145);
nor U18341 (N_18341,N_13199,N_13075);
nand U18342 (N_18342,N_14750,N_15277);
nand U18343 (N_18343,N_12721,N_14868);
nor U18344 (N_18344,N_12074,N_12818);
nor U18345 (N_18345,N_14806,N_12071);
and U18346 (N_18346,N_14588,N_13237);
nor U18347 (N_18347,N_12537,N_15974);
and U18348 (N_18348,N_15763,N_13821);
or U18349 (N_18349,N_13779,N_12625);
nor U18350 (N_18350,N_15461,N_13285);
or U18351 (N_18351,N_14215,N_15443);
nor U18352 (N_18352,N_12576,N_15838);
nand U18353 (N_18353,N_13854,N_13213);
nor U18354 (N_18354,N_15494,N_13014);
nand U18355 (N_18355,N_14215,N_15108);
xnor U18356 (N_18356,N_12626,N_15729);
nor U18357 (N_18357,N_12461,N_12815);
or U18358 (N_18358,N_15027,N_12340);
nand U18359 (N_18359,N_13540,N_13537);
or U18360 (N_18360,N_12523,N_12347);
and U18361 (N_18361,N_13311,N_15211);
xor U18362 (N_18362,N_13179,N_14669);
or U18363 (N_18363,N_13945,N_12141);
or U18364 (N_18364,N_14490,N_14717);
nor U18365 (N_18365,N_13646,N_13189);
or U18366 (N_18366,N_12512,N_15761);
nand U18367 (N_18367,N_13612,N_14193);
nor U18368 (N_18368,N_13500,N_13492);
and U18369 (N_18369,N_14142,N_13543);
or U18370 (N_18370,N_14312,N_14229);
and U18371 (N_18371,N_15147,N_15383);
and U18372 (N_18372,N_15627,N_12137);
nor U18373 (N_18373,N_15826,N_15478);
or U18374 (N_18374,N_12784,N_12343);
and U18375 (N_18375,N_14944,N_15700);
and U18376 (N_18376,N_14642,N_12610);
and U18377 (N_18377,N_15817,N_14608);
nor U18378 (N_18378,N_13172,N_15233);
xor U18379 (N_18379,N_12703,N_12442);
or U18380 (N_18380,N_15747,N_14886);
or U18381 (N_18381,N_15751,N_15690);
or U18382 (N_18382,N_13731,N_12647);
nor U18383 (N_18383,N_15187,N_13967);
nor U18384 (N_18384,N_12219,N_13552);
nor U18385 (N_18385,N_13045,N_13660);
nand U18386 (N_18386,N_12928,N_14862);
and U18387 (N_18387,N_13521,N_14111);
xor U18388 (N_18388,N_12482,N_14967);
nand U18389 (N_18389,N_12106,N_15634);
or U18390 (N_18390,N_13097,N_14055);
nand U18391 (N_18391,N_15362,N_15208);
xor U18392 (N_18392,N_12911,N_15087);
and U18393 (N_18393,N_13032,N_12739);
nand U18394 (N_18394,N_13458,N_13843);
nor U18395 (N_18395,N_12505,N_15503);
xnor U18396 (N_18396,N_13178,N_12468);
and U18397 (N_18397,N_14991,N_15318);
or U18398 (N_18398,N_14526,N_14177);
and U18399 (N_18399,N_14188,N_15921);
nand U18400 (N_18400,N_13080,N_12858);
nand U18401 (N_18401,N_15490,N_12351);
or U18402 (N_18402,N_12815,N_14896);
nor U18403 (N_18403,N_15811,N_13740);
nor U18404 (N_18404,N_12002,N_14879);
or U18405 (N_18405,N_15006,N_13020);
nand U18406 (N_18406,N_15187,N_13803);
xor U18407 (N_18407,N_15087,N_13601);
or U18408 (N_18408,N_15936,N_13011);
nand U18409 (N_18409,N_14349,N_12163);
and U18410 (N_18410,N_15389,N_14570);
or U18411 (N_18411,N_13092,N_15633);
or U18412 (N_18412,N_13432,N_14738);
nand U18413 (N_18413,N_15898,N_15703);
and U18414 (N_18414,N_12854,N_15109);
nand U18415 (N_18415,N_13895,N_14754);
nand U18416 (N_18416,N_15290,N_14288);
nor U18417 (N_18417,N_12981,N_15436);
nor U18418 (N_18418,N_15352,N_15409);
nor U18419 (N_18419,N_15749,N_14390);
nand U18420 (N_18420,N_12753,N_13066);
and U18421 (N_18421,N_15111,N_13417);
nor U18422 (N_18422,N_13278,N_13058);
xor U18423 (N_18423,N_14021,N_13772);
nand U18424 (N_18424,N_13578,N_13409);
nor U18425 (N_18425,N_15338,N_14802);
and U18426 (N_18426,N_15950,N_15483);
nor U18427 (N_18427,N_13506,N_12919);
nor U18428 (N_18428,N_13267,N_14413);
nand U18429 (N_18429,N_12038,N_13261);
and U18430 (N_18430,N_13802,N_15209);
nor U18431 (N_18431,N_13128,N_13015);
xor U18432 (N_18432,N_13994,N_12259);
or U18433 (N_18433,N_12816,N_14698);
and U18434 (N_18434,N_12706,N_14313);
nand U18435 (N_18435,N_12413,N_13887);
and U18436 (N_18436,N_12070,N_15103);
xor U18437 (N_18437,N_12456,N_15423);
and U18438 (N_18438,N_13940,N_12826);
nor U18439 (N_18439,N_13791,N_12596);
and U18440 (N_18440,N_14026,N_15378);
nand U18441 (N_18441,N_15876,N_13569);
nor U18442 (N_18442,N_15596,N_14845);
and U18443 (N_18443,N_15871,N_13617);
nand U18444 (N_18444,N_13438,N_15205);
xor U18445 (N_18445,N_14902,N_13654);
nor U18446 (N_18446,N_15553,N_14146);
nand U18447 (N_18447,N_12186,N_14860);
or U18448 (N_18448,N_12343,N_14595);
and U18449 (N_18449,N_14509,N_13260);
nor U18450 (N_18450,N_13007,N_14590);
nor U18451 (N_18451,N_13573,N_15676);
nor U18452 (N_18452,N_13384,N_15269);
or U18453 (N_18453,N_12269,N_13803);
xnor U18454 (N_18454,N_15681,N_13579);
xnor U18455 (N_18455,N_14183,N_15290);
and U18456 (N_18456,N_12321,N_15239);
nand U18457 (N_18457,N_13661,N_14124);
xnor U18458 (N_18458,N_15090,N_15032);
nand U18459 (N_18459,N_13226,N_15257);
or U18460 (N_18460,N_12068,N_14231);
and U18461 (N_18461,N_15133,N_13049);
nand U18462 (N_18462,N_12238,N_13989);
nor U18463 (N_18463,N_12181,N_12589);
or U18464 (N_18464,N_14990,N_12269);
nor U18465 (N_18465,N_12193,N_14607);
nor U18466 (N_18466,N_12893,N_14744);
nand U18467 (N_18467,N_14632,N_15127);
xnor U18468 (N_18468,N_13516,N_14756);
nand U18469 (N_18469,N_14120,N_15244);
and U18470 (N_18470,N_13110,N_15989);
nor U18471 (N_18471,N_12903,N_15271);
nor U18472 (N_18472,N_14989,N_15158);
nor U18473 (N_18473,N_14478,N_15112);
or U18474 (N_18474,N_12909,N_14961);
nor U18475 (N_18475,N_12512,N_13597);
or U18476 (N_18476,N_15581,N_14372);
nor U18477 (N_18477,N_14425,N_13980);
or U18478 (N_18478,N_13579,N_14999);
and U18479 (N_18479,N_12097,N_15453);
nand U18480 (N_18480,N_13296,N_12759);
or U18481 (N_18481,N_14064,N_15666);
or U18482 (N_18482,N_15654,N_13728);
nand U18483 (N_18483,N_14638,N_14817);
nand U18484 (N_18484,N_12059,N_15227);
nor U18485 (N_18485,N_13740,N_12001);
nor U18486 (N_18486,N_12909,N_14391);
and U18487 (N_18487,N_15832,N_15530);
and U18488 (N_18488,N_13186,N_14340);
nand U18489 (N_18489,N_14399,N_12347);
nand U18490 (N_18490,N_12213,N_14265);
or U18491 (N_18491,N_14258,N_12517);
and U18492 (N_18492,N_13156,N_12046);
and U18493 (N_18493,N_12131,N_15241);
nand U18494 (N_18494,N_13110,N_14703);
and U18495 (N_18495,N_13585,N_14156);
or U18496 (N_18496,N_13970,N_12816);
and U18497 (N_18497,N_15488,N_12532);
nor U18498 (N_18498,N_14901,N_14719);
and U18499 (N_18499,N_13380,N_13189);
nand U18500 (N_18500,N_15710,N_12211);
xnor U18501 (N_18501,N_13801,N_14076);
nand U18502 (N_18502,N_13027,N_12627);
xor U18503 (N_18503,N_13998,N_14697);
or U18504 (N_18504,N_14110,N_13924);
and U18505 (N_18505,N_14491,N_14714);
nand U18506 (N_18506,N_15400,N_12084);
or U18507 (N_18507,N_12802,N_13487);
and U18508 (N_18508,N_14055,N_15319);
and U18509 (N_18509,N_13368,N_12294);
nand U18510 (N_18510,N_14493,N_14693);
or U18511 (N_18511,N_13978,N_15205);
or U18512 (N_18512,N_15422,N_15013);
or U18513 (N_18513,N_13654,N_12520);
nor U18514 (N_18514,N_15383,N_15704);
or U18515 (N_18515,N_12937,N_13165);
or U18516 (N_18516,N_15058,N_12564);
and U18517 (N_18517,N_12067,N_15984);
xor U18518 (N_18518,N_12014,N_13530);
nor U18519 (N_18519,N_14996,N_14186);
and U18520 (N_18520,N_14108,N_14694);
xnor U18521 (N_18521,N_13647,N_13546);
xnor U18522 (N_18522,N_14904,N_12593);
nor U18523 (N_18523,N_12263,N_12626);
nand U18524 (N_18524,N_14624,N_12683);
and U18525 (N_18525,N_15967,N_13200);
nor U18526 (N_18526,N_15861,N_14589);
nor U18527 (N_18527,N_13547,N_12524);
nand U18528 (N_18528,N_13774,N_15689);
xnor U18529 (N_18529,N_14679,N_12110);
xnor U18530 (N_18530,N_15101,N_12604);
nor U18531 (N_18531,N_12540,N_15196);
or U18532 (N_18532,N_15181,N_15109);
nor U18533 (N_18533,N_14659,N_12935);
nand U18534 (N_18534,N_15099,N_14857);
nand U18535 (N_18535,N_15867,N_13323);
nor U18536 (N_18536,N_15014,N_15004);
xnor U18537 (N_18537,N_12447,N_15054);
and U18538 (N_18538,N_15905,N_14173);
or U18539 (N_18539,N_12868,N_15534);
or U18540 (N_18540,N_15217,N_12282);
or U18541 (N_18541,N_15881,N_12346);
nor U18542 (N_18542,N_14085,N_13666);
or U18543 (N_18543,N_12644,N_14124);
nand U18544 (N_18544,N_14989,N_15384);
or U18545 (N_18545,N_14431,N_14173);
nor U18546 (N_18546,N_14049,N_15556);
or U18547 (N_18547,N_12682,N_14038);
nor U18548 (N_18548,N_13109,N_12635);
nor U18549 (N_18549,N_13287,N_12780);
or U18550 (N_18550,N_15396,N_12513);
nor U18551 (N_18551,N_15368,N_15758);
and U18552 (N_18552,N_12080,N_15044);
xor U18553 (N_18553,N_12176,N_14132);
nand U18554 (N_18554,N_14623,N_15017);
or U18555 (N_18555,N_15775,N_14393);
nor U18556 (N_18556,N_14445,N_12018);
nor U18557 (N_18557,N_15080,N_12829);
or U18558 (N_18558,N_14952,N_13790);
nand U18559 (N_18559,N_12485,N_15809);
and U18560 (N_18560,N_13835,N_15656);
and U18561 (N_18561,N_12914,N_13512);
and U18562 (N_18562,N_15241,N_15220);
or U18563 (N_18563,N_15188,N_15154);
or U18564 (N_18564,N_14444,N_13082);
and U18565 (N_18565,N_13031,N_13163);
nand U18566 (N_18566,N_15035,N_14523);
nand U18567 (N_18567,N_15011,N_12008);
or U18568 (N_18568,N_12558,N_13136);
and U18569 (N_18569,N_12230,N_13444);
xnor U18570 (N_18570,N_12554,N_15272);
or U18571 (N_18571,N_12859,N_12680);
nand U18572 (N_18572,N_14831,N_15291);
and U18573 (N_18573,N_12741,N_15553);
nor U18574 (N_18574,N_12676,N_15764);
or U18575 (N_18575,N_13983,N_15330);
and U18576 (N_18576,N_14254,N_12538);
and U18577 (N_18577,N_14843,N_13428);
nor U18578 (N_18578,N_12477,N_15379);
or U18579 (N_18579,N_12913,N_13460);
or U18580 (N_18580,N_15498,N_14810);
nand U18581 (N_18581,N_14789,N_13334);
nor U18582 (N_18582,N_14155,N_14835);
nor U18583 (N_18583,N_13896,N_13818);
and U18584 (N_18584,N_15137,N_15254);
nand U18585 (N_18585,N_14586,N_15416);
or U18586 (N_18586,N_12049,N_14549);
nand U18587 (N_18587,N_12004,N_13792);
or U18588 (N_18588,N_15551,N_12627);
and U18589 (N_18589,N_12026,N_12409);
and U18590 (N_18590,N_13300,N_13526);
or U18591 (N_18591,N_14331,N_12800);
nand U18592 (N_18592,N_14736,N_13282);
and U18593 (N_18593,N_14798,N_15478);
nor U18594 (N_18594,N_12277,N_13083);
and U18595 (N_18595,N_15266,N_15117);
or U18596 (N_18596,N_12166,N_12882);
nor U18597 (N_18597,N_14591,N_12388);
nor U18598 (N_18598,N_14941,N_13679);
or U18599 (N_18599,N_12995,N_13910);
nor U18600 (N_18600,N_12918,N_13541);
and U18601 (N_18601,N_14413,N_14167);
nor U18602 (N_18602,N_12118,N_14562);
xor U18603 (N_18603,N_15256,N_12390);
or U18604 (N_18604,N_15227,N_14496);
nand U18605 (N_18605,N_12684,N_15991);
nand U18606 (N_18606,N_14387,N_14129);
or U18607 (N_18607,N_13921,N_15487);
xnor U18608 (N_18608,N_13829,N_14177);
nand U18609 (N_18609,N_15200,N_15720);
and U18610 (N_18610,N_15856,N_13561);
nand U18611 (N_18611,N_13222,N_13839);
nand U18612 (N_18612,N_13266,N_14212);
nand U18613 (N_18613,N_14460,N_12545);
xor U18614 (N_18614,N_12064,N_14187);
and U18615 (N_18615,N_12444,N_14788);
nand U18616 (N_18616,N_13295,N_13336);
or U18617 (N_18617,N_14331,N_12067);
or U18618 (N_18618,N_14333,N_13080);
xnor U18619 (N_18619,N_12758,N_12291);
and U18620 (N_18620,N_12551,N_15810);
or U18621 (N_18621,N_15662,N_14149);
nor U18622 (N_18622,N_14912,N_15503);
or U18623 (N_18623,N_12720,N_12370);
nand U18624 (N_18624,N_15064,N_14559);
and U18625 (N_18625,N_13286,N_13678);
xnor U18626 (N_18626,N_14214,N_14978);
xnor U18627 (N_18627,N_12050,N_15098);
nand U18628 (N_18628,N_14394,N_12122);
or U18629 (N_18629,N_12253,N_15314);
nor U18630 (N_18630,N_14666,N_12555);
xnor U18631 (N_18631,N_14667,N_15575);
nor U18632 (N_18632,N_14434,N_13461);
and U18633 (N_18633,N_15923,N_15406);
and U18634 (N_18634,N_13009,N_14942);
nand U18635 (N_18635,N_12088,N_15326);
and U18636 (N_18636,N_14627,N_13219);
and U18637 (N_18637,N_15295,N_13939);
and U18638 (N_18638,N_14253,N_13407);
or U18639 (N_18639,N_12967,N_12625);
xnor U18640 (N_18640,N_12898,N_12755);
xor U18641 (N_18641,N_12995,N_15028);
nand U18642 (N_18642,N_14349,N_15886);
xor U18643 (N_18643,N_15556,N_15440);
xor U18644 (N_18644,N_13497,N_14500);
nor U18645 (N_18645,N_13845,N_15154);
and U18646 (N_18646,N_15994,N_12337);
nand U18647 (N_18647,N_14917,N_12649);
nand U18648 (N_18648,N_12270,N_12016);
nor U18649 (N_18649,N_15762,N_14135);
nand U18650 (N_18650,N_13708,N_13322);
or U18651 (N_18651,N_15296,N_13824);
nor U18652 (N_18652,N_12458,N_14789);
or U18653 (N_18653,N_13134,N_13779);
nand U18654 (N_18654,N_14198,N_12076);
and U18655 (N_18655,N_13585,N_14972);
nand U18656 (N_18656,N_13985,N_14844);
or U18657 (N_18657,N_13385,N_14582);
nand U18658 (N_18658,N_15178,N_14796);
or U18659 (N_18659,N_12111,N_12015);
or U18660 (N_18660,N_12633,N_13477);
xnor U18661 (N_18661,N_14329,N_15191);
nor U18662 (N_18662,N_14571,N_13428);
nand U18663 (N_18663,N_13704,N_12387);
nand U18664 (N_18664,N_13998,N_13068);
xor U18665 (N_18665,N_14472,N_14795);
xor U18666 (N_18666,N_12792,N_14181);
and U18667 (N_18667,N_15726,N_13582);
or U18668 (N_18668,N_12539,N_13197);
xnor U18669 (N_18669,N_15373,N_12591);
nor U18670 (N_18670,N_15736,N_15336);
nor U18671 (N_18671,N_12505,N_12798);
nor U18672 (N_18672,N_12466,N_14776);
xor U18673 (N_18673,N_13430,N_15785);
nand U18674 (N_18674,N_15599,N_12625);
nor U18675 (N_18675,N_12274,N_12065);
nor U18676 (N_18676,N_15084,N_14453);
nand U18677 (N_18677,N_12342,N_14619);
nand U18678 (N_18678,N_14208,N_13955);
or U18679 (N_18679,N_13250,N_14146);
or U18680 (N_18680,N_12855,N_15705);
nor U18681 (N_18681,N_14456,N_12804);
and U18682 (N_18682,N_14324,N_12873);
and U18683 (N_18683,N_12565,N_13621);
or U18684 (N_18684,N_15346,N_13637);
or U18685 (N_18685,N_12972,N_12084);
nand U18686 (N_18686,N_13393,N_12827);
and U18687 (N_18687,N_13130,N_15378);
and U18688 (N_18688,N_13664,N_14939);
or U18689 (N_18689,N_12845,N_13527);
nor U18690 (N_18690,N_13628,N_12476);
nor U18691 (N_18691,N_14800,N_12384);
and U18692 (N_18692,N_13632,N_15148);
or U18693 (N_18693,N_13511,N_14622);
xnor U18694 (N_18694,N_12858,N_15474);
or U18695 (N_18695,N_14357,N_15481);
nand U18696 (N_18696,N_12602,N_13796);
nand U18697 (N_18697,N_13038,N_14227);
nand U18698 (N_18698,N_15458,N_12824);
and U18699 (N_18699,N_14000,N_13747);
and U18700 (N_18700,N_12024,N_13709);
nand U18701 (N_18701,N_12428,N_13020);
nand U18702 (N_18702,N_15629,N_15377);
nand U18703 (N_18703,N_15845,N_15844);
or U18704 (N_18704,N_15687,N_13949);
and U18705 (N_18705,N_13696,N_15192);
or U18706 (N_18706,N_15218,N_15677);
and U18707 (N_18707,N_12093,N_15161);
or U18708 (N_18708,N_12447,N_12117);
nand U18709 (N_18709,N_14512,N_14684);
nand U18710 (N_18710,N_15474,N_12961);
nor U18711 (N_18711,N_12074,N_14670);
and U18712 (N_18712,N_12983,N_13080);
or U18713 (N_18713,N_12678,N_12016);
and U18714 (N_18714,N_12329,N_12421);
nor U18715 (N_18715,N_15362,N_12548);
and U18716 (N_18716,N_15939,N_14584);
and U18717 (N_18717,N_14391,N_12620);
or U18718 (N_18718,N_13098,N_12747);
nand U18719 (N_18719,N_13626,N_14050);
nand U18720 (N_18720,N_14081,N_12605);
nor U18721 (N_18721,N_12831,N_12372);
or U18722 (N_18722,N_13695,N_15344);
nor U18723 (N_18723,N_15040,N_12971);
nor U18724 (N_18724,N_14187,N_14525);
or U18725 (N_18725,N_12313,N_12949);
and U18726 (N_18726,N_12017,N_15106);
or U18727 (N_18727,N_14929,N_13339);
or U18728 (N_18728,N_12676,N_13580);
and U18729 (N_18729,N_15548,N_14918);
nor U18730 (N_18730,N_14071,N_12304);
or U18731 (N_18731,N_15003,N_13847);
nand U18732 (N_18732,N_12712,N_15167);
and U18733 (N_18733,N_14267,N_13471);
nand U18734 (N_18734,N_14249,N_14693);
xnor U18735 (N_18735,N_15127,N_13037);
nand U18736 (N_18736,N_13089,N_15869);
nand U18737 (N_18737,N_14248,N_15694);
nand U18738 (N_18738,N_15674,N_14748);
nand U18739 (N_18739,N_15848,N_14632);
xor U18740 (N_18740,N_12688,N_13151);
nor U18741 (N_18741,N_12964,N_13133);
and U18742 (N_18742,N_13316,N_13756);
nor U18743 (N_18743,N_14670,N_13154);
or U18744 (N_18744,N_12408,N_13996);
nor U18745 (N_18745,N_12526,N_13733);
nor U18746 (N_18746,N_15006,N_15462);
and U18747 (N_18747,N_15449,N_15227);
nor U18748 (N_18748,N_12913,N_13445);
nand U18749 (N_18749,N_14802,N_14617);
nand U18750 (N_18750,N_12033,N_15047);
and U18751 (N_18751,N_12828,N_14022);
or U18752 (N_18752,N_13825,N_13194);
nor U18753 (N_18753,N_12363,N_14297);
and U18754 (N_18754,N_12858,N_12339);
nor U18755 (N_18755,N_14563,N_14791);
xor U18756 (N_18756,N_15029,N_12367);
and U18757 (N_18757,N_12532,N_15875);
or U18758 (N_18758,N_13357,N_13273);
or U18759 (N_18759,N_13089,N_14975);
or U18760 (N_18760,N_13212,N_12585);
or U18761 (N_18761,N_15422,N_12343);
nand U18762 (N_18762,N_15208,N_14761);
nand U18763 (N_18763,N_13584,N_13779);
and U18764 (N_18764,N_12326,N_12941);
and U18765 (N_18765,N_14092,N_14001);
nand U18766 (N_18766,N_13294,N_13817);
or U18767 (N_18767,N_14736,N_13181);
xor U18768 (N_18768,N_14663,N_15163);
or U18769 (N_18769,N_13647,N_15178);
or U18770 (N_18770,N_14275,N_14528);
xor U18771 (N_18771,N_15088,N_15753);
xor U18772 (N_18772,N_12689,N_14213);
and U18773 (N_18773,N_15862,N_13123);
nor U18774 (N_18774,N_13828,N_15705);
nand U18775 (N_18775,N_12745,N_12764);
and U18776 (N_18776,N_12646,N_14442);
xnor U18777 (N_18777,N_12451,N_12892);
or U18778 (N_18778,N_14822,N_14612);
nand U18779 (N_18779,N_13155,N_13667);
nor U18780 (N_18780,N_13924,N_14469);
nand U18781 (N_18781,N_14247,N_14940);
nand U18782 (N_18782,N_14289,N_15501);
and U18783 (N_18783,N_12116,N_13744);
or U18784 (N_18784,N_15695,N_12429);
nor U18785 (N_18785,N_12107,N_12712);
or U18786 (N_18786,N_12235,N_15609);
nand U18787 (N_18787,N_15339,N_12784);
or U18788 (N_18788,N_12308,N_13870);
nand U18789 (N_18789,N_13305,N_14127);
or U18790 (N_18790,N_12701,N_12153);
or U18791 (N_18791,N_15381,N_14967);
or U18792 (N_18792,N_15533,N_12636);
or U18793 (N_18793,N_14542,N_12650);
xor U18794 (N_18794,N_12795,N_13546);
and U18795 (N_18795,N_14115,N_13920);
nand U18796 (N_18796,N_15551,N_12792);
and U18797 (N_18797,N_14861,N_12068);
or U18798 (N_18798,N_13385,N_15201);
nand U18799 (N_18799,N_12988,N_12696);
and U18800 (N_18800,N_14955,N_14047);
nor U18801 (N_18801,N_15210,N_12583);
nor U18802 (N_18802,N_13837,N_14199);
nand U18803 (N_18803,N_15946,N_13461);
nand U18804 (N_18804,N_15889,N_13206);
and U18805 (N_18805,N_12165,N_13456);
and U18806 (N_18806,N_15604,N_14142);
and U18807 (N_18807,N_12536,N_14562);
nand U18808 (N_18808,N_13379,N_13100);
nor U18809 (N_18809,N_13620,N_12416);
nor U18810 (N_18810,N_15408,N_12109);
or U18811 (N_18811,N_14202,N_12309);
and U18812 (N_18812,N_13057,N_12296);
or U18813 (N_18813,N_13991,N_12054);
or U18814 (N_18814,N_14124,N_14801);
and U18815 (N_18815,N_14245,N_13451);
or U18816 (N_18816,N_13145,N_14471);
nand U18817 (N_18817,N_13144,N_13883);
or U18818 (N_18818,N_12461,N_15780);
and U18819 (N_18819,N_13835,N_15082);
and U18820 (N_18820,N_15563,N_15269);
xnor U18821 (N_18821,N_15199,N_14540);
nor U18822 (N_18822,N_13510,N_15821);
nor U18823 (N_18823,N_14412,N_13526);
nand U18824 (N_18824,N_15344,N_12822);
nand U18825 (N_18825,N_14216,N_15983);
nor U18826 (N_18826,N_14492,N_15717);
nand U18827 (N_18827,N_12824,N_15360);
and U18828 (N_18828,N_14068,N_15530);
nor U18829 (N_18829,N_14710,N_14564);
and U18830 (N_18830,N_13398,N_15470);
or U18831 (N_18831,N_12268,N_14121);
or U18832 (N_18832,N_13633,N_12447);
and U18833 (N_18833,N_14720,N_14687);
nand U18834 (N_18834,N_15248,N_15093);
and U18835 (N_18835,N_14777,N_15124);
and U18836 (N_18836,N_15054,N_12535);
nand U18837 (N_18837,N_13723,N_13928);
and U18838 (N_18838,N_14916,N_14401);
or U18839 (N_18839,N_14196,N_12142);
and U18840 (N_18840,N_14284,N_14606);
nand U18841 (N_18841,N_14189,N_13565);
nand U18842 (N_18842,N_12219,N_13948);
nand U18843 (N_18843,N_15167,N_12488);
nand U18844 (N_18844,N_14840,N_15255);
and U18845 (N_18845,N_15382,N_14281);
nand U18846 (N_18846,N_12969,N_13426);
nand U18847 (N_18847,N_15451,N_12685);
nand U18848 (N_18848,N_12378,N_13044);
or U18849 (N_18849,N_14939,N_13952);
nor U18850 (N_18850,N_12564,N_13897);
and U18851 (N_18851,N_15874,N_14612);
or U18852 (N_18852,N_14312,N_14032);
nand U18853 (N_18853,N_14413,N_14268);
xor U18854 (N_18854,N_15872,N_15874);
nand U18855 (N_18855,N_14382,N_15318);
and U18856 (N_18856,N_12731,N_12897);
nand U18857 (N_18857,N_13013,N_12228);
nor U18858 (N_18858,N_15121,N_14911);
nand U18859 (N_18859,N_13591,N_13502);
nor U18860 (N_18860,N_13889,N_14778);
and U18861 (N_18861,N_14562,N_12469);
xnor U18862 (N_18862,N_12318,N_14434);
nor U18863 (N_18863,N_13321,N_14275);
nand U18864 (N_18864,N_13888,N_14644);
xnor U18865 (N_18865,N_13086,N_13863);
nor U18866 (N_18866,N_12818,N_12533);
nand U18867 (N_18867,N_14285,N_13742);
nor U18868 (N_18868,N_13231,N_12613);
and U18869 (N_18869,N_12142,N_14107);
nor U18870 (N_18870,N_14172,N_14620);
and U18871 (N_18871,N_14876,N_12538);
nor U18872 (N_18872,N_13475,N_14696);
nor U18873 (N_18873,N_15248,N_13316);
or U18874 (N_18874,N_13955,N_12753);
xor U18875 (N_18875,N_15777,N_12964);
and U18876 (N_18876,N_13146,N_13842);
xor U18877 (N_18877,N_15188,N_15993);
or U18878 (N_18878,N_14084,N_14633);
nor U18879 (N_18879,N_14211,N_15989);
nand U18880 (N_18880,N_14493,N_14749);
nand U18881 (N_18881,N_15565,N_13225);
and U18882 (N_18882,N_14644,N_12448);
or U18883 (N_18883,N_15582,N_15642);
xor U18884 (N_18884,N_13089,N_14694);
and U18885 (N_18885,N_14835,N_14218);
xor U18886 (N_18886,N_14029,N_12605);
or U18887 (N_18887,N_15813,N_14026);
nor U18888 (N_18888,N_14437,N_12823);
and U18889 (N_18889,N_15502,N_12827);
or U18890 (N_18890,N_15497,N_15318);
and U18891 (N_18891,N_15586,N_15049);
and U18892 (N_18892,N_14132,N_15763);
nor U18893 (N_18893,N_14988,N_14164);
and U18894 (N_18894,N_15169,N_15532);
or U18895 (N_18895,N_15624,N_15385);
nor U18896 (N_18896,N_14042,N_14313);
or U18897 (N_18897,N_12350,N_14437);
and U18898 (N_18898,N_12043,N_15832);
nor U18899 (N_18899,N_12028,N_13438);
xnor U18900 (N_18900,N_15548,N_14996);
nor U18901 (N_18901,N_14359,N_12637);
or U18902 (N_18902,N_13250,N_13361);
nand U18903 (N_18903,N_15386,N_14660);
nand U18904 (N_18904,N_13836,N_15059);
nor U18905 (N_18905,N_13584,N_12681);
xor U18906 (N_18906,N_15801,N_13861);
nand U18907 (N_18907,N_13309,N_15379);
nor U18908 (N_18908,N_13055,N_13364);
and U18909 (N_18909,N_14912,N_12676);
or U18910 (N_18910,N_15551,N_13744);
nor U18911 (N_18911,N_13009,N_13557);
or U18912 (N_18912,N_12917,N_14016);
or U18913 (N_18913,N_13712,N_13762);
nand U18914 (N_18914,N_12575,N_12417);
nor U18915 (N_18915,N_14676,N_15591);
nand U18916 (N_18916,N_15472,N_15513);
and U18917 (N_18917,N_12460,N_13378);
or U18918 (N_18918,N_14019,N_14447);
nand U18919 (N_18919,N_14758,N_13528);
nor U18920 (N_18920,N_14626,N_12682);
and U18921 (N_18921,N_12570,N_15842);
or U18922 (N_18922,N_13796,N_12277);
nor U18923 (N_18923,N_14223,N_13764);
and U18924 (N_18924,N_15693,N_14871);
nand U18925 (N_18925,N_12150,N_15192);
nand U18926 (N_18926,N_13180,N_12403);
or U18927 (N_18927,N_15500,N_13843);
or U18928 (N_18928,N_13210,N_15302);
or U18929 (N_18929,N_12898,N_14077);
nor U18930 (N_18930,N_13331,N_13951);
and U18931 (N_18931,N_14023,N_13710);
or U18932 (N_18932,N_12169,N_15930);
and U18933 (N_18933,N_12910,N_12539);
or U18934 (N_18934,N_13060,N_15310);
xnor U18935 (N_18935,N_12341,N_15185);
xor U18936 (N_18936,N_15419,N_14916);
nor U18937 (N_18937,N_14758,N_12412);
nand U18938 (N_18938,N_12707,N_13684);
or U18939 (N_18939,N_12535,N_13360);
or U18940 (N_18940,N_15023,N_12870);
and U18941 (N_18941,N_12870,N_12558);
nor U18942 (N_18942,N_15500,N_13536);
or U18943 (N_18943,N_12352,N_15110);
and U18944 (N_18944,N_13160,N_13939);
nand U18945 (N_18945,N_14378,N_15914);
and U18946 (N_18946,N_15750,N_13728);
nor U18947 (N_18947,N_15694,N_14619);
nand U18948 (N_18948,N_15026,N_12010);
or U18949 (N_18949,N_15297,N_13618);
nor U18950 (N_18950,N_13346,N_12991);
and U18951 (N_18951,N_15332,N_14570);
nand U18952 (N_18952,N_15839,N_15109);
or U18953 (N_18953,N_12948,N_14484);
nand U18954 (N_18954,N_13306,N_12075);
nor U18955 (N_18955,N_12729,N_14054);
or U18956 (N_18956,N_13036,N_13350);
and U18957 (N_18957,N_15525,N_12926);
nand U18958 (N_18958,N_15126,N_14195);
and U18959 (N_18959,N_15902,N_13021);
or U18960 (N_18960,N_12060,N_14807);
and U18961 (N_18961,N_15640,N_15841);
and U18962 (N_18962,N_15439,N_14023);
or U18963 (N_18963,N_14914,N_14843);
nand U18964 (N_18964,N_14251,N_15711);
nand U18965 (N_18965,N_13574,N_13852);
nand U18966 (N_18966,N_14387,N_12463);
xnor U18967 (N_18967,N_15978,N_14344);
xor U18968 (N_18968,N_15367,N_15737);
or U18969 (N_18969,N_15437,N_13421);
or U18970 (N_18970,N_14793,N_14857);
or U18971 (N_18971,N_12536,N_15803);
and U18972 (N_18972,N_12430,N_14162);
nor U18973 (N_18973,N_13482,N_13912);
and U18974 (N_18974,N_15794,N_15427);
xnor U18975 (N_18975,N_15071,N_14064);
and U18976 (N_18976,N_14180,N_12879);
and U18977 (N_18977,N_14627,N_13480);
and U18978 (N_18978,N_12220,N_12912);
or U18979 (N_18979,N_12067,N_12372);
nor U18980 (N_18980,N_14225,N_15285);
or U18981 (N_18981,N_12689,N_12861);
and U18982 (N_18982,N_15399,N_14634);
and U18983 (N_18983,N_14729,N_14681);
and U18984 (N_18984,N_14495,N_15735);
nor U18985 (N_18985,N_13863,N_15335);
nor U18986 (N_18986,N_15095,N_14209);
xnor U18987 (N_18987,N_15578,N_15577);
and U18988 (N_18988,N_13802,N_13859);
nand U18989 (N_18989,N_14467,N_14028);
nor U18990 (N_18990,N_15428,N_15436);
and U18991 (N_18991,N_15200,N_12044);
nand U18992 (N_18992,N_15768,N_14276);
and U18993 (N_18993,N_12381,N_15574);
nor U18994 (N_18994,N_14304,N_14052);
nor U18995 (N_18995,N_14609,N_13995);
or U18996 (N_18996,N_12399,N_15764);
nor U18997 (N_18997,N_13873,N_12461);
and U18998 (N_18998,N_15429,N_12384);
and U18999 (N_18999,N_15944,N_15379);
or U19000 (N_19000,N_14353,N_13364);
nand U19001 (N_19001,N_15152,N_13304);
or U19002 (N_19002,N_14448,N_12306);
xor U19003 (N_19003,N_13129,N_15678);
xor U19004 (N_19004,N_12792,N_14918);
nand U19005 (N_19005,N_13697,N_14422);
nand U19006 (N_19006,N_12410,N_13773);
nor U19007 (N_19007,N_12146,N_15577);
nand U19008 (N_19008,N_12935,N_14723);
or U19009 (N_19009,N_12279,N_13248);
nor U19010 (N_19010,N_13611,N_15500);
or U19011 (N_19011,N_15741,N_15259);
and U19012 (N_19012,N_15816,N_12338);
or U19013 (N_19013,N_13660,N_15271);
xnor U19014 (N_19014,N_15634,N_14557);
and U19015 (N_19015,N_14770,N_15978);
or U19016 (N_19016,N_14398,N_13728);
nand U19017 (N_19017,N_13255,N_13316);
and U19018 (N_19018,N_13909,N_12635);
or U19019 (N_19019,N_15814,N_12916);
nor U19020 (N_19020,N_12831,N_15651);
and U19021 (N_19021,N_12035,N_13244);
and U19022 (N_19022,N_14634,N_13513);
nand U19023 (N_19023,N_13973,N_12680);
xor U19024 (N_19024,N_13613,N_15281);
or U19025 (N_19025,N_12511,N_15165);
nand U19026 (N_19026,N_13779,N_13563);
nand U19027 (N_19027,N_12434,N_13195);
nor U19028 (N_19028,N_14433,N_13128);
and U19029 (N_19029,N_15787,N_15902);
or U19030 (N_19030,N_12450,N_15531);
nand U19031 (N_19031,N_12919,N_13229);
nand U19032 (N_19032,N_15695,N_12181);
nor U19033 (N_19033,N_14955,N_13222);
nor U19034 (N_19034,N_15272,N_14780);
and U19035 (N_19035,N_14724,N_15310);
and U19036 (N_19036,N_13605,N_15715);
nand U19037 (N_19037,N_13438,N_14955);
or U19038 (N_19038,N_15836,N_13363);
or U19039 (N_19039,N_13825,N_12401);
nand U19040 (N_19040,N_12780,N_14648);
and U19041 (N_19041,N_13395,N_14282);
and U19042 (N_19042,N_13160,N_15090);
nand U19043 (N_19043,N_14857,N_12280);
and U19044 (N_19044,N_13762,N_12322);
nor U19045 (N_19045,N_13901,N_12543);
nand U19046 (N_19046,N_14326,N_13677);
or U19047 (N_19047,N_13271,N_12411);
and U19048 (N_19048,N_12231,N_14972);
or U19049 (N_19049,N_13291,N_15666);
xor U19050 (N_19050,N_15954,N_15307);
nand U19051 (N_19051,N_12282,N_12229);
and U19052 (N_19052,N_12520,N_14517);
or U19053 (N_19053,N_13935,N_13774);
and U19054 (N_19054,N_14561,N_12762);
or U19055 (N_19055,N_13745,N_15536);
nor U19056 (N_19056,N_13996,N_12493);
or U19057 (N_19057,N_12849,N_12037);
nand U19058 (N_19058,N_15849,N_15449);
xnor U19059 (N_19059,N_15369,N_14542);
and U19060 (N_19060,N_15370,N_12257);
nand U19061 (N_19061,N_13781,N_12894);
nor U19062 (N_19062,N_15953,N_13536);
or U19063 (N_19063,N_12278,N_12647);
and U19064 (N_19064,N_14075,N_13966);
nor U19065 (N_19065,N_15147,N_12662);
nand U19066 (N_19066,N_15502,N_13853);
nand U19067 (N_19067,N_15334,N_13463);
nor U19068 (N_19068,N_13691,N_14370);
or U19069 (N_19069,N_12600,N_15636);
and U19070 (N_19070,N_15583,N_13272);
nor U19071 (N_19071,N_15497,N_15688);
xnor U19072 (N_19072,N_13226,N_13231);
and U19073 (N_19073,N_15365,N_15155);
and U19074 (N_19074,N_13852,N_15536);
nor U19075 (N_19075,N_15270,N_14481);
or U19076 (N_19076,N_14029,N_12436);
nor U19077 (N_19077,N_13611,N_13015);
or U19078 (N_19078,N_15980,N_13856);
nand U19079 (N_19079,N_15562,N_14560);
and U19080 (N_19080,N_13846,N_15047);
nand U19081 (N_19081,N_14398,N_12019);
nor U19082 (N_19082,N_12658,N_15362);
or U19083 (N_19083,N_12348,N_12693);
and U19084 (N_19084,N_14751,N_15630);
and U19085 (N_19085,N_13504,N_15244);
nand U19086 (N_19086,N_12011,N_12295);
and U19087 (N_19087,N_14015,N_15234);
or U19088 (N_19088,N_14404,N_12159);
nand U19089 (N_19089,N_15273,N_15292);
nor U19090 (N_19090,N_12558,N_13300);
nor U19091 (N_19091,N_13021,N_15610);
or U19092 (N_19092,N_12520,N_12977);
nor U19093 (N_19093,N_15687,N_14881);
nor U19094 (N_19094,N_15421,N_13486);
nor U19095 (N_19095,N_14502,N_13851);
nand U19096 (N_19096,N_14803,N_12058);
nor U19097 (N_19097,N_13740,N_15995);
nor U19098 (N_19098,N_15215,N_12979);
nand U19099 (N_19099,N_15643,N_14128);
nor U19100 (N_19100,N_12327,N_15076);
nand U19101 (N_19101,N_12404,N_14424);
and U19102 (N_19102,N_14645,N_13291);
nand U19103 (N_19103,N_12129,N_15133);
or U19104 (N_19104,N_15006,N_13016);
nor U19105 (N_19105,N_15639,N_12730);
nand U19106 (N_19106,N_15595,N_13485);
and U19107 (N_19107,N_14423,N_14387);
and U19108 (N_19108,N_14598,N_13361);
and U19109 (N_19109,N_14362,N_12471);
nor U19110 (N_19110,N_15354,N_12399);
nor U19111 (N_19111,N_12954,N_15349);
nand U19112 (N_19112,N_12780,N_12287);
nand U19113 (N_19113,N_13940,N_14135);
nor U19114 (N_19114,N_14870,N_13958);
xnor U19115 (N_19115,N_14705,N_12077);
or U19116 (N_19116,N_13412,N_13801);
nor U19117 (N_19117,N_13983,N_14960);
xor U19118 (N_19118,N_12041,N_14178);
nor U19119 (N_19119,N_14531,N_15098);
nor U19120 (N_19120,N_15455,N_14308);
nand U19121 (N_19121,N_15338,N_12580);
nand U19122 (N_19122,N_12393,N_12398);
and U19123 (N_19123,N_15155,N_15904);
or U19124 (N_19124,N_15952,N_12788);
nor U19125 (N_19125,N_14208,N_12185);
and U19126 (N_19126,N_13894,N_14009);
nand U19127 (N_19127,N_14324,N_13648);
nand U19128 (N_19128,N_12880,N_15292);
xor U19129 (N_19129,N_14873,N_13022);
nor U19130 (N_19130,N_15605,N_12123);
nor U19131 (N_19131,N_13449,N_13033);
xor U19132 (N_19132,N_15595,N_15760);
nand U19133 (N_19133,N_14339,N_14288);
nor U19134 (N_19134,N_13833,N_13816);
nand U19135 (N_19135,N_15235,N_14297);
nand U19136 (N_19136,N_13732,N_15984);
nor U19137 (N_19137,N_14278,N_15846);
or U19138 (N_19138,N_12808,N_13058);
nor U19139 (N_19139,N_12792,N_14133);
and U19140 (N_19140,N_13996,N_12870);
nor U19141 (N_19141,N_14007,N_15828);
and U19142 (N_19142,N_15076,N_12864);
xnor U19143 (N_19143,N_14116,N_12903);
nor U19144 (N_19144,N_14912,N_14586);
nand U19145 (N_19145,N_15094,N_13697);
xor U19146 (N_19146,N_15396,N_15510);
or U19147 (N_19147,N_13238,N_15945);
nand U19148 (N_19148,N_14285,N_15845);
or U19149 (N_19149,N_14002,N_15955);
or U19150 (N_19150,N_14696,N_13883);
or U19151 (N_19151,N_13806,N_15072);
nand U19152 (N_19152,N_14457,N_14608);
nor U19153 (N_19153,N_14942,N_15613);
or U19154 (N_19154,N_13353,N_13175);
nor U19155 (N_19155,N_14988,N_13145);
and U19156 (N_19156,N_12958,N_15417);
or U19157 (N_19157,N_12778,N_15860);
nor U19158 (N_19158,N_13827,N_12875);
nor U19159 (N_19159,N_13741,N_14333);
nor U19160 (N_19160,N_15169,N_14759);
nand U19161 (N_19161,N_14439,N_14186);
nor U19162 (N_19162,N_12821,N_12482);
nor U19163 (N_19163,N_14160,N_13477);
or U19164 (N_19164,N_14483,N_15740);
nand U19165 (N_19165,N_14519,N_12286);
or U19166 (N_19166,N_12013,N_13072);
nand U19167 (N_19167,N_12255,N_15121);
nand U19168 (N_19168,N_15311,N_15103);
nand U19169 (N_19169,N_12888,N_15711);
xor U19170 (N_19170,N_14011,N_13557);
nor U19171 (N_19171,N_14209,N_14964);
and U19172 (N_19172,N_12463,N_14588);
and U19173 (N_19173,N_12573,N_12622);
and U19174 (N_19174,N_13936,N_14680);
xor U19175 (N_19175,N_13312,N_12608);
nor U19176 (N_19176,N_14403,N_15447);
or U19177 (N_19177,N_15445,N_12360);
or U19178 (N_19178,N_15134,N_15888);
or U19179 (N_19179,N_15935,N_13997);
and U19180 (N_19180,N_15972,N_13799);
or U19181 (N_19181,N_14985,N_14362);
xor U19182 (N_19182,N_12661,N_12821);
xnor U19183 (N_19183,N_13124,N_13078);
and U19184 (N_19184,N_12766,N_12947);
nor U19185 (N_19185,N_15826,N_14237);
xor U19186 (N_19186,N_15460,N_12682);
nor U19187 (N_19187,N_15450,N_15401);
nor U19188 (N_19188,N_14776,N_14023);
nand U19189 (N_19189,N_12423,N_13551);
nand U19190 (N_19190,N_14499,N_13261);
nand U19191 (N_19191,N_13159,N_15941);
nor U19192 (N_19192,N_15461,N_15566);
xnor U19193 (N_19193,N_15303,N_14311);
nand U19194 (N_19194,N_12744,N_12894);
nand U19195 (N_19195,N_15644,N_13200);
or U19196 (N_19196,N_15046,N_12747);
nand U19197 (N_19197,N_13742,N_13943);
and U19198 (N_19198,N_13424,N_13415);
nor U19199 (N_19199,N_13789,N_14828);
nor U19200 (N_19200,N_14571,N_14185);
nor U19201 (N_19201,N_14813,N_13209);
nand U19202 (N_19202,N_15326,N_14491);
and U19203 (N_19203,N_12478,N_13851);
nor U19204 (N_19204,N_12383,N_14587);
and U19205 (N_19205,N_12316,N_14135);
nor U19206 (N_19206,N_12075,N_12216);
nand U19207 (N_19207,N_12977,N_15627);
nor U19208 (N_19208,N_15479,N_12942);
and U19209 (N_19209,N_13001,N_12462);
nand U19210 (N_19210,N_12289,N_13206);
and U19211 (N_19211,N_15639,N_12800);
nor U19212 (N_19212,N_15602,N_14293);
nand U19213 (N_19213,N_13367,N_15606);
or U19214 (N_19214,N_15604,N_13903);
or U19215 (N_19215,N_12572,N_12014);
nand U19216 (N_19216,N_12666,N_14113);
nand U19217 (N_19217,N_12556,N_13771);
or U19218 (N_19218,N_12537,N_13411);
nor U19219 (N_19219,N_13552,N_14977);
nand U19220 (N_19220,N_13402,N_14772);
and U19221 (N_19221,N_12572,N_12115);
and U19222 (N_19222,N_14982,N_14199);
nor U19223 (N_19223,N_12203,N_12666);
or U19224 (N_19224,N_13851,N_12544);
or U19225 (N_19225,N_12168,N_12467);
and U19226 (N_19226,N_15335,N_14434);
xnor U19227 (N_19227,N_14186,N_14862);
and U19228 (N_19228,N_13572,N_12410);
nor U19229 (N_19229,N_12320,N_12134);
xor U19230 (N_19230,N_13019,N_13027);
or U19231 (N_19231,N_13361,N_12426);
nor U19232 (N_19232,N_14299,N_14327);
xnor U19233 (N_19233,N_13651,N_15573);
xor U19234 (N_19234,N_12335,N_15084);
nor U19235 (N_19235,N_12257,N_15316);
nand U19236 (N_19236,N_14281,N_13088);
and U19237 (N_19237,N_13051,N_13424);
nor U19238 (N_19238,N_12640,N_14687);
or U19239 (N_19239,N_15233,N_14629);
nand U19240 (N_19240,N_15304,N_14424);
nor U19241 (N_19241,N_14097,N_12354);
nor U19242 (N_19242,N_13910,N_14084);
xor U19243 (N_19243,N_12081,N_15658);
and U19244 (N_19244,N_15441,N_14220);
and U19245 (N_19245,N_13160,N_15150);
nor U19246 (N_19246,N_15844,N_13267);
nand U19247 (N_19247,N_13054,N_14909);
and U19248 (N_19248,N_15708,N_12144);
and U19249 (N_19249,N_15817,N_14284);
xor U19250 (N_19250,N_13162,N_15369);
nor U19251 (N_19251,N_15093,N_14719);
and U19252 (N_19252,N_15896,N_13000);
or U19253 (N_19253,N_13312,N_15650);
or U19254 (N_19254,N_13700,N_12949);
xnor U19255 (N_19255,N_15888,N_12165);
or U19256 (N_19256,N_13233,N_13218);
and U19257 (N_19257,N_13590,N_13088);
and U19258 (N_19258,N_14060,N_15550);
and U19259 (N_19259,N_14950,N_12973);
nand U19260 (N_19260,N_14409,N_13579);
nand U19261 (N_19261,N_12614,N_15070);
nand U19262 (N_19262,N_15504,N_15540);
nor U19263 (N_19263,N_14990,N_14908);
nor U19264 (N_19264,N_15857,N_15930);
and U19265 (N_19265,N_14547,N_13120);
nand U19266 (N_19266,N_12186,N_12924);
nor U19267 (N_19267,N_13504,N_15616);
nor U19268 (N_19268,N_14655,N_14816);
and U19269 (N_19269,N_13794,N_13477);
or U19270 (N_19270,N_15900,N_13735);
or U19271 (N_19271,N_13150,N_14100);
nand U19272 (N_19272,N_14371,N_14653);
nor U19273 (N_19273,N_14330,N_13455);
nor U19274 (N_19274,N_14394,N_12863);
or U19275 (N_19275,N_12567,N_12476);
nand U19276 (N_19276,N_14790,N_12143);
xor U19277 (N_19277,N_12832,N_12114);
nand U19278 (N_19278,N_13073,N_15384);
xnor U19279 (N_19279,N_15206,N_15780);
nand U19280 (N_19280,N_14076,N_12871);
nor U19281 (N_19281,N_14525,N_12610);
nand U19282 (N_19282,N_15073,N_15253);
or U19283 (N_19283,N_14490,N_15613);
and U19284 (N_19284,N_13933,N_13091);
nor U19285 (N_19285,N_13997,N_15292);
xor U19286 (N_19286,N_14772,N_13841);
xnor U19287 (N_19287,N_15371,N_14106);
nand U19288 (N_19288,N_14939,N_15891);
or U19289 (N_19289,N_12294,N_15266);
and U19290 (N_19290,N_13488,N_14496);
nor U19291 (N_19291,N_15109,N_14140);
and U19292 (N_19292,N_14878,N_14708);
nand U19293 (N_19293,N_14122,N_13564);
or U19294 (N_19294,N_15759,N_15222);
nor U19295 (N_19295,N_15499,N_14612);
or U19296 (N_19296,N_13879,N_14512);
or U19297 (N_19297,N_12808,N_14003);
or U19298 (N_19298,N_14021,N_12577);
and U19299 (N_19299,N_15498,N_14563);
or U19300 (N_19300,N_12746,N_15692);
or U19301 (N_19301,N_14816,N_12444);
nand U19302 (N_19302,N_14066,N_13908);
nor U19303 (N_19303,N_15638,N_12355);
nor U19304 (N_19304,N_14603,N_15969);
or U19305 (N_19305,N_13499,N_13045);
xor U19306 (N_19306,N_14595,N_12685);
xnor U19307 (N_19307,N_13441,N_15134);
nand U19308 (N_19308,N_12138,N_15621);
xnor U19309 (N_19309,N_12220,N_13694);
or U19310 (N_19310,N_12052,N_12253);
or U19311 (N_19311,N_12755,N_15908);
nor U19312 (N_19312,N_14497,N_13771);
nor U19313 (N_19313,N_13974,N_12310);
and U19314 (N_19314,N_13512,N_15073);
nand U19315 (N_19315,N_12078,N_15891);
or U19316 (N_19316,N_15338,N_15850);
and U19317 (N_19317,N_14330,N_12459);
nor U19318 (N_19318,N_14989,N_13629);
nor U19319 (N_19319,N_14686,N_15437);
nand U19320 (N_19320,N_12591,N_12621);
nand U19321 (N_19321,N_15692,N_15782);
nor U19322 (N_19322,N_15604,N_15483);
xor U19323 (N_19323,N_13190,N_12513);
or U19324 (N_19324,N_15698,N_15226);
or U19325 (N_19325,N_15953,N_13224);
and U19326 (N_19326,N_12967,N_12717);
xor U19327 (N_19327,N_15579,N_15205);
and U19328 (N_19328,N_12150,N_13027);
nor U19329 (N_19329,N_15511,N_14369);
xnor U19330 (N_19330,N_13560,N_15375);
or U19331 (N_19331,N_12753,N_14278);
nor U19332 (N_19332,N_12748,N_12337);
or U19333 (N_19333,N_15965,N_15361);
nor U19334 (N_19334,N_14543,N_12556);
nor U19335 (N_19335,N_14821,N_14689);
nor U19336 (N_19336,N_13178,N_15966);
nor U19337 (N_19337,N_12577,N_15354);
and U19338 (N_19338,N_14390,N_12921);
or U19339 (N_19339,N_13850,N_15164);
or U19340 (N_19340,N_15481,N_15952);
nor U19341 (N_19341,N_13173,N_14663);
nand U19342 (N_19342,N_15679,N_12223);
or U19343 (N_19343,N_12822,N_13167);
nand U19344 (N_19344,N_12873,N_15427);
or U19345 (N_19345,N_15106,N_15014);
nor U19346 (N_19346,N_13739,N_12327);
nor U19347 (N_19347,N_14945,N_13102);
nand U19348 (N_19348,N_12406,N_14124);
or U19349 (N_19349,N_15014,N_14711);
and U19350 (N_19350,N_15977,N_15832);
nand U19351 (N_19351,N_13839,N_13672);
nand U19352 (N_19352,N_15717,N_13725);
nor U19353 (N_19353,N_12129,N_13007);
xnor U19354 (N_19354,N_14110,N_13188);
nand U19355 (N_19355,N_14211,N_12725);
and U19356 (N_19356,N_12654,N_15999);
and U19357 (N_19357,N_13675,N_13463);
nand U19358 (N_19358,N_14022,N_14762);
nor U19359 (N_19359,N_13841,N_15012);
nor U19360 (N_19360,N_14558,N_12636);
or U19361 (N_19361,N_15127,N_15589);
nor U19362 (N_19362,N_13553,N_13531);
or U19363 (N_19363,N_15198,N_13448);
or U19364 (N_19364,N_14569,N_14054);
nor U19365 (N_19365,N_13192,N_12323);
or U19366 (N_19366,N_14430,N_14819);
nand U19367 (N_19367,N_13761,N_13401);
and U19368 (N_19368,N_14064,N_13730);
nand U19369 (N_19369,N_14481,N_15188);
nor U19370 (N_19370,N_14938,N_13647);
and U19371 (N_19371,N_13192,N_14920);
or U19372 (N_19372,N_14020,N_15071);
or U19373 (N_19373,N_14212,N_13119);
nor U19374 (N_19374,N_12133,N_12695);
and U19375 (N_19375,N_14567,N_15940);
nand U19376 (N_19376,N_14655,N_13172);
and U19377 (N_19377,N_14201,N_13044);
and U19378 (N_19378,N_12505,N_14760);
nor U19379 (N_19379,N_13311,N_15942);
nand U19380 (N_19380,N_12365,N_14862);
xnor U19381 (N_19381,N_12397,N_14860);
and U19382 (N_19382,N_12912,N_12094);
nand U19383 (N_19383,N_13289,N_12200);
nor U19384 (N_19384,N_15737,N_12207);
and U19385 (N_19385,N_15254,N_14030);
nor U19386 (N_19386,N_12778,N_14849);
nor U19387 (N_19387,N_14614,N_12617);
nand U19388 (N_19388,N_14359,N_13630);
nand U19389 (N_19389,N_14107,N_13905);
nor U19390 (N_19390,N_15384,N_14418);
xnor U19391 (N_19391,N_13098,N_13933);
nor U19392 (N_19392,N_12130,N_15946);
nand U19393 (N_19393,N_12629,N_13547);
nor U19394 (N_19394,N_13732,N_15369);
nand U19395 (N_19395,N_13393,N_15821);
and U19396 (N_19396,N_13032,N_13764);
nand U19397 (N_19397,N_13879,N_12646);
nor U19398 (N_19398,N_14813,N_12049);
nand U19399 (N_19399,N_13079,N_14318);
or U19400 (N_19400,N_12934,N_12439);
and U19401 (N_19401,N_12886,N_12629);
nand U19402 (N_19402,N_15348,N_15636);
or U19403 (N_19403,N_14050,N_12820);
nand U19404 (N_19404,N_12056,N_12188);
nor U19405 (N_19405,N_12859,N_15841);
nor U19406 (N_19406,N_15225,N_14029);
and U19407 (N_19407,N_15336,N_12945);
or U19408 (N_19408,N_15809,N_13512);
nor U19409 (N_19409,N_12405,N_14289);
nor U19410 (N_19410,N_12035,N_15823);
nand U19411 (N_19411,N_12166,N_14088);
or U19412 (N_19412,N_12267,N_13494);
or U19413 (N_19413,N_13848,N_14342);
and U19414 (N_19414,N_14939,N_13571);
nor U19415 (N_19415,N_13541,N_15446);
xnor U19416 (N_19416,N_15821,N_15138);
nor U19417 (N_19417,N_15335,N_14409);
or U19418 (N_19418,N_12462,N_15281);
and U19419 (N_19419,N_12156,N_13499);
or U19420 (N_19420,N_13225,N_15316);
nand U19421 (N_19421,N_13355,N_13715);
nor U19422 (N_19422,N_13029,N_14742);
and U19423 (N_19423,N_14291,N_15904);
nor U19424 (N_19424,N_14798,N_15292);
and U19425 (N_19425,N_14414,N_15248);
or U19426 (N_19426,N_14040,N_12325);
nor U19427 (N_19427,N_15488,N_15078);
and U19428 (N_19428,N_12508,N_12412);
or U19429 (N_19429,N_15604,N_12199);
and U19430 (N_19430,N_14208,N_15957);
nand U19431 (N_19431,N_14278,N_14060);
nand U19432 (N_19432,N_12133,N_12859);
and U19433 (N_19433,N_12796,N_15629);
xor U19434 (N_19434,N_14381,N_12018);
nor U19435 (N_19435,N_13706,N_12497);
or U19436 (N_19436,N_14868,N_13109);
nand U19437 (N_19437,N_12875,N_15639);
or U19438 (N_19438,N_13745,N_13200);
nand U19439 (N_19439,N_15130,N_12731);
xor U19440 (N_19440,N_12412,N_14860);
nor U19441 (N_19441,N_15685,N_14243);
or U19442 (N_19442,N_12573,N_12914);
or U19443 (N_19443,N_13828,N_12367);
nor U19444 (N_19444,N_15562,N_13061);
nor U19445 (N_19445,N_13648,N_12094);
nor U19446 (N_19446,N_14667,N_15725);
or U19447 (N_19447,N_15667,N_14476);
nor U19448 (N_19448,N_13385,N_14044);
and U19449 (N_19449,N_12658,N_13946);
or U19450 (N_19450,N_14422,N_14712);
xnor U19451 (N_19451,N_15108,N_15824);
and U19452 (N_19452,N_15347,N_12067);
nor U19453 (N_19453,N_14743,N_15048);
and U19454 (N_19454,N_12412,N_15015);
nor U19455 (N_19455,N_14248,N_15778);
and U19456 (N_19456,N_15288,N_13761);
nand U19457 (N_19457,N_13903,N_13487);
or U19458 (N_19458,N_14215,N_15013);
nand U19459 (N_19459,N_15259,N_14432);
or U19460 (N_19460,N_15493,N_15153);
nor U19461 (N_19461,N_13512,N_12780);
nand U19462 (N_19462,N_15832,N_13689);
nor U19463 (N_19463,N_13496,N_13469);
nor U19464 (N_19464,N_15767,N_14763);
nand U19465 (N_19465,N_14082,N_15544);
or U19466 (N_19466,N_12978,N_13821);
nand U19467 (N_19467,N_12107,N_12898);
nand U19468 (N_19468,N_14358,N_12947);
or U19469 (N_19469,N_14651,N_13817);
and U19470 (N_19470,N_13094,N_15581);
and U19471 (N_19471,N_15835,N_12003);
xnor U19472 (N_19472,N_13902,N_15428);
nor U19473 (N_19473,N_15710,N_13260);
nand U19474 (N_19474,N_13425,N_12699);
xnor U19475 (N_19475,N_14862,N_13761);
nand U19476 (N_19476,N_14410,N_14638);
nand U19477 (N_19477,N_12925,N_12263);
and U19478 (N_19478,N_14930,N_14152);
xnor U19479 (N_19479,N_15609,N_14608);
nand U19480 (N_19480,N_12246,N_13244);
or U19481 (N_19481,N_12639,N_15175);
or U19482 (N_19482,N_12717,N_12719);
xnor U19483 (N_19483,N_13749,N_15017);
and U19484 (N_19484,N_14861,N_15830);
nand U19485 (N_19485,N_15367,N_13281);
and U19486 (N_19486,N_12667,N_15690);
nor U19487 (N_19487,N_12419,N_12713);
and U19488 (N_19488,N_14355,N_12675);
and U19489 (N_19489,N_13845,N_12809);
and U19490 (N_19490,N_14367,N_14675);
and U19491 (N_19491,N_13113,N_15716);
nand U19492 (N_19492,N_14337,N_12547);
and U19493 (N_19493,N_12417,N_12568);
and U19494 (N_19494,N_13576,N_12388);
nand U19495 (N_19495,N_12436,N_13579);
or U19496 (N_19496,N_13891,N_14713);
nor U19497 (N_19497,N_13700,N_15908);
nor U19498 (N_19498,N_12371,N_12233);
nor U19499 (N_19499,N_13744,N_13957);
or U19500 (N_19500,N_15044,N_15614);
and U19501 (N_19501,N_15584,N_14956);
nand U19502 (N_19502,N_15793,N_15630);
nand U19503 (N_19503,N_15527,N_13192);
nor U19504 (N_19504,N_14641,N_13330);
and U19505 (N_19505,N_14556,N_13205);
nand U19506 (N_19506,N_14692,N_12252);
nor U19507 (N_19507,N_12348,N_13769);
nand U19508 (N_19508,N_13019,N_12131);
or U19509 (N_19509,N_14488,N_14833);
or U19510 (N_19510,N_15714,N_13000);
and U19511 (N_19511,N_14466,N_14916);
or U19512 (N_19512,N_12801,N_14838);
and U19513 (N_19513,N_13937,N_13695);
nor U19514 (N_19514,N_12991,N_12543);
nand U19515 (N_19515,N_13321,N_15214);
nor U19516 (N_19516,N_14321,N_14301);
nand U19517 (N_19517,N_15395,N_15161);
and U19518 (N_19518,N_14195,N_15285);
or U19519 (N_19519,N_12331,N_12361);
nand U19520 (N_19520,N_15981,N_14527);
nor U19521 (N_19521,N_12053,N_13876);
nand U19522 (N_19522,N_13475,N_12459);
or U19523 (N_19523,N_14414,N_15050);
nand U19524 (N_19524,N_15514,N_14073);
nand U19525 (N_19525,N_14853,N_12412);
and U19526 (N_19526,N_13510,N_15412);
nand U19527 (N_19527,N_14671,N_15474);
or U19528 (N_19528,N_14902,N_13231);
and U19529 (N_19529,N_13716,N_12078);
or U19530 (N_19530,N_14182,N_14397);
and U19531 (N_19531,N_12850,N_14363);
nor U19532 (N_19532,N_12695,N_12377);
nor U19533 (N_19533,N_14115,N_14630);
nand U19534 (N_19534,N_12328,N_13978);
nand U19535 (N_19535,N_12140,N_15862);
nor U19536 (N_19536,N_12193,N_15129);
and U19537 (N_19537,N_12764,N_12143);
nor U19538 (N_19538,N_13523,N_15943);
nor U19539 (N_19539,N_15719,N_14849);
nand U19540 (N_19540,N_13825,N_12492);
nand U19541 (N_19541,N_13241,N_12720);
or U19542 (N_19542,N_14868,N_13332);
nor U19543 (N_19543,N_15196,N_15041);
nand U19544 (N_19544,N_14569,N_13681);
or U19545 (N_19545,N_15782,N_12355);
nand U19546 (N_19546,N_14611,N_15997);
or U19547 (N_19547,N_14343,N_12363);
or U19548 (N_19548,N_15807,N_13305);
nand U19549 (N_19549,N_15954,N_13873);
nand U19550 (N_19550,N_12169,N_14945);
xor U19551 (N_19551,N_13956,N_12102);
nor U19552 (N_19552,N_12113,N_12907);
nor U19553 (N_19553,N_13425,N_13884);
nand U19554 (N_19554,N_12845,N_15064);
nor U19555 (N_19555,N_15666,N_12739);
or U19556 (N_19556,N_12982,N_14185);
nor U19557 (N_19557,N_13013,N_14449);
and U19558 (N_19558,N_13205,N_15188);
nor U19559 (N_19559,N_14678,N_15447);
or U19560 (N_19560,N_12529,N_14662);
and U19561 (N_19561,N_12040,N_12400);
xor U19562 (N_19562,N_14226,N_12296);
nand U19563 (N_19563,N_13667,N_14632);
or U19564 (N_19564,N_12102,N_12144);
xor U19565 (N_19565,N_15733,N_13128);
nor U19566 (N_19566,N_13687,N_13457);
or U19567 (N_19567,N_15323,N_13742);
and U19568 (N_19568,N_15390,N_13970);
nor U19569 (N_19569,N_14947,N_13737);
nor U19570 (N_19570,N_14085,N_13686);
xnor U19571 (N_19571,N_12081,N_15730);
nor U19572 (N_19572,N_13403,N_13970);
nor U19573 (N_19573,N_14161,N_12480);
nor U19574 (N_19574,N_12216,N_12771);
nor U19575 (N_19575,N_13774,N_12593);
nor U19576 (N_19576,N_14462,N_15112);
and U19577 (N_19577,N_13687,N_12877);
nor U19578 (N_19578,N_14001,N_15559);
nand U19579 (N_19579,N_13722,N_15520);
nor U19580 (N_19580,N_12381,N_14481);
and U19581 (N_19581,N_12634,N_13703);
nor U19582 (N_19582,N_14195,N_15000);
nor U19583 (N_19583,N_13800,N_12199);
nand U19584 (N_19584,N_13002,N_12827);
or U19585 (N_19585,N_14848,N_13506);
xor U19586 (N_19586,N_12460,N_13546);
and U19587 (N_19587,N_14235,N_12178);
and U19588 (N_19588,N_13170,N_14468);
nor U19589 (N_19589,N_14058,N_15451);
and U19590 (N_19590,N_12491,N_13893);
or U19591 (N_19591,N_15586,N_13070);
or U19592 (N_19592,N_14091,N_13644);
or U19593 (N_19593,N_14495,N_12461);
or U19594 (N_19594,N_15926,N_12016);
and U19595 (N_19595,N_14148,N_14353);
xnor U19596 (N_19596,N_13983,N_15211);
or U19597 (N_19597,N_12663,N_12177);
or U19598 (N_19598,N_14352,N_12537);
and U19599 (N_19599,N_14247,N_15620);
or U19600 (N_19600,N_13327,N_14537);
nand U19601 (N_19601,N_12346,N_15899);
and U19602 (N_19602,N_13211,N_15045);
nand U19603 (N_19603,N_12151,N_14007);
nor U19604 (N_19604,N_13721,N_13696);
or U19605 (N_19605,N_12616,N_15351);
nor U19606 (N_19606,N_15854,N_13826);
and U19607 (N_19607,N_15299,N_15036);
and U19608 (N_19608,N_15194,N_14653);
and U19609 (N_19609,N_14025,N_15399);
nand U19610 (N_19610,N_12089,N_12177);
and U19611 (N_19611,N_12441,N_15408);
nand U19612 (N_19612,N_12222,N_15673);
and U19613 (N_19613,N_12365,N_12559);
or U19614 (N_19614,N_15710,N_14443);
nand U19615 (N_19615,N_12497,N_12242);
or U19616 (N_19616,N_13424,N_13455);
or U19617 (N_19617,N_15202,N_15200);
nand U19618 (N_19618,N_13168,N_13939);
and U19619 (N_19619,N_13878,N_12453);
nand U19620 (N_19620,N_13040,N_15466);
and U19621 (N_19621,N_13457,N_15665);
nand U19622 (N_19622,N_13521,N_13051);
xnor U19623 (N_19623,N_13997,N_12737);
nand U19624 (N_19624,N_15574,N_12058);
nand U19625 (N_19625,N_13341,N_13684);
and U19626 (N_19626,N_12159,N_14029);
nor U19627 (N_19627,N_14287,N_12609);
nand U19628 (N_19628,N_13380,N_13993);
nor U19629 (N_19629,N_13720,N_14993);
xnor U19630 (N_19630,N_14861,N_13525);
or U19631 (N_19631,N_12581,N_15386);
nand U19632 (N_19632,N_13796,N_15927);
nor U19633 (N_19633,N_12478,N_12184);
xnor U19634 (N_19634,N_15554,N_14602);
or U19635 (N_19635,N_14627,N_13481);
and U19636 (N_19636,N_13914,N_13648);
nand U19637 (N_19637,N_13629,N_15852);
and U19638 (N_19638,N_13960,N_13411);
and U19639 (N_19639,N_12980,N_14370);
nand U19640 (N_19640,N_13587,N_14011);
nor U19641 (N_19641,N_13242,N_14569);
nand U19642 (N_19642,N_14069,N_13453);
and U19643 (N_19643,N_14307,N_14572);
and U19644 (N_19644,N_14386,N_12504);
or U19645 (N_19645,N_15047,N_13880);
nor U19646 (N_19646,N_15733,N_14770);
or U19647 (N_19647,N_15401,N_15384);
and U19648 (N_19648,N_14309,N_15674);
and U19649 (N_19649,N_13565,N_15433);
or U19650 (N_19650,N_13125,N_14867);
nand U19651 (N_19651,N_12266,N_13633);
and U19652 (N_19652,N_13901,N_14107);
and U19653 (N_19653,N_13930,N_13351);
nor U19654 (N_19654,N_13069,N_12843);
or U19655 (N_19655,N_15487,N_12588);
or U19656 (N_19656,N_15430,N_13932);
or U19657 (N_19657,N_15419,N_14270);
nor U19658 (N_19658,N_13896,N_13822);
and U19659 (N_19659,N_12825,N_12767);
nor U19660 (N_19660,N_15776,N_13290);
xnor U19661 (N_19661,N_12112,N_14681);
xnor U19662 (N_19662,N_14316,N_14219);
or U19663 (N_19663,N_14664,N_12697);
and U19664 (N_19664,N_13516,N_13678);
and U19665 (N_19665,N_15185,N_14067);
nor U19666 (N_19666,N_13657,N_12687);
nor U19667 (N_19667,N_15538,N_13830);
nand U19668 (N_19668,N_14973,N_12985);
nor U19669 (N_19669,N_13943,N_15068);
and U19670 (N_19670,N_13516,N_15130);
nand U19671 (N_19671,N_12725,N_12678);
nand U19672 (N_19672,N_14594,N_14849);
and U19673 (N_19673,N_12537,N_13617);
nand U19674 (N_19674,N_13342,N_14666);
xor U19675 (N_19675,N_15719,N_12096);
and U19676 (N_19676,N_15319,N_13605);
nand U19677 (N_19677,N_13265,N_13260);
and U19678 (N_19678,N_15913,N_14459);
and U19679 (N_19679,N_13863,N_15299);
nor U19680 (N_19680,N_13571,N_14019);
and U19681 (N_19681,N_12558,N_15274);
nand U19682 (N_19682,N_15040,N_12883);
and U19683 (N_19683,N_15349,N_12984);
xnor U19684 (N_19684,N_15031,N_13083);
nor U19685 (N_19685,N_15870,N_14194);
xor U19686 (N_19686,N_12646,N_14591);
or U19687 (N_19687,N_14589,N_12492);
nand U19688 (N_19688,N_12919,N_14021);
nand U19689 (N_19689,N_13048,N_15719);
nor U19690 (N_19690,N_14872,N_15536);
or U19691 (N_19691,N_12194,N_12046);
xnor U19692 (N_19692,N_15582,N_14249);
or U19693 (N_19693,N_14922,N_15357);
or U19694 (N_19694,N_15999,N_12613);
and U19695 (N_19695,N_15800,N_12100);
or U19696 (N_19696,N_15335,N_12625);
or U19697 (N_19697,N_15920,N_13867);
and U19698 (N_19698,N_12025,N_12758);
or U19699 (N_19699,N_15472,N_12338);
nand U19700 (N_19700,N_15830,N_15617);
nand U19701 (N_19701,N_12043,N_14571);
nor U19702 (N_19702,N_13997,N_14627);
or U19703 (N_19703,N_12248,N_14378);
nor U19704 (N_19704,N_12996,N_15829);
and U19705 (N_19705,N_13076,N_15653);
nand U19706 (N_19706,N_15021,N_14574);
nor U19707 (N_19707,N_13642,N_14201);
xor U19708 (N_19708,N_13143,N_12868);
or U19709 (N_19709,N_15042,N_14701);
or U19710 (N_19710,N_14294,N_15388);
nor U19711 (N_19711,N_14415,N_15472);
and U19712 (N_19712,N_13500,N_12476);
and U19713 (N_19713,N_15576,N_12740);
nor U19714 (N_19714,N_14672,N_14864);
or U19715 (N_19715,N_13343,N_12343);
nor U19716 (N_19716,N_12119,N_15759);
and U19717 (N_19717,N_12679,N_13868);
or U19718 (N_19718,N_14547,N_15716);
nor U19719 (N_19719,N_15670,N_15935);
or U19720 (N_19720,N_14318,N_13906);
nor U19721 (N_19721,N_15982,N_15595);
nand U19722 (N_19722,N_13236,N_14968);
xnor U19723 (N_19723,N_12417,N_15936);
nor U19724 (N_19724,N_12987,N_13807);
nand U19725 (N_19725,N_12803,N_15884);
xor U19726 (N_19726,N_12213,N_13193);
nor U19727 (N_19727,N_15723,N_15625);
xnor U19728 (N_19728,N_12140,N_13145);
nor U19729 (N_19729,N_12303,N_14212);
and U19730 (N_19730,N_15133,N_15760);
or U19731 (N_19731,N_15536,N_13193);
or U19732 (N_19732,N_15729,N_13438);
nor U19733 (N_19733,N_12646,N_12769);
nor U19734 (N_19734,N_15323,N_13027);
nand U19735 (N_19735,N_14624,N_15934);
and U19736 (N_19736,N_12600,N_14968);
or U19737 (N_19737,N_14547,N_12154);
xnor U19738 (N_19738,N_13286,N_13461);
or U19739 (N_19739,N_12859,N_14434);
xor U19740 (N_19740,N_12000,N_15001);
and U19741 (N_19741,N_14200,N_15154);
nor U19742 (N_19742,N_12949,N_12228);
nand U19743 (N_19743,N_12801,N_13407);
or U19744 (N_19744,N_15289,N_15546);
nand U19745 (N_19745,N_12125,N_12463);
nand U19746 (N_19746,N_15584,N_14247);
or U19747 (N_19747,N_14886,N_15881);
nor U19748 (N_19748,N_15626,N_15311);
nor U19749 (N_19749,N_13339,N_12592);
nor U19750 (N_19750,N_14499,N_13405);
nor U19751 (N_19751,N_15488,N_14470);
or U19752 (N_19752,N_15898,N_15205);
xor U19753 (N_19753,N_14964,N_15886);
or U19754 (N_19754,N_12999,N_13704);
nand U19755 (N_19755,N_13180,N_14971);
xnor U19756 (N_19756,N_13864,N_14895);
or U19757 (N_19757,N_15773,N_14315);
nor U19758 (N_19758,N_14350,N_15122);
nand U19759 (N_19759,N_13844,N_13313);
and U19760 (N_19760,N_13488,N_13000);
xor U19761 (N_19761,N_14378,N_14461);
xor U19762 (N_19762,N_13706,N_13442);
or U19763 (N_19763,N_13779,N_15424);
nor U19764 (N_19764,N_13750,N_13733);
and U19765 (N_19765,N_13151,N_14828);
nor U19766 (N_19766,N_13793,N_12633);
and U19767 (N_19767,N_13046,N_15135);
nand U19768 (N_19768,N_12231,N_14437);
nand U19769 (N_19769,N_15104,N_14535);
nand U19770 (N_19770,N_13747,N_13974);
nor U19771 (N_19771,N_14025,N_13584);
nor U19772 (N_19772,N_15138,N_14497);
and U19773 (N_19773,N_12410,N_13286);
nand U19774 (N_19774,N_15689,N_13536);
nand U19775 (N_19775,N_14717,N_15183);
and U19776 (N_19776,N_12972,N_12889);
nand U19777 (N_19777,N_12875,N_14147);
nor U19778 (N_19778,N_12383,N_13170);
or U19779 (N_19779,N_12952,N_15390);
nor U19780 (N_19780,N_12444,N_15614);
nand U19781 (N_19781,N_12593,N_12704);
and U19782 (N_19782,N_12030,N_15326);
nand U19783 (N_19783,N_13850,N_12198);
or U19784 (N_19784,N_14571,N_12489);
nand U19785 (N_19785,N_13928,N_14400);
nand U19786 (N_19786,N_12252,N_13672);
nand U19787 (N_19787,N_15085,N_15413);
or U19788 (N_19788,N_13954,N_12624);
nand U19789 (N_19789,N_12535,N_14049);
and U19790 (N_19790,N_15706,N_12201);
nor U19791 (N_19791,N_12279,N_13334);
nand U19792 (N_19792,N_15536,N_14605);
or U19793 (N_19793,N_14516,N_14414);
nand U19794 (N_19794,N_15640,N_13493);
xnor U19795 (N_19795,N_15693,N_13566);
or U19796 (N_19796,N_12671,N_15287);
or U19797 (N_19797,N_14670,N_12591);
nand U19798 (N_19798,N_12301,N_14423);
nor U19799 (N_19799,N_13986,N_13942);
xor U19800 (N_19800,N_15271,N_12879);
or U19801 (N_19801,N_15658,N_14964);
and U19802 (N_19802,N_15878,N_14042);
nor U19803 (N_19803,N_14844,N_14232);
and U19804 (N_19804,N_14095,N_12275);
xnor U19805 (N_19805,N_12907,N_13051);
or U19806 (N_19806,N_14892,N_14579);
and U19807 (N_19807,N_13732,N_14174);
nand U19808 (N_19808,N_14263,N_12596);
or U19809 (N_19809,N_12096,N_14330);
nand U19810 (N_19810,N_14329,N_15663);
nor U19811 (N_19811,N_13971,N_13287);
and U19812 (N_19812,N_12251,N_14526);
nand U19813 (N_19813,N_15620,N_13728);
or U19814 (N_19814,N_12142,N_15790);
or U19815 (N_19815,N_12637,N_13931);
or U19816 (N_19816,N_13156,N_14249);
or U19817 (N_19817,N_15852,N_12154);
nor U19818 (N_19818,N_13407,N_14634);
or U19819 (N_19819,N_12951,N_12235);
nand U19820 (N_19820,N_12216,N_15402);
or U19821 (N_19821,N_14850,N_14359);
nand U19822 (N_19822,N_12333,N_13587);
nor U19823 (N_19823,N_12456,N_15053);
nand U19824 (N_19824,N_12857,N_13217);
nor U19825 (N_19825,N_15329,N_12699);
nand U19826 (N_19826,N_13113,N_14693);
nor U19827 (N_19827,N_14459,N_12705);
nand U19828 (N_19828,N_15127,N_13615);
or U19829 (N_19829,N_14538,N_15762);
and U19830 (N_19830,N_15046,N_14206);
or U19831 (N_19831,N_14498,N_13331);
nand U19832 (N_19832,N_14745,N_14572);
xor U19833 (N_19833,N_13922,N_15476);
nand U19834 (N_19834,N_13754,N_15019);
nand U19835 (N_19835,N_12694,N_12149);
or U19836 (N_19836,N_12649,N_12301);
nand U19837 (N_19837,N_13233,N_15896);
nand U19838 (N_19838,N_12006,N_14626);
nor U19839 (N_19839,N_14972,N_12088);
and U19840 (N_19840,N_12571,N_15477);
or U19841 (N_19841,N_14089,N_14661);
or U19842 (N_19842,N_13687,N_15197);
nor U19843 (N_19843,N_14328,N_12645);
and U19844 (N_19844,N_12506,N_15227);
or U19845 (N_19845,N_13095,N_15536);
and U19846 (N_19846,N_15269,N_15683);
and U19847 (N_19847,N_15663,N_12599);
xnor U19848 (N_19848,N_14798,N_14153);
and U19849 (N_19849,N_15995,N_12680);
or U19850 (N_19850,N_15038,N_13637);
nand U19851 (N_19851,N_14910,N_13824);
and U19852 (N_19852,N_15506,N_15855);
or U19853 (N_19853,N_13344,N_13398);
nor U19854 (N_19854,N_13168,N_14190);
and U19855 (N_19855,N_15796,N_15280);
or U19856 (N_19856,N_12156,N_12627);
or U19857 (N_19857,N_14655,N_15355);
and U19858 (N_19858,N_15060,N_15322);
nor U19859 (N_19859,N_12607,N_12345);
and U19860 (N_19860,N_12793,N_14872);
nand U19861 (N_19861,N_14025,N_14895);
or U19862 (N_19862,N_15616,N_14330);
nor U19863 (N_19863,N_13324,N_13946);
or U19864 (N_19864,N_14199,N_14622);
nor U19865 (N_19865,N_13244,N_13886);
nand U19866 (N_19866,N_15883,N_13707);
and U19867 (N_19867,N_12193,N_13914);
and U19868 (N_19868,N_13262,N_14112);
nand U19869 (N_19869,N_14082,N_15406);
nor U19870 (N_19870,N_14305,N_14998);
and U19871 (N_19871,N_14156,N_15111);
nor U19872 (N_19872,N_13359,N_13859);
or U19873 (N_19873,N_14439,N_15980);
nand U19874 (N_19874,N_12361,N_13652);
and U19875 (N_19875,N_15502,N_13525);
nor U19876 (N_19876,N_13565,N_13962);
nor U19877 (N_19877,N_14162,N_12273);
nand U19878 (N_19878,N_14572,N_12511);
nor U19879 (N_19879,N_13426,N_15502);
and U19880 (N_19880,N_15551,N_14704);
nor U19881 (N_19881,N_13531,N_14811);
and U19882 (N_19882,N_13677,N_15642);
and U19883 (N_19883,N_12083,N_15502);
nand U19884 (N_19884,N_12189,N_15783);
nor U19885 (N_19885,N_12806,N_13254);
and U19886 (N_19886,N_13263,N_12784);
and U19887 (N_19887,N_13679,N_12399);
or U19888 (N_19888,N_14359,N_13115);
or U19889 (N_19889,N_14761,N_14061);
or U19890 (N_19890,N_14072,N_12462);
nor U19891 (N_19891,N_13076,N_14388);
nor U19892 (N_19892,N_15478,N_15661);
nand U19893 (N_19893,N_14565,N_14823);
nand U19894 (N_19894,N_15185,N_13973);
nand U19895 (N_19895,N_13791,N_12738);
nor U19896 (N_19896,N_13849,N_13113);
nand U19897 (N_19897,N_14308,N_13719);
nor U19898 (N_19898,N_15642,N_15277);
or U19899 (N_19899,N_13479,N_12071);
nand U19900 (N_19900,N_15042,N_15420);
nand U19901 (N_19901,N_14807,N_15405);
or U19902 (N_19902,N_14649,N_15127);
or U19903 (N_19903,N_13361,N_15118);
nand U19904 (N_19904,N_12659,N_12147);
nor U19905 (N_19905,N_12306,N_13492);
or U19906 (N_19906,N_12589,N_13007);
nand U19907 (N_19907,N_15393,N_13233);
nor U19908 (N_19908,N_15450,N_12824);
nand U19909 (N_19909,N_15772,N_14943);
nor U19910 (N_19910,N_13568,N_15943);
nand U19911 (N_19911,N_15103,N_15084);
and U19912 (N_19912,N_13516,N_12095);
or U19913 (N_19913,N_13287,N_15840);
nor U19914 (N_19914,N_12282,N_14305);
nand U19915 (N_19915,N_15551,N_13455);
and U19916 (N_19916,N_12396,N_14253);
nand U19917 (N_19917,N_12821,N_13018);
and U19918 (N_19918,N_15595,N_13909);
and U19919 (N_19919,N_13133,N_14297);
or U19920 (N_19920,N_12126,N_12957);
or U19921 (N_19921,N_15042,N_13666);
nor U19922 (N_19922,N_12706,N_13706);
nand U19923 (N_19923,N_12220,N_14638);
nand U19924 (N_19924,N_13039,N_14388);
and U19925 (N_19925,N_14555,N_12541);
nor U19926 (N_19926,N_13124,N_13801);
nor U19927 (N_19927,N_13823,N_15540);
nand U19928 (N_19928,N_13509,N_15655);
nand U19929 (N_19929,N_12481,N_15918);
and U19930 (N_19930,N_13782,N_15990);
and U19931 (N_19931,N_12360,N_13718);
or U19932 (N_19932,N_12811,N_12742);
nand U19933 (N_19933,N_15232,N_14408);
nor U19934 (N_19934,N_14388,N_13887);
nor U19935 (N_19935,N_12074,N_12417);
nand U19936 (N_19936,N_15036,N_15022);
and U19937 (N_19937,N_13396,N_15617);
nor U19938 (N_19938,N_15831,N_14475);
and U19939 (N_19939,N_13511,N_12628);
nand U19940 (N_19940,N_14266,N_13694);
and U19941 (N_19941,N_15533,N_12460);
nor U19942 (N_19942,N_15056,N_14220);
nand U19943 (N_19943,N_15785,N_15482);
or U19944 (N_19944,N_15176,N_13398);
and U19945 (N_19945,N_15736,N_12081);
xnor U19946 (N_19946,N_14793,N_13178);
or U19947 (N_19947,N_12529,N_12982);
xor U19948 (N_19948,N_12602,N_13506);
nor U19949 (N_19949,N_12496,N_15538);
or U19950 (N_19950,N_15997,N_12097);
and U19951 (N_19951,N_12597,N_15748);
nor U19952 (N_19952,N_13175,N_12981);
or U19953 (N_19953,N_12552,N_12557);
or U19954 (N_19954,N_14728,N_14337);
or U19955 (N_19955,N_12361,N_13989);
or U19956 (N_19956,N_15501,N_13285);
xnor U19957 (N_19957,N_13961,N_15346);
nand U19958 (N_19958,N_12689,N_12008);
nor U19959 (N_19959,N_13073,N_15484);
nor U19960 (N_19960,N_14395,N_15246);
nor U19961 (N_19961,N_13760,N_13723);
or U19962 (N_19962,N_13079,N_13598);
and U19963 (N_19963,N_15891,N_14270);
nand U19964 (N_19964,N_13788,N_14779);
nand U19965 (N_19965,N_14235,N_12988);
and U19966 (N_19966,N_14886,N_15128);
and U19967 (N_19967,N_12421,N_14060);
nand U19968 (N_19968,N_12255,N_14348);
nor U19969 (N_19969,N_12358,N_12885);
nand U19970 (N_19970,N_15378,N_14604);
nand U19971 (N_19971,N_12818,N_13918);
and U19972 (N_19972,N_14812,N_13069);
nand U19973 (N_19973,N_13661,N_14460);
xnor U19974 (N_19974,N_15439,N_12308);
or U19975 (N_19975,N_13926,N_12607);
or U19976 (N_19976,N_15677,N_14644);
nor U19977 (N_19977,N_12867,N_12044);
and U19978 (N_19978,N_12400,N_12106);
and U19979 (N_19979,N_14127,N_14783);
nor U19980 (N_19980,N_14200,N_14861);
nand U19981 (N_19981,N_14624,N_15160);
xor U19982 (N_19982,N_14577,N_13646);
nor U19983 (N_19983,N_14357,N_15773);
nor U19984 (N_19984,N_15015,N_15000);
xor U19985 (N_19985,N_12300,N_15266);
or U19986 (N_19986,N_14227,N_14062);
xnor U19987 (N_19987,N_15966,N_14890);
nor U19988 (N_19988,N_14379,N_14128);
nor U19989 (N_19989,N_13739,N_14665);
and U19990 (N_19990,N_15578,N_14474);
nor U19991 (N_19991,N_14697,N_13595);
nor U19992 (N_19992,N_14087,N_15533);
nor U19993 (N_19993,N_14791,N_15958);
nor U19994 (N_19994,N_15670,N_13733);
nor U19995 (N_19995,N_15622,N_14259);
nand U19996 (N_19996,N_13082,N_13900);
or U19997 (N_19997,N_14091,N_14119);
nand U19998 (N_19998,N_14505,N_15359);
or U19999 (N_19999,N_12450,N_12715);
nand UO_0 (O_0,N_18081,N_19755);
nor UO_1 (O_1,N_17237,N_17514);
and UO_2 (O_2,N_18126,N_16285);
nand UO_3 (O_3,N_17895,N_17108);
nand UO_4 (O_4,N_16789,N_19383);
nand UO_5 (O_5,N_16640,N_18349);
and UO_6 (O_6,N_17711,N_16979);
nor UO_7 (O_7,N_18446,N_16700);
nand UO_8 (O_8,N_19039,N_19047);
nand UO_9 (O_9,N_17433,N_19532);
and UO_10 (O_10,N_16553,N_16248);
nor UO_11 (O_11,N_19964,N_18336);
and UO_12 (O_12,N_19548,N_17678);
xnor UO_13 (O_13,N_19369,N_18186);
and UO_14 (O_14,N_18756,N_18686);
nor UO_15 (O_15,N_19052,N_19857);
nand UO_16 (O_16,N_19965,N_16103);
and UO_17 (O_17,N_17194,N_18688);
nand UO_18 (O_18,N_17291,N_19577);
or UO_19 (O_19,N_19542,N_17821);
nand UO_20 (O_20,N_16606,N_18922);
nor UO_21 (O_21,N_19404,N_16554);
nand UO_22 (O_22,N_17894,N_18045);
nor UO_23 (O_23,N_19635,N_18465);
or UO_24 (O_24,N_17335,N_18084);
nor UO_25 (O_25,N_18943,N_18921);
nand UO_26 (O_26,N_16311,N_18521);
and UO_27 (O_27,N_18280,N_16119);
or UO_28 (O_28,N_19596,N_17191);
or UO_29 (O_29,N_17540,N_18674);
nand UO_30 (O_30,N_17892,N_17208);
or UO_31 (O_31,N_17575,N_16550);
or UO_32 (O_32,N_16888,N_18005);
nor UO_33 (O_33,N_17284,N_19817);
and UO_34 (O_34,N_16824,N_19924);
nor UO_35 (O_35,N_16936,N_17765);
xor UO_36 (O_36,N_16319,N_16404);
nor UO_37 (O_37,N_18170,N_19425);
or UO_38 (O_38,N_17304,N_16942);
or UO_39 (O_39,N_17382,N_16494);
or UO_40 (O_40,N_19630,N_19076);
and UO_41 (O_41,N_18393,N_18306);
xnor UO_42 (O_42,N_18789,N_19767);
nand UO_43 (O_43,N_16926,N_19267);
xnor UO_44 (O_44,N_19847,N_19095);
or UO_45 (O_45,N_17622,N_17705);
xor UO_46 (O_46,N_16410,N_19364);
xor UO_47 (O_47,N_18980,N_18665);
nand UO_48 (O_48,N_16289,N_19725);
nand UO_49 (O_49,N_17756,N_16143);
nor UO_50 (O_50,N_18050,N_19862);
xnor UO_51 (O_51,N_17239,N_19412);
and UO_52 (O_52,N_17695,N_19141);
and UO_53 (O_53,N_17630,N_19509);
or UO_54 (O_54,N_17671,N_17613);
nor UO_55 (O_55,N_18405,N_18817);
nand UO_56 (O_56,N_16215,N_16266);
and UO_57 (O_57,N_18365,N_18046);
or UO_58 (O_58,N_16397,N_17295);
nand UO_59 (O_59,N_16389,N_17258);
and UO_60 (O_60,N_17449,N_16296);
and UO_61 (O_61,N_16474,N_18790);
nand UO_62 (O_62,N_17360,N_19950);
nor UO_63 (O_63,N_19982,N_17328);
xor UO_64 (O_64,N_17991,N_16676);
nand UO_65 (O_65,N_18488,N_16370);
or UO_66 (O_66,N_17617,N_19322);
or UO_67 (O_67,N_18165,N_17901);
and UO_68 (O_68,N_17105,N_18262);
nand UO_69 (O_69,N_17660,N_19539);
xnor UO_70 (O_70,N_19108,N_17106);
xnor UO_71 (O_71,N_16769,N_16573);
and UO_72 (O_72,N_18968,N_19538);
or UO_73 (O_73,N_17672,N_19703);
nand UO_74 (O_74,N_18531,N_18734);
and UO_75 (O_75,N_16548,N_18088);
and UO_76 (O_76,N_18244,N_18399);
or UO_77 (O_77,N_17791,N_16866);
and UO_78 (O_78,N_18568,N_19759);
nor UO_79 (O_79,N_17324,N_16533);
xor UO_80 (O_80,N_16287,N_19525);
or UO_81 (O_81,N_19714,N_17506);
nor UO_82 (O_82,N_19443,N_18408);
or UO_83 (O_83,N_17859,N_19062);
and UO_84 (O_84,N_18588,N_16278);
nor UO_85 (O_85,N_18497,N_19566);
and UO_86 (O_86,N_18247,N_19331);
nor UO_87 (O_87,N_17550,N_16381);
and UO_88 (O_88,N_19956,N_18845);
nor UO_89 (O_89,N_17992,N_19027);
and UO_90 (O_90,N_18600,N_16250);
nand UO_91 (O_91,N_19861,N_16368);
nor UO_92 (O_92,N_17225,N_19968);
and UO_93 (O_93,N_17307,N_19022);
and UO_94 (O_94,N_16727,N_16605);
nand UO_95 (O_95,N_16575,N_16298);
and UO_96 (O_96,N_19988,N_18622);
and UO_97 (O_97,N_17840,N_17042);
nor UO_98 (O_98,N_16776,N_19488);
xor UO_99 (O_99,N_18551,N_16168);
or UO_100 (O_100,N_18353,N_16637);
nor UO_101 (O_101,N_17132,N_16986);
and UO_102 (O_102,N_16037,N_17511);
nor UO_103 (O_103,N_16642,N_18499);
and UO_104 (O_104,N_17077,N_18270);
and UO_105 (O_105,N_18636,N_16171);
or UO_106 (O_106,N_17940,N_19136);
nand UO_107 (O_107,N_19065,N_19948);
xnor UO_108 (O_108,N_17252,N_17885);
or UO_109 (O_109,N_19233,N_19049);
and UO_110 (O_110,N_19389,N_19892);
and UO_111 (O_111,N_16693,N_19563);
nor UO_112 (O_112,N_18206,N_19201);
or UO_113 (O_113,N_16929,N_17217);
and UO_114 (O_114,N_19117,N_19588);
and UO_115 (O_115,N_19453,N_17156);
nor UO_116 (O_116,N_17569,N_19698);
or UO_117 (O_117,N_19876,N_18683);
or UO_118 (O_118,N_17771,N_16204);
xor UO_119 (O_119,N_16188,N_17586);
or UO_120 (O_120,N_16797,N_17845);
nor UO_121 (O_121,N_16648,N_18424);
xnor UO_122 (O_122,N_17679,N_18664);
or UO_123 (O_123,N_17313,N_19820);
nand UO_124 (O_124,N_17759,N_19655);
nor UO_125 (O_125,N_17111,N_16763);
nand UO_126 (O_126,N_16105,N_19316);
or UO_127 (O_127,N_16387,N_17928);
or UO_128 (O_128,N_18212,N_17911);
or UO_129 (O_129,N_16326,N_19646);
nand UO_130 (O_130,N_17245,N_16601);
nor UO_131 (O_131,N_19942,N_16990);
nand UO_132 (O_132,N_17530,N_16898);
nor UO_133 (O_133,N_17603,N_19937);
and UO_134 (O_134,N_17084,N_17648);
nand UO_135 (O_135,N_18708,N_16257);
or UO_136 (O_136,N_19806,N_19301);
nor UO_137 (O_137,N_17721,N_18208);
or UO_138 (O_138,N_17097,N_16277);
and UO_139 (O_139,N_19702,N_17170);
and UO_140 (O_140,N_19273,N_16492);
nor UO_141 (O_141,N_17834,N_16411);
or UO_142 (O_142,N_19976,N_19887);
and UO_143 (O_143,N_17027,N_19911);
and UO_144 (O_144,N_17762,N_19585);
or UO_145 (O_145,N_16344,N_18461);
nor UO_146 (O_146,N_17137,N_17329);
nor UO_147 (O_147,N_16187,N_19036);
and UO_148 (O_148,N_16645,N_16226);
or UO_149 (O_149,N_18007,N_17471);
or UO_150 (O_150,N_16270,N_16292);
nand UO_151 (O_151,N_18555,N_19710);
nand UO_152 (O_152,N_18112,N_17456);
or UO_153 (O_153,N_18854,N_18750);
and UO_154 (O_154,N_19692,N_17776);
nand UO_155 (O_155,N_16371,N_19991);
or UO_156 (O_156,N_16200,N_17800);
nand UO_157 (O_157,N_19489,N_18073);
and UO_158 (O_158,N_18233,N_16682);
and UO_159 (O_159,N_18389,N_19208);
and UO_160 (O_160,N_18275,N_19206);
and UO_161 (O_161,N_19159,N_16881);
nor UO_162 (O_162,N_16546,N_16123);
and UO_163 (O_163,N_16707,N_16619);
nor UO_164 (O_164,N_16140,N_17260);
or UO_165 (O_165,N_16733,N_19699);
xnor UO_166 (O_166,N_18856,N_18070);
xor UO_167 (O_167,N_17167,N_18456);
or UO_168 (O_168,N_18362,N_16816);
and UO_169 (O_169,N_18550,N_17333);
or UO_170 (O_170,N_18787,N_17924);
nor UO_171 (O_171,N_17409,N_17350);
xor UO_172 (O_172,N_18114,N_16767);
and UO_173 (O_173,N_17107,N_17234);
nand UO_174 (O_174,N_19465,N_19707);
or UO_175 (O_175,N_19652,N_18272);
nor UO_176 (O_176,N_17383,N_19504);
or UO_177 (O_177,N_19665,N_16151);
nor UO_178 (O_178,N_18091,N_19860);
nor UO_179 (O_179,N_19713,N_18742);
nand UO_180 (O_180,N_16194,N_19120);
and UO_181 (O_181,N_19505,N_19954);
or UO_182 (O_182,N_17717,N_18455);
or UO_183 (O_183,N_17615,N_16668);
nand UO_184 (O_184,N_19602,N_17024);
and UO_185 (O_185,N_17726,N_17598);
nor UO_186 (O_186,N_18137,N_18462);
nor UO_187 (O_187,N_19407,N_18643);
and UO_188 (O_188,N_19545,N_16872);
or UO_189 (O_189,N_17311,N_18816);
and UO_190 (O_190,N_19546,N_19734);
or UO_191 (O_191,N_16953,N_19782);
nand UO_192 (O_192,N_17680,N_17031);
and UO_193 (O_193,N_17581,N_16070);
nor UO_194 (O_194,N_17308,N_17957);
nor UO_195 (O_195,N_16909,N_19105);
nand UO_196 (O_196,N_19793,N_16305);
nand UO_197 (O_197,N_19157,N_16076);
or UO_198 (O_198,N_16930,N_18694);
and UO_199 (O_199,N_16440,N_17210);
xnor UO_200 (O_200,N_18868,N_19653);
or UO_201 (O_201,N_17677,N_19321);
nor UO_202 (O_202,N_17782,N_17715);
and UO_203 (O_203,N_19448,N_19902);
nor UO_204 (O_204,N_17416,N_16906);
or UO_205 (O_205,N_18530,N_19753);
nor UO_206 (O_206,N_18189,N_19612);
or UO_207 (O_207,N_17698,N_17642);
nand UO_208 (O_208,N_18449,N_17430);
and UO_209 (O_209,N_19520,N_17766);
and UO_210 (O_210,N_17742,N_16832);
nor UO_211 (O_211,N_18298,N_16181);
xnor UO_212 (O_212,N_19003,N_16283);
and UO_213 (O_213,N_18809,N_17921);
nand UO_214 (O_214,N_19871,N_17257);
nand UO_215 (O_215,N_16599,N_16850);
nor UO_216 (O_216,N_16656,N_19720);
xnor UO_217 (O_217,N_17690,N_18532);
or UO_218 (O_218,N_17701,N_16290);
nor UO_219 (O_219,N_19867,N_17922);
xor UO_220 (O_220,N_19006,N_18970);
nor UO_221 (O_221,N_16473,N_16272);
nor UO_222 (O_222,N_19016,N_18235);
xor UO_223 (O_223,N_16975,N_17270);
and UO_224 (O_224,N_19040,N_19382);
nor UO_225 (O_225,N_18028,N_16674);
and UO_226 (O_226,N_18518,N_16026);
nor UO_227 (O_227,N_18426,N_18257);
and UO_228 (O_228,N_19373,N_18130);
and UO_229 (O_229,N_19107,N_16003);
nor UO_230 (O_230,N_17244,N_18769);
and UO_231 (O_231,N_18351,N_19730);
nor UO_232 (O_232,N_18895,N_17301);
nand UO_233 (O_233,N_18493,N_16350);
nand UO_234 (O_234,N_19439,N_19058);
nand UO_235 (O_235,N_17422,N_16454);
or UO_236 (O_236,N_19018,N_18295);
nand UO_237 (O_237,N_16995,N_17638);
xor UO_238 (O_238,N_16125,N_17413);
or UO_239 (O_239,N_17253,N_17875);
or UO_240 (O_240,N_19132,N_18867);
nand UO_241 (O_241,N_17990,N_17028);
nand UO_242 (O_242,N_18898,N_18011);
and UO_243 (O_243,N_16329,N_18229);
and UO_244 (O_244,N_19353,N_16099);
nand UO_245 (O_245,N_16600,N_16147);
and UO_246 (O_246,N_19952,N_19712);
xnor UO_247 (O_247,N_17224,N_17129);
and UO_248 (O_248,N_18710,N_16328);
nand UO_249 (O_249,N_19474,N_18090);
nor UO_250 (O_250,N_17853,N_18690);
nor UO_251 (O_251,N_16716,N_18754);
nor UO_252 (O_252,N_18181,N_18955);
nor UO_253 (O_253,N_19078,N_18207);
xnor UO_254 (O_254,N_16303,N_16864);
nand UO_255 (O_255,N_17976,N_16249);
and UO_256 (O_256,N_16386,N_17869);
nand UO_257 (O_257,N_17139,N_19926);
nor UO_258 (O_258,N_19181,N_18069);
xnor UO_259 (O_259,N_19481,N_16138);
nor UO_260 (O_260,N_16241,N_17819);
or UO_261 (O_261,N_18989,N_18603);
or UO_262 (O_262,N_16762,N_18075);
or UO_263 (O_263,N_16061,N_18318);
xor UO_264 (O_264,N_16524,N_16703);
and UO_265 (O_265,N_19145,N_18025);
nor UO_266 (O_266,N_18167,N_17793);
and UO_267 (O_267,N_17101,N_18434);
nor UO_268 (O_268,N_19930,N_18528);
and UO_269 (O_269,N_17442,N_16702);
and UO_270 (O_270,N_16876,N_17861);
or UO_271 (O_271,N_17355,N_16396);
or UO_272 (O_272,N_16378,N_19342);
and UO_273 (O_273,N_17346,N_17386);
or UO_274 (O_274,N_19754,N_18241);
and UO_275 (O_275,N_19330,N_19413);
xor UO_276 (O_276,N_17798,N_19056);
xnor UO_277 (O_277,N_19537,N_17220);
or UO_278 (O_278,N_17979,N_16192);
nand UO_279 (O_279,N_18000,N_19437);
and UO_280 (O_280,N_18038,N_18156);
nor UO_281 (O_281,N_18277,N_16587);
xor UO_282 (O_282,N_18224,N_19882);
xnor UO_283 (O_283,N_17482,N_17578);
nor UO_284 (O_284,N_18127,N_17956);
and UO_285 (O_285,N_19417,N_19900);
nor UO_286 (O_286,N_18273,N_16581);
nor UO_287 (O_287,N_16654,N_19051);
xnor UO_288 (O_288,N_17149,N_17938);
and UO_289 (O_289,N_18216,N_17264);
and UO_290 (O_290,N_18804,N_16114);
or UO_291 (O_291,N_17792,N_16346);
and UO_292 (O_292,N_18220,N_17009);
nor UO_293 (O_293,N_16110,N_19262);
nor UO_294 (O_294,N_17851,N_19883);
nand UO_295 (O_295,N_19476,N_18705);
nor UO_296 (O_296,N_19866,N_19220);
or UO_297 (O_297,N_17288,N_16176);
nand UO_298 (O_298,N_19628,N_18847);
xnor UO_299 (O_299,N_16155,N_16617);
nand UO_300 (O_300,N_17119,N_16013);
nand UO_301 (O_301,N_16288,N_17532);
or UO_302 (O_302,N_19651,N_19282);
nand UO_303 (O_303,N_16039,N_17183);
xor UO_304 (O_304,N_17808,N_19418);
and UO_305 (O_305,N_16803,N_19294);
xnor UO_306 (O_306,N_18391,N_18429);
or UO_307 (O_307,N_18320,N_16837);
nand UO_308 (O_308,N_17681,N_16994);
nor UO_309 (O_309,N_16996,N_18770);
nor UO_310 (O_310,N_19312,N_16313);
and UO_311 (O_311,N_17246,N_16603);
or UO_312 (O_312,N_16771,N_17344);
or UO_313 (O_313,N_16031,N_16661);
or UO_314 (O_314,N_18513,N_16914);
nand UO_315 (O_315,N_17040,N_16376);
nand UO_316 (O_316,N_17145,N_19172);
nand UO_317 (O_317,N_17152,N_16775);
or UO_318 (O_318,N_18481,N_18991);
nand UO_319 (O_319,N_19490,N_17395);
nand UO_320 (O_320,N_18155,N_16385);
nor UO_321 (O_321,N_19089,N_18982);
nand UO_322 (O_322,N_19271,N_16567);
nor UO_323 (O_323,N_19432,N_19020);
and UO_324 (O_324,N_19281,N_17790);
nor UO_325 (O_325,N_17038,N_16349);
and UO_326 (O_326,N_16591,N_19480);
and UO_327 (O_327,N_19696,N_17354);
and UO_328 (O_328,N_17973,N_17655);
and UO_329 (O_329,N_17459,N_18059);
or UO_330 (O_330,N_17987,N_17531);
or UO_331 (O_331,N_19973,N_18524);
and UO_332 (O_332,N_17589,N_17647);
or UO_333 (O_333,N_16858,N_16500);
nand UO_334 (O_334,N_18163,N_19263);
or UO_335 (O_335,N_18077,N_17188);
nand UO_336 (O_336,N_18733,N_19960);
nand UO_337 (O_337,N_16819,N_17135);
nor UO_338 (O_338,N_18193,N_16590);
and UO_339 (O_339,N_19589,N_17880);
xnor UO_340 (O_340,N_17146,N_18923);
and UO_341 (O_341,N_16859,N_18667);
and UO_342 (O_342,N_17666,N_19915);
or UO_343 (O_343,N_18080,N_17610);
nand UO_344 (O_344,N_17474,N_16046);
or UO_345 (O_345,N_17855,N_19365);
or UO_346 (O_346,N_16878,N_17803);
nor UO_347 (O_347,N_18617,N_19673);
or UO_348 (O_348,N_19739,N_18271);
or UO_349 (O_349,N_17890,N_18511);
nor UO_350 (O_350,N_17187,N_19641);
nor UO_351 (O_351,N_17047,N_18748);
xor UO_352 (O_352,N_19344,N_19317);
nand UO_353 (O_353,N_19958,N_17450);
or UO_354 (O_354,N_17525,N_18930);
and UO_355 (O_355,N_19656,N_16294);
and UO_356 (O_356,N_16425,N_16414);
or UO_357 (O_357,N_17545,N_18221);
or UO_358 (O_358,N_19977,N_17657);
or UO_359 (O_359,N_17127,N_17952);
nor UO_360 (O_360,N_16948,N_18027);
or UO_361 (O_361,N_19547,N_19324);
and UO_362 (O_362,N_18442,N_18700);
nor UO_363 (O_363,N_18715,N_18466);
nand UO_364 (O_364,N_16416,N_16467);
nor UO_365 (O_365,N_16615,N_18594);
or UO_366 (O_366,N_17891,N_16274);
nand UO_367 (O_367,N_16282,N_18650);
or UO_368 (O_368,N_19202,N_19446);
nor UO_369 (O_369,N_18213,N_16088);
and UO_370 (O_370,N_18065,N_17661);
and UO_371 (O_371,N_17917,N_19303);
and UO_372 (O_372,N_19463,N_17561);
or UO_373 (O_373,N_17585,N_18978);
or UO_374 (O_374,N_19278,N_16132);
nand UO_375 (O_375,N_17989,N_18385);
or UO_376 (O_376,N_16195,N_19593);
nand UO_377 (O_377,N_19099,N_16565);
xor UO_378 (O_378,N_18299,N_17888);
nor UO_379 (O_379,N_19530,N_19811);
nor UO_380 (O_380,N_18157,N_17420);
or UO_381 (O_381,N_17142,N_18198);
nand UO_382 (O_382,N_17763,N_19522);
and UO_383 (O_383,N_19460,N_16644);
nand UO_384 (O_384,N_17758,N_17261);
nor UO_385 (O_385,N_16985,N_19815);
or UO_386 (O_386,N_19744,N_18463);
xnor UO_387 (O_387,N_16822,N_19287);
or UO_388 (O_388,N_19875,N_18624);
nand UO_389 (O_389,N_19125,N_17085);
nor UO_390 (O_390,N_19347,N_18338);
or UO_391 (O_391,N_16256,N_19116);
nand UO_392 (O_392,N_16890,N_16972);
or UO_393 (O_393,N_16649,N_19097);
and UO_394 (O_394,N_17876,N_19598);
nand UO_395 (O_395,N_19388,N_18605);
or UO_396 (O_396,N_19776,N_17724);
or UO_397 (O_397,N_16388,N_18645);
nor UO_398 (O_398,N_19378,N_16631);
xor UO_399 (O_399,N_16920,N_19729);
nor UO_400 (O_400,N_17778,N_17637);
or UO_401 (O_401,N_18041,N_18939);
nand UO_402 (O_402,N_16937,N_18593);
or UO_403 (O_403,N_18337,N_17203);
and UO_404 (O_404,N_16475,N_16534);
nand UO_405 (O_405,N_16430,N_16586);
nor UO_406 (O_406,N_19803,N_17315);
xnor UO_407 (O_407,N_16987,N_18334);
and UO_408 (O_408,N_18510,N_19986);
or UO_409 (O_409,N_16163,N_19715);
nand UO_410 (O_410,N_16894,N_19493);
or UO_411 (O_411,N_19023,N_17838);
or UO_412 (O_412,N_17802,N_17983);
nor UO_413 (O_413,N_17478,N_16040);
xnor UO_414 (O_414,N_19786,N_18110);
nor UO_415 (O_415,N_18109,N_18347);
nor UO_416 (O_416,N_16398,N_18933);
and UO_417 (O_417,N_18205,N_16400);
and UO_418 (O_418,N_16744,N_18788);
nor UO_419 (O_419,N_18872,N_18899);
and UO_420 (O_420,N_19310,N_19224);
nor UO_421 (O_421,N_16889,N_16805);
nand UO_422 (O_422,N_18527,N_17612);
nand UO_423 (O_423,N_18776,N_16363);
and UO_424 (O_424,N_17011,N_18192);
or UO_425 (O_425,N_19138,N_18494);
and UO_426 (O_426,N_17697,N_18243);
nor UO_427 (O_427,N_17927,N_18698);
or UO_428 (O_428,N_18514,N_19349);
nor UO_429 (O_429,N_18687,N_18765);
nor UO_430 (O_430,N_16186,N_17556);
or UO_431 (O_431,N_19524,N_17968);
nor UO_432 (O_432,N_17863,N_17043);
and UO_433 (O_433,N_19156,N_17624);
nand UO_434 (O_434,N_17889,N_18714);
nor UO_435 (O_435,N_18726,N_18693);
xnor UO_436 (O_436,N_19916,N_19470);
or UO_437 (O_437,N_16549,N_17494);
or UO_438 (O_438,N_17186,N_17345);
nand UO_439 (O_439,N_17963,N_19780);
nor UO_440 (O_440,N_19377,N_16976);
and UO_441 (O_441,N_16836,N_19581);
and UO_442 (O_442,N_17384,N_16459);
and UO_443 (O_443,N_17879,N_19836);
nand UO_444 (O_444,N_17300,N_17691);
or UO_445 (O_445,N_18533,N_16035);
nor UO_446 (O_446,N_18954,N_16052);
and UO_447 (O_447,N_18730,N_16510);
nor UO_448 (O_448,N_17981,N_19716);
or UO_449 (O_449,N_16897,N_16687);
nand UO_450 (O_450,N_16112,N_17664);
nor UO_451 (O_451,N_19864,N_16596);
or UO_452 (O_452,N_16813,N_16232);
and UO_453 (O_453,N_17507,N_19726);
nor UO_454 (O_454,N_17848,N_19629);
or UO_455 (O_455,N_17099,N_16471);
or UO_456 (O_456,N_16323,N_16347);
nor UO_457 (O_457,N_19605,N_16185);
and UO_458 (O_458,N_16267,N_19048);
nor UO_459 (O_459,N_17683,N_19077);
or UO_460 (O_460,N_17219,N_17935);
nor UO_461 (O_461,N_19781,N_19697);
nor UO_462 (O_462,N_19093,N_19469);
or UO_463 (O_463,N_17251,N_19863);
or UO_464 (O_464,N_16028,N_17702);
nor UO_465 (O_465,N_16564,N_16952);
and UO_466 (O_466,N_17296,N_16765);
nor UO_467 (O_467,N_16810,N_19770);
nor UO_468 (O_468,N_17314,N_19005);
nor UO_469 (O_469,N_19936,N_17951);
nor UO_470 (O_470,N_16932,N_16020);
nand UO_471 (O_471,N_17760,N_17465);
nand UO_472 (O_472,N_16074,N_19167);
xnor UO_473 (O_473,N_17144,N_18346);
nor UO_474 (O_474,N_18696,N_18253);
nand UO_475 (O_475,N_17232,N_19237);
nor UO_476 (O_476,N_19434,N_19010);
or UO_477 (O_477,N_19209,N_16958);
xor UO_478 (O_478,N_17523,N_18701);
nor UO_479 (O_479,N_18369,N_18321);
nand UO_480 (O_480,N_17841,N_16097);
and UO_481 (O_481,N_19719,N_19814);
or UO_482 (O_482,N_19462,N_17480);
or UO_483 (O_483,N_16133,N_19442);
nand UO_484 (O_484,N_17723,N_19468);
and UO_485 (O_485,N_16954,N_19517);
nand UO_486 (O_486,N_17440,N_16579);
or UO_487 (O_487,N_19225,N_16998);
xor UO_488 (O_488,N_19992,N_16563);
and UO_489 (O_489,N_18093,N_18880);
nand UO_490 (O_490,N_17066,N_18095);
xor UO_491 (O_491,N_18994,N_16286);
or UO_492 (O_492,N_19559,N_17055);
nor UO_493 (O_493,N_18464,N_18116);
and UO_494 (O_494,N_17982,N_16746);
nand UO_495 (O_495,N_18419,N_18468);
or UO_496 (O_496,N_18004,N_17839);
xor UO_497 (O_497,N_18222,N_18613);
or UO_498 (O_498,N_17072,N_17153);
and UO_499 (O_499,N_16583,N_18471);
or UO_500 (O_500,N_16424,N_17905);
and UO_501 (O_501,N_16915,N_16800);
nor UO_502 (O_502,N_17562,N_17950);
and UO_503 (O_503,N_18897,N_17403);
and UO_504 (O_504,N_18626,N_18797);
nor UO_505 (O_505,N_17421,N_18874);
and UO_506 (O_506,N_19631,N_16247);
nand UO_507 (O_507,N_18678,N_18340);
or UO_508 (O_508,N_18819,N_18996);
nor UO_509 (O_509,N_16055,N_16390);
and UO_510 (O_510,N_19241,N_18060);
and UO_511 (O_511,N_17215,N_18252);
xnor UO_512 (O_512,N_17263,N_17755);
and UO_513 (O_513,N_19269,N_17813);
nor UO_514 (O_514,N_18906,N_18438);
nor UO_515 (O_515,N_17423,N_17732);
and UO_516 (O_516,N_17505,N_19399);
and UO_517 (O_517,N_16310,N_17971);
and UO_518 (O_518,N_19199,N_16019);
or UO_519 (O_519,N_18240,N_19826);
nor UO_520 (O_520,N_19454,N_18210);
xor UO_521 (O_521,N_18835,N_19821);
nand UO_522 (O_522,N_17667,N_18736);
or UO_523 (O_523,N_17273,N_18894);
nor UO_524 (O_524,N_19210,N_18618);
nand UO_525 (O_525,N_16023,N_19638);
or UO_526 (O_526,N_17305,N_18546);
nand UO_527 (O_527,N_16011,N_18376);
and UO_528 (O_528,N_16271,N_16945);
xnor UO_529 (O_529,N_18443,N_16093);
nor UO_530 (O_530,N_19473,N_19649);
nand UO_531 (O_531,N_18875,N_19946);
or UO_532 (O_532,N_19002,N_17495);
nand UO_533 (O_533,N_17125,N_18542);
xor UO_534 (O_534,N_18781,N_16616);
or UO_535 (O_535,N_18607,N_17795);
and UO_536 (O_536,N_19115,N_17443);
and UO_537 (O_537,N_17538,N_17102);
or UO_538 (O_538,N_17593,N_17543);
or UO_539 (O_539,N_16757,N_17150);
xor UO_540 (O_540,N_16508,N_17236);
or UO_541 (O_541,N_18201,N_16253);
nand UO_542 (O_542,N_18843,N_16208);
nor UO_543 (O_543,N_17512,N_16276);
nand UO_544 (O_544,N_16852,N_16478);
nor UO_545 (O_545,N_16623,N_16206);
and UO_546 (O_546,N_16753,N_16219);
and UO_547 (O_547,N_18526,N_18713);
nor UO_548 (O_548,N_16718,N_17508);
or UO_549 (O_549,N_19034,N_18689);
nand UO_550 (O_550,N_18256,N_19009);
nor UO_551 (O_551,N_19091,N_18260);
or UO_552 (O_552,N_18406,N_19403);
nor UO_553 (O_553,N_18265,N_16887);
xnor UO_554 (O_554,N_17407,N_19771);
and UO_555 (O_555,N_19919,N_16320);
or UO_556 (O_556,N_16060,N_17608);
nor UO_557 (O_557,N_16094,N_16448);
xor UO_558 (O_558,N_18317,N_17051);
or UO_559 (O_559,N_16496,N_18910);
xor UO_560 (O_560,N_16056,N_17729);
xor UO_561 (O_561,N_16008,N_17623);
nand UO_562 (O_562,N_19429,N_18782);
nor UO_563 (O_563,N_19030,N_18883);
nor UO_564 (O_564,N_16051,N_17906);
and UO_565 (O_565,N_17584,N_19375);
nor UO_566 (O_566,N_18332,N_16264);
nor UO_567 (O_567,N_19738,N_16221);
nand UO_568 (O_568,N_17275,N_17736);
xnor UO_569 (O_569,N_19614,N_16610);
nor UO_570 (O_570,N_18545,N_18458);
nand UO_571 (O_571,N_17656,N_19044);
and UO_572 (O_572,N_18250,N_18761);
nor UO_573 (O_573,N_18935,N_18869);
nor UO_574 (O_574,N_17445,N_19122);
or UO_575 (O_575,N_19801,N_18274);
or UO_576 (O_576,N_18361,N_16823);
or UO_577 (O_577,N_17124,N_19511);
or UO_578 (O_578,N_16725,N_17424);
nor UO_579 (O_579,N_18836,N_17477);
nor UO_580 (O_580,N_19644,N_18640);
xor UO_581 (O_581,N_17323,N_19292);
and UO_582 (O_582,N_16875,N_19562);
and UO_583 (O_583,N_17768,N_18865);
nand UO_584 (O_584,N_17118,N_18834);
and UO_585 (O_585,N_18026,N_17343);
or UO_586 (O_586,N_16284,N_18925);
and UO_587 (O_587,N_19072,N_17425);
nand UO_588 (O_588,N_19711,N_16189);
nor UO_589 (O_589,N_19672,N_18905);
and UO_590 (O_590,N_19586,N_19339);
nand UO_591 (O_591,N_19890,N_18581);
xor UO_592 (O_592,N_17117,N_16443);
and UO_593 (O_593,N_17643,N_19623);
nor UO_594 (O_594,N_19749,N_17280);
nand UO_595 (O_595,N_16708,N_17369);
nand UO_596 (O_596,N_18352,N_17073);
or UO_597 (O_597,N_17165,N_17180);
or UO_598 (O_598,N_19250,N_16857);
and UO_599 (O_599,N_17856,N_18557);
nor UO_600 (O_600,N_18234,N_16362);
nor UO_601 (O_601,N_19833,N_18312);
nor UO_602 (O_602,N_16205,N_17340);
or UO_603 (O_603,N_18969,N_18722);
xnor UO_604 (O_604,N_19239,N_16526);
and UO_605 (O_605,N_17943,N_18998);
and UO_606 (O_606,N_16721,N_17114);
nor UO_607 (O_607,N_16308,N_17601);
nor UO_608 (O_608,N_17387,N_17826);
nand UO_609 (O_609,N_17233,N_17048);
or UO_610 (O_610,N_16774,N_19428);
xnor UO_611 (O_611,N_19531,N_18928);
nor UO_612 (O_612,N_18635,N_17378);
and UO_613 (O_613,N_18048,N_19571);
xor UO_614 (O_614,N_17392,N_19405);
and UO_615 (O_615,N_16259,N_19798);
nor UO_616 (O_616,N_19285,N_18398);
xnor UO_617 (O_617,N_19110,N_16820);
nor UO_618 (O_618,N_18537,N_16821);
nand UO_619 (O_619,N_19574,N_18268);
xor UO_620 (O_620,N_17984,N_17198);
and UO_621 (O_621,N_16848,N_18759);
nor UO_622 (O_622,N_18074,N_17035);
or UO_623 (O_623,N_18942,N_18380);
nand UO_624 (O_624,N_17130,N_18440);
or UO_625 (O_625,N_18363,N_16519);
or UO_626 (O_626,N_18737,N_19193);
nor UO_627 (O_627,N_18658,N_16992);
or UO_628 (O_628,N_16847,N_16704);
xnor UO_629 (O_629,N_18183,N_19501);
nand UO_630 (O_630,N_16938,N_17214);
nand UO_631 (O_631,N_17999,N_17205);
and UO_632 (O_632,N_19791,N_19679);
nand UO_633 (O_633,N_19244,N_19773);
and UO_634 (O_634,N_18484,N_19971);
or UO_635 (O_635,N_17241,N_18936);
nor UO_636 (O_636,N_19234,N_17809);
nor UO_637 (O_637,N_19541,N_17560);
and UO_638 (O_638,N_16604,N_18450);
nand UO_639 (O_639,N_19521,N_18122);
nand UO_640 (O_640,N_17278,N_16392);
nand UO_641 (O_641,N_19098,N_17089);
and UO_642 (O_642,N_16651,N_16729);
nand UO_643 (O_643,N_17558,N_19374);
or UO_644 (O_644,N_17347,N_16799);
and UO_645 (O_645,N_16190,N_19580);
nand UO_646 (O_646,N_19483,N_19012);
or UO_647 (O_647,N_17769,N_19996);
nand UO_648 (O_648,N_19852,N_17158);
nand UO_649 (O_649,N_18747,N_18573);
and UO_650 (O_650,N_16925,N_16469);
nor UO_651 (O_651,N_19691,N_17713);
and UO_652 (O_652,N_19315,N_16067);
and UO_653 (O_653,N_16355,N_19379);
nor UO_654 (O_654,N_18926,N_19735);
or UO_655 (O_655,N_16353,N_18832);
xnor UO_656 (O_656,N_18432,N_16491);
xor UO_657 (O_657,N_19227,N_18685);
nand UO_658 (O_658,N_16968,N_18255);
nor UO_659 (O_659,N_19160,N_17285);
and UO_660 (O_660,N_16941,N_18258);
xor UO_661 (O_661,N_16622,N_16214);
xor UO_662 (O_662,N_17607,N_17751);
xor UO_663 (O_663,N_17337,N_17003);
or UO_664 (O_664,N_18591,N_16113);
nand UO_665 (O_665,N_17907,N_19560);
and UO_666 (O_666,N_17216,N_17184);
and UO_667 (O_667,N_16470,N_18485);
and UO_668 (O_668,N_17019,N_16201);
nor UO_669 (O_669,N_16300,N_17393);
and UO_670 (O_670,N_18719,N_16665);
or UO_671 (O_671,N_17448,N_18435);
nand UO_672 (O_672,N_18496,N_18779);
xnor UO_673 (O_673,N_17515,N_17962);
and UO_674 (O_674,N_16678,N_19878);
nand UO_675 (O_675,N_16910,N_16173);
and UO_676 (O_676,N_18578,N_18864);
and UO_677 (O_677,N_18548,N_17854);
nand UO_678 (O_678,N_17402,N_17269);
or UO_679 (O_679,N_16903,N_19829);
and UO_680 (O_680,N_16543,N_16463);
or UO_681 (O_681,N_17616,N_16408);
and UO_682 (O_682,N_17959,N_18927);
nand UO_683 (O_683,N_19824,N_18911);
nor UO_684 (O_684,N_16580,N_18669);
nor UO_685 (O_685,N_16139,N_19688);
nand UO_686 (O_686,N_19124,N_16928);
nor UO_687 (O_687,N_18813,N_17923);
nor UO_688 (O_688,N_18961,N_18392);
or UO_689 (O_689,N_17719,N_17013);
nor UO_690 (O_690,N_16688,N_17867);
nand UO_691 (O_691,N_18717,N_16679);
xor UO_692 (O_692,N_19283,N_17485);
nand UO_693 (O_693,N_18749,N_17912);
and UO_694 (O_694,N_18242,N_19280);
and UO_695 (O_695,N_16135,N_16541);
or UO_696 (O_696,N_18439,N_16742);
xor UO_697 (O_697,N_18731,N_16666);
and UO_698 (O_698,N_18129,N_17415);
and UO_699 (O_699,N_18330,N_16379);
and UO_700 (O_700,N_19935,N_19290);
and UO_701 (O_701,N_19819,N_17772);
nand UO_702 (O_702,N_16516,N_19215);
and UO_703 (O_703,N_16983,N_17811);
and UO_704 (O_704,N_17010,N_16366);
nand UO_705 (O_705,N_16658,N_17519);
and UO_706 (O_706,N_17436,N_16464);
nand UO_707 (O_707,N_17083,N_18901);
or UO_708 (O_708,N_19908,N_16050);
or UO_709 (O_709,N_19544,N_19543);
or UO_710 (O_710,N_18055,N_16833);
and UO_711 (O_711,N_17426,N_17176);
and UO_712 (O_712,N_19119,N_16418);
nand UO_713 (O_713,N_19479,N_19358);
and UO_714 (O_714,N_17722,N_19758);
nand UO_715 (O_715,N_16962,N_17002);
nand UO_716 (O_716,N_18047,N_17588);
or UO_717 (O_717,N_17356,N_19506);
nor UO_718 (O_718,N_18087,N_19668);
and UO_719 (O_719,N_17945,N_19645);
or UO_720 (O_720,N_19254,N_16017);
and UO_721 (O_721,N_17592,N_18409);
nand UO_722 (O_722,N_17609,N_16770);
and UO_723 (O_723,N_18326,N_19804);
nand UO_724 (O_724,N_16988,N_17949);
and UO_725 (O_725,N_17394,N_16569);
or UO_726 (O_726,N_18849,N_18786);
nand UO_727 (O_727,N_18670,N_19396);
nor UO_728 (O_728,N_19038,N_16034);
or UO_729 (O_729,N_19477,N_17529);
and UO_730 (O_730,N_16760,N_17513);
nand UO_731 (O_731,N_19650,N_19904);
nor UO_732 (O_732,N_19445,N_19300);
or UO_733 (O_733,N_16981,N_16831);
xnor UO_734 (O_734,N_16068,N_19969);
nand UO_735 (O_735,N_18725,N_19808);
or UO_736 (O_736,N_17272,N_19173);
or UO_737 (O_737,N_18540,N_19880);
or UO_738 (O_738,N_19575,N_18711);
nand UO_739 (O_739,N_16860,N_16455);
and UO_740 (O_740,N_19957,N_19226);
or UO_741 (O_741,N_18311,N_16342);
and UO_742 (O_742,N_17277,N_17625);
nor UO_743 (O_743,N_18308,N_19212);
or UO_744 (O_744,N_17684,N_18625);
or UO_745 (O_745,N_16227,N_19305);
and UO_746 (O_746,N_16511,N_17104);
or UO_747 (O_747,N_18947,N_16949);
nand UO_748 (O_748,N_18795,N_18076);
xnor UO_749 (O_749,N_17937,N_16562);
nor UO_750 (O_750,N_16045,N_18178);
nor UO_751 (O_751,N_16672,N_19296);
and UO_752 (O_752,N_19029,N_17235);
nand UO_753 (O_753,N_17226,N_16217);
nor UO_754 (O_754,N_18628,N_19799);
xnor UO_755 (O_755,N_17499,N_16786);
nor UO_756 (O_756,N_19390,N_17113);
nor UO_757 (O_757,N_18842,N_16814);
and UO_758 (O_758,N_19247,N_17348);
nand UO_759 (O_759,N_16846,N_19340);
nor UO_760 (O_760,N_19456,N_18861);
xnor UO_761 (O_761,N_18313,N_18422);
xor UO_762 (O_762,N_18291,N_19102);
xor UO_763 (O_763,N_17404,N_18881);
nand UO_764 (O_764,N_19906,N_18354);
nand UO_765 (O_765,N_19599,N_19348);
nor UO_766 (O_766,N_19825,N_16111);
xor UO_767 (O_767,N_17397,N_16293);
nor UO_768 (O_768,N_18327,N_19211);
nand UO_769 (O_769,N_19884,N_19410);
nor UO_770 (O_770,N_16375,N_18003);
or UO_771 (O_771,N_19080,N_16620);
xor UO_772 (O_772,N_17553,N_19914);
nand UO_773 (O_773,N_18886,N_17455);
or UO_774 (O_774,N_16939,N_17915);
nor UO_775 (O_775,N_19872,N_18079);
or UO_776 (O_776,N_19740,N_17720);
nor UO_777 (O_777,N_18611,N_19750);
or UO_778 (O_778,N_17831,N_16009);
or UO_779 (O_779,N_19139,N_19561);
or UO_780 (O_780,N_17534,N_18831);
or UO_781 (O_781,N_17696,N_19855);
and UO_782 (O_782,N_18039,N_19041);
or UO_783 (O_783,N_16445,N_17627);
nand UO_784 (O_784,N_16497,N_19219);
and UO_785 (O_785,N_17265,N_17712);
and UO_786 (O_786,N_19395,N_18992);
nand UO_787 (O_787,N_18774,N_19360);
nand UO_788 (O_788,N_19721,N_17227);
and UO_789 (O_789,N_17242,N_17873);
and UO_790 (O_790,N_18608,N_17116);
or UO_791 (O_791,N_16384,N_19709);
nand UO_792 (O_792,N_17998,N_16957);
nor UO_793 (O_793,N_19831,N_18592);
and UO_794 (O_794,N_19268,N_18314);
nand UO_795 (O_795,N_18553,N_16595);
nor UO_796 (O_796,N_17368,N_16213);
nor UO_797 (O_797,N_18489,N_16900);
and UO_798 (O_798,N_17088,N_17868);
nor UO_799 (O_799,N_18507,N_17091);
nor UO_800 (O_800,N_18445,N_17993);
or UO_801 (O_801,N_17706,N_16291);
nand UO_802 (O_802,N_19221,N_17230);
or UO_803 (O_803,N_19944,N_19014);
xnor UO_804 (O_804,N_19564,N_17218);
or UO_805 (O_805,N_18976,N_18929);
or UO_806 (O_806,N_17925,N_17385);
or UO_807 (O_807,N_18575,N_18105);
nand UO_808 (O_808,N_16199,N_19177);
or UO_809 (O_809,N_19279,N_19747);
or UO_810 (O_810,N_19079,N_18018);
nor UO_811 (O_811,N_19500,N_19433);
nand UO_812 (O_812,N_17844,N_18784);
nor UO_813 (O_813,N_17614,N_17883);
nand UO_814 (O_814,N_19587,N_18436);
or UO_815 (O_815,N_17632,N_19457);
or UO_816 (O_816,N_16130,N_17542);
nand UO_817 (O_817,N_17972,N_16627);
or UO_818 (O_818,N_18760,N_19854);
nor UO_819 (O_819,N_18128,N_17852);
or UO_820 (O_820,N_18467,N_19176);
nand UO_821 (O_821,N_16458,N_17703);
and UO_822 (O_822,N_17602,N_16172);
nor UO_823 (O_823,N_18671,N_18078);
and UO_824 (O_824,N_19194,N_17427);
and UO_825 (O_825,N_19949,N_18194);
nor UO_826 (O_826,N_17029,N_16372);
and UO_827 (O_827,N_16409,N_17639);
nor UO_828 (O_828,N_18197,N_16489);
nand UO_829 (O_829,N_19970,N_16621);
xnor UO_830 (O_830,N_19497,N_19775);
or UO_831 (O_831,N_17098,N_16480);
nand UO_832 (O_832,N_19535,N_16946);
and UO_833 (O_833,N_19810,N_18475);
nand UO_834 (O_834,N_19015,N_17823);
or UO_835 (O_835,N_19461,N_19533);
or UO_836 (O_836,N_19514,N_16184);
and UO_837 (O_837,N_17974,N_19858);
nor UO_838 (O_838,N_17457,N_16295);
and UO_839 (O_839,N_17299,N_16490);
or UO_840 (O_840,N_18297,N_17700);
or UO_841 (O_841,N_16856,N_16102);
nand UO_842 (O_842,N_16802,N_16481);
nand UO_843 (O_843,N_19526,N_17688);
nand UO_844 (O_844,N_19430,N_18615);
xor UO_845 (O_845,N_18166,N_16809);
nand UO_846 (O_846,N_17189,N_19891);
nor UO_847 (O_847,N_16844,N_19178);
or UO_848 (O_848,N_17367,N_16749);
or UO_849 (O_849,N_17522,N_16345);
and UO_850 (O_850,N_16895,N_19795);
nor UO_851 (O_851,N_19632,N_17770);
and UO_852 (O_852,N_16505,N_17162);
and UO_853 (O_853,N_18099,N_16539);
and UO_854 (O_854,N_16525,N_17122);
and UO_855 (O_855,N_17967,N_19001);
or UO_856 (O_856,N_19367,N_16545);
xor UO_857 (O_857,N_17590,N_16498);
nand UO_858 (O_858,N_17338,N_16065);
nand UO_859 (O_859,N_17200,N_16183);
nand UO_860 (O_860,N_18814,N_19724);
nand UO_861 (O_861,N_17250,N_17641);
nor UO_862 (O_862,N_19667,N_18900);
nor UO_863 (O_863,N_19678,N_16835);
xor UO_864 (O_864,N_17022,N_19203);
nor UO_865 (O_865,N_19085,N_19843);
nand UO_866 (O_866,N_17502,N_16210);
nor UO_867 (O_867,N_17710,N_16748);
nand UO_868 (O_868,N_18599,N_18302);
and UO_869 (O_869,N_17650,N_17049);
or UO_870 (O_870,N_17842,N_18219);
or UO_871 (O_871,N_18638,N_19313);
nand UO_872 (O_872,N_19299,N_17884);
or UO_873 (O_873,N_17363,N_19731);
and UO_874 (O_874,N_18453,N_19888);
nand UO_875 (O_875,N_18967,N_18447);
xor UO_876 (O_876,N_18972,N_18388);
and UO_877 (O_877,N_18469,N_19555);
nor UO_878 (O_878,N_19654,N_19974);
and UO_879 (O_879,N_17953,N_18431);
and UO_880 (O_880,N_19472,N_16231);
and UO_881 (O_881,N_17302,N_17896);
or UO_882 (O_882,N_16817,N_17767);
and UO_883 (O_883,N_19214,N_19467);
nand UO_884 (O_884,N_19736,N_19466);
nor UO_885 (O_885,N_18741,N_17396);
nand UO_886 (O_886,N_16309,N_18682);
nand UO_887 (O_887,N_16059,N_16152);
and UO_888 (O_888,N_19264,N_19475);
or UO_889 (O_889,N_17785,N_18877);
nor UO_890 (O_890,N_19333,N_18254);
and UO_891 (O_891,N_16795,N_16403);
nand UO_892 (O_892,N_18147,N_19984);
or UO_893 (O_893,N_18534,N_19081);
and UO_894 (O_894,N_16120,N_19198);
nor UO_895 (O_895,N_19071,N_18261);
xnor UO_896 (O_896,N_18430,N_16237);
nor UO_897 (O_897,N_18892,N_17539);
nor UO_898 (O_898,N_19807,N_19622);
and UO_899 (O_899,N_16585,N_19147);
nor UO_900 (O_900,N_19998,N_19143);
and UO_901 (O_901,N_17306,N_18509);
or UO_902 (O_902,N_18149,N_16904);
nor UO_903 (O_903,N_19955,N_17605);
nand UO_904 (O_904,N_19573,N_18724);
and UO_905 (O_905,N_18034,N_19394);
or UO_906 (O_906,N_19994,N_18914);
and UO_907 (O_907,N_19912,N_18887);
nor UO_908 (O_908,N_17492,N_17599);
nand UO_909 (O_909,N_19380,N_17916);
nor UO_910 (O_910,N_16960,N_16646);
nor UO_911 (O_911,N_19695,N_18637);
nor UO_912 (O_912,N_16150,N_19837);
and UO_913 (O_913,N_17362,N_19536);
nand UO_914 (O_914,N_16843,N_18322);
or UO_915 (O_915,N_19742,N_17373);
and UO_916 (O_916,N_17379,N_17966);
nor UO_917 (O_917,N_19187,N_18523);
nor UO_918 (O_918,N_17282,N_16436);
xor UO_919 (O_919,N_16365,N_19823);
and UO_920 (O_920,N_16710,N_16148);
xnor UO_921 (O_921,N_19057,N_16279);
nand UO_922 (O_922,N_19676,N_17052);
or UO_923 (O_923,N_18358,N_19757);
xor UO_924 (O_924,N_17359,N_18479);
nor UO_925 (O_925,N_19017,N_19200);
or UO_926 (O_926,N_18062,N_19832);
nand UO_927 (O_927,N_16811,N_16449);
or UO_928 (O_928,N_19059,N_18762);
and UO_929 (O_929,N_17157,N_16499);
and UO_930 (O_930,N_16512,N_17342);
or UO_931 (O_931,N_18042,N_16777);
nand UO_932 (O_932,N_17110,N_17567);
nand UO_933 (O_933,N_16025,N_17503);
or UO_934 (O_934,N_17061,N_17846);
xor UO_935 (O_935,N_17281,N_16923);
or UO_936 (O_936,N_17169,N_16033);
xnor UO_937 (O_937,N_17675,N_18934);
or UO_938 (O_938,N_16572,N_16632);
and UO_939 (O_939,N_18560,N_19594);
nor UO_940 (O_940,N_16592,N_16713);
or UO_941 (O_941,N_18283,N_17435);
nand UO_942 (O_942,N_19420,N_18949);
and UO_943 (O_943,N_16391,N_17279);
nor UO_944 (O_944,N_18173,N_17004);
and UO_945 (O_945,N_16696,N_19849);
and UO_946 (O_946,N_16951,N_17053);
or UO_947 (O_947,N_17518,N_17160);
nand UO_948 (O_948,N_16212,N_16109);
nand UO_949 (O_949,N_19308,N_19070);
nand UO_950 (O_950,N_18888,N_17065);
nor UO_951 (O_951,N_17570,N_17310);
and UO_952 (O_952,N_19838,N_19779);
and UO_953 (O_953,N_16427,N_18656);
and UO_954 (O_954,N_16115,N_19999);
xnor UO_955 (O_955,N_16063,N_17773);
nand UO_956 (O_956,N_19363,N_18415);
nand UO_957 (O_957,N_18629,N_18401);
nand UO_958 (O_958,N_19008,N_16142);
or UO_959 (O_959,N_16338,N_18675);
and UO_960 (O_960,N_17468,N_18344);
xor UO_961 (O_961,N_19249,N_17274);
nor UO_962 (O_962,N_18597,N_18703);
and UO_963 (O_963,N_19835,N_17400);
nand UO_964 (O_964,N_17716,N_17902);
and UO_965 (O_965,N_16413,N_17636);
nand UO_966 (O_966,N_18350,N_19778);
or UO_967 (O_967,N_16827,N_18660);
nand UO_968 (O_968,N_17995,N_17744);
and UO_969 (O_969,N_18476,N_19518);
and UO_970 (O_970,N_19223,N_19304);
nand UO_971 (O_971,N_17332,N_17580);
or UO_972 (O_972,N_17961,N_19685);
and UO_973 (O_973,N_18619,N_16224);
and UO_974 (O_974,N_16327,N_19192);
or UO_975 (O_975,N_18985,N_17541);
xor UO_976 (O_976,N_17417,N_16167);
xnor UO_977 (O_977,N_18576,N_16529);
nand UO_978 (O_978,N_18177,N_19554);
and UO_979 (O_979,N_19298,N_18536);
nand UO_980 (O_980,N_19664,N_18753);
and UO_981 (O_981,N_17837,N_17527);
nand UO_982 (O_982,N_18851,N_19397);
nor UO_983 (O_983,N_18846,N_18200);
nand UO_984 (O_984,N_18850,N_17576);
and UO_985 (O_985,N_16577,N_19671);
nor UO_986 (O_986,N_18579,N_16451);
nor UO_987 (O_987,N_18554,N_19082);
nand UO_988 (O_988,N_19659,N_18785);
or UO_989 (O_989,N_18100,N_18567);
nor UO_990 (O_990,N_19604,N_16164);
and UO_991 (O_991,N_19687,N_17936);
nand UO_992 (O_992,N_17640,N_17996);
nand UO_993 (O_993,N_19550,N_18552);
xor UO_994 (O_994,N_16438,N_18120);
nor UO_995 (O_995,N_16796,N_16862);
xnor UO_996 (O_996,N_18172,N_18217);
and UO_997 (O_997,N_19218,N_19818);
nand UO_998 (O_998,N_16724,N_17262);
and UO_999 (O_999,N_19496,N_17497);
nand UO_1000 (O_1000,N_16081,N_19945);
nor UO_1001 (O_1001,N_17645,N_16884);
or UO_1002 (O_1002,N_19963,N_16069);
nor UO_1003 (O_1003,N_16791,N_16940);
or UO_1004 (O_1004,N_18135,N_19100);
nand UO_1005 (O_1005,N_19953,N_18966);
nand UO_1006 (O_1006,N_18032,N_16502);
and UO_1007 (O_1007,N_16318,N_16664);
or UO_1008 (O_1008,N_18556,N_19609);
and UO_1009 (O_1009,N_16229,N_17249);
nor UO_1010 (O_1010,N_16179,N_19393);
or UO_1011 (O_1011,N_16918,N_18621);
nor UO_1012 (O_1012,N_19591,N_19341);
or UO_1013 (O_1013,N_16901,N_17644);
and UO_1014 (O_1014,N_18366,N_16166);
nand UO_1015 (O_1015,N_18908,N_17948);
nor UO_1016 (O_1016,N_16412,N_17411);
nand UO_1017 (O_1017,N_16690,N_17123);
and UO_1018 (O_1018,N_18500,N_16466);
or UO_1019 (O_1019,N_18044,N_17794);
or UO_1020 (O_1020,N_18950,N_18639);
nand UO_1021 (O_1021,N_18492,N_18793);
or UO_1022 (O_1022,N_16000,N_18359);
nor UO_1023 (O_1023,N_17805,N_16107);
nand UO_1024 (O_1024,N_18182,N_18245);
or UO_1025 (O_1025,N_17910,N_19031);
nand UO_1026 (O_1026,N_17223,N_17095);
and UO_1027 (O_1027,N_16126,N_16380);
and UO_1028 (O_1028,N_16568,N_17112);
or UO_1029 (O_1029,N_19675,N_17546);
or UO_1030 (O_1030,N_16657,N_17994);
xor UO_1031 (O_1031,N_17060,N_17212);
nor UO_1032 (O_1032,N_17806,N_19370);
or UO_1033 (O_1033,N_19484,N_16405);
nand UO_1034 (O_1034,N_17658,N_18662);
nand UO_1035 (O_1035,N_17231,N_16950);
nor UO_1036 (O_1036,N_19295,N_19288);
nor UO_1037 (O_1037,N_18378,N_18974);
nor UO_1038 (O_1038,N_18416,N_18778);
nand UO_1039 (O_1039,N_16908,N_18627);
nand UO_1040 (O_1040,N_16306,N_18838);
or UO_1041 (O_1041,N_16907,N_19552);
nand UO_1042 (O_1042,N_19063,N_18783);
nor UO_1043 (O_1043,N_17488,N_18858);
nand UO_1044 (O_1044,N_17410,N_17070);
nor UO_1045 (O_1045,N_19235,N_16504);
xor UO_1046 (O_1046,N_18990,N_16235);
nor UO_1047 (O_1047,N_17012,N_18549);
nand UO_1048 (O_1048,N_17018,N_17080);
nor UO_1049 (O_1049,N_16608,N_18477);
and UO_1050 (O_1050,N_16768,N_16161);
xor UO_1051 (O_1051,N_16528,N_18057);
or UO_1052 (O_1052,N_18944,N_18986);
and UO_1053 (O_1053,N_17978,N_19674);
and UO_1054 (O_1054,N_16441,N_19032);
and UO_1055 (O_1055,N_17676,N_18483);
nor UO_1056 (O_1056,N_16825,N_17857);
and UO_1057 (O_1057,N_17611,N_16536);
nor UO_1058 (O_1058,N_16268,N_18367);
or UO_1059 (O_1059,N_19961,N_17201);
xor UO_1060 (O_1060,N_16242,N_18125);
or UO_1061 (O_1061,N_18889,N_18891);
nor UO_1062 (O_1062,N_19449,N_16312);
nand UO_1063 (O_1063,N_19788,N_16394);
and UO_1064 (O_1064,N_19979,N_17412);
or UO_1065 (O_1065,N_19745,N_16255);
or UO_1066 (O_1066,N_17473,N_18587);
nand UO_1067 (O_1067,N_19639,N_19495);
and UO_1068 (O_1068,N_16030,N_17093);
nor UO_1069 (O_1069,N_16912,N_19028);
or UO_1070 (O_1070,N_18098,N_18641);
or UO_1071 (O_1071,N_17536,N_16574);
and UO_1072 (O_1072,N_17006,N_18410);
nor UO_1073 (O_1073,N_17900,N_16683);
or UO_1074 (O_1074,N_17401,N_16609);
nand UO_1075 (O_1075,N_17163,N_18855);
or UO_1076 (O_1076,N_19359,N_18150);
and UO_1077 (O_1077,N_18924,N_19640);
nor UO_1078 (O_1078,N_16518,N_19371);
or UO_1079 (O_1079,N_18238,N_18251);
and UO_1080 (O_1080,N_18916,N_17591);
xnor UO_1081 (O_1081,N_18757,N_19236);
nand UO_1082 (O_1082,N_17434,N_17339);
xor UO_1083 (O_1083,N_16450,N_18952);
or UO_1084 (O_1084,N_19302,N_19794);
nand UO_1085 (O_1085,N_16273,N_16961);
nor UO_1086 (O_1086,N_19990,N_16741);
nand UO_1087 (O_1087,N_19144,N_18472);
or UO_1088 (O_1088,N_18052,N_19850);
or UO_1089 (O_1089,N_16576,N_18024);
nand UO_1090 (O_1090,N_18964,N_16080);
nor UO_1091 (O_1091,N_16728,N_17484);
or UO_1092 (O_1092,N_19568,N_19106);
nand UO_1093 (O_1093,N_18403,N_16705);
nor UO_1094 (O_1094,N_17481,N_19238);
xnor UO_1095 (O_1095,N_19101,N_18586);
nor UO_1096 (O_1096,N_18885,N_18063);
nor UO_1097 (O_1097,N_18681,N_16993);
nor UO_1098 (O_1098,N_16263,N_18290);
or UO_1099 (O_1099,N_16629,N_16626);
nand UO_1100 (O_1100,N_18386,N_17725);
or UO_1101 (O_1101,N_16756,N_18743);
nor UO_1102 (O_1102,N_17932,N_18333);
nor UO_1103 (O_1103,N_16758,N_19681);
and UO_1104 (O_1104,N_19216,N_19603);
or UO_1105 (O_1105,N_19648,N_19338);
nor UO_1106 (O_1106,N_19291,N_18803);
or UO_1107 (O_1107,N_19401,N_18919);
or UO_1108 (O_1108,N_19025,N_17571);
nand UO_1109 (O_1109,N_17406,N_16254);
nor UO_1110 (O_1110,N_16322,N_16307);
and UO_1111 (O_1111,N_17801,N_17033);
and UO_1112 (O_1112,N_16160,N_16487);
nand UO_1113 (O_1113,N_18066,N_17380);
xnor UO_1114 (O_1114,N_17824,N_18879);
and UO_1115 (O_1115,N_19307,N_16002);
nand UO_1116 (O_1116,N_19777,N_17516);
nor UO_1117 (O_1117,N_19805,N_18729);
nand UO_1118 (O_1118,N_19572,N_17960);
xor UO_1119 (O_1119,N_19846,N_18239);
nor UO_1120 (O_1120,N_19096,N_19419);
and UO_1121 (O_1121,N_16735,N_16560);
xnor UO_1122 (O_1122,N_18535,N_16612);
xor UO_1123 (O_1123,N_18574,N_18853);
nor UO_1124 (O_1124,N_17843,N_17044);
nand UO_1125 (O_1125,N_16461,N_16625);
nand UO_1126 (O_1126,N_17320,N_19402);
nor UO_1127 (O_1127,N_19148,N_17860);
xnor UO_1128 (O_1128,N_19796,N_19075);
or UO_1129 (O_1129,N_19723,N_17847);
and UO_1130 (O_1130,N_18132,N_18138);
nor UO_1131 (O_1131,N_17881,N_16246);
nor UO_1132 (O_1132,N_18230,N_18562);
nand UO_1133 (O_1133,N_17439,N_18630);
nor UO_1134 (O_1134,N_19180,N_18706);
nor UO_1135 (O_1135,N_19131,N_18292);
or UO_1136 (O_1136,N_18202,N_19155);
nand UO_1137 (O_1137,N_19328,N_17204);
or UO_1138 (O_1138,N_17493,N_18732);
or UO_1139 (O_1139,N_17254,N_16108);
nand UO_1140 (O_1140,N_17822,N_19789);
xor UO_1141 (O_1141,N_19813,N_17781);
xnor UO_1142 (O_1142,N_18822,N_19343);
xnor UO_1143 (O_1143,N_18646,N_16882);
nand UO_1144 (O_1144,N_19708,N_16265);
and UO_1145 (O_1145,N_16706,N_18644);
or UO_1146 (O_1146,N_19240,N_19137);
nand UO_1147 (O_1147,N_19932,N_16144);
nor UO_1148 (O_1148,N_17565,N_16083);
or UO_1149 (O_1149,N_18596,N_16527);
nand UO_1150 (O_1150,N_18516,N_19959);
and UO_1151 (O_1151,N_16540,N_18984);
and UO_1152 (O_1152,N_16401,N_18859);
nor UO_1153 (O_1153,N_17229,N_19074);
and UO_1154 (O_1154,N_19761,N_16149);
xor UO_1155 (O_1155,N_19765,N_16764);
nand UO_1156 (O_1156,N_18805,N_16077);
or UO_1157 (O_1157,N_18580,N_17920);
nor UO_1158 (O_1158,N_19812,N_16369);
nand UO_1159 (O_1159,N_19873,N_18584);
or UO_1160 (O_1160,N_19229,N_18720);
and UO_1161 (O_1161,N_16896,N_18267);
nor UO_1162 (O_1162,N_16779,N_19094);
nand UO_1163 (O_1163,N_16236,N_18131);
or UO_1164 (O_1164,N_18746,N_18355);
and UO_1165 (O_1165,N_18412,N_17312);
nor UO_1166 (O_1166,N_17199,N_17140);
or UO_1167 (O_1167,N_17243,N_17292);
nand UO_1168 (O_1168,N_19376,N_18946);
xor UO_1169 (O_1169,N_19877,N_18123);
or UO_1170 (O_1170,N_19424,N_18697);
xnor UO_1171 (O_1171,N_17689,N_16978);
or UO_1172 (O_1172,N_19326,N_16542);
and UO_1173 (O_1173,N_19337,N_17665);
and UO_1174 (O_1174,N_18857,N_19231);
and UO_1175 (O_1175,N_18296,N_18852);
or UO_1176 (O_1176,N_18821,N_18505);
nand UO_1177 (O_1177,N_16129,N_16044);
and UO_1178 (O_1178,N_19921,N_16738);
xor UO_1179 (O_1179,N_17934,N_19064);
nand UO_1180 (O_1180,N_17461,N_18187);
and UO_1181 (O_1181,N_17076,N_18266);
nand UO_1182 (O_1182,N_19046,N_16750);
nand UO_1183 (O_1183,N_16761,N_16169);
and UO_1184 (O_1184,N_18563,N_17092);
nand UO_1185 (O_1185,N_19232,N_16838);
nand UO_1186 (O_1186,N_19284,N_18610);
or UO_1187 (O_1187,N_18772,N_16422);
xnor UO_1188 (O_1188,N_19940,N_16054);
and UO_1189 (O_1189,N_16535,N_16509);
and UO_1190 (O_1190,N_16871,N_18962);
nor UO_1191 (O_1191,N_19459,N_19896);
nand UO_1192 (O_1192,N_16336,N_18411);
xnor UO_1193 (O_1193,N_17628,N_17816);
nand UO_1194 (O_1194,N_16209,N_17750);
nand UO_1195 (O_1195,N_18965,N_17898);
nand UO_1196 (O_1196,N_16180,N_16084);
nand UO_1197 (O_1197,N_17182,N_18953);
and UO_1198 (O_1198,N_19700,N_16588);
or UO_1199 (O_1199,N_19111,N_19516);
nor UO_1200 (O_1200,N_18480,N_18829);
nor UO_1201 (O_1201,N_17001,N_17939);
nor UO_1202 (O_1202,N_18884,N_19634);
nand UO_1203 (O_1203,N_16038,N_19925);
nand UO_1204 (O_1204,N_17371,N_18841);
xor UO_1205 (O_1205,N_16302,N_19486);
or UO_1206 (O_1206,N_19728,N_17704);
and UO_1207 (O_1207,N_19195,N_18395);
nand UO_1208 (O_1208,N_17914,N_16428);
nor UO_1209 (O_1209,N_18941,N_19318);
or UO_1210 (O_1210,N_17662,N_17414);
or UO_1211 (O_1211,N_19578,N_17501);
nor UO_1212 (O_1212,N_16685,N_16955);
nand UO_1213 (O_1213,N_19625,N_18634);
or UO_1214 (O_1214,N_19112,N_18566);
nand UO_1215 (O_1215,N_18360,N_19109);
or UO_1216 (O_1216,N_16321,N_19508);
and UO_1217 (O_1217,N_19004,N_18752);
nor UO_1218 (O_1218,N_19722,N_17786);
or UO_1219 (O_1219,N_19182,N_19158);
and UO_1220 (O_1220,N_17829,N_17428);
and UO_1221 (O_1221,N_17357,N_18995);
and UO_1222 (O_1222,N_18651,N_18668);
or UO_1223 (O_1223,N_18828,N_16343);
nand UO_1224 (O_1224,N_19993,N_17600);
and UO_1225 (O_1225,N_19007,N_19763);
nand UO_1226 (O_1226,N_16772,N_17454);
xor UO_1227 (O_1227,N_16297,N_17366);
nand UO_1228 (O_1228,N_16694,N_18820);
nand UO_1229 (O_1229,N_16522,N_18666);
nand UO_1230 (O_1230,N_17682,N_16095);
nand UO_1231 (O_1231,N_16334,N_16476);
xor UO_1232 (O_1232,N_19217,N_16162);
and UO_1233 (O_1233,N_17669,N_17086);
nor UO_1234 (O_1234,N_16855,N_19929);
nand UO_1235 (O_1235,N_17737,N_19966);
and UO_1236 (O_1236,N_16557,N_18659);
nor UO_1237 (O_1237,N_19170,N_16740);
or UO_1238 (O_1238,N_17178,N_16048);
or UO_1239 (O_1239,N_18791,N_19320);
and UO_1240 (O_1240,N_19683,N_17289);
nor UO_1241 (O_1241,N_16202,N_17965);
or UO_1242 (O_1242,N_19903,N_16722);
and UO_1243 (O_1243,N_18382,N_19253);
or UO_1244 (O_1244,N_19188,N_19478);
nand UO_1245 (O_1245,N_18633,N_16304);
or UO_1246 (O_1246,N_18692,N_16778);
and UO_1247 (O_1247,N_18191,N_19764);
and UO_1248 (O_1248,N_16087,N_16073);
and UO_1249 (O_1249,N_16790,N_19690);
nor UO_1250 (O_1250,N_17564,N_17574);
or UO_1251 (O_1251,N_18802,N_19540);
or UO_1252 (O_1252,N_17376,N_18529);
or UO_1253 (O_1253,N_18751,N_17820);
xnor UO_1254 (O_1254,N_16356,N_16062);
nor UO_1255 (O_1255,N_16773,N_18539);
nor UO_1256 (O_1256,N_19161,N_16830);
xnor UO_1257 (O_1257,N_19899,N_19943);
xor UO_1258 (O_1258,N_18577,N_19894);
nor UO_1259 (O_1259,N_17818,N_16671);
nand UO_1260 (O_1260,N_18807,N_17835);
xor UO_1261 (O_1261,N_16924,N_17141);
and UO_1262 (O_1262,N_18823,N_18214);
or UO_1263 (O_1263,N_17577,N_18142);
nand UO_1264 (O_1264,N_18310,N_16116);
or UO_1265 (O_1265,N_16117,N_16667);
nand UO_1266 (O_1266,N_19704,N_17020);
nand UO_1267 (O_1267,N_16611,N_19037);
and UO_1268 (O_1268,N_17904,N_18655);
and UO_1269 (O_1269,N_18913,N_17151);
xor UO_1270 (O_1270,N_18810,N_16337);
and UO_1271 (O_1271,N_18343,N_17195);
nor UO_1272 (O_1272,N_16922,N_19947);
and UO_1273 (O_1273,N_17727,N_17761);
and UO_1274 (O_1274,N_17621,N_16980);
or UO_1275 (O_1275,N_18796,N_19103);
nor UO_1276 (O_1276,N_18798,N_16692);
nor UO_1277 (O_1277,N_19499,N_16477);
and UO_1278 (O_1278,N_19345,N_16853);
or UO_1279 (O_1279,N_19748,N_17797);
nor UO_1280 (O_1280,N_18543,N_16106);
or UO_1281 (O_1281,N_16806,N_17408);
nor UO_1282 (O_1282,N_19168,N_16589);
nor UO_1283 (O_1283,N_16442,N_19306);
nor UO_1284 (O_1284,N_16032,N_16460);
or UO_1285 (O_1285,N_19104,N_17365);
or UO_1286 (O_1286,N_16943,N_18491);
and UO_1287 (O_1287,N_18342,N_19352);
or UO_1288 (O_1288,N_18309,N_17372);
nand UO_1289 (O_1289,N_19934,N_17479);
and UO_1290 (O_1290,N_16316,N_17476);
or UO_1291 (O_1291,N_19842,N_18108);
nand UO_1292 (O_1292,N_17202,N_17147);
or UO_1293 (O_1293,N_19175,N_19576);
or UO_1294 (O_1294,N_16417,N_18704);
and UO_1295 (O_1295,N_19928,N_19797);
nand UO_1296 (O_1296,N_16423,N_18226);
xor UO_1297 (O_1297,N_16406,N_19260);
or UO_1298 (O_1298,N_18402,N_19415);
nor UO_1299 (O_1299,N_17874,N_18677);
nand UO_1300 (O_1300,N_19515,N_17743);
nor UO_1301 (O_1301,N_16154,N_19408);
and UO_1302 (O_1302,N_19431,N_18482);
nor UO_1303 (O_1303,N_18728,N_17817);
nor UO_1304 (O_1304,N_16325,N_17780);
and UO_1305 (O_1305,N_18818,N_18699);
nor UO_1306 (O_1306,N_16747,N_18287);
nor UO_1307 (O_1307,N_18179,N_18775);
nor UO_1308 (O_1308,N_16244,N_18133);
xor UO_1309 (O_1309,N_19752,N_18709);
and UO_1310 (O_1310,N_17050,N_16354);
xnor UO_1311 (O_1311,N_16012,N_19529);
nand UO_1312 (O_1312,N_18602,N_17490);
nor UO_1313 (O_1313,N_17659,N_17958);
and UO_1314 (O_1314,N_17133,N_19204);
nand UO_1315 (O_1315,N_18691,N_18195);
and UO_1316 (O_1316,N_16357,N_16719);
nor UO_1317 (O_1317,N_18975,N_16421);
and UO_1318 (O_1318,N_18826,N_18508);
nor UO_1319 (O_1319,N_18945,N_16684);
and UO_1320 (O_1320,N_18293,N_16377);
nand UO_1321 (O_1321,N_19633,N_19905);
and UO_1322 (O_1322,N_16794,N_16407);
or UO_1323 (O_1323,N_16812,N_16331);
nand UO_1324 (O_1324,N_19066,N_17559);
nand UO_1325 (O_1325,N_19897,N_19595);
nand UO_1326 (O_1326,N_19045,N_17926);
nor UO_1327 (O_1327,N_19931,N_18473);
nor UO_1328 (O_1328,N_18673,N_16507);
nand UO_1329 (O_1329,N_17882,N_17303);
and UO_1330 (O_1330,N_19258,N_18278);
or UO_1331 (O_1331,N_17980,N_16828);
nand UO_1332 (O_1332,N_17458,N_17126);
xnor UO_1333 (O_1333,N_18547,N_19350);
nor UO_1334 (O_1334,N_16419,N_17858);
or UO_1335 (O_1335,N_18013,N_16571);
and UO_1336 (O_1336,N_18425,N_17259);
nand UO_1337 (O_1337,N_17286,N_18368);
nor UO_1338 (O_1338,N_19026,N_18357);
nor UO_1339 (O_1339,N_16709,N_16788);
or UO_1340 (O_1340,N_16997,N_16669);
nor UO_1341 (O_1341,N_16717,N_16453);
or UO_1342 (O_1342,N_17464,N_17207);
xor UO_1343 (O_1343,N_16826,N_17524);
or UO_1344 (O_1344,N_18848,N_19325);
and UO_1345 (O_1345,N_18979,N_17810);
or UO_1346 (O_1346,N_19769,N_18301);
nand UO_1347 (O_1347,N_18335,N_16515);
and UO_1348 (O_1348,N_19135,N_17975);
and UO_1349 (O_1349,N_16239,N_18839);
nand UO_1350 (O_1350,N_19381,N_17877);
and UO_1351 (O_1351,N_19523,N_19118);
nand UO_1352 (O_1352,N_18030,N_18263);
nor UO_1353 (O_1353,N_19487,N_16196);
nor UO_1354 (O_1354,N_19309,N_16374);
and UO_1355 (O_1355,N_18957,N_18623);
nand UO_1356 (O_1356,N_16699,N_16006);
or UO_1357 (O_1357,N_16432,N_16096);
xnor UO_1358 (O_1358,N_19257,N_19387);
or UO_1359 (O_1359,N_18223,N_19939);
xnor UO_1360 (O_1360,N_19828,N_18215);
nor UO_1361 (O_1361,N_16999,N_18680);
nand UO_1362 (O_1362,N_16402,N_16933);
xnor UO_1363 (O_1363,N_17161,N_17500);
nand UO_1364 (O_1364,N_19069,N_19332);
and UO_1365 (O_1365,N_16049,N_16815);
nand UO_1366 (O_1366,N_18679,N_18134);
and UO_1367 (O_1367,N_18282,N_16468);
or UO_1368 (O_1368,N_16570,N_17673);
nand UO_1369 (O_1369,N_18373,N_17419);
or UO_1370 (O_1370,N_16010,N_17646);
and UO_1371 (O_1371,N_18487,N_19314);
nand UO_1372 (O_1372,N_19055,N_16663);
nor UO_1373 (O_1373,N_18938,N_18049);
and UO_1374 (O_1374,N_16818,N_17318);
or UO_1375 (O_1375,N_16004,N_17381);
xnor UO_1376 (O_1376,N_18907,N_18723);
or UO_1377 (O_1377,N_17327,N_16919);
or UO_1378 (O_1378,N_16382,N_18356);
nand UO_1379 (O_1379,N_17707,N_16170);
or UO_1380 (O_1380,N_19869,N_16849);
xor UO_1381 (O_1381,N_17977,N_18154);
nor UO_1382 (O_1382,N_17930,N_16137);
nand UO_1383 (O_1383,N_19455,N_19583);
nand UO_1384 (O_1384,N_16399,N_16444);
nand UO_1385 (O_1385,N_18364,N_16916);
nor UO_1386 (O_1386,N_17446,N_16367);
nor UO_1387 (O_1387,N_19121,N_19790);
nor UO_1388 (O_1388,N_16269,N_18956);
and UO_1389 (O_1389,N_19146,N_16804);
nor UO_1390 (O_1390,N_19967,N_16493);
nor UO_1391 (O_1391,N_16911,N_18609);
nor UO_1392 (O_1392,N_19422,N_17784);
and UO_1393 (O_1393,N_18433,N_18303);
or UO_1394 (O_1394,N_19851,N_17463);
or UO_1395 (O_1395,N_19701,N_17466);
xor UO_1396 (O_1396,N_18504,N_16538);
nor UO_1397 (O_1397,N_19151,N_19447);
and UO_1398 (O_1398,N_17309,N_18288);
nand UO_1399 (O_1399,N_19556,N_18876);
and UO_1400 (O_1400,N_19092,N_17668);
and UO_1401 (O_1401,N_18873,N_18768);
and UO_1402 (O_1402,N_17276,N_19737);
nor UO_1403 (O_1403,N_17374,N_16670);
nand UO_1404 (O_1404,N_17032,N_17814);
and UO_1405 (O_1405,N_19013,N_17067);
nand UO_1406 (O_1406,N_16485,N_18175);
nor UO_1407 (O_1407,N_19975,N_18478);
nand UO_1408 (O_1408,N_16520,N_19610);
nand UO_1409 (O_1409,N_19086,N_18794);
and UO_1410 (O_1410,N_16447,N_17298);
nor UO_1411 (O_1411,N_16361,N_19907);
and UO_1412 (O_1412,N_16793,N_18246);
or UO_1413 (O_1413,N_16638,N_18506);
or UO_1414 (O_1414,N_17193,N_16042);
and UO_1415 (O_1415,N_17566,N_17266);
and UO_1416 (O_1416,N_17753,N_18159);
nor UO_1417 (O_1417,N_18870,N_17866);
xnor UO_1418 (O_1418,N_18196,N_19123);
nand UO_1419 (O_1419,N_18844,N_19677);
and UO_1420 (O_1420,N_16556,N_16211);
xor UO_1421 (O_1421,N_18374,N_19870);
or UO_1422 (O_1422,N_18316,N_19073);
or UO_1423 (O_1423,N_17316,N_18519);
nor UO_1424 (O_1424,N_17015,N_16332);
and UO_1425 (O_1425,N_16635,N_19482);
or UO_1426 (O_1426,N_18199,N_17509);
and UO_1427 (O_1427,N_16207,N_19043);
nand UO_1428 (O_1428,N_19270,N_19980);
or UO_1429 (O_1429,N_17913,N_16544);
nor UO_1430 (O_1430,N_17557,N_17815);
or UO_1431 (O_1431,N_16079,N_18276);
nor UO_1432 (O_1432,N_19800,N_16158);
and UO_1433 (O_1433,N_19406,N_19492);
nand UO_1434 (O_1434,N_19392,N_16364);
nand UO_1435 (O_1435,N_16299,N_18428);
or UO_1436 (O_1436,N_17063,N_16488);
or UO_1437 (O_1437,N_17933,N_19859);
nor UO_1438 (O_1438,N_19140,N_17764);
xnor UO_1439 (O_1439,N_16203,N_18740);
nor UO_1440 (O_1440,N_16868,N_19705);
nand UO_1441 (O_1441,N_16532,N_18218);
nor UO_1442 (O_1442,N_17074,N_18305);
or UO_1443 (O_1443,N_17941,N_18648);
and UO_1444 (O_1444,N_19627,N_18565);
and UO_1445 (O_1445,N_19879,N_16439);
nand UO_1446 (O_1446,N_18232,N_18571);
nand UO_1447 (O_1447,N_17336,N_19663);
or UO_1448 (O_1448,N_17897,N_19174);
and UO_1449 (O_1449,N_18019,N_16015);
xor UO_1450 (O_1450,N_19228,N_17804);
or UO_1451 (O_1451,N_16218,N_19361);
nand UO_1452 (O_1452,N_17267,N_18180);
or UO_1453 (O_1453,N_18525,N_18015);
or UO_1454 (O_1454,N_17918,N_18231);
nand UO_1455 (O_1455,N_16193,N_18390);
nand UO_1456 (O_1456,N_17196,N_18387);
nor UO_1457 (O_1457,N_16314,N_17447);
and UO_1458 (O_1458,N_19230,N_19391);
and UO_1459 (O_1459,N_16873,N_18824);
and UO_1460 (O_1460,N_18016,N_17228);
nor UO_1461 (O_1461,N_18037,N_16090);
nor UO_1462 (O_1462,N_18119,N_19164);
and UO_1463 (O_1463,N_16879,N_19067);
nand UO_1464 (O_1464,N_18490,N_16874);
and UO_1465 (O_1465,N_17172,N_19751);
and UO_1466 (O_1466,N_16977,N_18115);
or UO_1467 (O_1467,N_17255,N_19372);
or UO_1468 (O_1468,N_17535,N_18418);
nor UO_1469 (O_1469,N_17452,N_17268);
nor UO_1470 (O_1470,N_19185,N_18649);
nor UO_1471 (O_1471,N_19611,N_16174);
nor UO_1472 (O_1472,N_16014,N_18094);
nor UO_1473 (O_1473,N_16517,N_16141);
nor UO_1474 (O_1474,N_16462,N_16969);
and UO_1475 (O_1475,N_18085,N_19527);
nor UO_1476 (O_1476,N_17064,N_19743);
and UO_1477 (O_1477,N_16521,N_18777);
nor UO_1478 (O_1478,N_18815,N_19427);
nand UO_1479 (O_1479,N_17947,N_17555);
nor UO_1480 (O_1480,N_19266,N_17573);
nand UO_1481 (O_1481,N_18517,N_17057);
or UO_1482 (O_1482,N_16089,N_19608);
or UO_1483 (O_1483,N_18383,N_18606);
or UO_1484 (O_1484,N_19885,N_18375);
nor UO_1485 (O_1485,N_17674,N_19149);
and UO_1486 (O_1486,N_16971,N_18169);
nor UO_1487 (O_1487,N_19243,N_19987);
nor UO_1488 (O_1488,N_19841,N_16234);
and UO_1489 (O_1489,N_18808,N_16555);
or UO_1490 (O_1490,N_19166,N_18800);
or UO_1491 (O_1491,N_17131,N_19809);
xnor UO_1492 (O_1492,N_17714,N_16792);
xnor UO_1493 (O_1493,N_16146,N_19909);
or UO_1494 (O_1494,N_18324,N_18190);
or UO_1495 (O_1495,N_16578,N_16383);
nor UO_1496 (O_1496,N_16100,N_16134);
nand UO_1497 (O_1497,N_17431,N_18862);
nor UO_1498 (O_1498,N_16333,N_18893);
and UO_1499 (O_1499,N_18460,N_19848);
or UO_1500 (O_1500,N_17517,N_18890);
and UO_1501 (O_1501,N_19242,N_17171);
nand UO_1502 (O_1502,N_19033,N_18716);
nor UO_1503 (O_1503,N_17293,N_17483);
or UO_1504 (O_1504,N_17830,N_19423);
nand UO_1505 (O_1505,N_18092,N_19647);
or UO_1506 (O_1506,N_18647,N_16131);
nand UO_1507 (O_1507,N_16808,N_17487);
xnor UO_1508 (O_1508,N_16435,N_19197);
nor UO_1509 (O_1509,N_17748,N_16001);
nor UO_1510 (O_1510,N_18932,N_18161);
nor UO_1511 (O_1511,N_16974,N_19019);
xnor UO_1512 (O_1512,N_16913,N_16128);
nor UO_1513 (O_1513,N_17192,N_16472);
and UO_1514 (O_1514,N_17687,N_17597);
nand UO_1515 (O_1515,N_18068,N_17807);
or UO_1516 (O_1516,N_19222,N_17179);
and UO_1517 (O_1517,N_18948,N_18400);
nor UO_1518 (O_1518,N_18773,N_19989);
or UO_1519 (O_1519,N_17796,N_18146);
nand UO_1520 (O_1520,N_18101,N_16091);
and UO_1521 (O_1521,N_17256,N_16281);
xnor UO_1522 (O_1522,N_16513,N_19205);
or UO_1523 (O_1523,N_19451,N_19920);
or UO_1524 (O_1524,N_16483,N_18999);
nor UO_1525 (O_1525,N_16630,N_17496);
and UO_1526 (O_1526,N_19822,N_17173);
or UO_1527 (O_1527,N_19601,N_19087);
or UO_1528 (O_1528,N_19613,N_17903);
nand UO_1529 (O_1529,N_19248,N_19637);
or UO_1530 (O_1530,N_18512,N_18237);
nand UO_1531 (O_1531,N_19191,N_19830);
nand UO_1532 (O_1532,N_18228,N_18522);
and UO_1533 (O_1533,N_17240,N_17016);
nor UO_1534 (O_1534,N_17041,N_18158);
and UO_1535 (O_1535,N_17985,N_18448);
nor UO_1536 (O_1536,N_16841,N_17197);
nand UO_1537 (O_1537,N_19421,N_17120);
nand UO_1538 (O_1538,N_16301,N_19584);
and UO_1539 (O_1539,N_19068,N_17741);
and UO_1540 (O_1540,N_18799,N_17206);
or UO_1541 (O_1541,N_16973,N_19126);
and UO_1542 (O_1542,N_18225,N_17510);
nand UO_1543 (O_1543,N_19355,N_16854);
or UO_1544 (O_1544,N_18140,N_16252);
and UO_1545 (O_1545,N_16752,N_18702);
nor UO_1546 (O_1546,N_19133,N_16829);
nand UO_1547 (O_1547,N_17159,N_18441);
nor UO_1548 (O_1548,N_17886,N_19272);
and UO_1549 (O_1549,N_18558,N_16092);
or UO_1550 (O_1550,N_18811,N_19357);
nand UO_1551 (O_1551,N_19901,N_18501);
or UO_1552 (O_1552,N_17121,N_16636);
xnor UO_1553 (O_1553,N_16851,N_19265);
or UO_1554 (O_1554,N_19196,N_16845);
or UO_1555 (O_1555,N_16883,N_18515);
or UO_1556 (O_1556,N_16415,N_17685);
nor UO_1557 (O_1557,N_18589,N_17045);
xor UO_1558 (O_1558,N_17997,N_17017);
nor UO_1559 (O_1559,N_18345,N_17828);
nand UO_1560 (O_1560,N_19784,N_16547);
nor UO_1561 (O_1561,N_16339,N_18102);
and UO_1562 (O_1562,N_16021,N_18248);
and UO_1563 (O_1563,N_17460,N_19772);
xnor UO_1564 (O_1564,N_17211,N_16593);
nand UO_1565 (O_1565,N_17654,N_16431);
nand UO_1566 (O_1566,N_18470,N_16641);
nor UO_1567 (O_1567,N_17109,N_18097);
nand UO_1568 (O_1568,N_17787,N_18912);
nor UO_1569 (O_1569,N_19746,N_18341);
nor UO_1570 (O_1570,N_17046,N_16197);
or UO_1571 (O_1571,N_16902,N_17467);
xor UO_1572 (O_1572,N_19927,N_17899);
and UO_1573 (O_1573,N_16261,N_16393);
nor UO_1574 (O_1574,N_17008,N_17054);
nand UO_1575 (O_1575,N_16275,N_19293);
nor UO_1576 (O_1576,N_17596,N_19756);
or UO_1577 (O_1577,N_17528,N_17619);
nor UO_1578 (O_1578,N_17825,N_16551);
nand UO_1579 (O_1579,N_17168,N_16905);
nand UO_1580 (O_1580,N_19398,N_18920);
nor UO_1581 (O_1581,N_18394,N_16798);
nand UO_1582 (O_1582,N_17635,N_18707);
nor UO_1583 (O_1583,N_18083,N_19615);
nor UO_1584 (O_1584,N_16157,N_17491);
or UO_1585 (O_1585,N_16842,N_16022);
xnor UO_1586 (O_1586,N_19972,N_18866);
nor UO_1587 (O_1587,N_16351,N_17330);
nor UO_1588 (O_1588,N_17030,N_18143);
nand UO_1589 (O_1589,N_18963,N_16618);
or UO_1590 (O_1590,N_16784,N_18329);
nor UO_1591 (O_1591,N_16689,N_18279);
nand UO_1592 (O_1592,N_18096,N_18502);
nand UO_1593 (O_1593,N_17872,N_16558);
and UO_1594 (O_1594,N_17136,N_17321);
xor UO_1595 (O_1595,N_19621,N_18339);
or UO_1596 (O_1596,N_19528,N_18285);
or UO_1597 (O_1597,N_16064,N_18833);
or UO_1598 (O_1598,N_19995,N_18372);
and UO_1599 (O_1599,N_19150,N_17175);
nand UO_1600 (O_1600,N_17143,N_18904);
and UO_1601 (O_1601,N_16686,N_17734);
xnor UO_1602 (O_1602,N_19050,N_16711);
nor UO_1603 (O_1603,N_17096,N_17544);
nor UO_1604 (O_1604,N_19189,N_19436);
and UO_1605 (O_1605,N_16230,N_19035);
and UO_1606 (O_1606,N_19452,N_17709);
and UO_1607 (O_1607,N_19114,N_19733);
and UO_1608 (O_1608,N_17836,N_17128);
and UO_1609 (O_1609,N_17537,N_17364);
nand UO_1610 (O_1610,N_16944,N_18806);
and UO_1611 (O_1611,N_16175,N_18561);
or UO_1612 (O_1612,N_17014,N_18421);
xnor UO_1613 (O_1613,N_17747,N_16597);
and UO_1614 (O_1614,N_18758,N_17865);
or UO_1615 (O_1615,N_18017,N_16484);
and UO_1616 (O_1616,N_19297,N_18381);
or UO_1617 (O_1617,N_18569,N_19718);
or UO_1618 (O_1618,N_19435,N_19534);
nor UO_1619 (O_1619,N_18269,N_19512);
nor UO_1620 (O_1620,N_17594,N_19329);
and UO_1621 (O_1621,N_17572,N_18878);
nand UO_1622 (O_1622,N_19913,N_17358);
nand UO_1623 (O_1623,N_17733,N_16251);
nand UO_1624 (O_1624,N_19184,N_19334);
nor UO_1625 (O_1625,N_19385,N_19213);
or UO_1626 (O_1626,N_16743,N_17370);
nor UO_1627 (O_1627,N_17634,N_18168);
xnor UO_1628 (O_1628,N_19670,N_19245);
and UO_1629 (O_1629,N_19624,N_16085);
and UO_1630 (O_1630,N_18454,N_19600);
nor UO_1631 (O_1631,N_19152,N_18918);
xor UO_1632 (O_1632,N_16101,N_17069);
and UO_1633 (O_1633,N_17862,N_16523);
nor UO_1634 (O_1634,N_16057,N_17418);
nor UO_1635 (O_1635,N_17317,N_19354);
nand UO_1636 (O_1636,N_16965,N_17075);
and UO_1637 (O_1637,N_17353,N_17322);
or UO_1638 (O_1638,N_18735,N_16970);
nor UO_1639 (O_1639,N_17663,N_19275);
or UO_1640 (O_1640,N_19130,N_18118);
or UO_1641 (O_1641,N_19416,N_16177);
xnor UO_1642 (O_1642,N_17247,N_18631);
or UO_1643 (O_1643,N_19513,N_18058);
nor UO_1644 (O_1644,N_16602,N_17325);
and UO_1645 (O_1645,N_16712,N_16701);
nand UO_1646 (O_1646,N_16681,N_19579);
nand UO_1647 (O_1647,N_19941,N_17908);
nor UO_1648 (O_1648,N_19868,N_17470);
nor UO_1649 (O_1649,N_19551,N_16240);
nand UO_1650 (O_1650,N_19567,N_18396);
and UO_1651 (O_1651,N_17595,N_18020);
and UO_1652 (O_1652,N_19785,N_18801);
xnor UO_1653 (O_1653,N_19251,N_18616);
nor UO_1654 (O_1654,N_17520,N_16122);
nor UO_1655 (O_1655,N_19618,N_18745);
or UO_1656 (O_1656,N_18564,N_19323);
xor UO_1657 (O_1657,N_16877,N_18654);
or UO_1658 (O_1658,N_17399,N_19327);
and UO_1659 (O_1659,N_16647,N_16456);
nor UO_1660 (O_1660,N_16839,N_16662);
nand UO_1661 (O_1661,N_18541,N_16869);
and UO_1662 (O_1662,N_18583,N_16759);
and UO_1663 (O_1663,N_18023,N_17779);
xnor UO_1664 (O_1664,N_16673,N_16677);
xnor UO_1665 (O_1665,N_17438,N_16781);
nand UO_1666 (O_1666,N_16027,N_17812);
nor UO_1667 (O_1667,N_18495,N_19582);
and UO_1668 (O_1668,N_19274,N_19689);
or UO_1669 (O_1669,N_19162,N_17036);
nor UO_1670 (O_1670,N_18022,N_16018);
and UO_1671 (O_1671,N_18721,N_17563);
and UO_1672 (O_1672,N_17451,N_19440);
xor UO_1673 (O_1673,N_17633,N_16082);
and UO_1674 (O_1674,N_18236,N_19917);
and UO_1675 (O_1675,N_17349,N_16675);
or UO_1676 (O_1676,N_17728,N_19792);
and UO_1677 (O_1677,N_19693,N_17942);
and UO_1678 (O_1678,N_18061,N_18837);
nand UO_1679 (O_1679,N_17283,N_16104);
nand UO_1680 (O_1680,N_16024,N_17059);
nor UO_1681 (O_1681,N_18960,N_19346);
or UO_1682 (O_1682,N_16341,N_19666);
and UO_1683 (O_1683,N_17181,N_16956);
or UO_1684 (O_1684,N_16561,N_16754);
and UO_1685 (O_1685,N_18684,N_18103);
nand UO_1686 (O_1686,N_18827,N_18909);
nand UO_1687 (O_1687,N_16238,N_19414);
nor UO_1688 (O_1688,N_18153,N_17547);
and UO_1689 (O_1689,N_16071,N_16434);
nand UO_1690 (O_1690,N_18882,N_18029);
or UO_1691 (O_1691,N_19839,N_17909);
nor UO_1692 (O_1692,N_18176,N_19464);
and UO_1693 (O_1693,N_19485,N_17475);
xor UO_1694 (O_1694,N_16652,N_18319);
nor UO_1695 (O_1695,N_19154,N_16005);
nand UO_1696 (O_1696,N_16552,N_17731);
nand UO_1697 (O_1697,N_16807,N_16041);
xor UO_1698 (O_1698,N_18582,N_17037);
xnor UO_1699 (O_1699,N_19169,N_18304);
or UO_1700 (O_1700,N_19165,N_16989);
or UO_1701 (O_1701,N_19335,N_19368);
nor UO_1702 (O_1702,N_18323,N_19840);
nor UO_1703 (O_1703,N_16991,N_18653);
or UO_1704 (O_1704,N_16893,N_16047);
nand UO_1705 (O_1705,N_16245,N_17290);
and UO_1706 (O_1706,N_19142,N_17068);
nor UO_1707 (O_1707,N_18451,N_19411);
nand UO_1708 (O_1708,N_19827,N_16880);
and UO_1709 (O_1709,N_18370,N_16766);
nor UO_1710 (O_1710,N_17287,N_19276);
nand UO_1711 (O_1711,N_16165,N_19626);
or UO_1712 (O_1712,N_18286,N_19289);
nor UO_1713 (O_1713,N_17718,N_16745);
nand UO_1714 (O_1714,N_17071,N_16225);
and UO_1715 (O_1715,N_18211,N_19983);
nor UO_1716 (O_1716,N_16198,N_17271);
and UO_1717 (O_1717,N_19856,N_19507);
nand UO_1718 (O_1718,N_17453,N_16506);
nand UO_1719 (O_1719,N_19519,N_18040);
nand UO_1720 (O_1720,N_16967,N_16885);
nand UO_1721 (O_1721,N_19163,N_16178);
or UO_1722 (O_1722,N_17174,N_18371);
and UO_1723 (O_1723,N_19458,N_17100);
nor UO_1724 (O_1724,N_19766,N_19042);
or UO_1725 (O_1725,N_16530,N_18840);
xor UO_1726 (O_1726,N_19669,N_16963);
and UO_1727 (O_1727,N_19569,N_18067);
or UO_1728 (O_1728,N_19409,N_18404);
and UO_1729 (O_1729,N_18744,N_17154);
nor UO_1730 (O_1730,N_18590,N_18767);
nand UO_1731 (O_1731,N_16655,N_16982);
or UO_1732 (O_1732,N_17388,N_16495);
xnor UO_1733 (O_1733,N_17699,N_19682);
and UO_1734 (O_1734,N_18486,N_16566);
nand UO_1735 (O_1735,N_19351,N_18498);
nor UO_1736 (O_1736,N_19802,N_16121);
and UO_1737 (O_1737,N_17248,N_16324);
nand UO_1738 (O_1738,N_19021,N_17871);
and UO_1739 (O_1739,N_19889,N_17775);
and UO_1740 (O_1740,N_16222,N_16594);
nand UO_1741 (O_1741,N_18348,N_18174);
and UO_1742 (O_1742,N_17148,N_17087);
nand UO_1743 (O_1743,N_18054,N_16643);
xnor UO_1744 (O_1744,N_19024,N_16737);
nand UO_1745 (O_1745,N_16360,N_16861);
and UO_1746 (O_1746,N_18672,N_18053);
and UO_1747 (O_1747,N_17740,N_16075);
and UO_1748 (O_1748,N_17023,N_19259);
nand UO_1749 (O_1749,N_17670,N_17739);
or UO_1750 (O_1750,N_18009,N_17081);
or UO_1751 (O_1751,N_18006,N_17964);
nand UO_1752 (O_1752,N_19910,N_16934);
xnor UO_1753 (O_1753,N_18988,N_18259);
nor UO_1754 (O_1754,N_18294,N_18632);
nor UO_1755 (O_1755,N_18397,N_17090);
or UO_1756 (O_1756,N_19874,N_19636);
and UO_1757 (O_1757,N_17361,N_17352);
nand UO_1758 (O_1758,N_19444,N_19853);
xor UO_1759 (O_1759,N_17489,N_19207);
or UO_1760 (O_1760,N_17757,N_16782);
nor UO_1761 (O_1761,N_16373,N_19922);
and UO_1762 (O_1762,N_18452,N_18188);
xnor UO_1763 (O_1763,N_16613,N_17390);
and UO_1764 (O_1764,N_19183,N_17548);
and UO_1765 (O_1765,N_18981,N_18151);
nand UO_1766 (O_1766,N_18307,N_19502);
and UO_1767 (O_1767,N_18755,N_17878);
or UO_1768 (O_1768,N_17526,N_18612);
and UO_1769 (O_1769,N_16680,N_17377);
nand UO_1770 (O_1770,N_17021,N_16614);
xnor UO_1771 (O_1771,N_19844,N_17551);
nand UO_1772 (O_1772,N_19060,N_19190);
nand UO_1773 (O_1773,N_16124,N_19286);
or UO_1774 (O_1774,N_16607,N_16628);
or UO_1775 (O_1775,N_16066,N_18538);
xnor UO_1776 (O_1776,N_19686,N_18300);
nand UO_1777 (O_1777,N_17079,N_18164);
or UO_1778 (O_1778,N_16870,N_18033);
or UO_1779 (O_1779,N_16352,N_17341);
and UO_1780 (O_1780,N_19565,N_16650);
and UO_1781 (O_1781,N_17604,N_16755);
and UO_1782 (O_1782,N_18595,N_16136);
or UO_1783 (O_1783,N_19951,N_16036);
nand UO_1784 (O_1784,N_17606,N_16917);
nor UO_1785 (O_1785,N_19732,N_18601);
and UO_1786 (O_1786,N_18570,N_17653);
nor UO_1787 (O_1787,N_16465,N_17429);
or UO_1788 (O_1788,N_19893,N_17000);
nand UO_1789 (O_1789,N_18203,N_17693);
or UO_1790 (O_1790,N_17504,N_16098);
nor UO_1791 (O_1791,N_19186,N_19774);
or UO_1792 (O_1792,N_18917,N_17294);
nand UO_1793 (O_1793,N_16127,N_17552);
and UO_1794 (O_1794,N_18204,N_18328);
nand UO_1795 (O_1795,N_16280,N_19918);
nor UO_1796 (O_1796,N_16639,N_17469);
nor UO_1797 (O_1797,N_19881,N_19336);
or UO_1798 (O_1798,N_16016,N_18407);
and UO_1799 (O_1799,N_17893,N_17752);
and UO_1800 (O_1800,N_16258,N_16043);
and UO_1801 (O_1801,N_16220,N_17094);
or UO_1802 (O_1802,N_19441,N_18289);
nor UO_1803 (O_1803,N_19816,N_16358);
xor UO_1804 (O_1804,N_17521,N_16486);
and UO_1805 (O_1805,N_18951,N_16029);
or UO_1806 (O_1806,N_17062,N_19886);
or UO_1807 (O_1807,N_17652,N_18185);
or UO_1808 (O_1808,N_19553,N_16559);
nor UO_1809 (O_1809,N_18227,N_18021);
nor UO_1810 (O_1810,N_17686,N_19471);
nand UO_1811 (O_1811,N_17164,N_18863);
nand UO_1812 (O_1812,N_16731,N_16715);
and UO_1813 (O_1813,N_16457,N_18585);
nor UO_1814 (O_1814,N_16243,N_17007);
or UO_1815 (O_1815,N_17708,N_16053);
nor UO_1816 (O_1816,N_19438,N_19981);
xor UO_1817 (O_1817,N_18325,N_18712);
and UO_1818 (O_1818,N_18825,N_17849);
xor UO_1819 (O_1819,N_17988,N_16886);
nor UO_1820 (O_1820,N_18427,N_17754);
nor UO_1821 (O_1821,N_18071,N_19962);
or UO_1822 (O_1822,N_17774,N_18064);
or UO_1823 (O_1823,N_18763,N_17631);
or UO_1824 (O_1824,N_19129,N_17238);
nor UO_1825 (O_1825,N_17929,N_16959);
or UO_1826 (O_1826,N_18642,N_18764);
nor UO_1827 (O_1827,N_17213,N_19083);
xor UO_1828 (O_1828,N_19494,N_18695);
or UO_1829 (O_1829,N_16531,N_16153);
nand UO_1830 (O_1830,N_16582,N_19727);
nor UO_1831 (O_1831,N_16159,N_18284);
xnor UO_1832 (O_1832,N_16726,N_18676);
nand UO_1833 (O_1833,N_17437,N_17039);
nand UO_1834 (O_1834,N_18437,N_16317);
xor UO_1835 (O_1835,N_16086,N_17498);
nand UO_1836 (O_1836,N_17986,N_18940);
nor UO_1837 (O_1837,N_19503,N_16863);
nand UO_1838 (O_1838,N_18958,N_19246);
or UO_1839 (O_1839,N_19898,N_16429);
or UO_1840 (O_1840,N_17919,N_19366);
and UO_1841 (O_1841,N_18973,N_18036);
nand UO_1842 (O_1842,N_19171,N_19179);
nand UO_1843 (O_1843,N_19694,N_17115);
or UO_1844 (O_1844,N_18993,N_18124);
or UO_1845 (O_1845,N_19088,N_17103);
nor UO_1846 (O_1846,N_16514,N_17138);
and UO_1847 (O_1847,N_16479,N_19657);
and UO_1848 (O_1848,N_18001,N_16624);
nor UO_1849 (O_1849,N_18264,N_18031);
nand UO_1850 (O_1850,N_16078,N_18014);
or UO_1851 (O_1851,N_16899,N_17931);
nand UO_1852 (O_1852,N_18043,N_19660);
and UO_1853 (O_1853,N_17005,N_16340);
or UO_1854 (O_1854,N_19680,N_17887);
nand UO_1855 (O_1855,N_17955,N_17331);
nor UO_1856 (O_1856,N_19997,N_18184);
or UO_1857 (O_1857,N_16315,N_17432);
nand UO_1858 (O_1858,N_16118,N_16191);
xnor UO_1859 (O_1859,N_18089,N_18766);
nand UO_1860 (O_1860,N_18117,N_17833);
nand UO_1861 (O_1861,N_18459,N_16921);
nand UO_1862 (O_1862,N_18987,N_16634);
xor UO_1863 (O_1863,N_19978,N_18051);
nor UO_1864 (O_1864,N_19985,N_18915);
nor UO_1865 (O_1865,N_18420,N_19127);
nor UO_1866 (O_1866,N_16751,N_16867);
and UO_1867 (O_1867,N_17389,N_17777);
and UO_1868 (O_1868,N_17783,N_16395);
and UO_1869 (O_1869,N_16697,N_17472);
xor UO_1870 (O_1870,N_17799,N_19783);
nand UO_1871 (O_1871,N_19762,N_18209);
nor UO_1872 (O_1872,N_18379,N_17398);
or UO_1873 (O_1873,N_19617,N_18559);
or UO_1874 (O_1874,N_16426,N_18072);
xor UO_1875 (O_1875,N_19607,N_19592);
xnor UO_1876 (O_1876,N_19895,N_17554);
nor UO_1877 (O_1877,N_19923,N_19549);
xnor UO_1878 (O_1878,N_18902,N_16228);
or UO_1879 (O_1879,N_18111,N_18983);
xnor UO_1880 (O_1880,N_18971,N_19558);
xor UO_1881 (O_1881,N_18136,N_18107);
nand UO_1882 (O_1882,N_16927,N_19356);
nor UO_1883 (O_1883,N_18663,N_16840);
nand UO_1884 (O_1884,N_18661,N_17620);
or UO_1885 (O_1885,N_17746,N_16182);
or UO_1886 (O_1886,N_16964,N_17789);
and UO_1887 (O_1887,N_16783,N_16714);
or UO_1888 (O_1888,N_18414,N_18780);
xor UO_1889 (O_1889,N_17735,N_19084);
or UO_1890 (O_1890,N_16736,N_17946);
nand UO_1891 (O_1891,N_19386,N_19590);
nand UO_1892 (O_1892,N_16216,N_19658);
and UO_1893 (O_1893,N_18010,N_18738);
xnor UO_1894 (O_1894,N_19620,N_19261);
nand UO_1895 (O_1895,N_17351,N_17222);
nor UO_1896 (O_1896,N_17462,N_16935);
and UO_1897 (O_1897,N_19717,N_16446);
or UO_1898 (O_1898,N_18377,N_16233);
and UO_1899 (O_1899,N_19134,N_16984);
or UO_1900 (O_1900,N_18896,N_18413);
nand UO_1901 (O_1901,N_19845,N_18139);
xnor UO_1902 (O_1902,N_16720,N_19384);
nor UO_1903 (O_1903,N_19760,N_16420);
xor UO_1904 (O_1904,N_19256,N_18249);
nor UO_1905 (O_1905,N_18056,N_18281);
and UO_1906 (O_1906,N_18086,N_18520);
and UO_1907 (O_1907,N_17058,N_17209);
or UO_1908 (O_1908,N_16359,N_19255);
nand UO_1909 (O_1909,N_16734,N_18162);
or UO_1910 (O_1910,N_18860,N_19706);
nor UO_1911 (O_1911,N_17969,N_16007);
nor UO_1912 (O_1912,N_16785,N_18417);
nand UO_1913 (O_1913,N_18444,N_19362);
xnor UO_1914 (O_1914,N_17549,N_17582);
nand UO_1915 (O_1915,N_19834,N_17649);
nand UO_1916 (O_1916,N_18121,N_17730);
or UO_1917 (O_1917,N_16653,N_16633);
nor UO_1918 (O_1918,N_17326,N_16891);
nand UO_1919 (O_1919,N_17970,N_18035);
and UO_1920 (O_1920,N_18315,N_18457);
nor UO_1921 (O_1921,N_19933,N_18544);
nand UO_1922 (O_1922,N_17334,N_16659);
nor UO_1923 (O_1923,N_17444,N_17221);
nor UO_1924 (O_1924,N_19252,N_19113);
xnor UO_1925 (O_1925,N_16966,N_16501);
nand UO_1926 (O_1926,N_16598,N_17034);
nand UO_1927 (O_1927,N_19311,N_17694);
nand UO_1928 (O_1928,N_16698,N_16503);
and UO_1929 (O_1929,N_18423,N_19684);
nor UO_1930 (O_1930,N_18598,N_16058);
or UO_1931 (O_1931,N_17788,N_17391);
nor UO_1932 (O_1932,N_17692,N_18012);
nand UO_1933 (O_1933,N_17749,N_19557);
and UO_1934 (O_1934,N_17026,N_16865);
xor UO_1935 (O_1935,N_18171,N_18082);
xnor UO_1936 (O_1936,N_16730,N_18572);
or UO_1937 (O_1937,N_16801,N_17618);
nor UO_1938 (O_1938,N_19938,N_19011);
nor UO_1939 (O_1939,N_17375,N_19616);
nor UO_1940 (O_1940,N_18997,N_18144);
xor UO_1941 (O_1941,N_17587,N_17297);
nand UO_1942 (O_1942,N_16787,N_17870);
or UO_1943 (O_1943,N_16780,N_17319);
and UO_1944 (O_1944,N_18792,N_17405);
or UO_1945 (O_1945,N_18871,N_16348);
and UO_1946 (O_1946,N_18718,N_19128);
or UO_1947 (O_1947,N_16156,N_18739);
nor UO_1948 (O_1948,N_18145,N_18903);
and UO_1949 (O_1949,N_18104,N_16330);
nor UO_1950 (O_1950,N_16072,N_16335);
nand UO_1951 (O_1951,N_18002,N_19000);
nor UO_1952 (O_1952,N_18959,N_16452);
nor UO_1953 (O_1953,N_19606,N_18152);
and UO_1954 (O_1954,N_19570,N_17082);
and UO_1955 (O_1955,N_19053,N_19661);
nand UO_1956 (O_1956,N_16537,N_16931);
nor UO_1957 (O_1957,N_17850,N_16482);
nand UO_1958 (O_1958,N_19153,N_16691);
and UO_1959 (O_1959,N_17944,N_16145);
nor UO_1960 (O_1960,N_19787,N_18812);
nand UO_1961 (O_1961,N_18384,N_17827);
or UO_1962 (O_1962,N_18503,N_19643);
nor UO_1963 (O_1963,N_17056,N_18771);
and UO_1964 (O_1964,N_17441,N_16584);
nand UO_1965 (O_1965,N_16437,N_19426);
nand UO_1966 (O_1966,N_17579,N_16260);
nor UO_1967 (O_1967,N_19450,N_19642);
and UO_1968 (O_1968,N_19319,N_16947);
nor UO_1969 (O_1969,N_19510,N_18620);
nand UO_1970 (O_1970,N_16739,N_18331);
xor UO_1971 (O_1971,N_17078,N_18106);
nor UO_1972 (O_1972,N_17832,N_17134);
xor UO_1973 (O_1973,N_17486,N_16433);
xor UO_1974 (O_1974,N_19054,N_16262);
nand UO_1975 (O_1975,N_17166,N_18008);
nor UO_1976 (O_1976,N_17568,N_16834);
and UO_1977 (O_1977,N_19662,N_17738);
nor UO_1978 (O_1978,N_17025,N_17745);
and UO_1979 (O_1979,N_17626,N_19865);
xnor UO_1980 (O_1980,N_17177,N_18614);
or UO_1981 (O_1981,N_18160,N_16723);
nand UO_1982 (O_1982,N_17185,N_17651);
xor UO_1983 (O_1983,N_18113,N_17190);
nand UO_1984 (O_1984,N_19741,N_19090);
and UO_1985 (O_1985,N_16732,N_17533);
or UO_1986 (O_1986,N_19498,N_18652);
and UO_1987 (O_1987,N_16660,N_18727);
nor UO_1988 (O_1988,N_18657,N_17583);
and UO_1989 (O_1989,N_18830,N_16223);
nand UO_1990 (O_1990,N_16892,N_18604);
or UO_1991 (O_1991,N_18931,N_17864);
and UO_1992 (O_1992,N_18937,N_19597);
and UO_1993 (O_1993,N_18977,N_17954);
xor UO_1994 (O_1994,N_18141,N_19400);
or UO_1995 (O_1995,N_19619,N_18474);
nand UO_1996 (O_1996,N_17629,N_19768);
nor UO_1997 (O_1997,N_17155,N_16695);
nand UO_1998 (O_1998,N_18148,N_19491);
and UO_1999 (O_1999,N_19277,N_19061);
nor UO_2000 (O_2000,N_19819,N_17195);
and UO_2001 (O_2001,N_19390,N_18418);
or UO_2002 (O_2002,N_16417,N_17087);
xnor UO_2003 (O_2003,N_19323,N_16062);
and UO_2004 (O_2004,N_16857,N_18392);
or UO_2005 (O_2005,N_16601,N_18934);
and UO_2006 (O_2006,N_19769,N_16359);
xnor UO_2007 (O_2007,N_18748,N_16716);
nand UO_2008 (O_2008,N_19207,N_19677);
nor UO_2009 (O_2009,N_17747,N_17010);
nor UO_2010 (O_2010,N_16262,N_19911);
xor UO_2011 (O_2011,N_16684,N_17159);
xnor UO_2012 (O_2012,N_17994,N_17393);
and UO_2013 (O_2013,N_16646,N_17487);
nor UO_2014 (O_2014,N_18914,N_16904);
or UO_2015 (O_2015,N_16683,N_19259);
nand UO_2016 (O_2016,N_17665,N_16767);
nor UO_2017 (O_2017,N_19420,N_18244);
nand UO_2018 (O_2018,N_19367,N_16806);
and UO_2019 (O_2019,N_16715,N_16960);
xnor UO_2020 (O_2020,N_18847,N_18179);
nand UO_2021 (O_2021,N_17080,N_16147);
or UO_2022 (O_2022,N_19090,N_19117);
nand UO_2023 (O_2023,N_16046,N_16829);
or UO_2024 (O_2024,N_19583,N_17354);
or UO_2025 (O_2025,N_16920,N_17170);
nor UO_2026 (O_2026,N_18119,N_17332);
nand UO_2027 (O_2027,N_16855,N_17895);
nand UO_2028 (O_2028,N_19822,N_19151);
nor UO_2029 (O_2029,N_16287,N_17572);
xnor UO_2030 (O_2030,N_18436,N_17139);
nand UO_2031 (O_2031,N_18337,N_17048);
nor UO_2032 (O_2032,N_16244,N_19794);
nand UO_2033 (O_2033,N_16626,N_19561);
nor UO_2034 (O_2034,N_18269,N_18136);
or UO_2035 (O_2035,N_19833,N_18669);
nor UO_2036 (O_2036,N_19735,N_18948);
nand UO_2037 (O_2037,N_16254,N_17847);
and UO_2038 (O_2038,N_18354,N_17512);
nor UO_2039 (O_2039,N_16037,N_16358);
nand UO_2040 (O_2040,N_16163,N_16962);
and UO_2041 (O_2041,N_17256,N_17671);
or UO_2042 (O_2042,N_19999,N_16325);
or UO_2043 (O_2043,N_18393,N_16529);
and UO_2044 (O_2044,N_16686,N_18839);
or UO_2045 (O_2045,N_18720,N_16406);
nor UO_2046 (O_2046,N_18987,N_18141);
xor UO_2047 (O_2047,N_18222,N_18750);
xnor UO_2048 (O_2048,N_19648,N_19831);
or UO_2049 (O_2049,N_16715,N_19552);
nor UO_2050 (O_2050,N_17495,N_17352);
and UO_2051 (O_2051,N_16912,N_17271);
and UO_2052 (O_2052,N_19495,N_16510);
nor UO_2053 (O_2053,N_16781,N_18807);
nor UO_2054 (O_2054,N_16534,N_19114);
nor UO_2055 (O_2055,N_19587,N_18697);
and UO_2056 (O_2056,N_16962,N_16235);
nor UO_2057 (O_2057,N_17858,N_19684);
and UO_2058 (O_2058,N_19682,N_17294);
or UO_2059 (O_2059,N_17071,N_17007);
or UO_2060 (O_2060,N_18139,N_17864);
nor UO_2061 (O_2061,N_18315,N_17207);
xnor UO_2062 (O_2062,N_16056,N_19967);
nor UO_2063 (O_2063,N_19458,N_16389);
nor UO_2064 (O_2064,N_17836,N_17047);
or UO_2065 (O_2065,N_19709,N_19750);
and UO_2066 (O_2066,N_19605,N_19405);
nand UO_2067 (O_2067,N_18206,N_18560);
or UO_2068 (O_2068,N_19596,N_18199);
xor UO_2069 (O_2069,N_17789,N_17571);
or UO_2070 (O_2070,N_17106,N_16838);
or UO_2071 (O_2071,N_19446,N_18058);
nand UO_2072 (O_2072,N_19365,N_17611);
or UO_2073 (O_2073,N_19519,N_19493);
nand UO_2074 (O_2074,N_16301,N_19809);
nand UO_2075 (O_2075,N_18940,N_19831);
or UO_2076 (O_2076,N_17132,N_16553);
or UO_2077 (O_2077,N_17147,N_17696);
nor UO_2078 (O_2078,N_16068,N_19700);
nand UO_2079 (O_2079,N_16108,N_19211);
nor UO_2080 (O_2080,N_17246,N_16601);
nor UO_2081 (O_2081,N_17541,N_17007);
and UO_2082 (O_2082,N_19984,N_17985);
and UO_2083 (O_2083,N_16967,N_16905);
xnor UO_2084 (O_2084,N_19182,N_17305);
and UO_2085 (O_2085,N_19487,N_19167);
and UO_2086 (O_2086,N_18547,N_18551);
nor UO_2087 (O_2087,N_18515,N_19347);
and UO_2088 (O_2088,N_17113,N_18532);
and UO_2089 (O_2089,N_18629,N_17154);
nor UO_2090 (O_2090,N_19452,N_18770);
and UO_2091 (O_2091,N_19299,N_19095);
or UO_2092 (O_2092,N_18491,N_16033);
nand UO_2093 (O_2093,N_17331,N_17231);
nor UO_2094 (O_2094,N_16359,N_16239);
xnor UO_2095 (O_2095,N_19086,N_16325);
and UO_2096 (O_2096,N_17264,N_16642);
or UO_2097 (O_2097,N_16063,N_19637);
or UO_2098 (O_2098,N_18969,N_18492);
or UO_2099 (O_2099,N_18481,N_19998);
nand UO_2100 (O_2100,N_18845,N_18468);
and UO_2101 (O_2101,N_17515,N_19302);
and UO_2102 (O_2102,N_19582,N_18684);
or UO_2103 (O_2103,N_17144,N_19906);
or UO_2104 (O_2104,N_19053,N_16397);
or UO_2105 (O_2105,N_18160,N_16670);
or UO_2106 (O_2106,N_18666,N_17736);
xnor UO_2107 (O_2107,N_18374,N_18270);
nand UO_2108 (O_2108,N_19485,N_16186);
nand UO_2109 (O_2109,N_17778,N_19511);
and UO_2110 (O_2110,N_16349,N_17519);
nand UO_2111 (O_2111,N_16331,N_19477);
nor UO_2112 (O_2112,N_19586,N_18424);
or UO_2113 (O_2113,N_18849,N_16991);
or UO_2114 (O_2114,N_19196,N_18664);
and UO_2115 (O_2115,N_18775,N_17308);
and UO_2116 (O_2116,N_18327,N_18800);
and UO_2117 (O_2117,N_17435,N_17043);
or UO_2118 (O_2118,N_17591,N_16302);
or UO_2119 (O_2119,N_16836,N_16699);
nor UO_2120 (O_2120,N_17007,N_19529);
or UO_2121 (O_2121,N_16419,N_19067);
nor UO_2122 (O_2122,N_16146,N_17551);
nand UO_2123 (O_2123,N_16694,N_16453);
and UO_2124 (O_2124,N_19492,N_18086);
or UO_2125 (O_2125,N_17496,N_16716);
or UO_2126 (O_2126,N_18216,N_18518);
and UO_2127 (O_2127,N_18249,N_18851);
and UO_2128 (O_2128,N_18508,N_16289);
and UO_2129 (O_2129,N_19115,N_19433);
and UO_2130 (O_2130,N_19959,N_18559);
nand UO_2131 (O_2131,N_19303,N_18850);
nand UO_2132 (O_2132,N_19526,N_18833);
and UO_2133 (O_2133,N_17939,N_17864);
and UO_2134 (O_2134,N_17940,N_18086);
and UO_2135 (O_2135,N_18205,N_19468);
or UO_2136 (O_2136,N_18384,N_17047);
or UO_2137 (O_2137,N_17117,N_18044);
or UO_2138 (O_2138,N_19695,N_18505);
nand UO_2139 (O_2139,N_16063,N_16179);
nor UO_2140 (O_2140,N_18796,N_16896);
xor UO_2141 (O_2141,N_17350,N_18272);
or UO_2142 (O_2142,N_19489,N_18529);
nor UO_2143 (O_2143,N_17107,N_17353);
or UO_2144 (O_2144,N_17286,N_18942);
nand UO_2145 (O_2145,N_19899,N_19270);
and UO_2146 (O_2146,N_17954,N_19248);
nand UO_2147 (O_2147,N_19888,N_17010);
or UO_2148 (O_2148,N_16978,N_16039);
or UO_2149 (O_2149,N_16858,N_19666);
or UO_2150 (O_2150,N_17822,N_16735);
or UO_2151 (O_2151,N_18676,N_17696);
or UO_2152 (O_2152,N_18658,N_16741);
nor UO_2153 (O_2153,N_16864,N_19611);
and UO_2154 (O_2154,N_17882,N_16381);
nand UO_2155 (O_2155,N_18669,N_18222);
and UO_2156 (O_2156,N_17612,N_19027);
nand UO_2157 (O_2157,N_18203,N_16764);
xor UO_2158 (O_2158,N_17485,N_18971);
nand UO_2159 (O_2159,N_18998,N_16907);
xnor UO_2160 (O_2160,N_17775,N_18312);
and UO_2161 (O_2161,N_19715,N_18420);
or UO_2162 (O_2162,N_17588,N_18180);
or UO_2163 (O_2163,N_16570,N_16824);
and UO_2164 (O_2164,N_17379,N_17504);
and UO_2165 (O_2165,N_19584,N_17195);
nor UO_2166 (O_2166,N_16821,N_16636);
and UO_2167 (O_2167,N_17851,N_17110);
and UO_2168 (O_2168,N_18369,N_17435);
nor UO_2169 (O_2169,N_17374,N_17595);
nand UO_2170 (O_2170,N_16686,N_16936);
nor UO_2171 (O_2171,N_16440,N_16385);
nor UO_2172 (O_2172,N_17084,N_18734);
or UO_2173 (O_2173,N_19214,N_19165);
xnor UO_2174 (O_2174,N_16614,N_17679);
and UO_2175 (O_2175,N_19437,N_17684);
or UO_2176 (O_2176,N_19639,N_19470);
or UO_2177 (O_2177,N_17791,N_16044);
or UO_2178 (O_2178,N_19037,N_17636);
nor UO_2179 (O_2179,N_17905,N_19678);
nor UO_2180 (O_2180,N_19386,N_17578);
nor UO_2181 (O_2181,N_16624,N_16011);
and UO_2182 (O_2182,N_18029,N_16911);
and UO_2183 (O_2183,N_16893,N_19786);
or UO_2184 (O_2184,N_16985,N_17910);
nor UO_2185 (O_2185,N_16162,N_19612);
or UO_2186 (O_2186,N_17399,N_17827);
and UO_2187 (O_2187,N_16786,N_16348);
and UO_2188 (O_2188,N_19636,N_19892);
or UO_2189 (O_2189,N_19319,N_17911);
and UO_2190 (O_2190,N_19984,N_16307);
xor UO_2191 (O_2191,N_17883,N_18279);
or UO_2192 (O_2192,N_16330,N_16487);
nor UO_2193 (O_2193,N_16835,N_16882);
nand UO_2194 (O_2194,N_16907,N_16996);
or UO_2195 (O_2195,N_17440,N_19436);
nor UO_2196 (O_2196,N_19961,N_18591);
nand UO_2197 (O_2197,N_17535,N_16195);
and UO_2198 (O_2198,N_17999,N_19553);
nand UO_2199 (O_2199,N_16787,N_19257);
xor UO_2200 (O_2200,N_16668,N_16735);
nor UO_2201 (O_2201,N_16886,N_17319);
nor UO_2202 (O_2202,N_19987,N_19947);
and UO_2203 (O_2203,N_17970,N_19591);
or UO_2204 (O_2204,N_18513,N_19190);
or UO_2205 (O_2205,N_19632,N_18120);
and UO_2206 (O_2206,N_16839,N_18393);
nor UO_2207 (O_2207,N_16280,N_16727);
xor UO_2208 (O_2208,N_17524,N_19394);
xnor UO_2209 (O_2209,N_17154,N_18726);
nand UO_2210 (O_2210,N_18793,N_18911);
nand UO_2211 (O_2211,N_16225,N_17795);
or UO_2212 (O_2212,N_19503,N_19618);
nand UO_2213 (O_2213,N_17279,N_19260);
or UO_2214 (O_2214,N_19316,N_17751);
nand UO_2215 (O_2215,N_17732,N_18657);
nand UO_2216 (O_2216,N_16182,N_19189);
or UO_2217 (O_2217,N_16326,N_17025);
and UO_2218 (O_2218,N_18410,N_16494);
nor UO_2219 (O_2219,N_17257,N_16552);
nand UO_2220 (O_2220,N_17956,N_18945);
and UO_2221 (O_2221,N_16619,N_17648);
nand UO_2222 (O_2222,N_18424,N_16443);
or UO_2223 (O_2223,N_16747,N_17134);
or UO_2224 (O_2224,N_19382,N_19031);
or UO_2225 (O_2225,N_19146,N_19577);
or UO_2226 (O_2226,N_17671,N_17665);
or UO_2227 (O_2227,N_16970,N_17194);
and UO_2228 (O_2228,N_16300,N_18588);
xnor UO_2229 (O_2229,N_18399,N_16774);
and UO_2230 (O_2230,N_19095,N_19896);
or UO_2231 (O_2231,N_19857,N_17596);
and UO_2232 (O_2232,N_18364,N_19185);
nand UO_2233 (O_2233,N_18221,N_16658);
nand UO_2234 (O_2234,N_19372,N_19797);
or UO_2235 (O_2235,N_18696,N_19791);
xnor UO_2236 (O_2236,N_16860,N_17124);
nand UO_2237 (O_2237,N_19264,N_17151);
nor UO_2238 (O_2238,N_17680,N_17807);
or UO_2239 (O_2239,N_18059,N_17907);
and UO_2240 (O_2240,N_16766,N_19677);
and UO_2241 (O_2241,N_17640,N_18251);
and UO_2242 (O_2242,N_19227,N_17183);
xnor UO_2243 (O_2243,N_16223,N_17512);
nor UO_2244 (O_2244,N_18371,N_18975);
xnor UO_2245 (O_2245,N_16782,N_17408);
and UO_2246 (O_2246,N_17134,N_17844);
nand UO_2247 (O_2247,N_16765,N_16722);
nor UO_2248 (O_2248,N_18972,N_19401);
nor UO_2249 (O_2249,N_16732,N_19457);
nor UO_2250 (O_2250,N_18431,N_19887);
nand UO_2251 (O_2251,N_19462,N_19953);
and UO_2252 (O_2252,N_17956,N_16062);
nand UO_2253 (O_2253,N_16396,N_19869);
or UO_2254 (O_2254,N_18916,N_19296);
nor UO_2255 (O_2255,N_16721,N_17968);
and UO_2256 (O_2256,N_17077,N_19939);
nor UO_2257 (O_2257,N_16517,N_18092);
and UO_2258 (O_2258,N_16616,N_16335);
or UO_2259 (O_2259,N_19008,N_19393);
nand UO_2260 (O_2260,N_16080,N_16828);
or UO_2261 (O_2261,N_17958,N_19243);
nor UO_2262 (O_2262,N_19723,N_17193);
or UO_2263 (O_2263,N_17137,N_16329);
nor UO_2264 (O_2264,N_19900,N_17247);
nand UO_2265 (O_2265,N_17992,N_17288);
and UO_2266 (O_2266,N_17161,N_17425);
and UO_2267 (O_2267,N_17727,N_17690);
nand UO_2268 (O_2268,N_16088,N_17005);
nand UO_2269 (O_2269,N_16779,N_16314);
xnor UO_2270 (O_2270,N_19944,N_19566);
and UO_2271 (O_2271,N_16950,N_16528);
or UO_2272 (O_2272,N_19615,N_19717);
and UO_2273 (O_2273,N_18392,N_16100);
nor UO_2274 (O_2274,N_17889,N_17018);
and UO_2275 (O_2275,N_17089,N_16435);
nor UO_2276 (O_2276,N_16906,N_19678);
xnor UO_2277 (O_2277,N_17044,N_17425);
nand UO_2278 (O_2278,N_19032,N_17668);
or UO_2279 (O_2279,N_19701,N_19966);
nor UO_2280 (O_2280,N_17727,N_18898);
and UO_2281 (O_2281,N_19123,N_19552);
or UO_2282 (O_2282,N_17981,N_16868);
and UO_2283 (O_2283,N_18512,N_17678);
and UO_2284 (O_2284,N_19682,N_16199);
nand UO_2285 (O_2285,N_19774,N_18458);
nand UO_2286 (O_2286,N_16628,N_19147);
nand UO_2287 (O_2287,N_16361,N_16292);
or UO_2288 (O_2288,N_18453,N_17573);
nand UO_2289 (O_2289,N_16487,N_17167);
nand UO_2290 (O_2290,N_16405,N_19719);
or UO_2291 (O_2291,N_19970,N_17734);
nor UO_2292 (O_2292,N_17787,N_16239);
or UO_2293 (O_2293,N_19501,N_16476);
nor UO_2294 (O_2294,N_18784,N_18362);
xnor UO_2295 (O_2295,N_19189,N_17178);
nand UO_2296 (O_2296,N_19385,N_16639);
nor UO_2297 (O_2297,N_19736,N_18671);
or UO_2298 (O_2298,N_19202,N_19832);
and UO_2299 (O_2299,N_17329,N_19391);
nor UO_2300 (O_2300,N_19153,N_19203);
or UO_2301 (O_2301,N_18972,N_17775);
or UO_2302 (O_2302,N_19075,N_16332);
nor UO_2303 (O_2303,N_19557,N_18007);
nor UO_2304 (O_2304,N_16019,N_19303);
and UO_2305 (O_2305,N_16268,N_18119);
or UO_2306 (O_2306,N_17887,N_17815);
nand UO_2307 (O_2307,N_17170,N_16908);
or UO_2308 (O_2308,N_19496,N_17035);
or UO_2309 (O_2309,N_19000,N_18081);
nor UO_2310 (O_2310,N_19385,N_17744);
nand UO_2311 (O_2311,N_18163,N_18398);
and UO_2312 (O_2312,N_19112,N_17157);
or UO_2313 (O_2313,N_18695,N_17662);
or UO_2314 (O_2314,N_18128,N_19396);
and UO_2315 (O_2315,N_19704,N_18957);
and UO_2316 (O_2316,N_19181,N_17211);
nor UO_2317 (O_2317,N_17271,N_19806);
and UO_2318 (O_2318,N_19025,N_16965);
and UO_2319 (O_2319,N_16598,N_17427);
and UO_2320 (O_2320,N_16306,N_19429);
nor UO_2321 (O_2321,N_19044,N_17339);
nor UO_2322 (O_2322,N_17043,N_19099);
and UO_2323 (O_2323,N_18775,N_17154);
or UO_2324 (O_2324,N_18227,N_16103);
or UO_2325 (O_2325,N_18727,N_19910);
nor UO_2326 (O_2326,N_19943,N_17942);
nor UO_2327 (O_2327,N_19821,N_17484);
nand UO_2328 (O_2328,N_16706,N_18166);
and UO_2329 (O_2329,N_17216,N_16007);
and UO_2330 (O_2330,N_18243,N_17238);
nor UO_2331 (O_2331,N_17808,N_19394);
or UO_2332 (O_2332,N_16499,N_18644);
xnor UO_2333 (O_2333,N_17560,N_19294);
nand UO_2334 (O_2334,N_18377,N_19791);
nand UO_2335 (O_2335,N_19973,N_16769);
and UO_2336 (O_2336,N_16013,N_16477);
or UO_2337 (O_2337,N_16060,N_16214);
nor UO_2338 (O_2338,N_16637,N_16571);
nor UO_2339 (O_2339,N_19303,N_18160);
or UO_2340 (O_2340,N_16873,N_16703);
xor UO_2341 (O_2341,N_19553,N_18636);
nand UO_2342 (O_2342,N_16907,N_19985);
nor UO_2343 (O_2343,N_17841,N_16600);
nand UO_2344 (O_2344,N_16979,N_17219);
or UO_2345 (O_2345,N_17949,N_17755);
and UO_2346 (O_2346,N_18005,N_19571);
nor UO_2347 (O_2347,N_19153,N_17175);
or UO_2348 (O_2348,N_17298,N_17033);
xor UO_2349 (O_2349,N_17075,N_16707);
or UO_2350 (O_2350,N_19462,N_17268);
and UO_2351 (O_2351,N_16816,N_17812);
nor UO_2352 (O_2352,N_17049,N_16697);
and UO_2353 (O_2353,N_19098,N_16075);
or UO_2354 (O_2354,N_18702,N_18936);
and UO_2355 (O_2355,N_18105,N_19154);
nor UO_2356 (O_2356,N_16532,N_18461);
and UO_2357 (O_2357,N_17232,N_17361);
or UO_2358 (O_2358,N_17230,N_16414);
and UO_2359 (O_2359,N_19053,N_19775);
or UO_2360 (O_2360,N_18996,N_17726);
xnor UO_2361 (O_2361,N_19955,N_16898);
xor UO_2362 (O_2362,N_17504,N_19727);
and UO_2363 (O_2363,N_16182,N_17791);
xor UO_2364 (O_2364,N_16119,N_17892);
or UO_2365 (O_2365,N_19274,N_17018);
nor UO_2366 (O_2366,N_16471,N_16095);
xor UO_2367 (O_2367,N_19880,N_18348);
and UO_2368 (O_2368,N_18306,N_19377);
nand UO_2369 (O_2369,N_16972,N_16504);
or UO_2370 (O_2370,N_17010,N_19255);
and UO_2371 (O_2371,N_17376,N_17131);
and UO_2372 (O_2372,N_18844,N_16317);
nor UO_2373 (O_2373,N_18892,N_19188);
xor UO_2374 (O_2374,N_17904,N_19439);
nor UO_2375 (O_2375,N_19378,N_17180);
or UO_2376 (O_2376,N_16978,N_17238);
nor UO_2377 (O_2377,N_19409,N_18425);
nor UO_2378 (O_2378,N_18545,N_16953);
and UO_2379 (O_2379,N_18482,N_19862);
nand UO_2380 (O_2380,N_18322,N_16801);
nor UO_2381 (O_2381,N_17951,N_17000);
nand UO_2382 (O_2382,N_19717,N_18619);
nand UO_2383 (O_2383,N_16858,N_16198);
nor UO_2384 (O_2384,N_18171,N_19025);
xnor UO_2385 (O_2385,N_19236,N_17344);
nor UO_2386 (O_2386,N_19415,N_18097);
and UO_2387 (O_2387,N_17104,N_19014);
nor UO_2388 (O_2388,N_18077,N_18067);
nor UO_2389 (O_2389,N_18571,N_18125);
or UO_2390 (O_2390,N_19358,N_16476);
xnor UO_2391 (O_2391,N_19484,N_18192);
nor UO_2392 (O_2392,N_17735,N_18631);
or UO_2393 (O_2393,N_18348,N_16444);
nor UO_2394 (O_2394,N_19826,N_17610);
and UO_2395 (O_2395,N_18235,N_16288);
and UO_2396 (O_2396,N_17447,N_17110);
and UO_2397 (O_2397,N_18842,N_18789);
or UO_2398 (O_2398,N_19436,N_19373);
xnor UO_2399 (O_2399,N_18472,N_19483);
nor UO_2400 (O_2400,N_17001,N_19490);
and UO_2401 (O_2401,N_18819,N_18240);
nor UO_2402 (O_2402,N_16959,N_19020);
or UO_2403 (O_2403,N_16427,N_17767);
nand UO_2404 (O_2404,N_19515,N_19309);
nor UO_2405 (O_2405,N_17349,N_17762);
nor UO_2406 (O_2406,N_17254,N_19453);
or UO_2407 (O_2407,N_19072,N_19383);
nand UO_2408 (O_2408,N_17350,N_16227);
and UO_2409 (O_2409,N_16331,N_17830);
and UO_2410 (O_2410,N_16416,N_19575);
and UO_2411 (O_2411,N_18009,N_18556);
nor UO_2412 (O_2412,N_18609,N_19451);
xor UO_2413 (O_2413,N_19072,N_18677);
or UO_2414 (O_2414,N_16956,N_18231);
nor UO_2415 (O_2415,N_17265,N_16549);
or UO_2416 (O_2416,N_18630,N_19057);
nand UO_2417 (O_2417,N_18287,N_18216);
xor UO_2418 (O_2418,N_17507,N_18960);
nor UO_2419 (O_2419,N_17040,N_19629);
xor UO_2420 (O_2420,N_17864,N_17693);
or UO_2421 (O_2421,N_18760,N_19139);
xor UO_2422 (O_2422,N_19081,N_19714);
xor UO_2423 (O_2423,N_16600,N_16921);
or UO_2424 (O_2424,N_19255,N_17236);
nor UO_2425 (O_2425,N_16842,N_19698);
and UO_2426 (O_2426,N_18660,N_17380);
xor UO_2427 (O_2427,N_16585,N_18559);
xor UO_2428 (O_2428,N_16614,N_16390);
nor UO_2429 (O_2429,N_19385,N_16250);
and UO_2430 (O_2430,N_16980,N_18272);
or UO_2431 (O_2431,N_19077,N_18037);
or UO_2432 (O_2432,N_18084,N_19423);
nand UO_2433 (O_2433,N_17872,N_17797);
and UO_2434 (O_2434,N_19645,N_18438);
nor UO_2435 (O_2435,N_17726,N_17328);
xnor UO_2436 (O_2436,N_18375,N_17696);
xnor UO_2437 (O_2437,N_16647,N_18460);
nand UO_2438 (O_2438,N_18007,N_18588);
or UO_2439 (O_2439,N_19625,N_17870);
nor UO_2440 (O_2440,N_19025,N_16665);
and UO_2441 (O_2441,N_17496,N_16513);
nand UO_2442 (O_2442,N_19946,N_17421);
and UO_2443 (O_2443,N_16464,N_16937);
and UO_2444 (O_2444,N_16526,N_16786);
or UO_2445 (O_2445,N_16260,N_18280);
and UO_2446 (O_2446,N_17431,N_16057);
or UO_2447 (O_2447,N_16416,N_17032);
and UO_2448 (O_2448,N_19201,N_16497);
xor UO_2449 (O_2449,N_19796,N_17022);
nand UO_2450 (O_2450,N_16358,N_18373);
or UO_2451 (O_2451,N_17427,N_18205);
nand UO_2452 (O_2452,N_18725,N_19194);
nor UO_2453 (O_2453,N_19349,N_16899);
and UO_2454 (O_2454,N_17373,N_18240);
and UO_2455 (O_2455,N_16365,N_16805);
nand UO_2456 (O_2456,N_17202,N_18376);
nor UO_2457 (O_2457,N_19153,N_18588);
nand UO_2458 (O_2458,N_17412,N_17068);
and UO_2459 (O_2459,N_18804,N_18797);
nand UO_2460 (O_2460,N_17288,N_17928);
and UO_2461 (O_2461,N_19994,N_17834);
nor UO_2462 (O_2462,N_16993,N_19934);
xnor UO_2463 (O_2463,N_18495,N_18636);
or UO_2464 (O_2464,N_16969,N_16662);
nand UO_2465 (O_2465,N_17634,N_18505);
nand UO_2466 (O_2466,N_16659,N_18127);
and UO_2467 (O_2467,N_18111,N_18973);
or UO_2468 (O_2468,N_19454,N_17705);
or UO_2469 (O_2469,N_16072,N_19664);
and UO_2470 (O_2470,N_18640,N_16546);
nor UO_2471 (O_2471,N_17202,N_17586);
nand UO_2472 (O_2472,N_18414,N_16521);
or UO_2473 (O_2473,N_19154,N_16791);
nand UO_2474 (O_2474,N_18056,N_16708);
nor UO_2475 (O_2475,N_16702,N_19363);
nor UO_2476 (O_2476,N_19312,N_17981);
or UO_2477 (O_2477,N_18594,N_18197);
or UO_2478 (O_2478,N_18669,N_19814);
or UO_2479 (O_2479,N_17170,N_18575);
and UO_2480 (O_2480,N_17551,N_16196);
or UO_2481 (O_2481,N_16093,N_19945);
nor UO_2482 (O_2482,N_18008,N_19555);
nor UO_2483 (O_2483,N_16967,N_16761);
nand UO_2484 (O_2484,N_19002,N_19132);
nand UO_2485 (O_2485,N_19341,N_18778);
xor UO_2486 (O_2486,N_17194,N_19094);
nand UO_2487 (O_2487,N_19372,N_16554);
and UO_2488 (O_2488,N_17153,N_19557);
nand UO_2489 (O_2489,N_19879,N_17748);
or UO_2490 (O_2490,N_16139,N_19292);
nor UO_2491 (O_2491,N_19980,N_16266);
or UO_2492 (O_2492,N_17649,N_18687);
or UO_2493 (O_2493,N_19146,N_16812);
or UO_2494 (O_2494,N_19079,N_19010);
and UO_2495 (O_2495,N_17868,N_17192);
nor UO_2496 (O_2496,N_16831,N_17304);
nor UO_2497 (O_2497,N_16705,N_17661);
and UO_2498 (O_2498,N_17304,N_18614);
or UO_2499 (O_2499,N_16891,N_16511);
endmodule