module basic_500_3000_500_15_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_456,In_466);
or U1 (N_1,In_34,In_245);
xnor U2 (N_2,In_122,In_329);
and U3 (N_3,In_318,In_485);
or U4 (N_4,In_379,In_109);
nand U5 (N_5,In_413,In_461);
or U6 (N_6,In_41,In_417);
xnor U7 (N_7,In_277,In_436);
nor U8 (N_8,In_175,In_20);
nor U9 (N_9,In_234,In_160);
nor U10 (N_10,In_278,In_150);
xnor U11 (N_11,In_377,In_163);
and U12 (N_12,In_274,In_405);
nor U13 (N_13,In_83,In_291);
nor U14 (N_14,In_451,In_438);
nand U15 (N_15,In_486,In_434);
nand U16 (N_16,In_401,In_197);
or U17 (N_17,In_216,In_478);
xor U18 (N_18,In_115,In_237);
and U19 (N_19,In_118,In_67);
or U20 (N_20,In_10,In_136);
xnor U21 (N_21,In_49,In_431);
and U22 (N_22,In_368,In_251);
nand U23 (N_23,In_345,In_476);
xor U24 (N_24,In_263,In_288);
or U25 (N_25,In_130,In_71);
or U26 (N_26,In_298,In_125);
or U27 (N_27,In_454,In_248);
and U28 (N_28,In_443,In_164);
xor U29 (N_29,In_52,In_471);
or U30 (N_30,In_70,In_75);
nor U31 (N_31,In_2,In_186);
xor U32 (N_32,In_78,In_259);
xnor U33 (N_33,In_138,In_499);
xnor U34 (N_34,In_273,In_388);
xnor U35 (N_35,In_296,In_312);
nor U36 (N_36,In_253,In_261);
nand U37 (N_37,In_211,In_103);
or U38 (N_38,In_85,In_12);
nand U39 (N_39,In_188,In_190);
nor U40 (N_40,In_168,In_382);
nand U41 (N_41,In_383,In_204);
nor U42 (N_42,In_223,In_120);
or U43 (N_43,In_409,In_489);
and U44 (N_44,In_285,In_445);
and U45 (N_45,In_441,In_244);
xnor U46 (N_46,In_214,In_220);
or U47 (N_47,In_422,In_171);
nor U48 (N_48,In_396,In_384);
nand U49 (N_49,In_336,In_60);
nand U50 (N_50,In_437,In_102);
nor U51 (N_51,In_309,In_153);
nor U52 (N_52,In_411,In_386);
or U53 (N_53,In_367,In_348);
or U54 (N_54,In_217,In_205);
xnor U55 (N_55,In_300,In_177);
or U56 (N_56,In_361,In_252);
nand U57 (N_57,In_28,In_135);
nand U58 (N_58,In_77,In_376);
and U59 (N_59,In_134,In_420);
nand U60 (N_60,In_292,In_126);
nand U61 (N_61,In_395,In_293);
nor U62 (N_62,In_50,In_254);
and U63 (N_63,In_290,In_82);
nand U64 (N_64,In_469,In_106);
nor U65 (N_65,In_453,In_342);
xor U66 (N_66,In_452,In_282);
nand U67 (N_67,In_375,In_6);
or U68 (N_68,In_464,In_428);
and U69 (N_69,In_210,In_22);
nand U70 (N_70,In_238,In_398);
nor U71 (N_71,In_66,In_228);
nand U72 (N_72,In_340,In_180);
nor U73 (N_73,In_195,In_224);
or U74 (N_74,In_33,In_266);
nor U75 (N_75,In_355,In_286);
nand U76 (N_76,In_412,In_81);
or U77 (N_77,In_322,In_497);
nand U78 (N_78,In_491,In_250);
nor U79 (N_79,In_119,In_337);
nand U80 (N_80,In_339,In_13);
nand U81 (N_81,In_196,In_95);
or U82 (N_82,In_440,In_231);
or U83 (N_83,In_112,In_241);
xnor U84 (N_84,In_225,In_206);
nand U85 (N_85,In_279,In_145);
nor U86 (N_86,In_107,In_1);
xor U87 (N_87,In_25,In_450);
nand U88 (N_88,In_213,In_144);
and U89 (N_89,In_155,In_467);
xnor U90 (N_90,In_363,In_264);
or U91 (N_91,In_269,In_470);
or U92 (N_92,In_64,In_421);
nand U93 (N_93,In_330,In_480);
nor U94 (N_94,In_57,In_56);
xor U95 (N_95,In_127,In_492);
nor U96 (N_96,In_46,In_31);
nand U97 (N_97,In_68,In_199);
or U98 (N_98,In_179,In_321);
nand U99 (N_99,In_418,In_100);
and U100 (N_100,In_43,In_323);
xor U101 (N_101,In_404,In_272);
or U102 (N_102,In_47,In_333);
nor U103 (N_103,In_209,In_283);
nand U104 (N_104,In_15,In_86);
or U105 (N_105,In_328,In_27);
nor U106 (N_106,In_419,In_258);
or U107 (N_107,In_232,In_99);
and U108 (N_108,In_458,In_390);
and U109 (N_109,In_462,In_23);
and U110 (N_110,In_7,In_346);
nor U111 (N_111,In_69,In_334);
nor U112 (N_112,In_161,In_166);
nand U113 (N_113,In_202,In_146);
and U114 (N_114,In_131,In_308);
nor U115 (N_115,In_38,In_235);
xor U116 (N_116,In_193,In_257);
nor U117 (N_117,In_357,In_327);
xnor U118 (N_118,In_117,In_203);
and U119 (N_119,In_488,In_490);
or U120 (N_120,In_275,In_148);
nand U121 (N_121,In_219,In_426);
nand U122 (N_122,In_97,In_455);
or U123 (N_123,In_59,In_178);
or U124 (N_124,In_316,In_242);
nor U125 (N_125,In_63,In_372);
nor U126 (N_126,In_304,In_381);
or U127 (N_127,In_303,In_365);
nand U128 (N_128,In_37,In_65);
nor U129 (N_129,In_61,In_435);
or U130 (N_130,In_236,In_305);
xnor U131 (N_131,In_306,In_449);
nand U132 (N_132,In_338,In_494);
nand U133 (N_133,In_265,In_108);
nor U134 (N_134,In_19,In_4);
nor U135 (N_135,In_463,In_8);
and U136 (N_136,In_0,In_9);
and U137 (N_137,In_430,In_331);
xnor U138 (N_138,In_101,In_392);
nand U139 (N_139,In_397,In_221);
nor U140 (N_140,In_156,In_320);
nand U141 (N_141,In_55,In_287);
and U142 (N_142,In_18,In_89);
nand U143 (N_143,In_62,In_256);
and U144 (N_144,In_457,In_201);
or U145 (N_145,In_198,In_170);
nor U146 (N_146,In_72,In_351);
nand U147 (N_147,In_157,In_200);
and U148 (N_148,In_189,In_468);
nand U149 (N_149,In_326,In_165);
xnor U150 (N_150,In_226,In_162);
or U151 (N_151,In_460,In_92);
and U152 (N_152,In_123,In_240);
or U153 (N_153,In_76,In_104);
nand U154 (N_154,In_344,In_378);
nor U155 (N_155,In_30,In_358);
nor U156 (N_156,In_174,In_482);
and U157 (N_157,In_16,In_359);
or U158 (N_158,In_80,In_270);
or U159 (N_159,In_280,In_385);
nor U160 (N_160,In_284,In_110);
nor U161 (N_161,In_315,In_268);
or U162 (N_162,In_410,In_387);
xnor U163 (N_163,In_427,In_227);
xor U164 (N_164,In_32,In_429);
and U165 (N_165,In_230,In_142);
nor U166 (N_166,In_302,In_187);
or U167 (N_167,In_369,In_400);
or U168 (N_168,In_447,In_111);
and U169 (N_169,In_373,In_352);
nor U170 (N_170,In_218,In_424);
nor U171 (N_171,In_94,In_140);
or U172 (N_172,In_116,In_121);
or U173 (N_173,In_191,In_79);
nand U174 (N_174,In_347,In_408);
nor U175 (N_175,In_26,In_474);
nand U176 (N_176,In_173,In_393);
or U177 (N_177,In_185,In_212);
nand U178 (N_178,In_364,In_335);
nor U179 (N_179,In_149,In_132);
nor U180 (N_180,In_262,In_483);
nor U181 (N_181,In_35,In_406);
nand U182 (N_182,In_407,In_113);
nor U183 (N_183,In_446,In_444);
or U184 (N_184,In_152,In_93);
or U185 (N_185,In_301,In_24);
and U186 (N_186,In_143,In_487);
xnor U187 (N_187,In_133,In_247);
xor U188 (N_188,In_433,In_51);
xor U189 (N_189,In_481,In_394);
xor U190 (N_190,In_495,In_439);
nand U191 (N_191,In_249,In_432);
nor U192 (N_192,In_29,In_98);
nor U193 (N_193,In_313,In_229);
nor U194 (N_194,In_317,In_39);
nor U195 (N_195,In_14,In_389);
or U196 (N_196,In_183,In_151);
nor U197 (N_197,In_307,In_36);
or U198 (N_198,In_260,In_194);
nor U199 (N_199,In_128,In_356);
xnor U200 (N_200,N_116,N_146);
and U201 (N_201,In_129,N_27);
xnor U202 (N_202,N_75,N_44);
and U203 (N_203,N_150,In_448);
nand U204 (N_204,In_475,In_215);
and U205 (N_205,N_170,N_194);
or U206 (N_206,In_479,N_91);
nand U207 (N_207,N_20,N_195);
xor U208 (N_208,In_90,N_46);
nor U209 (N_209,N_74,In_222);
nor U210 (N_210,N_85,N_161);
nor U211 (N_211,N_100,In_414);
nand U212 (N_212,In_182,N_143);
or U213 (N_213,In_325,In_271);
nor U214 (N_214,In_208,N_16);
nor U215 (N_215,N_56,N_139);
or U216 (N_216,N_133,In_294);
and U217 (N_217,N_165,N_190);
xnor U218 (N_218,N_148,In_310);
xnor U219 (N_219,N_60,N_186);
or U220 (N_220,N_121,N_42);
or U221 (N_221,N_154,N_199);
and U222 (N_222,In_416,N_107);
nor U223 (N_223,N_2,In_289);
nor U224 (N_224,N_40,N_164);
and U225 (N_225,In_484,N_31);
or U226 (N_226,N_113,N_112);
xor U227 (N_227,In_276,In_91);
nor U228 (N_228,N_160,In_181);
nand U229 (N_229,In_399,N_115);
and U230 (N_230,N_159,N_106);
or U231 (N_231,In_44,N_54);
nand U232 (N_232,N_0,N_34);
xor U233 (N_233,N_55,N_39);
nand U234 (N_234,In_53,N_180);
and U235 (N_235,In_442,In_366);
nand U236 (N_236,N_38,In_243);
nor U237 (N_237,In_281,N_9);
nand U238 (N_238,In_124,N_76);
or U239 (N_239,In_341,N_128);
or U240 (N_240,N_48,N_123);
xnor U241 (N_241,N_145,N_33);
and U242 (N_242,N_108,N_96);
xnor U243 (N_243,N_64,N_131);
xor U244 (N_244,N_169,N_189);
nor U245 (N_245,N_144,N_111);
or U246 (N_246,N_187,N_1);
nand U247 (N_247,N_177,N_35);
or U248 (N_248,N_78,N_3);
or U249 (N_249,In_88,In_459);
nor U250 (N_250,In_21,N_93);
or U251 (N_251,N_7,In_477);
nor U252 (N_252,In_360,N_166);
and U253 (N_253,In_87,N_72);
or U254 (N_254,N_71,N_36);
nor U255 (N_255,N_153,N_124);
and U256 (N_256,N_43,N_191);
and U257 (N_257,N_162,N_30);
nand U258 (N_258,N_21,In_362);
nand U259 (N_259,N_151,N_126);
or U260 (N_260,N_197,N_156);
or U261 (N_261,In_391,N_32);
nand U262 (N_262,N_19,N_65);
nor U263 (N_263,N_97,N_185);
xor U264 (N_264,In_299,N_141);
and U265 (N_265,N_152,N_5);
and U266 (N_266,N_127,N_61);
or U267 (N_267,In_207,N_105);
and U268 (N_268,N_193,N_13);
and U269 (N_269,In_233,In_267);
nand U270 (N_270,N_12,In_167);
xnor U271 (N_271,In_402,N_171);
nor U272 (N_272,N_125,N_79);
xnor U273 (N_273,In_473,N_22);
nand U274 (N_274,N_119,N_69);
nand U275 (N_275,N_49,In_48);
and U276 (N_276,In_295,N_86);
and U277 (N_277,In_311,N_10);
xnor U278 (N_278,In_147,In_154);
nor U279 (N_279,In_139,In_169);
nor U280 (N_280,N_14,N_135);
or U281 (N_281,N_47,N_155);
nand U282 (N_282,N_110,N_176);
or U283 (N_283,N_41,N_62);
nand U284 (N_284,In_255,In_380);
or U285 (N_285,N_58,N_45);
or U286 (N_286,In_5,N_95);
or U287 (N_287,In_176,N_140);
and U288 (N_288,In_493,In_465);
xor U289 (N_289,N_23,N_109);
nor U290 (N_290,N_67,In_350);
or U291 (N_291,In_96,In_84);
nand U292 (N_292,In_403,N_174);
xnor U293 (N_293,In_45,In_114);
xor U294 (N_294,In_137,In_246);
xnor U295 (N_295,N_25,N_17);
xnor U296 (N_296,In_73,In_354);
and U297 (N_297,In_74,N_102);
or U298 (N_298,N_172,In_472);
xnor U299 (N_299,N_28,N_101);
nor U300 (N_300,N_15,In_58);
or U301 (N_301,N_122,In_40);
xor U302 (N_302,N_120,N_129);
nor U303 (N_303,N_68,N_114);
nor U304 (N_304,N_88,In_319);
and U305 (N_305,N_138,N_53);
xor U306 (N_306,In_54,N_163);
xnor U307 (N_307,In_158,In_159);
and U308 (N_308,In_297,N_103);
and U309 (N_309,N_188,In_498);
nor U310 (N_310,In_425,In_11);
nor U311 (N_311,N_92,N_90);
and U312 (N_312,N_157,N_63);
or U313 (N_313,In_371,N_178);
nor U314 (N_314,N_181,In_184);
nand U315 (N_315,N_184,In_374);
and U316 (N_316,N_37,N_168);
nand U317 (N_317,In_349,In_415);
or U318 (N_318,N_82,N_70);
xnor U319 (N_319,N_149,N_83);
or U320 (N_320,N_130,In_141);
xor U321 (N_321,N_136,N_198);
or U322 (N_322,In_17,N_26);
nor U323 (N_323,In_172,N_175);
xor U324 (N_324,N_11,N_104);
or U325 (N_325,In_353,N_51);
nor U326 (N_326,In_42,N_59);
or U327 (N_327,In_239,In_3);
and U328 (N_328,In_332,In_343);
or U329 (N_329,N_57,N_6);
or U330 (N_330,N_158,N_182);
and U331 (N_331,In_324,N_167);
nor U332 (N_332,In_496,N_99);
nor U333 (N_333,In_314,N_73);
or U334 (N_334,In_423,N_24);
nand U335 (N_335,N_192,N_29);
nand U336 (N_336,N_147,N_142);
nor U337 (N_337,N_98,N_137);
or U338 (N_338,N_50,N_87);
and U339 (N_339,N_8,N_183);
or U340 (N_340,N_118,N_52);
nand U341 (N_341,In_192,N_134);
nor U342 (N_342,N_89,N_80);
nor U343 (N_343,In_370,N_196);
nand U344 (N_344,N_117,N_81);
nor U345 (N_345,N_18,N_66);
and U346 (N_346,N_94,N_84);
or U347 (N_347,N_173,N_132);
xor U348 (N_348,N_179,N_77);
and U349 (N_349,In_105,N_4);
nand U350 (N_350,In_53,N_89);
nand U351 (N_351,In_311,N_92);
or U352 (N_352,N_176,N_127);
nor U353 (N_353,N_168,N_88);
nor U354 (N_354,N_99,N_178);
nand U355 (N_355,In_192,In_243);
and U356 (N_356,In_332,N_49);
nand U357 (N_357,N_30,N_70);
nand U358 (N_358,N_54,N_19);
nand U359 (N_359,N_28,N_138);
xnor U360 (N_360,N_20,In_114);
xnor U361 (N_361,In_243,N_31);
xnor U362 (N_362,N_151,N_38);
xor U363 (N_363,In_172,N_6);
and U364 (N_364,In_343,N_54);
nand U365 (N_365,In_325,N_113);
or U366 (N_366,In_299,N_35);
or U367 (N_367,N_90,N_88);
nor U368 (N_368,In_239,N_36);
nor U369 (N_369,In_353,N_95);
xor U370 (N_370,N_90,N_53);
xnor U371 (N_371,N_190,N_68);
or U372 (N_372,N_60,In_21);
or U373 (N_373,N_38,N_170);
or U374 (N_374,N_56,In_294);
xor U375 (N_375,N_197,In_281);
nor U376 (N_376,N_85,In_360);
xor U377 (N_377,In_415,N_102);
and U378 (N_378,N_48,N_13);
nor U379 (N_379,N_160,In_459);
nand U380 (N_380,N_137,N_18);
or U381 (N_381,N_153,N_3);
nand U382 (N_382,N_106,N_116);
nor U383 (N_383,N_184,In_58);
and U384 (N_384,N_12,N_68);
nor U385 (N_385,In_295,N_22);
xnor U386 (N_386,N_199,N_77);
nand U387 (N_387,N_47,In_3);
or U388 (N_388,In_139,N_113);
or U389 (N_389,N_114,N_75);
xor U390 (N_390,In_184,N_96);
nand U391 (N_391,N_183,N_128);
nand U392 (N_392,In_87,N_80);
xor U393 (N_393,N_124,N_6);
nor U394 (N_394,N_101,N_113);
nand U395 (N_395,N_26,In_370);
and U396 (N_396,In_310,N_144);
xor U397 (N_397,N_41,In_158);
nor U398 (N_398,In_496,N_120);
xor U399 (N_399,N_102,In_124);
and U400 (N_400,N_328,N_302);
nor U401 (N_401,N_329,N_232);
or U402 (N_402,N_306,N_287);
or U403 (N_403,N_259,N_363);
nor U404 (N_404,N_298,N_360);
or U405 (N_405,N_338,N_258);
xor U406 (N_406,N_309,N_289);
and U407 (N_407,N_372,N_355);
nand U408 (N_408,N_273,N_245);
nand U409 (N_409,N_284,N_205);
xnor U410 (N_410,N_223,N_394);
nor U411 (N_411,N_263,N_251);
xnor U412 (N_412,N_391,N_236);
and U413 (N_413,N_250,N_216);
nand U414 (N_414,N_370,N_343);
and U415 (N_415,N_203,N_359);
xnor U416 (N_416,N_340,N_345);
xor U417 (N_417,N_330,N_277);
nor U418 (N_418,N_389,N_367);
xor U419 (N_419,N_204,N_297);
nor U420 (N_420,N_206,N_352);
nor U421 (N_421,N_230,N_247);
and U422 (N_422,N_293,N_260);
xor U423 (N_423,N_386,N_325);
or U424 (N_424,N_337,N_333);
and U425 (N_425,N_208,N_242);
nor U426 (N_426,N_272,N_321);
or U427 (N_427,N_384,N_257);
xnor U428 (N_428,N_335,N_323);
and U429 (N_429,N_219,N_399);
or U430 (N_430,N_326,N_336);
xor U431 (N_431,N_305,N_397);
nor U432 (N_432,N_375,N_374);
xor U433 (N_433,N_316,N_310);
nor U434 (N_434,N_320,N_356);
and U435 (N_435,N_248,N_369);
or U436 (N_436,N_342,N_240);
xor U437 (N_437,N_261,N_292);
xor U438 (N_438,N_221,N_393);
nor U439 (N_439,N_398,N_392);
and U440 (N_440,N_243,N_349);
or U441 (N_441,N_315,N_358);
and U442 (N_442,N_226,N_202);
nor U443 (N_443,N_331,N_201);
or U444 (N_444,N_312,N_295);
and U445 (N_445,N_220,N_213);
and U446 (N_446,N_353,N_318);
xnor U447 (N_447,N_217,N_225);
nand U448 (N_448,N_278,N_354);
xnor U449 (N_449,N_218,N_211);
or U450 (N_450,N_348,N_314);
and U451 (N_451,N_373,N_256);
and U452 (N_452,N_366,N_351);
xnor U453 (N_453,N_347,N_299);
and U454 (N_454,N_276,N_327);
and U455 (N_455,N_210,N_291);
xor U456 (N_456,N_269,N_296);
nor U457 (N_457,N_364,N_266);
nand U458 (N_458,N_332,N_301);
nand U459 (N_459,N_241,N_308);
nand U460 (N_460,N_362,N_311);
nand U461 (N_461,N_304,N_357);
or U462 (N_462,N_285,N_267);
and U463 (N_463,N_227,N_281);
and U464 (N_464,N_390,N_239);
xor U465 (N_465,N_265,N_317);
nand U466 (N_466,N_324,N_365);
xor U467 (N_467,N_300,N_290);
and U468 (N_468,N_381,N_379);
and U469 (N_469,N_307,N_280);
or U470 (N_470,N_229,N_344);
xor U471 (N_471,N_253,N_222);
and U472 (N_472,N_255,N_234);
nor U473 (N_473,N_282,N_212);
nor U474 (N_474,N_233,N_249);
or U475 (N_475,N_224,N_254);
xnor U476 (N_476,N_380,N_275);
and U477 (N_477,N_268,N_322);
nand U478 (N_478,N_283,N_341);
nor U479 (N_479,N_368,N_319);
and U480 (N_480,N_383,N_228);
and U481 (N_481,N_252,N_334);
or U482 (N_482,N_396,N_388);
xnor U483 (N_483,N_238,N_346);
and U484 (N_484,N_279,N_274);
or U485 (N_485,N_288,N_387);
nor U486 (N_486,N_262,N_264);
and U487 (N_487,N_271,N_246);
and U488 (N_488,N_361,N_235);
or U489 (N_489,N_303,N_377);
or U490 (N_490,N_313,N_270);
xnor U491 (N_491,N_214,N_207);
nand U492 (N_492,N_231,N_385);
xnor U493 (N_493,N_339,N_382);
nand U494 (N_494,N_200,N_350);
nand U495 (N_495,N_215,N_237);
nand U496 (N_496,N_294,N_376);
and U497 (N_497,N_286,N_244);
or U498 (N_498,N_371,N_395);
and U499 (N_499,N_378,N_209);
and U500 (N_500,N_275,N_331);
nor U501 (N_501,N_265,N_301);
xnor U502 (N_502,N_326,N_206);
or U503 (N_503,N_354,N_250);
nand U504 (N_504,N_393,N_202);
and U505 (N_505,N_292,N_229);
or U506 (N_506,N_204,N_257);
nor U507 (N_507,N_297,N_390);
or U508 (N_508,N_270,N_383);
xnor U509 (N_509,N_355,N_232);
and U510 (N_510,N_360,N_243);
and U511 (N_511,N_259,N_347);
nand U512 (N_512,N_251,N_368);
nand U513 (N_513,N_285,N_259);
nor U514 (N_514,N_264,N_265);
or U515 (N_515,N_390,N_394);
nor U516 (N_516,N_320,N_377);
nor U517 (N_517,N_261,N_281);
or U518 (N_518,N_292,N_221);
and U519 (N_519,N_273,N_215);
and U520 (N_520,N_244,N_287);
xnor U521 (N_521,N_240,N_303);
nor U522 (N_522,N_383,N_333);
nand U523 (N_523,N_319,N_330);
nand U524 (N_524,N_235,N_203);
nand U525 (N_525,N_291,N_200);
or U526 (N_526,N_270,N_346);
and U527 (N_527,N_255,N_289);
and U528 (N_528,N_205,N_340);
nand U529 (N_529,N_242,N_332);
and U530 (N_530,N_228,N_311);
nor U531 (N_531,N_262,N_256);
nor U532 (N_532,N_234,N_357);
or U533 (N_533,N_239,N_201);
or U534 (N_534,N_376,N_248);
xnor U535 (N_535,N_217,N_252);
nand U536 (N_536,N_272,N_362);
nand U537 (N_537,N_324,N_233);
or U538 (N_538,N_266,N_390);
or U539 (N_539,N_223,N_386);
or U540 (N_540,N_302,N_354);
or U541 (N_541,N_365,N_309);
nand U542 (N_542,N_240,N_225);
nor U543 (N_543,N_285,N_230);
xnor U544 (N_544,N_388,N_209);
or U545 (N_545,N_276,N_301);
and U546 (N_546,N_247,N_264);
and U547 (N_547,N_281,N_203);
xnor U548 (N_548,N_247,N_297);
xnor U549 (N_549,N_387,N_304);
or U550 (N_550,N_371,N_320);
xnor U551 (N_551,N_282,N_293);
xnor U552 (N_552,N_292,N_368);
xnor U553 (N_553,N_287,N_337);
or U554 (N_554,N_299,N_226);
nor U555 (N_555,N_251,N_230);
nand U556 (N_556,N_295,N_343);
or U557 (N_557,N_236,N_381);
and U558 (N_558,N_395,N_311);
or U559 (N_559,N_323,N_262);
and U560 (N_560,N_237,N_227);
nor U561 (N_561,N_341,N_369);
and U562 (N_562,N_220,N_297);
and U563 (N_563,N_384,N_392);
nor U564 (N_564,N_350,N_358);
and U565 (N_565,N_209,N_333);
and U566 (N_566,N_319,N_266);
xor U567 (N_567,N_347,N_295);
and U568 (N_568,N_397,N_235);
and U569 (N_569,N_323,N_312);
xor U570 (N_570,N_249,N_359);
nor U571 (N_571,N_261,N_323);
nor U572 (N_572,N_212,N_327);
and U573 (N_573,N_314,N_380);
nor U574 (N_574,N_281,N_204);
and U575 (N_575,N_351,N_260);
nand U576 (N_576,N_277,N_295);
nand U577 (N_577,N_287,N_297);
nor U578 (N_578,N_307,N_266);
and U579 (N_579,N_368,N_254);
nand U580 (N_580,N_343,N_329);
or U581 (N_581,N_372,N_277);
nand U582 (N_582,N_372,N_353);
xnor U583 (N_583,N_338,N_202);
and U584 (N_584,N_287,N_313);
nor U585 (N_585,N_387,N_382);
xnor U586 (N_586,N_388,N_314);
or U587 (N_587,N_255,N_230);
and U588 (N_588,N_315,N_394);
nand U589 (N_589,N_259,N_398);
nand U590 (N_590,N_363,N_346);
or U591 (N_591,N_211,N_375);
nor U592 (N_592,N_272,N_349);
or U593 (N_593,N_311,N_284);
nand U594 (N_594,N_312,N_383);
xnor U595 (N_595,N_271,N_321);
nor U596 (N_596,N_282,N_378);
nor U597 (N_597,N_237,N_223);
nor U598 (N_598,N_308,N_356);
and U599 (N_599,N_388,N_272);
xnor U600 (N_600,N_504,N_558);
nor U601 (N_601,N_466,N_505);
nand U602 (N_602,N_525,N_544);
and U603 (N_603,N_489,N_553);
or U604 (N_604,N_542,N_408);
or U605 (N_605,N_592,N_404);
nand U606 (N_606,N_599,N_537);
nand U607 (N_607,N_502,N_469);
and U608 (N_608,N_467,N_483);
nand U609 (N_609,N_453,N_516);
nand U610 (N_610,N_501,N_488);
or U611 (N_611,N_456,N_557);
or U612 (N_612,N_470,N_519);
and U613 (N_613,N_433,N_491);
and U614 (N_614,N_430,N_411);
nor U615 (N_615,N_462,N_442);
and U616 (N_616,N_548,N_431);
xor U617 (N_617,N_515,N_568);
xnor U618 (N_618,N_561,N_421);
nor U619 (N_619,N_407,N_448);
xor U620 (N_620,N_596,N_485);
nand U621 (N_621,N_582,N_460);
xnor U622 (N_622,N_447,N_465);
nor U623 (N_623,N_487,N_598);
xor U624 (N_624,N_597,N_538);
xnor U625 (N_625,N_590,N_472);
xor U626 (N_626,N_550,N_532);
or U627 (N_627,N_530,N_443);
nand U628 (N_628,N_595,N_498);
nor U629 (N_629,N_438,N_570);
nor U630 (N_630,N_520,N_593);
nor U631 (N_631,N_510,N_482);
nor U632 (N_632,N_468,N_589);
nand U633 (N_633,N_416,N_400);
or U634 (N_634,N_512,N_534);
and U635 (N_635,N_409,N_507);
xor U636 (N_636,N_587,N_403);
or U637 (N_637,N_560,N_423);
xnor U638 (N_638,N_577,N_439);
nand U639 (N_639,N_526,N_486);
nor U640 (N_640,N_559,N_574);
nand U641 (N_641,N_579,N_541);
and U642 (N_642,N_464,N_435);
xnor U643 (N_643,N_424,N_406);
and U644 (N_644,N_440,N_539);
nand U645 (N_645,N_585,N_573);
or U646 (N_646,N_506,N_563);
and U647 (N_647,N_549,N_543);
or U648 (N_648,N_503,N_444);
nand U649 (N_649,N_449,N_547);
and U650 (N_650,N_521,N_584);
xor U651 (N_651,N_591,N_478);
and U652 (N_652,N_546,N_556);
xor U653 (N_653,N_567,N_422);
xnor U654 (N_654,N_441,N_452);
nand U655 (N_655,N_566,N_459);
nor U656 (N_656,N_564,N_457);
or U657 (N_657,N_454,N_490);
nor U658 (N_658,N_523,N_445);
and U659 (N_659,N_474,N_476);
xor U660 (N_660,N_426,N_594);
or U661 (N_661,N_529,N_481);
nand U662 (N_662,N_509,N_545);
or U663 (N_663,N_401,N_463);
nand U664 (N_664,N_533,N_496);
nand U665 (N_665,N_493,N_450);
xor U666 (N_666,N_475,N_495);
nand U667 (N_667,N_571,N_536);
nand U668 (N_668,N_517,N_551);
or U669 (N_669,N_461,N_513);
nor U670 (N_670,N_569,N_473);
xor U671 (N_671,N_522,N_511);
and U672 (N_672,N_555,N_436);
or U673 (N_673,N_576,N_554);
nor U674 (N_674,N_514,N_583);
xnor U675 (N_675,N_471,N_497);
and U676 (N_676,N_484,N_413);
or U677 (N_677,N_432,N_477);
and U678 (N_678,N_578,N_425);
xor U679 (N_679,N_580,N_572);
nor U680 (N_680,N_494,N_588);
nor U681 (N_681,N_586,N_427);
nand U682 (N_682,N_518,N_434);
xnor U683 (N_683,N_552,N_499);
nor U684 (N_684,N_437,N_540);
nor U685 (N_685,N_575,N_429);
xor U686 (N_686,N_508,N_428);
nand U687 (N_687,N_527,N_535);
and U688 (N_688,N_565,N_417);
and U689 (N_689,N_415,N_479);
xor U690 (N_690,N_562,N_405);
nand U691 (N_691,N_524,N_446);
nand U692 (N_692,N_418,N_458);
nor U693 (N_693,N_528,N_581);
and U694 (N_694,N_420,N_451);
nor U695 (N_695,N_419,N_455);
or U696 (N_696,N_480,N_414);
or U697 (N_697,N_410,N_402);
nand U698 (N_698,N_531,N_500);
nand U699 (N_699,N_492,N_412);
xor U700 (N_700,N_400,N_461);
or U701 (N_701,N_462,N_457);
or U702 (N_702,N_446,N_562);
and U703 (N_703,N_550,N_405);
or U704 (N_704,N_503,N_596);
nor U705 (N_705,N_423,N_486);
xnor U706 (N_706,N_497,N_526);
nand U707 (N_707,N_597,N_450);
nor U708 (N_708,N_415,N_587);
xor U709 (N_709,N_412,N_407);
or U710 (N_710,N_435,N_539);
and U711 (N_711,N_583,N_426);
xnor U712 (N_712,N_579,N_533);
xor U713 (N_713,N_530,N_504);
nor U714 (N_714,N_498,N_586);
nand U715 (N_715,N_498,N_594);
xnor U716 (N_716,N_457,N_547);
xor U717 (N_717,N_502,N_423);
and U718 (N_718,N_585,N_592);
xnor U719 (N_719,N_591,N_540);
nand U720 (N_720,N_492,N_497);
and U721 (N_721,N_592,N_536);
or U722 (N_722,N_408,N_459);
nor U723 (N_723,N_519,N_427);
nand U724 (N_724,N_502,N_498);
nor U725 (N_725,N_544,N_426);
nand U726 (N_726,N_581,N_597);
xor U727 (N_727,N_488,N_430);
nor U728 (N_728,N_507,N_458);
or U729 (N_729,N_555,N_425);
nor U730 (N_730,N_408,N_525);
nor U731 (N_731,N_508,N_420);
xnor U732 (N_732,N_491,N_406);
or U733 (N_733,N_403,N_412);
or U734 (N_734,N_583,N_498);
xor U735 (N_735,N_542,N_553);
or U736 (N_736,N_468,N_414);
xnor U737 (N_737,N_498,N_578);
or U738 (N_738,N_442,N_551);
nand U739 (N_739,N_493,N_587);
and U740 (N_740,N_483,N_403);
and U741 (N_741,N_573,N_478);
xnor U742 (N_742,N_578,N_559);
and U743 (N_743,N_512,N_540);
nand U744 (N_744,N_528,N_580);
xnor U745 (N_745,N_573,N_525);
nor U746 (N_746,N_578,N_469);
or U747 (N_747,N_468,N_508);
and U748 (N_748,N_413,N_490);
nor U749 (N_749,N_423,N_437);
xor U750 (N_750,N_482,N_449);
xor U751 (N_751,N_412,N_572);
or U752 (N_752,N_586,N_481);
xnor U753 (N_753,N_421,N_455);
nand U754 (N_754,N_545,N_423);
nor U755 (N_755,N_486,N_444);
and U756 (N_756,N_510,N_416);
or U757 (N_757,N_553,N_436);
nor U758 (N_758,N_563,N_559);
nor U759 (N_759,N_526,N_507);
or U760 (N_760,N_579,N_409);
xnor U761 (N_761,N_444,N_484);
and U762 (N_762,N_565,N_416);
and U763 (N_763,N_543,N_585);
nand U764 (N_764,N_454,N_421);
and U765 (N_765,N_533,N_425);
xor U766 (N_766,N_567,N_403);
or U767 (N_767,N_444,N_418);
nor U768 (N_768,N_419,N_409);
nand U769 (N_769,N_486,N_454);
and U770 (N_770,N_505,N_494);
nor U771 (N_771,N_543,N_480);
or U772 (N_772,N_585,N_504);
xnor U773 (N_773,N_457,N_490);
and U774 (N_774,N_565,N_479);
nand U775 (N_775,N_588,N_478);
and U776 (N_776,N_469,N_443);
nor U777 (N_777,N_424,N_425);
nor U778 (N_778,N_532,N_519);
xor U779 (N_779,N_493,N_552);
and U780 (N_780,N_458,N_524);
nor U781 (N_781,N_517,N_445);
nor U782 (N_782,N_575,N_511);
nand U783 (N_783,N_536,N_480);
and U784 (N_784,N_564,N_546);
nand U785 (N_785,N_542,N_554);
or U786 (N_786,N_515,N_412);
xor U787 (N_787,N_549,N_461);
xnor U788 (N_788,N_534,N_416);
and U789 (N_789,N_576,N_403);
and U790 (N_790,N_584,N_460);
nand U791 (N_791,N_485,N_533);
nor U792 (N_792,N_439,N_473);
or U793 (N_793,N_569,N_434);
xor U794 (N_794,N_528,N_540);
xnor U795 (N_795,N_565,N_570);
nand U796 (N_796,N_559,N_528);
nor U797 (N_797,N_472,N_453);
and U798 (N_798,N_534,N_453);
nand U799 (N_799,N_547,N_559);
nand U800 (N_800,N_601,N_656);
or U801 (N_801,N_772,N_713);
and U802 (N_802,N_724,N_762);
nor U803 (N_803,N_658,N_785);
and U804 (N_804,N_799,N_739);
and U805 (N_805,N_605,N_639);
or U806 (N_806,N_721,N_789);
and U807 (N_807,N_759,N_659);
and U808 (N_808,N_657,N_682);
xnor U809 (N_809,N_680,N_685);
nor U810 (N_810,N_632,N_697);
and U811 (N_811,N_769,N_652);
nand U812 (N_812,N_613,N_780);
xnor U813 (N_813,N_717,N_760);
xor U814 (N_814,N_642,N_770);
xnor U815 (N_815,N_757,N_678);
nand U816 (N_816,N_705,N_608);
and U817 (N_817,N_715,N_662);
xor U818 (N_818,N_718,N_790);
nand U819 (N_819,N_764,N_774);
or U820 (N_820,N_787,N_712);
nand U821 (N_821,N_624,N_687);
xnor U822 (N_822,N_795,N_767);
nor U823 (N_823,N_738,N_618);
xor U824 (N_824,N_711,N_645);
or U825 (N_825,N_775,N_619);
xor U826 (N_826,N_644,N_729);
nand U827 (N_827,N_754,N_751);
xnor U828 (N_828,N_796,N_782);
nand U829 (N_829,N_643,N_666);
xor U830 (N_830,N_627,N_742);
nand U831 (N_831,N_731,N_607);
nand U832 (N_832,N_745,N_623);
or U833 (N_833,N_675,N_725);
nor U834 (N_834,N_730,N_647);
xnor U835 (N_835,N_690,N_655);
nand U836 (N_836,N_746,N_600);
nor U837 (N_837,N_773,N_777);
nand U838 (N_838,N_736,N_735);
xor U839 (N_839,N_755,N_784);
xnor U840 (N_840,N_737,N_653);
or U841 (N_841,N_603,N_696);
nor U842 (N_842,N_793,N_750);
or U843 (N_843,N_672,N_708);
xnor U844 (N_844,N_681,N_701);
nand U845 (N_845,N_710,N_707);
nor U846 (N_846,N_640,N_691);
nand U847 (N_847,N_779,N_783);
or U848 (N_848,N_612,N_676);
or U849 (N_849,N_694,N_693);
nand U850 (N_850,N_668,N_788);
or U851 (N_851,N_634,N_641);
or U852 (N_852,N_752,N_768);
and U853 (N_853,N_765,N_650);
xor U854 (N_854,N_610,N_669);
nand U855 (N_855,N_665,N_631);
xnor U856 (N_856,N_673,N_741);
xor U857 (N_857,N_671,N_625);
or U858 (N_858,N_615,N_748);
xor U859 (N_859,N_700,N_633);
xor U860 (N_860,N_649,N_776);
xnor U861 (N_861,N_740,N_753);
nor U862 (N_862,N_706,N_763);
and U863 (N_863,N_670,N_621);
and U864 (N_864,N_756,N_728);
nor U865 (N_865,N_609,N_660);
xor U866 (N_866,N_692,N_626);
xnor U867 (N_867,N_630,N_704);
or U868 (N_868,N_698,N_635);
nor U869 (N_869,N_661,N_646);
or U870 (N_870,N_747,N_792);
nand U871 (N_871,N_688,N_617);
and U872 (N_872,N_667,N_614);
or U873 (N_873,N_714,N_722);
or U874 (N_874,N_604,N_791);
nand U875 (N_875,N_628,N_719);
or U876 (N_876,N_794,N_766);
or U877 (N_877,N_723,N_771);
or U878 (N_878,N_651,N_629);
and U879 (N_879,N_622,N_648);
nor U880 (N_880,N_786,N_744);
and U881 (N_881,N_720,N_636);
or U882 (N_882,N_709,N_606);
nand U883 (N_883,N_781,N_743);
or U884 (N_884,N_758,N_664);
xnor U885 (N_885,N_695,N_616);
nand U886 (N_886,N_702,N_749);
and U887 (N_887,N_732,N_637);
and U888 (N_888,N_686,N_761);
or U889 (N_889,N_734,N_674);
and U890 (N_890,N_677,N_727);
xor U891 (N_891,N_726,N_611);
and U892 (N_892,N_683,N_797);
nor U893 (N_893,N_654,N_663);
and U894 (N_894,N_798,N_684);
nor U895 (N_895,N_733,N_716);
nor U896 (N_896,N_679,N_689);
or U897 (N_897,N_699,N_638);
or U898 (N_898,N_778,N_620);
nand U899 (N_899,N_703,N_602);
nand U900 (N_900,N_626,N_724);
and U901 (N_901,N_675,N_607);
xor U902 (N_902,N_612,N_671);
nor U903 (N_903,N_602,N_754);
or U904 (N_904,N_733,N_735);
or U905 (N_905,N_684,N_627);
nor U906 (N_906,N_603,N_650);
nor U907 (N_907,N_678,N_734);
xor U908 (N_908,N_604,N_675);
xor U909 (N_909,N_791,N_640);
xor U910 (N_910,N_657,N_660);
nor U911 (N_911,N_702,N_681);
and U912 (N_912,N_604,N_676);
nand U913 (N_913,N_691,N_707);
or U914 (N_914,N_668,N_745);
xor U915 (N_915,N_771,N_741);
nand U916 (N_916,N_798,N_758);
nor U917 (N_917,N_675,N_766);
xor U918 (N_918,N_799,N_633);
xor U919 (N_919,N_639,N_723);
nor U920 (N_920,N_626,N_793);
xnor U921 (N_921,N_767,N_727);
and U922 (N_922,N_796,N_662);
and U923 (N_923,N_649,N_788);
xnor U924 (N_924,N_661,N_685);
xnor U925 (N_925,N_775,N_701);
xor U926 (N_926,N_739,N_666);
or U927 (N_927,N_679,N_775);
nand U928 (N_928,N_606,N_655);
nand U929 (N_929,N_782,N_674);
or U930 (N_930,N_694,N_715);
or U931 (N_931,N_740,N_738);
and U932 (N_932,N_674,N_743);
xnor U933 (N_933,N_683,N_698);
nor U934 (N_934,N_727,N_620);
nor U935 (N_935,N_669,N_711);
or U936 (N_936,N_762,N_726);
nand U937 (N_937,N_603,N_618);
and U938 (N_938,N_735,N_698);
xnor U939 (N_939,N_749,N_755);
xnor U940 (N_940,N_603,N_726);
or U941 (N_941,N_665,N_688);
or U942 (N_942,N_680,N_612);
xnor U943 (N_943,N_797,N_634);
nor U944 (N_944,N_736,N_707);
and U945 (N_945,N_710,N_783);
or U946 (N_946,N_765,N_753);
nand U947 (N_947,N_735,N_602);
nand U948 (N_948,N_600,N_682);
and U949 (N_949,N_727,N_718);
nor U950 (N_950,N_716,N_743);
or U951 (N_951,N_622,N_744);
nor U952 (N_952,N_658,N_698);
or U953 (N_953,N_656,N_762);
and U954 (N_954,N_779,N_786);
nand U955 (N_955,N_731,N_688);
xor U956 (N_956,N_774,N_759);
nand U957 (N_957,N_604,N_666);
nand U958 (N_958,N_653,N_799);
nand U959 (N_959,N_650,N_702);
xnor U960 (N_960,N_675,N_669);
or U961 (N_961,N_724,N_718);
and U962 (N_962,N_629,N_746);
and U963 (N_963,N_623,N_750);
xor U964 (N_964,N_681,N_666);
or U965 (N_965,N_708,N_602);
or U966 (N_966,N_672,N_742);
nand U967 (N_967,N_728,N_706);
nand U968 (N_968,N_675,N_670);
xor U969 (N_969,N_755,N_663);
nor U970 (N_970,N_669,N_690);
xor U971 (N_971,N_687,N_639);
and U972 (N_972,N_756,N_790);
and U973 (N_973,N_663,N_691);
xnor U974 (N_974,N_746,N_761);
and U975 (N_975,N_796,N_764);
or U976 (N_976,N_723,N_687);
nor U977 (N_977,N_619,N_705);
nand U978 (N_978,N_622,N_792);
xor U979 (N_979,N_658,N_776);
nor U980 (N_980,N_665,N_650);
or U981 (N_981,N_610,N_715);
or U982 (N_982,N_674,N_603);
and U983 (N_983,N_737,N_661);
and U984 (N_984,N_703,N_692);
nand U985 (N_985,N_640,N_670);
and U986 (N_986,N_680,N_652);
and U987 (N_987,N_760,N_689);
xnor U988 (N_988,N_656,N_702);
and U989 (N_989,N_763,N_640);
nand U990 (N_990,N_752,N_740);
and U991 (N_991,N_712,N_790);
and U992 (N_992,N_789,N_762);
or U993 (N_993,N_681,N_760);
or U994 (N_994,N_628,N_602);
and U995 (N_995,N_779,N_643);
or U996 (N_996,N_620,N_711);
xor U997 (N_997,N_760,N_615);
nand U998 (N_998,N_708,N_620);
xor U999 (N_999,N_740,N_680);
xor U1000 (N_1000,N_905,N_998);
xnor U1001 (N_1001,N_851,N_988);
nand U1002 (N_1002,N_857,N_999);
xor U1003 (N_1003,N_963,N_838);
nor U1004 (N_1004,N_990,N_884);
or U1005 (N_1005,N_898,N_880);
or U1006 (N_1006,N_814,N_934);
and U1007 (N_1007,N_842,N_890);
nand U1008 (N_1008,N_991,N_907);
and U1009 (N_1009,N_887,N_825);
xor U1010 (N_1010,N_941,N_967);
and U1011 (N_1011,N_989,N_981);
xor U1012 (N_1012,N_863,N_942);
or U1013 (N_1013,N_860,N_859);
xor U1014 (N_1014,N_913,N_858);
and U1015 (N_1015,N_918,N_980);
xor U1016 (N_1016,N_984,N_804);
and U1017 (N_1017,N_911,N_985);
nor U1018 (N_1018,N_862,N_928);
xnor U1019 (N_1019,N_886,N_937);
xor U1020 (N_1020,N_925,N_875);
xor U1021 (N_1021,N_943,N_926);
nor U1022 (N_1022,N_915,N_930);
nand U1023 (N_1023,N_801,N_805);
or U1024 (N_1024,N_826,N_994);
and U1025 (N_1025,N_881,N_807);
xnor U1026 (N_1026,N_987,N_960);
and U1027 (N_1027,N_955,N_818);
and U1028 (N_1028,N_840,N_982);
or U1029 (N_1029,N_876,N_891);
or U1030 (N_1030,N_979,N_836);
or U1031 (N_1031,N_929,N_953);
nand U1032 (N_1032,N_817,N_920);
xor U1033 (N_1033,N_885,N_909);
xnor U1034 (N_1034,N_802,N_971);
or U1035 (N_1035,N_945,N_902);
or U1036 (N_1036,N_978,N_908);
nand U1037 (N_1037,N_868,N_973);
and U1038 (N_1038,N_914,N_888);
nor U1039 (N_1039,N_970,N_883);
xnor U1040 (N_1040,N_869,N_940);
nand U1041 (N_1041,N_837,N_931);
or U1042 (N_1042,N_892,N_927);
xor U1043 (N_1043,N_816,N_889);
and U1044 (N_1044,N_904,N_924);
nor U1045 (N_1045,N_959,N_812);
xor U1046 (N_1046,N_993,N_906);
and U1047 (N_1047,N_835,N_871);
or U1048 (N_1048,N_939,N_899);
nor U1049 (N_1049,N_882,N_867);
or U1050 (N_1050,N_811,N_800);
nor U1051 (N_1051,N_965,N_828);
nor U1052 (N_1052,N_852,N_810);
and U1053 (N_1053,N_846,N_841);
nand U1054 (N_1054,N_866,N_827);
and U1055 (N_1055,N_831,N_933);
nor U1056 (N_1056,N_870,N_854);
nor U1057 (N_1057,N_865,N_947);
or U1058 (N_1058,N_822,N_845);
nand U1059 (N_1059,N_895,N_901);
nand U1060 (N_1060,N_820,N_938);
nor U1061 (N_1061,N_954,N_900);
nand U1062 (N_1062,N_855,N_958);
and U1063 (N_1063,N_917,N_986);
and U1064 (N_1064,N_806,N_861);
and U1065 (N_1065,N_815,N_808);
and U1066 (N_1066,N_824,N_952);
nor U1067 (N_1067,N_919,N_847);
nand U1068 (N_1068,N_813,N_946);
nand U1069 (N_1069,N_864,N_830);
xor U1070 (N_1070,N_894,N_976);
nand U1071 (N_1071,N_916,N_848);
or U1072 (N_1072,N_833,N_983);
nand U1073 (N_1073,N_856,N_956);
xnor U1074 (N_1074,N_995,N_877);
nor U1075 (N_1075,N_932,N_975);
nor U1076 (N_1076,N_873,N_910);
xor U1077 (N_1077,N_957,N_922);
and U1078 (N_1078,N_974,N_893);
or U1079 (N_1079,N_950,N_962);
xnor U1080 (N_1080,N_921,N_896);
or U1081 (N_1081,N_879,N_944);
nand U1082 (N_1082,N_843,N_969);
or U1083 (N_1083,N_966,N_897);
xnor U1084 (N_1084,N_935,N_809);
nand U1085 (N_1085,N_936,N_949);
xnor U1086 (N_1086,N_912,N_951);
nand U1087 (N_1087,N_839,N_834);
nor U1088 (N_1088,N_903,N_823);
and U1089 (N_1089,N_948,N_850);
nand U1090 (N_1090,N_844,N_849);
or U1091 (N_1091,N_972,N_997);
or U1092 (N_1092,N_977,N_878);
xnor U1093 (N_1093,N_853,N_964);
or U1094 (N_1094,N_961,N_996);
and U1095 (N_1095,N_803,N_829);
nor U1096 (N_1096,N_874,N_923);
and U1097 (N_1097,N_819,N_872);
nand U1098 (N_1098,N_992,N_968);
nor U1099 (N_1099,N_832,N_821);
nor U1100 (N_1100,N_963,N_826);
or U1101 (N_1101,N_984,N_945);
nand U1102 (N_1102,N_958,N_969);
xnor U1103 (N_1103,N_998,N_831);
nand U1104 (N_1104,N_802,N_978);
xor U1105 (N_1105,N_822,N_909);
or U1106 (N_1106,N_845,N_982);
nand U1107 (N_1107,N_913,N_952);
and U1108 (N_1108,N_921,N_962);
nand U1109 (N_1109,N_827,N_917);
or U1110 (N_1110,N_872,N_999);
xor U1111 (N_1111,N_937,N_854);
nor U1112 (N_1112,N_815,N_871);
and U1113 (N_1113,N_818,N_893);
xor U1114 (N_1114,N_873,N_977);
nand U1115 (N_1115,N_924,N_873);
xnor U1116 (N_1116,N_985,N_946);
nand U1117 (N_1117,N_941,N_932);
nand U1118 (N_1118,N_800,N_812);
or U1119 (N_1119,N_950,N_875);
and U1120 (N_1120,N_981,N_993);
or U1121 (N_1121,N_806,N_808);
xnor U1122 (N_1122,N_979,N_908);
or U1123 (N_1123,N_881,N_823);
or U1124 (N_1124,N_912,N_864);
and U1125 (N_1125,N_908,N_906);
nor U1126 (N_1126,N_957,N_867);
nand U1127 (N_1127,N_972,N_988);
nand U1128 (N_1128,N_838,N_825);
nor U1129 (N_1129,N_849,N_889);
xnor U1130 (N_1130,N_825,N_920);
and U1131 (N_1131,N_929,N_830);
or U1132 (N_1132,N_905,N_848);
nand U1133 (N_1133,N_896,N_992);
or U1134 (N_1134,N_870,N_816);
nand U1135 (N_1135,N_826,N_834);
and U1136 (N_1136,N_913,N_800);
nor U1137 (N_1137,N_907,N_835);
or U1138 (N_1138,N_856,N_894);
nor U1139 (N_1139,N_960,N_976);
or U1140 (N_1140,N_874,N_974);
nand U1141 (N_1141,N_924,N_814);
nand U1142 (N_1142,N_826,N_857);
or U1143 (N_1143,N_894,N_997);
or U1144 (N_1144,N_981,N_804);
xnor U1145 (N_1145,N_857,N_934);
and U1146 (N_1146,N_805,N_815);
nor U1147 (N_1147,N_863,N_932);
nor U1148 (N_1148,N_831,N_949);
nor U1149 (N_1149,N_857,N_850);
nor U1150 (N_1150,N_802,N_965);
or U1151 (N_1151,N_822,N_998);
nor U1152 (N_1152,N_816,N_930);
and U1153 (N_1153,N_910,N_981);
or U1154 (N_1154,N_836,N_924);
nor U1155 (N_1155,N_965,N_917);
nor U1156 (N_1156,N_806,N_914);
nand U1157 (N_1157,N_901,N_957);
xor U1158 (N_1158,N_837,N_844);
and U1159 (N_1159,N_907,N_971);
nor U1160 (N_1160,N_801,N_844);
xor U1161 (N_1161,N_870,N_960);
and U1162 (N_1162,N_889,N_934);
xor U1163 (N_1163,N_945,N_813);
xor U1164 (N_1164,N_871,N_849);
xor U1165 (N_1165,N_937,N_846);
and U1166 (N_1166,N_922,N_986);
nor U1167 (N_1167,N_961,N_875);
nor U1168 (N_1168,N_909,N_942);
and U1169 (N_1169,N_910,N_855);
nand U1170 (N_1170,N_982,N_974);
nand U1171 (N_1171,N_854,N_882);
and U1172 (N_1172,N_811,N_831);
nand U1173 (N_1173,N_811,N_820);
nand U1174 (N_1174,N_956,N_889);
nand U1175 (N_1175,N_915,N_877);
nor U1176 (N_1176,N_843,N_967);
nand U1177 (N_1177,N_856,N_837);
nand U1178 (N_1178,N_898,N_839);
or U1179 (N_1179,N_819,N_903);
nand U1180 (N_1180,N_869,N_812);
and U1181 (N_1181,N_989,N_841);
xnor U1182 (N_1182,N_920,N_824);
and U1183 (N_1183,N_813,N_835);
nor U1184 (N_1184,N_944,N_838);
and U1185 (N_1185,N_942,N_888);
and U1186 (N_1186,N_963,N_975);
or U1187 (N_1187,N_837,N_894);
xnor U1188 (N_1188,N_919,N_967);
nand U1189 (N_1189,N_917,N_968);
and U1190 (N_1190,N_819,N_834);
and U1191 (N_1191,N_996,N_905);
or U1192 (N_1192,N_882,N_887);
nand U1193 (N_1193,N_903,N_910);
and U1194 (N_1194,N_929,N_986);
xor U1195 (N_1195,N_881,N_992);
nand U1196 (N_1196,N_910,N_950);
xor U1197 (N_1197,N_816,N_912);
nand U1198 (N_1198,N_969,N_955);
or U1199 (N_1199,N_983,N_968);
xor U1200 (N_1200,N_1027,N_1046);
nor U1201 (N_1201,N_1013,N_1037);
or U1202 (N_1202,N_1001,N_1169);
and U1203 (N_1203,N_1092,N_1049);
nand U1204 (N_1204,N_1002,N_1156);
nor U1205 (N_1205,N_1026,N_1053);
and U1206 (N_1206,N_1189,N_1091);
or U1207 (N_1207,N_1021,N_1059);
or U1208 (N_1208,N_1118,N_1006);
or U1209 (N_1209,N_1095,N_1184);
nor U1210 (N_1210,N_1179,N_1009);
or U1211 (N_1211,N_1115,N_1025);
or U1212 (N_1212,N_1031,N_1044);
nand U1213 (N_1213,N_1066,N_1061);
and U1214 (N_1214,N_1101,N_1097);
and U1215 (N_1215,N_1183,N_1083);
or U1216 (N_1216,N_1073,N_1187);
nor U1217 (N_1217,N_1034,N_1174);
and U1218 (N_1218,N_1022,N_1018);
nand U1219 (N_1219,N_1178,N_1191);
and U1220 (N_1220,N_1136,N_1087);
xnor U1221 (N_1221,N_1148,N_1131);
nand U1222 (N_1222,N_1122,N_1020);
or U1223 (N_1223,N_1003,N_1150);
xnor U1224 (N_1224,N_1065,N_1038);
and U1225 (N_1225,N_1126,N_1051);
or U1226 (N_1226,N_1029,N_1048);
or U1227 (N_1227,N_1124,N_1058);
nor U1228 (N_1228,N_1099,N_1193);
xnor U1229 (N_1229,N_1180,N_1098);
nand U1230 (N_1230,N_1088,N_1120);
and U1231 (N_1231,N_1069,N_1154);
nor U1232 (N_1232,N_1062,N_1196);
or U1233 (N_1233,N_1141,N_1149);
nor U1234 (N_1234,N_1032,N_1171);
nor U1235 (N_1235,N_1033,N_1060);
and U1236 (N_1236,N_1004,N_1017);
nand U1237 (N_1237,N_1078,N_1163);
nor U1238 (N_1238,N_1182,N_1079);
nand U1239 (N_1239,N_1166,N_1103);
nand U1240 (N_1240,N_1143,N_1068);
or U1241 (N_1241,N_1192,N_1094);
and U1242 (N_1242,N_1076,N_1176);
or U1243 (N_1243,N_1137,N_1056);
or U1244 (N_1244,N_1090,N_1121);
xor U1245 (N_1245,N_1071,N_1190);
nand U1246 (N_1246,N_1055,N_1105);
nor U1247 (N_1247,N_1028,N_1085);
xor U1248 (N_1248,N_1123,N_1146);
or U1249 (N_1249,N_1015,N_1138);
xor U1250 (N_1250,N_1024,N_1054);
nand U1251 (N_1251,N_1042,N_1080);
nor U1252 (N_1252,N_1112,N_1145);
xor U1253 (N_1253,N_1139,N_1165);
nand U1254 (N_1254,N_1064,N_1155);
and U1255 (N_1255,N_1096,N_1142);
nor U1256 (N_1256,N_1070,N_1030);
nand U1257 (N_1257,N_1185,N_1111);
and U1258 (N_1258,N_1159,N_1110);
nor U1259 (N_1259,N_1106,N_1160);
nor U1260 (N_1260,N_1041,N_1140);
and U1261 (N_1261,N_1116,N_1161);
and U1262 (N_1262,N_1102,N_1043);
nor U1263 (N_1263,N_1132,N_1152);
nand U1264 (N_1264,N_1074,N_1082);
or U1265 (N_1265,N_1127,N_1075);
xor U1266 (N_1266,N_1036,N_1005);
xnor U1267 (N_1267,N_1072,N_1147);
nand U1268 (N_1268,N_1084,N_1113);
or U1269 (N_1269,N_1129,N_1135);
xor U1270 (N_1270,N_1063,N_1186);
nor U1271 (N_1271,N_1057,N_1039);
nand U1272 (N_1272,N_1012,N_1130);
or U1273 (N_1273,N_1119,N_1162);
nor U1274 (N_1274,N_1107,N_1047);
and U1275 (N_1275,N_1194,N_1023);
nand U1276 (N_1276,N_1164,N_1195);
nor U1277 (N_1277,N_1168,N_1198);
nand U1278 (N_1278,N_1077,N_1016);
nor U1279 (N_1279,N_1114,N_1007);
nand U1280 (N_1280,N_1011,N_1167);
and U1281 (N_1281,N_1081,N_1067);
or U1282 (N_1282,N_1104,N_1125);
and U1283 (N_1283,N_1117,N_1175);
xor U1284 (N_1284,N_1108,N_1153);
or U1285 (N_1285,N_1158,N_1014);
and U1286 (N_1286,N_1008,N_1086);
and U1287 (N_1287,N_1109,N_1093);
and U1288 (N_1288,N_1100,N_1172);
and U1289 (N_1289,N_1019,N_1050);
and U1290 (N_1290,N_1199,N_1089);
nor U1291 (N_1291,N_1010,N_1170);
nor U1292 (N_1292,N_1173,N_1045);
nor U1293 (N_1293,N_1188,N_1181);
nor U1294 (N_1294,N_1035,N_1128);
xor U1295 (N_1295,N_1157,N_1000);
and U1296 (N_1296,N_1134,N_1133);
and U1297 (N_1297,N_1052,N_1197);
nand U1298 (N_1298,N_1144,N_1151);
nor U1299 (N_1299,N_1040,N_1177);
xor U1300 (N_1300,N_1032,N_1096);
xnor U1301 (N_1301,N_1108,N_1152);
nor U1302 (N_1302,N_1061,N_1108);
nand U1303 (N_1303,N_1042,N_1112);
nand U1304 (N_1304,N_1064,N_1154);
xor U1305 (N_1305,N_1126,N_1133);
nor U1306 (N_1306,N_1001,N_1040);
and U1307 (N_1307,N_1128,N_1194);
and U1308 (N_1308,N_1118,N_1095);
or U1309 (N_1309,N_1092,N_1175);
or U1310 (N_1310,N_1058,N_1012);
or U1311 (N_1311,N_1096,N_1198);
nor U1312 (N_1312,N_1083,N_1071);
nand U1313 (N_1313,N_1063,N_1154);
xor U1314 (N_1314,N_1089,N_1166);
nand U1315 (N_1315,N_1126,N_1146);
and U1316 (N_1316,N_1125,N_1059);
nand U1317 (N_1317,N_1114,N_1148);
nand U1318 (N_1318,N_1135,N_1150);
nor U1319 (N_1319,N_1126,N_1122);
xnor U1320 (N_1320,N_1061,N_1055);
nor U1321 (N_1321,N_1000,N_1024);
or U1322 (N_1322,N_1125,N_1026);
nor U1323 (N_1323,N_1196,N_1109);
and U1324 (N_1324,N_1025,N_1175);
nor U1325 (N_1325,N_1171,N_1042);
nor U1326 (N_1326,N_1173,N_1085);
nor U1327 (N_1327,N_1047,N_1119);
nand U1328 (N_1328,N_1089,N_1063);
nor U1329 (N_1329,N_1071,N_1014);
and U1330 (N_1330,N_1133,N_1148);
xor U1331 (N_1331,N_1133,N_1041);
xnor U1332 (N_1332,N_1063,N_1037);
and U1333 (N_1333,N_1044,N_1095);
and U1334 (N_1334,N_1013,N_1147);
xor U1335 (N_1335,N_1135,N_1147);
nor U1336 (N_1336,N_1080,N_1046);
xor U1337 (N_1337,N_1185,N_1193);
xor U1338 (N_1338,N_1016,N_1095);
and U1339 (N_1339,N_1195,N_1018);
xor U1340 (N_1340,N_1066,N_1121);
nand U1341 (N_1341,N_1119,N_1055);
nor U1342 (N_1342,N_1075,N_1109);
xor U1343 (N_1343,N_1136,N_1014);
nand U1344 (N_1344,N_1141,N_1073);
and U1345 (N_1345,N_1175,N_1021);
nand U1346 (N_1346,N_1142,N_1037);
or U1347 (N_1347,N_1043,N_1025);
nor U1348 (N_1348,N_1066,N_1030);
xor U1349 (N_1349,N_1029,N_1109);
xor U1350 (N_1350,N_1057,N_1198);
nand U1351 (N_1351,N_1000,N_1152);
or U1352 (N_1352,N_1033,N_1075);
nand U1353 (N_1353,N_1059,N_1090);
and U1354 (N_1354,N_1099,N_1027);
nand U1355 (N_1355,N_1041,N_1151);
and U1356 (N_1356,N_1189,N_1135);
xor U1357 (N_1357,N_1040,N_1062);
or U1358 (N_1358,N_1099,N_1144);
nor U1359 (N_1359,N_1051,N_1123);
nand U1360 (N_1360,N_1060,N_1053);
and U1361 (N_1361,N_1068,N_1193);
xor U1362 (N_1362,N_1159,N_1073);
xor U1363 (N_1363,N_1091,N_1108);
and U1364 (N_1364,N_1189,N_1092);
or U1365 (N_1365,N_1015,N_1074);
and U1366 (N_1366,N_1142,N_1023);
xor U1367 (N_1367,N_1138,N_1067);
and U1368 (N_1368,N_1150,N_1045);
or U1369 (N_1369,N_1153,N_1005);
nor U1370 (N_1370,N_1044,N_1098);
nor U1371 (N_1371,N_1183,N_1153);
xnor U1372 (N_1372,N_1180,N_1017);
and U1373 (N_1373,N_1148,N_1109);
nor U1374 (N_1374,N_1076,N_1170);
xor U1375 (N_1375,N_1023,N_1077);
nor U1376 (N_1376,N_1191,N_1137);
xor U1377 (N_1377,N_1003,N_1015);
and U1378 (N_1378,N_1015,N_1109);
xor U1379 (N_1379,N_1062,N_1051);
nor U1380 (N_1380,N_1005,N_1126);
nand U1381 (N_1381,N_1177,N_1159);
xor U1382 (N_1382,N_1128,N_1013);
and U1383 (N_1383,N_1188,N_1047);
or U1384 (N_1384,N_1024,N_1115);
and U1385 (N_1385,N_1007,N_1018);
nor U1386 (N_1386,N_1067,N_1073);
xor U1387 (N_1387,N_1079,N_1074);
or U1388 (N_1388,N_1140,N_1171);
nand U1389 (N_1389,N_1142,N_1155);
or U1390 (N_1390,N_1195,N_1066);
xnor U1391 (N_1391,N_1054,N_1175);
nand U1392 (N_1392,N_1114,N_1022);
xnor U1393 (N_1393,N_1161,N_1008);
or U1394 (N_1394,N_1122,N_1125);
nor U1395 (N_1395,N_1022,N_1078);
or U1396 (N_1396,N_1041,N_1123);
or U1397 (N_1397,N_1082,N_1064);
and U1398 (N_1398,N_1000,N_1037);
or U1399 (N_1399,N_1107,N_1098);
nand U1400 (N_1400,N_1281,N_1274);
or U1401 (N_1401,N_1299,N_1385);
nor U1402 (N_1402,N_1354,N_1217);
or U1403 (N_1403,N_1267,N_1209);
nor U1404 (N_1404,N_1329,N_1263);
nor U1405 (N_1405,N_1357,N_1353);
and U1406 (N_1406,N_1365,N_1356);
nand U1407 (N_1407,N_1204,N_1202);
nand U1408 (N_1408,N_1320,N_1399);
xnor U1409 (N_1409,N_1344,N_1250);
nand U1410 (N_1410,N_1283,N_1397);
nand U1411 (N_1411,N_1291,N_1215);
xnor U1412 (N_1412,N_1296,N_1386);
xor U1413 (N_1413,N_1301,N_1315);
or U1414 (N_1414,N_1242,N_1312);
or U1415 (N_1415,N_1280,N_1286);
or U1416 (N_1416,N_1245,N_1335);
xor U1417 (N_1417,N_1359,N_1216);
nand U1418 (N_1418,N_1232,N_1363);
and U1419 (N_1419,N_1393,N_1225);
nor U1420 (N_1420,N_1241,N_1364);
xor U1421 (N_1421,N_1278,N_1224);
nand U1422 (N_1422,N_1307,N_1244);
or U1423 (N_1423,N_1268,N_1310);
nor U1424 (N_1424,N_1265,N_1379);
nand U1425 (N_1425,N_1302,N_1297);
and U1426 (N_1426,N_1380,N_1208);
xor U1427 (N_1427,N_1340,N_1201);
xnor U1428 (N_1428,N_1259,N_1270);
nand U1429 (N_1429,N_1279,N_1210);
nand U1430 (N_1430,N_1228,N_1309);
nor U1431 (N_1431,N_1377,N_1257);
nand U1432 (N_1432,N_1346,N_1308);
or U1433 (N_1433,N_1237,N_1262);
xor U1434 (N_1434,N_1375,N_1321);
nand U1435 (N_1435,N_1243,N_1369);
nand U1436 (N_1436,N_1342,N_1230);
nand U1437 (N_1437,N_1395,N_1254);
xnor U1438 (N_1438,N_1205,N_1366);
or U1439 (N_1439,N_1390,N_1227);
xor U1440 (N_1440,N_1392,N_1258);
nand U1441 (N_1441,N_1349,N_1277);
nand U1442 (N_1442,N_1388,N_1298);
xnor U1443 (N_1443,N_1371,N_1347);
nor U1444 (N_1444,N_1269,N_1367);
nor U1445 (N_1445,N_1213,N_1292);
and U1446 (N_1446,N_1207,N_1287);
nand U1447 (N_1447,N_1285,N_1255);
and U1448 (N_1448,N_1361,N_1239);
and U1449 (N_1449,N_1249,N_1222);
and U1450 (N_1450,N_1317,N_1341);
or U1451 (N_1451,N_1331,N_1384);
nor U1452 (N_1452,N_1373,N_1294);
xor U1453 (N_1453,N_1271,N_1398);
and U1454 (N_1454,N_1251,N_1260);
nor U1455 (N_1455,N_1305,N_1328);
and U1456 (N_1456,N_1229,N_1374);
nor U1457 (N_1457,N_1330,N_1368);
nor U1458 (N_1458,N_1389,N_1355);
nor U1459 (N_1459,N_1226,N_1358);
and U1460 (N_1460,N_1236,N_1326);
nor U1461 (N_1461,N_1334,N_1360);
nor U1462 (N_1462,N_1246,N_1345);
nand U1463 (N_1463,N_1219,N_1333);
nor U1464 (N_1464,N_1240,N_1289);
or U1465 (N_1465,N_1235,N_1275);
xnor U1466 (N_1466,N_1221,N_1276);
nor U1467 (N_1467,N_1378,N_1247);
xor U1468 (N_1468,N_1256,N_1382);
nor U1469 (N_1469,N_1206,N_1212);
and U1470 (N_1470,N_1322,N_1314);
nand U1471 (N_1471,N_1383,N_1273);
nand U1472 (N_1472,N_1253,N_1327);
nand U1473 (N_1473,N_1282,N_1352);
or U1474 (N_1474,N_1372,N_1200);
xnor U1475 (N_1475,N_1348,N_1223);
or U1476 (N_1476,N_1376,N_1214);
or U1477 (N_1477,N_1233,N_1304);
nand U1478 (N_1478,N_1338,N_1303);
nor U1479 (N_1479,N_1284,N_1211);
nand U1480 (N_1480,N_1306,N_1325);
xor U1481 (N_1481,N_1351,N_1391);
or U1482 (N_1482,N_1316,N_1323);
nor U1483 (N_1483,N_1266,N_1252);
nor U1484 (N_1484,N_1220,N_1264);
and U1485 (N_1485,N_1324,N_1381);
nand U1486 (N_1486,N_1231,N_1288);
nor U1487 (N_1487,N_1218,N_1295);
xnor U1488 (N_1488,N_1336,N_1238);
xnor U1489 (N_1489,N_1313,N_1203);
nand U1490 (N_1490,N_1248,N_1337);
or U1491 (N_1491,N_1290,N_1332);
and U1492 (N_1492,N_1261,N_1339);
and U1493 (N_1493,N_1350,N_1293);
nor U1494 (N_1494,N_1370,N_1318);
xor U1495 (N_1495,N_1387,N_1272);
or U1496 (N_1496,N_1311,N_1394);
and U1497 (N_1497,N_1362,N_1343);
or U1498 (N_1498,N_1319,N_1396);
and U1499 (N_1499,N_1234,N_1300);
nor U1500 (N_1500,N_1388,N_1346);
nor U1501 (N_1501,N_1254,N_1271);
xnor U1502 (N_1502,N_1347,N_1399);
xor U1503 (N_1503,N_1215,N_1370);
nand U1504 (N_1504,N_1315,N_1265);
xnor U1505 (N_1505,N_1356,N_1363);
nor U1506 (N_1506,N_1357,N_1302);
and U1507 (N_1507,N_1332,N_1352);
and U1508 (N_1508,N_1233,N_1391);
or U1509 (N_1509,N_1384,N_1388);
nor U1510 (N_1510,N_1230,N_1253);
and U1511 (N_1511,N_1377,N_1329);
nand U1512 (N_1512,N_1322,N_1270);
and U1513 (N_1513,N_1296,N_1226);
nor U1514 (N_1514,N_1381,N_1338);
or U1515 (N_1515,N_1367,N_1206);
and U1516 (N_1516,N_1391,N_1239);
xnor U1517 (N_1517,N_1258,N_1254);
or U1518 (N_1518,N_1264,N_1242);
nand U1519 (N_1519,N_1294,N_1291);
nand U1520 (N_1520,N_1296,N_1287);
xnor U1521 (N_1521,N_1349,N_1363);
nor U1522 (N_1522,N_1242,N_1223);
and U1523 (N_1523,N_1274,N_1224);
xnor U1524 (N_1524,N_1214,N_1375);
and U1525 (N_1525,N_1371,N_1379);
nor U1526 (N_1526,N_1395,N_1315);
nor U1527 (N_1527,N_1227,N_1374);
and U1528 (N_1528,N_1392,N_1305);
or U1529 (N_1529,N_1253,N_1351);
xor U1530 (N_1530,N_1339,N_1349);
xor U1531 (N_1531,N_1276,N_1393);
nand U1532 (N_1532,N_1346,N_1303);
nor U1533 (N_1533,N_1342,N_1341);
nor U1534 (N_1534,N_1291,N_1354);
and U1535 (N_1535,N_1312,N_1371);
nor U1536 (N_1536,N_1256,N_1351);
xnor U1537 (N_1537,N_1343,N_1254);
or U1538 (N_1538,N_1208,N_1205);
or U1539 (N_1539,N_1302,N_1381);
nor U1540 (N_1540,N_1319,N_1264);
nand U1541 (N_1541,N_1293,N_1314);
nand U1542 (N_1542,N_1224,N_1320);
and U1543 (N_1543,N_1281,N_1395);
nor U1544 (N_1544,N_1364,N_1396);
nand U1545 (N_1545,N_1340,N_1324);
nand U1546 (N_1546,N_1204,N_1390);
xnor U1547 (N_1547,N_1309,N_1285);
and U1548 (N_1548,N_1280,N_1203);
nand U1549 (N_1549,N_1273,N_1375);
and U1550 (N_1550,N_1355,N_1381);
or U1551 (N_1551,N_1322,N_1356);
and U1552 (N_1552,N_1334,N_1293);
and U1553 (N_1553,N_1325,N_1339);
nor U1554 (N_1554,N_1349,N_1357);
xnor U1555 (N_1555,N_1252,N_1274);
xnor U1556 (N_1556,N_1263,N_1226);
nand U1557 (N_1557,N_1223,N_1344);
and U1558 (N_1558,N_1283,N_1307);
and U1559 (N_1559,N_1206,N_1329);
and U1560 (N_1560,N_1273,N_1390);
and U1561 (N_1561,N_1326,N_1310);
xnor U1562 (N_1562,N_1349,N_1218);
nor U1563 (N_1563,N_1251,N_1277);
or U1564 (N_1564,N_1252,N_1289);
nand U1565 (N_1565,N_1227,N_1332);
nand U1566 (N_1566,N_1381,N_1349);
and U1567 (N_1567,N_1313,N_1311);
and U1568 (N_1568,N_1277,N_1255);
nor U1569 (N_1569,N_1241,N_1333);
nand U1570 (N_1570,N_1217,N_1254);
and U1571 (N_1571,N_1213,N_1296);
xor U1572 (N_1572,N_1216,N_1295);
and U1573 (N_1573,N_1368,N_1393);
nor U1574 (N_1574,N_1377,N_1244);
nor U1575 (N_1575,N_1359,N_1268);
nor U1576 (N_1576,N_1318,N_1269);
nand U1577 (N_1577,N_1391,N_1263);
xnor U1578 (N_1578,N_1288,N_1311);
xnor U1579 (N_1579,N_1297,N_1389);
xor U1580 (N_1580,N_1267,N_1275);
xnor U1581 (N_1581,N_1351,N_1393);
or U1582 (N_1582,N_1391,N_1200);
and U1583 (N_1583,N_1311,N_1310);
xor U1584 (N_1584,N_1338,N_1208);
nor U1585 (N_1585,N_1254,N_1380);
or U1586 (N_1586,N_1299,N_1297);
or U1587 (N_1587,N_1225,N_1307);
nand U1588 (N_1588,N_1291,N_1247);
or U1589 (N_1589,N_1275,N_1341);
nor U1590 (N_1590,N_1358,N_1300);
or U1591 (N_1591,N_1331,N_1222);
and U1592 (N_1592,N_1345,N_1285);
nor U1593 (N_1593,N_1380,N_1384);
nor U1594 (N_1594,N_1269,N_1231);
nand U1595 (N_1595,N_1353,N_1267);
nor U1596 (N_1596,N_1352,N_1296);
and U1597 (N_1597,N_1212,N_1205);
or U1598 (N_1598,N_1262,N_1327);
nand U1599 (N_1599,N_1293,N_1355);
or U1600 (N_1600,N_1515,N_1556);
and U1601 (N_1601,N_1590,N_1406);
nor U1602 (N_1602,N_1518,N_1433);
xnor U1603 (N_1603,N_1534,N_1510);
xnor U1604 (N_1604,N_1582,N_1593);
nand U1605 (N_1605,N_1524,N_1455);
and U1606 (N_1606,N_1527,N_1559);
and U1607 (N_1607,N_1594,N_1564);
or U1608 (N_1608,N_1544,N_1588);
nand U1609 (N_1609,N_1494,N_1554);
nor U1610 (N_1610,N_1415,N_1408);
or U1611 (N_1611,N_1569,N_1597);
and U1612 (N_1612,N_1472,N_1499);
and U1613 (N_1613,N_1540,N_1439);
xnor U1614 (N_1614,N_1587,N_1574);
xor U1615 (N_1615,N_1501,N_1427);
nor U1616 (N_1616,N_1589,N_1416);
and U1617 (N_1617,N_1419,N_1407);
nor U1618 (N_1618,N_1467,N_1577);
nor U1619 (N_1619,N_1557,N_1443);
and U1620 (N_1620,N_1478,N_1424);
and U1621 (N_1621,N_1592,N_1461);
nand U1622 (N_1622,N_1521,N_1573);
nor U1623 (N_1623,N_1413,N_1579);
xnor U1624 (N_1624,N_1532,N_1476);
xnor U1625 (N_1625,N_1570,N_1481);
nand U1626 (N_1626,N_1418,N_1500);
or U1627 (N_1627,N_1450,N_1549);
xnor U1628 (N_1628,N_1405,N_1451);
or U1629 (N_1629,N_1580,N_1517);
nor U1630 (N_1630,N_1487,N_1551);
xor U1631 (N_1631,N_1462,N_1565);
and U1632 (N_1632,N_1493,N_1447);
xnor U1633 (N_1633,N_1507,N_1548);
and U1634 (N_1634,N_1545,N_1585);
and U1635 (N_1635,N_1552,N_1446);
or U1636 (N_1636,N_1411,N_1508);
and U1637 (N_1637,N_1420,N_1509);
xor U1638 (N_1638,N_1529,N_1505);
or U1639 (N_1639,N_1452,N_1536);
nand U1640 (N_1640,N_1562,N_1488);
xor U1641 (N_1641,N_1444,N_1463);
nand U1642 (N_1642,N_1595,N_1578);
nand U1643 (N_1643,N_1563,N_1550);
or U1644 (N_1644,N_1586,N_1568);
xnor U1645 (N_1645,N_1566,N_1437);
nor U1646 (N_1646,N_1464,N_1560);
nor U1647 (N_1647,N_1471,N_1543);
xnor U1648 (N_1648,N_1449,N_1403);
xor U1649 (N_1649,N_1466,N_1438);
nand U1650 (N_1650,N_1504,N_1440);
or U1651 (N_1651,N_1465,N_1489);
nand U1652 (N_1652,N_1567,N_1538);
or U1653 (N_1653,N_1409,N_1547);
nand U1654 (N_1654,N_1520,N_1445);
nand U1655 (N_1655,N_1474,N_1404);
xor U1656 (N_1656,N_1441,N_1460);
nand U1657 (N_1657,N_1486,N_1583);
xor U1658 (N_1658,N_1533,N_1470);
and U1659 (N_1659,N_1485,N_1414);
and U1660 (N_1660,N_1448,N_1581);
or U1661 (N_1661,N_1459,N_1410);
xor U1662 (N_1662,N_1596,N_1442);
or U1663 (N_1663,N_1571,N_1513);
nand U1664 (N_1664,N_1553,N_1599);
and U1665 (N_1665,N_1541,N_1400);
or U1666 (N_1666,N_1435,N_1456);
nor U1667 (N_1667,N_1561,N_1555);
and U1668 (N_1668,N_1576,N_1512);
nor U1669 (N_1669,N_1469,N_1482);
nor U1670 (N_1670,N_1425,N_1572);
nand U1671 (N_1671,N_1598,N_1480);
nor U1672 (N_1672,N_1496,N_1483);
nand U1673 (N_1673,N_1584,N_1523);
and U1674 (N_1674,N_1475,N_1436);
nand U1675 (N_1675,N_1511,N_1422);
and U1676 (N_1676,N_1495,N_1522);
or U1677 (N_1677,N_1490,N_1498);
or U1678 (N_1678,N_1531,N_1497);
or U1679 (N_1679,N_1492,N_1454);
or U1680 (N_1680,N_1434,N_1539);
nand U1681 (N_1681,N_1412,N_1401);
nand U1682 (N_1682,N_1421,N_1546);
and U1683 (N_1683,N_1591,N_1506);
nor U1684 (N_1684,N_1432,N_1468);
nor U1685 (N_1685,N_1473,N_1519);
nand U1686 (N_1686,N_1428,N_1484);
or U1687 (N_1687,N_1503,N_1491);
or U1688 (N_1688,N_1402,N_1525);
and U1689 (N_1689,N_1516,N_1453);
and U1690 (N_1690,N_1457,N_1575);
xnor U1691 (N_1691,N_1479,N_1502);
nor U1692 (N_1692,N_1535,N_1558);
or U1693 (N_1693,N_1417,N_1431);
xor U1694 (N_1694,N_1429,N_1528);
nand U1695 (N_1695,N_1514,N_1526);
nand U1696 (N_1696,N_1530,N_1477);
nand U1697 (N_1697,N_1458,N_1430);
nor U1698 (N_1698,N_1426,N_1537);
nor U1699 (N_1699,N_1542,N_1423);
or U1700 (N_1700,N_1513,N_1439);
and U1701 (N_1701,N_1596,N_1507);
or U1702 (N_1702,N_1503,N_1564);
and U1703 (N_1703,N_1503,N_1401);
or U1704 (N_1704,N_1441,N_1419);
nand U1705 (N_1705,N_1585,N_1487);
or U1706 (N_1706,N_1461,N_1544);
and U1707 (N_1707,N_1401,N_1545);
xnor U1708 (N_1708,N_1552,N_1510);
nor U1709 (N_1709,N_1508,N_1424);
or U1710 (N_1710,N_1499,N_1577);
xnor U1711 (N_1711,N_1509,N_1406);
and U1712 (N_1712,N_1506,N_1470);
xor U1713 (N_1713,N_1446,N_1525);
nor U1714 (N_1714,N_1540,N_1511);
nand U1715 (N_1715,N_1597,N_1559);
and U1716 (N_1716,N_1536,N_1445);
nor U1717 (N_1717,N_1486,N_1558);
nand U1718 (N_1718,N_1487,N_1507);
nand U1719 (N_1719,N_1467,N_1489);
nor U1720 (N_1720,N_1474,N_1566);
nand U1721 (N_1721,N_1506,N_1564);
nor U1722 (N_1722,N_1583,N_1570);
and U1723 (N_1723,N_1565,N_1468);
or U1724 (N_1724,N_1461,N_1454);
or U1725 (N_1725,N_1470,N_1588);
and U1726 (N_1726,N_1478,N_1493);
nand U1727 (N_1727,N_1489,N_1444);
xnor U1728 (N_1728,N_1487,N_1503);
xnor U1729 (N_1729,N_1563,N_1551);
xnor U1730 (N_1730,N_1515,N_1490);
or U1731 (N_1731,N_1422,N_1408);
and U1732 (N_1732,N_1525,N_1537);
xor U1733 (N_1733,N_1407,N_1569);
nor U1734 (N_1734,N_1482,N_1522);
or U1735 (N_1735,N_1544,N_1545);
nand U1736 (N_1736,N_1438,N_1570);
or U1737 (N_1737,N_1446,N_1417);
nor U1738 (N_1738,N_1546,N_1410);
or U1739 (N_1739,N_1466,N_1450);
nand U1740 (N_1740,N_1456,N_1541);
and U1741 (N_1741,N_1577,N_1490);
and U1742 (N_1742,N_1557,N_1450);
nor U1743 (N_1743,N_1403,N_1585);
nor U1744 (N_1744,N_1540,N_1455);
nor U1745 (N_1745,N_1481,N_1449);
nor U1746 (N_1746,N_1471,N_1594);
nand U1747 (N_1747,N_1469,N_1417);
nor U1748 (N_1748,N_1574,N_1591);
or U1749 (N_1749,N_1447,N_1500);
or U1750 (N_1750,N_1413,N_1542);
nor U1751 (N_1751,N_1416,N_1575);
or U1752 (N_1752,N_1502,N_1469);
xnor U1753 (N_1753,N_1418,N_1411);
or U1754 (N_1754,N_1432,N_1539);
nor U1755 (N_1755,N_1566,N_1524);
or U1756 (N_1756,N_1517,N_1463);
and U1757 (N_1757,N_1404,N_1472);
nor U1758 (N_1758,N_1486,N_1508);
xnor U1759 (N_1759,N_1526,N_1400);
and U1760 (N_1760,N_1518,N_1427);
nor U1761 (N_1761,N_1484,N_1552);
or U1762 (N_1762,N_1599,N_1501);
or U1763 (N_1763,N_1493,N_1509);
and U1764 (N_1764,N_1424,N_1540);
nand U1765 (N_1765,N_1495,N_1408);
nand U1766 (N_1766,N_1526,N_1421);
nand U1767 (N_1767,N_1541,N_1523);
nand U1768 (N_1768,N_1403,N_1481);
and U1769 (N_1769,N_1492,N_1517);
nor U1770 (N_1770,N_1595,N_1516);
or U1771 (N_1771,N_1572,N_1560);
xor U1772 (N_1772,N_1456,N_1540);
or U1773 (N_1773,N_1491,N_1415);
xnor U1774 (N_1774,N_1595,N_1506);
xnor U1775 (N_1775,N_1495,N_1437);
and U1776 (N_1776,N_1487,N_1543);
and U1777 (N_1777,N_1452,N_1488);
nand U1778 (N_1778,N_1548,N_1435);
xor U1779 (N_1779,N_1557,N_1492);
xnor U1780 (N_1780,N_1414,N_1541);
xor U1781 (N_1781,N_1510,N_1554);
xnor U1782 (N_1782,N_1502,N_1406);
nand U1783 (N_1783,N_1551,N_1472);
nor U1784 (N_1784,N_1405,N_1481);
and U1785 (N_1785,N_1538,N_1486);
xor U1786 (N_1786,N_1579,N_1531);
nor U1787 (N_1787,N_1539,N_1529);
nor U1788 (N_1788,N_1496,N_1561);
or U1789 (N_1789,N_1443,N_1534);
nor U1790 (N_1790,N_1548,N_1452);
nor U1791 (N_1791,N_1450,N_1480);
and U1792 (N_1792,N_1558,N_1420);
nor U1793 (N_1793,N_1520,N_1578);
and U1794 (N_1794,N_1441,N_1527);
and U1795 (N_1795,N_1568,N_1557);
xnor U1796 (N_1796,N_1569,N_1413);
nand U1797 (N_1797,N_1565,N_1438);
or U1798 (N_1798,N_1483,N_1417);
nor U1799 (N_1799,N_1428,N_1567);
nor U1800 (N_1800,N_1775,N_1719);
nand U1801 (N_1801,N_1689,N_1777);
nor U1802 (N_1802,N_1746,N_1743);
or U1803 (N_1803,N_1625,N_1774);
and U1804 (N_1804,N_1616,N_1609);
xor U1805 (N_1805,N_1704,N_1659);
xnor U1806 (N_1806,N_1601,N_1748);
and U1807 (N_1807,N_1769,N_1607);
and U1808 (N_1808,N_1685,N_1669);
or U1809 (N_1809,N_1720,N_1649);
and U1810 (N_1810,N_1631,N_1718);
and U1811 (N_1811,N_1650,N_1670);
xor U1812 (N_1812,N_1660,N_1683);
nand U1813 (N_1813,N_1796,N_1657);
xor U1814 (N_1814,N_1639,N_1733);
nor U1815 (N_1815,N_1641,N_1768);
nand U1816 (N_1816,N_1739,N_1725);
or U1817 (N_1817,N_1687,N_1658);
or U1818 (N_1818,N_1716,N_1765);
or U1819 (N_1819,N_1708,N_1622);
nand U1820 (N_1820,N_1723,N_1643);
nand U1821 (N_1821,N_1766,N_1724);
and U1822 (N_1822,N_1737,N_1706);
or U1823 (N_1823,N_1705,N_1792);
nor U1824 (N_1824,N_1773,N_1675);
and U1825 (N_1825,N_1744,N_1754);
nor U1826 (N_1826,N_1624,N_1656);
nor U1827 (N_1827,N_1772,N_1612);
and U1828 (N_1828,N_1654,N_1617);
or U1829 (N_1829,N_1789,N_1700);
xor U1830 (N_1830,N_1721,N_1647);
nand U1831 (N_1831,N_1699,N_1740);
nand U1832 (N_1832,N_1608,N_1782);
nor U1833 (N_1833,N_1715,N_1735);
and U1834 (N_1834,N_1759,N_1613);
xor U1835 (N_1835,N_1637,N_1666);
nand U1836 (N_1836,N_1747,N_1711);
xnor U1837 (N_1837,N_1651,N_1696);
xnor U1838 (N_1838,N_1640,N_1606);
nor U1839 (N_1839,N_1776,N_1729);
nand U1840 (N_1840,N_1620,N_1652);
or U1841 (N_1841,N_1684,N_1605);
or U1842 (N_1842,N_1672,N_1757);
xor U1843 (N_1843,N_1794,N_1630);
nor U1844 (N_1844,N_1667,N_1686);
nor U1845 (N_1845,N_1779,N_1603);
nand U1846 (N_1846,N_1626,N_1663);
nor U1847 (N_1847,N_1703,N_1741);
nor U1848 (N_1848,N_1694,N_1784);
or U1849 (N_1849,N_1634,N_1791);
nor U1850 (N_1850,N_1752,N_1758);
xor U1851 (N_1851,N_1714,N_1677);
nor U1852 (N_1852,N_1635,N_1600);
nand U1853 (N_1853,N_1780,N_1653);
and U1854 (N_1854,N_1786,N_1762);
and U1855 (N_1855,N_1668,N_1695);
or U1856 (N_1856,N_1763,N_1665);
nand U1857 (N_1857,N_1798,N_1795);
and U1858 (N_1858,N_1764,N_1638);
and U1859 (N_1859,N_1745,N_1664);
or U1860 (N_1860,N_1730,N_1726);
nor U1861 (N_1861,N_1661,N_1679);
and U1862 (N_1862,N_1755,N_1749);
xnor U1863 (N_1863,N_1628,N_1770);
nand U1864 (N_1864,N_1648,N_1691);
nor U1865 (N_1865,N_1619,N_1604);
and U1866 (N_1866,N_1710,N_1627);
or U1867 (N_1867,N_1781,N_1693);
and U1868 (N_1868,N_1676,N_1688);
and U1869 (N_1869,N_1602,N_1633);
or U1870 (N_1870,N_1732,N_1731);
nor U1871 (N_1871,N_1671,N_1698);
nand U1872 (N_1872,N_1680,N_1785);
or U1873 (N_1873,N_1790,N_1799);
nor U1874 (N_1874,N_1728,N_1692);
nand U1875 (N_1875,N_1707,N_1761);
nor U1876 (N_1876,N_1615,N_1655);
xnor U1877 (N_1877,N_1709,N_1778);
xor U1878 (N_1878,N_1610,N_1690);
nor U1879 (N_1879,N_1673,N_1760);
or U1880 (N_1880,N_1623,N_1646);
nand U1881 (N_1881,N_1621,N_1793);
or U1882 (N_1882,N_1797,N_1697);
and U1883 (N_1883,N_1788,N_1662);
nor U1884 (N_1884,N_1645,N_1701);
nand U1885 (N_1885,N_1674,N_1727);
and U1886 (N_1886,N_1632,N_1787);
or U1887 (N_1887,N_1722,N_1713);
or U1888 (N_1888,N_1642,N_1678);
and U1889 (N_1889,N_1618,N_1629);
nor U1890 (N_1890,N_1682,N_1751);
and U1891 (N_1891,N_1702,N_1736);
and U1892 (N_1892,N_1611,N_1767);
or U1893 (N_1893,N_1783,N_1742);
nor U1894 (N_1894,N_1644,N_1753);
nand U1895 (N_1895,N_1771,N_1717);
xor U1896 (N_1896,N_1712,N_1738);
nand U1897 (N_1897,N_1750,N_1636);
xor U1898 (N_1898,N_1681,N_1614);
and U1899 (N_1899,N_1734,N_1756);
nor U1900 (N_1900,N_1682,N_1686);
or U1901 (N_1901,N_1783,N_1748);
or U1902 (N_1902,N_1668,N_1759);
and U1903 (N_1903,N_1777,N_1745);
or U1904 (N_1904,N_1753,N_1702);
or U1905 (N_1905,N_1690,N_1614);
nand U1906 (N_1906,N_1614,N_1687);
nand U1907 (N_1907,N_1765,N_1631);
nor U1908 (N_1908,N_1711,N_1785);
or U1909 (N_1909,N_1769,N_1755);
nor U1910 (N_1910,N_1600,N_1722);
nor U1911 (N_1911,N_1779,N_1712);
or U1912 (N_1912,N_1722,N_1752);
or U1913 (N_1913,N_1746,N_1722);
nor U1914 (N_1914,N_1697,N_1620);
or U1915 (N_1915,N_1656,N_1609);
and U1916 (N_1916,N_1690,N_1667);
and U1917 (N_1917,N_1740,N_1607);
nor U1918 (N_1918,N_1698,N_1768);
nand U1919 (N_1919,N_1678,N_1633);
nand U1920 (N_1920,N_1643,N_1647);
nand U1921 (N_1921,N_1602,N_1798);
and U1922 (N_1922,N_1728,N_1769);
nand U1923 (N_1923,N_1682,N_1798);
nand U1924 (N_1924,N_1617,N_1677);
and U1925 (N_1925,N_1671,N_1798);
nand U1926 (N_1926,N_1647,N_1660);
nand U1927 (N_1927,N_1603,N_1777);
or U1928 (N_1928,N_1779,N_1748);
and U1929 (N_1929,N_1796,N_1798);
or U1930 (N_1930,N_1697,N_1674);
or U1931 (N_1931,N_1621,N_1610);
or U1932 (N_1932,N_1795,N_1678);
nor U1933 (N_1933,N_1736,N_1651);
and U1934 (N_1934,N_1635,N_1709);
or U1935 (N_1935,N_1779,N_1796);
nor U1936 (N_1936,N_1629,N_1756);
nand U1937 (N_1937,N_1642,N_1644);
and U1938 (N_1938,N_1694,N_1642);
nand U1939 (N_1939,N_1751,N_1797);
or U1940 (N_1940,N_1716,N_1745);
nand U1941 (N_1941,N_1646,N_1693);
xor U1942 (N_1942,N_1626,N_1631);
or U1943 (N_1943,N_1785,N_1733);
nand U1944 (N_1944,N_1733,N_1710);
and U1945 (N_1945,N_1649,N_1653);
nand U1946 (N_1946,N_1764,N_1776);
nor U1947 (N_1947,N_1722,N_1788);
nor U1948 (N_1948,N_1719,N_1761);
nand U1949 (N_1949,N_1680,N_1782);
and U1950 (N_1950,N_1732,N_1605);
nor U1951 (N_1951,N_1782,N_1633);
nand U1952 (N_1952,N_1649,N_1794);
and U1953 (N_1953,N_1787,N_1700);
and U1954 (N_1954,N_1788,N_1646);
or U1955 (N_1955,N_1777,N_1700);
xor U1956 (N_1956,N_1787,N_1786);
nand U1957 (N_1957,N_1701,N_1743);
and U1958 (N_1958,N_1633,N_1769);
nand U1959 (N_1959,N_1684,N_1792);
nand U1960 (N_1960,N_1617,N_1711);
nor U1961 (N_1961,N_1614,N_1621);
or U1962 (N_1962,N_1662,N_1705);
and U1963 (N_1963,N_1795,N_1661);
nor U1964 (N_1964,N_1787,N_1617);
or U1965 (N_1965,N_1658,N_1739);
or U1966 (N_1966,N_1706,N_1608);
xnor U1967 (N_1967,N_1724,N_1712);
or U1968 (N_1968,N_1745,N_1791);
nand U1969 (N_1969,N_1627,N_1755);
nor U1970 (N_1970,N_1686,N_1735);
nor U1971 (N_1971,N_1664,N_1799);
or U1972 (N_1972,N_1679,N_1762);
and U1973 (N_1973,N_1618,N_1685);
nand U1974 (N_1974,N_1738,N_1682);
nor U1975 (N_1975,N_1652,N_1701);
nor U1976 (N_1976,N_1795,N_1792);
or U1977 (N_1977,N_1606,N_1704);
and U1978 (N_1978,N_1773,N_1767);
and U1979 (N_1979,N_1777,N_1705);
or U1980 (N_1980,N_1720,N_1687);
nor U1981 (N_1981,N_1733,N_1654);
or U1982 (N_1982,N_1629,N_1692);
or U1983 (N_1983,N_1743,N_1754);
xor U1984 (N_1984,N_1700,N_1712);
nor U1985 (N_1985,N_1765,N_1782);
or U1986 (N_1986,N_1753,N_1617);
xnor U1987 (N_1987,N_1639,N_1600);
and U1988 (N_1988,N_1648,N_1781);
xnor U1989 (N_1989,N_1790,N_1641);
nand U1990 (N_1990,N_1799,N_1693);
nor U1991 (N_1991,N_1611,N_1736);
or U1992 (N_1992,N_1783,N_1736);
nand U1993 (N_1993,N_1761,N_1694);
nand U1994 (N_1994,N_1779,N_1655);
or U1995 (N_1995,N_1655,N_1719);
and U1996 (N_1996,N_1709,N_1609);
nand U1997 (N_1997,N_1671,N_1696);
xnor U1998 (N_1998,N_1663,N_1729);
xnor U1999 (N_1999,N_1748,N_1732);
nor U2000 (N_2000,N_1905,N_1814);
and U2001 (N_2001,N_1994,N_1952);
or U2002 (N_2002,N_1978,N_1899);
nor U2003 (N_2003,N_1927,N_1837);
xnor U2004 (N_2004,N_1818,N_1971);
or U2005 (N_2005,N_1801,N_1925);
xnor U2006 (N_2006,N_1888,N_1937);
and U2007 (N_2007,N_1909,N_1900);
nor U2008 (N_2008,N_1895,N_1924);
nor U2009 (N_2009,N_1896,N_1991);
or U2010 (N_2010,N_1945,N_1889);
nand U2011 (N_2011,N_1988,N_1806);
nor U2012 (N_2012,N_1975,N_1853);
xor U2013 (N_2013,N_1823,N_1831);
nand U2014 (N_2014,N_1923,N_1965);
and U2015 (N_2015,N_1892,N_1826);
xnor U2016 (N_2016,N_1860,N_1986);
nor U2017 (N_2017,N_1939,N_1890);
nor U2018 (N_2018,N_1829,N_1990);
nor U2019 (N_2019,N_1879,N_1805);
xnor U2020 (N_2020,N_1867,N_1874);
nand U2021 (N_2021,N_1836,N_1861);
xnor U2022 (N_2022,N_1834,N_1989);
or U2023 (N_2023,N_1838,N_1910);
or U2024 (N_2024,N_1967,N_1920);
xnor U2025 (N_2025,N_1998,N_1815);
and U2026 (N_2026,N_1865,N_1893);
nor U2027 (N_2027,N_1811,N_1949);
xor U2028 (N_2028,N_1907,N_1983);
and U2029 (N_2029,N_1908,N_1946);
xnor U2030 (N_2030,N_1847,N_1809);
nand U2031 (N_2031,N_1891,N_1824);
nand U2032 (N_2032,N_1850,N_1821);
and U2033 (N_2033,N_1864,N_1901);
nand U2034 (N_2034,N_1881,N_1858);
xor U2035 (N_2035,N_1997,N_1995);
and U2036 (N_2036,N_1869,N_1944);
xnor U2037 (N_2037,N_1820,N_1996);
or U2038 (N_2038,N_1825,N_1974);
and U2039 (N_2039,N_1929,N_1857);
or U2040 (N_2040,N_1954,N_1849);
nand U2041 (N_2041,N_1916,N_1856);
or U2042 (N_2042,N_1948,N_1958);
nor U2043 (N_2043,N_1898,N_1915);
nor U2044 (N_2044,N_1933,N_1928);
nor U2045 (N_2045,N_1813,N_1982);
xor U2046 (N_2046,N_1886,N_1979);
or U2047 (N_2047,N_1819,N_1804);
or U2048 (N_2048,N_1943,N_1951);
nor U2049 (N_2049,N_1887,N_1941);
nand U2050 (N_2050,N_1832,N_1984);
or U2051 (N_2051,N_1873,N_1992);
nor U2052 (N_2052,N_1852,N_1816);
nand U2053 (N_2053,N_1977,N_1976);
nor U2054 (N_2054,N_1914,N_1935);
xnor U2055 (N_2055,N_1833,N_1968);
nand U2056 (N_2056,N_1848,N_1859);
and U2057 (N_2057,N_1930,N_1962);
or U2058 (N_2058,N_1999,N_1885);
nand U2059 (N_2059,N_1808,N_1956);
xor U2060 (N_2060,N_1980,N_1972);
and U2061 (N_2061,N_1830,N_1803);
or U2062 (N_2062,N_1877,N_1917);
or U2063 (N_2063,N_1871,N_1827);
xnor U2064 (N_2064,N_1966,N_1851);
xnor U2065 (N_2065,N_1953,N_1985);
nor U2066 (N_2066,N_1955,N_1846);
nand U2067 (N_2067,N_1940,N_1903);
nand U2068 (N_2068,N_1921,N_1942);
nand U2069 (N_2069,N_1936,N_1922);
or U2070 (N_2070,N_1842,N_1835);
and U2071 (N_2071,N_1841,N_1960);
and U2072 (N_2072,N_1911,N_1840);
xor U2073 (N_2073,N_1904,N_1918);
xor U2074 (N_2074,N_1931,N_1828);
nand U2075 (N_2075,N_1963,N_1810);
or U2076 (N_2076,N_1938,N_1969);
and U2077 (N_2077,N_1872,N_1913);
nand U2078 (N_2078,N_1854,N_1973);
and U2079 (N_2079,N_1894,N_1875);
nor U2080 (N_2080,N_1926,N_1855);
and U2081 (N_2081,N_1883,N_1987);
nor U2082 (N_2082,N_1959,N_1868);
and U2083 (N_2083,N_1897,N_1934);
xnor U2084 (N_2084,N_1802,N_1932);
xnor U2085 (N_2085,N_1844,N_1961);
nor U2086 (N_2086,N_1884,N_1957);
xor U2087 (N_2087,N_1843,N_1970);
xor U2088 (N_2088,N_1947,N_1870);
nor U2089 (N_2089,N_1993,N_1812);
nor U2090 (N_2090,N_1839,N_1919);
xor U2091 (N_2091,N_1981,N_1878);
or U2092 (N_2092,N_1822,N_1880);
nand U2093 (N_2093,N_1866,N_1906);
nor U2094 (N_2094,N_1807,N_1800);
nand U2095 (N_2095,N_1862,N_1964);
nand U2096 (N_2096,N_1912,N_1817);
xor U2097 (N_2097,N_1882,N_1902);
or U2098 (N_2098,N_1950,N_1876);
and U2099 (N_2099,N_1845,N_1863);
and U2100 (N_2100,N_1952,N_1984);
nand U2101 (N_2101,N_1994,N_1929);
nand U2102 (N_2102,N_1847,N_1887);
nor U2103 (N_2103,N_1840,N_1993);
xor U2104 (N_2104,N_1874,N_1831);
nor U2105 (N_2105,N_1984,N_1801);
and U2106 (N_2106,N_1856,N_1897);
nor U2107 (N_2107,N_1924,N_1966);
nor U2108 (N_2108,N_1833,N_1898);
xor U2109 (N_2109,N_1915,N_1986);
nand U2110 (N_2110,N_1859,N_1829);
nand U2111 (N_2111,N_1973,N_1920);
or U2112 (N_2112,N_1870,N_1929);
nor U2113 (N_2113,N_1832,N_1962);
xor U2114 (N_2114,N_1893,N_1927);
xor U2115 (N_2115,N_1931,N_1822);
and U2116 (N_2116,N_1898,N_1933);
or U2117 (N_2117,N_1910,N_1878);
and U2118 (N_2118,N_1813,N_1867);
xnor U2119 (N_2119,N_1802,N_1936);
nor U2120 (N_2120,N_1867,N_1845);
xor U2121 (N_2121,N_1973,N_1864);
nand U2122 (N_2122,N_1923,N_1953);
and U2123 (N_2123,N_1894,N_1977);
nand U2124 (N_2124,N_1806,N_1982);
nand U2125 (N_2125,N_1995,N_1884);
or U2126 (N_2126,N_1821,N_1802);
xnor U2127 (N_2127,N_1915,N_1813);
or U2128 (N_2128,N_1833,N_1959);
or U2129 (N_2129,N_1917,N_1881);
and U2130 (N_2130,N_1811,N_1957);
nor U2131 (N_2131,N_1998,N_1964);
and U2132 (N_2132,N_1955,N_1968);
nand U2133 (N_2133,N_1962,N_1831);
nor U2134 (N_2134,N_1963,N_1936);
or U2135 (N_2135,N_1840,N_1989);
xor U2136 (N_2136,N_1844,N_1926);
or U2137 (N_2137,N_1817,N_1914);
xnor U2138 (N_2138,N_1974,N_1949);
or U2139 (N_2139,N_1856,N_1888);
nor U2140 (N_2140,N_1930,N_1947);
and U2141 (N_2141,N_1987,N_1912);
or U2142 (N_2142,N_1990,N_1903);
and U2143 (N_2143,N_1888,N_1827);
and U2144 (N_2144,N_1980,N_1990);
nand U2145 (N_2145,N_1827,N_1945);
nand U2146 (N_2146,N_1846,N_1810);
nor U2147 (N_2147,N_1917,N_1855);
or U2148 (N_2148,N_1910,N_1913);
nand U2149 (N_2149,N_1993,N_1921);
nor U2150 (N_2150,N_1910,N_1872);
nand U2151 (N_2151,N_1924,N_1834);
or U2152 (N_2152,N_1828,N_1988);
nor U2153 (N_2153,N_1828,N_1999);
nand U2154 (N_2154,N_1871,N_1817);
or U2155 (N_2155,N_1996,N_1929);
or U2156 (N_2156,N_1981,N_1991);
nor U2157 (N_2157,N_1976,N_1862);
xor U2158 (N_2158,N_1871,N_1965);
nand U2159 (N_2159,N_1945,N_1964);
nor U2160 (N_2160,N_1994,N_1845);
nor U2161 (N_2161,N_1940,N_1849);
nand U2162 (N_2162,N_1971,N_1896);
and U2163 (N_2163,N_1930,N_1845);
nand U2164 (N_2164,N_1979,N_1924);
nor U2165 (N_2165,N_1960,N_1961);
nor U2166 (N_2166,N_1925,N_1962);
xor U2167 (N_2167,N_1914,N_1837);
nand U2168 (N_2168,N_1869,N_1934);
nand U2169 (N_2169,N_1878,N_1822);
or U2170 (N_2170,N_1832,N_1849);
xnor U2171 (N_2171,N_1963,N_1856);
or U2172 (N_2172,N_1959,N_1846);
and U2173 (N_2173,N_1980,N_1800);
xor U2174 (N_2174,N_1970,N_1823);
nor U2175 (N_2175,N_1888,N_1835);
or U2176 (N_2176,N_1969,N_1894);
nand U2177 (N_2177,N_1950,N_1879);
and U2178 (N_2178,N_1943,N_1822);
xor U2179 (N_2179,N_1839,N_1970);
nor U2180 (N_2180,N_1864,N_1980);
or U2181 (N_2181,N_1965,N_1960);
or U2182 (N_2182,N_1929,N_1935);
or U2183 (N_2183,N_1830,N_1998);
xor U2184 (N_2184,N_1850,N_1907);
nand U2185 (N_2185,N_1808,N_1940);
nor U2186 (N_2186,N_1831,N_1869);
or U2187 (N_2187,N_1985,N_1942);
nor U2188 (N_2188,N_1972,N_1882);
and U2189 (N_2189,N_1949,N_1962);
and U2190 (N_2190,N_1888,N_1806);
nand U2191 (N_2191,N_1918,N_1947);
nand U2192 (N_2192,N_1936,N_1875);
xor U2193 (N_2193,N_1856,N_1823);
nand U2194 (N_2194,N_1933,N_1945);
nand U2195 (N_2195,N_1805,N_1849);
xnor U2196 (N_2196,N_1823,N_1920);
xnor U2197 (N_2197,N_1917,N_1934);
nand U2198 (N_2198,N_1877,N_1827);
and U2199 (N_2199,N_1808,N_1876);
and U2200 (N_2200,N_2167,N_2110);
nor U2201 (N_2201,N_2081,N_2149);
and U2202 (N_2202,N_2057,N_2100);
xnor U2203 (N_2203,N_2131,N_2150);
and U2204 (N_2204,N_2111,N_2055);
nand U2205 (N_2205,N_2127,N_2122);
and U2206 (N_2206,N_2034,N_2152);
nand U2207 (N_2207,N_2168,N_2171);
or U2208 (N_2208,N_2113,N_2075);
nor U2209 (N_2209,N_2030,N_2071);
and U2210 (N_2210,N_2078,N_2040);
nor U2211 (N_2211,N_2069,N_2107);
xor U2212 (N_2212,N_2160,N_2199);
nor U2213 (N_2213,N_2129,N_2039);
nand U2214 (N_2214,N_2197,N_2137);
xor U2215 (N_2215,N_2102,N_2095);
and U2216 (N_2216,N_2195,N_2181);
or U2217 (N_2217,N_2001,N_2067);
xnor U2218 (N_2218,N_2130,N_2196);
and U2219 (N_2219,N_2024,N_2105);
and U2220 (N_2220,N_2025,N_2052);
nor U2221 (N_2221,N_2178,N_2112);
or U2222 (N_2222,N_2064,N_2161);
nor U2223 (N_2223,N_2033,N_2177);
nor U2224 (N_2224,N_2104,N_2188);
and U2225 (N_2225,N_2094,N_2097);
nor U2226 (N_2226,N_2162,N_2174);
nor U2227 (N_2227,N_2074,N_2054);
and U2228 (N_2228,N_2012,N_2151);
or U2229 (N_2229,N_2096,N_2009);
nor U2230 (N_2230,N_2089,N_2079);
nand U2231 (N_2231,N_2027,N_2043);
xor U2232 (N_2232,N_2017,N_2041);
nand U2233 (N_2233,N_2124,N_2092);
xor U2234 (N_2234,N_2141,N_2116);
and U2235 (N_2235,N_2190,N_2179);
or U2236 (N_2236,N_2106,N_2060);
nor U2237 (N_2237,N_2066,N_2077);
nor U2238 (N_2238,N_2144,N_2063);
nor U2239 (N_2239,N_2090,N_2032);
or U2240 (N_2240,N_2046,N_2065);
xor U2241 (N_2241,N_2068,N_2047);
nor U2242 (N_2242,N_2015,N_2053);
or U2243 (N_2243,N_2083,N_2058);
or U2244 (N_2244,N_2008,N_2029);
nor U2245 (N_2245,N_2087,N_2010);
nor U2246 (N_2246,N_2136,N_2082);
or U2247 (N_2247,N_2133,N_2147);
or U2248 (N_2248,N_2016,N_2134);
xnor U2249 (N_2249,N_2125,N_2042);
or U2250 (N_2250,N_2050,N_2021);
nor U2251 (N_2251,N_2123,N_2182);
nand U2252 (N_2252,N_2093,N_2038);
nand U2253 (N_2253,N_2132,N_2080);
nor U2254 (N_2254,N_2004,N_2186);
or U2255 (N_2255,N_2026,N_2164);
nor U2256 (N_2256,N_2166,N_2155);
nand U2257 (N_2257,N_2076,N_2194);
nor U2258 (N_2258,N_2165,N_2121);
nor U2259 (N_2259,N_2035,N_2098);
xnor U2260 (N_2260,N_2014,N_2062);
or U2261 (N_2261,N_2051,N_2189);
nor U2262 (N_2262,N_2118,N_2006);
nor U2263 (N_2263,N_2101,N_2139);
or U2264 (N_2264,N_2193,N_2045);
or U2265 (N_2265,N_2114,N_2091);
nor U2266 (N_2266,N_2085,N_2005);
and U2267 (N_2267,N_2138,N_2018);
nor U2268 (N_2268,N_2146,N_2037);
nand U2269 (N_2269,N_2140,N_2048);
xor U2270 (N_2270,N_2011,N_2070);
nor U2271 (N_2271,N_2023,N_2099);
or U2272 (N_2272,N_2135,N_2145);
nand U2273 (N_2273,N_2013,N_2183);
xor U2274 (N_2274,N_2153,N_2180);
and U2275 (N_2275,N_2031,N_2154);
and U2276 (N_2276,N_2156,N_2044);
nand U2277 (N_2277,N_2003,N_2109);
nor U2278 (N_2278,N_2128,N_2192);
xor U2279 (N_2279,N_2163,N_2120);
xor U2280 (N_2280,N_2028,N_2172);
and U2281 (N_2281,N_2198,N_2036);
nand U2282 (N_2282,N_2115,N_2173);
and U2283 (N_2283,N_2148,N_2000);
and U2284 (N_2284,N_2191,N_2002);
or U2285 (N_2285,N_2061,N_2059);
and U2286 (N_2286,N_2084,N_2108);
xnor U2287 (N_2287,N_2157,N_2126);
xnor U2288 (N_2288,N_2103,N_2073);
nor U2289 (N_2289,N_2020,N_2072);
and U2290 (N_2290,N_2056,N_2184);
nor U2291 (N_2291,N_2176,N_2169);
or U2292 (N_2292,N_2019,N_2022);
nor U2293 (N_2293,N_2117,N_2086);
nor U2294 (N_2294,N_2159,N_2175);
and U2295 (N_2295,N_2187,N_2143);
xnor U2296 (N_2296,N_2158,N_2088);
xor U2297 (N_2297,N_2119,N_2049);
and U2298 (N_2298,N_2185,N_2142);
nor U2299 (N_2299,N_2170,N_2007);
and U2300 (N_2300,N_2186,N_2176);
nand U2301 (N_2301,N_2140,N_2025);
nor U2302 (N_2302,N_2136,N_2077);
xnor U2303 (N_2303,N_2104,N_2069);
xnor U2304 (N_2304,N_2045,N_2081);
and U2305 (N_2305,N_2146,N_2160);
nor U2306 (N_2306,N_2018,N_2023);
and U2307 (N_2307,N_2126,N_2196);
xor U2308 (N_2308,N_2154,N_2049);
and U2309 (N_2309,N_2173,N_2024);
nor U2310 (N_2310,N_2001,N_2091);
xnor U2311 (N_2311,N_2028,N_2004);
nand U2312 (N_2312,N_2032,N_2075);
nand U2313 (N_2313,N_2040,N_2177);
nor U2314 (N_2314,N_2047,N_2032);
nor U2315 (N_2315,N_2124,N_2100);
nand U2316 (N_2316,N_2170,N_2164);
nor U2317 (N_2317,N_2162,N_2141);
nor U2318 (N_2318,N_2065,N_2178);
or U2319 (N_2319,N_2052,N_2007);
and U2320 (N_2320,N_2022,N_2198);
and U2321 (N_2321,N_2162,N_2017);
xor U2322 (N_2322,N_2143,N_2130);
nor U2323 (N_2323,N_2155,N_2169);
nor U2324 (N_2324,N_2107,N_2147);
and U2325 (N_2325,N_2028,N_2182);
and U2326 (N_2326,N_2010,N_2121);
and U2327 (N_2327,N_2092,N_2166);
and U2328 (N_2328,N_2031,N_2004);
xor U2329 (N_2329,N_2118,N_2159);
nor U2330 (N_2330,N_2041,N_2138);
nor U2331 (N_2331,N_2058,N_2009);
or U2332 (N_2332,N_2077,N_2045);
xor U2333 (N_2333,N_2092,N_2040);
or U2334 (N_2334,N_2154,N_2061);
xnor U2335 (N_2335,N_2032,N_2150);
xor U2336 (N_2336,N_2051,N_2033);
xor U2337 (N_2337,N_2006,N_2125);
or U2338 (N_2338,N_2107,N_2016);
nand U2339 (N_2339,N_2023,N_2054);
xor U2340 (N_2340,N_2058,N_2103);
or U2341 (N_2341,N_2195,N_2134);
nand U2342 (N_2342,N_2063,N_2179);
nand U2343 (N_2343,N_2120,N_2133);
nand U2344 (N_2344,N_2122,N_2070);
or U2345 (N_2345,N_2056,N_2071);
nand U2346 (N_2346,N_2037,N_2199);
nand U2347 (N_2347,N_2117,N_2186);
nand U2348 (N_2348,N_2177,N_2064);
xnor U2349 (N_2349,N_2039,N_2030);
or U2350 (N_2350,N_2081,N_2161);
xor U2351 (N_2351,N_2042,N_2198);
xor U2352 (N_2352,N_2100,N_2115);
nand U2353 (N_2353,N_2034,N_2014);
nor U2354 (N_2354,N_2143,N_2091);
or U2355 (N_2355,N_2163,N_2027);
and U2356 (N_2356,N_2031,N_2111);
xnor U2357 (N_2357,N_2028,N_2083);
or U2358 (N_2358,N_2138,N_2043);
nand U2359 (N_2359,N_2139,N_2037);
nor U2360 (N_2360,N_2154,N_2122);
nor U2361 (N_2361,N_2134,N_2053);
nor U2362 (N_2362,N_2134,N_2179);
or U2363 (N_2363,N_2034,N_2068);
and U2364 (N_2364,N_2138,N_2147);
xnor U2365 (N_2365,N_2088,N_2043);
nand U2366 (N_2366,N_2125,N_2187);
xor U2367 (N_2367,N_2178,N_2199);
or U2368 (N_2368,N_2044,N_2005);
nor U2369 (N_2369,N_2008,N_2086);
or U2370 (N_2370,N_2128,N_2050);
nor U2371 (N_2371,N_2185,N_2165);
or U2372 (N_2372,N_2141,N_2068);
xnor U2373 (N_2373,N_2039,N_2195);
and U2374 (N_2374,N_2046,N_2168);
or U2375 (N_2375,N_2117,N_2172);
or U2376 (N_2376,N_2037,N_2067);
or U2377 (N_2377,N_2076,N_2162);
and U2378 (N_2378,N_2086,N_2178);
xnor U2379 (N_2379,N_2039,N_2077);
nand U2380 (N_2380,N_2175,N_2071);
nand U2381 (N_2381,N_2001,N_2100);
nand U2382 (N_2382,N_2185,N_2055);
or U2383 (N_2383,N_2158,N_2196);
nand U2384 (N_2384,N_2059,N_2008);
xnor U2385 (N_2385,N_2165,N_2119);
xor U2386 (N_2386,N_2108,N_2065);
nor U2387 (N_2387,N_2119,N_2039);
nor U2388 (N_2388,N_2142,N_2149);
and U2389 (N_2389,N_2007,N_2084);
and U2390 (N_2390,N_2139,N_2111);
xnor U2391 (N_2391,N_2118,N_2174);
xor U2392 (N_2392,N_2015,N_2167);
xnor U2393 (N_2393,N_2093,N_2146);
xnor U2394 (N_2394,N_2122,N_2074);
or U2395 (N_2395,N_2166,N_2160);
nand U2396 (N_2396,N_2042,N_2112);
xnor U2397 (N_2397,N_2137,N_2011);
or U2398 (N_2398,N_2032,N_2194);
xor U2399 (N_2399,N_2021,N_2170);
and U2400 (N_2400,N_2277,N_2284);
or U2401 (N_2401,N_2287,N_2214);
nor U2402 (N_2402,N_2220,N_2372);
nor U2403 (N_2403,N_2245,N_2371);
and U2404 (N_2404,N_2259,N_2393);
xnor U2405 (N_2405,N_2240,N_2255);
nor U2406 (N_2406,N_2385,N_2300);
nand U2407 (N_2407,N_2293,N_2201);
and U2408 (N_2408,N_2331,N_2225);
or U2409 (N_2409,N_2213,N_2263);
and U2410 (N_2410,N_2378,N_2320);
nand U2411 (N_2411,N_2328,N_2250);
nand U2412 (N_2412,N_2272,N_2370);
or U2413 (N_2413,N_2342,N_2376);
or U2414 (N_2414,N_2206,N_2265);
nand U2415 (N_2415,N_2207,N_2337);
nand U2416 (N_2416,N_2353,N_2347);
nand U2417 (N_2417,N_2308,N_2382);
or U2418 (N_2418,N_2394,N_2398);
xor U2419 (N_2419,N_2235,N_2262);
and U2420 (N_2420,N_2319,N_2325);
xor U2421 (N_2421,N_2222,N_2321);
or U2422 (N_2422,N_2266,N_2291);
and U2423 (N_2423,N_2358,N_2362);
or U2424 (N_2424,N_2384,N_2396);
or U2425 (N_2425,N_2399,N_2256);
xnor U2426 (N_2426,N_2269,N_2279);
xnor U2427 (N_2427,N_2217,N_2379);
nand U2428 (N_2428,N_2258,N_2289);
and U2429 (N_2429,N_2387,N_2373);
xor U2430 (N_2430,N_2200,N_2286);
nor U2431 (N_2431,N_2390,N_2381);
and U2432 (N_2432,N_2233,N_2314);
xor U2433 (N_2433,N_2309,N_2202);
nand U2434 (N_2434,N_2208,N_2231);
and U2435 (N_2435,N_2303,N_2251);
nand U2436 (N_2436,N_2330,N_2299);
nand U2437 (N_2437,N_2365,N_2356);
nor U2438 (N_2438,N_2329,N_2311);
nor U2439 (N_2439,N_2275,N_2268);
nand U2440 (N_2440,N_2361,N_2210);
nand U2441 (N_2441,N_2282,N_2351);
and U2442 (N_2442,N_2271,N_2360);
or U2443 (N_2443,N_2260,N_2334);
nand U2444 (N_2444,N_2344,N_2230);
xor U2445 (N_2445,N_2312,N_2333);
xor U2446 (N_2446,N_2267,N_2313);
and U2447 (N_2447,N_2305,N_2310);
or U2448 (N_2448,N_2315,N_2288);
and U2449 (N_2449,N_2335,N_2332);
or U2450 (N_2450,N_2204,N_2248);
nand U2451 (N_2451,N_2323,N_2211);
and U2452 (N_2452,N_2343,N_2366);
and U2453 (N_2453,N_2237,N_2339);
or U2454 (N_2454,N_2395,N_2397);
xor U2455 (N_2455,N_2292,N_2252);
nand U2456 (N_2456,N_2254,N_2226);
nor U2457 (N_2457,N_2290,N_2285);
nand U2458 (N_2458,N_2242,N_2340);
nand U2459 (N_2459,N_2354,N_2297);
xor U2460 (N_2460,N_2257,N_2380);
nor U2461 (N_2461,N_2280,N_2249);
nand U2462 (N_2462,N_2236,N_2229);
and U2463 (N_2463,N_2244,N_2246);
xnor U2464 (N_2464,N_2368,N_2324);
nor U2465 (N_2465,N_2295,N_2261);
and U2466 (N_2466,N_2363,N_2274);
and U2467 (N_2467,N_2228,N_2221);
and U2468 (N_2468,N_2307,N_2349);
xor U2469 (N_2469,N_2346,N_2345);
xnor U2470 (N_2470,N_2238,N_2318);
and U2471 (N_2471,N_2364,N_2209);
xor U2472 (N_2472,N_2316,N_2224);
xnor U2473 (N_2473,N_2278,N_2388);
nor U2474 (N_2474,N_2392,N_2216);
nand U2475 (N_2475,N_2281,N_2391);
nor U2476 (N_2476,N_2317,N_2212);
and U2477 (N_2477,N_2296,N_2386);
xor U2478 (N_2478,N_2270,N_2227);
or U2479 (N_2479,N_2276,N_2348);
nor U2480 (N_2480,N_2383,N_2302);
or U2481 (N_2481,N_2369,N_2306);
nand U2482 (N_2482,N_2389,N_2322);
and U2483 (N_2483,N_2352,N_2273);
and U2484 (N_2484,N_2377,N_2374);
or U2485 (N_2485,N_2338,N_2203);
nor U2486 (N_2486,N_2367,N_2327);
or U2487 (N_2487,N_2304,N_2223);
and U2488 (N_2488,N_2243,N_2234);
xor U2489 (N_2489,N_2232,N_2264);
xnor U2490 (N_2490,N_2283,N_2301);
nor U2491 (N_2491,N_2326,N_2359);
or U2492 (N_2492,N_2375,N_2205);
nand U2493 (N_2493,N_2239,N_2357);
nor U2494 (N_2494,N_2341,N_2219);
nor U2495 (N_2495,N_2247,N_2215);
or U2496 (N_2496,N_2298,N_2218);
nor U2497 (N_2497,N_2355,N_2241);
or U2498 (N_2498,N_2294,N_2253);
or U2499 (N_2499,N_2350,N_2336);
and U2500 (N_2500,N_2384,N_2205);
and U2501 (N_2501,N_2355,N_2318);
or U2502 (N_2502,N_2290,N_2393);
and U2503 (N_2503,N_2374,N_2241);
nor U2504 (N_2504,N_2389,N_2204);
nand U2505 (N_2505,N_2252,N_2256);
nand U2506 (N_2506,N_2236,N_2339);
nor U2507 (N_2507,N_2218,N_2303);
nor U2508 (N_2508,N_2338,N_2206);
nor U2509 (N_2509,N_2237,N_2330);
and U2510 (N_2510,N_2219,N_2220);
nor U2511 (N_2511,N_2207,N_2394);
nand U2512 (N_2512,N_2222,N_2268);
or U2513 (N_2513,N_2334,N_2213);
nand U2514 (N_2514,N_2309,N_2283);
and U2515 (N_2515,N_2288,N_2352);
xor U2516 (N_2516,N_2296,N_2233);
nand U2517 (N_2517,N_2206,N_2349);
nor U2518 (N_2518,N_2242,N_2206);
or U2519 (N_2519,N_2347,N_2283);
xor U2520 (N_2520,N_2277,N_2341);
and U2521 (N_2521,N_2365,N_2204);
or U2522 (N_2522,N_2283,N_2285);
xor U2523 (N_2523,N_2201,N_2238);
nand U2524 (N_2524,N_2301,N_2252);
and U2525 (N_2525,N_2358,N_2268);
nor U2526 (N_2526,N_2362,N_2207);
nand U2527 (N_2527,N_2238,N_2321);
xor U2528 (N_2528,N_2355,N_2275);
xor U2529 (N_2529,N_2265,N_2327);
or U2530 (N_2530,N_2333,N_2268);
and U2531 (N_2531,N_2249,N_2233);
nand U2532 (N_2532,N_2269,N_2368);
or U2533 (N_2533,N_2333,N_2338);
or U2534 (N_2534,N_2240,N_2216);
xor U2535 (N_2535,N_2342,N_2238);
nor U2536 (N_2536,N_2284,N_2213);
or U2537 (N_2537,N_2232,N_2255);
nand U2538 (N_2538,N_2276,N_2352);
nor U2539 (N_2539,N_2282,N_2303);
nand U2540 (N_2540,N_2255,N_2380);
and U2541 (N_2541,N_2361,N_2317);
xor U2542 (N_2542,N_2292,N_2267);
xor U2543 (N_2543,N_2384,N_2299);
nor U2544 (N_2544,N_2313,N_2340);
nand U2545 (N_2545,N_2276,N_2216);
nand U2546 (N_2546,N_2225,N_2398);
nand U2547 (N_2547,N_2217,N_2348);
nor U2548 (N_2548,N_2339,N_2252);
nor U2549 (N_2549,N_2383,N_2346);
xnor U2550 (N_2550,N_2257,N_2223);
or U2551 (N_2551,N_2347,N_2275);
or U2552 (N_2552,N_2256,N_2367);
nand U2553 (N_2553,N_2315,N_2274);
or U2554 (N_2554,N_2354,N_2286);
nor U2555 (N_2555,N_2284,N_2301);
or U2556 (N_2556,N_2218,N_2209);
and U2557 (N_2557,N_2312,N_2380);
xnor U2558 (N_2558,N_2209,N_2397);
or U2559 (N_2559,N_2244,N_2258);
xor U2560 (N_2560,N_2219,N_2354);
xor U2561 (N_2561,N_2308,N_2217);
nand U2562 (N_2562,N_2231,N_2228);
or U2563 (N_2563,N_2206,N_2238);
nand U2564 (N_2564,N_2332,N_2358);
nor U2565 (N_2565,N_2394,N_2329);
xor U2566 (N_2566,N_2320,N_2336);
nor U2567 (N_2567,N_2294,N_2279);
nand U2568 (N_2568,N_2286,N_2213);
nor U2569 (N_2569,N_2300,N_2367);
nor U2570 (N_2570,N_2351,N_2355);
or U2571 (N_2571,N_2210,N_2291);
and U2572 (N_2572,N_2306,N_2351);
nand U2573 (N_2573,N_2384,N_2337);
nand U2574 (N_2574,N_2202,N_2227);
and U2575 (N_2575,N_2258,N_2223);
xnor U2576 (N_2576,N_2214,N_2224);
nand U2577 (N_2577,N_2352,N_2357);
nor U2578 (N_2578,N_2266,N_2322);
xor U2579 (N_2579,N_2296,N_2261);
nor U2580 (N_2580,N_2219,N_2206);
nand U2581 (N_2581,N_2342,N_2335);
nor U2582 (N_2582,N_2303,N_2362);
nand U2583 (N_2583,N_2377,N_2294);
or U2584 (N_2584,N_2214,N_2280);
nand U2585 (N_2585,N_2344,N_2371);
and U2586 (N_2586,N_2238,N_2202);
xor U2587 (N_2587,N_2279,N_2203);
nor U2588 (N_2588,N_2366,N_2320);
or U2589 (N_2589,N_2361,N_2260);
nand U2590 (N_2590,N_2271,N_2367);
nand U2591 (N_2591,N_2288,N_2219);
and U2592 (N_2592,N_2220,N_2283);
xnor U2593 (N_2593,N_2348,N_2306);
xor U2594 (N_2594,N_2382,N_2201);
xnor U2595 (N_2595,N_2260,N_2209);
and U2596 (N_2596,N_2368,N_2263);
or U2597 (N_2597,N_2335,N_2325);
xnor U2598 (N_2598,N_2280,N_2315);
or U2599 (N_2599,N_2240,N_2261);
nor U2600 (N_2600,N_2509,N_2408);
xnor U2601 (N_2601,N_2537,N_2595);
or U2602 (N_2602,N_2433,N_2470);
nand U2603 (N_2603,N_2542,N_2524);
or U2604 (N_2604,N_2425,N_2518);
and U2605 (N_2605,N_2449,N_2448);
nand U2606 (N_2606,N_2547,N_2516);
nor U2607 (N_2607,N_2406,N_2461);
and U2608 (N_2608,N_2441,N_2454);
nor U2609 (N_2609,N_2522,N_2426);
nand U2610 (N_2610,N_2498,N_2440);
nor U2611 (N_2611,N_2418,N_2576);
nor U2612 (N_2612,N_2479,N_2584);
nand U2613 (N_2613,N_2413,N_2581);
and U2614 (N_2614,N_2520,N_2558);
nor U2615 (N_2615,N_2499,N_2519);
and U2616 (N_2616,N_2421,N_2415);
nand U2617 (N_2617,N_2561,N_2510);
xnor U2618 (N_2618,N_2599,N_2540);
nand U2619 (N_2619,N_2432,N_2469);
nand U2620 (N_2620,N_2551,N_2525);
nor U2621 (N_2621,N_2500,N_2563);
nor U2622 (N_2622,N_2577,N_2564);
nor U2623 (N_2623,N_2445,N_2405);
or U2624 (N_2624,N_2492,N_2553);
and U2625 (N_2625,N_2447,N_2471);
xor U2626 (N_2626,N_2452,N_2503);
nand U2627 (N_2627,N_2538,N_2586);
and U2628 (N_2628,N_2434,N_2552);
xnor U2629 (N_2629,N_2526,N_2407);
and U2630 (N_2630,N_2589,N_2568);
and U2631 (N_2631,N_2569,N_2462);
nand U2632 (N_2632,N_2481,N_2442);
and U2633 (N_2633,N_2478,N_2596);
and U2634 (N_2634,N_2513,N_2570);
or U2635 (N_2635,N_2468,N_2456);
xor U2636 (N_2636,N_2429,N_2531);
xnor U2637 (N_2637,N_2411,N_2475);
nand U2638 (N_2638,N_2582,N_2453);
nor U2639 (N_2639,N_2420,N_2501);
and U2640 (N_2640,N_2450,N_2556);
nand U2641 (N_2641,N_2549,N_2508);
and U2642 (N_2642,N_2439,N_2419);
nor U2643 (N_2643,N_2567,N_2505);
nor U2644 (N_2644,N_2463,N_2428);
xor U2645 (N_2645,N_2400,N_2459);
nor U2646 (N_2646,N_2457,N_2517);
nor U2647 (N_2647,N_2528,N_2521);
nor U2648 (N_2648,N_2446,N_2482);
xor U2649 (N_2649,N_2476,N_2473);
nand U2650 (N_2650,N_2597,N_2490);
and U2651 (N_2651,N_2583,N_2571);
or U2652 (N_2652,N_2485,N_2417);
nor U2653 (N_2653,N_2491,N_2423);
and U2654 (N_2654,N_2580,N_2474);
xor U2655 (N_2655,N_2507,N_2545);
xor U2656 (N_2656,N_2557,N_2430);
nand U2657 (N_2657,N_2451,N_2532);
or U2658 (N_2658,N_2541,N_2493);
and U2659 (N_2659,N_2458,N_2533);
nand U2660 (N_2660,N_2497,N_2578);
xnor U2661 (N_2661,N_2495,N_2486);
and U2662 (N_2662,N_2554,N_2594);
nor U2663 (N_2663,N_2550,N_2435);
xor U2664 (N_2664,N_2467,N_2483);
xor U2665 (N_2665,N_2422,N_2555);
or U2666 (N_2666,N_2424,N_2504);
xnor U2667 (N_2667,N_2527,N_2466);
xor U2668 (N_2668,N_2588,N_2511);
nor U2669 (N_2669,N_2562,N_2573);
and U2670 (N_2670,N_2514,N_2480);
or U2671 (N_2671,N_2494,N_2592);
xnor U2672 (N_2672,N_2414,N_2598);
nor U2673 (N_2673,N_2401,N_2437);
or U2674 (N_2674,N_2487,N_2529);
nand U2675 (N_2675,N_2410,N_2412);
nand U2676 (N_2676,N_2534,N_2515);
and U2677 (N_2677,N_2523,N_2587);
and U2678 (N_2678,N_2465,N_2489);
xnor U2679 (N_2679,N_2512,N_2460);
and U2680 (N_2680,N_2548,N_2464);
xnor U2681 (N_2681,N_2593,N_2402);
nor U2682 (N_2682,N_2560,N_2575);
and U2683 (N_2683,N_2472,N_2496);
xor U2684 (N_2684,N_2591,N_2543);
xor U2685 (N_2685,N_2403,N_2502);
xor U2686 (N_2686,N_2565,N_2409);
nand U2687 (N_2687,N_2544,N_2436);
nand U2688 (N_2688,N_2416,N_2579);
nor U2689 (N_2689,N_2590,N_2566);
nor U2690 (N_2690,N_2404,N_2535);
and U2691 (N_2691,N_2431,N_2506);
xnor U2692 (N_2692,N_2530,N_2539);
xor U2693 (N_2693,N_2455,N_2536);
and U2694 (N_2694,N_2559,N_2438);
or U2695 (N_2695,N_2585,N_2488);
or U2696 (N_2696,N_2572,N_2484);
nor U2697 (N_2697,N_2574,N_2427);
and U2698 (N_2698,N_2546,N_2477);
nand U2699 (N_2699,N_2444,N_2443);
xnor U2700 (N_2700,N_2594,N_2551);
and U2701 (N_2701,N_2589,N_2583);
and U2702 (N_2702,N_2472,N_2527);
nor U2703 (N_2703,N_2570,N_2530);
nor U2704 (N_2704,N_2531,N_2573);
xnor U2705 (N_2705,N_2496,N_2568);
nand U2706 (N_2706,N_2520,N_2567);
nand U2707 (N_2707,N_2534,N_2568);
nand U2708 (N_2708,N_2428,N_2557);
nand U2709 (N_2709,N_2591,N_2555);
nand U2710 (N_2710,N_2456,N_2417);
nor U2711 (N_2711,N_2539,N_2535);
nand U2712 (N_2712,N_2471,N_2412);
or U2713 (N_2713,N_2563,N_2525);
nor U2714 (N_2714,N_2580,N_2553);
xnor U2715 (N_2715,N_2567,N_2420);
and U2716 (N_2716,N_2407,N_2442);
xnor U2717 (N_2717,N_2469,N_2419);
xnor U2718 (N_2718,N_2467,N_2587);
and U2719 (N_2719,N_2444,N_2543);
xor U2720 (N_2720,N_2423,N_2449);
nand U2721 (N_2721,N_2517,N_2450);
xor U2722 (N_2722,N_2405,N_2458);
nor U2723 (N_2723,N_2469,N_2463);
and U2724 (N_2724,N_2483,N_2578);
nor U2725 (N_2725,N_2519,N_2526);
nor U2726 (N_2726,N_2432,N_2471);
or U2727 (N_2727,N_2456,N_2489);
xor U2728 (N_2728,N_2558,N_2570);
or U2729 (N_2729,N_2478,N_2576);
and U2730 (N_2730,N_2419,N_2536);
or U2731 (N_2731,N_2439,N_2441);
and U2732 (N_2732,N_2437,N_2470);
nor U2733 (N_2733,N_2557,N_2435);
and U2734 (N_2734,N_2462,N_2506);
xnor U2735 (N_2735,N_2488,N_2544);
xnor U2736 (N_2736,N_2538,N_2437);
or U2737 (N_2737,N_2555,N_2477);
xor U2738 (N_2738,N_2459,N_2426);
or U2739 (N_2739,N_2576,N_2487);
and U2740 (N_2740,N_2529,N_2463);
and U2741 (N_2741,N_2493,N_2571);
nand U2742 (N_2742,N_2542,N_2443);
nor U2743 (N_2743,N_2527,N_2533);
or U2744 (N_2744,N_2519,N_2560);
nand U2745 (N_2745,N_2448,N_2546);
xnor U2746 (N_2746,N_2512,N_2502);
nor U2747 (N_2747,N_2501,N_2459);
or U2748 (N_2748,N_2447,N_2481);
xnor U2749 (N_2749,N_2424,N_2517);
and U2750 (N_2750,N_2474,N_2514);
xnor U2751 (N_2751,N_2477,N_2418);
nand U2752 (N_2752,N_2406,N_2403);
or U2753 (N_2753,N_2542,N_2579);
nand U2754 (N_2754,N_2578,N_2506);
or U2755 (N_2755,N_2561,N_2567);
xnor U2756 (N_2756,N_2413,N_2402);
nor U2757 (N_2757,N_2576,N_2503);
nand U2758 (N_2758,N_2522,N_2444);
nor U2759 (N_2759,N_2484,N_2496);
or U2760 (N_2760,N_2447,N_2539);
or U2761 (N_2761,N_2543,N_2420);
xor U2762 (N_2762,N_2489,N_2434);
xnor U2763 (N_2763,N_2538,N_2404);
xnor U2764 (N_2764,N_2472,N_2432);
and U2765 (N_2765,N_2503,N_2572);
or U2766 (N_2766,N_2452,N_2426);
nand U2767 (N_2767,N_2571,N_2485);
and U2768 (N_2768,N_2478,N_2466);
nand U2769 (N_2769,N_2518,N_2550);
nor U2770 (N_2770,N_2546,N_2460);
or U2771 (N_2771,N_2573,N_2520);
xnor U2772 (N_2772,N_2511,N_2563);
and U2773 (N_2773,N_2467,N_2535);
and U2774 (N_2774,N_2434,N_2535);
and U2775 (N_2775,N_2565,N_2477);
nor U2776 (N_2776,N_2425,N_2468);
or U2777 (N_2777,N_2516,N_2403);
or U2778 (N_2778,N_2492,N_2551);
or U2779 (N_2779,N_2493,N_2579);
xor U2780 (N_2780,N_2519,N_2426);
xor U2781 (N_2781,N_2598,N_2403);
or U2782 (N_2782,N_2458,N_2450);
nand U2783 (N_2783,N_2461,N_2589);
nor U2784 (N_2784,N_2518,N_2484);
or U2785 (N_2785,N_2492,N_2504);
nor U2786 (N_2786,N_2462,N_2409);
and U2787 (N_2787,N_2464,N_2533);
and U2788 (N_2788,N_2493,N_2425);
and U2789 (N_2789,N_2415,N_2538);
and U2790 (N_2790,N_2409,N_2552);
or U2791 (N_2791,N_2541,N_2412);
nor U2792 (N_2792,N_2582,N_2467);
xnor U2793 (N_2793,N_2596,N_2545);
nand U2794 (N_2794,N_2546,N_2421);
nor U2795 (N_2795,N_2505,N_2464);
or U2796 (N_2796,N_2596,N_2454);
nand U2797 (N_2797,N_2537,N_2522);
nand U2798 (N_2798,N_2463,N_2425);
or U2799 (N_2799,N_2468,N_2476);
xnor U2800 (N_2800,N_2710,N_2792);
or U2801 (N_2801,N_2654,N_2791);
nor U2802 (N_2802,N_2779,N_2731);
nand U2803 (N_2803,N_2711,N_2608);
nor U2804 (N_2804,N_2647,N_2646);
and U2805 (N_2805,N_2768,N_2741);
nand U2806 (N_2806,N_2715,N_2604);
and U2807 (N_2807,N_2753,N_2697);
nand U2808 (N_2808,N_2784,N_2764);
nand U2809 (N_2809,N_2755,N_2648);
nor U2810 (N_2810,N_2609,N_2698);
and U2811 (N_2811,N_2651,N_2650);
nor U2812 (N_2812,N_2720,N_2781);
nor U2813 (N_2813,N_2636,N_2645);
or U2814 (N_2814,N_2771,N_2670);
nor U2815 (N_2815,N_2610,N_2727);
xnor U2816 (N_2816,N_2740,N_2726);
xor U2817 (N_2817,N_2713,N_2666);
nor U2818 (N_2818,N_2621,N_2649);
xnor U2819 (N_2819,N_2744,N_2663);
or U2820 (N_2820,N_2657,N_2765);
nor U2821 (N_2821,N_2702,N_2742);
and U2822 (N_2822,N_2746,N_2766);
or U2823 (N_2823,N_2605,N_2619);
nor U2824 (N_2824,N_2681,N_2637);
and U2825 (N_2825,N_2616,N_2736);
or U2826 (N_2826,N_2738,N_2695);
and U2827 (N_2827,N_2793,N_2614);
or U2828 (N_2828,N_2712,N_2709);
xnor U2829 (N_2829,N_2603,N_2794);
nor U2830 (N_2830,N_2734,N_2620);
nand U2831 (N_2831,N_2611,N_2725);
xor U2832 (N_2832,N_2658,N_2788);
nor U2833 (N_2833,N_2661,N_2703);
xor U2834 (N_2834,N_2743,N_2628);
and U2835 (N_2835,N_2707,N_2721);
nand U2836 (N_2836,N_2680,N_2659);
xor U2837 (N_2837,N_2686,N_2769);
nor U2838 (N_2838,N_2653,N_2683);
nand U2839 (N_2839,N_2652,N_2691);
or U2840 (N_2840,N_2722,N_2679);
nor U2841 (N_2841,N_2730,N_2799);
and U2842 (N_2842,N_2701,N_2618);
xor U2843 (N_2843,N_2719,N_2797);
xnor U2844 (N_2844,N_2789,N_2600);
nor U2845 (N_2845,N_2762,N_2717);
or U2846 (N_2846,N_2641,N_2625);
and U2847 (N_2847,N_2623,N_2700);
or U2848 (N_2848,N_2633,N_2728);
or U2849 (N_2849,N_2758,N_2639);
nor U2850 (N_2850,N_2796,N_2682);
or U2851 (N_2851,N_2677,N_2732);
or U2852 (N_2852,N_2662,N_2748);
nor U2853 (N_2853,N_2737,N_2782);
nand U2854 (N_2854,N_2723,N_2607);
nor U2855 (N_2855,N_2631,N_2676);
and U2856 (N_2856,N_2774,N_2626);
nor U2857 (N_2857,N_2783,N_2729);
nand U2858 (N_2858,N_2638,N_2747);
xnor U2859 (N_2859,N_2724,N_2750);
and U2860 (N_2860,N_2798,N_2675);
or U2861 (N_2861,N_2643,N_2671);
or U2862 (N_2862,N_2790,N_2690);
and U2863 (N_2863,N_2776,N_2640);
xor U2864 (N_2864,N_2622,N_2669);
nor U2865 (N_2865,N_2673,N_2775);
or U2866 (N_2866,N_2688,N_2795);
nor U2867 (N_2867,N_2696,N_2787);
xor U2868 (N_2868,N_2693,N_2668);
nor U2869 (N_2869,N_2627,N_2694);
and U2870 (N_2870,N_2718,N_2759);
nor U2871 (N_2871,N_2642,N_2763);
or U2872 (N_2872,N_2678,N_2689);
nor U2873 (N_2873,N_2606,N_2687);
nand U2874 (N_2874,N_2692,N_2786);
nand U2875 (N_2875,N_2601,N_2767);
or U2876 (N_2876,N_2770,N_2735);
xnor U2877 (N_2877,N_2716,N_2635);
xor U2878 (N_2878,N_2706,N_2602);
or U2879 (N_2879,N_2632,N_2704);
xor U2880 (N_2880,N_2685,N_2667);
or U2881 (N_2881,N_2778,N_2615);
nor U2882 (N_2882,N_2705,N_2777);
and U2883 (N_2883,N_2664,N_2644);
xnor U2884 (N_2884,N_2772,N_2660);
or U2885 (N_2885,N_2634,N_2612);
and U2886 (N_2886,N_2617,N_2752);
or U2887 (N_2887,N_2757,N_2624);
and U2888 (N_2888,N_2684,N_2785);
xnor U2889 (N_2889,N_2751,N_2754);
xor U2890 (N_2890,N_2745,N_2780);
or U2891 (N_2891,N_2761,N_2630);
nand U2892 (N_2892,N_2674,N_2665);
or U2893 (N_2893,N_2656,N_2655);
and U2894 (N_2894,N_2708,N_2613);
or U2895 (N_2895,N_2739,N_2699);
xor U2896 (N_2896,N_2760,N_2749);
and U2897 (N_2897,N_2714,N_2672);
xor U2898 (N_2898,N_2733,N_2629);
nor U2899 (N_2899,N_2756,N_2773);
xnor U2900 (N_2900,N_2649,N_2749);
nand U2901 (N_2901,N_2732,N_2747);
nand U2902 (N_2902,N_2647,N_2774);
or U2903 (N_2903,N_2708,N_2701);
xnor U2904 (N_2904,N_2718,N_2749);
and U2905 (N_2905,N_2600,N_2773);
and U2906 (N_2906,N_2690,N_2711);
or U2907 (N_2907,N_2715,N_2668);
and U2908 (N_2908,N_2760,N_2705);
xor U2909 (N_2909,N_2679,N_2665);
or U2910 (N_2910,N_2641,N_2782);
and U2911 (N_2911,N_2647,N_2762);
xor U2912 (N_2912,N_2630,N_2624);
and U2913 (N_2913,N_2741,N_2646);
nor U2914 (N_2914,N_2614,N_2794);
nor U2915 (N_2915,N_2697,N_2659);
or U2916 (N_2916,N_2604,N_2621);
or U2917 (N_2917,N_2687,N_2623);
xor U2918 (N_2918,N_2633,N_2797);
xnor U2919 (N_2919,N_2752,N_2658);
xor U2920 (N_2920,N_2716,N_2678);
or U2921 (N_2921,N_2772,N_2705);
xor U2922 (N_2922,N_2749,N_2601);
nor U2923 (N_2923,N_2764,N_2754);
nor U2924 (N_2924,N_2649,N_2795);
nand U2925 (N_2925,N_2673,N_2701);
or U2926 (N_2926,N_2709,N_2696);
xor U2927 (N_2927,N_2715,N_2730);
and U2928 (N_2928,N_2676,N_2775);
or U2929 (N_2929,N_2642,N_2670);
xor U2930 (N_2930,N_2765,N_2699);
nand U2931 (N_2931,N_2616,N_2657);
nand U2932 (N_2932,N_2643,N_2730);
nor U2933 (N_2933,N_2621,N_2697);
and U2934 (N_2934,N_2606,N_2605);
or U2935 (N_2935,N_2760,N_2609);
or U2936 (N_2936,N_2634,N_2604);
xnor U2937 (N_2937,N_2795,N_2626);
and U2938 (N_2938,N_2770,N_2602);
and U2939 (N_2939,N_2675,N_2633);
nor U2940 (N_2940,N_2716,N_2653);
nand U2941 (N_2941,N_2739,N_2630);
or U2942 (N_2942,N_2639,N_2695);
xor U2943 (N_2943,N_2661,N_2746);
xor U2944 (N_2944,N_2656,N_2722);
nand U2945 (N_2945,N_2732,N_2607);
nor U2946 (N_2946,N_2698,N_2671);
or U2947 (N_2947,N_2691,N_2758);
xnor U2948 (N_2948,N_2636,N_2726);
nand U2949 (N_2949,N_2665,N_2644);
nor U2950 (N_2950,N_2739,N_2777);
and U2951 (N_2951,N_2688,N_2648);
xor U2952 (N_2952,N_2777,N_2635);
or U2953 (N_2953,N_2695,N_2697);
and U2954 (N_2954,N_2786,N_2746);
nor U2955 (N_2955,N_2765,N_2678);
nor U2956 (N_2956,N_2703,N_2634);
xor U2957 (N_2957,N_2727,N_2730);
xnor U2958 (N_2958,N_2742,N_2757);
xnor U2959 (N_2959,N_2608,N_2650);
and U2960 (N_2960,N_2797,N_2651);
and U2961 (N_2961,N_2635,N_2751);
or U2962 (N_2962,N_2664,N_2695);
nor U2963 (N_2963,N_2648,N_2745);
xor U2964 (N_2964,N_2648,N_2652);
xor U2965 (N_2965,N_2703,N_2640);
nand U2966 (N_2966,N_2613,N_2783);
and U2967 (N_2967,N_2630,N_2786);
or U2968 (N_2968,N_2610,N_2638);
nand U2969 (N_2969,N_2775,N_2708);
nand U2970 (N_2970,N_2773,N_2784);
nand U2971 (N_2971,N_2704,N_2665);
nand U2972 (N_2972,N_2720,N_2711);
nand U2973 (N_2973,N_2679,N_2744);
xor U2974 (N_2974,N_2683,N_2638);
xor U2975 (N_2975,N_2727,N_2798);
nand U2976 (N_2976,N_2755,N_2734);
xor U2977 (N_2977,N_2716,N_2743);
or U2978 (N_2978,N_2631,N_2733);
nand U2979 (N_2979,N_2619,N_2699);
xnor U2980 (N_2980,N_2734,N_2780);
nand U2981 (N_2981,N_2784,N_2709);
nand U2982 (N_2982,N_2796,N_2748);
and U2983 (N_2983,N_2738,N_2692);
nand U2984 (N_2984,N_2603,N_2633);
and U2985 (N_2985,N_2639,N_2611);
nand U2986 (N_2986,N_2721,N_2732);
xor U2987 (N_2987,N_2767,N_2768);
and U2988 (N_2988,N_2775,N_2790);
nand U2989 (N_2989,N_2640,N_2771);
xor U2990 (N_2990,N_2614,N_2785);
nand U2991 (N_2991,N_2712,N_2670);
xnor U2992 (N_2992,N_2648,N_2617);
nor U2993 (N_2993,N_2652,N_2627);
xnor U2994 (N_2994,N_2648,N_2692);
xnor U2995 (N_2995,N_2701,N_2672);
nor U2996 (N_2996,N_2615,N_2669);
and U2997 (N_2997,N_2634,N_2765);
nor U2998 (N_2998,N_2704,N_2771);
xor U2999 (N_2999,N_2602,N_2649);
nand UO_0 (O_0,N_2983,N_2815);
or UO_1 (O_1,N_2900,N_2909);
xor UO_2 (O_2,N_2810,N_2883);
xor UO_3 (O_3,N_2886,N_2826);
and UO_4 (O_4,N_2821,N_2920);
xnor UO_5 (O_5,N_2857,N_2823);
xnor UO_6 (O_6,N_2880,N_2865);
xor UO_7 (O_7,N_2972,N_2879);
and UO_8 (O_8,N_2847,N_2873);
nor UO_9 (O_9,N_2811,N_2991);
xnor UO_10 (O_10,N_2867,N_2852);
nand UO_11 (O_11,N_2966,N_2968);
nor UO_12 (O_12,N_2990,N_2955);
xnor UO_13 (O_13,N_2925,N_2965);
nor UO_14 (O_14,N_2984,N_2914);
nor UO_15 (O_15,N_2932,N_2871);
or UO_16 (O_16,N_2818,N_2878);
and UO_17 (O_17,N_2926,N_2970);
or UO_18 (O_18,N_2858,N_2927);
xnor UO_19 (O_19,N_2830,N_2866);
xnor UO_20 (O_20,N_2902,N_2829);
xnor UO_21 (O_21,N_2989,N_2947);
xor UO_22 (O_22,N_2868,N_2837);
and UO_23 (O_23,N_2800,N_2953);
nor UO_24 (O_24,N_2940,N_2802);
xnor UO_25 (O_25,N_2828,N_2934);
or UO_26 (O_26,N_2835,N_2892);
and UO_27 (O_27,N_2938,N_2889);
and UO_28 (O_28,N_2844,N_2849);
or UO_29 (O_29,N_2806,N_2998);
xor UO_30 (O_30,N_2807,N_2924);
nand UO_31 (O_31,N_2971,N_2999);
or UO_32 (O_32,N_2948,N_2916);
xnor UO_33 (O_33,N_2822,N_2859);
or UO_34 (O_34,N_2872,N_2840);
nand UO_35 (O_35,N_2988,N_2855);
xnor UO_36 (O_36,N_2995,N_2931);
xor UO_37 (O_37,N_2817,N_2856);
nor UO_38 (O_38,N_2864,N_2941);
or UO_39 (O_39,N_2922,N_2959);
xnor UO_40 (O_40,N_2910,N_2804);
nor UO_41 (O_41,N_2895,N_2994);
xor UO_42 (O_42,N_2997,N_2976);
nor UO_43 (O_43,N_2893,N_2903);
nand UO_44 (O_44,N_2936,N_2901);
or UO_45 (O_45,N_2846,N_2967);
xnor UO_46 (O_46,N_2906,N_2841);
xor UO_47 (O_47,N_2853,N_2980);
xnor UO_48 (O_48,N_2833,N_2969);
nand UO_49 (O_49,N_2961,N_2861);
nand UO_50 (O_50,N_2915,N_2993);
or UO_51 (O_51,N_2843,N_2929);
or UO_52 (O_52,N_2836,N_2952);
xor UO_53 (O_53,N_2918,N_2928);
xnor UO_54 (O_54,N_2816,N_2832);
nor UO_55 (O_55,N_2819,N_2912);
and UO_56 (O_56,N_2875,N_2874);
nor UO_57 (O_57,N_2831,N_2882);
or UO_58 (O_58,N_2986,N_2884);
nor UO_59 (O_59,N_2950,N_2813);
nor UO_60 (O_60,N_2923,N_2917);
or UO_61 (O_61,N_2851,N_2919);
nand UO_62 (O_62,N_2964,N_2981);
or UO_63 (O_63,N_2803,N_2907);
or UO_64 (O_64,N_2942,N_2979);
and UO_65 (O_65,N_2860,N_2809);
nor UO_66 (O_66,N_2845,N_2982);
or UO_67 (O_67,N_2962,N_2992);
or UO_68 (O_68,N_2820,N_2911);
and UO_69 (O_69,N_2812,N_2869);
xor UO_70 (O_70,N_2904,N_2954);
and UO_71 (O_71,N_2963,N_2949);
nand UO_72 (O_72,N_2905,N_2943);
nor UO_73 (O_73,N_2877,N_2935);
or UO_74 (O_74,N_2985,N_2854);
nand UO_75 (O_75,N_2987,N_2978);
xor UO_76 (O_76,N_2881,N_2974);
or UO_77 (O_77,N_2946,N_2825);
nand UO_78 (O_78,N_2862,N_2956);
nor UO_79 (O_79,N_2977,N_2898);
nor UO_80 (O_80,N_2891,N_2839);
nand UO_81 (O_81,N_2908,N_2930);
or UO_82 (O_82,N_2951,N_2899);
or UO_83 (O_83,N_2827,N_2885);
or UO_84 (O_84,N_2824,N_2973);
and UO_85 (O_85,N_2834,N_2894);
nor UO_86 (O_86,N_2933,N_2848);
and UO_87 (O_87,N_2975,N_2913);
or UO_88 (O_88,N_2838,N_2960);
and UO_89 (O_89,N_2801,N_2896);
or UO_90 (O_90,N_2996,N_2814);
nor UO_91 (O_91,N_2887,N_2870);
nand UO_92 (O_92,N_2850,N_2945);
xnor UO_93 (O_93,N_2958,N_2937);
xnor UO_94 (O_94,N_2808,N_2939);
and UO_95 (O_95,N_2863,N_2876);
xor UO_96 (O_96,N_2897,N_2921);
xnor UO_97 (O_97,N_2890,N_2805);
xor UO_98 (O_98,N_2888,N_2944);
nor UO_99 (O_99,N_2842,N_2957);
nor UO_100 (O_100,N_2840,N_2858);
and UO_101 (O_101,N_2915,N_2893);
or UO_102 (O_102,N_2909,N_2908);
xnor UO_103 (O_103,N_2810,N_2880);
nor UO_104 (O_104,N_2967,N_2871);
nor UO_105 (O_105,N_2987,N_2879);
nand UO_106 (O_106,N_2813,N_2857);
and UO_107 (O_107,N_2956,N_2868);
and UO_108 (O_108,N_2810,N_2814);
xor UO_109 (O_109,N_2806,N_2844);
xor UO_110 (O_110,N_2802,N_2957);
nor UO_111 (O_111,N_2818,N_2969);
xor UO_112 (O_112,N_2987,N_2881);
xor UO_113 (O_113,N_2857,N_2835);
or UO_114 (O_114,N_2967,N_2971);
nand UO_115 (O_115,N_2807,N_2870);
or UO_116 (O_116,N_2925,N_2841);
nor UO_117 (O_117,N_2806,N_2849);
and UO_118 (O_118,N_2814,N_2950);
or UO_119 (O_119,N_2909,N_2847);
nor UO_120 (O_120,N_2949,N_2961);
and UO_121 (O_121,N_2958,N_2816);
nor UO_122 (O_122,N_2958,N_2890);
or UO_123 (O_123,N_2832,N_2976);
xnor UO_124 (O_124,N_2989,N_2984);
and UO_125 (O_125,N_2986,N_2858);
and UO_126 (O_126,N_2855,N_2953);
nor UO_127 (O_127,N_2874,N_2932);
nand UO_128 (O_128,N_2811,N_2916);
or UO_129 (O_129,N_2876,N_2950);
nand UO_130 (O_130,N_2985,N_2895);
and UO_131 (O_131,N_2991,N_2949);
nand UO_132 (O_132,N_2923,N_2899);
and UO_133 (O_133,N_2924,N_2872);
or UO_134 (O_134,N_2947,N_2958);
and UO_135 (O_135,N_2908,N_2974);
and UO_136 (O_136,N_2932,N_2925);
or UO_137 (O_137,N_2938,N_2871);
and UO_138 (O_138,N_2833,N_2850);
nand UO_139 (O_139,N_2978,N_2891);
or UO_140 (O_140,N_2823,N_2838);
xor UO_141 (O_141,N_2890,N_2860);
or UO_142 (O_142,N_2983,N_2881);
and UO_143 (O_143,N_2902,N_2826);
and UO_144 (O_144,N_2816,N_2868);
nand UO_145 (O_145,N_2930,N_2844);
nand UO_146 (O_146,N_2833,N_2865);
nor UO_147 (O_147,N_2966,N_2918);
and UO_148 (O_148,N_2827,N_2888);
xnor UO_149 (O_149,N_2820,N_2816);
nor UO_150 (O_150,N_2917,N_2857);
or UO_151 (O_151,N_2869,N_2928);
xor UO_152 (O_152,N_2950,N_2846);
or UO_153 (O_153,N_2998,N_2846);
nor UO_154 (O_154,N_2934,N_2978);
nand UO_155 (O_155,N_2802,N_2847);
or UO_156 (O_156,N_2975,N_2966);
and UO_157 (O_157,N_2826,N_2891);
xor UO_158 (O_158,N_2912,N_2851);
nor UO_159 (O_159,N_2972,N_2831);
or UO_160 (O_160,N_2959,N_2977);
nor UO_161 (O_161,N_2855,N_2937);
and UO_162 (O_162,N_2809,N_2847);
nand UO_163 (O_163,N_2831,N_2912);
and UO_164 (O_164,N_2894,N_2911);
or UO_165 (O_165,N_2984,N_2834);
xnor UO_166 (O_166,N_2863,N_2858);
and UO_167 (O_167,N_2960,N_2803);
and UO_168 (O_168,N_2881,N_2954);
nand UO_169 (O_169,N_2879,N_2844);
nor UO_170 (O_170,N_2859,N_2871);
nand UO_171 (O_171,N_2864,N_2838);
and UO_172 (O_172,N_2822,N_2957);
and UO_173 (O_173,N_2888,N_2994);
and UO_174 (O_174,N_2920,N_2918);
nor UO_175 (O_175,N_2975,N_2815);
nor UO_176 (O_176,N_2912,N_2892);
nor UO_177 (O_177,N_2942,N_2801);
nand UO_178 (O_178,N_2956,N_2978);
nand UO_179 (O_179,N_2931,N_2919);
or UO_180 (O_180,N_2817,N_2804);
or UO_181 (O_181,N_2903,N_2974);
and UO_182 (O_182,N_2935,N_2852);
and UO_183 (O_183,N_2907,N_2824);
nor UO_184 (O_184,N_2920,N_2948);
xor UO_185 (O_185,N_2853,N_2911);
xnor UO_186 (O_186,N_2810,N_2881);
nor UO_187 (O_187,N_2928,N_2805);
nor UO_188 (O_188,N_2957,N_2803);
or UO_189 (O_189,N_2921,N_2813);
xnor UO_190 (O_190,N_2914,N_2833);
xor UO_191 (O_191,N_2992,N_2837);
nor UO_192 (O_192,N_2991,N_2851);
nor UO_193 (O_193,N_2975,N_2988);
or UO_194 (O_194,N_2862,N_2918);
or UO_195 (O_195,N_2802,N_2939);
and UO_196 (O_196,N_2810,N_2821);
nand UO_197 (O_197,N_2808,N_2902);
or UO_198 (O_198,N_2849,N_2901);
nand UO_199 (O_199,N_2909,N_2813);
nand UO_200 (O_200,N_2980,N_2883);
xnor UO_201 (O_201,N_2955,N_2931);
or UO_202 (O_202,N_2944,N_2833);
nand UO_203 (O_203,N_2805,N_2860);
xnor UO_204 (O_204,N_2860,N_2996);
and UO_205 (O_205,N_2998,N_2864);
xnor UO_206 (O_206,N_2927,N_2951);
nand UO_207 (O_207,N_2827,N_2802);
xnor UO_208 (O_208,N_2996,N_2806);
xnor UO_209 (O_209,N_2874,N_2809);
nand UO_210 (O_210,N_2841,N_2983);
nor UO_211 (O_211,N_2844,N_2966);
nand UO_212 (O_212,N_2974,N_2863);
nand UO_213 (O_213,N_2913,N_2881);
xor UO_214 (O_214,N_2906,N_2813);
or UO_215 (O_215,N_2919,N_2856);
nor UO_216 (O_216,N_2919,N_2812);
xor UO_217 (O_217,N_2908,N_2963);
xor UO_218 (O_218,N_2897,N_2982);
or UO_219 (O_219,N_2919,N_2984);
nor UO_220 (O_220,N_2806,N_2868);
and UO_221 (O_221,N_2847,N_2905);
or UO_222 (O_222,N_2928,N_2822);
and UO_223 (O_223,N_2898,N_2991);
or UO_224 (O_224,N_2861,N_2951);
nand UO_225 (O_225,N_2914,N_2997);
nand UO_226 (O_226,N_2811,N_2945);
xor UO_227 (O_227,N_2880,N_2824);
nand UO_228 (O_228,N_2825,N_2985);
and UO_229 (O_229,N_2877,N_2879);
or UO_230 (O_230,N_2954,N_2988);
xor UO_231 (O_231,N_2942,N_2943);
and UO_232 (O_232,N_2800,N_2933);
and UO_233 (O_233,N_2890,N_2910);
nor UO_234 (O_234,N_2935,N_2837);
or UO_235 (O_235,N_2882,N_2929);
and UO_236 (O_236,N_2896,N_2805);
nand UO_237 (O_237,N_2886,N_2883);
xnor UO_238 (O_238,N_2994,N_2826);
nor UO_239 (O_239,N_2886,N_2837);
nor UO_240 (O_240,N_2910,N_2994);
and UO_241 (O_241,N_2897,N_2959);
xor UO_242 (O_242,N_2872,N_2936);
or UO_243 (O_243,N_2969,N_2806);
and UO_244 (O_244,N_2917,N_2959);
xor UO_245 (O_245,N_2951,N_2818);
or UO_246 (O_246,N_2820,N_2842);
nand UO_247 (O_247,N_2976,N_2828);
or UO_248 (O_248,N_2808,N_2910);
xor UO_249 (O_249,N_2874,N_2931);
or UO_250 (O_250,N_2821,N_2942);
and UO_251 (O_251,N_2918,N_2968);
nand UO_252 (O_252,N_2865,N_2923);
or UO_253 (O_253,N_2979,N_2995);
nand UO_254 (O_254,N_2930,N_2994);
or UO_255 (O_255,N_2867,N_2821);
nor UO_256 (O_256,N_2892,N_2909);
or UO_257 (O_257,N_2834,N_2865);
nand UO_258 (O_258,N_2992,N_2806);
and UO_259 (O_259,N_2835,N_2948);
nor UO_260 (O_260,N_2977,N_2936);
nand UO_261 (O_261,N_2937,N_2902);
nor UO_262 (O_262,N_2970,N_2856);
nand UO_263 (O_263,N_2845,N_2910);
and UO_264 (O_264,N_2902,N_2947);
and UO_265 (O_265,N_2838,N_2867);
or UO_266 (O_266,N_2985,N_2957);
xnor UO_267 (O_267,N_2977,N_2882);
and UO_268 (O_268,N_2808,N_2963);
nor UO_269 (O_269,N_2996,N_2822);
xnor UO_270 (O_270,N_2931,N_2866);
or UO_271 (O_271,N_2958,N_2959);
nor UO_272 (O_272,N_2997,N_2934);
nor UO_273 (O_273,N_2845,N_2942);
and UO_274 (O_274,N_2941,N_2867);
xor UO_275 (O_275,N_2952,N_2964);
nand UO_276 (O_276,N_2981,N_2941);
nand UO_277 (O_277,N_2993,N_2834);
nor UO_278 (O_278,N_2888,N_2998);
nand UO_279 (O_279,N_2946,N_2822);
and UO_280 (O_280,N_2954,N_2834);
and UO_281 (O_281,N_2821,N_2851);
and UO_282 (O_282,N_2982,N_2948);
xor UO_283 (O_283,N_2907,N_2827);
nand UO_284 (O_284,N_2975,N_2931);
xnor UO_285 (O_285,N_2801,N_2867);
nand UO_286 (O_286,N_2804,N_2816);
or UO_287 (O_287,N_2900,N_2978);
nor UO_288 (O_288,N_2804,N_2846);
xor UO_289 (O_289,N_2903,N_2975);
nor UO_290 (O_290,N_2883,N_2806);
or UO_291 (O_291,N_2828,N_2930);
xor UO_292 (O_292,N_2915,N_2839);
and UO_293 (O_293,N_2969,N_2897);
nor UO_294 (O_294,N_2929,N_2856);
xor UO_295 (O_295,N_2873,N_2885);
and UO_296 (O_296,N_2956,N_2927);
and UO_297 (O_297,N_2871,N_2874);
or UO_298 (O_298,N_2924,N_2864);
or UO_299 (O_299,N_2907,N_2968);
nand UO_300 (O_300,N_2894,N_2945);
xor UO_301 (O_301,N_2995,N_2847);
xor UO_302 (O_302,N_2856,N_2860);
nor UO_303 (O_303,N_2960,N_2864);
nand UO_304 (O_304,N_2895,N_2954);
or UO_305 (O_305,N_2817,N_2921);
nand UO_306 (O_306,N_2842,N_2824);
and UO_307 (O_307,N_2990,N_2918);
nand UO_308 (O_308,N_2875,N_2977);
xor UO_309 (O_309,N_2985,N_2950);
and UO_310 (O_310,N_2958,N_2801);
xnor UO_311 (O_311,N_2859,N_2854);
xor UO_312 (O_312,N_2945,N_2973);
nand UO_313 (O_313,N_2803,N_2984);
nand UO_314 (O_314,N_2811,N_2816);
nand UO_315 (O_315,N_2929,N_2921);
nand UO_316 (O_316,N_2953,N_2886);
or UO_317 (O_317,N_2978,N_2880);
and UO_318 (O_318,N_2860,N_2895);
nand UO_319 (O_319,N_2970,N_2937);
xor UO_320 (O_320,N_2962,N_2873);
nand UO_321 (O_321,N_2836,N_2983);
or UO_322 (O_322,N_2908,N_2835);
and UO_323 (O_323,N_2839,N_2905);
and UO_324 (O_324,N_2983,N_2921);
nor UO_325 (O_325,N_2894,N_2985);
xnor UO_326 (O_326,N_2979,N_2855);
nand UO_327 (O_327,N_2970,N_2981);
and UO_328 (O_328,N_2818,N_2889);
or UO_329 (O_329,N_2854,N_2981);
nor UO_330 (O_330,N_2906,N_2925);
nand UO_331 (O_331,N_2984,N_2986);
xnor UO_332 (O_332,N_2833,N_2866);
nor UO_333 (O_333,N_2918,N_2907);
nand UO_334 (O_334,N_2856,N_2903);
and UO_335 (O_335,N_2866,N_2945);
xor UO_336 (O_336,N_2922,N_2881);
nor UO_337 (O_337,N_2812,N_2908);
or UO_338 (O_338,N_2931,N_2850);
or UO_339 (O_339,N_2930,N_2839);
nor UO_340 (O_340,N_2950,N_2856);
and UO_341 (O_341,N_2822,N_2837);
nor UO_342 (O_342,N_2947,N_2982);
and UO_343 (O_343,N_2962,N_2951);
xnor UO_344 (O_344,N_2827,N_2818);
and UO_345 (O_345,N_2890,N_2983);
xnor UO_346 (O_346,N_2846,N_2839);
nor UO_347 (O_347,N_2991,N_2820);
nand UO_348 (O_348,N_2881,N_2886);
nor UO_349 (O_349,N_2917,N_2983);
xor UO_350 (O_350,N_2920,N_2926);
xor UO_351 (O_351,N_2970,N_2892);
nand UO_352 (O_352,N_2942,N_2896);
nor UO_353 (O_353,N_2867,N_2913);
xnor UO_354 (O_354,N_2818,N_2846);
nand UO_355 (O_355,N_2979,N_2937);
nor UO_356 (O_356,N_2934,N_2890);
xor UO_357 (O_357,N_2868,N_2989);
nand UO_358 (O_358,N_2890,N_2914);
xor UO_359 (O_359,N_2989,N_2979);
and UO_360 (O_360,N_2840,N_2969);
nor UO_361 (O_361,N_2994,N_2917);
or UO_362 (O_362,N_2941,N_2820);
xor UO_363 (O_363,N_2987,N_2869);
nand UO_364 (O_364,N_2931,N_2949);
and UO_365 (O_365,N_2922,N_2966);
nor UO_366 (O_366,N_2886,N_2936);
or UO_367 (O_367,N_2861,N_2903);
and UO_368 (O_368,N_2824,N_2918);
nor UO_369 (O_369,N_2855,N_2907);
nand UO_370 (O_370,N_2869,N_2942);
and UO_371 (O_371,N_2934,N_2885);
and UO_372 (O_372,N_2905,N_2946);
nor UO_373 (O_373,N_2982,N_2959);
and UO_374 (O_374,N_2885,N_2944);
or UO_375 (O_375,N_2989,N_2933);
nand UO_376 (O_376,N_2843,N_2953);
nand UO_377 (O_377,N_2824,N_2863);
nand UO_378 (O_378,N_2941,N_2958);
nand UO_379 (O_379,N_2854,N_2901);
nor UO_380 (O_380,N_2946,N_2971);
nor UO_381 (O_381,N_2806,N_2929);
nand UO_382 (O_382,N_2991,N_2819);
xnor UO_383 (O_383,N_2950,N_2919);
and UO_384 (O_384,N_2973,N_2842);
or UO_385 (O_385,N_2927,N_2811);
and UO_386 (O_386,N_2892,N_2895);
xor UO_387 (O_387,N_2955,N_2921);
nor UO_388 (O_388,N_2869,N_2930);
and UO_389 (O_389,N_2812,N_2877);
nor UO_390 (O_390,N_2864,N_2927);
xor UO_391 (O_391,N_2990,N_2871);
or UO_392 (O_392,N_2843,N_2971);
nor UO_393 (O_393,N_2922,N_2896);
nor UO_394 (O_394,N_2906,N_2885);
nand UO_395 (O_395,N_2844,N_2936);
nand UO_396 (O_396,N_2882,N_2950);
nand UO_397 (O_397,N_2999,N_2961);
or UO_398 (O_398,N_2962,N_2921);
nor UO_399 (O_399,N_2853,N_2890);
nand UO_400 (O_400,N_2814,N_2894);
nor UO_401 (O_401,N_2968,N_2960);
or UO_402 (O_402,N_2974,N_2873);
xor UO_403 (O_403,N_2969,N_2814);
nand UO_404 (O_404,N_2800,N_2897);
nor UO_405 (O_405,N_2821,N_2883);
nand UO_406 (O_406,N_2883,N_2956);
or UO_407 (O_407,N_2883,N_2837);
or UO_408 (O_408,N_2846,N_2986);
nand UO_409 (O_409,N_2892,N_2978);
nor UO_410 (O_410,N_2902,N_2801);
or UO_411 (O_411,N_2995,N_2825);
or UO_412 (O_412,N_2847,N_2845);
xnor UO_413 (O_413,N_2916,N_2883);
xnor UO_414 (O_414,N_2993,N_2886);
and UO_415 (O_415,N_2987,N_2807);
nor UO_416 (O_416,N_2944,N_2844);
xnor UO_417 (O_417,N_2933,N_2871);
nor UO_418 (O_418,N_2844,N_2918);
nor UO_419 (O_419,N_2889,N_2883);
and UO_420 (O_420,N_2989,N_2985);
or UO_421 (O_421,N_2894,N_2959);
or UO_422 (O_422,N_2954,N_2920);
or UO_423 (O_423,N_2917,N_2957);
xnor UO_424 (O_424,N_2835,N_2938);
xnor UO_425 (O_425,N_2977,N_2845);
and UO_426 (O_426,N_2871,N_2919);
and UO_427 (O_427,N_2904,N_2992);
nand UO_428 (O_428,N_2896,N_2858);
xor UO_429 (O_429,N_2928,N_2944);
xor UO_430 (O_430,N_2853,N_2846);
and UO_431 (O_431,N_2869,N_2863);
nand UO_432 (O_432,N_2875,N_2954);
or UO_433 (O_433,N_2949,N_2877);
or UO_434 (O_434,N_2887,N_2988);
nand UO_435 (O_435,N_2822,N_2983);
xor UO_436 (O_436,N_2839,N_2898);
xnor UO_437 (O_437,N_2883,N_2812);
nor UO_438 (O_438,N_2940,N_2880);
nand UO_439 (O_439,N_2870,N_2810);
nor UO_440 (O_440,N_2984,N_2966);
nand UO_441 (O_441,N_2874,N_2837);
nand UO_442 (O_442,N_2807,N_2904);
xor UO_443 (O_443,N_2850,N_2915);
nor UO_444 (O_444,N_2830,N_2900);
nor UO_445 (O_445,N_2967,N_2896);
xor UO_446 (O_446,N_2901,N_2927);
nand UO_447 (O_447,N_2880,N_2877);
xnor UO_448 (O_448,N_2828,N_2905);
nand UO_449 (O_449,N_2919,N_2820);
nand UO_450 (O_450,N_2919,N_2864);
nand UO_451 (O_451,N_2893,N_2921);
or UO_452 (O_452,N_2944,N_2899);
and UO_453 (O_453,N_2852,N_2926);
nor UO_454 (O_454,N_2901,N_2843);
and UO_455 (O_455,N_2990,N_2811);
or UO_456 (O_456,N_2946,N_2982);
or UO_457 (O_457,N_2994,N_2865);
or UO_458 (O_458,N_2880,N_2905);
or UO_459 (O_459,N_2897,N_2812);
nor UO_460 (O_460,N_2857,N_2815);
nor UO_461 (O_461,N_2880,N_2847);
and UO_462 (O_462,N_2934,N_2872);
or UO_463 (O_463,N_2841,N_2854);
or UO_464 (O_464,N_2998,N_2844);
xnor UO_465 (O_465,N_2922,N_2879);
nor UO_466 (O_466,N_2890,N_2953);
or UO_467 (O_467,N_2853,N_2845);
and UO_468 (O_468,N_2811,N_2842);
nand UO_469 (O_469,N_2972,N_2814);
and UO_470 (O_470,N_2988,N_2925);
and UO_471 (O_471,N_2820,N_2863);
and UO_472 (O_472,N_2995,N_2854);
xor UO_473 (O_473,N_2851,N_2885);
xor UO_474 (O_474,N_2976,N_2859);
and UO_475 (O_475,N_2820,N_2818);
or UO_476 (O_476,N_2839,N_2874);
nand UO_477 (O_477,N_2820,N_2938);
and UO_478 (O_478,N_2981,N_2804);
nand UO_479 (O_479,N_2885,N_2956);
xnor UO_480 (O_480,N_2845,N_2848);
xnor UO_481 (O_481,N_2960,N_2816);
nand UO_482 (O_482,N_2966,N_2917);
and UO_483 (O_483,N_2953,N_2958);
nor UO_484 (O_484,N_2928,N_2982);
nand UO_485 (O_485,N_2811,N_2845);
nand UO_486 (O_486,N_2820,N_2862);
xnor UO_487 (O_487,N_2844,N_2997);
and UO_488 (O_488,N_2904,N_2836);
nor UO_489 (O_489,N_2871,N_2970);
nand UO_490 (O_490,N_2977,N_2958);
nor UO_491 (O_491,N_2881,N_2840);
xor UO_492 (O_492,N_2822,N_2810);
or UO_493 (O_493,N_2931,N_2827);
and UO_494 (O_494,N_2856,N_2901);
and UO_495 (O_495,N_2873,N_2825);
or UO_496 (O_496,N_2803,N_2992);
and UO_497 (O_497,N_2903,N_2967);
nand UO_498 (O_498,N_2901,N_2860);
and UO_499 (O_499,N_2834,N_2887);
endmodule