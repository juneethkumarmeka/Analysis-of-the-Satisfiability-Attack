module basic_500_3000_500_15_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_67,In_473);
and U1 (N_1,In_25,In_455);
and U2 (N_2,In_161,In_418);
nand U3 (N_3,In_322,In_163);
xor U4 (N_4,In_485,In_118);
and U5 (N_5,In_413,In_3);
nand U6 (N_6,In_289,In_444);
nand U7 (N_7,In_198,In_35);
or U8 (N_8,In_157,In_23);
nor U9 (N_9,In_63,In_184);
nor U10 (N_10,In_371,In_320);
and U11 (N_11,In_292,In_471);
or U12 (N_12,In_120,In_366);
or U13 (N_13,In_260,In_158);
or U14 (N_14,In_297,In_137);
nand U15 (N_15,In_1,In_79);
nor U16 (N_16,In_486,In_232);
nor U17 (N_17,In_469,In_385);
nand U18 (N_18,In_380,In_150);
nor U19 (N_19,In_328,In_41);
and U20 (N_20,In_337,In_99);
and U21 (N_21,In_262,In_356);
nand U22 (N_22,In_64,In_465);
or U23 (N_23,In_110,In_340);
nand U24 (N_24,In_296,In_325);
or U25 (N_25,In_362,In_414);
nor U26 (N_26,In_56,In_330);
or U27 (N_27,In_182,In_169);
nor U28 (N_28,In_281,In_111);
nor U29 (N_29,In_311,In_131);
or U30 (N_30,In_482,In_445);
and U31 (N_31,In_172,In_404);
or U32 (N_32,In_399,In_442);
nand U33 (N_33,In_238,In_176);
and U34 (N_34,In_321,In_152);
nand U35 (N_35,In_87,In_217);
nor U36 (N_36,In_353,In_187);
and U37 (N_37,In_211,In_171);
nand U38 (N_38,In_141,In_31);
nand U39 (N_39,In_419,In_436);
nor U40 (N_40,In_167,In_367);
or U41 (N_41,In_364,In_22);
or U42 (N_42,In_140,In_345);
and U43 (N_43,In_4,In_411);
nor U44 (N_44,In_253,In_219);
or U45 (N_45,In_74,In_178);
nor U46 (N_46,In_375,In_492);
nor U47 (N_47,In_452,In_153);
or U48 (N_48,In_11,In_271);
nor U49 (N_49,In_410,In_477);
nor U50 (N_50,In_72,In_218);
or U51 (N_51,In_123,In_180);
or U52 (N_52,In_236,In_9);
and U53 (N_53,In_258,In_332);
and U54 (N_54,In_96,In_261);
and U55 (N_55,In_208,In_193);
nor U56 (N_56,In_323,In_498);
and U57 (N_57,In_499,In_82);
and U58 (N_58,In_472,In_339);
nor U59 (N_59,In_183,In_464);
or U60 (N_60,In_144,In_265);
xnor U61 (N_61,In_34,In_421);
and U62 (N_62,In_359,In_426);
nor U63 (N_63,In_57,In_300);
nor U64 (N_64,In_448,In_207);
or U65 (N_65,In_268,In_173);
or U66 (N_66,In_495,In_13);
or U67 (N_67,In_346,In_372);
nand U68 (N_68,In_494,In_122);
and U69 (N_69,In_331,In_308);
and U70 (N_70,In_14,In_68);
nor U71 (N_71,In_139,In_350);
nor U72 (N_72,In_407,In_59);
and U73 (N_73,In_454,In_203);
and U74 (N_74,In_453,In_192);
nor U75 (N_75,In_347,In_391);
nor U76 (N_76,In_143,In_97);
nor U77 (N_77,In_46,In_389);
nand U78 (N_78,In_269,In_303);
or U79 (N_79,In_12,In_306);
nor U80 (N_80,In_263,In_428);
or U81 (N_81,In_257,In_388);
nor U82 (N_82,In_133,In_291);
nor U83 (N_83,In_222,In_149);
nor U84 (N_84,In_361,In_138);
nor U85 (N_85,In_231,In_147);
nand U86 (N_86,In_316,In_496);
nand U87 (N_87,In_483,In_216);
and U88 (N_88,In_73,In_27);
or U89 (N_89,In_66,In_225);
nand U90 (N_90,In_33,In_435);
nand U91 (N_91,In_80,In_415);
and U92 (N_92,In_287,In_214);
nor U93 (N_93,In_199,In_466);
and U94 (N_94,In_497,In_313);
or U95 (N_95,In_181,In_145);
nor U96 (N_96,In_201,In_318);
or U97 (N_97,In_405,In_94);
or U98 (N_98,In_427,In_294);
and U99 (N_99,In_85,In_491);
and U100 (N_100,In_451,In_44);
and U101 (N_101,In_69,In_26);
nor U102 (N_102,In_83,In_425);
nand U103 (N_103,In_305,In_342);
nor U104 (N_104,In_283,In_196);
nand U105 (N_105,In_127,In_100);
nand U106 (N_106,In_285,In_103);
and U107 (N_107,In_241,In_159);
nand U108 (N_108,In_278,In_395);
nor U109 (N_109,In_351,In_107);
nand U110 (N_110,In_259,In_186);
or U111 (N_111,In_90,In_459);
nand U112 (N_112,In_280,In_106);
or U113 (N_113,In_0,In_156);
nor U114 (N_114,In_252,In_130);
or U115 (N_115,In_16,In_476);
or U116 (N_116,In_277,In_195);
and U117 (N_117,In_368,In_490);
nor U118 (N_118,In_148,In_406);
nor U119 (N_119,In_95,In_117);
and U120 (N_120,In_166,In_71);
or U121 (N_121,In_125,In_124);
and U122 (N_122,In_250,In_88);
nor U123 (N_123,In_478,In_333);
nor U124 (N_124,In_164,In_51);
and U125 (N_125,In_417,In_461);
nand U126 (N_126,In_481,In_474);
nand U127 (N_127,In_105,In_228);
or U128 (N_128,In_457,In_432);
or U129 (N_129,In_394,In_55);
nand U130 (N_130,In_112,In_142);
and U131 (N_131,In_443,In_370);
or U132 (N_132,In_2,In_319);
and U133 (N_133,In_273,In_215);
and U134 (N_134,In_488,In_403);
nand U135 (N_135,In_61,In_266);
nor U136 (N_136,In_28,In_248);
or U137 (N_137,In_191,In_160);
and U138 (N_138,In_449,In_352);
or U139 (N_139,In_376,In_37);
or U140 (N_140,In_212,In_204);
or U141 (N_141,In_47,In_48);
nand U142 (N_142,In_479,In_98);
nand U143 (N_143,In_363,In_200);
xor U144 (N_144,In_326,In_240);
nand U145 (N_145,In_402,In_116);
or U146 (N_146,In_274,In_447);
and U147 (N_147,In_54,In_121);
nor U148 (N_148,In_396,In_36);
nor U149 (N_149,In_489,In_17);
nand U150 (N_150,In_202,In_315);
and U151 (N_151,In_354,In_119);
or U152 (N_152,In_314,In_256);
nor U153 (N_153,In_423,In_302);
nand U154 (N_154,In_18,In_179);
nor U155 (N_155,In_102,In_190);
nor U156 (N_156,In_234,In_21);
or U157 (N_157,In_440,In_189);
nor U158 (N_158,In_185,In_8);
and U159 (N_159,In_358,In_329);
nand U160 (N_160,In_335,In_114);
xnor U161 (N_161,In_272,In_374);
nand U162 (N_162,In_456,In_438);
and U163 (N_163,In_397,In_60);
nand U164 (N_164,In_101,In_227);
nor U165 (N_165,In_40,In_378);
nand U166 (N_166,In_434,In_175);
or U167 (N_167,In_43,In_424);
nor U168 (N_168,In_484,In_386);
nand U169 (N_169,In_249,In_151);
and U170 (N_170,In_188,In_134);
and U171 (N_171,In_229,In_53);
nand U172 (N_172,In_267,In_230);
or U173 (N_173,In_298,In_460);
or U174 (N_174,In_6,In_246);
and U175 (N_175,In_282,In_15);
nand U176 (N_176,In_70,In_416);
and U177 (N_177,In_392,In_220);
and U178 (N_178,In_480,In_341);
nor U179 (N_179,In_429,In_19);
xnor U180 (N_180,In_467,In_221);
and U181 (N_181,In_324,In_462);
and U182 (N_182,In_334,In_242);
nor U183 (N_183,In_412,In_433);
or U184 (N_184,In_194,In_365);
nor U185 (N_185,In_463,In_113);
and U186 (N_186,In_20,In_146);
or U187 (N_187,In_369,In_84);
and U188 (N_188,In_45,In_154);
or U189 (N_189,In_487,In_468);
nand U190 (N_190,In_128,In_210);
or U191 (N_191,In_81,In_309);
nor U192 (N_192,In_49,In_244);
nor U193 (N_193,In_77,In_93);
nor U194 (N_194,In_129,In_408);
nor U195 (N_195,In_243,In_286);
or U196 (N_196,In_30,In_39);
and U197 (N_197,In_270,In_205);
nand U198 (N_198,In_177,In_317);
xor U199 (N_199,In_360,In_247);
nor U200 (N_200,N_184,N_108);
and U201 (N_201,N_46,In_115);
and U202 (N_202,N_69,N_85);
nand U203 (N_203,N_188,N_111);
or U204 (N_204,N_3,In_239);
and U205 (N_205,N_38,N_47);
xor U206 (N_206,N_35,In_162);
and U207 (N_207,In_295,In_336);
and U208 (N_208,In_379,N_187);
nor U209 (N_209,N_83,N_0);
and U210 (N_210,N_80,In_223);
and U211 (N_211,N_197,N_75);
nand U212 (N_212,In_155,In_381);
or U213 (N_213,N_63,N_37);
and U214 (N_214,N_32,N_150);
nor U215 (N_215,N_152,N_164);
nor U216 (N_216,In_255,In_275);
nand U217 (N_217,N_15,N_89);
and U218 (N_218,In_89,N_42);
or U219 (N_219,N_186,N_168);
nor U220 (N_220,N_24,N_29);
nand U221 (N_221,In_126,N_16);
or U222 (N_222,N_76,In_450);
nor U223 (N_223,N_122,N_10);
and U224 (N_224,In_304,N_78);
or U225 (N_225,N_178,N_56);
and U226 (N_226,In_58,N_128);
and U227 (N_227,N_171,N_86);
nand U228 (N_228,N_182,In_279);
nor U229 (N_229,N_130,N_14);
nor U230 (N_230,In_135,In_5);
or U231 (N_231,N_17,In_344);
and U232 (N_232,N_88,N_191);
nor U233 (N_233,N_174,N_157);
and U234 (N_234,N_121,In_206);
nor U235 (N_235,N_31,In_470);
or U236 (N_236,N_146,In_86);
and U237 (N_237,N_7,In_233);
nor U238 (N_238,N_161,N_57);
nor U239 (N_239,In_245,N_93);
or U240 (N_240,N_50,In_393);
nand U241 (N_241,N_94,N_199);
nand U242 (N_242,In_197,N_68);
nor U243 (N_243,In_446,N_156);
or U244 (N_244,N_153,N_170);
or U245 (N_245,N_166,N_21);
nand U246 (N_246,In_355,In_431);
nand U247 (N_247,In_109,In_288);
nand U248 (N_248,In_276,N_2);
nor U249 (N_249,N_11,In_338);
nor U250 (N_250,N_142,N_72);
nand U251 (N_251,N_81,N_34);
and U252 (N_252,N_192,In_290);
and U253 (N_253,N_95,In_398);
or U254 (N_254,In_390,In_493);
nor U255 (N_255,In_29,In_382);
or U256 (N_256,N_52,N_101);
or U257 (N_257,N_79,N_43);
nand U258 (N_258,N_6,In_458);
or U259 (N_259,N_145,N_129);
and U260 (N_260,In_400,N_20);
and U261 (N_261,N_99,N_112);
nor U262 (N_262,N_148,In_373);
and U263 (N_263,In_430,In_213);
or U264 (N_264,N_109,N_74);
and U265 (N_265,N_139,In_136);
nand U266 (N_266,N_8,N_127);
or U267 (N_267,N_97,N_123);
nor U268 (N_268,In_32,N_5);
and U269 (N_269,In_420,N_58);
or U270 (N_270,In_254,In_42);
nand U271 (N_271,N_159,N_117);
nor U272 (N_272,N_60,N_177);
nor U273 (N_273,N_92,N_90);
and U274 (N_274,In_422,N_110);
nor U275 (N_275,In_174,N_71);
nor U276 (N_276,In_357,N_96);
nand U277 (N_277,In_312,N_67);
or U278 (N_278,N_66,N_158);
nand U279 (N_279,N_160,In_293);
nand U280 (N_280,N_106,N_82);
nand U281 (N_281,N_61,N_180);
nand U282 (N_282,N_40,N_126);
or U283 (N_283,N_39,In_75);
and U284 (N_284,N_91,N_183);
and U285 (N_285,In_384,In_349);
or U286 (N_286,In_38,N_19);
nand U287 (N_287,N_113,N_100);
nand U288 (N_288,N_9,N_167);
and U289 (N_289,N_194,N_22);
and U290 (N_290,In_52,N_132);
nor U291 (N_291,N_62,In_92);
and U292 (N_292,In_441,In_76);
and U293 (N_293,N_172,N_54);
nand U294 (N_294,N_143,N_135);
nor U295 (N_295,N_163,N_103);
and U296 (N_296,In_251,N_149);
and U297 (N_297,N_51,N_53);
nand U298 (N_298,N_45,In_7);
nor U299 (N_299,In_235,N_84);
or U300 (N_300,N_162,In_264);
or U301 (N_301,In_165,In_439);
or U302 (N_302,N_136,In_307);
nand U303 (N_303,In_284,N_176);
nand U304 (N_304,In_401,In_168);
nor U305 (N_305,N_147,N_144);
nand U306 (N_306,In_104,In_327);
nand U307 (N_307,N_1,N_190);
or U308 (N_308,N_64,In_310);
nor U309 (N_309,N_131,N_124);
nor U310 (N_310,In_377,N_175);
and U311 (N_311,N_138,In_224);
or U312 (N_312,N_102,N_195);
nor U313 (N_313,N_70,In_475);
or U314 (N_314,N_115,N_119);
and U315 (N_315,N_151,N_116);
nand U316 (N_316,In_383,N_196);
and U317 (N_317,N_59,N_137);
and U318 (N_318,N_118,N_105);
nand U319 (N_319,N_36,N_154);
or U320 (N_320,N_193,N_41);
and U321 (N_321,N_13,N_155);
and U322 (N_322,In_65,N_125);
nand U323 (N_323,N_65,In_343);
nand U324 (N_324,N_12,N_87);
nor U325 (N_325,In_209,N_169);
nand U326 (N_326,N_26,N_120);
or U327 (N_327,N_140,N_18);
and U328 (N_328,In_301,N_73);
nor U329 (N_329,In_132,N_28);
nor U330 (N_330,N_49,N_98);
and U331 (N_331,N_107,N_44);
nand U332 (N_332,In_170,N_33);
nor U333 (N_333,In_108,N_185);
or U334 (N_334,N_55,N_181);
nor U335 (N_335,In_226,In_62);
nor U336 (N_336,N_133,N_30);
nand U337 (N_337,N_114,In_10);
nand U338 (N_338,In_237,In_50);
nor U339 (N_339,In_437,N_165);
nand U340 (N_340,In_78,N_77);
or U341 (N_341,N_4,N_198);
or U342 (N_342,In_409,N_141);
nand U343 (N_343,In_91,N_48);
and U344 (N_344,N_173,N_23);
and U345 (N_345,N_27,N_189);
or U346 (N_346,N_104,N_25);
and U347 (N_347,In_299,N_134);
nand U348 (N_348,In_387,In_348);
nor U349 (N_349,N_179,In_24);
nor U350 (N_350,In_470,In_276);
and U351 (N_351,N_85,N_45);
nor U352 (N_352,In_251,In_312);
and U353 (N_353,In_29,N_164);
nand U354 (N_354,In_38,N_76);
xnor U355 (N_355,In_390,In_206);
and U356 (N_356,N_181,In_5);
or U357 (N_357,N_39,N_148);
or U358 (N_358,In_233,In_235);
nand U359 (N_359,N_35,In_450);
and U360 (N_360,In_104,In_409);
nor U361 (N_361,N_16,In_91);
and U362 (N_362,N_106,N_140);
nor U363 (N_363,In_226,N_22);
nand U364 (N_364,N_185,In_381);
nand U365 (N_365,In_295,N_180);
nand U366 (N_366,In_162,N_117);
nand U367 (N_367,N_129,N_53);
nor U368 (N_368,N_81,In_379);
and U369 (N_369,N_138,N_113);
and U370 (N_370,In_422,N_42);
or U371 (N_371,N_75,In_422);
and U372 (N_372,N_136,In_132);
or U373 (N_373,N_4,N_21);
or U374 (N_374,In_284,N_47);
and U375 (N_375,In_437,N_194);
and U376 (N_376,N_191,N_173);
nor U377 (N_377,N_175,N_148);
nor U378 (N_378,N_51,In_310);
or U379 (N_379,N_36,N_137);
and U380 (N_380,N_195,N_88);
or U381 (N_381,N_19,In_165);
or U382 (N_382,In_65,In_343);
nand U383 (N_383,N_187,In_401);
nand U384 (N_384,N_56,N_187);
nand U385 (N_385,N_91,In_29);
and U386 (N_386,In_377,N_44);
nand U387 (N_387,N_44,In_50);
and U388 (N_388,N_90,N_12);
and U389 (N_389,In_162,N_74);
or U390 (N_390,In_38,N_184);
nand U391 (N_391,In_301,N_144);
or U392 (N_392,N_56,In_108);
and U393 (N_393,N_138,In_383);
nor U394 (N_394,N_79,N_98);
and U395 (N_395,In_383,In_65);
xnor U396 (N_396,N_151,N_141);
nor U397 (N_397,N_14,In_245);
nand U398 (N_398,N_161,N_0);
or U399 (N_399,N_88,In_29);
nor U400 (N_400,N_215,N_255);
or U401 (N_401,N_367,N_276);
or U402 (N_402,N_204,N_241);
nor U403 (N_403,N_294,N_214);
nor U404 (N_404,N_351,N_232);
nor U405 (N_405,N_311,N_314);
or U406 (N_406,N_397,N_243);
and U407 (N_407,N_343,N_331);
and U408 (N_408,N_315,N_258);
xnor U409 (N_409,N_309,N_233);
and U410 (N_410,N_247,N_285);
and U411 (N_411,N_270,N_272);
or U412 (N_412,N_226,N_235);
nor U413 (N_413,N_395,N_332);
and U414 (N_414,N_213,N_236);
or U415 (N_415,N_288,N_375);
or U416 (N_416,N_246,N_324);
and U417 (N_417,N_269,N_290);
or U418 (N_418,N_257,N_363);
nor U419 (N_419,N_326,N_302);
nor U420 (N_420,N_387,N_208);
and U421 (N_421,N_299,N_330);
or U422 (N_422,N_220,N_229);
or U423 (N_423,N_383,N_200);
and U424 (N_424,N_202,N_225);
or U425 (N_425,N_273,N_211);
and U426 (N_426,N_339,N_237);
and U427 (N_427,N_371,N_364);
or U428 (N_428,N_318,N_266);
nor U429 (N_429,N_353,N_389);
nor U430 (N_430,N_267,N_312);
or U431 (N_431,N_335,N_386);
nor U432 (N_432,N_295,N_377);
and U433 (N_433,N_316,N_238);
nand U434 (N_434,N_240,N_223);
nor U435 (N_435,N_370,N_323);
or U436 (N_436,N_352,N_345);
or U437 (N_437,N_210,N_313);
nand U438 (N_438,N_256,N_212);
and U439 (N_439,N_360,N_291);
and U440 (N_440,N_337,N_340);
nand U441 (N_441,N_262,N_336);
and U442 (N_442,N_399,N_362);
or U443 (N_443,N_317,N_254);
or U444 (N_444,N_310,N_384);
or U445 (N_445,N_242,N_279);
or U446 (N_446,N_260,N_306);
nand U447 (N_447,N_329,N_278);
nor U448 (N_448,N_251,N_393);
nand U449 (N_449,N_286,N_224);
and U450 (N_450,N_327,N_245);
nand U451 (N_451,N_265,N_358);
nor U452 (N_452,N_320,N_271);
or U453 (N_453,N_268,N_366);
nor U454 (N_454,N_390,N_275);
nor U455 (N_455,N_297,N_325);
and U456 (N_456,N_391,N_359);
nor U457 (N_457,N_304,N_388);
nor U458 (N_458,N_322,N_378);
nand U459 (N_459,N_250,N_303);
or U460 (N_460,N_209,N_300);
and U461 (N_461,N_218,N_356);
nand U462 (N_462,N_355,N_374);
nand U463 (N_463,N_376,N_350);
xnor U464 (N_464,N_228,N_369);
and U465 (N_465,N_347,N_239);
nor U466 (N_466,N_394,N_365);
or U467 (N_467,N_298,N_227);
nand U468 (N_468,N_342,N_287);
and U469 (N_469,N_321,N_249);
or U470 (N_470,N_274,N_207);
nor U471 (N_471,N_382,N_296);
nand U472 (N_472,N_305,N_283);
and U473 (N_473,N_392,N_289);
nand U474 (N_474,N_252,N_346);
nand U475 (N_475,N_277,N_284);
or U476 (N_476,N_248,N_354);
nand U477 (N_477,N_338,N_398);
nor U478 (N_478,N_231,N_201);
nor U479 (N_479,N_244,N_219);
and U480 (N_480,N_333,N_349);
nor U481 (N_481,N_301,N_253);
nand U482 (N_482,N_222,N_216);
and U483 (N_483,N_206,N_368);
nand U484 (N_484,N_334,N_319);
or U485 (N_485,N_307,N_281);
or U486 (N_486,N_282,N_230);
or U487 (N_487,N_259,N_357);
nand U488 (N_488,N_308,N_234);
nand U489 (N_489,N_373,N_264);
and U490 (N_490,N_203,N_348);
and U491 (N_491,N_361,N_217);
or U492 (N_492,N_380,N_341);
nor U493 (N_493,N_263,N_379);
nor U494 (N_494,N_221,N_205);
nand U495 (N_495,N_293,N_385);
or U496 (N_496,N_328,N_280);
nor U497 (N_497,N_344,N_372);
nor U498 (N_498,N_381,N_396);
or U499 (N_499,N_292,N_261);
or U500 (N_500,N_268,N_228);
and U501 (N_501,N_251,N_359);
or U502 (N_502,N_271,N_268);
and U503 (N_503,N_377,N_233);
and U504 (N_504,N_281,N_200);
or U505 (N_505,N_307,N_201);
or U506 (N_506,N_271,N_296);
nand U507 (N_507,N_342,N_312);
nor U508 (N_508,N_284,N_374);
nor U509 (N_509,N_223,N_269);
or U510 (N_510,N_243,N_296);
and U511 (N_511,N_216,N_261);
nand U512 (N_512,N_383,N_219);
nand U513 (N_513,N_340,N_208);
and U514 (N_514,N_398,N_221);
or U515 (N_515,N_353,N_378);
nand U516 (N_516,N_228,N_202);
xor U517 (N_517,N_303,N_389);
or U518 (N_518,N_393,N_390);
or U519 (N_519,N_386,N_237);
or U520 (N_520,N_231,N_271);
and U521 (N_521,N_276,N_379);
and U522 (N_522,N_246,N_205);
and U523 (N_523,N_330,N_392);
and U524 (N_524,N_281,N_399);
nand U525 (N_525,N_297,N_216);
nand U526 (N_526,N_382,N_357);
nor U527 (N_527,N_360,N_357);
nand U528 (N_528,N_386,N_204);
or U529 (N_529,N_325,N_358);
and U530 (N_530,N_373,N_271);
or U531 (N_531,N_386,N_242);
nor U532 (N_532,N_377,N_243);
and U533 (N_533,N_397,N_244);
nand U534 (N_534,N_217,N_257);
nand U535 (N_535,N_362,N_350);
nand U536 (N_536,N_209,N_390);
and U537 (N_537,N_203,N_334);
nor U538 (N_538,N_276,N_324);
or U539 (N_539,N_332,N_323);
or U540 (N_540,N_380,N_204);
and U541 (N_541,N_366,N_337);
nor U542 (N_542,N_316,N_212);
and U543 (N_543,N_365,N_371);
nor U544 (N_544,N_386,N_378);
or U545 (N_545,N_238,N_352);
nand U546 (N_546,N_257,N_205);
nand U547 (N_547,N_396,N_257);
or U548 (N_548,N_273,N_304);
or U549 (N_549,N_302,N_376);
and U550 (N_550,N_347,N_212);
and U551 (N_551,N_277,N_359);
or U552 (N_552,N_268,N_229);
and U553 (N_553,N_282,N_368);
nand U554 (N_554,N_219,N_374);
nand U555 (N_555,N_204,N_238);
and U556 (N_556,N_302,N_299);
or U557 (N_557,N_335,N_311);
or U558 (N_558,N_337,N_257);
nand U559 (N_559,N_347,N_209);
and U560 (N_560,N_216,N_334);
and U561 (N_561,N_371,N_385);
and U562 (N_562,N_357,N_234);
nor U563 (N_563,N_316,N_243);
and U564 (N_564,N_299,N_284);
nor U565 (N_565,N_209,N_228);
nor U566 (N_566,N_345,N_204);
or U567 (N_567,N_340,N_385);
nand U568 (N_568,N_213,N_232);
nand U569 (N_569,N_234,N_275);
or U570 (N_570,N_279,N_229);
and U571 (N_571,N_321,N_208);
and U572 (N_572,N_213,N_352);
or U573 (N_573,N_387,N_211);
nand U574 (N_574,N_218,N_241);
nor U575 (N_575,N_235,N_322);
nor U576 (N_576,N_354,N_361);
nand U577 (N_577,N_377,N_346);
and U578 (N_578,N_386,N_347);
nand U579 (N_579,N_266,N_297);
and U580 (N_580,N_348,N_301);
and U581 (N_581,N_395,N_280);
nand U582 (N_582,N_274,N_264);
nand U583 (N_583,N_241,N_352);
nand U584 (N_584,N_205,N_383);
nand U585 (N_585,N_321,N_295);
nand U586 (N_586,N_241,N_297);
and U587 (N_587,N_365,N_272);
and U588 (N_588,N_264,N_341);
and U589 (N_589,N_326,N_321);
or U590 (N_590,N_367,N_334);
and U591 (N_591,N_249,N_302);
or U592 (N_592,N_305,N_317);
and U593 (N_593,N_286,N_245);
or U594 (N_594,N_375,N_342);
nand U595 (N_595,N_246,N_222);
and U596 (N_596,N_376,N_217);
or U597 (N_597,N_377,N_315);
or U598 (N_598,N_218,N_261);
and U599 (N_599,N_248,N_257);
nor U600 (N_600,N_534,N_422);
nor U601 (N_601,N_495,N_549);
and U602 (N_602,N_492,N_577);
nand U603 (N_603,N_465,N_563);
xnor U604 (N_604,N_571,N_505);
nand U605 (N_605,N_565,N_559);
nand U606 (N_606,N_483,N_436);
and U607 (N_607,N_451,N_456);
nor U608 (N_608,N_567,N_543);
and U609 (N_609,N_455,N_583);
or U610 (N_610,N_546,N_588);
nor U611 (N_611,N_569,N_568);
and U612 (N_612,N_501,N_516);
and U613 (N_613,N_503,N_452);
nand U614 (N_614,N_586,N_410);
nand U615 (N_615,N_470,N_494);
or U616 (N_616,N_497,N_475);
nand U617 (N_617,N_551,N_426);
or U618 (N_618,N_482,N_599);
and U619 (N_619,N_485,N_498);
and U620 (N_620,N_581,N_467);
nor U621 (N_621,N_463,N_420);
or U622 (N_622,N_520,N_572);
and U623 (N_623,N_474,N_526);
and U624 (N_624,N_449,N_518);
nor U625 (N_625,N_421,N_461);
nor U626 (N_626,N_542,N_530);
nor U627 (N_627,N_537,N_595);
nand U628 (N_628,N_418,N_533);
and U629 (N_629,N_448,N_491);
and U630 (N_630,N_517,N_499);
xnor U631 (N_631,N_400,N_489);
nor U632 (N_632,N_472,N_545);
nand U633 (N_633,N_576,N_578);
or U634 (N_634,N_579,N_427);
and U635 (N_635,N_442,N_525);
nor U636 (N_636,N_538,N_444);
and U637 (N_637,N_473,N_447);
or U638 (N_638,N_566,N_423);
and U639 (N_639,N_478,N_540);
nor U640 (N_640,N_587,N_511);
nand U641 (N_641,N_573,N_419);
nand U642 (N_642,N_531,N_407);
nor U643 (N_643,N_584,N_412);
nand U644 (N_644,N_589,N_481);
nor U645 (N_645,N_469,N_594);
and U646 (N_646,N_443,N_405);
or U647 (N_647,N_408,N_413);
and U648 (N_648,N_561,N_560);
and U649 (N_649,N_502,N_440);
and U650 (N_650,N_552,N_479);
nor U651 (N_651,N_532,N_541);
nor U652 (N_652,N_570,N_425);
or U653 (N_653,N_460,N_555);
or U654 (N_654,N_429,N_593);
and U655 (N_655,N_580,N_445);
nand U656 (N_656,N_486,N_450);
and U657 (N_657,N_441,N_477);
and U658 (N_658,N_564,N_519);
nor U659 (N_659,N_496,N_500);
or U660 (N_660,N_428,N_487);
nand U661 (N_661,N_459,N_480);
nor U662 (N_662,N_454,N_508);
or U663 (N_663,N_527,N_597);
nor U664 (N_664,N_528,N_431);
nand U665 (N_665,N_513,N_522);
nor U666 (N_666,N_403,N_401);
xnor U667 (N_667,N_514,N_507);
and U668 (N_668,N_493,N_509);
nand U669 (N_669,N_510,N_464);
and U670 (N_670,N_548,N_590);
nor U671 (N_671,N_432,N_515);
nand U672 (N_672,N_506,N_575);
nor U673 (N_673,N_458,N_402);
nand U674 (N_674,N_466,N_434);
and U675 (N_675,N_462,N_471);
nand U676 (N_676,N_535,N_435);
and U677 (N_677,N_490,N_598);
or U678 (N_678,N_453,N_512);
nand U679 (N_679,N_437,N_484);
and U680 (N_680,N_457,N_592);
and U681 (N_681,N_424,N_562);
nor U682 (N_682,N_411,N_406);
nand U683 (N_683,N_438,N_416);
nor U684 (N_684,N_529,N_574);
or U685 (N_685,N_536,N_556);
and U686 (N_686,N_585,N_468);
nor U687 (N_687,N_523,N_539);
or U688 (N_688,N_415,N_544);
nor U689 (N_689,N_404,N_591);
nand U690 (N_690,N_553,N_414);
or U691 (N_691,N_596,N_521);
or U692 (N_692,N_547,N_524);
or U693 (N_693,N_557,N_439);
nand U694 (N_694,N_558,N_409);
nor U695 (N_695,N_433,N_446);
nand U696 (N_696,N_476,N_417);
nand U697 (N_697,N_582,N_488);
and U698 (N_698,N_504,N_554);
nor U699 (N_699,N_430,N_550);
nand U700 (N_700,N_507,N_479);
and U701 (N_701,N_466,N_531);
nand U702 (N_702,N_548,N_467);
or U703 (N_703,N_492,N_522);
and U704 (N_704,N_492,N_506);
nor U705 (N_705,N_575,N_489);
nand U706 (N_706,N_592,N_569);
nand U707 (N_707,N_559,N_521);
or U708 (N_708,N_520,N_432);
nand U709 (N_709,N_594,N_457);
or U710 (N_710,N_405,N_433);
and U711 (N_711,N_534,N_526);
and U712 (N_712,N_580,N_577);
or U713 (N_713,N_475,N_551);
nor U714 (N_714,N_419,N_590);
and U715 (N_715,N_526,N_561);
and U716 (N_716,N_493,N_523);
nand U717 (N_717,N_559,N_415);
nor U718 (N_718,N_591,N_482);
and U719 (N_719,N_448,N_519);
nand U720 (N_720,N_426,N_418);
nor U721 (N_721,N_553,N_454);
and U722 (N_722,N_467,N_439);
nand U723 (N_723,N_412,N_488);
nand U724 (N_724,N_580,N_456);
nand U725 (N_725,N_460,N_445);
or U726 (N_726,N_443,N_552);
nand U727 (N_727,N_496,N_433);
or U728 (N_728,N_524,N_582);
and U729 (N_729,N_593,N_507);
and U730 (N_730,N_436,N_559);
and U731 (N_731,N_426,N_543);
nor U732 (N_732,N_425,N_407);
nand U733 (N_733,N_485,N_449);
nor U734 (N_734,N_534,N_543);
nand U735 (N_735,N_454,N_564);
nand U736 (N_736,N_597,N_491);
or U737 (N_737,N_585,N_587);
nand U738 (N_738,N_488,N_421);
or U739 (N_739,N_531,N_593);
and U740 (N_740,N_539,N_405);
nor U741 (N_741,N_476,N_535);
nor U742 (N_742,N_429,N_431);
or U743 (N_743,N_539,N_506);
or U744 (N_744,N_548,N_589);
nand U745 (N_745,N_493,N_561);
or U746 (N_746,N_505,N_445);
nand U747 (N_747,N_512,N_475);
or U748 (N_748,N_531,N_504);
xor U749 (N_749,N_598,N_526);
nor U750 (N_750,N_599,N_566);
nand U751 (N_751,N_437,N_529);
nand U752 (N_752,N_543,N_472);
nor U753 (N_753,N_503,N_565);
nand U754 (N_754,N_482,N_443);
nand U755 (N_755,N_551,N_467);
nor U756 (N_756,N_527,N_557);
or U757 (N_757,N_477,N_420);
nor U758 (N_758,N_577,N_588);
and U759 (N_759,N_495,N_410);
nand U760 (N_760,N_445,N_523);
nand U761 (N_761,N_586,N_594);
xnor U762 (N_762,N_421,N_486);
and U763 (N_763,N_554,N_404);
nand U764 (N_764,N_505,N_514);
nand U765 (N_765,N_519,N_525);
nor U766 (N_766,N_564,N_511);
and U767 (N_767,N_526,N_559);
nand U768 (N_768,N_430,N_537);
or U769 (N_769,N_547,N_500);
nor U770 (N_770,N_488,N_526);
nand U771 (N_771,N_591,N_442);
nand U772 (N_772,N_535,N_579);
and U773 (N_773,N_428,N_494);
or U774 (N_774,N_441,N_458);
and U775 (N_775,N_435,N_463);
or U776 (N_776,N_474,N_495);
or U777 (N_777,N_416,N_454);
or U778 (N_778,N_543,N_514);
and U779 (N_779,N_412,N_453);
or U780 (N_780,N_478,N_457);
nand U781 (N_781,N_408,N_425);
and U782 (N_782,N_517,N_401);
and U783 (N_783,N_522,N_443);
xor U784 (N_784,N_508,N_479);
nor U785 (N_785,N_464,N_566);
nor U786 (N_786,N_554,N_533);
nand U787 (N_787,N_572,N_574);
nand U788 (N_788,N_416,N_588);
nor U789 (N_789,N_520,N_545);
nand U790 (N_790,N_416,N_597);
nor U791 (N_791,N_475,N_526);
and U792 (N_792,N_435,N_447);
nand U793 (N_793,N_455,N_544);
nand U794 (N_794,N_425,N_424);
or U795 (N_795,N_504,N_469);
or U796 (N_796,N_569,N_562);
or U797 (N_797,N_441,N_502);
or U798 (N_798,N_408,N_561);
and U799 (N_799,N_436,N_576);
nor U800 (N_800,N_688,N_746);
and U801 (N_801,N_669,N_797);
nor U802 (N_802,N_676,N_614);
nor U803 (N_803,N_613,N_640);
nand U804 (N_804,N_634,N_728);
and U805 (N_805,N_641,N_606);
or U806 (N_806,N_712,N_715);
or U807 (N_807,N_758,N_781);
nor U808 (N_808,N_629,N_760);
nand U809 (N_809,N_770,N_733);
and U810 (N_810,N_796,N_779);
and U811 (N_811,N_674,N_735);
nand U812 (N_812,N_671,N_668);
nand U813 (N_813,N_780,N_659);
nor U814 (N_814,N_710,N_711);
and U815 (N_815,N_620,N_705);
or U816 (N_816,N_719,N_682);
nor U817 (N_817,N_689,N_684);
or U818 (N_818,N_720,N_789);
and U819 (N_819,N_722,N_605);
nor U820 (N_820,N_698,N_651);
nand U821 (N_821,N_607,N_601);
xor U822 (N_822,N_612,N_602);
or U823 (N_823,N_649,N_673);
or U824 (N_824,N_622,N_691);
nand U825 (N_825,N_771,N_670);
and U826 (N_826,N_677,N_600);
nor U827 (N_827,N_617,N_791);
and U828 (N_828,N_655,N_616);
or U829 (N_829,N_724,N_794);
nor U830 (N_830,N_665,N_738);
nand U831 (N_831,N_757,N_666);
and U832 (N_832,N_660,N_654);
nor U833 (N_833,N_662,N_609);
or U834 (N_834,N_775,N_639);
or U835 (N_835,N_747,N_690);
nor U836 (N_836,N_793,N_798);
or U837 (N_837,N_648,N_740);
nor U838 (N_838,N_663,N_604);
and U839 (N_839,N_736,N_784);
and U840 (N_840,N_632,N_743);
nand U841 (N_841,N_618,N_672);
or U842 (N_842,N_696,N_795);
nand U843 (N_843,N_638,N_699);
or U844 (N_844,N_658,N_764);
and U845 (N_845,N_717,N_767);
or U846 (N_846,N_765,N_748);
or U847 (N_847,N_643,N_610);
or U848 (N_848,N_652,N_753);
nor U849 (N_849,N_644,N_692);
nand U850 (N_850,N_704,N_636);
nor U851 (N_851,N_630,N_786);
or U852 (N_852,N_637,N_642);
nor U853 (N_853,N_777,N_678);
nand U854 (N_854,N_608,N_754);
nand U855 (N_855,N_667,N_725);
and U856 (N_856,N_683,N_737);
or U857 (N_857,N_730,N_721);
nor U858 (N_858,N_751,N_729);
nor U859 (N_859,N_621,N_783);
and U860 (N_860,N_706,N_656);
nor U861 (N_861,N_633,N_686);
nand U862 (N_862,N_619,N_664);
nor U863 (N_863,N_734,N_774);
xor U864 (N_864,N_693,N_661);
or U865 (N_865,N_776,N_708);
nand U866 (N_866,N_650,N_713);
nand U867 (N_867,N_623,N_718);
and U868 (N_868,N_726,N_731);
nor U869 (N_869,N_657,N_752);
nand U870 (N_870,N_785,N_756);
nand U871 (N_871,N_768,N_700);
nor U872 (N_872,N_714,N_709);
nor U873 (N_873,N_697,N_799);
nand U874 (N_874,N_707,N_628);
or U875 (N_875,N_626,N_723);
or U876 (N_876,N_761,N_687);
and U877 (N_877,N_759,N_755);
or U878 (N_878,N_675,N_741);
and U879 (N_879,N_742,N_744);
and U880 (N_880,N_635,N_762);
and U881 (N_881,N_716,N_750);
nand U882 (N_882,N_763,N_782);
nand U883 (N_883,N_611,N_645);
and U884 (N_884,N_615,N_778);
or U885 (N_885,N_745,N_772);
nor U886 (N_886,N_681,N_624);
and U887 (N_887,N_701,N_680);
nor U888 (N_888,N_732,N_694);
or U889 (N_889,N_727,N_627);
or U890 (N_890,N_749,N_647);
and U891 (N_891,N_769,N_679);
or U892 (N_892,N_625,N_685);
nand U893 (N_893,N_703,N_773);
or U894 (N_894,N_646,N_702);
nor U895 (N_895,N_787,N_603);
nor U896 (N_896,N_792,N_766);
or U897 (N_897,N_739,N_788);
or U898 (N_898,N_631,N_790);
and U899 (N_899,N_653,N_695);
nor U900 (N_900,N_703,N_781);
and U901 (N_901,N_672,N_736);
and U902 (N_902,N_742,N_699);
or U903 (N_903,N_601,N_672);
nand U904 (N_904,N_637,N_792);
nor U905 (N_905,N_654,N_692);
nor U906 (N_906,N_696,N_651);
and U907 (N_907,N_612,N_639);
and U908 (N_908,N_733,N_669);
and U909 (N_909,N_605,N_735);
and U910 (N_910,N_710,N_725);
xor U911 (N_911,N_765,N_655);
nand U912 (N_912,N_746,N_690);
nand U913 (N_913,N_702,N_758);
nand U914 (N_914,N_605,N_636);
nand U915 (N_915,N_600,N_653);
or U916 (N_916,N_653,N_767);
nor U917 (N_917,N_771,N_745);
and U918 (N_918,N_642,N_658);
or U919 (N_919,N_767,N_722);
nor U920 (N_920,N_661,N_680);
or U921 (N_921,N_717,N_689);
or U922 (N_922,N_672,N_746);
or U923 (N_923,N_682,N_779);
and U924 (N_924,N_776,N_672);
and U925 (N_925,N_682,N_600);
nand U926 (N_926,N_646,N_661);
and U927 (N_927,N_744,N_759);
and U928 (N_928,N_701,N_681);
nand U929 (N_929,N_628,N_682);
nor U930 (N_930,N_724,N_690);
nand U931 (N_931,N_609,N_782);
nand U932 (N_932,N_758,N_632);
nor U933 (N_933,N_712,N_764);
and U934 (N_934,N_728,N_759);
nor U935 (N_935,N_775,N_787);
nor U936 (N_936,N_689,N_754);
nor U937 (N_937,N_776,N_636);
nor U938 (N_938,N_642,N_755);
or U939 (N_939,N_728,N_638);
and U940 (N_940,N_782,N_648);
or U941 (N_941,N_715,N_627);
and U942 (N_942,N_739,N_726);
nand U943 (N_943,N_794,N_660);
nand U944 (N_944,N_762,N_675);
or U945 (N_945,N_690,N_756);
or U946 (N_946,N_636,N_653);
nand U947 (N_947,N_614,N_697);
and U948 (N_948,N_741,N_732);
nand U949 (N_949,N_605,N_770);
and U950 (N_950,N_626,N_695);
nand U951 (N_951,N_779,N_775);
nor U952 (N_952,N_667,N_605);
or U953 (N_953,N_761,N_657);
and U954 (N_954,N_711,N_669);
or U955 (N_955,N_791,N_719);
and U956 (N_956,N_676,N_606);
or U957 (N_957,N_780,N_623);
and U958 (N_958,N_657,N_616);
nor U959 (N_959,N_623,N_617);
or U960 (N_960,N_784,N_664);
nor U961 (N_961,N_637,N_775);
or U962 (N_962,N_799,N_745);
and U963 (N_963,N_758,N_616);
nand U964 (N_964,N_623,N_767);
nand U965 (N_965,N_741,N_740);
and U966 (N_966,N_747,N_609);
nor U967 (N_967,N_616,N_727);
nor U968 (N_968,N_609,N_768);
nor U969 (N_969,N_617,N_645);
nor U970 (N_970,N_735,N_658);
and U971 (N_971,N_693,N_773);
nor U972 (N_972,N_758,N_645);
or U973 (N_973,N_679,N_722);
and U974 (N_974,N_665,N_763);
and U975 (N_975,N_742,N_639);
nor U976 (N_976,N_792,N_746);
or U977 (N_977,N_702,N_622);
nor U978 (N_978,N_743,N_681);
nand U979 (N_979,N_722,N_665);
or U980 (N_980,N_603,N_713);
and U981 (N_981,N_654,N_621);
nor U982 (N_982,N_613,N_717);
or U983 (N_983,N_790,N_687);
and U984 (N_984,N_751,N_695);
or U985 (N_985,N_747,N_684);
and U986 (N_986,N_720,N_621);
and U987 (N_987,N_776,N_790);
or U988 (N_988,N_655,N_719);
or U989 (N_989,N_784,N_601);
or U990 (N_990,N_627,N_673);
nor U991 (N_991,N_729,N_645);
nand U992 (N_992,N_659,N_768);
nor U993 (N_993,N_663,N_632);
and U994 (N_994,N_791,N_717);
and U995 (N_995,N_753,N_701);
nor U996 (N_996,N_615,N_758);
and U997 (N_997,N_787,N_612);
and U998 (N_998,N_611,N_617);
nand U999 (N_999,N_721,N_677);
nor U1000 (N_1000,N_915,N_805);
nand U1001 (N_1001,N_816,N_935);
and U1002 (N_1002,N_891,N_876);
nor U1003 (N_1003,N_908,N_812);
and U1004 (N_1004,N_830,N_834);
or U1005 (N_1005,N_965,N_859);
xnor U1006 (N_1006,N_942,N_836);
and U1007 (N_1007,N_845,N_977);
or U1008 (N_1008,N_870,N_962);
nor U1009 (N_1009,N_903,N_994);
and U1010 (N_1010,N_945,N_852);
or U1011 (N_1011,N_877,N_824);
nor U1012 (N_1012,N_932,N_807);
or U1013 (N_1013,N_989,N_963);
nand U1014 (N_1014,N_966,N_810);
or U1015 (N_1015,N_858,N_895);
nand U1016 (N_1016,N_857,N_811);
or U1017 (N_1017,N_803,N_919);
or U1018 (N_1018,N_955,N_889);
or U1019 (N_1019,N_841,N_862);
and U1020 (N_1020,N_801,N_918);
or U1021 (N_1021,N_867,N_960);
nor U1022 (N_1022,N_986,N_866);
nor U1023 (N_1023,N_818,N_890);
and U1024 (N_1024,N_980,N_847);
or U1025 (N_1025,N_938,N_827);
and U1026 (N_1026,N_846,N_887);
nand U1027 (N_1027,N_865,N_843);
nor U1028 (N_1028,N_815,N_911);
nand U1029 (N_1029,N_853,N_927);
nor U1030 (N_1030,N_828,N_849);
nor U1031 (N_1031,N_995,N_900);
nor U1032 (N_1032,N_928,N_924);
and U1033 (N_1033,N_978,N_822);
or U1034 (N_1034,N_892,N_825);
nor U1035 (N_1035,N_952,N_861);
or U1036 (N_1036,N_976,N_893);
and U1037 (N_1037,N_930,N_957);
nand U1038 (N_1038,N_884,N_883);
nand U1039 (N_1039,N_850,N_913);
and U1040 (N_1040,N_979,N_988);
and U1041 (N_1041,N_910,N_808);
nand U1042 (N_1042,N_868,N_814);
and U1043 (N_1043,N_837,N_821);
nand U1044 (N_1044,N_982,N_956);
or U1045 (N_1045,N_964,N_842);
and U1046 (N_1046,N_992,N_909);
xor U1047 (N_1047,N_885,N_813);
nand U1048 (N_1048,N_937,N_898);
and U1049 (N_1049,N_855,N_971);
nand U1050 (N_1050,N_806,N_901);
and U1051 (N_1051,N_925,N_838);
or U1052 (N_1052,N_894,N_974);
nand U1053 (N_1053,N_904,N_993);
nor U1054 (N_1054,N_880,N_922);
or U1055 (N_1055,N_871,N_998);
and U1056 (N_1056,N_888,N_947);
nand U1057 (N_1057,N_882,N_899);
nand U1058 (N_1058,N_829,N_864);
or U1059 (N_1059,N_987,N_886);
or U1060 (N_1060,N_860,N_800);
nand U1061 (N_1061,N_950,N_851);
and U1062 (N_1062,N_940,N_840);
nand U1063 (N_1063,N_905,N_968);
nand U1064 (N_1064,N_999,N_873);
nand U1065 (N_1065,N_949,N_934);
and U1066 (N_1066,N_975,N_972);
and U1067 (N_1067,N_959,N_951);
nand U1068 (N_1068,N_958,N_809);
or U1069 (N_1069,N_984,N_819);
or U1070 (N_1070,N_869,N_991);
and U1071 (N_1071,N_990,N_946);
nor U1072 (N_1072,N_826,N_969);
nor U1073 (N_1073,N_933,N_902);
and U1074 (N_1074,N_896,N_961);
nor U1075 (N_1075,N_844,N_944);
or U1076 (N_1076,N_879,N_878);
or U1077 (N_1077,N_856,N_916);
and U1078 (N_1078,N_875,N_920);
and U1079 (N_1079,N_917,N_897);
or U1080 (N_1080,N_823,N_907);
xnor U1081 (N_1081,N_874,N_848);
or U1082 (N_1082,N_929,N_996);
or U1083 (N_1083,N_832,N_835);
nor U1084 (N_1084,N_931,N_863);
or U1085 (N_1085,N_981,N_833);
nand U1086 (N_1086,N_802,N_926);
and U1087 (N_1087,N_872,N_854);
nand U1088 (N_1088,N_906,N_881);
and U1089 (N_1089,N_954,N_912);
nor U1090 (N_1090,N_985,N_970);
nand U1091 (N_1091,N_923,N_953);
or U1092 (N_1092,N_941,N_921);
or U1093 (N_1093,N_804,N_997);
and U1094 (N_1094,N_948,N_983);
nand U1095 (N_1095,N_831,N_820);
or U1096 (N_1096,N_817,N_939);
nand U1097 (N_1097,N_839,N_943);
nor U1098 (N_1098,N_967,N_914);
xnor U1099 (N_1099,N_973,N_936);
and U1100 (N_1100,N_873,N_800);
and U1101 (N_1101,N_871,N_978);
or U1102 (N_1102,N_934,N_898);
nand U1103 (N_1103,N_995,N_872);
nor U1104 (N_1104,N_990,N_934);
or U1105 (N_1105,N_890,N_919);
nor U1106 (N_1106,N_871,N_869);
nor U1107 (N_1107,N_940,N_979);
nor U1108 (N_1108,N_928,N_882);
and U1109 (N_1109,N_959,N_927);
or U1110 (N_1110,N_826,N_817);
nor U1111 (N_1111,N_814,N_960);
nand U1112 (N_1112,N_978,N_894);
nand U1113 (N_1113,N_836,N_809);
nand U1114 (N_1114,N_943,N_846);
or U1115 (N_1115,N_804,N_890);
or U1116 (N_1116,N_944,N_924);
nor U1117 (N_1117,N_835,N_951);
or U1118 (N_1118,N_939,N_913);
nand U1119 (N_1119,N_841,N_973);
or U1120 (N_1120,N_985,N_811);
and U1121 (N_1121,N_994,N_947);
and U1122 (N_1122,N_815,N_959);
nand U1123 (N_1123,N_910,N_945);
nor U1124 (N_1124,N_909,N_856);
and U1125 (N_1125,N_821,N_975);
nand U1126 (N_1126,N_827,N_824);
nor U1127 (N_1127,N_909,N_918);
nor U1128 (N_1128,N_914,N_989);
nand U1129 (N_1129,N_932,N_851);
nand U1130 (N_1130,N_810,N_957);
nor U1131 (N_1131,N_984,N_998);
and U1132 (N_1132,N_838,N_938);
nand U1133 (N_1133,N_939,N_955);
or U1134 (N_1134,N_854,N_877);
nor U1135 (N_1135,N_830,N_803);
nand U1136 (N_1136,N_878,N_980);
or U1137 (N_1137,N_968,N_939);
nand U1138 (N_1138,N_853,N_849);
and U1139 (N_1139,N_983,N_809);
nand U1140 (N_1140,N_954,N_995);
or U1141 (N_1141,N_930,N_852);
or U1142 (N_1142,N_990,N_811);
and U1143 (N_1143,N_826,N_849);
nor U1144 (N_1144,N_953,N_848);
nand U1145 (N_1145,N_842,N_894);
and U1146 (N_1146,N_860,N_937);
nand U1147 (N_1147,N_918,N_806);
nand U1148 (N_1148,N_963,N_939);
or U1149 (N_1149,N_857,N_997);
nor U1150 (N_1150,N_823,N_893);
nor U1151 (N_1151,N_900,N_819);
or U1152 (N_1152,N_969,N_967);
nand U1153 (N_1153,N_994,N_992);
nor U1154 (N_1154,N_837,N_950);
and U1155 (N_1155,N_992,N_947);
nor U1156 (N_1156,N_982,N_868);
nor U1157 (N_1157,N_988,N_856);
nand U1158 (N_1158,N_858,N_861);
nand U1159 (N_1159,N_897,N_971);
or U1160 (N_1160,N_936,N_934);
and U1161 (N_1161,N_849,N_971);
nand U1162 (N_1162,N_827,N_864);
xnor U1163 (N_1163,N_900,N_952);
nand U1164 (N_1164,N_870,N_996);
nor U1165 (N_1165,N_849,N_972);
and U1166 (N_1166,N_956,N_990);
or U1167 (N_1167,N_809,N_822);
nand U1168 (N_1168,N_803,N_903);
and U1169 (N_1169,N_826,N_925);
and U1170 (N_1170,N_845,N_816);
or U1171 (N_1171,N_950,N_880);
and U1172 (N_1172,N_842,N_885);
or U1173 (N_1173,N_969,N_909);
and U1174 (N_1174,N_820,N_813);
and U1175 (N_1175,N_917,N_848);
or U1176 (N_1176,N_872,N_886);
nor U1177 (N_1177,N_916,N_950);
nand U1178 (N_1178,N_900,N_890);
or U1179 (N_1179,N_874,N_995);
nand U1180 (N_1180,N_969,N_813);
nor U1181 (N_1181,N_806,N_973);
nor U1182 (N_1182,N_897,N_802);
or U1183 (N_1183,N_936,N_940);
nor U1184 (N_1184,N_897,N_809);
and U1185 (N_1185,N_943,N_815);
nand U1186 (N_1186,N_933,N_931);
nor U1187 (N_1187,N_873,N_939);
nor U1188 (N_1188,N_860,N_850);
nand U1189 (N_1189,N_929,N_900);
or U1190 (N_1190,N_988,N_941);
or U1191 (N_1191,N_848,N_948);
and U1192 (N_1192,N_943,N_909);
and U1193 (N_1193,N_910,N_883);
nor U1194 (N_1194,N_880,N_991);
nor U1195 (N_1195,N_902,N_942);
xor U1196 (N_1196,N_981,N_964);
and U1197 (N_1197,N_804,N_904);
nor U1198 (N_1198,N_955,N_972);
nand U1199 (N_1199,N_872,N_975);
nor U1200 (N_1200,N_1156,N_1103);
and U1201 (N_1201,N_1013,N_1018);
nor U1202 (N_1202,N_1023,N_1074);
nand U1203 (N_1203,N_1169,N_1077);
nor U1204 (N_1204,N_1067,N_1057);
nand U1205 (N_1205,N_1170,N_1040);
and U1206 (N_1206,N_1028,N_1066);
nor U1207 (N_1207,N_1145,N_1106);
nor U1208 (N_1208,N_1070,N_1085);
nor U1209 (N_1209,N_1093,N_1186);
and U1210 (N_1210,N_1008,N_1026);
nor U1211 (N_1211,N_1150,N_1165);
nand U1212 (N_1212,N_1116,N_1138);
nor U1213 (N_1213,N_1081,N_1166);
nor U1214 (N_1214,N_1094,N_1131);
and U1215 (N_1215,N_1000,N_1174);
nand U1216 (N_1216,N_1126,N_1161);
or U1217 (N_1217,N_1083,N_1104);
nor U1218 (N_1218,N_1095,N_1089);
or U1219 (N_1219,N_1086,N_1019);
nor U1220 (N_1220,N_1115,N_1012);
or U1221 (N_1221,N_1049,N_1198);
or U1222 (N_1222,N_1167,N_1146);
and U1223 (N_1223,N_1180,N_1031);
and U1224 (N_1224,N_1082,N_1188);
nand U1225 (N_1225,N_1105,N_1114);
and U1226 (N_1226,N_1118,N_1035);
or U1227 (N_1227,N_1171,N_1024);
and U1228 (N_1228,N_1032,N_1047);
nand U1229 (N_1229,N_1060,N_1042);
and U1230 (N_1230,N_1014,N_1176);
nor U1231 (N_1231,N_1058,N_1157);
nor U1232 (N_1232,N_1109,N_1052);
nor U1233 (N_1233,N_1092,N_1133);
or U1234 (N_1234,N_1111,N_1005);
and U1235 (N_1235,N_1080,N_1182);
and U1236 (N_1236,N_1117,N_1079);
and U1237 (N_1237,N_1053,N_1159);
nor U1238 (N_1238,N_1048,N_1020);
nor U1239 (N_1239,N_1078,N_1168);
or U1240 (N_1240,N_1143,N_1129);
nand U1241 (N_1241,N_1055,N_1050);
nand U1242 (N_1242,N_1073,N_1144);
nand U1243 (N_1243,N_1072,N_1027);
nor U1244 (N_1244,N_1181,N_1041);
and U1245 (N_1245,N_1099,N_1172);
and U1246 (N_1246,N_1090,N_1160);
and U1247 (N_1247,N_1148,N_1179);
or U1248 (N_1248,N_1110,N_1021);
nand U1249 (N_1249,N_1107,N_1075);
nor U1250 (N_1250,N_1100,N_1098);
or U1251 (N_1251,N_1065,N_1178);
nor U1252 (N_1252,N_1033,N_1022);
nand U1253 (N_1253,N_1154,N_1124);
nand U1254 (N_1254,N_1096,N_1007);
and U1255 (N_1255,N_1162,N_1069);
nor U1256 (N_1256,N_1010,N_1113);
nor U1257 (N_1257,N_1149,N_1009);
nand U1258 (N_1258,N_1061,N_1068);
and U1259 (N_1259,N_1137,N_1046);
or U1260 (N_1260,N_1054,N_1043);
nand U1261 (N_1261,N_1038,N_1119);
nand U1262 (N_1262,N_1130,N_1199);
and U1263 (N_1263,N_1025,N_1128);
and U1264 (N_1264,N_1158,N_1136);
and U1265 (N_1265,N_1039,N_1191);
nor U1266 (N_1266,N_1123,N_1011);
and U1267 (N_1267,N_1192,N_1037);
nand U1268 (N_1268,N_1036,N_1101);
and U1269 (N_1269,N_1064,N_1132);
and U1270 (N_1270,N_1140,N_1108);
nand U1271 (N_1271,N_1134,N_1189);
nand U1272 (N_1272,N_1051,N_1177);
or U1273 (N_1273,N_1001,N_1063);
or U1274 (N_1274,N_1183,N_1127);
nor U1275 (N_1275,N_1121,N_1002);
and U1276 (N_1276,N_1006,N_1097);
xor U1277 (N_1277,N_1196,N_1084);
or U1278 (N_1278,N_1190,N_1112);
or U1279 (N_1279,N_1059,N_1135);
or U1280 (N_1280,N_1015,N_1102);
or U1281 (N_1281,N_1045,N_1152);
nor U1282 (N_1282,N_1184,N_1029);
and U1283 (N_1283,N_1016,N_1030);
nand U1284 (N_1284,N_1197,N_1122);
and U1285 (N_1285,N_1017,N_1004);
nand U1286 (N_1286,N_1034,N_1044);
or U1287 (N_1287,N_1163,N_1125);
and U1288 (N_1288,N_1155,N_1062);
nor U1289 (N_1289,N_1147,N_1195);
or U1290 (N_1290,N_1139,N_1056);
or U1291 (N_1291,N_1175,N_1185);
nor U1292 (N_1292,N_1071,N_1164);
nor U1293 (N_1293,N_1142,N_1088);
or U1294 (N_1294,N_1194,N_1120);
nand U1295 (N_1295,N_1076,N_1187);
or U1296 (N_1296,N_1003,N_1193);
nand U1297 (N_1297,N_1151,N_1153);
nor U1298 (N_1298,N_1173,N_1087);
nor U1299 (N_1299,N_1141,N_1091);
nor U1300 (N_1300,N_1093,N_1115);
and U1301 (N_1301,N_1039,N_1171);
and U1302 (N_1302,N_1031,N_1084);
or U1303 (N_1303,N_1186,N_1171);
and U1304 (N_1304,N_1012,N_1022);
nand U1305 (N_1305,N_1052,N_1144);
and U1306 (N_1306,N_1073,N_1095);
nand U1307 (N_1307,N_1073,N_1167);
or U1308 (N_1308,N_1146,N_1030);
nor U1309 (N_1309,N_1170,N_1101);
and U1310 (N_1310,N_1095,N_1087);
or U1311 (N_1311,N_1128,N_1125);
and U1312 (N_1312,N_1041,N_1110);
nand U1313 (N_1313,N_1107,N_1071);
or U1314 (N_1314,N_1100,N_1164);
nor U1315 (N_1315,N_1062,N_1197);
and U1316 (N_1316,N_1020,N_1115);
and U1317 (N_1317,N_1157,N_1197);
or U1318 (N_1318,N_1126,N_1113);
nor U1319 (N_1319,N_1124,N_1079);
nor U1320 (N_1320,N_1175,N_1075);
or U1321 (N_1321,N_1192,N_1117);
or U1322 (N_1322,N_1015,N_1156);
and U1323 (N_1323,N_1052,N_1119);
or U1324 (N_1324,N_1128,N_1113);
or U1325 (N_1325,N_1093,N_1075);
nand U1326 (N_1326,N_1085,N_1186);
nand U1327 (N_1327,N_1166,N_1051);
or U1328 (N_1328,N_1107,N_1035);
or U1329 (N_1329,N_1100,N_1196);
nor U1330 (N_1330,N_1158,N_1073);
and U1331 (N_1331,N_1155,N_1042);
or U1332 (N_1332,N_1110,N_1036);
or U1333 (N_1333,N_1140,N_1080);
nor U1334 (N_1334,N_1136,N_1163);
nand U1335 (N_1335,N_1023,N_1091);
and U1336 (N_1336,N_1189,N_1198);
nor U1337 (N_1337,N_1152,N_1083);
and U1338 (N_1338,N_1137,N_1092);
nand U1339 (N_1339,N_1098,N_1090);
nand U1340 (N_1340,N_1199,N_1192);
nand U1341 (N_1341,N_1059,N_1142);
or U1342 (N_1342,N_1024,N_1005);
or U1343 (N_1343,N_1047,N_1003);
nor U1344 (N_1344,N_1065,N_1004);
or U1345 (N_1345,N_1146,N_1076);
nand U1346 (N_1346,N_1120,N_1190);
or U1347 (N_1347,N_1101,N_1116);
nor U1348 (N_1348,N_1129,N_1131);
and U1349 (N_1349,N_1111,N_1045);
or U1350 (N_1350,N_1064,N_1180);
and U1351 (N_1351,N_1057,N_1035);
and U1352 (N_1352,N_1176,N_1115);
or U1353 (N_1353,N_1130,N_1029);
nand U1354 (N_1354,N_1016,N_1011);
nand U1355 (N_1355,N_1177,N_1161);
nand U1356 (N_1356,N_1039,N_1079);
and U1357 (N_1357,N_1005,N_1000);
and U1358 (N_1358,N_1081,N_1087);
xnor U1359 (N_1359,N_1118,N_1030);
xnor U1360 (N_1360,N_1167,N_1039);
or U1361 (N_1361,N_1060,N_1162);
nor U1362 (N_1362,N_1151,N_1191);
or U1363 (N_1363,N_1009,N_1045);
or U1364 (N_1364,N_1146,N_1072);
nor U1365 (N_1365,N_1179,N_1067);
nand U1366 (N_1366,N_1042,N_1039);
nor U1367 (N_1367,N_1033,N_1094);
nand U1368 (N_1368,N_1033,N_1137);
and U1369 (N_1369,N_1021,N_1142);
or U1370 (N_1370,N_1187,N_1097);
nor U1371 (N_1371,N_1149,N_1038);
nor U1372 (N_1372,N_1025,N_1181);
nand U1373 (N_1373,N_1171,N_1049);
or U1374 (N_1374,N_1124,N_1131);
or U1375 (N_1375,N_1076,N_1047);
or U1376 (N_1376,N_1057,N_1165);
nor U1377 (N_1377,N_1095,N_1065);
or U1378 (N_1378,N_1033,N_1070);
or U1379 (N_1379,N_1069,N_1068);
and U1380 (N_1380,N_1117,N_1162);
or U1381 (N_1381,N_1136,N_1186);
nor U1382 (N_1382,N_1020,N_1141);
and U1383 (N_1383,N_1094,N_1008);
xor U1384 (N_1384,N_1080,N_1033);
nor U1385 (N_1385,N_1124,N_1031);
or U1386 (N_1386,N_1050,N_1181);
xor U1387 (N_1387,N_1088,N_1023);
and U1388 (N_1388,N_1111,N_1164);
nand U1389 (N_1389,N_1180,N_1124);
or U1390 (N_1390,N_1075,N_1038);
or U1391 (N_1391,N_1126,N_1015);
or U1392 (N_1392,N_1125,N_1157);
and U1393 (N_1393,N_1153,N_1100);
nand U1394 (N_1394,N_1099,N_1076);
or U1395 (N_1395,N_1173,N_1159);
nor U1396 (N_1396,N_1008,N_1088);
nor U1397 (N_1397,N_1167,N_1134);
nor U1398 (N_1398,N_1130,N_1109);
and U1399 (N_1399,N_1092,N_1100);
nand U1400 (N_1400,N_1220,N_1279);
nand U1401 (N_1401,N_1337,N_1222);
or U1402 (N_1402,N_1308,N_1287);
nor U1403 (N_1403,N_1320,N_1376);
or U1404 (N_1404,N_1254,N_1204);
nand U1405 (N_1405,N_1206,N_1328);
nand U1406 (N_1406,N_1330,N_1208);
and U1407 (N_1407,N_1327,N_1353);
or U1408 (N_1408,N_1202,N_1250);
and U1409 (N_1409,N_1262,N_1394);
and U1410 (N_1410,N_1349,N_1372);
nand U1411 (N_1411,N_1243,N_1303);
or U1412 (N_1412,N_1340,N_1368);
and U1413 (N_1413,N_1313,N_1384);
or U1414 (N_1414,N_1241,N_1276);
nor U1415 (N_1415,N_1295,N_1288);
nand U1416 (N_1416,N_1234,N_1316);
nand U1417 (N_1417,N_1351,N_1341);
nand U1418 (N_1418,N_1321,N_1214);
or U1419 (N_1419,N_1378,N_1331);
nand U1420 (N_1420,N_1293,N_1240);
nor U1421 (N_1421,N_1246,N_1280);
nor U1422 (N_1422,N_1348,N_1286);
or U1423 (N_1423,N_1312,N_1231);
nor U1424 (N_1424,N_1297,N_1257);
nor U1425 (N_1425,N_1223,N_1289);
nor U1426 (N_1426,N_1264,N_1339);
or U1427 (N_1427,N_1318,N_1356);
nand U1428 (N_1428,N_1375,N_1290);
or U1429 (N_1429,N_1385,N_1211);
and U1430 (N_1430,N_1212,N_1294);
nand U1431 (N_1431,N_1338,N_1256);
or U1432 (N_1432,N_1233,N_1228);
and U1433 (N_1433,N_1267,N_1363);
or U1434 (N_1434,N_1362,N_1298);
or U1435 (N_1435,N_1205,N_1332);
or U1436 (N_1436,N_1392,N_1207);
and U1437 (N_1437,N_1358,N_1329);
nor U1438 (N_1438,N_1357,N_1258);
or U1439 (N_1439,N_1277,N_1317);
nor U1440 (N_1440,N_1309,N_1377);
or U1441 (N_1441,N_1324,N_1344);
nor U1442 (N_1442,N_1229,N_1311);
and U1443 (N_1443,N_1373,N_1350);
nor U1444 (N_1444,N_1304,N_1379);
or U1445 (N_1445,N_1374,N_1307);
nand U1446 (N_1446,N_1355,N_1301);
or U1447 (N_1447,N_1370,N_1315);
nand U1448 (N_1448,N_1371,N_1354);
nand U1449 (N_1449,N_1352,N_1346);
nor U1450 (N_1450,N_1360,N_1269);
and U1451 (N_1451,N_1299,N_1333);
and U1452 (N_1452,N_1284,N_1382);
and U1453 (N_1453,N_1255,N_1268);
nor U1454 (N_1454,N_1227,N_1215);
or U1455 (N_1455,N_1336,N_1386);
nand U1456 (N_1456,N_1281,N_1248);
nor U1457 (N_1457,N_1380,N_1226);
or U1458 (N_1458,N_1365,N_1235);
or U1459 (N_1459,N_1273,N_1369);
or U1460 (N_1460,N_1251,N_1390);
nor U1461 (N_1461,N_1249,N_1391);
nand U1462 (N_1462,N_1213,N_1245);
nand U1463 (N_1463,N_1291,N_1275);
and U1464 (N_1464,N_1325,N_1396);
and U1465 (N_1465,N_1210,N_1236);
or U1466 (N_1466,N_1201,N_1237);
or U1467 (N_1467,N_1319,N_1217);
nand U1468 (N_1468,N_1398,N_1230);
or U1469 (N_1469,N_1219,N_1395);
or U1470 (N_1470,N_1224,N_1218);
or U1471 (N_1471,N_1239,N_1263);
or U1472 (N_1472,N_1306,N_1361);
nand U1473 (N_1473,N_1343,N_1314);
and U1474 (N_1474,N_1272,N_1259);
and U1475 (N_1475,N_1225,N_1393);
nor U1476 (N_1476,N_1326,N_1238);
nand U1477 (N_1477,N_1359,N_1367);
or U1478 (N_1478,N_1285,N_1265);
and U1479 (N_1479,N_1302,N_1381);
or U1480 (N_1480,N_1203,N_1266);
nand U1481 (N_1481,N_1305,N_1261);
or U1482 (N_1482,N_1242,N_1221);
nor U1483 (N_1483,N_1271,N_1283);
nand U1484 (N_1484,N_1260,N_1342);
or U1485 (N_1485,N_1252,N_1389);
and U1486 (N_1486,N_1282,N_1399);
and U1487 (N_1487,N_1310,N_1364);
and U1488 (N_1488,N_1345,N_1232);
and U1489 (N_1489,N_1322,N_1397);
or U1490 (N_1490,N_1387,N_1278);
or U1491 (N_1491,N_1347,N_1334);
or U1492 (N_1492,N_1244,N_1253);
and U1493 (N_1493,N_1388,N_1200);
or U1494 (N_1494,N_1383,N_1323);
and U1495 (N_1495,N_1270,N_1335);
or U1496 (N_1496,N_1366,N_1300);
nand U1497 (N_1497,N_1216,N_1274);
nand U1498 (N_1498,N_1209,N_1247);
nand U1499 (N_1499,N_1292,N_1296);
nor U1500 (N_1500,N_1284,N_1337);
or U1501 (N_1501,N_1223,N_1279);
and U1502 (N_1502,N_1228,N_1326);
nand U1503 (N_1503,N_1253,N_1363);
or U1504 (N_1504,N_1346,N_1342);
or U1505 (N_1505,N_1287,N_1303);
nor U1506 (N_1506,N_1206,N_1216);
nand U1507 (N_1507,N_1351,N_1261);
nor U1508 (N_1508,N_1245,N_1209);
nor U1509 (N_1509,N_1311,N_1279);
or U1510 (N_1510,N_1373,N_1353);
or U1511 (N_1511,N_1328,N_1374);
or U1512 (N_1512,N_1265,N_1266);
and U1513 (N_1513,N_1305,N_1283);
nor U1514 (N_1514,N_1331,N_1395);
nand U1515 (N_1515,N_1380,N_1313);
nor U1516 (N_1516,N_1286,N_1361);
and U1517 (N_1517,N_1229,N_1363);
and U1518 (N_1518,N_1227,N_1345);
and U1519 (N_1519,N_1358,N_1306);
nor U1520 (N_1520,N_1253,N_1333);
nor U1521 (N_1521,N_1310,N_1248);
or U1522 (N_1522,N_1329,N_1366);
nor U1523 (N_1523,N_1376,N_1362);
nand U1524 (N_1524,N_1360,N_1266);
nor U1525 (N_1525,N_1398,N_1345);
nor U1526 (N_1526,N_1313,N_1225);
nor U1527 (N_1527,N_1209,N_1377);
or U1528 (N_1528,N_1380,N_1275);
and U1529 (N_1529,N_1392,N_1380);
or U1530 (N_1530,N_1229,N_1271);
and U1531 (N_1531,N_1373,N_1253);
nand U1532 (N_1532,N_1312,N_1232);
nor U1533 (N_1533,N_1312,N_1341);
and U1534 (N_1534,N_1306,N_1293);
nand U1535 (N_1535,N_1360,N_1346);
or U1536 (N_1536,N_1376,N_1307);
or U1537 (N_1537,N_1391,N_1245);
or U1538 (N_1538,N_1381,N_1351);
or U1539 (N_1539,N_1235,N_1335);
nor U1540 (N_1540,N_1358,N_1322);
or U1541 (N_1541,N_1287,N_1328);
nand U1542 (N_1542,N_1320,N_1367);
nand U1543 (N_1543,N_1378,N_1247);
or U1544 (N_1544,N_1348,N_1212);
or U1545 (N_1545,N_1335,N_1381);
nand U1546 (N_1546,N_1231,N_1307);
and U1547 (N_1547,N_1278,N_1301);
or U1548 (N_1548,N_1277,N_1379);
and U1549 (N_1549,N_1352,N_1250);
nor U1550 (N_1550,N_1255,N_1211);
and U1551 (N_1551,N_1261,N_1226);
nand U1552 (N_1552,N_1330,N_1240);
and U1553 (N_1553,N_1334,N_1382);
or U1554 (N_1554,N_1296,N_1355);
nor U1555 (N_1555,N_1270,N_1389);
and U1556 (N_1556,N_1230,N_1338);
nand U1557 (N_1557,N_1227,N_1275);
nand U1558 (N_1558,N_1206,N_1219);
nor U1559 (N_1559,N_1362,N_1244);
and U1560 (N_1560,N_1284,N_1338);
or U1561 (N_1561,N_1214,N_1257);
and U1562 (N_1562,N_1280,N_1273);
or U1563 (N_1563,N_1314,N_1338);
nand U1564 (N_1564,N_1209,N_1248);
nor U1565 (N_1565,N_1268,N_1277);
nor U1566 (N_1566,N_1202,N_1214);
nor U1567 (N_1567,N_1395,N_1362);
or U1568 (N_1568,N_1328,N_1394);
nor U1569 (N_1569,N_1384,N_1244);
nand U1570 (N_1570,N_1383,N_1213);
nor U1571 (N_1571,N_1368,N_1353);
and U1572 (N_1572,N_1309,N_1394);
or U1573 (N_1573,N_1216,N_1254);
nand U1574 (N_1574,N_1375,N_1373);
nand U1575 (N_1575,N_1245,N_1253);
or U1576 (N_1576,N_1353,N_1291);
or U1577 (N_1577,N_1230,N_1203);
or U1578 (N_1578,N_1314,N_1242);
or U1579 (N_1579,N_1282,N_1378);
and U1580 (N_1580,N_1389,N_1239);
nor U1581 (N_1581,N_1346,N_1319);
and U1582 (N_1582,N_1277,N_1382);
nand U1583 (N_1583,N_1219,N_1345);
nand U1584 (N_1584,N_1260,N_1387);
nor U1585 (N_1585,N_1255,N_1326);
or U1586 (N_1586,N_1355,N_1263);
or U1587 (N_1587,N_1363,N_1328);
nand U1588 (N_1588,N_1267,N_1281);
and U1589 (N_1589,N_1355,N_1369);
or U1590 (N_1590,N_1307,N_1241);
or U1591 (N_1591,N_1261,N_1218);
nand U1592 (N_1592,N_1372,N_1242);
or U1593 (N_1593,N_1251,N_1329);
or U1594 (N_1594,N_1374,N_1261);
nand U1595 (N_1595,N_1340,N_1255);
and U1596 (N_1596,N_1249,N_1223);
nor U1597 (N_1597,N_1237,N_1355);
nand U1598 (N_1598,N_1340,N_1228);
or U1599 (N_1599,N_1325,N_1330);
nor U1600 (N_1600,N_1543,N_1456);
or U1601 (N_1601,N_1575,N_1499);
and U1602 (N_1602,N_1412,N_1465);
and U1603 (N_1603,N_1559,N_1497);
and U1604 (N_1604,N_1410,N_1420);
and U1605 (N_1605,N_1523,N_1562);
nand U1606 (N_1606,N_1544,N_1529);
nand U1607 (N_1607,N_1560,N_1443);
or U1608 (N_1608,N_1549,N_1405);
nand U1609 (N_1609,N_1589,N_1563);
nor U1610 (N_1610,N_1434,N_1453);
and U1611 (N_1611,N_1561,N_1422);
nand U1612 (N_1612,N_1579,N_1552);
nor U1613 (N_1613,N_1598,N_1502);
or U1614 (N_1614,N_1492,N_1429);
nor U1615 (N_1615,N_1483,N_1512);
or U1616 (N_1616,N_1490,N_1546);
nor U1617 (N_1617,N_1468,N_1461);
or U1618 (N_1618,N_1557,N_1566);
nand U1619 (N_1619,N_1573,N_1572);
nand U1620 (N_1620,N_1431,N_1510);
or U1621 (N_1621,N_1505,N_1592);
or U1622 (N_1622,N_1463,N_1467);
and U1623 (N_1623,N_1588,N_1577);
or U1624 (N_1624,N_1508,N_1484);
nand U1625 (N_1625,N_1582,N_1433);
and U1626 (N_1626,N_1509,N_1516);
nand U1627 (N_1627,N_1578,N_1511);
and U1628 (N_1628,N_1556,N_1459);
and U1629 (N_1629,N_1481,N_1406);
or U1630 (N_1630,N_1494,N_1548);
nor U1631 (N_1631,N_1518,N_1547);
and U1632 (N_1632,N_1574,N_1480);
nand U1633 (N_1633,N_1555,N_1527);
nor U1634 (N_1634,N_1435,N_1569);
nand U1635 (N_1635,N_1554,N_1482);
nor U1636 (N_1636,N_1571,N_1413);
or U1637 (N_1637,N_1564,N_1414);
nor U1638 (N_1638,N_1530,N_1583);
and U1639 (N_1639,N_1436,N_1584);
nand U1640 (N_1640,N_1596,N_1507);
or U1641 (N_1641,N_1477,N_1446);
nor U1642 (N_1642,N_1424,N_1432);
and U1643 (N_1643,N_1421,N_1528);
nor U1644 (N_1644,N_1464,N_1500);
and U1645 (N_1645,N_1550,N_1407);
nor U1646 (N_1646,N_1545,N_1402);
and U1647 (N_1647,N_1444,N_1495);
nand U1648 (N_1648,N_1452,N_1531);
nand U1649 (N_1649,N_1400,N_1417);
nand U1650 (N_1650,N_1441,N_1491);
nand U1651 (N_1651,N_1401,N_1440);
or U1652 (N_1652,N_1580,N_1462);
or U1653 (N_1653,N_1551,N_1524);
nand U1654 (N_1654,N_1455,N_1472);
and U1655 (N_1655,N_1597,N_1568);
or U1656 (N_1656,N_1447,N_1594);
nor U1657 (N_1657,N_1515,N_1487);
nand U1658 (N_1658,N_1590,N_1478);
and U1659 (N_1659,N_1586,N_1513);
nor U1660 (N_1660,N_1471,N_1595);
and U1661 (N_1661,N_1411,N_1454);
nor U1662 (N_1662,N_1520,N_1542);
nand U1663 (N_1663,N_1504,N_1427);
nand U1664 (N_1664,N_1591,N_1489);
or U1665 (N_1665,N_1522,N_1576);
and U1666 (N_1666,N_1458,N_1448);
nand U1667 (N_1667,N_1526,N_1460);
and U1668 (N_1668,N_1419,N_1532);
and U1669 (N_1669,N_1476,N_1585);
nand U1670 (N_1670,N_1470,N_1506);
and U1671 (N_1671,N_1537,N_1498);
and U1672 (N_1672,N_1485,N_1442);
nand U1673 (N_1673,N_1449,N_1514);
and U1674 (N_1674,N_1540,N_1474);
nand U1675 (N_1675,N_1565,N_1418);
and U1676 (N_1676,N_1593,N_1539);
and U1677 (N_1677,N_1533,N_1415);
nor U1678 (N_1678,N_1445,N_1581);
and U1679 (N_1679,N_1501,N_1469);
nand U1680 (N_1680,N_1541,N_1479);
nand U1681 (N_1681,N_1521,N_1486);
or U1682 (N_1682,N_1517,N_1475);
or U1683 (N_1683,N_1599,N_1493);
nand U1684 (N_1684,N_1525,N_1538);
nor U1685 (N_1685,N_1553,N_1437);
and U1686 (N_1686,N_1408,N_1519);
or U1687 (N_1687,N_1570,N_1503);
or U1688 (N_1688,N_1496,N_1567);
and U1689 (N_1689,N_1416,N_1536);
and U1690 (N_1690,N_1404,N_1450);
or U1691 (N_1691,N_1535,N_1409);
nand U1692 (N_1692,N_1473,N_1558);
and U1693 (N_1693,N_1430,N_1403);
nor U1694 (N_1694,N_1451,N_1587);
nand U1695 (N_1695,N_1438,N_1425);
and U1696 (N_1696,N_1534,N_1439);
and U1697 (N_1697,N_1428,N_1423);
nand U1698 (N_1698,N_1488,N_1466);
nor U1699 (N_1699,N_1426,N_1457);
or U1700 (N_1700,N_1504,N_1597);
nand U1701 (N_1701,N_1498,N_1459);
or U1702 (N_1702,N_1483,N_1549);
and U1703 (N_1703,N_1407,N_1525);
nor U1704 (N_1704,N_1541,N_1516);
and U1705 (N_1705,N_1422,N_1416);
and U1706 (N_1706,N_1496,N_1507);
or U1707 (N_1707,N_1567,N_1553);
or U1708 (N_1708,N_1447,N_1468);
and U1709 (N_1709,N_1455,N_1581);
and U1710 (N_1710,N_1585,N_1404);
or U1711 (N_1711,N_1522,N_1586);
nand U1712 (N_1712,N_1438,N_1428);
xor U1713 (N_1713,N_1405,N_1417);
and U1714 (N_1714,N_1444,N_1558);
and U1715 (N_1715,N_1564,N_1557);
nand U1716 (N_1716,N_1582,N_1593);
nand U1717 (N_1717,N_1515,N_1456);
or U1718 (N_1718,N_1452,N_1552);
and U1719 (N_1719,N_1401,N_1531);
nor U1720 (N_1720,N_1507,N_1451);
or U1721 (N_1721,N_1546,N_1521);
and U1722 (N_1722,N_1459,N_1589);
or U1723 (N_1723,N_1414,N_1527);
nor U1724 (N_1724,N_1564,N_1501);
nor U1725 (N_1725,N_1576,N_1557);
nor U1726 (N_1726,N_1455,N_1538);
and U1727 (N_1727,N_1577,N_1479);
and U1728 (N_1728,N_1521,N_1501);
and U1729 (N_1729,N_1504,N_1554);
and U1730 (N_1730,N_1468,N_1546);
nand U1731 (N_1731,N_1412,N_1452);
or U1732 (N_1732,N_1489,N_1437);
and U1733 (N_1733,N_1561,N_1428);
and U1734 (N_1734,N_1431,N_1462);
nand U1735 (N_1735,N_1595,N_1487);
or U1736 (N_1736,N_1587,N_1419);
nand U1737 (N_1737,N_1516,N_1470);
or U1738 (N_1738,N_1516,N_1432);
and U1739 (N_1739,N_1477,N_1542);
nand U1740 (N_1740,N_1432,N_1461);
nand U1741 (N_1741,N_1502,N_1431);
nor U1742 (N_1742,N_1460,N_1471);
nor U1743 (N_1743,N_1463,N_1419);
and U1744 (N_1744,N_1588,N_1496);
or U1745 (N_1745,N_1542,N_1424);
or U1746 (N_1746,N_1454,N_1405);
nand U1747 (N_1747,N_1535,N_1588);
nor U1748 (N_1748,N_1526,N_1490);
nand U1749 (N_1749,N_1428,N_1402);
or U1750 (N_1750,N_1567,N_1492);
nor U1751 (N_1751,N_1416,N_1463);
nand U1752 (N_1752,N_1588,N_1501);
or U1753 (N_1753,N_1435,N_1578);
or U1754 (N_1754,N_1415,N_1518);
nand U1755 (N_1755,N_1416,N_1597);
and U1756 (N_1756,N_1443,N_1425);
nand U1757 (N_1757,N_1423,N_1535);
nor U1758 (N_1758,N_1429,N_1451);
or U1759 (N_1759,N_1543,N_1446);
nand U1760 (N_1760,N_1539,N_1495);
or U1761 (N_1761,N_1550,N_1452);
nand U1762 (N_1762,N_1450,N_1453);
or U1763 (N_1763,N_1422,N_1479);
and U1764 (N_1764,N_1449,N_1542);
nor U1765 (N_1765,N_1578,N_1529);
and U1766 (N_1766,N_1514,N_1500);
nor U1767 (N_1767,N_1429,N_1422);
nand U1768 (N_1768,N_1404,N_1475);
and U1769 (N_1769,N_1499,N_1411);
nor U1770 (N_1770,N_1585,N_1597);
nor U1771 (N_1771,N_1468,N_1581);
and U1772 (N_1772,N_1547,N_1494);
and U1773 (N_1773,N_1527,N_1479);
and U1774 (N_1774,N_1430,N_1559);
and U1775 (N_1775,N_1408,N_1507);
nand U1776 (N_1776,N_1467,N_1490);
and U1777 (N_1777,N_1489,N_1421);
nor U1778 (N_1778,N_1439,N_1496);
or U1779 (N_1779,N_1454,N_1574);
and U1780 (N_1780,N_1417,N_1503);
nor U1781 (N_1781,N_1585,N_1440);
and U1782 (N_1782,N_1578,N_1468);
nor U1783 (N_1783,N_1565,N_1482);
nor U1784 (N_1784,N_1548,N_1584);
or U1785 (N_1785,N_1464,N_1591);
nand U1786 (N_1786,N_1401,N_1447);
and U1787 (N_1787,N_1504,N_1576);
nand U1788 (N_1788,N_1549,N_1558);
and U1789 (N_1789,N_1442,N_1588);
and U1790 (N_1790,N_1571,N_1417);
nor U1791 (N_1791,N_1597,N_1542);
nor U1792 (N_1792,N_1461,N_1458);
nand U1793 (N_1793,N_1517,N_1434);
or U1794 (N_1794,N_1455,N_1439);
or U1795 (N_1795,N_1409,N_1461);
nor U1796 (N_1796,N_1555,N_1442);
nand U1797 (N_1797,N_1585,N_1439);
and U1798 (N_1798,N_1415,N_1432);
nor U1799 (N_1799,N_1419,N_1599);
and U1800 (N_1800,N_1649,N_1777);
xor U1801 (N_1801,N_1755,N_1642);
nor U1802 (N_1802,N_1726,N_1632);
nand U1803 (N_1803,N_1651,N_1616);
or U1804 (N_1804,N_1779,N_1699);
nor U1805 (N_1805,N_1684,N_1712);
and U1806 (N_1806,N_1687,N_1697);
or U1807 (N_1807,N_1607,N_1770);
nor U1808 (N_1808,N_1794,N_1667);
nor U1809 (N_1809,N_1764,N_1768);
and U1810 (N_1810,N_1652,N_1724);
or U1811 (N_1811,N_1705,N_1692);
or U1812 (N_1812,N_1782,N_1745);
nand U1813 (N_1813,N_1661,N_1798);
and U1814 (N_1814,N_1716,N_1714);
or U1815 (N_1815,N_1696,N_1657);
or U1816 (N_1816,N_1763,N_1690);
nor U1817 (N_1817,N_1614,N_1709);
or U1818 (N_1818,N_1743,N_1753);
nand U1819 (N_1819,N_1767,N_1695);
and U1820 (N_1820,N_1731,N_1671);
nand U1821 (N_1821,N_1660,N_1707);
nor U1822 (N_1822,N_1757,N_1759);
and U1823 (N_1823,N_1674,N_1778);
nor U1824 (N_1824,N_1682,N_1703);
or U1825 (N_1825,N_1676,N_1750);
and U1826 (N_1826,N_1738,N_1748);
nand U1827 (N_1827,N_1694,N_1787);
and U1828 (N_1828,N_1605,N_1740);
nor U1829 (N_1829,N_1710,N_1762);
nor U1830 (N_1830,N_1776,N_1735);
and U1831 (N_1831,N_1727,N_1631);
nand U1832 (N_1832,N_1622,N_1636);
and U1833 (N_1833,N_1720,N_1633);
nor U1834 (N_1834,N_1683,N_1639);
and U1835 (N_1835,N_1698,N_1702);
or U1836 (N_1836,N_1733,N_1788);
nand U1837 (N_1837,N_1734,N_1773);
or U1838 (N_1838,N_1608,N_1637);
nor U1839 (N_1839,N_1715,N_1744);
nor U1840 (N_1840,N_1749,N_1623);
and U1841 (N_1841,N_1677,N_1789);
and U1842 (N_1842,N_1672,N_1790);
nor U1843 (N_1843,N_1793,N_1719);
or U1844 (N_1844,N_1747,N_1602);
or U1845 (N_1845,N_1601,N_1693);
nand U1846 (N_1846,N_1603,N_1626);
or U1847 (N_1847,N_1739,N_1795);
nand U1848 (N_1848,N_1722,N_1700);
xor U1849 (N_1849,N_1769,N_1765);
and U1850 (N_1850,N_1647,N_1675);
nor U1851 (N_1851,N_1756,N_1713);
and U1852 (N_1852,N_1600,N_1766);
and U1853 (N_1853,N_1730,N_1729);
and U1854 (N_1854,N_1617,N_1644);
and U1855 (N_1855,N_1742,N_1783);
nor U1856 (N_1856,N_1685,N_1641);
and U1857 (N_1857,N_1717,N_1658);
and U1858 (N_1858,N_1797,N_1654);
nand U1859 (N_1859,N_1728,N_1721);
nand U1860 (N_1860,N_1725,N_1781);
nand U1861 (N_1861,N_1799,N_1792);
nor U1862 (N_1862,N_1772,N_1691);
or U1863 (N_1863,N_1610,N_1686);
or U1864 (N_1864,N_1746,N_1643);
nor U1865 (N_1865,N_1665,N_1760);
and U1866 (N_1866,N_1638,N_1680);
nor U1867 (N_1867,N_1718,N_1784);
nand U1868 (N_1868,N_1736,N_1774);
nand U1869 (N_1869,N_1741,N_1678);
or U1870 (N_1870,N_1785,N_1621);
nand U1871 (N_1871,N_1648,N_1663);
and U1872 (N_1872,N_1612,N_1668);
and U1873 (N_1873,N_1619,N_1689);
or U1874 (N_1874,N_1655,N_1723);
nor U1875 (N_1875,N_1701,N_1673);
nor U1876 (N_1876,N_1625,N_1791);
nand U1877 (N_1877,N_1761,N_1662);
or U1878 (N_1878,N_1618,N_1620);
nor U1879 (N_1879,N_1606,N_1650);
nand U1880 (N_1880,N_1635,N_1627);
nor U1881 (N_1881,N_1737,N_1615);
nand U1882 (N_1882,N_1634,N_1664);
nor U1883 (N_1883,N_1624,N_1796);
or U1884 (N_1884,N_1670,N_1604);
or U1885 (N_1885,N_1708,N_1659);
or U1886 (N_1886,N_1688,N_1706);
nand U1887 (N_1887,N_1775,N_1629);
or U1888 (N_1888,N_1780,N_1704);
nand U1889 (N_1889,N_1640,N_1628);
nand U1890 (N_1890,N_1771,N_1630);
and U1891 (N_1891,N_1681,N_1656);
nor U1892 (N_1892,N_1613,N_1752);
nand U1893 (N_1893,N_1751,N_1758);
or U1894 (N_1894,N_1679,N_1786);
nand U1895 (N_1895,N_1611,N_1669);
nor U1896 (N_1896,N_1609,N_1653);
nand U1897 (N_1897,N_1732,N_1754);
nor U1898 (N_1898,N_1666,N_1646);
nor U1899 (N_1899,N_1711,N_1645);
and U1900 (N_1900,N_1699,N_1666);
nand U1901 (N_1901,N_1639,N_1791);
nand U1902 (N_1902,N_1694,N_1796);
nor U1903 (N_1903,N_1737,N_1680);
nand U1904 (N_1904,N_1689,N_1628);
and U1905 (N_1905,N_1666,N_1638);
nand U1906 (N_1906,N_1616,N_1722);
nand U1907 (N_1907,N_1638,N_1783);
nand U1908 (N_1908,N_1771,N_1689);
and U1909 (N_1909,N_1771,N_1739);
and U1910 (N_1910,N_1769,N_1744);
or U1911 (N_1911,N_1657,N_1784);
nor U1912 (N_1912,N_1627,N_1743);
nor U1913 (N_1913,N_1675,N_1676);
nand U1914 (N_1914,N_1605,N_1793);
and U1915 (N_1915,N_1710,N_1676);
nor U1916 (N_1916,N_1783,N_1619);
or U1917 (N_1917,N_1604,N_1715);
or U1918 (N_1918,N_1632,N_1713);
nor U1919 (N_1919,N_1650,N_1613);
nand U1920 (N_1920,N_1738,N_1742);
or U1921 (N_1921,N_1779,N_1619);
nor U1922 (N_1922,N_1785,N_1713);
nor U1923 (N_1923,N_1669,N_1782);
or U1924 (N_1924,N_1602,N_1757);
nor U1925 (N_1925,N_1799,N_1751);
nor U1926 (N_1926,N_1781,N_1619);
or U1927 (N_1927,N_1619,N_1736);
or U1928 (N_1928,N_1720,N_1682);
and U1929 (N_1929,N_1678,N_1613);
nor U1930 (N_1930,N_1720,N_1740);
nand U1931 (N_1931,N_1717,N_1657);
nand U1932 (N_1932,N_1653,N_1710);
nand U1933 (N_1933,N_1698,N_1675);
and U1934 (N_1934,N_1637,N_1613);
nand U1935 (N_1935,N_1771,N_1606);
and U1936 (N_1936,N_1747,N_1670);
nand U1937 (N_1937,N_1751,N_1730);
nand U1938 (N_1938,N_1639,N_1648);
or U1939 (N_1939,N_1717,N_1649);
nor U1940 (N_1940,N_1792,N_1779);
and U1941 (N_1941,N_1628,N_1696);
nand U1942 (N_1942,N_1742,N_1637);
and U1943 (N_1943,N_1601,N_1758);
or U1944 (N_1944,N_1767,N_1685);
nand U1945 (N_1945,N_1648,N_1756);
nand U1946 (N_1946,N_1653,N_1620);
and U1947 (N_1947,N_1725,N_1603);
nor U1948 (N_1948,N_1661,N_1765);
nor U1949 (N_1949,N_1669,N_1693);
nand U1950 (N_1950,N_1769,N_1793);
xor U1951 (N_1951,N_1738,N_1769);
nor U1952 (N_1952,N_1765,N_1757);
nand U1953 (N_1953,N_1736,N_1780);
nor U1954 (N_1954,N_1702,N_1694);
and U1955 (N_1955,N_1747,N_1711);
or U1956 (N_1956,N_1771,N_1758);
and U1957 (N_1957,N_1794,N_1681);
nor U1958 (N_1958,N_1731,N_1614);
nor U1959 (N_1959,N_1620,N_1786);
and U1960 (N_1960,N_1656,N_1754);
and U1961 (N_1961,N_1642,N_1628);
and U1962 (N_1962,N_1792,N_1651);
or U1963 (N_1963,N_1692,N_1654);
and U1964 (N_1964,N_1744,N_1639);
nand U1965 (N_1965,N_1675,N_1747);
and U1966 (N_1966,N_1709,N_1609);
nand U1967 (N_1967,N_1664,N_1733);
nand U1968 (N_1968,N_1775,N_1798);
nor U1969 (N_1969,N_1755,N_1656);
or U1970 (N_1970,N_1754,N_1654);
or U1971 (N_1971,N_1768,N_1603);
and U1972 (N_1972,N_1637,N_1601);
and U1973 (N_1973,N_1703,N_1679);
and U1974 (N_1974,N_1743,N_1644);
nand U1975 (N_1975,N_1767,N_1715);
nand U1976 (N_1976,N_1698,N_1755);
and U1977 (N_1977,N_1640,N_1635);
nand U1978 (N_1978,N_1758,N_1794);
nand U1979 (N_1979,N_1731,N_1718);
nand U1980 (N_1980,N_1631,N_1626);
nand U1981 (N_1981,N_1675,N_1662);
nand U1982 (N_1982,N_1654,N_1775);
and U1983 (N_1983,N_1701,N_1672);
nand U1984 (N_1984,N_1703,N_1726);
nand U1985 (N_1985,N_1717,N_1724);
nor U1986 (N_1986,N_1746,N_1726);
and U1987 (N_1987,N_1775,N_1694);
and U1988 (N_1988,N_1733,N_1637);
nand U1989 (N_1989,N_1799,N_1794);
nand U1990 (N_1990,N_1665,N_1610);
or U1991 (N_1991,N_1678,N_1714);
or U1992 (N_1992,N_1613,N_1664);
and U1993 (N_1993,N_1707,N_1619);
and U1994 (N_1994,N_1638,N_1611);
nor U1995 (N_1995,N_1635,N_1682);
and U1996 (N_1996,N_1765,N_1668);
and U1997 (N_1997,N_1718,N_1732);
or U1998 (N_1998,N_1713,N_1656);
nand U1999 (N_1999,N_1655,N_1604);
nor U2000 (N_2000,N_1810,N_1901);
and U2001 (N_2001,N_1986,N_1809);
or U2002 (N_2002,N_1814,N_1918);
and U2003 (N_2003,N_1840,N_1822);
and U2004 (N_2004,N_1849,N_1939);
or U2005 (N_2005,N_1862,N_1837);
and U2006 (N_2006,N_1905,N_1916);
nand U2007 (N_2007,N_1854,N_1988);
and U2008 (N_2008,N_1953,N_1893);
or U2009 (N_2009,N_1925,N_1870);
nor U2010 (N_2010,N_1895,N_1864);
nor U2011 (N_2011,N_1920,N_1890);
nand U2012 (N_2012,N_1894,N_1931);
or U2013 (N_2013,N_1872,N_1947);
nor U2014 (N_2014,N_1891,N_1929);
or U2015 (N_2015,N_1892,N_1844);
and U2016 (N_2016,N_1961,N_1818);
nand U2017 (N_2017,N_1817,N_1990);
nor U2018 (N_2018,N_1982,N_1908);
and U2019 (N_2019,N_1806,N_1911);
nand U2020 (N_2020,N_1820,N_1977);
nor U2021 (N_2021,N_1847,N_1996);
and U2022 (N_2022,N_1898,N_1968);
or U2023 (N_2023,N_1955,N_1994);
or U2024 (N_2024,N_1976,N_1811);
nor U2025 (N_2025,N_1960,N_1980);
and U2026 (N_2026,N_1924,N_1951);
nand U2027 (N_2027,N_1825,N_1850);
xor U2028 (N_2028,N_1867,N_1950);
or U2029 (N_2029,N_1896,N_1903);
and U2030 (N_2030,N_1804,N_1910);
nand U2031 (N_2031,N_1860,N_1832);
and U2032 (N_2032,N_1937,N_1859);
nand U2033 (N_2033,N_1846,N_1882);
and U2034 (N_2034,N_1812,N_1973);
nor U2035 (N_2035,N_1971,N_1970);
and U2036 (N_2036,N_1871,N_1841);
or U2037 (N_2037,N_1866,N_1800);
and U2038 (N_2038,N_1972,N_1808);
nor U2039 (N_2039,N_1992,N_1865);
nand U2040 (N_2040,N_1965,N_1946);
or U2041 (N_2041,N_1828,N_1874);
and U2042 (N_2042,N_1926,N_1909);
nand U2043 (N_2043,N_1873,N_1858);
and U2044 (N_2044,N_1824,N_1885);
or U2045 (N_2045,N_1819,N_1984);
nor U2046 (N_2046,N_1801,N_1839);
nand U2047 (N_2047,N_1944,N_1821);
and U2048 (N_2048,N_1881,N_1975);
and U2049 (N_2049,N_1948,N_1834);
and U2050 (N_2050,N_1845,N_1987);
nor U2051 (N_2051,N_1836,N_1856);
nor U2052 (N_2052,N_1998,N_1938);
or U2053 (N_2053,N_1989,N_1848);
nor U2054 (N_2054,N_1857,N_1978);
nand U2055 (N_2055,N_1981,N_1863);
or U2056 (N_2056,N_1922,N_1805);
or U2057 (N_2057,N_1803,N_1843);
or U2058 (N_2058,N_1967,N_1949);
nor U2059 (N_2059,N_1974,N_1927);
nor U2060 (N_2060,N_1838,N_1879);
nand U2061 (N_2061,N_1969,N_1983);
or U2062 (N_2062,N_1878,N_1868);
nor U2063 (N_2063,N_1889,N_1830);
nor U2064 (N_2064,N_1993,N_1919);
or U2065 (N_2065,N_1827,N_1935);
nand U2066 (N_2066,N_1876,N_1835);
and U2067 (N_2067,N_1963,N_1952);
and U2068 (N_2068,N_1934,N_1979);
nor U2069 (N_2069,N_1831,N_1900);
and U2070 (N_2070,N_1997,N_1855);
or U2071 (N_2071,N_1884,N_1906);
and U2072 (N_2072,N_1807,N_1962);
nand U2073 (N_2073,N_1958,N_1802);
nor U2074 (N_2074,N_1833,N_1959);
nand U2075 (N_2075,N_1851,N_1930);
nand U2076 (N_2076,N_1928,N_1936);
nor U2077 (N_2077,N_1914,N_1912);
and U2078 (N_2078,N_1941,N_1823);
nand U2079 (N_2079,N_1957,N_1877);
or U2080 (N_2080,N_1964,N_1815);
or U2081 (N_2081,N_1853,N_1888);
nor U2082 (N_2082,N_1917,N_1933);
nand U2083 (N_2083,N_1932,N_1897);
or U2084 (N_2084,N_1875,N_1943);
and U2085 (N_2085,N_1829,N_1880);
nor U2086 (N_2086,N_1869,N_1813);
xnor U2087 (N_2087,N_1985,N_1945);
nand U2088 (N_2088,N_1904,N_1883);
and U2089 (N_2089,N_1995,N_1956);
or U2090 (N_2090,N_1991,N_1942);
nor U2091 (N_2091,N_1999,N_1921);
nor U2092 (N_2092,N_1940,N_1923);
and U2093 (N_2093,N_1816,N_1887);
nand U2094 (N_2094,N_1852,N_1907);
or U2095 (N_2095,N_1902,N_1954);
nor U2096 (N_2096,N_1826,N_1899);
nor U2097 (N_2097,N_1842,N_1913);
and U2098 (N_2098,N_1915,N_1861);
and U2099 (N_2099,N_1966,N_1886);
nor U2100 (N_2100,N_1996,N_1946);
and U2101 (N_2101,N_1965,N_1951);
or U2102 (N_2102,N_1882,N_1907);
nand U2103 (N_2103,N_1802,N_1894);
or U2104 (N_2104,N_1896,N_1920);
and U2105 (N_2105,N_1824,N_1902);
or U2106 (N_2106,N_1926,N_1870);
and U2107 (N_2107,N_1988,N_1869);
nand U2108 (N_2108,N_1885,N_1843);
or U2109 (N_2109,N_1941,N_1963);
nor U2110 (N_2110,N_1818,N_1819);
nor U2111 (N_2111,N_1857,N_1838);
and U2112 (N_2112,N_1903,N_1980);
and U2113 (N_2113,N_1973,N_1925);
and U2114 (N_2114,N_1928,N_1940);
nor U2115 (N_2115,N_1961,N_1938);
or U2116 (N_2116,N_1801,N_1994);
or U2117 (N_2117,N_1938,N_1920);
and U2118 (N_2118,N_1975,N_1970);
and U2119 (N_2119,N_1871,N_1848);
nor U2120 (N_2120,N_1801,N_1842);
nand U2121 (N_2121,N_1866,N_1875);
xor U2122 (N_2122,N_1877,N_1941);
nand U2123 (N_2123,N_1860,N_1852);
nand U2124 (N_2124,N_1943,N_1877);
nand U2125 (N_2125,N_1814,N_1835);
or U2126 (N_2126,N_1902,N_1837);
nand U2127 (N_2127,N_1811,N_1834);
nor U2128 (N_2128,N_1944,N_1950);
and U2129 (N_2129,N_1946,N_1801);
nor U2130 (N_2130,N_1890,N_1805);
nand U2131 (N_2131,N_1882,N_1912);
or U2132 (N_2132,N_1979,N_1990);
nor U2133 (N_2133,N_1811,N_1861);
and U2134 (N_2134,N_1881,N_1839);
nor U2135 (N_2135,N_1861,N_1821);
and U2136 (N_2136,N_1983,N_1839);
or U2137 (N_2137,N_1805,N_1863);
nand U2138 (N_2138,N_1801,N_1840);
nor U2139 (N_2139,N_1908,N_1926);
or U2140 (N_2140,N_1997,N_1840);
nor U2141 (N_2141,N_1977,N_1922);
nor U2142 (N_2142,N_1966,N_1962);
and U2143 (N_2143,N_1963,N_1926);
nor U2144 (N_2144,N_1837,N_1918);
and U2145 (N_2145,N_1958,N_1910);
or U2146 (N_2146,N_1922,N_1810);
nand U2147 (N_2147,N_1989,N_1900);
or U2148 (N_2148,N_1845,N_1946);
nor U2149 (N_2149,N_1913,N_1907);
and U2150 (N_2150,N_1806,N_1973);
nand U2151 (N_2151,N_1822,N_1856);
nand U2152 (N_2152,N_1849,N_1909);
or U2153 (N_2153,N_1837,N_1885);
nand U2154 (N_2154,N_1871,N_1831);
nand U2155 (N_2155,N_1995,N_1941);
nor U2156 (N_2156,N_1990,N_1810);
nand U2157 (N_2157,N_1956,N_1907);
or U2158 (N_2158,N_1893,N_1854);
nand U2159 (N_2159,N_1879,N_1815);
nor U2160 (N_2160,N_1973,N_1841);
nand U2161 (N_2161,N_1809,N_1931);
nor U2162 (N_2162,N_1860,N_1917);
nand U2163 (N_2163,N_1858,N_1979);
nor U2164 (N_2164,N_1951,N_1887);
and U2165 (N_2165,N_1851,N_1849);
nand U2166 (N_2166,N_1984,N_1977);
or U2167 (N_2167,N_1822,N_1971);
nor U2168 (N_2168,N_1880,N_1959);
nor U2169 (N_2169,N_1992,N_1859);
and U2170 (N_2170,N_1958,N_1963);
nand U2171 (N_2171,N_1961,N_1911);
nor U2172 (N_2172,N_1851,N_1960);
nand U2173 (N_2173,N_1924,N_1909);
nor U2174 (N_2174,N_1865,N_1868);
nand U2175 (N_2175,N_1827,N_1920);
and U2176 (N_2176,N_1866,N_1987);
nand U2177 (N_2177,N_1832,N_1950);
nand U2178 (N_2178,N_1897,N_1977);
nand U2179 (N_2179,N_1812,N_1902);
nand U2180 (N_2180,N_1980,N_1910);
nor U2181 (N_2181,N_1805,N_1964);
nand U2182 (N_2182,N_1867,N_1972);
and U2183 (N_2183,N_1822,N_1930);
nor U2184 (N_2184,N_1828,N_1823);
nand U2185 (N_2185,N_1907,N_1804);
nor U2186 (N_2186,N_1864,N_1983);
nand U2187 (N_2187,N_1807,N_1955);
or U2188 (N_2188,N_1940,N_1942);
or U2189 (N_2189,N_1835,N_1844);
nand U2190 (N_2190,N_1917,N_1915);
and U2191 (N_2191,N_1928,N_1976);
nor U2192 (N_2192,N_1984,N_1855);
nand U2193 (N_2193,N_1848,N_1886);
and U2194 (N_2194,N_1821,N_1839);
nor U2195 (N_2195,N_1820,N_1991);
xnor U2196 (N_2196,N_1862,N_1883);
nor U2197 (N_2197,N_1882,N_1967);
nand U2198 (N_2198,N_1911,N_1919);
nor U2199 (N_2199,N_1997,N_1839);
or U2200 (N_2200,N_2105,N_2055);
nand U2201 (N_2201,N_2136,N_2109);
xnor U2202 (N_2202,N_2038,N_2159);
or U2203 (N_2203,N_2131,N_2069);
nor U2204 (N_2204,N_2047,N_2006);
nand U2205 (N_2205,N_2106,N_2120);
nor U2206 (N_2206,N_2165,N_2097);
or U2207 (N_2207,N_2128,N_2023);
nor U2208 (N_2208,N_2124,N_2086);
nor U2209 (N_2209,N_2091,N_2149);
or U2210 (N_2210,N_2166,N_2169);
and U2211 (N_2211,N_2014,N_2044);
nand U2212 (N_2212,N_2087,N_2154);
or U2213 (N_2213,N_2019,N_2049);
or U2214 (N_2214,N_2092,N_2164);
or U2215 (N_2215,N_2057,N_2155);
nand U2216 (N_2216,N_2017,N_2041);
nand U2217 (N_2217,N_2065,N_2093);
and U2218 (N_2218,N_2193,N_2148);
nor U2219 (N_2219,N_2002,N_2113);
nand U2220 (N_2220,N_2170,N_2103);
nand U2221 (N_2221,N_2062,N_2110);
or U2222 (N_2222,N_2009,N_2172);
nor U2223 (N_2223,N_2024,N_2050);
nor U2224 (N_2224,N_2130,N_2146);
nor U2225 (N_2225,N_2151,N_2081);
nand U2226 (N_2226,N_2080,N_2001);
and U2227 (N_2227,N_2076,N_2084);
or U2228 (N_2228,N_2075,N_2039);
nand U2229 (N_2229,N_2101,N_2175);
nor U2230 (N_2230,N_2085,N_2178);
and U2231 (N_2231,N_2192,N_2063);
nor U2232 (N_2232,N_2000,N_2071);
nor U2233 (N_2233,N_2189,N_2121);
or U2234 (N_2234,N_2020,N_2135);
nand U2235 (N_2235,N_2045,N_2030);
nand U2236 (N_2236,N_2174,N_2031);
nor U2237 (N_2237,N_2122,N_2168);
or U2238 (N_2238,N_2051,N_2138);
and U2239 (N_2239,N_2025,N_2162);
and U2240 (N_2240,N_2104,N_2013);
or U2241 (N_2241,N_2005,N_2177);
or U2242 (N_2242,N_2119,N_2056);
nand U2243 (N_2243,N_2052,N_2118);
or U2244 (N_2244,N_2107,N_2141);
nor U2245 (N_2245,N_2046,N_2067);
and U2246 (N_2246,N_2018,N_2197);
nand U2247 (N_2247,N_2117,N_2043);
xnor U2248 (N_2248,N_2072,N_2026);
nor U2249 (N_2249,N_2012,N_2035);
nor U2250 (N_2250,N_2060,N_2089);
and U2251 (N_2251,N_2161,N_2042);
nand U2252 (N_2252,N_2028,N_2132);
nor U2253 (N_2253,N_2088,N_2129);
or U2254 (N_2254,N_2167,N_2112);
and U2255 (N_2255,N_2139,N_2079);
and U2256 (N_2256,N_2143,N_2094);
nand U2257 (N_2257,N_2163,N_2077);
and U2258 (N_2258,N_2029,N_2115);
or U2259 (N_2259,N_2082,N_2054);
or U2260 (N_2260,N_2066,N_2040);
or U2261 (N_2261,N_2007,N_2058);
nor U2262 (N_2262,N_2083,N_2059);
and U2263 (N_2263,N_2156,N_2195);
or U2264 (N_2264,N_2183,N_2036);
and U2265 (N_2265,N_2003,N_2199);
nand U2266 (N_2266,N_2090,N_2158);
and U2267 (N_2267,N_2179,N_2140);
or U2268 (N_2268,N_2116,N_2171);
or U2269 (N_2269,N_2098,N_2188);
and U2270 (N_2270,N_2078,N_2111);
nor U2271 (N_2271,N_2181,N_2187);
or U2272 (N_2272,N_2191,N_2037);
nand U2273 (N_2273,N_2185,N_2182);
or U2274 (N_2274,N_2176,N_2074);
nand U2275 (N_2275,N_2150,N_2095);
or U2276 (N_2276,N_2016,N_2021);
nor U2277 (N_2277,N_2198,N_2033);
nor U2278 (N_2278,N_2142,N_2190);
nor U2279 (N_2279,N_2196,N_2137);
and U2280 (N_2280,N_2061,N_2125);
or U2281 (N_2281,N_2015,N_2004);
nand U2282 (N_2282,N_2186,N_2010);
or U2283 (N_2283,N_2068,N_2160);
nor U2284 (N_2284,N_2184,N_2008);
nor U2285 (N_2285,N_2053,N_2133);
nor U2286 (N_2286,N_2034,N_2070);
and U2287 (N_2287,N_2064,N_2127);
nand U2288 (N_2288,N_2180,N_2152);
or U2289 (N_2289,N_2173,N_2145);
nand U2290 (N_2290,N_2022,N_2126);
or U2291 (N_2291,N_2134,N_2123);
nor U2292 (N_2292,N_2144,N_2157);
xnor U2293 (N_2293,N_2100,N_2147);
nand U2294 (N_2294,N_2032,N_2194);
or U2295 (N_2295,N_2099,N_2108);
and U2296 (N_2296,N_2027,N_2102);
nand U2297 (N_2297,N_2114,N_2073);
nand U2298 (N_2298,N_2011,N_2153);
and U2299 (N_2299,N_2048,N_2096);
and U2300 (N_2300,N_2043,N_2006);
nor U2301 (N_2301,N_2078,N_2076);
nor U2302 (N_2302,N_2139,N_2166);
and U2303 (N_2303,N_2079,N_2017);
nand U2304 (N_2304,N_2118,N_2167);
and U2305 (N_2305,N_2053,N_2151);
nor U2306 (N_2306,N_2114,N_2116);
and U2307 (N_2307,N_2140,N_2038);
and U2308 (N_2308,N_2074,N_2128);
nand U2309 (N_2309,N_2179,N_2121);
and U2310 (N_2310,N_2052,N_2057);
xnor U2311 (N_2311,N_2057,N_2038);
nand U2312 (N_2312,N_2048,N_2057);
and U2313 (N_2313,N_2118,N_2134);
and U2314 (N_2314,N_2096,N_2057);
or U2315 (N_2315,N_2082,N_2084);
nor U2316 (N_2316,N_2129,N_2189);
or U2317 (N_2317,N_2102,N_2014);
nor U2318 (N_2318,N_2103,N_2044);
and U2319 (N_2319,N_2108,N_2009);
nand U2320 (N_2320,N_2165,N_2001);
and U2321 (N_2321,N_2189,N_2096);
nor U2322 (N_2322,N_2120,N_2070);
nor U2323 (N_2323,N_2064,N_2120);
and U2324 (N_2324,N_2148,N_2156);
nand U2325 (N_2325,N_2083,N_2011);
and U2326 (N_2326,N_2175,N_2166);
and U2327 (N_2327,N_2017,N_2066);
nand U2328 (N_2328,N_2154,N_2108);
xnor U2329 (N_2329,N_2096,N_2050);
and U2330 (N_2330,N_2027,N_2074);
nand U2331 (N_2331,N_2132,N_2138);
nor U2332 (N_2332,N_2169,N_2059);
and U2333 (N_2333,N_2110,N_2096);
nand U2334 (N_2334,N_2184,N_2104);
nor U2335 (N_2335,N_2176,N_2068);
nand U2336 (N_2336,N_2159,N_2158);
and U2337 (N_2337,N_2198,N_2038);
and U2338 (N_2338,N_2075,N_2018);
nor U2339 (N_2339,N_2027,N_2082);
or U2340 (N_2340,N_2123,N_2078);
and U2341 (N_2341,N_2003,N_2005);
nor U2342 (N_2342,N_2067,N_2178);
and U2343 (N_2343,N_2090,N_2030);
nand U2344 (N_2344,N_2133,N_2194);
nor U2345 (N_2345,N_2120,N_2038);
nor U2346 (N_2346,N_2178,N_2145);
and U2347 (N_2347,N_2067,N_2164);
nand U2348 (N_2348,N_2144,N_2073);
or U2349 (N_2349,N_2092,N_2031);
nor U2350 (N_2350,N_2142,N_2084);
nor U2351 (N_2351,N_2075,N_2059);
nand U2352 (N_2352,N_2158,N_2083);
nor U2353 (N_2353,N_2100,N_2132);
nand U2354 (N_2354,N_2052,N_2189);
nand U2355 (N_2355,N_2171,N_2123);
or U2356 (N_2356,N_2187,N_2153);
nor U2357 (N_2357,N_2048,N_2169);
and U2358 (N_2358,N_2017,N_2028);
and U2359 (N_2359,N_2075,N_2190);
and U2360 (N_2360,N_2035,N_2072);
nor U2361 (N_2361,N_2195,N_2007);
or U2362 (N_2362,N_2190,N_2039);
nor U2363 (N_2363,N_2006,N_2087);
xnor U2364 (N_2364,N_2002,N_2051);
and U2365 (N_2365,N_2092,N_2175);
nand U2366 (N_2366,N_2174,N_2109);
or U2367 (N_2367,N_2074,N_2116);
nor U2368 (N_2368,N_2165,N_2114);
nand U2369 (N_2369,N_2187,N_2166);
and U2370 (N_2370,N_2020,N_2033);
nor U2371 (N_2371,N_2188,N_2103);
or U2372 (N_2372,N_2152,N_2150);
nor U2373 (N_2373,N_2092,N_2183);
and U2374 (N_2374,N_2050,N_2056);
and U2375 (N_2375,N_2157,N_2093);
or U2376 (N_2376,N_2183,N_2047);
nor U2377 (N_2377,N_2004,N_2082);
nand U2378 (N_2378,N_2114,N_2045);
nand U2379 (N_2379,N_2130,N_2048);
or U2380 (N_2380,N_2100,N_2077);
nor U2381 (N_2381,N_2009,N_2128);
nand U2382 (N_2382,N_2053,N_2085);
nor U2383 (N_2383,N_2175,N_2197);
nor U2384 (N_2384,N_2182,N_2130);
nor U2385 (N_2385,N_2198,N_2081);
or U2386 (N_2386,N_2088,N_2064);
nor U2387 (N_2387,N_2144,N_2001);
or U2388 (N_2388,N_2042,N_2188);
nor U2389 (N_2389,N_2196,N_2097);
and U2390 (N_2390,N_2108,N_2170);
nand U2391 (N_2391,N_2106,N_2064);
and U2392 (N_2392,N_2016,N_2075);
and U2393 (N_2393,N_2118,N_2181);
and U2394 (N_2394,N_2073,N_2078);
nand U2395 (N_2395,N_2065,N_2118);
nand U2396 (N_2396,N_2046,N_2129);
and U2397 (N_2397,N_2184,N_2126);
nor U2398 (N_2398,N_2038,N_2142);
nand U2399 (N_2399,N_2146,N_2149);
nand U2400 (N_2400,N_2311,N_2293);
and U2401 (N_2401,N_2325,N_2349);
nand U2402 (N_2402,N_2228,N_2300);
or U2403 (N_2403,N_2298,N_2370);
and U2404 (N_2404,N_2316,N_2253);
and U2405 (N_2405,N_2200,N_2202);
nor U2406 (N_2406,N_2248,N_2303);
and U2407 (N_2407,N_2317,N_2352);
or U2408 (N_2408,N_2267,N_2231);
or U2409 (N_2409,N_2206,N_2251);
or U2410 (N_2410,N_2380,N_2302);
nand U2411 (N_2411,N_2334,N_2338);
and U2412 (N_2412,N_2333,N_2262);
and U2413 (N_2413,N_2233,N_2383);
nand U2414 (N_2414,N_2250,N_2376);
or U2415 (N_2415,N_2244,N_2256);
and U2416 (N_2416,N_2221,N_2324);
or U2417 (N_2417,N_2345,N_2222);
or U2418 (N_2418,N_2315,N_2290);
nor U2419 (N_2419,N_2319,N_2393);
and U2420 (N_2420,N_2268,N_2361);
nor U2421 (N_2421,N_2309,N_2214);
or U2422 (N_2422,N_2378,N_2332);
nor U2423 (N_2423,N_2218,N_2275);
or U2424 (N_2424,N_2314,N_2264);
nor U2425 (N_2425,N_2364,N_2320);
or U2426 (N_2426,N_2367,N_2346);
xnor U2427 (N_2427,N_2295,N_2273);
or U2428 (N_2428,N_2296,N_2201);
or U2429 (N_2429,N_2260,N_2212);
nand U2430 (N_2430,N_2365,N_2271);
nor U2431 (N_2431,N_2209,N_2318);
and U2432 (N_2432,N_2213,N_2342);
nand U2433 (N_2433,N_2203,N_2355);
nand U2434 (N_2434,N_2226,N_2341);
or U2435 (N_2435,N_2286,N_2255);
or U2436 (N_2436,N_2230,N_2258);
or U2437 (N_2437,N_2284,N_2232);
or U2438 (N_2438,N_2220,N_2374);
and U2439 (N_2439,N_2216,N_2350);
or U2440 (N_2440,N_2331,N_2327);
nand U2441 (N_2441,N_2347,N_2301);
and U2442 (N_2442,N_2257,N_2348);
or U2443 (N_2443,N_2240,N_2289);
nand U2444 (N_2444,N_2351,N_2217);
and U2445 (N_2445,N_2340,N_2373);
and U2446 (N_2446,N_2357,N_2292);
or U2447 (N_2447,N_2313,N_2358);
or U2448 (N_2448,N_2278,N_2363);
and U2449 (N_2449,N_2238,N_2252);
and U2450 (N_2450,N_2321,N_2369);
or U2451 (N_2451,N_2368,N_2283);
and U2452 (N_2452,N_2398,N_2390);
or U2453 (N_2453,N_2245,N_2395);
nor U2454 (N_2454,N_2328,N_2263);
and U2455 (N_2455,N_2353,N_2297);
and U2456 (N_2456,N_2287,N_2385);
or U2457 (N_2457,N_2359,N_2239);
and U2458 (N_2458,N_2205,N_2396);
and U2459 (N_2459,N_2241,N_2399);
and U2460 (N_2460,N_2323,N_2277);
or U2461 (N_2461,N_2266,N_2386);
or U2462 (N_2462,N_2227,N_2392);
and U2463 (N_2463,N_2261,N_2215);
and U2464 (N_2464,N_2326,N_2308);
nor U2465 (N_2465,N_2279,N_2387);
nand U2466 (N_2466,N_2372,N_2339);
nand U2467 (N_2467,N_2354,N_2322);
nor U2468 (N_2468,N_2281,N_2285);
nor U2469 (N_2469,N_2288,N_2237);
and U2470 (N_2470,N_2280,N_2247);
or U2471 (N_2471,N_2259,N_2336);
nor U2472 (N_2472,N_2377,N_2305);
nor U2473 (N_2473,N_2330,N_2304);
nand U2474 (N_2474,N_2208,N_2270);
nand U2475 (N_2475,N_2379,N_2389);
nor U2476 (N_2476,N_2223,N_2356);
or U2477 (N_2477,N_2224,N_2344);
or U2478 (N_2478,N_2272,N_2312);
or U2479 (N_2479,N_2211,N_2242);
nor U2480 (N_2480,N_2360,N_2210);
or U2481 (N_2481,N_2249,N_2384);
and U2482 (N_2482,N_2307,N_2362);
and U2483 (N_2483,N_2306,N_2265);
or U2484 (N_2484,N_2343,N_2276);
or U2485 (N_2485,N_2207,N_2235);
or U2486 (N_2486,N_2254,N_2382);
xor U2487 (N_2487,N_2391,N_2371);
nor U2488 (N_2488,N_2204,N_2335);
and U2489 (N_2489,N_2234,N_2269);
nand U2490 (N_2490,N_2225,N_2388);
or U2491 (N_2491,N_2299,N_2397);
nand U2492 (N_2492,N_2291,N_2394);
nand U2493 (N_2493,N_2243,N_2366);
and U2494 (N_2494,N_2375,N_2381);
nand U2495 (N_2495,N_2229,N_2236);
or U2496 (N_2496,N_2329,N_2219);
nor U2497 (N_2497,N_2310,N_2246);
or U2498 (N_2498,N_2274,N_2282);
nor U2499 (N_2499,N_2337,N_2294);
nand U2500 (N_2500,N_2298,N_2387);
nor U2501 (N_2501,N_2293,N_2396);
or U2502 (N_2502,N_2335,N_2365);
and U2503 (N_2503,N_2328,N_2241);
or U2504 (N_2504,N_2354,N_2346);
and U2505 (N_2505,N_2227,N_2209);
and U2506 (N_2506,N_2302,N_2269);
nand U2507 (N_2507,N_2259,N_2224);
nand U2508 (N_2508,N_2277,N_2267);
nand U2509 (N_2509,N_2274,N_2305);
nor U2510 (N_2510,N_2399,N_2363);
and U2511 (N_2511,N_2204,N_2381);
or U2512 (N_2512,N_2349,N_2224);
and U2513 (N_2513,N_2346,N_2278);
and U2514 (N_2514,N_2270,N_2350);
nand U2515 (N_2515,N_2283,N_2353);
or U2516 (N_2516,N_2357,N_2310);
and U2517 (N_2517,N_2290,N_2353);
and U2518 (N_2518,N_2276,N_2341);
nor U2519 (N_2519,N_2292,N_2308);
nor U2520 (N_2520,N_2230,N_2330);
and U2521 (N_2521,N_2394,N_2206);
nor U2522 (N_2522,N_2279,N_2386);
nand U2523 (N_2523,N_2380,N_2244);
nand U2524 (N_2524,N_2291,N_2339);
or U2525 (N_2525,N_2212,N_2238);
or U2526 (N_2526,N_2242,N_2273);
nor U2527 (N_2527,N_2399,N_2362);
nand U2528 (N_2528,N_2241,N_2363);
nor U2529 (N_2529,N_2383,N_2374);
nand U2530 (N_2530,N_2335,N_2287);
and U2531 (N_2531,N_2328,N_2262);
or U2532 (N_2532,N_2279,N_2366);
and U2533 (N_2533,N_2397,N_2200);
nand U2534 (N_2534,N_2383,N_2320);
nor U2535 (N_2535,N_2368,N_2296);
nor U2536 (N_2536,N_2217,N_2235);
and U2537 (N_2537,N_2276,N_2371);
or U2538 (N_2538,N_2336,N_2223);
and U2539 (N_2539,N_2344,N_2288);
and U2540 (N_2540,N_2287,N_2387);
nand U2541 (N_2541,N_2303,N_2317);
and U2542 (N_2542,N_2235,N_2316);
and U2543 (N_2543,N_2379,N_2306);
nor U2544 (N_2544,N_2382,N_2375);
and U2545 (N_2545,N_2373,N_2376);
nand U2546 (N_2546,N_2356,N_2256);
and U2547 (N_2547,N_2348,N_2268);
and U2548 (N_2548,N_2256,N_2323);
and U2549 (N_2549,N_2290,N_2202);
and U2550 (N_2550,N_2225,N_2275);
and U2551 (N_2551,N_2217,N_2288);
and U2552 (N_2552,N_2240,N_2397);
nand U2553 (N_2553,N_2389,N_2331);
or U2554 (N_2554,N_2390,N_2366);
and U2555 (N_2555,N_2317,N_2211);
and U2556 (N_2556,N_2237,N_2250);
and U2557 (N_2557,N_2294,N_2361);
nor U2558 (N_2558,N_2284,N_2398);
nand U2559 (N_2559,N_2399,N_2217);
or U2560 (N_2560,N_2307,N_2232);
nand U2561 (N_2561,N_2375,N_2276);
and U2562 (N_2562,N_2200,N_2209);
nor U2563 (N_2563,N_2328,N_2326);
nand U2564 (N_2564,N_2268,N_2310);
or U2565 (N_2565,N_2321,N_2343);
and U2566 (N_2566,N_2311,N_2365);
nor U2567 (N_2567,N_2388,N_2245);
or U2568 (N_2568,N_2387,N_2356);
and U2569 (N_2569,N_2226,N_2300);
nor U2570 (N_2570,N_2331,N_2359);
or U2571 (N_2571,N_2247,N_2309);
nand U2572 (N_2572,N_2304,N_2208);
and U2573 (N_2573,N_2226,N_2258);
nor U2574 (N_2574,N_2332,N_2203);
and U2575 (N_2575,N_2371,N_2330);
and U2576 (N_2576,N_2336,N_2241);
xnor U2577 (N_2577,N_2301,N_2368);
nor U2578 (N_2578,N_2235,N_2334);
or U2579 (N_2579,N_2348,N_2364);
nor U2580 (N_2580,N_2338,N_2360);
and U2581 (N_2581,N_2393,N_2372);
and U2582 (N_2582,N_2255,N_2257);
or U2583 (N_2583,N_2398,N_2256);
and U2584 (N_2584,N_2387,N_2352);
or U2585 (N_2585,N_2237,N_2345);
and U2586 (N_2586,N_2325,N_2311);
or U2587 (N_2587,N_2350,N_2373);
and U2588 (N_2588,N_2234,N_2384);
and U2589 (N_2589,N_2201,N_2207);
nor U2590 (N_2590,N_2363,N_2235);
nor U2591 (N_2591,N_2247,N_2327);
or U2592 (N_2592,N_2376,N_2263);
and U2593 (N_2593,N_2310,N_2276);
and U2594 (N_2594,N_2288,N_2282);
nand U2595 (N_2595,N_2225,N_2321);
nand U2596 (N_2596,N_2220,N_2324);
nor U2597 (N_2597,N_2261,N_2332);
and U2598 (N_2598,N_2347,N_2346);
nor U2599 (N_2599,N_2263,N_2220);
or U2600 (N_2600,N_2432,N_2494);
nor U2601 (N_2601,N_2582,N_2529);
nand U2602 (N_2602,N_2497,N_2403);
and U2603 (N_2603,N_2566,N_2577);
and U2604 (N_2604,N_2507,N_2477);
nor U2605 (N_2605,N_2446,N_2524);
xor U2606 (N_2606,N_2579,N_2487);
nor U2607 (N_2607,N_2453,N_2418);
or U2608 (N_2608,N_2421,N_2549);
and U2609 (N_2609,N_2483,N_2423);
or U2610 (N_2610,N_2503,N_2542);
and U2611 (N_2611,N_2518,N_2415);
nor U2612 (N_2612,N_2468,N_2545);
and U2613 (N_2613,N_2541,N_2420);
or U2614 (N_2614,N_2580,N_2523);
nor U2615 (N_2615,N_2561,N_2401);
nand U2616 (N_2616,N_2419,N_2445);
nor U2617 (N_2617,N_2478,N_2409);
nand U2618 (N_2618,N_2571,N_2526);
nor U2619 (N_2619,N_2572,N_2551);
nor U2620 (N_2620,N_2443,N_2560);
nand U2621 (N_2621,N_2575,N_2540);
xnor U2622 (N_2622,N_2476,N_2546);
and U2623 (N_2623,N_2480,N_2597);
nor U2624 (N_2624,N_2431,N_2511);
and U2625 (N_2625,N_2408,N_2563);
nor U2626 (N_2626,N_2467,N_2590);
or U2627 (N_2627,N_2469,N_2485);
xor U2628 (N_2628,N_2417,N_2425);
nor U2629 (N_2629,N_2500,N_2530);
or U2630 (N_2630,N_2581,N_2589);
or U2631 (N_2631,N_2525,N_2498);
nand U2632 (N_2632,N_2486,N_2558);
or U2633 (N_2633,N_2488,N_2442);
nor U2634 (N_2634,N_2439,N_2547);
nor U2635 (N_2635,N_2471,N_2510);
or U2636 (N_2636,N_2538,N_2482);
nor U2637 (N_2637,N_2521,N_2465);
or U2638 (N_2638,N_2461,N_2474);
nand U2639 (N_2639,N_2475,N_2596);
nor U2640 (N_2640,N_2522,N_2457);
and U2641 (N_2641,N_2472,N_2552);
nand U2642 (N_2642,N_2501,N_2490);
nand U2643 (N_2643,N_2506,N_2406);
nand U2644 (N_2644,N_2422,N_2481);
and U2645 (N_2645,N_2407,N_2584);
and U2646 (N_2646,N_2496,N_2412);
nand U2647 (N_2647,N_2489,N_2533);
or U2648 (N_2648,N_2514,N_2585);
and U2649 (N_2649,N_2413,N_2502);
and U2650 (N_2650,N_2554,N_2414);
nand U2651 (N_2651,N_2583,N_2527);
and U2652 (N_2652,N_2405,N_2567);
nor U2653 (N_2653,N_2534,N_2550);
nor U2654 (N_2654,N_2555,N_2404);
nor U2655 (N_2655,N_2433,N_2557);
nand U2656 (N_2656,N_2451,N_2536);
nor U2657 (N_2657,N_2479,N_2499);
and U2658 (N_2658,N_2473,N_2576);
and U2659 (N_2659,N_2456,N_2400);
nand U2660 (N_2660,N_2447,N_2569);
nor U2661 (N_2661,N_2444,N_2508);
and U2662 (N_2662,N_2568,N_2449);
and U2663 (N_2663,N_2428,N_2460);
or U2664 (N_2664,N_2435,N_2519);
nor U2665 (N_2665,N_2458,N_2573);
and U2666 (N_2666,N_2565,N_2470);
nand U2667 (N_2667,N_2416,N_2484);
and U2668 (N_2668,N_2429,N_2504);
nor U2669 (N_2669,N_2532,N_2448);
or U2670 (N_2670,N_2462,N_2559);
or U2671 (N_2671,N_2426,N_2593);
and U2672 (N_2672,N_2440,N_2513);
and U2673 (N_2673,N_2517,N_2556);
or U2674 (N_2674,N_2492,N_2537);
or U2675 (N_2675,N_2570,N_2539);
and U2676 (N_2676,N_2466,N_2450);
nand U2677 (N_2677,N_2544,N_2535);
nor U2678 (N_2678,N_2594,N_2553);
and U2679 (N_2679,N_2410,N_2454);
nor U2680 (N_2680,N_2588,N_2528);
and U2681 (N_2681,N_2512,N_2509);
nand U2682 (N_2682,N_2595,N_2437);
or U2683 (N_2683,N_2438,N_2586);
nand U2684 (N_2684,N_2402,N_2452);
and U2685 (N_2685,N_2520,N_2411);
and U2686 (N_2686,N_2587,N_2543);
nor U2687 (N_2687,N_2430,N_2455);
and U2688 (N_2688,N_2441,N_2531);
nand U2689 (N_2689,N_2434,N_2578);
or U2690 (N_2690,N_2591,N_2598);
nand U2691 (N_2691,N_2592,N_2599);
and U2692 (N_2692,N_2516,N_2548);
nor U2693 (N_2693,N_2505,N_2562);
and U2694 (N_2694,N_2459,N_2493);
nor U2695 (N_2695,N_2427,N_2464);
and U2696 (N_2696,N_2564,N_2436);
and U2697 (N_2697,N_2515,N_2424);
and U2698 (N_2698,N_2491,N_2574);
and U2699 (N_2699,N_2495,N_2463);
and U2700 (N_2700,N_2504,N_2591);
nor U2701 (N_2701,N_2583,N_2565);
nand U2702 (N_2702,N_2422,N_2474);
or U2703 (N_2703,N_2426,N_2442);
nand U2704 (N_2704,N_2403,N_2488);
nand U2705 (N_2705,N_2405,N_2498);
nand U2706 (N_2706,N_2473,N_2468);
nand U2707 (N_2707,N_2550,N_2429);
or U2708 (N_2708,N_2525,N_2528);
and U2709 (N_2709,N_2425,N_2451);
nand U2710 (N_2710,N_2568,N_2490);
and U2711 (N_2711,N_2456,N_2448);
nor U2712 (N_2712,N_2521,N_2440);
nand U2713 (N_2713,N_2572,N_2511);
nor U2714 (N_2714,N_2403,N_2547);
and U2715 (N_2715,N_2407,N_2491);
nand U2716 (N_2716,N_2400,N_2552);
and U2717 (N_2717,N_2467,N_2405);
or U2718 (N_2718,N_2530,N_2540);
nand U2719 (N_2719,N_2579,N_2581);
and U2720 (N_2720,N_2496,N_2581);
or U2721 (N_2721,N_2531,N_2482);
or U2722 (N_2722,N_2579,N_2441);
or U2723 (N_2723,N_2473,N_2417);
nor U2724 (N_2724,N_2477,N_2536);
or U2725 (N_2725,N_2506,N_2535);
and U2726 (N_2726,N_2483,N_2492);
nand U2727 (N_2727,N_2556,N_2445);
and U2728 (N_2728,N_2487,N_2457);
and U2729 (N_2729,N_2524,N_2501);
nor U2730 (N_2730,N_2427,N_2483);
nand U2731 (N_2731,N_2427,N_2522);
nand U2732 (N_2732,N_2574,N_2460);
nand U2733 (N_2733,N_2547,N_2498);
or U2734 (N_2734,N_2437,N_2438);
nand U2735 (N_2735,N_2567,N_2494);
and U2736 (N_2736,N_2453,N_2410);
or U2737 (N_2737,N_2539,N_2534);
nand U2738 (N_2738,N_2451,N_2436);
and U2739 (N_2739,N_2406,N_2474);
or U2740 (N_2740,N_2520,N_2565);
nand U2741 (N_2741,N_2526,N_2424);
and U2742 (N_2742,N_2525,N_2563);
or U2743 (N_2743,N_2564,N_2583);
nor U2744 (N_2744,N_2543,N_2447);
or U2745 (N_2745,N_2440,N_2486);
or U2746 (N_2746,N_2440,N_2527);
or U2747 (N_2747,N_2447,N_2504);
nor U2748 (N_2748,N_2444,N_2488);
and U2749 (N_2749,N_2498,N_2561);
and U2750 (N_2750,N_2406,N_2488);
nand U2751 (N_2751,N_2502,N_2461);
or U2752 (N_2752,N_2576,N_2438);
or U2753 (N_2753,N_2555,N_2510);
nand U2754 (N_2754,N_2563,N_2403);
or U2755 (N_2755,N_2594,N_2462);
and U2756 (N_2756,N_2499,N_2493);
or U2757 (N_2757,N_2537,N_2516);
nand U2758 (N_2758,N_2452,N_2472);
nor U2759 (N_2759,N_2532,N_2579);
or U2760 (N_2760,N_2466,N_2507);
and U2761 (N_2761,N_2509,N_2577);
nor U2762 (N_2762,N_2467,N_2456);
or U2763 (N_2763,N_2435,N_2569);
or U2764 (N_2764,N_2511,N_2545);
or U2765 (N_2765,N_2518,N_2559);
and U2766 (N_2766,N_2527,N_2560);
and U2767 (N_2767,N_2475,N_2518);
nor U2768 (N_2768,N_2486,N_2420);
or U2769 (N_2769,N_2417,N_2492);
or U2770 (N_2770,N_2496,N_2558);
nor U2771 (N_2771,N_2580,N_2540);
nor U2772 (N_2772,N_2559,N_2597);
nor U2773 (N_2773,N_2454,N_2513);
nor U2774 (N_2774,N_2446,N_2543);
nor U2775 (N_2775,N_2469,N_2475);
nand U2776 (N_2776,N_2578,N_2596);
or U2777 (N_2777,N_2458,N_2554);
or U2778 (N_2778,N_2515,N_2442);
or U2779 (N_2779,N_2410,N_2425);
nor U2780 (N_2780,N_2515,N_2563);
nand U2781 (N_2781,N_2563,N_2443);
nor U2782 (N_2782,N_2402,N_2531);
or U2783 (N_2783,N_2592,N_2491);
nor U2784 (N_2784,N_2433,N_2554);
nor U2785 (N_2785,N_2506,N_2503);
or U2786 (N_2786,N_2427,N_2500);
and U2787 (N_2787,N_2415,N_2559);
nor U2788 (N_2788,N_2535,N_2404);
and U2789 (N_2789,N_2550,N_2599);
nand U2790 (N_2790,N_2549,N_2485);
or U2791 (N_2791,N_2553,N_2561);
and U2792 (N_2792,N_2401,N_2505);
nand U2793 (N_2793,N_2401,N_2403);
nand U2794 (N_2794,N_2564,N_2571);
nor U2795 (N_2795,N_2438,N_2582);
or U2796 (N_2796,N_2462,N_2489);
nor U2797 (N_2797,N_2464,N_2485);
nand U2798 (N_2798,N_2496,N_2481);
and U2799 (N_2799,N_2526,N_2496);
nor U2800 (N_2800,N_2799,N_2643);
nand U2801 (N_2801,N_2683,N_2708);
or U2802 (N_2802,N_2775,N_2611);
nand U2803 (N_2803,N_2658,N_2759);
or U2804 (N_2804,N_2652,N_2665);
nor U2805 (N_2805,N_2688,N_2711);
and U2806 (N_2806,N_2614,N_2679);
or U2807 (N_2807,N_2649,N_2748);
or U2808 (N_2808,N_2603,N_2756);
nor U2809 (N_2809,N_2636,N_2639);
nand U2810 (N_2810,N_2776,N_2735);
and U2811 (N_2811,N_2684,N_2678);
nand U2812 (N_2812,N_2761,N_2731);
nor U2813 (N_2813,N_2606,N_2618);
nor U2814 (N_2814,N_2703,N_2721);
nand U2815 (N_2815,N_2734,N_2720);
and U2816 (N_2816,N_2637,N_2647);
nand U2817 (N_2817,N_2604,N_2763);
or U2818 (N_2818,N_2728,N_2737);
nand U2819 (N_2819,N_2723,N_2749);
or U2820 (N_2820,N_2693,N_2659);
nor U2821 (N_2821,N_2713,N_2782);
or U2822 (N_2822,N_2628,N_2709);
and U2823 (N_2823,N_2692,N_2675);
nor U2824 (N_2824,N_2668,N_2778);
or U2825 (N_2825,N_2654,N_2690);
nor U2826 (N_2826,N_2741,N_2793);
and U2827 (N_2827,N_2797,N_2780);
and U2828 (N_2828,N_2784,N_2712);
nor U2829 (N_2829,N_2733,N_2794);
or U2830 (N_2830,N_2661,N_2626);
or U2831 (N_2831,N_2791,N_2754);
or U2832 (N_2832,N_2732,N_2624);
nor U2833 (N_2833,N_2673,N_2601);
or U2834 (N_2834,N_2613,N_2669);
nor U2835 (N_2835,N_2788,N_2621);
or U2836 (N_2836,N_2750,N_2736);
nor U2837 (N_2837,N_2722,N_2605);
and U2838 (N_2838,N_2642,N_2698);
and U2839 (N_2839,N_2770,N_2702);
nor U2840 (N_2840,N_2699,N_2660);
and U2841 (N_2841,N_2646,N_2676);
nor U2842 (N_2842,N_2789,N_2796);
nand U2843 (N_2843,N_2706,N_2694);
or U2844 (N_2844,N_2757,N_2747);
or U2845 (N_2845,N_2630,N_2769);
or U2846 (N_2846,N_2657,N_2622);
or U2847 (N_2847,N_2725,N_2633);
and U2848 (N_2848,N_2704,N_2777);
and U2849 (N_2849,N_2663,N_2655);
nor U2850 (N_2850,N_2715,N_2612);
and U2851 (N_2851,N_2689,N_2714);
nor U2852 (N_2852,N_2765,N_2701);
nand U2853 (N_2853,N_2771,N_2792);
and U2854 (N_2854,N_2650,N_2766);
or U2855 (N_2855,N_2798,N_2726);
and U2856 (N_2856,N_2753,N_2609);
nor U2857 (N_2857,N_2695,N_2783);
nor U2858 (N_2858,N_2615,N_2674);
and U2859 (N_2859,N_2719,N_2610);
or U2860 (N_2860,N_2607,N_2632);
nand U2861 (N_2861,N_2629,N_2785);
and U2862 (N_2862,N_2696,N_2682);
and U2863 (N_2863,N_2755,N_2667);
or U2864 (N_2864,N_2730,N_2627);
or U2865 (N_2865,N_2746,N_2751);
and U2866 (N_2866,N_2640,N_2631);
or U2867 (N_2867,N_2727,N_2638);
or U2868 (N_2868,N_2758,N_2772);
or U2869 (N_2869,N_2710,N_2623);
nand U2870 (N_2870,N_2705,N_2790);
or U2871 (N_2871,N_2795,N_2681);
nor U2872 (N_2872,N_2620,N_2760);
and U2873 (N_2873,N_2666,N_2762);
or U2874 (N_2874,N_2724,N_2764);
and U2875 (N_2875,N_2738,N_2648);
and U2876 (N_2876,N_2656,N_2729);
or U2877 (N_2877,N_2619,N_2644);
and U2878 (N_2878,N_2743,N_2779);
or U2879 (N_2879,N_2602,N_2740);
nor U2880 (N_2880,N_2685,N_2600);
or U2881 (N_2881,N_2691,N_2641);
nor U2882 (N_2882,N_2625,N_2707);
nand U2883 (N_2883,N_2745,N_2671);
nand U2884 (N_2884,N_2774,N_2677);
and U2885 (N_2885,N_2645,N_2752);
nor U2886 (N_2886,N_2635,N_2744);
xor U2887 (N_2887,N_2767,N_2653);
nor U2888 (N_2888,N_2680,N_2739);
nor U2889 (N_2889,N_2718,N_2742);
nor U2890 (N_2890,N_2697,N_2687);
and U2891 (N_2891,N_2768,N_2700);
nand U2892 (N_2892,N_2662,N_2651);
nand U2893 (N_2893,N_2716,N_2616);
nor U2894 (N_2894,N_2786,N_2773);
nand U2895 (N_2895,N_2686,N_2617);
nand U2896 (N_2896,N_2672,N_2781);
and U2897 (N_2897,N_2670,N_2634);
or U2898 (N_2898,N_2717,N_2787);
nor U2899 (N_2899,N_2608,N_2664);
nand U2900 (N_2900,N_2641,N_2785);
nand U2901 (N_2901,N_2774,N_2787);
nand U2902 (N_2902,N_2673,N_2664);
nor U2903 (N_2903,N_2670,N_2629);
nor U2904 (N_2904,N_2651,N_2653);
or U2905 (N_2905,N_2779,N_2719);
or U2906 (N_2906,N_2608,N_2662);
nand U2907 (N_2907,N_2688,N_2775);
nand U2908 (N_2908,N_2710,N_2767);
and U2909 (N_2909,N_2613,N_2663);
or U2910 (N_2910,N_2776,N_2711);
or U2911 (N_2911,N_2691,N_2782);
and U2912 (N_2912,N_2682,N_2760);
or U2913 (N_2913,N_2733,N_2795);
or U2914 (N_2914,N_2715,N_2692);
or U2915 (N_2915,N_2749,N_2671);
or U2916 (N_2916,N_2680,N_2691);
or U2917 (N_2917,N_2715,N_2663);
or U2918 (N_2918,N_2637,N_2730);
or U2919 (N_2919,N_2644,N_2744);
nor U2920 (N_2920,N_2620,N_2726);
and U2921 (N_2921,N_2659,N_2638);
and U2922 (N_2922,N_2747,N_2601);
or U2923 (N_2923,N_2669,N_2606);
nand U2924 (N_2924,N_2768,N_2776);
and U2925 (N_2925,N_2668,N_2613);
or U2926 (N_2926,N_2695,N_2651);
nor U2927 (N_2927,N_2673,N_2704);
nand U2928 (N_2928,N_2673,N_2768);
nor U2929 (N_2929,N_2605,N_2652);
or U2930 (N_2930,N_2643,N_2719);
or U2931 (N_2931,N_2706,N_2710);
and U2932 (N_2932,N_2649,N_2749);
and U2933 (N_2933,N_2788,N_2669);
and U2934 (N_2934,N_2689,N_2712);
nor U2935 (N_2935,N_2627,N_2659);
nand U2936 (N_2936,N_2688,N_2744);
and U2937 (N_2937,N_2748,N_2767);
and U2938 (N_2938,N_2778,N_2776);
nand U2939 (N_2939,N_2638,N_2766);
and U2940 (N_2940,N_2638,N_2720);
or U2941 (N_2941,N_2776,N_2649);
nand U2942 (N_2942,N_2732,N_2784);
and U2943 (N_2943,N_2740,N_2734);
or U2944 (N_2944,N_2673,N_2751);
nor U2945 (N_2945,N_2671,N_2634);
nor U2946 (N_2946,N_2698,N_2782);
nor U2947 (N_2947,N_2653,N_2684);
and U2948 (N_2948,N_2696,N_2643);
or U2949 (N_2949,N_2664,N_2633);
nor U2950 (N_2950,N_2793,N_2619);
and U2951 (N_2951,N_2632,N_2769);
nor U2952 (N_2952,N_2756,N_2669);
nor U2953 (N_2953,N_2665,N_2607);
or U2954 (N_2954,N_2690,N_2758);
nor U2955 (N_2955,N_2703,N_2740);
or U2956 (N_2956,N_2730,N_2756);
xor U2957 (N_2957,N_2634,N_2657);
and U2958 (N_2958,N_2756,N_2629);
nand U2959 (N_2959,N_2706,N_2648);
nand U2960 (N_2960,N_2768,N_2637);
and U2961 (N_2961,N_2679,N_2698);
nand U2962 (N_2962,N_2764,N_2608);
or U2963 (N_2963,N_2638,N_2680);
and U2964 (N_2964,N_2722,N_2693);
and U2965 (N_2965,N_2614,N_2639);
nor U2966 (N_2966,N_2631,N_2739);
and U2967 (N_2967,N_2624,N_2674);
and U2968 (N_2968,N_2668,N_2768);
nand U2969 (N_2969,N_2698,N_2759);
or U2970 (N_2970,N_2681,N_2759);
nand U2971 (N_2971,N_2718,N_2723);
nand U2972 (N_2972,N_2775,N_2640);
and U2973 (N_2973,N_2762,N_2722);
nand U2974 (N_2974,N_2650,N_2630);
nor U2975 (N_2975,N_2619,N_2704);
nor U2976 (N_2976,N_2680,N_2791);
and U2977 (N_2977,N_2753,N_2688);
nand U2978 (N_2978,N_2669,N_2740);
or U2979 (N_2979,N_2663,N_2781);
nor U2980 (N_2980,N_2765,N_2735);
and U2981 (N_2981,N_2694,N_2751);
nor U2982 (N_2982,N_2778,N_2631);
nor U2983 (N_2983,N_2661,N_2657);
and U2984 (N_2984,N_2651,N_2776);
or U2985 (N_2985,N_2735,N_2794);
and U2986 (N_2986,N_2608,N_2723);
nor U2987 (N_2987,N_2669,N_2751);
nand U2988 (N_2988,N_2790,N_2754);
and U2989 (N_2989,N_2702,N_2627);
and U2990 (N_2990,N_2723,N_2663);
nand U2991 (N_2991,N_2689,N_2693);
or U2992 (N_2992,N_2602,N_2635);
nor U2993 (N_2993,N_2736,N_2707);
nand U2994 (N_2994,N_2600,N_2635);
nor U2995 (N_2995,N_2620,N_2600);
nor U2996 (N_2996,N_2679,N_2706);
xor U2997 (N_2997,N_2691,N_2703);
or U2998 (N_2998,N_2794,N_2796);
or U2999 (N_2999,N_2614,N_2738);
and UO_0 (O_0,N_2842,N_2988);
nor UO_1 (O_1,N_2948,N_2981);
and UO_2 (O_2,N_2863,N_2921);
or UO_3 (O_3,N_2986,N_2915);
nor UO_4 (O_4,N_2928,N_2958);
nand UO_5 (O_5,N_2949,N_2972);
nand UO_6 (O_6,N_2936,N_2809);
or UO_7 (O_7,N_2849,N_2998);
or UO_8 (O_8,N_2860,N_2858);
nand UO_9 (O_9,N_2956,N_2957);
nor UO_10 (O_10,N_2942,N_2944);
or UO_11 (O_11,N_2910,N_2883);
or UO_12 (O_12,N_2843,N_2870);
nor UO_13 (O_13,N_2966,N_2806);
and UO_14 (O_14,N_2840,N_2821);
xor UO_15 (O_15,N_2969,N_2962);
and UO_16 (O_16,N_2879,N_2898);
nand UO_17 (O_17,N_2947,N_2827);
or UO_18 (O_18,N_2831,N_2976);
nand UO_19 (O_19,N_2970,N_2838);
and UO_20 (O_20,N_2923,N_2886);
nand UO_21 (O_21,N_2903,N_2920);
nand UO_22 (O_22,N_2866,N_2971);
nand UO_23 (O_23,N_2933,N_2989);
nand UO_24 (O_24,N_2867,N_2983);
nand UO_25 (O_25,N_2985,N_2816);
or UO_26 (O_26,N_2907,N_2808);
and UO_27 (O_27,N_2980,N_2908);
or UO_28 (O_28,N_2946,N_2984);
nor UO_29 (O_29,N_2803,N_2869);
nor UO_30 (O_30,N_2832,N_2825);
and UO_31 (O_31,N_2881,N_2927);
nor UO_32 (O_32,N_2995,N_2887);
nand UO_33 (O_33,N_2974,N_2990);
and UO_34 (O_34,N_2823,N_2819);
nor UO_35 (O_35,N_2895,N_2905);
nand UO_36 (O_36,N_2978,N_2929);
nand UO_37 (O_37,N_2902,N_2973);
or UO_38 (O_38,N_2826,N_2961);
nand UO_39 (O_39,N_2967,N_2951);
nor UO_40 (O_40,N_2937,N_2800);
nand UO_41 (O_41,N_2926,N_2913);
or UO_42 (O_42,N_2914,N_2837);
nand UO_43 (O_43,N_2943,N_2896);
or UO_44 (O_44,N_2959,N_2977);
or UO_45 (O_45,N_2934,N_2924);
and UO_46 (O_46,N_2954,N_2993);
nand UO_47 (O_47,N_2804,N_2939);
or UO_48 (O_48,N_2868,N_2857);
nor UO_49 (O_49,N_2996,N_2856);
and UO_50 (O_50,N_2829,N_2982);
nor UO_51 (O_51,N_2815,N_2952);
and UO_52 (O_52,N_2963,N_2814);
nor UO_53 (O_53,N_2906,N_2911);
nor UO_54 (O_54,N_2859,N_2953);
nand UO_55 (O_55,N_2925,N_2917);
and UO_56 (O_56,N_2964,N_2830);
and UO_57 (O_57,N_2885,N_2930);
nand UO_58 (O_58,N_2877,N_2817);
nor UO_59 (O_59,N_2992,N_2897);
and UO_60 (O_60,N_2892,N_2997);
nor UO_61 (O_61,N_2965,N_2848);
nand UO_62 (O_62,N_2802,N_2894);
nor UO_63 (O_63,N_2873,N_2852);
or UO_64 (O_64,N_2899,N_2880);
or UO_65 (O_65,N_2871,N_2882);
and UO_66 (O_66,N_2844,N_2813);
nor UO_67 (O_67,N_2812,N_2909);
nor UO_68 (O_68,N_2855,N_2900);
nor UO_69 (O_69,N_2841,N_2945);
nand UO_70 (O_70,N_2938,N_2834);
or UO_71 (O_71,N_2847,N_2893);
or UO_72 (O_72,N_2805,N_2884);
nor UO_73 (O_73,N_2822,N_2864);
nor UO_74 (O_74,N_2968,N_2820);
and UO_75 (O_75,N_2828,N_2904);
or UO_76 (O_76,N_2918,N_2960);
and UO_77 (O_77,N_2801,N_2874);
or UO_78 (O_78,N_2807,N_2850);
nor UO_79 (O_79,N_2811,N_2935);
and UO_80 (O_80,N_2916,N_2833);
and UO_81 (O_81,N_2861,N_2865);
nand UO_82 (O_82,N_2846,N_2999);
nand UO_83 (O_83,N_2975,N_2818);
and UO_84 (O_84,N_2891,N_2955);
nand UO_85 (O_85,N_2872,N_2890);
and UO_86 (O_86,N_2876,N_2888);
nand UO_87 (O_87,N_2875,N_2851);
and UO_88 (O_88,N_2950,N_2889);
nand UO_89 (O_89,N_2810,N_2835);
nor UO_90 (O_90,N_2931,N_2987);
nand UO_91 (O_91,N_2932,N_2901);
nor UO_92 (O_92,N_2854,N_2836);
and UO_93 (O_93,N_2912,N_2878);
or UO_94 (O_94,N_2824,N_2991);
and UO_95 (O_95,N_2862,N_2853);
nor UO_96 (O_96,N_2941,N_2839);
nor UO_97 (O_97,N_2922,N_2919);
nand UO_98 (O_98,N_2994,N_2845);
and UO_99 (O_99,N_2940,N_2979);
or UO_100 (O_100,N_2937,N_2825);
or UO_101 (O_101,N_2899,N_2991);
nor UO_102 (O_102,N_2972,N_2894);
and UO_103 (O_103,N_2970,N_2896);
nand UO_104 (O_104,N_2875,N_2959);
and UO_105 (O_105,N_2960,N_2887);
or UO_106 (O_106,N_2883,N_2949);
nand UO_107 (O_107,N_2940,N_2824);
nand UO_108 (O_108,N_2942,N_2812);
nor UO_109 (O_109,N_2870,N_2928);
and UO_110 (O_110,N_2848,N_2861);
nand UO_111 (O_111,N_2940,N_2952);
or UO_112 (O_112,N_2842,N_2997);
nand UO_113 (O_113,N_2914,N_2945);
nand UO_114 (O_114,N_2821,N_2870);
or UO_115 (O_115,N_2842,N_2883);
nand UO_116 (O_116,N_2916,N_2841);
or UO_117 (O_117,N_2846,N_2825);
and UO_118 (O_118,N_2936,N_2915);
and UO_119 (O_119,N_2983,N_2846);
or UO_120 (O_120,N_2813,N_2892);
and UO_121 (O_121,N_2980,N_2887);
or UO_122 (O_122,N_2948,N_2851);
nand UO_123 (O_123,N_2852,N_2932);
nand UO_124 (O_124,N_2981,N_2985);
nand UO_125 (O_125,N_2891,N_2849);
and UO_126 (O_126,N_2859,N_2990);
nand UO_127 (O_127,N_2915,N_2970);
nand UO_128 (O_128,N_2835,N_2883);
nor UO_129 (O_129,N_2838,N_2866);
nor UO_130 (O_130,N_2937,N_2917);
nor UO_131 (O_131,N_2808,N_2922);
or UO_132 (O_132,N_2878,N_2890);
nand UO_133 (O_133,N_2873,N_2817);
and UO_134 (O_134,N_2927,N_2873);
or UO_135 (O_135,N_2907,N_2842);
or UO_136 (O_136,N_2962,N_2994);
or UO_137 (O_137,N_2979,N_2844);
and UO_138 (O_138,N_2966,N_2922);
and UO_139 (O_139,N_2947,N_2874);
or UO_140 (O_140,N_2894,N_2940);
nor UO_141 (O_141,N_2882,N_2938);
nand UO_142 (O_142,N_2882,N_2915);
or UO_143 (O_143,N_2828,N_2834);
nand UO_144 (O_144,N_2958,N_2907);
nor UO_145 (O_145,N_2836,N_2815);
nand UO_146 (O_146,N_2908,N_2843);
nor UO_147 (O_147,N_2982,N_2889);
nor UO_148 (O_148,N_2941,N_2970);
nand UO_149 (O_149,N_2983,N_2862);
nor UO_150 (O_150,N_2987,N_2939);
nand UO_151 (O_151,N_2906,N_2926);
and UO_152 (O_152,N_2982,N_2823);
nor UO_153 (O_153,N_2975,N_2890);
nand UO_154 (O_154,N_2833,N_2868);
and UO_155 (O_155,N_2899,N_2916);
nand UO_156 (O_156,N_2898,N_2808);
or UO_157 (O_157,N_2900,N_2975);
or UO_158 (O_158,N_2846,N_2981);
or UO_159 (O_159,N_2952,N_2862);
or UO_160 (O_160,N_2837,N_2802);
and UO_161 (O_161,N_2807,N_2966);
and UO_162 (O_162,N_2937,N_2871);
and UO_163 (O_163,N_2827,N_2812);
or UO_164 (O_164,N_2892,N_2929);
or UO_165 (O_165,N_2889,N_2879);
nand UO_166 (O_166,N_2983,N_2945);
nor UO_167 (O_167,N_2923,N_2839);
or UO_168 (O_168,N_2952,N_2928);
nand UO_169 (O_169,N_2930,N_2817);
nand UO_170 (O_170,N_2801,N_2996);
nand UO_171 (O_171,N_2866,N_2874);
and UO_172 (O_172,N_2897,N_2808);
nor UO_173 (O_173,N_2926,N_2928);
and UO_174 (O_174,N_2932,N_2854);
or UO_175 (O_175,N_2898,N_2904);
nor UO_176 (O_176,N_2894,N_2884);
and UO_177 (O_177,N_2883,N_2907);
nor UO_178 (O_178,N_2847,N_2960);
or UO_179 (O_179,N_2950,N_2852);
nor UO_180 (O_180,N_2873,N_2980);
nand UO_181 (O_181,N_2865,N_2910);
nor UO_182 (O_182,N_2887,N_2872);
or UO_183 (O_183,N_2890,N_2829);
xnor UO_184 (O_184,N_2852,N_2900);
nand UO_185 (O_185,N_2915,N_2847);
and UO_186 (O_186,N_2962,N_2948);
nor UO_187 (O_187,N_2821,N_2810);
and UO_188 (O_188,N_2858,N_2995);
or UO_189 (O_189,N_2948,N_2893);
nand UO_190 (O_190,N_2864,N_2833);
nor UO_191 (O_191,N_2990,N_2964);
and UO_192 (O_192,N_2867,N_2973);
nand UO_193 (O_193,N_2953,N_2845);
and UO_194 (O_194,N_2827,N_2879);
or UO_195 (O_195,N_2923,N_2860);
nor UO_196 (O_196,N_2854,N_2833);
and UO_197 (O_197,N_2964,N_2884);
nor UO_198 (O_198,N_2888,N_2942);
nor UO_199 (O_199,N_2901,N_2948);
nand UO_200 (O_200,N_2911,N_2837);
or UO_201 (O_201,N_2979,N_2970);
nand UO_202 (O_202,N_2878,N_2962);
nor UO_203 (O_203,N_2960,N_2925);
xnor UO_204 (O_204,N_2900,N_2968);
and UO_205 (O_205,N_2878,N_2860);
or UO_206 (O_206,N_2836,N_2812);
and UO_207 (O_207,N_2950,N_2987);
nand UO_208 (O_208,N_2800,N_2838);
nand UO_209 (O_209,N_2929,N_2974);
or UO_210 (O_210,N_2977,N_2805);
nand UO_211 (O_211,N_2872,N_2844);
and UO_212 (O_212,N_2833,N_2837);
or UO_213 (O_213,N_2922,N_2906);
nor UO_214 (O_214,N_2892,N_2903);
or UO_215 (O_215,N_2878,N_2873);
and UO_216 (O_216,N_2849,N_2820);
or UO_217 (O_217,N_2943,N_2960);
or UO_218 (O_218,N_2817,N_2801);
and UO_219 (O_219,N_2827,N_2952);
nand UO_220 (O_220,N_2825,N_2998);
and UO_221 (O_221,N_2904,N_2894);
or UO_222 (O_222,N_2900,N_2874);
or UO_223 (O_223,N_2877,N_2911);
nor UO_224 (O_224,N_2968,N_2981);
and UO_225 (O_225,N_2908,N_2931);
nor UO_226 (O_226,N_2892,N_2832);
and UO_227 (O_227,N_2889,N_2813);
or UO_228 (O_228,N_2923,N_2903);
nor UO_229 (O_229,N_2825,N_2877);
and UO_230 (O_230,N_2935,N_2965);
nand UO_231 (O_231,N_2939,N_2889);
nand UO_232 (O_232,N_2973,N_2811);
and UO_233 (O_233,N_2953,N_2914);
or UO_234 (O_234,N_2857,N_2848);
nor UO_235 (O_235,N_2914,N_2920);
and UO_236 (O_236,N_2850,N_2983);
xor UO_237 (O_237,N_2999,N_2984);
and UO_238 (O_238,N_2848,N_2817);
nor UO_239 (O_239,N_2917,N_2953);
or UO_240 (O_240,N_2987,N_2824);
or UO_241 (O_241,N_2839,N_2881);
nor UO_242 (O_242,N_2845,N_2827);
or UO_243 (O_243,N_2874,N_2910);
and UO_244 (O_244,N_2996,N_2988);
or UO_245 (O_245,N_2857,N_2942);
or UO_246 (O_246,N_2827,N_2806);
nand UO_247 (O_247,N_2942,N_2865);
nand UO_248 (O_248,N_2920,N_2899);
nand UO_249 (O_249,N_2924,N_2819);
and UO_250 (O_250,N_2956,N_2960);
and UO_251 (O_251,N_2941,N_2836);
or UO_252 (O_252,N_2876,N_2853);
nor UO_253 (O_253,N_2811,N_2839);
and UO_254 (O_254,N_2980,N_2830);
nor UO_255 (O_255,N_2987,N_2968);
nand UO_256 (O_256,N_2812,N_2816);
nand UO_257 (O_257,N_2827,N_2841);
nand UO_258 (O_258,N_2927,N_2848);
or UO_259 (O_259,N_2876,N_2910);
or UO_260 (O_260,N_2859,N_2857);
nand UO_261 (O_261,N_2847,N_2881);
nand UO_262 (O_262,N_2930,N_2928);
or UO_263 (O_263,N_2995,N_2906);
nor UO_264 (O_264,N_2822,N_2857);
and UO_265 (O_265,N_2922,N_2874);
nand UO_266 (O_266,N_2882,N_2909);
or UO_267 (O_267,N_2857,N_2932);
or UO_268 (O_268,N_2842,N_2962);
nor UO_269 (O_269,N_2888,N_2868);
nand UO_270 (O_270,N_2843,N_2987);
and UO_271 (O_271,N_2916,N_2863);
nor UO_272 (O_272,N_2807,N_2808);
and UO_273 (O_273,N_2807,N_2945);
and UO_274 (O_274,N_2933,N_2855);
nor UO_275 (O_275,N_2819,N_2851);
nand UO_276 (O_276,N_2828,N_2984);
nand UO_277 (O_277,N_2918,N_2856);
or UO_278 (O_278,N_2985,N_2867);
nor UO_279 (O_279,N_2848,N_2993);
nand UO_280 (O_280,N_2807,N_2866);
nor UO_281 (O_281,N_2884,N_2864);
nor UO_282 (O_282,N_2954,N_2839);
nor UO_283 (O_283,N_2831,N_2917);
nor UO_284 (O_284,N_2908,N_2936);
nand UO_285 (O_285,N_2914,N_2882);
and UO_286 (O_286,N_2849,N_2902);
or UO_287 (O_287,N_2911,N_2961);
and UO_288 (O_288,N_2964,N_2856);
and UO_289 (O_289,N_2852,N_2938);
nor UO_290 (O_290,N_2961,N_2925);
nor UO_291 (O_291,N_2827,N_2908);
or UO_292 (O_292,N_2999,N_2934);
nand UO_293 (O_293,N_2827,N_2877);
and UO_294 (O_294,N_2855,N_2810);
nor UO_295 (O_295,N_2905,N_2818);
and UO_296 (O_296,N_2997,N_2955);
or UO_297 (O_297,N_2993,N_2802);
or UO_298 (O_298,N_2914,N_2984);
and UO_299 (O_299,N_2863,N_2869);
or UO_300 (O_300,N_2951,N_2870);
nand UO_301 (O_301,N_2938,N_2922);
nor UO_302 (O_302,N_2878,N_2844);
nand UO_303 (O_303,N_2815,N_2850);
nand UO_304 (O_304,N_2995,N_2951);
nor UO_305 (O_305,N_2840,N_2999);
and UO_306 (O_306,N_2823,N_2838);
nand UO_307 (O_307,N_2964,N_2888);
nand UO_308 (O_308,N_2854,N_2888);
nand UO_309 (O_309,N_2870,N_2828);
or UO_310 (O_310,N_2827,N_2824);
nor UO_311 (O_311,N_2972,N_2981);
nand UO_312 (O_312,N_2969,N_2863);
xor UO_313 (O_313,N_2865,N_2883);
nand UO_314 (O_314,N_2818,N_2833);
nand UO_315 (O_315,N_2827,N_2809);
and UO_316 (O_316,N_2894,N_2840);
nand UO_317 (O_317,N_2855,N_2958);
and UO_318 (O_318,N_2841,N_2964);
nand UO_319 (O_319,N_2934,N_2903);
nand UO_320 (O_320,N_2987,N_2937);
and UO_321 (O_321,N_2809,N_2826);
or UO_322 (O_322,N_2914,N_2902);
nand UO_323 (O_323,N_2897,N_2991);
nand UO_324 (O_324,N_2965,N_2883);
nor UO_325 (O_325,N_2847,N_2921);
nor UO_326 (O_326,N_2818,N_2853);
or UO_327 (O_327,N_2931,N_2915);
or UO_328 (O_328,N_2887,N_2949);
or UO_329 (O_329,N_2940,N_2810);
nor UO_330 (O_330,N_2895,N_2856);
nor UO_331 (O_331,N_2863,N_2923);
or UO_332 (O_332,N_2842,N_2873);
and UO_333 (O_333,N_2973,N_2856);
nand UO_334 (O_334,N_2805,N_2892);
nor UO_335 (O_335,N_2844,N_2851);
or UO_336 (O_336,N_2937,N_2851);
nand UO_337 (O_337,N_2802,N_2967);
nor UO_338 (O_338,N_2810,N_2953);
or UO_339 (O_339,N_2943,N_2880);
nand UO_340 (O_340,N_2954,N_2964);
and UO_341 (O_341,N_2978,N_2825);
and UO_342 (O_342,N_2969,N_2999);
nor UO_343 (O_343,N_2916,N_2882);
nor UO_344 (O_344,N_2886,N_2917);
nand UO_345 (O_345,N_2821,N_2879);
and UO_346 (O_346,N_2804,N_2940);
nand UO_347 (O_347,N_2959,N_2800);
nand UO_348 (O_348,N_2884,N_2898);
nor UO_349 (O_349,N_2987,N_2906);
nand UO_350 (O_350,N_2813,N_2828);
and UO_351 (O_351,N_2942,N_2844);
nor UO_352 (O_352,N_2849,N_2856);
or UO_353 (O_353,N_2986,N_2843);
nor UO_354 (O_354,N_2947,N_2881);
nor UO_355 (O_355,N_2828,N_2905);
and UO_356 (O_356,N_2825,N_2943);
or UO_357 (O_357,N_2883,N_2804);
or UO_358 (O_358,N_2856,N_2909);
nand UO_359 (O_359,N_2841,N_2956);
nand UO_360 (O_360,N_2919,N_2867);
or UO_361 (O_361,N_2919,N_2950);
and UO_362 (O_362,N_2974,N_2970);
nor UO_363 (O_363,N_2829,N_2949);
or UO_364 (O_364,N_2813,N_2827);
and UO_365 (O_365,N_2997,N_2945);
nand UO_366 (O_366,N_2857,N_2910);
nor UO_367 (O_367,N_2830,N_2829);
nor UO_368 (O_368,N_2812,N_2842);
and UO_369 (O_369,N_2953,N_2820);
or UO_370 (O_370,N_2953,N_2919);
nor UO_371 (O_371,N_2982,N_2890);
nand UO_372 (O_372,N_2988,N_2995);
or UO_373 (O_373,N_2893,N_2808);
nor UO_374 (O_374,N_2999,N_2898);
nor UO_375 (O_375,N_2893,N_2890);
nor UO_376 (O_376,N_2989,N_2904);
nand UO_377 (O_377,N_2861,N_2947);
or UO_378 (O_378,N_2830,N_2976);
and UO_379 (O_379,N_2877,N_2886);
xor UO_380 (O_380,N_2985,N_2945);
or UO_381 (O_381,N_2947,N_2851);
or UO_382 (O_382,N_2874,N_2992);
or UO_383 (O_383,N_2898,N_2801);
or UO_384 (O_384,N_2898,N_2825);
or UO_385 (O_385,N_2838,N_2966);
nand UO_386 (O_386,N_2810,N_2833);
or UO_387 (O_387,N_2800,N_2812);
nand UO_388 (O_388,N_2885,N_2923);
nor UO_389 (O_389,N_2915,N_2867);
or UO_390 (O_390,N_2863,N_2854);
or UO_391 (O_391,N_2850,N_2829);
nand UO_392 (O_392,N_2884,N_2827);
and UO_393 (O_393,N_2913,N_2909);
nor UO_394 (O_394,N_2901,N_2907);
and UO_395 (O_395,N_2892,N_2822);
nand UO_396 (O_396,N_2922,N_2860);
nor UO_397 (O_397,N_2959,N_2931);
or UO_398 (O_398,N_2837,N_2897);
nand UO_399 (O_399,N_2903,N_2993);
or UO_400 (O_400,N_2804,N_2890);
and UO_401 (O_401,N_2864,N_2910);
or UO_402 (O_402,N_2800,N_2826);
or UO_403 (O_403,N_2935,N_2936);
nand UO_404 (O_404,N_2959,N_2929);
and UO_405 (O_405,N_2949,N_2872);
or UO_406 (O_406,N_2825,N_2985);
and UO_407 (O_407,N_2851,N_2878);
xnor UO_408 (O_408,N_2974,N_2870);
nor UO_409 (O_409,N_2863,N_2880);
nand UO_410 (O_410,N_2976,N_2809);
nand UO_411 (O_411,N_2834,N_2973);
nand UO_412 (O_412,N_2801,N_2859);
nand UO_413 (O_413,N_2949,N_2964);
nand UO_414 (O_414,N_2826,N_2900);
nand UO_415 (O_415,N_2846,N_2907);
nand UO_416 (O_416,N_2918,N_2975);
nor UO_417 (O_417,N_2985,N_2888);
nor UO_418 (O_418,N_2935,N_2987);
and UO_419 (O_419,N_2957,N_2990);
nand UO_420 (O_420,N_2825,N_2823);
and UO_421 (O_421,N_2939,N_2861);
or UO_422 (O_422,N_2808,N_2987);
nand UO_423 (O_423,N_2905,N_2966);
nor UO_424 (O_424,N_2908,N_2905);
and UO_425 (O_425,N_2821,N_2977);
or UO_426 (O_426,N_2896,N_2859);
and UO_427 (O_427,N_2832,N_2991);
or UO_428 (O_428,N_2984,N_2934);
and UO_429 (O_429,N_2863,N_2913);
nor UO_430 (O_430,N_2955,N_2817);
nand UO_431 (O_431,N_2829,N_2869);
nor UO_432 (O_432,N_2842,N_2845);
and UO_433 (O_433,N_2845,N_2802);
nand UO_434 (O_434,N_2917,N_2918);
or UO_435 (O_435,N_2981,N_2936);
nand UO_436 (O_436,N_2922,N_2803);
and UO_437 (O_437,N_2844,N_2801);
and UO_438 (O_438,N_2813,N_2878);
or UO_439 (O_439,N_2805,N_2898);
nand UO_440 (O_440,N_2816,N_2840);
or UO_441 (O_441,N_2963,N_2822);
and UO_442 (O_442,N_2962,N_2952);
or UO_443 (O_443,N_2958,N_2988);
nand UO_444 (O_444,N_2889,N_2956);
nand UO_445 (O_445,N_2986,N_2803);
nand UO_446 (O_446,N_2991,N_2952);
and UO_447 (O_447,N_2843,N_2873);
or UO_448 (O_448,N_2891,N_2811);
or UO_449 (O_449,N_2894,N_2842);
and UO_450 (O_450,N_2918,N_2876);
nand UO_451 (O_451,N_2943,N_2863);
and UO_452 (O_452,N_2982,N_2944);
nand UO_453 (O_453,N_2814,N_2834);
nor UO_454 (O_454,N_2909,N_2965);
and UO_455 (O_455,N_2898,N_2905);
or UO_456 (O_456,N_2942,N_2935);
nand UO_457 (O_457,N_2876,N_2817);
or UO_458 (O_458,N_2884,N_2886);
and UO_459 (O_459,N_2897,N_2928);
nor UO_460 (O_460,N_2824,N_2932);
or UO_461 (O_461,N_2989,N_2980);
or UO_462 (O_462,N_2950,N_2880);
or UO_463 (O_463,N_2809,N_2859);
and UO_464 (O_464,N_2906,N_2901);
and UO_465 (O_465,N_2891,N_2911);
nand UO_466 (O_466,N_2903,N_2998);
nor UO_467 (O_467,N_2857,N_2852);
nor UO_468 (O_468,N_2953,N_2857);
and UO_469 (O_469,N_2959,N_2817);
or UO_470 (O_470,N_2920,N_2882);
or UO_471 (O_471,N_2867,N_2949);
nand UO_472 (O_472,N_2933,N_2927);
and UO_473 (O_473,N_2826,N_2895);
nand UO_474 (O_474,N_2861,N_2824);
and UO_475 (O_475,N_2895,N_2865);
nand UO_476 (O_476,N_2813,N_2845);
nand UO_477 (O_477,N_2930,N_2874);
nand UO_478 (O_478,N_2970,N_2950);
and UO_479 (O_479,N_2873,N_2805);
nor UO_480 (O_480,N_2955,N_2946);
or UO_481 (O_481,N_2833,N_2989);
nand UO_482 (O_482,N_2812,N_2864);
nand UO_483 (O_483,N_2825,N_2892);
nand UO_484 (O_484,N_2963,N_2866);
and UO_485 (O_485,N_2825,N_2850);
or UO_486 (O_486,N_2869,N_2819);
nor UO_487 (O_487,N_2933,N_2813);
nor UO_488 (O_488,N_2989,N_2944);
or UO_489 (O_489,N_2864,N_2859);
nor UO_490 (O_490,N_2814,N_2857);
and UO_491 (O_491,N_2989,N_2912);
or UO_492 (O_492,N_2913,N_2897);
or UO_493 (O_493,N_2959,N_2803);
or UO_494 (O_494,N_2963,N_2982);
or UO_495 (O_495,N_2928,N_2927);
or UO_496 (O_496,N_2912,N_2865);
or UO_497 (O_497,N_2906,N_2930);
nor UO_498 (O_498,N_2926,N_2947);
or UO_499 (O_499,N_2820,N_2966);
endmodule