module basic_1500_15000_2000_10_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_428,In_26);
xnor U1 (N_1,In_1030,In_1037);
nand U2 (N_2,In_745,In_988);
and U3 (N_3,In_122,In_959);
or U4 (N_4,In_429,In_1467);
and U5 (N_5,In_362,In_928);
and U6 (N_6,In_767,In_1209);
nand U7 (N_7,In_222,In_1066);
xnor U8 (N_8,In_1052,In_72);
nor U9 (N_9,In_1130,In_843);
nand U10 (N_10,In_366,In_1286);
or U11 (N_11,In_391,In_1299);
or U12 (N_12,In_215,In_1447);
and U13 (N_13,In_639,In_941);
nand U14 (N_14,In_858,In_191);
nor U15 (N_15,In_857,In_560);
nand U16 (N_16,In_906,In_138);
xnor U17 (N_17,In_165,In_544);
or U18 (N_18,In_826,In_650);
nand U19 (N_19,In_1256,In_19);
nand U20 (N_20,In_266,In_1494);
or U21 (N_21,In_438,In_606);
xnor U22 (N_22,In_822,In_267);
nor U23 (N_23,In_351,In_404);
nand U24 (N_24,In_761,In_164);
or U25 (N_25,In_442,In_1336);
nor U26 (N_26,In_1108,In_622);
or U27 (N_27,In_672,In_981);
nor U28 (N_28,In_798,In_61);
or U29 (N_29,In_794,In_514);
xor U30 (N_30,In_640,In_345);
and U31 (N_31,In_596,In_756);
and U32 (N_32,In_809,In_851);
and U33 (N_33,In_616,In_179);
or U34 (N_34,In_28,In_239);
nor U35 (N_35,In_1045,In_293);
and U36 (N_36,In_445,In_291);
or U37 (N_37,In_1344,In_4);
or U38 (N_38,In_8,In_854);
or U39 (N_39,In_464,In_1451);
xor U40 (N_40,In_970,In_577);
and U41 (N_41,In_1269,In_1355);
and U42 (N_42,In_168,In_286);
or U43 (N_43,In_787,In_1144);
or U44 (N_44,In_855,In_1207);
or U45 (N_45,In_754,In_1409);
nand U46 (N_46,In_212,In_55);
xnor U47 (N_47,In_17,In_475);
nand U48 (N_48,In_1487,In_227);
xor U49 (N_49,In_872,In_1078);
or U50 (N_50,In_1230,In_1035);
or U51 (N_51,In_1290,In_1339);
xor U52 (N_52,In_354,In_1154);
or U53 (N_53,In_1488,In_1081);
nand U54 (N_54,In_434,In_943);
nor U55 (N_55,In_541,In_1410);
or U56 (N_56,In_1386,In_820);
nor U57 (N_57,In_340,In_387);
and U58 (N_58,In_1322,In_1497);
and U59 (N_59,In_1429,In_611);
or U60 (N_60,In_935,In_671);
and U61 (N_61,In_125,In_1004);
and U62 (N_62,In_751,In_727);
and U63 (N_63,In_600,In_282);
nor U64 (N_64,In_627,In_1448);
nor U65 (N_65,In_556,In_1117);
nand U66 (N_66,In_88,In_372);
xnor U67 (N_67,In_1316,In_54);
nor U68 (N_68,In_251,In_807);
or U69 (N_69,In_41,In_626);
xor U70 (N_70,In_1060,In_695);
nand U71 (N_71,In_1319,In_137);
nand U72 (N_72,In_95,In_1405);
nand U73 (N_73,In_50,In_355);
xor U74 (N_74,In_476,In_1398);
xor U75 (N_75,In_849,In_702);
or U76 (N_76,In_1164,In_489);
nand U77 (N_77,In_1153,In_1026);
or U78 (N_78,In_927,In_205);
and U79 (N_79,In_269,In_642);
and U80 (N_80,In_457,In_264);
nor U81 (N_81,In_97,In_9);
and U82 (N_82,In_1080,In_1271);
nor U83 (N_83,In_121,In_1303);
xor U84 (N_84,In_410,In_583);
nor U85 (N_85,In_505,In_1359);
nor U86 (N_86,In_1137,In_1238);
and U87 (N_87,In_675,In_1456);
xnor U88 (N_88,In_896,In_590);
nand U89 (N_89,In_1222,In_460);
nor U90 (N_90,In_631,In_484);
xnor U91 (N_91,In_522,In_224);
xnor U92 (N_92,In_257,In_1219);
xnor U93 (N_93,In_552,In_1250);
nor U94 (N_94,In_220,In_237);
nor U95 (N_95,In_1289,In_833);
nand U96 (N_96,In_539,In_525);
nand U97 (N_97,In_922,In_791);
nor U98 (N_98,In_677,In_120);
and U99 (N_99,In_1146,In_29);
or U100 (N_100,In_1466,In_130);
and U101 (N_101,In_1446,In_1454);
or U102 (N_102,In_380,In_868);
nor U103 (N_103,In_1380,In_46);
nor U104 (N_104,In_945,In_548);
nand U105 (N_105,In_1313,In_306);
xnor U106 (N_106,In_1426,In_501);
or U107 (N_107,In_808,In_1321);
nor U108 (N_108,In_836,In_1485);
nor U109 (N_109,In_1318,In_870);
or U110 (N_110,In_721,In_737);
nand U111 (N_111,In_0,In_1183);
nand U112 (N_112,In_646,In_343);
or U113 (N_113,In_1277,In_443);
nor U114 (N_114,In_914,In_993);
xor U115 (N_115,In_1096,In_243);
and U116 (N_116,In_1295,In_85);
and U117 (N_117,In_507,In_1275);
xor U118 (N_118,In_952,In_705);
xnor U119 (N_119,In_571,In_153);
nor U120 (N_120,In_1082,In_834);
xor U121 (N_121,In_465,In_1388);
xnor U122 (N_122,In_272,In_845);
nor U123 (N_123,In_1261,In_816);
nand U124 (N_124,In_995,In_270);
nand U125 (N_125,In_180,In_304);
nor U126 (N_126,In_1053,In_1079);
or U127 (N_127,In_316,In_889);
or U128 (N_128,In_666,In_888);
nand U129 (N_129,In_1370,In_608);
nand U130 (N_130,In_1057,In_759);
nand U131 (N_131,In_667,In_789);
and U132 (N_132,In_815,In_618);
xor U133 (N_133,In_1330,In_158);
or U134 (N_134,In_1367,In_924);
nand U135 (N_135,In_149,In_1465);
and U136 (N_136,In_1036,In_312);
and U137 (N_137,In_772,In_714);
nor U138 (N_138,In_152,In_1092);
nor U139 (N_139,In_1283,In_1457);
xnor U140 (N_140,In_925,In_1481);
nor U141 (N_141,In_1043,In_542);
and U142 (N_142,In_1323,In_73);
nor U143 (N_143,In_207,In_1157);
and U144 (N_144,In_1297,In_853);
and U145 (N_145,In_632,In_1291);
xor U146 (N_146,In_591,In_910);
nand U147 (N_147,In_575,In_271);
nand U148 (N_148,In_169,In_938);
or U149 (N_149,In_568,In_102);
xnor U150 (N_150,In_1018,In_486);
nor U151 (N_151,In_334,In_133);
nor U152 (N_152,In_16,In_711);
or U153 (N_153,In_1101,In_1471);
nand U154 (N_154,In_1002,In_746);
or U155 (N_155,In_792,In_592);
xor U156 (N_156,In_109,In_1384);
and U157 (N_157,In_1039,In_161);
and U158 (N_158,In_1416,In_975);
or U159 (N_159,In_339,In_688);
nor U160 (N_160,In_131,In_1302);
xor U161 (N_161,In_374,In_942);
or U162 (N_162,In_520,In_1421);
nand U163 (N_163,In_308,In_1047);
and U164 (N_164,In_708,In_90);
and U165 (N_165,In_613,In_936);
and U166 (N_166,In_838,In_232);
and U167 (N_167,In_314,In_821);
nor U168 (N_168,In_796,In_1423);
or U169 (N_169,In_297,In_1362);
or U170 (N_170,In_115,In_456);
xnor U171 (N_171,In_1473,In_684);
and U172 (N_172,In_288,In_368);
or U173 (N_173,In_1309,In_1202);
nor U174 (N_174,In_1048,In_722);
or U175 (N_175,In_1265,In_1213);
nor U176 (N_176,In_1008,In_225);
or U177 (N_177,In_1203,In_1194);
nand U178 (N_178,In_1055,In_416);
nand U179 (N_179,In_1218,In_444);
or U180 (N_180,In_965,In_1169);
and U181 (N_181,In_1149,In_256);
nand U182 (N_182,In_884,In_1034);
nor U183 (N_183,In_1105,In_69);
nor U184 (N_184,In_344,In_142);
and U185 (N_185,In_946,In_806);
xor U186 (N_186,In_863,In_1244);
nand U187 (N_187,In_189,In_1170);
and U188 (N_188,In_1143,In_253);
or U189 (N_189,In_1050,In_1412);
nand U190 (N_190,In_283,In_804);
xnor U191 (N_191,In_811,In_861);
nor U192 (N_192,In_1148,In_1484);
nor U193 (N_193,In_181,In_1326);
nor U194 (N_194,In_837,In_116);
nand U195 (N_195,In_766,In_782);
and U196 (N_196,In_1252,In_147);
xnor U197 (N_197,In_1356,In_567);
xnor U198 (N_198,In_1311,In_1434);
or U199 (N_199,In_1347,In_87);
nand U200 (N_200,In_96,In_537);
xnor U201 (N_201,In_209,In_315);
nor U202 (N_202,In_479,In_1425);
or U203 (N_203,In_917,In_176);
nor U204 (N_204,In_1178,In_1254);
or U205 (N_205,In_1097,In_883);
nand U206 (N_206,In_483,In_94);
nand U207 (N_207,In_1072,In_1064);
and U208 (N_208,In_163,In_657);
xor U209 (N_209,In_157,In_1025);
nand U210 (N_210,In_1001,In_154);
xor U211 (N_211,In_648,In_1490);
nand U212 (N_212,In_686,In_1159);
or U213 (N_213,In_1099,In_342);
xnor U214 (N_214,In_1285,In_1021);
and U215 (N_215,In_565,In_185);
xnor U216 (N_216,In_907,In_1100);
nand U217 (N_217,In_1006,In_871);
nor U218 (N_218,In_747,In_403);
and U219 (N_219,In_1427,In_134);
xor U220 (N_220,In_958,In_1468);
nand U221 (N_221,In_1185,In_1401);
nor U222 (N_222,In_1433,In_1011);
nor U223 (N_223,In_738,In_182);
xor U224 (N_224,In_586,In_835);
nor U225 (N_225,In_503,In_370);
nand U226 (N_226,In_1361,In_1126);
nand U227 (N_227,In_126,In_247);
and U228 (N_228,In_985,In_1246);
or U229 (N_229,In_1436,In_614);
nand U230 (N_230,In_71,In_890);
xor U231 (N_231,In_118,In_188);
nor U232 (N_232,In_1288,In_84);
nor U233 (N_233,In_956,In_661);
and U234 (N_234,In_459,In_244);
nand U235 (N_235,In_1061,In_7);
xnor U236 (N_236,In_1404,In_1113);
or U237 (N_237,In_1206,In_867);
and U238 (N_238,In_1327,In_660);
and U239 (N_239,In_1414,In_976);
nand U240 (N_240,In_972,In_690);
nor U241 (N_241,In_1226,In_1287);
and U242 (N_242,In_211,In_1116);
nand U243 (N_243,In_712,In_322);
and U244 (N_244,In_670,In_1134);
and U245 (N_245,In_319,In_107);
xnor U246 (N_246,In_1478,In_1158);
xor U247 (N_247,In_1237,In_1095);
nand U248 (N_248,In_700,In_1348);
xnor U249 (N_249,In_18,In_1279);
nor U250 (N_250,In_148,In_612);
nand U251 (N_251,In_653,In_1138);
xnor U252 (N_252,In_1332,In_234);
and U253 (N_253,In_703,In_1071);
nor U254 (N_254,In_681,In_966);
or U255 (N_255,In_758,In_1027);
nand U256 (N_256,In_1231,In_418);
and U257 (N_257,In_1142,In_453);
nor U258 (N_258,In_1073,In_621);
and U259 (N_259,In_974,In_1306);
xor U260 (N_260,In_783,In_1443);
nor U261 (N_261,In_1266,In_21);
nor U262 (N_262,In_630,In_146);
and U263 (N_263,In_129,In_452);
nand U264 (N_264,In_659,In_1349);
nand U265 (N_265,In_114,In_760);
and U266 (N_266,In_335,In_338);
nor U267 (N_267,In_1442,In_229);
nor U268 (N_268,In_573,In_35);
nor U269 (N_269,In_1151,In_799);
nor U270 (N_270,In_433,In_423);
or U271 (N_271,In_619,In_228);
and U272 (N_272,In_101,In_27);
nor U273 (N_273,In_170,In_276);
nand U274 (N_274,In_356,In_183);
and U275 (N_275,In_67,In_647);
and U276 (N_276,In_1475,In_1314);
xor U277 (N_277,In_104,In_823);
and U278 (N_278,In_1119,In_358);
nor U279 (N_279,In_674,In_519);
and U280 (N_280,In_446,In_382);
and U281 (N_281,In_512,In_1184);
nand U282 (N_282,In_500,In_866);
xnor U283 (N_283,In_1028,In_202);
nor U284 (N_284,In_1051,In_1007);
and U285 (N_285,In_1086,In_255);
or U286 (N_286,In_1,In_401);
nand U287 (N_287,In_879,In_719);
or U288 (N_288,In_878,In_1109);
or U289 (N_289,In_1450,In_414);
or U290 (N_290,In_634,In_1139);
or U291 (N_291,In_47,In_1310);
nand U292 (N_292,In_1233,In_645);
or U293 (N_293,In_814,In_296);
nor U294 (N_294,In_683,In_40);
or U295 (N_295,In_658,In_625);
xnor U296 (N_296,In_1341,In_388);
nor U297 (N_297,In_1013,In_623);
and U298 (N_298,In_1373,In_848);
or U299 (N_299,In_390,In_605);
xnor U300 (N_300,In_1147,In_1088);
nand U301 (N_301,In_939,In_49);
xnor U302 (N_302,In_880,In_1223);
or U303 (N_303,In_376,In_466);
xor U304 (N_304,In_1249,In_558);
and U305 (N_305,In_369,In_847);
nor U306 (N_306,In_499,In_698);
nor U307 (N_307,In_1338,In_1198);
or U308 (N_308,In_184,In_844);
or U309 (N_309,In_160,In_1489);
nand U310 (N_310,In_770,In_1400);
and U311 (N_311,In_1133,In_1128);
xor U312 (N_312,In_470,In_513);
or U313 (N_313,In_1188,In_68);
nor U314 (N_314,In_805,In_1225);
nor U315 (N_315,In_1365,In_908);
or U316 (N_316,In_492,In_1385);
or U317 (N_317,In_1014,In_381);
nand U318 (N_318,In_864,In_34);
xnor U319 (N_319,In_1351,In_216);
and U320 (N_320,In_36,In_1483);
xor U321 (N_321,In_1167,In_143);
nor U322 (N_322,In_1363,In_1089);
nor U323 (N_323,In_1123,In_641);
xnor U324 (N_324,In_827,In_1301);
xnor U325 (N_325,In_655,In_912);
xor U326 (N_326,In_321,In_915);
nor U327 (N_327,In_669,In_526);
or U328 (N_328,In_1360,In_1476);
and U329 (N_329,In_564,In_607);
xnor U330 (N_330,In_693,In_206);
and U331 (N_331,In_1017,In_258);
nor U332 (N_332,In_458,In_236);
nor U333 (N_333,In_1160,In_285);
or U334 (N_334,In_123,In_764);
xor U335 (N_335,In_37,In_620);
nand U336 (N_336,In_1276,In_287);
nand U337 (N_337,In_529,In_733);
and U338 (N_338,In_1415,In_1091);
or U339 (N_339,In_1189,In_451);
and U340 (N_340,In_1190,In_64);
and U341 (N_341,In_740,In_579);
nand U342 (N_342,In_420,In_396);
nor U343 (N_343,In_441,In_59);
xor U344 (N_344,In_1217,In_74);
xnor U345 (N_345,In_327,In_469);
nand U346 (N_346,In_1371,In_145);
or U347 (N_347,In_60,In_472);
or U348 (N_348,In_80,In_682);
nor U349 (N_349,In_455,In_1215);
nor U350 (N_350,In_547,In_533);
and U351 (N_351,In_1156,In_395);
nand U352 (N_352,In_99,In_856);
or U353 (N_353,In_569,In_1245);
nor U354 (N_354,In_1182,In_361);
nand U355 (N_355,In_832,In_259);
nor U356 (N_356,In_629,In_110);
xnor U357 (N_357,In_869,In_748);
nor U358 (N_358,In_409,In_117);
xor U359 (N_359,In_1077,In_106);
and U360 (N_360,In_144,In_481);
xnor U361 (N_361,In_1369,In_437);
nor U362 (N_362,In_1281,In_730);
nor U363 (N_363,In_940,In_128);
nor U364 (N_364,In_706,In_1232);
and U365 (N_365,In_819,In_1255);
nor U366 (N_366,In_986,In_151);
nor U367 (N_367,In_491,In_33);
or U368 (N_368,In_502,In_707);
nand U369 (N_369,In_790,In_1391);
xor U370 (N_370,In_709,In_400);
or U371 (N_371,In_589,In_894);
xor U372 (N_372,In_566,In_635);
nand U373 (N_373,In_12,In_633);
nand U374 (N_374,In_495,In_20);
nand U375 (N_375,In_732,In_1304);
nand U376 (N_376,In_493,In_48);
nor U377 (N_377,In_349,In_1059);
xnor U378 (N_378,In_1305,In_167);
nor U379 (N_379,In_1431,In_1235);
nand U380 (N_380,In_219,In_417);
or U381 (N_381,In_885,In_75);
or U382 (N_382,In_517,In_478);
xnor U383 (N_383,In_379,In_824);
or U384 (N_384,In_331,In_425);
xor U385 (N_385,In_1062,In_213);
xnor U386 (N_386,In_1176,In_3);
or U387 (N_387,In_994,In_462);
nor U388 (N_388,In_411,In_1343);
nand U389 (N_389,In_393,In_535);
and U390 (N_390,In_1441,In_1162);
and U391 (N_391,In_628,In_454);
nand U392 (N_392,In_1397,In_802);
nand U393 (N_393,In_1383,In_421);
and U394 (N_394,In_250,In_779);
and U395 (N_395,In_341,In_1406);
and U396 (N_396,In_1140,In_1111);
nand U397 (N_397,In_743,In_662);
xor U398 (N_398,In_178,In_685);
and U399 (N_399,In_1382,In_431);
nor U400 (N_400,In_773,In_1272);
or U401 (N_401,In_201,In_598);
nor U402 (N_402,In_1324,In_412);
nand U403 (N_403,In_728,In_637);
or U404 (N_404,In_221,In_1440);
nor U405 (N_405,In_930,In_1122);
nand U406 (N_406,In_768,In_960);
nand U407 (N_407,In_1296,In_999);
or U408 (N_408,In_1392,In_1381);
xnor U409 (N_409,In_447,In_638);
nor U410 (N_410,In_303,In_691);
nor U411 (N_411,In_177,In_531);
and U412 (N_412,In_1396,In_1469);
nand U413 (N_413,In_696,In_617);
or U414 (N_414,In_367,In_310);
xnor U415 (N_415,In_62,In_1201);
xor U416 (N_416,In_595,In_1093);
nor U417 (N_417,In_1307,In_1461);
xnor U418 (N_418,In_755,In_488);
or U419 (N_419,In_839,In_172);
or U420 (N_420,In_254,In_136);
nand U421 (N_421,In_496,In_1449);
nand U422 (N_422,In_150,In_53);
or U423 (N_423,In_31,In_1046);
nor U424 (N_424,In_916,In_725);
xor U425 (N_425,In_1248,In_311);
and U426 (N_426,In_1419,In_800);
xor U427 (N_427,In_903,In_511);
nand U428 (N_428,In_402,In_1438);
and U429 (N_429,In_676,In_93);
or U430 (N_430,In_195,In_1023);
or U431 (N_431,In_874,In_1395);
and U432 (N_432,In_920,In_1264);
nand U433 (N_433,In_235,In_597);
nor U434 (N_434,In_1110,In_828);
and U435 (N_435,In_487,In_1204);
xor U436 (N_436,In_1236,In_801);
and U437 (N_437,In_162,In_1458);
nor U438 (N_438,In_1177,In_570);
nand U439 (N_439,In_694,In_1181);
nand U440 (N_440,In_375,In_1453);
and U441 (N_441,In_204,In_249);
nand U442 (N_442,In_947,In_25);
xnor U443 (N_443,In_1049,In_1056);
or U444 (N_444,In_1486,In_1376);
and U445 (N_445,In_260,In_1357);
nand U446 (N_446,In_860,In_1462);
or U447 (N_447,In_1090,In_226);
xor U448 (N_448,In_983,In_1267);
xnor U449 (N_449,In_105,In_357);
nand U450 (N_450,In_371,In_1003);
and U451 (N_451,In_298,In_127);
xnor U452 (N_452,In_724,In_174);
or U453 (N_453,In_406,In_534);
and U454 (N_454,In_1477,In_913);
xnor U455 (N_455,In_951,In_1352);
xor U456 (N_456,In_1127,In_63);
or U457 (N_457,In_987,In_902);
or U458 (N_458,In_1432,In_919);
or U459 (N_459,In_899,In_1372);
and U460 (N_460,In_692,In_1328);
nor U461 (N_461,In_576,In_262);
xnor U462 (N_462,In_92,In_1174);
or U463 (N_463,In_978,In_527);
or U464 (N_464,In_261,In_1179);
nor U465 (N_465,In_1358,In_777);
or U466 (N_466,In_1260,In_599);
or U467 (N_467,In_578,In_448);
nand U468 (N_468,In_273,In_24);
nor U469 (N_469,In_1019,In_1455);
or U470 (N_470,In_1076,In_399);
nor U471 (N_471,In_450,In_233);
nor U472 (N_472,In_223,In_731);
nor U473 (N_473,In_294,In_984);
nand U474 (N_474,In_1041,In_1075);
or U475 (N_475,In_318,In_1196);
nor U476 (N_476,In_38,In_1479);
nand U477 (N_477,In_803,In_726);
and U478 (N_478,In_968,In_1408);
or U479 (N_479,In_1242,In_574);
xor U480 (N_480,In_697,In_1439);
nor U481 (N_481,In_739,In_540);
nor U482 (N_482,In_1038,In_715);
or U483 (N_483,In_1239,In_1069);
xor U484 (N_484,In_408,In_463);
nor U485 (N_485,In_818,In_347);
nand U486 (N_486,In_435,In_196);
nor U487 (N_487,In_430,In_780);
nor U488 (N_488,In_1054,In_957);
nand U489 (N_489,In_736,In_680);
nor U490 (N_490,In_769,In_506);
nor U491 (N_491,In_1437,In_352);
or U492 (N_492,In_1350,In_841);
nor U493 (N_493,In_208,In_649);
or U494 (N_494,In_654,In_39);
nor U495 (N_495,In_86,In_461);
and U496 (N_496,In_893,In_320);
nor U497 (N_497,In_328,In_246);
nand U498 (N_498,In_82,In_643);
or U499 (N_499,In_1166,In_1084);
or U500 (N_500,In_1087,In_830);
xor U501 (N_501,In_664,In_330);
xor U502 (N_502,In_1379,In_1197);
xnor U503 (N_503,In_407,In_426);
xor U504 (N_504,In_1042,In_929);
nor U505 (N_505,In_842,In_384);
nand U506 (N_506,In_1474,In_1375);
and U507 (N_507,In_509,In_603);
or U508 (N_508,In_278,In_744);
or U509 (N_509,In_268,In_651);
nor U510 (N_510,In_1459,In_141);
nor U511 (N_511,In_497,In_909);
xnor U512 (N_512,In_1083,In_1234);
xnor U513 (N_513,In_840,In_346);
or U514 (N_514,In_543,In_504);
nand U515 (N_515,In_582,In_741);
xor U516 (N_516,In_385,In_515);
or U517 (N_517,In_111,In_325);
nor U518 (N_518,In_963,In_873);
and U519 (N_519,In_786,In_333);
nand U520 (N_520,In_81,In_1435);
or U521 (N_521,In_13,In_1152);
nor U522 (N_522,In_1107,In_1320);
nand U523 (N_523,In_610,In_1165);
nand U524 (N_524,In_898,In_1470);
and U525 (N_525,In_1221,In_1121);
xor U526 (N_526,In_1227,In_1102);
xnor U527 (N_527,In_79,In_490);
nand U528 (N_528,In_581,In_1329);
xnor U529 (N_529,In_217,In_781);
nand U530 (N_530,In_594,In_301);
or U531 (N_531,In_1141,In_187);
nand U532 (N_532,In_365,In_895);
nor U533 (N_533,In_336,In_440);
xnor U534 (N_534,In_1012,In_580);
xnor U535 (N_535,In_1390,In_1132);
xnor U536 (N_536,In_1262,In_359);
nand U537 (N_537,In_1333,In_1106);
nand U538 (N_538,In_1498,In_887);
nand U539 (N_539,In_471,In_1491);
xor U540 (N_540,In_585,In_1192);
and U541 (N_541,In_831,In_723);
or U542 (N_542,In_1292,In_882);
or U543 (N_543,In_601,In_1407);
nand U544 (N_544,In_265,In_1029);
and U545 (N_545,In_295,In_241);
nor U546 (N_546,In_1496,In_485);
xor U547 (N_547,In_139,In_494);
or U548 (N_548,In_198,In_200);
xor U549 (N_549,In_1005,In_765);
and U550 (N_550,In_113,In_348);
xor U551 (N_551,In_238,In_977);
and U552 (N_552,In_1331,In_186);
xnor U553 (N_553,In_10,In_91);
xor U554 (N_554,In_735,In_317);
xnor U555 (N_555,In_193,In_1070);
or U556 (N_556,In_1195,In_778);
nand U557 (N_557,In_1411,In_1253);
or U558 (N_558,In_1335,In_1135);
xor U559 (N_559,In_518,In_663);
nor U560 (N_560,In_656,In_124);
or U561 (N_561,In_949,In_242);
and U562 (N_562,In_716,In_1031);
or U563 (N_563,In_810,In_742);
or U564 (N_564,In_1464,In_713);
or U565 (N_565,In_1085,In_422);
nand U566 (N_566,In_135,In_83);
and U567 (N_567,In_587,In_1240);
or U568 (N_568,In_22,In_852);
and U569 (N_569,In_156,In_51);
nor U570 (N_570,In_112,In_508);
xnor U571 (N_571,In_1460,In_1346);
or U572 (N_572,In_1020,In_1228);
or U573 (N_573,In_829,In_274);
or U574 (N_574,In_1430,In_679);
nand U575 (N_575,In_757,In_926);
nand U576 (N_576,In_2,In_103);
or U577 (N_577,In_1120,In_729);
xnor U578 (N_578,In_389,In_1150);
nand U579 (N_579,In_1000,In_1200);
and U580 (N_580,In_538,In_1191);
and U581 (N_581,In_1280,In_971);
nor U582 (N_582,In_932,In_14);
nand U583 (N_583,In_119,In_1241);
or U584 (N_584,In_65,In_350);
nor U585 (N_585,In_275,In_689);
xor U586 (N_586,In_1337,In_1180);
nand U587 (N_587,In_326,In_214);
xor U588 (N_588,In_1342,In_1294);
nor U589 (N_589,In_1393,In_644);
nor U590 (N_590,In_1312,In_950);
nand U591 (N_591,In_424,In_1044);
xor U592 (N_592,In_797,In_1161);
and U593 (N_593,In_948,In_329);
nor U594 (N_594,In_378,In_862);
nor U595 (N_595,In_886,In_1251);
nor U596 (N_596,In_1317,In_1145);
and U597 (N_597,In_850,In_877);
nand U598 (N_598,In_252,In_159);
or U599 (N_599,In_918,In_953);
nand U600 (N_600,In_140,In_1354);
xnor U601 (N_601,In_588,In_1278);
nand U602 (N_602,In_394,In_1172);
nor U603 (N_603,In_155,In_218);
or U604 (N_604,In_66,In_57);
nand U605 (N_605,In_762,In_1131);
xnor U606 (N_606,In_332,In_752);
nand U607 (N_607,In_1499,In_473);
nor U608 (N_608,In_996,In_546);
and U609 (N_609,In_545,In_549);
xor U610 (N_610,In_901,In_231);
xor U611 (N_611,In_277,In_876);
xnor U612 (N_612,In_45,In_194);
nor U613 (N_613,In_56,In_1444);
nor U614 (N_614,In_528,In_687);
or U615 (N_615,In_413,In_900);
nor U616 (N_616,In_309,In_427);
or U617 (N_617,In_1199,In_58);
xor U618 (N_618,In_1186,In_609);
and U619 (N_619,In_550,In_510);
nand U620 (N_620,In_175,In_1094);
nor U621 (N_621,In_1284,In_1273);
nor U622 (N_622,In_812,In_480);
and U623 (N_623,In_1472,In_962);
or U624 (N_624,In_717,In_530);
xnor U625 (N_625,In_673,In_1205);
or U626 (N_626,In_991,In_1058);
or U627 (N_627,In_108,In_1293);
or U628 (N_628,In_1104,In_905);
nand U629 (N_629,In_665,In_1125);
nand U630 (N_630,In_1402,In_967);
xor U631 (N_631,In_383,In_1024);
nand U632 (N_632,In_360,In_199);
and U633 (N_633,In_937,In_1345);
and U634 (N_634,In_432,In_43);
or U635 (N_635,In_190,In_1243);
xnor U636 (N_636,In_793,In_1155);
nor U637 (N_637,In_1065,In_551);
nor U638 (N_638,In_1211,In_1282);
nand U639 (N_639,In_584,In_559);
nor U640 (N_640,In_523,In_1308);
nor U641 (N_641,In_76,In_1315);
and U642 (N_642,In_1399,In_1016);
nor U643 (N_643,In_6,In_795);
nor U644 (N_644,In_468,In_436);
or U645 (N_645,In_881,In_1368);
or U646 (N_646,In_944,In_825);
nor U647 (N_647,In_290,In_498);
nor U648 (N_648,In_562,In_100);
xnor U649 (N_649,In_1263,In_1413);
nand U650 (N_650,In_284,In_15);
nor U651 (N_651,In_532,In_720);
nand U652 (N_652,In_668,In_313);
or U653 (N_653,In_230,In_1214);
and U654 (N_654,In_210,In_516);
nand U655 (N_655,In_11,In_771);
nor U656 (N_656,In_363,In_323);
or U657 (N_657,In_954,In_324);
xor U658 (N_658,In_1208,In_775);
and U659 (N_659,In_1366,In_1010);
xnor U660 (N_660,In_192,In_1229);
nand U661 (N_661,In_1257,In_553);
and U662 (N_662,In_1364,In_1298);
and U663 (N_663,In_373,In_602);
nand U664 (N_664,In_1103,In_5);
nand U665 (N_665,In_23,In_30);
or U666 (N_666,In_1258,In_561);
nor U667 (N_667,In_305,In_593);
or U668 (N_668,In_197,In_969);
and U669 (N_669,In_405,In_788);
nor U670 (N_670,In_1212,In_1374);
xor U671 (N_671,In_1074,In_132);
or U672 (N_672,In_245,In_964);
nand U673 (N_673,In_1175,In_1022);
xnor U674 (N_674,In_652,In_1124);
nor U675 (N_675,In_1033,In_1334);
xor U676 (N_676,In_701,In_1171);
or U677 (N_677,In_1492,In_933);
and U678 (N_678,In_699,In_992);
and U679 (N_679,In_1187,In_989);
nand U680 (N_680,In_1463,In_1224);
nand U681 (N_681,In_572,In_281);
xnor U682 (N_682,In_1389,In_1118);
nor U683 (N_683,In_439,In_248);
and U684 (N_684,In_307,In_536);
nand U685 (N_685,In_785,In_979);
nand U686 (N_686,In_449,In_1216);
nor U687 (N_687,In_718,In_1115);
xor U688 (N_688,In_474,In_750);
or U689 (N_689,In_982,In_280);
nor U690 (N_690,In_1340,In_955);
nand U691 (N_691,In_70,In_904);
nor U692 (N_692,In_1445,In_1495);
xnor U693 (N_693,In_1268,In_467);
xor U694 (N_694,In_1387,In_1325);
nor U695 (N_695,In_44,In_921);
or U696 (N_696,In_1210,In_98);
nand U697 (N_697,In_279,In_1063);
xnor U698 (N_698,In_1452,In_911);
nand U699 (N_699,In_1136,In_392);
xnor U700 (N_700,In_1068,In_302);
nand U701 (N_701,In_1067,In_1378);
or U702 (N_702,In_171,In_203);
nand U703 (N_703,In_624,In_42);
and U704 (N_704,In_753,In_710);
nand U705 (N_705,In_1173,In_813);
nand U706 (N_706,In_923,In_1220);
nand U707 (N_707,In_846,In_865);
nor U708 (N_708,In_1420,In_89);
xor U709 (N_709,In_784,In_961);
nor U710 (N_710,In_1040,In_875);
nand U711 (N_711,In_1274,In_1163);
nor U712 (N_712,In_1098,In_1482);
or U713 (N_713,In_749,In_1424);
nand U714 (N_714,In_292,In_776);
xnor U715 (N_715,In_1403,In_166);
nor U716 (N_716,In_524,In_1193);
nor U717 (N_717,In_77,In_998);
xnor U718 (N_718,In_557,In_289);
and U719 (N_719,In_173,In_477);
nand U720 (N_720,In_364,In_859);
nand U721 (N_721,In_1428,In_973);
or U722 (N_722,In_897,In_353);
or U723 (N_723,In_337,In_1015);
nor U724 (N_724,In_774,In_704);
or U725 (N_725,In_734,In_554);
xnor U726 (N_726,In_1480,In_1129);
and U727 (N_727,In_482,In_1114);
and U728 (N_728,In_300,In_1493);
nand U729 (N_729,In_1300,In_78);
and U730 (N_730,In_1422,In_1032);
nor U731 (N_731,In_240,In_934);
and U732 (N_732,In_1112,In_763);
or U733 (N_733,In_1009,In_52);
nor U734 (N_734,In_1417,In_678);
nor U735 (N_735,In_636,In_1377);
or U736 (N_736,In_1394,In_891);
nor U737 (N_737,In_980,In_615);
xnor U738 (N_738,In_299,In_263);
nand U739 (N_739,In_1270,In_1353);
xor U740 (N_740,In_1259,In_1247);
nand U741 (N_741,In_521,In_1168);
nand U742 (N_742,In_604,In_415);
nand U743 (N_743,In_555,In_386);
nand U744 (N_744,In_563,In_997);
or U745 (N_745,In_817,In_398);
xnor U746 (N_746,In_419,In_377);
nor U747 (N_747,In_397,In_990);
xor U748 (N_748,In_1418,In_32);
xor U749 (N_749,In_931,In_892);
or U750 (N_750,In_1220,In_646);
and U751 (N_751,In_1014,In_255);
or U752 (N_752,In_959,In_1093);
xor U753 (N_753,In_276,In_902);
nor U754 (N_754,In_105,In_461);
nand U755 (N_755,In_1296,In_95);
or U756 (N_756,In_975,In_564);
xor U757 (N_757,In_649,In_1178);
nor U758 (N_758,In_704,In_1019);
xor U759 (N_759,In_471,In_87);
nand U760 (N_760,In_734,In_504);
xnor U761 (N_761,In_564,In_23);
nand U762 (N_762,In_1293,In_423);
and U763 (N_763,In_837,In_1137);
and U764 (N_764,In_761,In_389);
nor U765 (N_765,In_1120,In_165);
or U766 (N_766,In_823,In_524);
nand U767 (N_767,In_444,In_166);
nand U768 (N_768,In_543,In_1281);
nand U769 (N_769,In_1197,In_1028);
or U770 (N_770,In_1047,In_130);
and U771 (N_771,In_889,In_1485);
or U772 (N_772,In_944,In_1453);
and U773 (N_773,In_93,In_1462);
nand U774 (N_774,In_1,In_1361);
xor U775 (N_775,In_1276,In_1076);
nor U776 (N_776,In_626,In_1428);
or U777 (N_777,In_1022,In_484);
nor U778 (N_778,In_597,In_809);
xor U779 (N_779,In_357,In_1410);
nand U780 (N_780,In_827,In_35);
nand U781 (N_781,In_1236,In_1347);
nand U782 (N_782,In_20,In_27);
or U783 (N_783,In_292,In_1174);
and U784 (N_784,In_555,In_743);
and U785 (N_785,In_237,In_1302);
or U786 (N_786,In_1242,In_888);
or U787 (N_787,In_277,In_401);
or U788 (N_788,In_982,In_481);
and U789 (N_789,In_18,In_886);
xor U790 (N_790,In_372,In_48);
xnor U791 (N_791,In_44,In_759);
or U792 (N_792,In_905,In_1372);
nand U793 (N_793,In_1255,In_1052);
and U794 (N_794,In_124,In_1389);
and U795 (N_795,In_740,In_1342);
or U796 (N_796,In_1459,In_667);
nand U797 (N_797,In_856,In_1038);
and U798 (N_798,In_992,In_200);
xnor U799 (N_799,In_805,In_1108);
nor U800 (N_800,In_451,In_670);
nand U801 (N_801,In_41,In_790);
and U802 (N_802,In_476,In_771);
xor U803 (N_803,In_944,In_1465);
and U804 (N_804,In_1013,In_458);
nor U805 (N_805,In_1427,In_470);
nand U806 (N_806,In_1215,In_569);
xor U807 (N_807,In_398,In_13);
xor U808 (N_808,In_15,In_647);
nor U809 (N_809,In_845,In_1134);
and U810 (N_810,In_716,In_678);
nand U811 (N_811,In_976,In_1211);
xor U812 (N_812,In_1137,In_1181);
xnor U813 (N_813,In_261,In_218);
nand U814 (N_814,In_319,In_1029);
and U815 (N_815,In_531,In_257);
and U816 (N_816,In_1224,In_300);
or U817 (N_817,In_1008,In_706);
nand U818 (N_818,In_1152,In_252);
or U819 (N_819,In_1165,In_32);
xor U820 (N_820,In_653,In_787);
nor U821 (N_821,In_457,In_343);
and U822 (N_822,In_768,In_495);
xnor U823 (N_823,In_1371,In_1372);
and U824 (N_824,In_87,In_358);
and U825 (N_825,In_822,In_752);
and U826 (N_826,In_735,In_198);
nand U827 (N_827,In_1361,In_1458);
xor U828 (N_828,In_1082,In_1027);
xnor U829 (N_829,In_197,In_13);
or U830 (N_830,In_725,In_1020);
nor U831 (N_831,In_863,In_184);
nor U832 (N_832,In_393,In_1134);
or U833 (N_833,In_1192,In_1421);
and U834 (N_834,In_320,In_1042);
or U835 (N_835,In_102,In_1210);
or U836 (N_836,In_333,In_317);
or U837 (N_837,In_1231,In_1186);
nor U838 (N_838,In_770,In_717);
and U839 (N_839,In_248,In_380);
nor U840 (N_840,In_841,In_1011);
xnor U841 (N_841,In_571,In_549);
nand U842 (N_842,In_1338,In_1131);
and U843 (N_843,In_254,In_786);
or U844 (N_844,In_801,In_592);
and U845 (N_845,In_923,In_983);
and U846 (N_846,In_1361,In_626);
nand U847 (N_847,In_0,In_420);
xor U848 (N_848,In_426,In_1137);
nand U849 (N_849,In_919,In_69);
or U850 (N_850,In_927,In_1017);
nor U851 (N_851,In_199,In_1287);
and U852 (N_852,In_1066,In_795);
nand U853 (N_853,In_439,In_1067);
xnor U854 (N_854,In_1287,In_157);
or U855 (N_855,In_1051,In_1020);
or U856 (N_856,In_117,In_1470);
or U857 (N_857,In_1042,In_1260);
nor U858 (N_858,In_1325,In_346);
xor U859 (N_859,In_1074,In_855);
nand U860 (N_860,In_1175,In_8);
nand U861 (N_861,In_707,In_135);
and U862 (N_862,In_315,In_1028);
and U863 (N_863,In_1102,In_1363);
xor U864 (N_864,In_1422,In_109);
xor U865 (N_865,In_1410,In_851);
and U866 (N_866,In_1376,In_1231);
xor U867 (N_867,In_1355,In_155);
xor U868 (N_868,In_308,In_750);
or U869 (N_869,In_1355,In_916);
and U870 (N_870,In_812,In_829);
or U871 (N_871,In_233,In_166);
nor U872 (N_872,In_436,In_652);
nand U873 (N_873,In_689,In_22);
xor U874 (N_874,In_50,In_18);
or U875 (N_875,In_1310,In_23);
or U876 (N_876,In_365,In_585);
or U877 (N_877,In_22,In_1115);
nor U878 (N_878,In_1084,In_945);
or U879 (N_879,In_876,In_1039);
and U880 (N_880,In_453,In_848);
nor U881 (N_881,In_574,In_861);
and U882 (N_882,In_943,In_1214);
or U883 (N_883,In_478,In_499);
nor U884 (N_884,In_803,In_1384);
nor U885 (N_885,In_1482,In_62);
nand U886 (N_886,In_786,In_1337);
nand U887 (N_887,In_1377,In_977);
xnor U888 (N_888,In_293,In_128);
or U889 (N_889,In_930,In_1438);
xnor U890 (N_890,In_1109,In_75);
xor U891 (N_891,In_756,In_1312);
and U892 (N_892,In_145,In_1382);
nor U893 (N_893,In_1427,In_309);
and U894 (N_894,In_156,In_914);
xnor U895 (N_895,In_423,In_1028);
or U896 (N_896,In_362,In_81);
nand U897 (N_897,In_1117,In_863);
or U898 (N_898,In_447,In_618);
and U899 (N_899,In_724,In_1408);
xor U900 (N_900,In_946,In_496);
xnor U901 (N_901,In_383,In_1054);
nor U902 (N_902,In_1480,In_1283);
xnor U903 (N_903,In_1172,In_1332);
nand U904 (N_904,In_761,In_97);
or U905 (N_905,In_739,In_1323);
nor U906 (N_906,In_130,In_207);
nand U907 (N_907,In_599,In_1016);
nand U908 (N_908,In_885,In_105);
nand U909 (N_909,In_564,In_1349);
xor U910 (N_910,In_259,In_384);
xor U911 (N_911,In_1470,In_44);
and U912 (N_912,In_933,In_187);
or U913 (N_913,In_561,In_1325);
nor U914 (N_914,In_1394,In_1431);
or U915 (N_915,In_1421,In_1346);
xnor U916 (N_916,In_1333,In_1479);
nand U917 (N_917,In_789,In_540);
xnor U918 (N_918,In_939,In_1129);
or U919 (N_919,In_1300,In_887);
nor U920 (N_920,In_570,In_54);
and U921 (N_921,In_1018,In_1227);
and U922 (N_922,In_1096,In_1077);
and U923 (N_923,In_1248,In_397);
xor U924 (N_924,In_1441,In_1358);
nor U925 (N_925,In_1462,In_243);
or U926 (N_926,In_878,In_541);
nor U927 (N_927,In_447,In_579);
or U928 (N_928,In_239,In_456);
or U929 (N_929,In_879,In_1292);
nor U930 (N_930,In_1202,In_1311);
nor U931 (N_931,In_211,In_441);
nor U932 (N_932,In_288,In_86);
nor U933 (N_933,In_1070,In_707);
and U934 (N_934,In_839,In_924);
nand U935 (N_935,In_886,In_632);
nand U936 (N_936,In_1065,In_27);
xor U937 (N_937,In_41,In_725);
xor U938 (N_938,In_829,In_1071);
and U939 (N_939,In_621,In_365);
nand U940 (N_940,In_995,In_1295);
or U941 (N_941,In_1396,In_1056);
or U942 (N_942,In_1283,In_906);
and U943 (N_943,In_16,In_399);
nor U944 (N_944,In_1253,In_798);
or U945 (N_945,In_1421,In_1160);
or U946 (N_946,In_46,In_428);
xnor U947 (N_947,In_538,In_1454);
and U948 (N_948,In_1261,In_1032);
or U949 (N_949,In_156,In_717);
or U950 (N_950,In_49,In_1481);
or U951 (N_951,In_913,In_448);
nor U952 (N_952,In_1025,In_25);
and U953 (N_953,In_208,In_222);
xor U954 (N_954,In_1189,In_762);
nand U955 (N_955,In_440,In_808);
nor U956 (N_956,In_404,In_670);
nand U957 (N_957,In_451,In_762);
and U958 (N_958,In_1196,In_512);
xnor U959 (N_959,In_1252,In_1192);
or U960 (N_960,In_778,In_1353);
and U961 (N_961,In_365,In_43);
and U962 (N_962,In_816,In_1091);
nor U963 (N_963,In_1174,In_1316);
and U964 (N_964,In_1390,In_807);
or U965 (N_965,In_623,In_1421);
nor U966 (N_966,In_370,In_922);
nor U967 (N_967,In_1369,In_371);
nand U968 (N_968,In_473,In_1127);
nor U969 (N_969,In_673,In_38);
xnor U970 (N_970,In_1296,In_549);
xnor U971 (N_971,In_1130,In_180);
nor U972 (N_972,In_1220,In_700);
or U973 (N_973,In_552,In_894);
nand U974 (N_974,In_497,In_630);
and U975 (N_975,In_1345,In_321);
or U976 (N_976,In_905,In_1184);
nor U977 (N_977,In_186,In_1218);
or U978 (N_978,In_685,In_1036);
nor U979 (N_979,In_85,In_621);
or U980 (N_980,In_1023,In_76);
xor U981 (N_981,In_90,In_735);
nand U982 (N_982,In_1173,In_223);
or U983 (N_983,In_987,In_1413);
and U984 (N_984,In_935,In_1098);
xor U985 (N_985,In_191,In_294);
xor U986 (N_986,In_442,In_14);
or U987 (N_987,In_1481,In_1108);
or U988 (N_988,In_1213,In_1044);
nand U989 (N_989,In_18,In_332);
and U990 (N_990,In_292,In_569);
and U991 (N_991,In_104,In_616);
nor U992 (N_992,In_989,In_416);
xor U993 (N_993,In_567,In_393);
xor U994 (N_994,In_1018,In_8);
xor U995 (N_995,In_550,In_1473);
and U996 (N_996,In_365,In_481);
or U997 (N_997,In_160,In_1148);
and U998 (N_998,In_1087,In_1198);
nor U999 (N_999,In_1178,In_1369);
and U1000 (N_1000,In_828,In_388);
nand U1001 (N_1001,In_915,In_151);
nand U1002 (N_1002,In_1302,In_678);
or U1003 (N_1003,In_709,In_697);
nor U1004 (N_1004,In_480,In_182);
nor U1005 (N_1005,In_1030,In_702);
xor U1006 (N_1006,In_185,In_212);
xnor U1007 (N_1007,In_1051,In_230);
or U1008 (N_1008,In_509,In_380);
or U1009 (N_1009,In_1390,In_328);
xor U1010 (N_1010,In_1218,In_1328);
or U1011 (N_1011,In_986,In_723);
nor U1012 (N_1012,In_154,In_695);
xor U1013 (N_1013,In_1212,In_599);
and U1014 (N_1014,In_757,In_1158);
xnor U1015 (N_1015,In_216,In_737);
nand U1016 (N_1016,In_151,In_142);
nor U1017 (N_1017,In_1063,In_950);
or U1018 (N_1018,In_1352,In_427);
or U1019 (N_1019,In_1300,In_1229);
and U1020 (N_1020,In_639,In_110);
xor U1021 (N_1021,In_1422,In_100);
nand U1022 (N_1022,In_137,In_490);
and U1023 (N_1023,In_1286,In_645);
nor U1024 (N_1024,In_1381,In_1226);
and U1025 (N_1025,In_1449,In_1330);
nor U1026 (N_1026,In_593,In_821);
and U1027 (N_1027,In_666,In_1092);
or U1028 (N_1028,In_139,In_1228);
xor U1029 (N_1029,In_1474,In_572);
and U1030 (N_1030,In_353,In_1245);
and U1031 (N_1031,In_589,In_49);
nor U1032 (N_1032,In_118,In_1200);
nand U1033 (N_1033,In_14,In_935);
and U1034 (N_1034,In_452,In_155);
nand U1035 (N_1035,In_677,In_510);
xor U1036 (N_1036,In_929,In_654);
and U1037 (N_1037,In_877,In_520);
nor U1038 (N_1038,In_664,In_926);
and U1039 (N_1039,In_622,In_523);
nor U1040 (N_1040,In_1492,In_499);
nor U1041 (N_1041,In_803,In_991);
nand U1042 (N_1042,In_25,In_703);
or U1043 (N_1043,In_69,In_1441);
nor U1044 (N_1044,In_903,In_861);
xor U1045 (N_1045,In_11,In_686);
or U1046 (N_1046,In_73,In_187);
nor U1047 (N_1047,In_1184,In_1290);
nor U1048 (N_1048,In_741,In_1172);
xnor U1049 (N_1049,In_235,In_469);
and U1050 (N_1050,In_1203,In_1146);
nor U1051 (N_1051,In_478,In_759);
or U1052 (N_1052,In_1485,In_990);
and U1053 (N_1053,In_476,In_803);
and U1054 (N_1054,In_222,In_290);
nand U1055 (N_1055,In_415,In_617);
xor U1056 (N_1056,In_1058,In_914);
xnor U1057 (N_1057,In_112,In_137);
nor U1058 (N_1058,In_927,In_1386);
and U1059 (N_1059,In_1215,In_796);
or U1060 (N_1060,In_1484,In_655);
and U1061 (N_1061,In_769,In_267);
or U1062 (N_1062,In_287,In_939);
and U1063 (N_1063,In_1161,In_815);
or U1064 (N_1064,In_155,In_1157);
or U1065 (N_1065,In_1397,In_54);
nand U1066 (N_1066,In_1493,In_1058);
or U1067 (N_1067,In_640,In_761);
and U1068 (N_1068,In_1199,In_14);
or U1069 (N_1069,In_1331,In_994);
nor U1070 (N_1070,In_84,In_1157);
nor U1071 (N_1071,In_89,In_967);
nand U1072 (N_1072,In_679,In_1244);
nand U1073 (N_1073,In_1125,In_890);
xor U1074 (N_1074,In_530,In_12);
xnor U1075 (N_1075,In_575,In_169);
nor U1076 (N_1076,In_763,In_857);
nor U1077 (N_1077,In_386,In_1473);
xnor U1078 (N_1078,In_402,In_1184);
xor U1079 (N_1079,In_902,In_183);
nand U1080 (N_1080,In_54,In_1366);
nor U1081 (N_1081,In_96,In_1403);
xnor U1082 (N_1082,In_1466,In_1288);
and U1083 (N_1083,In_75,In_952);
and U1084 (N_1084,In_288,In_228);
xor U1085 (N_1085,In_166,In_75);
xor U1086 (N_1086,In_1138,In_9);
or U1087 (N_1087,In_799,In_940);
nand U1088 (N_1088,In_87,In_746);
or U1089 (N_1089,In_999,In_203);
or U1090 (N_1090,In_84,In_1394);
xor U1091 (N_1091,In_481,In_1437);
nand U1092 (N_1092,In_1135,In_1403);
nand U1093 (N_1093,In_484,In_1008);
xor U1094 (N_1094,In_783,In_26);
nor U1095 (N_1095,In_577,In_1399);
xnor U1096 (N_1096,In_1450,In_856);
or U1097 (N_1097,In_1419,In_650);
nand U1098 (N_1098,In_885,In_163);
and U1099 (N_1099,In_595,In_16);
nor U1100 (N_1100,In_754,In_1079);
nor U1101 (N_1101,In_969,In_1090);
or U1102 (N_1102,In_441,In_118);
nand U1103 (N_1103,In_1447,In_1343);
or U1104 (N_1104,In_60,In_172);
nand U1105 (N_1105,In_395,In_939);
or U1106 (N_1106,In_1469,In_549);
xor U1107 (N_1107,In_833,In_67);
and U1108 (N_1108,In_956,In_1154);
nor U1109 (N_1109,In_599,In_1166);
xor U1110 (N_1110,In_1212,In_1481);
nand U1111 (N_1111,In_416,In_165);
and U1112 (N_1112,In_1413,In_75);
xnor U1113 (N_1113,In_1113,In_108);
nand U1114 (N_1114,In_431,In_616);
or U1115 (N_1115,In_349,In_1318);
nand U1116 (N_1116,In_568,In_882);
xor U1117 (N_1117,In_416,In_1133);
xnor U1118 (N_1118,In_97,In_128);
or U1119 (N_1119,In_1314,In_1337);
xnor U1120 (N_1120,In_1392,In_178);
or U1121 (N_1121,In_730,In_922);
and U1122 (N_1122,In_229,In_530);
nor U1123 (N_1123,In_803,In_1183);
or U1124 (N_1124,In_1328,In_31);
nor U1125 (N_1125,In_1123,In_299);
nor U1126 (N_1126,In_1397,In_1429);
xnor U1127 (N_1127,In_180,In_366);
or U1128 (N_1128,In_573,In_1218);
nor U1129 (N_1129,In_57,In_767);
nand U1130 (N_1130,In_1282,In_1249);
nor U1131 (N_1131,In_765,In_1136);
nand U1132 (N_1132,In_643,In_932);
nor U1133 (N_1133,In_1098,In_82);
xnor U1134 (N_1134,In_784,In_1272);
or U1135 (N_1135,In_1120,In_152);
and U1136 (N_1136,In_217,In_1210);
nand U1137 (N_1137,In_1142,In_620);
nor U1138 (N_1138,In_1261,In_504);
and U1139 (N_1139,In_873,In_557);
xor U1140 (N_1140,In_1497,In_902);
nand U1141 (N_1141,In_1479,In_214);
nand U1142 (N_1142,In_1487,In_817);
nor U1143 (N_1143,In_451,In_154);
and U1144 (N_1144,In_169,In_1134);
and U1145 (N_1145,In_1422,In_145);
nor U1146 (N_1146,In_1235,In_532);
or U1147 (N_1147,In_413,In_373);
nor U1148 (N_1148,In_612,In_413);
xnor U1149 (N_1149,In_1199,In_1077);
and U1150 (N_1150,In_1160,In_610);
or U1151 (N_1151,In_1217,In_464);
or U1152 (N_1152,In_569,In_1083);
nand U1153 (N_1153,In_601,In_283);
nand U1154 (N_1154,In_1149,In_596);
nand U1155 (N_1155,In_926,In_298);
or U1156 (N_1156,In_11,In_64);
and U1157 (N_1157,In_780,In_53);
xnor U1158 (N_1158,In_1141,In_542);
xnor U1159 (N_1159,In_702,In_181);
xor U1160 (N_1160,In_1144,In_625);
or U1161 (N_1161,In_538,In_183);
and U1162 (N_1162,In_540,In_259);
xor U1163 (N_1163,In_805,In_251);
or U1164 (N_1164,In_286,In_1277);
nand U1165 (N_1165,In_686,In_1299);
nand U1166 (N_1166,In_628,In_36);
xnor U1167 (N_1167,In_1165,In_879);
or U1168 (N_1168,In_743,In_1301);
nand U1169 (N_1169,In_440,In_94);
xor U1170 (N_1170,In_797,In_400);
and U1171 (N_1171,In_1020,In_91);
and U1172 (N_1172,In_150,In_179);
nand U1173 (N_1173,In_1424,In_302);
nor U1174 (N_1174,In_198,In_1491);
and U1175 (N_1175,In_738,In_567);
nor U1176 (N_1176,In_1420,In_85);
or U1177 (N_1177,In_1240,In_1339);
and U1178 (N_1178,In_1390,In_936);
and U1179 (N_1179,In_751,In_1395);
or U1180 (N_1180,In_1344,In_1111);
nand U1181 (N_1181,In_1002,In_160);
nor U1182 (N_1182,In_1341,In_681);
xor U1183 (N_1183,In_1329,In_1034);
nor U1184 (N_1184,In_289,In_1428);
nor U1185 (N_1185,In_1337,In_1453);
nand U1186 (N_1186,In_136,In_1415);
nand U1187 (N_1187,In_220,In_621);
nand U1188 (N_1188,In_1343,In_1063);
nor U1189 (N_1189,In_746,In_141);
and U1190 (N_1190,In_1396,In_831);
nand U1191 (N_1191,In_269,In_513);
or U1192 (N_1192,In_941,In_1196);
and U1193 (N_1193,In_1334,In_245);
xor U1194 (N_1194,In_299,In_1164);
nand U1195 (N_1195,In_1485,In_696);
xnor U1196 (N_1196,In_647,In_631);
xor U1197 (N_1197,In_941,In_971);
xor U1198 (N_1198,In_15,In_740);
xor U1199 (N_1199,In_478,In_1370);
and U1200 (N_1200,In_501,In_139);
nor U1201 (N_1201,In_764,In_395);
xnor U1202 (N_1202,In_323,In_1043);
and U1203 (N_1203,In_1337,In_852);
nand U1204 (N_1204,In_635,In_77);
nand U1205 (N_1205,In_1454,In_327);
or U1206 (N_1206,In_542,In_359);
nor U1207 (N_1207,In_452,In_43);
nand U1208 (N_1208,In_301,In_225);
nand U1209 (N_1209,In_1408,In_616);
or U1210 (N_1210,In_285,In_139);
xor U1211 (N_1211,In_316,In_567);
nand U1212 (N_1212,In_547,In_732);
nor U1213 (N_1213,In_398,In_642);
nand U1214 (N_1214,In_1101,In_1317);
nand U1215 (N_1215,In_680,In_379);
or U1216 (N_1216,In_471,In_708);
xor U1217 (N_1217,In_795,In_1386);
nor U1218 (N_1218,In_958,In_812);
nor U1219 (N_1219,In_1212,In_324);
or U1220 (N_1220,In_451,In_1207);
nand U1221 (N_1221,In_1199,In_1042);
or U1222 (N_1222,In_390,In_1348);
xor U1223 (N_1223,In_976,In_296);
or U1224 (N_1224,In_1196,In_173);
xor U1225 (N_1225,In_102,In_1083);
or U1226 (N_1226,In_589,In_1209);
nor U1227 (N_1227,In_715,In_963);
nor U1228 (N_1228,In_1210,In_260);
or U1229 (N_1229,In_596,In_407);
nand U1230 (N_1230,In_595,In_1425);
and U1231 (N_1231,In_386,In_1218);
xnor U1232 (N_1232,In_569,In_1439);
xnor U1233 (N_1233,In_349,In_1159);
xnor U1234 (N_1234,In_673,In_884);
nand U1235 (N_1235,In_144,In_1165);
xor U1236 (N_1236,In_497,In_1133);
or U1237 (N_1237,In_908,In_298);
nor U1238 (N_1238,In_535,In_294);
xnor U1239 (N_1239,In_1026,In_435);
xor U1240 (N_1240,In_169,In_742);
and U1241 (N_1241,In_1340,In_102);
nor U1242 (N_1242,In_492,In_1280);
xor U1243 (N_1243,In_189,In_1467);
and U1244 (N_1244,In_304,In_439);
xnor U1245 (N_1245,In_36,In_1473);
or U1246 (N_1246,In_570,In_223);
xor U1247 (N_1247,In_454,In_1201);
and U1248 (N_1248,In_1171,In_461);
nand U1249 (N_1249,In_1393,In_1288);
xor U1250 (N_1250,In_412,In_10);
xor U1251 (N_1251,In_723,In_170);
xnor U1252 (N_1252,In_164,In_427);
or U1253 (N_1253,In_1169,In_509);
nand U1254 (N_1254,In_1107,In_482);
xor U1255 (N_1255,In_643,In_1040);
or U1256 (N_1256,In_1284,In_1035);
xnor U1257 (N_1257,In_455,In_443);
xor U1258 (N_1258,In_218,In_853);
nand U1259 (N_1259,In_1018,In_933);
or U1260 (N_1260,In_207,In_88);
or U1261 (N_1261,In_1123,In_795);
xnor U1262 (N_1262,In_350,In_339);
xor U1263 (N_1263,In_444,In_804);
nor U1264 (N_1264,In_526,In_1143);
or U1265 (N_1265,In_106,In_1427);
nand U1266 (N_1266,In_1469,In_239);
nand U1267 (N_1267,In_1263,In_1191);
and U1268 (N_1268,In_162,In_1018);
nor U1269 (N_1269,In_384,In_756);
nor U1270 (N_1270,In_1196,In_444);
xnor U1271 (N_1271,In_925,In_10);
or U1272 (N_1272,In_844,In_508);
nor U1273 (N_1273,In_56,In_1380);
or U1274 (N_1274,In_132,In_130);
and U1275 (N_1275,In_294,In_474);
nor U1276 (N_1276,In_1148,In_674);
nand U1277 (N_1277,In_480,In_1001);
and U1278 (N_1278,In_676,In_169);
nand U1279 (N_1279,In_1191,In_1056);
nor U1280 (N_1280,In_983,In_963);
xor U1281 (N_1281,In_457,In_1190);
or U1282 (N_1282,In_1364,In_1105);
xnor U1283 (N_1283,In_707,In_85);
and U1284 (N_1284,In_747,In_108);
xnor U1285 (N_1285,In_1349,In_150);
nor U1286 (N_1286,In_527,In_899);
xor U1287 (N_1287,In_1000,In_1029);
and U1288 (N_1288,In_768,In_1125);
xnor U1289 (N_1289,In_629,In_710);
or U1290 (N_1290,In_327,In_113);
or U1291 (N_1291,In_34,In_677);
and U1292 (N_1292,In_130,In_1360);
nand U1293 (N_1293,In_952,In_821);
xor U1294 (N_1294,In_1228,In_401);
xor U1295 (N_1295,In_865,In_881);
nand U1296 (N_1296,In_748,In_103);
nand U1297 (N_1297,In_697,In_46);
nor U1298 (N_1298,In_24,In_855);
xnor U1299 (N_1299,In_797,In_1487);
nand U1300 (N_1300,In_342,In_1045);
xnor U1301 (N_1301,In_880,In_236);
nand U1302 (N_1302,In_5,In_272);
and U1303 (N_1303,In_1064,In_6);
nor U1304 (N_1304,In_922,In_1056);
xnor U1305 (N_1305,In_901,In_1289);
xor U1306 (N_1306,In_157,In_314);
and U1307 (N_1307,In_662,In_778);
nor U1308 (N_1308,In_282,In_860);
nand U1309 (N_1309,In_216,In_1);
xor U1310 (N_1310,In_1269,In_422);
nor U1311 (N_1311,In_422,In_763);
or U1312 (N_1312,In_688,In_490);
nand U1313 (N_1313,In_440,In_766);
nor U1314 (N_1314,In_805,In_738);
xnor U1315 (N_1315,In_410,In_296);
xnor U1316 (N_1316,In_370,In_253);
and U1317 (N_1317,In_777,In_289);
nor U1318 (N_1318,In_575,In_1400);
xor U1319 (N_1319,In_1049,In_565);
nor U1320 (N_1320,In_937,In_825);
and U1321 (N_1321,In_1194,In_289);
xor U1322 (N_1322,In_722,In_1203);
nand U1323 (N_1323,In_963,In_81);
nand U1324 (N_1324,In_841,In_980);
nand U1325 (N_1325,In_996,In_135);
or U1326 (N_1326,In_320,In_798);
and U1327 (N_1327,In_1364,In_357);
and U1328 (N_1328,In_1279,In_1347);
nand U1329 (N_1329,In_291,In_144);
xor U1330 (N_1330,In_349,In_42);
nand U1331 (N_1331,In_345,In_1322);
and U1332 (N_1332,In_597,In_136);
nor U1333 (N_1333,In_721,In_1384);
nand U1334 (N_1334,In_1400,In_529);
xnor U1335 (N_1335,In_50,In_134);
nand U1336 (N_1336,In_1025,In_434);
and U1337 (N_1337,In_428,In_1315);
and U1338 (N_1338,In_833,In_1000);
nor U1339 (N_1339,In_1165,In_668);
xnor U1340 (N_1340,In_78,In_882);
nor U1341 (N_1341,In_534,In_1260);
xnor U1342 (N_1342,In_182,In_1167);
nand U1343 (N_1343,In_21,In_1275);
or U1344 (N_1344,In_329,In_1319);
xnor U1345 (N_1345,In_389,In_646);
or U1346 (N_1346,In_1261,In_1258);
xnor U1347 (N_1347,In_1255,In_566);
and U1348 (N_1348,In_1435,In_106);
or U1349 (N_1349,In_707,In_1038);
xnor U1350 (N_1350,In_1206,In_535);
and U1351 (N_1351,In_1269,In_1041);
nand U1352 (N_1352,In_399,In_1073);
and U1353 (N_1353,In_1421,In_1464);
or U1354 (N_1354,In_310,In_482);
or U1355 (N_1355,In_296,In_991);
xor U1356 (N_1356,In_1280,In_102);
or U1357 (N_1357,In_427,In_1439);
and U1358 (N_1358,In_622,In_575);
xor U1359 (N_1359,In_663,In_272);
and U1360 (N_1360,In_1189,In_1303);
nor U1361 (N_1361,In_977,In_279);
nand U1362 (N_1362,In_956,In_136);
xor U1363 (N_1363,In_1217,In_57);
nor U1364 (N_1364,In_930,In_870);
nor U1365 (N_1365,In_1289,In_86);
or U1366 (N_1366,In_458,In_201);
nand U1367 (N_1367,In_1007,In_855);
or U1368 (N_1368,In_1409,In_668);
nand U1369 (N_1369,In_607,In_1026);
xor U1370 (N_1370,In_271,In_1104);
nor U1371 (N_1371,In_63,In_709);
or U1372 (N_1372,In_889,In_1242);
nand U1373 (N_1373,In_723,In_1062);
nor U1374 (N_1374,In_734,In_1465);
nor U1375 (N_1375,In_1162,In_457);
and U1376 (N_1376,In_990,In_430);
nor U1377 (N_1377,In_1104,In_363);
xor U1378 (N_1378,In_873,In_312);
nand U1379 (N_1379,In_1290,In_1474);
or U1380 (N_1380,In_903,In_500);
or U1381 (N_1381,In_128,In_1017);
nor U1382 (N_1382,In_42,In_554);
and U1383 (N_1383,In_1353,In_1099);
xor U1384 (N_1384,In_644,In_1206);
and U1385 (N_1385,In_287,In_1271);
nand U1386 (N_1386,In_389,In_1174);
nor U1387 (N_1387,In_960,In_920);
nor U1388 (N_1388,In_146,In_68);
or U1389 (N_1389,In_949,In_32);
nand U1390 (N_1390,In_626,In_747);
and U1391 (N_1391,In_375,In_1012);
nand U1392 (N_1392,In_652,In_206);
nor U1393 (N_1393,In_884,In_854);
and U1394 (N_1394,In_743,In_228);
nand U1395 (N_1395,In_292,In_600);
nor U1396 (N_1396,In_1490,In_942);
and U1397 (N_1397,In_917,In_210);
xor U1398 (N_1398,In_871,In_708);
nand U1399 (N_1399,In_374,In_294);
xnor U1400 (N_1400,In_1416,In_283);
or U1401 (N_1401,In_940,In_323);
nand U1402 (N_1402,In_1401,In_1020);
and U1403 (N_1403,In_36,In_428);
or U1404 (N_1404,In_477,In_766);
or U1405 (N_1405,In_1247,In_1404);
and U1406 (N_1406,In_1,In_827);
and U1407 (N_1407,In_365,In_690);
nor U1408 (N_1408,In_638,In_781);
and U1409 (N_1409,In_1375,In_936);
nor U1410 (N_1410,In_1404,In_185);
nor U1411 (N_1411,In_474,In_599);
or U1412 (N_1412,In_1153,In_1131);
nor U1413 (N_1413,In_1229,In_1484);
nor U1414 (N_1414,In_616,In_1272);
or U1415 (N_1415,In_7,In_1219);
or U1416 (N_1416,In_531,In_874);
or U1417 (N_1417,In_446,In_744);
and U1418 (N_1418,In_392,In_111);
xor U1419 (N_1419,In_544,In_266);
xnor U1420 (N_1420,In_1395,In_388);
xnor U1421 (N_1421,In_797,In_1211);
and U1422 (N_1422,In_1188,In_903);
xor U1423 (N_1423,In_644,In_327);
and U1424 (N_1424,In_1357,In_1411);
and U1425 (N_1425,In_1163,In_934);
nor U1426 (N_1426,In_1454,In_940);
or U1427 (N_1427,In_136,In_1197);
xnor U1428 (N_1428,In_1316,In_1116);
xor U1429 (N_1429,In_1095,In_124);
or U1430 (N_1430,In_298,In_1221);
or U1431 (N_1431,In_778,In_1390);
or U1432 (N_1432,In_80,In_1273);
or U1433 (N_1433,In_1192,In_372);
nor U1434 (N_1434,In_70,In_175);
nand U1435 (N_1435,In_708,In_703);
nor U1436 (N_1436,In_219,In_174);
xnor U1437 (N_1437,In_169,In_1475);
nor U1438 (N_1438,In_876,In_224);
xnor U1439 (N_1439,In_26,In_1114);
nand U1440 (N_1440,In_105,In_1456);
and U1441 (N_1441,In_430,In_894);
xor U1442 (N_1442,In_120,In_1055);
xor U1443 (N_1443,In_189,In_1160);
nor U1444 (N_1444,In_428,In_1470);
and U1445 (N_1445,In_1442,In_1142);
xor U1446 (N_1446,In_1052,In_914);
or U1447 (N_1447,In_1307,In_1452);
nand U1448 (N_1448,In_1448,In_231);
nand U1449 (N_1449,In_1431,In_1243);
xor U1450 (N_1450,In_1171,In_663);
and U1451 (N_1451,In_1086,In_1301);
nand U1452 (N_1452,In_1242,In_296);
nor U1453 (N_1453,In_573,In_379);
and U1454 (N_1454,In_312,In_1092);
nor U1455 (N_1455,In_306,In_1005);
and U1456 (N_1456,In_174,In_859);
nand U1457 (N_1457,In_67,In_1022);
and U1458 (N_1458,In_407,In_1382);
nor U1459 (N_1459,In_521,In_697);
nand U1460 (N_1460,In_378,In_302);
xnor U1461 (N_1461,In_1427,In_444);
nand U1462 (N_1462,In_134,In_55);
nand U1463 (N_1463,In_1309,In_422);
nand U1464 (N_1464,In_316,In_838);
nand U1465 (N_1465,In_1198,In_1322);
nor U1466 (N_1466,In_1002,In_967);
nand U1467 (N_1467,In_659,In_1108);
xor U1468 (N_1468,In_940,In_706);
nand U1469 (N_1469,In_73,In_522);
and U1470 (N_1470,In_288,In_1496);
nor U1471 (N_1471,In_1461,In_1230);
xnor U1472 (N_1472,In_723,In_40);
nand U1473 (N_1473,In_1222,In_804);
nor U1474 (N_1474,In_74,In_223);
or U1475 (N_1475,In_780,In_1220);
or U1476 (N_1476,In_180,In_1191);
or U1477 (N_1477,In_518,In_1488);
nor U1478 (N_1478,In_185,In_232);
and U1479 (N_1479,In_1136,In_1314);
and U1480 (N_1480,In_791,In_940);
nor U1481 (N_1481,In_811,In_384);
nand U1482 (N_1482,In_7,In_498);
xor U1483 (N_1483,In_493,In_886);
nor U1484 (N_1484,In_611,In_27);
xnor U1485 (N_1485,In_711,In_842);
xor U1486 (N_1486,In_1395,In_265);
nand U1487 (N_1487,In_1092,In_229);
and U1488 (N_1488,In_709,In_567);
and U1489 (N_1489,In_934,In_772);
xor U1490 (N_1490,In_1070,In_1333);
nand U1491 (N_1491,In_1336,In_695);
nand U1492 (N_1492,In_864,In_1390);
nand U1493 (N_1493,In_219,In_491);
or U1494 (N_1494,In_623,In_859);
and U1495 (N_1495,In_62,In_598);
xnor U1496 (N_1496,In_1315,In_902);
or U1497 (N_1497,In_52,In_1424);
xnor U1498 (N_1498,In_810,In_491);
or U1499 (N_1499,In_1210,In_181);
nand U1500 (N_1500,N_1459,N_790);
or U1501 (N_1501,N_1329,N_812);
or U1502 (N_1502,N_373,N_372);
and U1503 (N_1503,N_1402,N_1371);
or U1504 (N_1504,N_9,N_152);
or U1505 (N_1505,N_1084,N_430);
xor U1506 (N_1506,N_573,N_231);
and U1507 (N_1507,N_214,N_1440);
xor U1508 (N_1508,N_1251,N_482);
nor U1509 (N_1509,N_1307,N_1314);
and U1510 (N_1510,N_851,N_1265);
or U1511 (N_1511,N_1190,N_676);
nand U1512 (N_1512,N_157,N_876);
nand U1513 (N_1513,N_888,N_234);
or U1514 (N_1514,N_864,N_1129);
xnor U1515 (N_1515,N_1349,N_654);
nor U1516 (N_1516,N_118,N_756);
nor U1517 (N_1517,N_959,N_636);
nand U1518 (N_1518,N_539,N_287);
or U1519 (N_1519,N_701,N_308);
or U1520 (N_1520,N_1107,N_167);
nand U1521 (N_1521,N_333,N_1237);
nand U1522 (N_1522,N_1000,N_562);
nor U1523 (N_1523,N_1487,N_1474);
and U1524 (N_1524,N_31,N_488);
or U1525 (N_1525,N_720,N_243);
nor U1526 (N_1526,N_613,N_906);
nand U1527 (N_1527,N_924,N_40);
and U1528 (N_1528,N_765,N_1390);
and U1529 (N_1529,N_69,N_615);
nor U1530 (N_1530,N_606,N_137);
nand U1531 (N_1531,N_1416,N_329);
and U1532 (N_1532,N_138,N_1014);
or U1533 (N_1533,N_1223,N_1127);
nor U1534 (N_1534,N_404,N_1472);
xnor U1535 (N_1535,N_650,N_1067);
or U1536 (N_1536,N_1478,N_737);
nand U1537 (N_1537,N_494,N_385);
nor U1538 (N_1538,N_1399,N_938);
nor U1539 (N_1539,N_1176,N_79);
nand U1540 (N_1540,N_810,N_1486);
nor U1541 (N_1541,N_409,N_692);
and U1542 (N_1542,N_403,N_191);
and U1543 (N_1543,N_967,N_1452);
nor U1544 (N_1544,N_658,N_1342);
or U1545 (N_1545,N_664,N_123);
xnor U1546 (N_1546,N_897,N_306);
xor U1547 (N_1547,N_1346,N_1137);
nor U1548 (N_1548,N_192,N_534);
xnor U1549 (N_1549,N_1493,N_608);
nand U1550 (N_1550,N_1445,N_437);
and U1551 (N_1551,N_1386,N_1248);
xor U1552 (N_1552,N_338,N_1074);
nand U1553 (N_1553,N_313,N_49);
or U1554 (N_1554,N_1116,N_297);
or U1555 (N_1555,N_1185,N_1164);
nand U1556 (N_1556,N_1088,N_1274);
and U1557 (N_1557,N_1035,N_408);
and U1558 (N_1558,N_947,N_697);
nand U1559 (N_1559,N_1173,N_1458);
and U1560 (N_1560,N_175,N_750);
and U1561 (N_1561,N_903,N_434);
xor U1562 (N_1562,N_945,N_954);
nand U1563 (N_1563,N_52,N_1213);
nand U1564 (N_1564,N_1049,N_1039);
or U1565 (N_1565,N_193,N_413);
xnor U1566 (N_1566,N_149,N_250);
xor U1567 (N_1567,N_693,N_295);
or U1568 (N_1568,N_1232,N_1465);
nand U1569 (N_1569,N_346,N_13);
and U1570 (N_1570,N_484,N_705);
or U1571 (N_1571,N_1269,N_600);
nand U1572 (N_1572,N_1241,N_1316);
xnor U1573 (N_1573,N_238,N_1080);
xnor U1574 (N_1574,N_28,N_619);
nor U1575 (N_1575,N_112,N_1043);
and U1576 (N_1576,N_163,N_305);
xor U1577 (N_1577,N_1455,N_223);
nand U1578 (N_1578,N_858,N_481);
nor U1579 (N_1579,N_64,N_8);
xnor U1580 (N_1580,N_883,N_828);
or U1581 (N_1581,N_1312,N_367);
xor U1582 (N_1582,N_68,N_104);
nand U1583 (N_1583,N_743,N_1192);
or U1584 (N_1584,N_1436,N_647);
nand U1585 (N_1585,N_337,N_1187);
nor U1586 (N_1586,N_1475,N_171);
or U1587 (N_1587,N_1271,N_953);
and U1588 (N_1588,N_140,N_462);
nor U1589 (N_1589,N_898,N_628);
nor U1590 (N_1590,N_563,N_1380);
or U1591 (N_1591,N_1453,N_1417);
or U1592 (N_1592,N_744,N_880);
xnor U1593 (N_1593,N_727,N_962);
nand U1594 (N_1594,N_801,N_90);
nor U1595 (N_1595,N_679,N_331);
or U1596 (N_1596,N_1471,N_646);
nor U1597 (N_1597,N_141,N_1047);
nand U1598 (N_1598,N_719,N_61);
nor U1599 (N_1599,N_882,N_296);
and U1600 (N_1600,N_82,N_70);
nor U1601 (N_1601,N_702,N_845);
nand U1602 (N_1602,N_1170,N_1369);
or U1603 (N_1603,N_1024,N_94);
xnor U1604 (N_1604,N_1351,N_454);
nor U1605 (N_1605,N_236,N_1256);
nand U1606 (N_1606,N_1037,N_1132);
or U1607 (N_1607,N_607,N_172);
nand U1608 (N_1608,N_46,N_1285);
xnor U1609 (N_1609,N_81,N_728);
xnor U1610 (N_1610,N_849,N_1154);
and U1611 (N_1611,N_211,N_1012);
and U1612 (N_1612,N_1169,N_505);
nand U1613 (N_1613,N_887,N_918);
and U1614 (N_1614,N_1076,N_759);
and U1615 (N_1615,N_922,N_377);
and U1616 (N_1616,N_616,N_1191);
and U1617 (N_1617,N_1004,N_1143);
xor U1618 (N_1618,N_1413,N_30);
and U1619 (N_1619,N_1336,N_354);
xnor U1620 (N_1620,N_785,N_17);
nor U1621 (N_1621,N_12,N_528);
or U1622 (N_1622,N_1398,N_753);
and U1623 (N_1623,N_361,N_1013);
or U1624 (N_1624,N_1003,N_1135);
nand U1625 (N_1625,N_1157,N_780);
nand U1626 (N_1626,N_1064,N_507);
xnor U1627 (N_1627,N_1199,N_821);
xnor U1628 (N_1628,N_1333,N_788);
nor U1629 (N_1629,N_325,N_978);
and U1630 (N_1630,N_1311,N_771);
xor U1631 (N_1631,N_937,N_1360);
nor U1632 (N_1632,N_799,N_427);
nand U1633 (N_1633,N_181,N_342);
nand U1634 (N_1634,N_165,N_435);
or U1635 (N_1635,N_240,N_509);
and U1636 (N_1636,N_1165,N_1480);
nand U1637 (N_1637,N_1022,N_264);
xnor U1638 (N_1638,N_548,N_134);
nor U1639 (N_1639,N_1308,N_1138);
nand U1640 (N_1640,N_1484,N_98);
nor U1641 (N_1641,N_402,N_519);
nand U1642 (N_1642,N_256,N_1068);
nand U1643 (N_1643,N_1332,N_424);
and U1644 (N_1644,N_718,N_1302);
and U1645 (N_1645,N_1492,N_699);
nand U1646 (N_1646,N_837,N_1432);
nor U1647 (N_1647,N_1298,N_514);
nand U1648 (N_1648,N_929,N_1429);
nor U1649 (N_1649,N_358,N_1077);
nor U1650 (N_1650,N_218,N_817);
xnor U1651 (N_1651,N_818,N_708);
xor U1652 (N_1652,N_29,N_805);
xnor U1653 (N_1653,N_969,N_1258);
xor U1654 (N_1654,N_441,N_700);
nor U1655 (N_1655,N_71,N_57);
or U1656 (N_1656,N_596,N_904);
nand U1657 (N_1657,N_836,N_204);
xnor U1658 (N_1658,N_767,N_1293);
xor U1659 (N_1659,N_1062,N_444);
xor U1660 (N_1660,N_419,N_1414);
nand U1661 (N_1661,N_109,N_198);
xnor U1662 (N_1662,N_1066,N_1409);
nor U1663 (N_1663,N_62,N_695);
xnor U1664 (N_1664,N_551,N_197);
nor U1665 (N_1665,N_580,N_589);
xor U1666 (N_1666,N_1427,N_988);
or U1667 (N_1667,N_84,N_1009);
and U1668 (N_1668,N_955,N_909);
nand U1669 (N_1669,N_1163,N_587);
nor U1670 (N_1670,N_283,N_986);
or U1671 (N_1671,N_1300,N_1488);
xnor U1672 (N_1672,N_545,N_850);
nand U1673 (N_1673,N_800,N_1352);
and U1674 (N_1674,N_1018,N_189);
nor U1675 (N_1675,N_544,N_660);
and U1676 (N_1676,N_455,N_91);
xor U1677 (N_1677,N_483,N_1379);
xor U1678 (N_1678,N_912,N_394);
and U1679 (N_1679,N_1085,N_1454);
and U1680 (N_1680,N_170,N_1181);
xor U1681 (N_1681,N_1194,N_339);
and U1682 (N_1682,N_1147,N_565);
or U1683 (N_1683,N_1099,N_696);
xnor U1684 (N_1684,N_1148,N_1410);
nor U1685 (N_1685,N_963,N_417);
xor U1686 (N_1686,N_526,N_943);
nand U1687 (N_1687,N_99,N_1082);
xor U1688 (N_1688,N_1162,N_226);
xor U1689 (N_1689,N_445,N_618);
nor U1690 (N_1690,N_1236,N_601);
xnor U1691 (N_1691,N_894,N_368);
and U1692 (N_1692,N_1255,N_128);
nand U1693 (N_1693,N_450,N_471);
nor U1694 (N_1694,N_286,N_210);
nor U1695 (N_1695,N_10,N_1441);
nand U1696 (N_1696,N_623,N_399);
nand U1697 (N_1697,N_973,N_1122);
and U1698 (N_1698,N_268,N_925);
or U1699 (N_1699,N_843,N_703);
xnor U1700 (N_1700,N_1463,N_1177);
nand U1701 (N_1701,N_795,N_410);
nand U1702 (N_1702,N_1396,N_652);
and U1703 (N_1703,N_89,N_1069);
nand U1704 (N_1704,N_835,N_1460);
or U1705 (N_1705,N_343,N_135);
and U1706 (N_1706,N_328,N_838);
nand U1707 (N_1707,N_841,N_578);
nor U1708 (N_1708,N_698,N_56);
or U1709 (N_1709,N_290,N_107);
and U1710 (N_1710,N_1304,N_14);
or U1711 (N_1711,N_1339,N_401);
or U1712 (N_1712,N_1276,N_979);
and U1713 (N_1713,N_561,N_1098);
nor U1714 (N_1714,N_645,N_1226);
or U1715 (N_1715,N_35,N_102);
nor U1716 (N_1716,N_1456,N_321);
or U1717 (N_1717,N_1244,N_823);
xnor U1718 (N_1718,N_443,N_1239);
nand U1719 (N_1719,N_1261,N_730);
nand U1720 (N_1720,N_365,N_100);
xnor U1721 (N_1721,N_375,N_1476);
xor U1722 (N_1722,N_690,N_914);
xor U1723 (N_1723,N_55,N_1221);
xnor U1724 (N_1724,N_1101,N_748);
nand U1725 (N_1725,N_133,N_557);
nand U1726 (N_1726,N_160,N_1384);
xor U1727 (N_1727,N_768,N_808);
or U1728 (N_1728,N_178,N_840);
or U1729 (N_1729,N_472,N_1033);
xnor U1730 (N_1730,N_220,N_1301);
or U1731 (N_1731,N_33,N_1395);
and U1732 (N_1732,N_1040,N_860);
xnor U1733 (N_1733,N_575,N_738);
or U1734 (N_1734,N_999,N_319);
xor U1735 (N_1735,N_677,N_617);
xnor U1736 (N_1736,N_60,N_680);
and U1737 (N_1737,N_1136,N_675);
xor U1738 (N_1738,N_1497,N_1407);
or U1739 (N_1739,N_1291,N_731);
nand U1740 (N_1740,N_1449,N_1100);
nor U1741 (N_1741,N_631,N_1128);
nand U1742 (N_1742,N_1087,N_47);
nand U1743 (N_1743,N_1016,N_96);
or U1744 (N_1744,N_792,N_1048);
and U1745 (N_1745,N_244,N_442);
and U1746 (N_1746,N_1113,N_276);
nor U1747 (N_1747,N_604,N_1482);
and U1748 (N_1748,N_948,N_714);
xnor U1749 (N_1749,N_1183,N_889);
nand U1750 (N_1750,N_1028,N_605);
nor U1751 (N_1751,N_1171,N_196);
or U1752 (N_1752,N_734,N_284);
or U1753 (N_1753,N_1249,N_383);
nor U1754 (N_1754,N_779,N_487);
and U1755 (N_1755,N_594,N_669);
or U1756 (N_1756,N_859,N_582);
nand U1757 (N_1757,N_848,N_942);
and U1758 (N_1758,N_387,N_230);
xor U1759 (N_1759,N_1315,N_1275);
nor U1760 (N_1760,N_298,N_350);
and U1761 (N_1761,N_1092,N_407);
nand U1762 (N_1762,N_5,N_438);
or U1763 (N_1763,N_501,N_1444);
and U1764 (N_1764,N_1485,N_148);
xor U1765 (N_1765,N_478,N_871);
nor U1766 (N_1766,N_1211,N_176);
and U1767 (N_1767,N_941,N_207);
xnor U1768 (N_1768,N_213,N_972);
nor U1769 (N_1769,N_50,N_1467);
or U1770 (N_1770,N_75,N_1240);
or U1771 (N_1771,N_374,N_725);
and U1772 (N_1772,N_219,N_715);
xor U1773 (N_1773,N_1038,N_1108);
nor U1774 (N_1774,N_1189,N_239);
or U1775 (N_1775,N_18,N_1010);
nand U1776 (N_1776,N_132,N_1153);
and U1777 (N_1777,N_547,N_691);
nand U1778 (N_1778,N_1005,N_525);
or U1779 (N_1779,N_511,N_1139);
nand U1780 (N_1780,N_120,N_1434);
or U1781 (N_1781,N_1144,N_156);
xor U1782 (N_1782,N_741,N_285);
nand U1783 (N_1783,N_1054,N_388);
nand U1784 (N_1784,N_406,N_166);
or U1785 (N_1785,N_119,N_568);
and U1786 (N_1786,N_1046,N_369);
xnor U1787 (N_1787,N_349,N_185);
nor U1788 (N_1788,N_844,N_1284);
or U1789 (N_1789,N_1124,N_41);
nor U1790 (N_1790,N_1309,N_1378);
and U1791 (N_1791,N_1201,N_891);
or U1792 (N_1792,N_726,N_827);
xor U1793 (N_1793,N_847,N_1155);
nand U1794 (N_1794,N_258,N_1096);
and U1795 (N_1795,N_1461,N_1104);
nand U1796 (N_1796,N_1063,N_627);
and U1797 (N_1797,N_262,N_278);
or U1798 (N_1798,N_1202,N_260);
and U1799 (N_1799,N_1123,N_710);
nand U1800 (N_1800,N_951,N_447);
xor U1801 (N_1801,N_59,N_322);
or U1802 (N_1802,N_1206,N_569);
xor U1803 (N_1803,N_63,N_155);
nor U1804 (N_1804,N_465,N_216);
nor U1805 (N_1805,N_486,N_630);
or U1806 (N_1806,N_635,N_1341);
nor U1807 (N_1807,N_1015,N_813);
or U1808 (N_1808,N_448,N_1151);
nor U1809 (N_1809,N_508,N_1426);
and U1810 (N_1810,N_921,N_225);
xor U1811 (N_1811,N_558,N_1400);
nand U1812 (N_1812,N_1119,N_892);
nand U1813 (N_1813,N_1140,N_742);
nand U1814 (N_1814,N_19,N_168);
and U1815 (N_1815,N_1045,N_497);
nor U1816 (N_1816,N_1093,N_745);
xor U1817 (N_1817,N_857,N_867);
and U1818 (N_1818,N_92,N_974);
xor U1819 (N_1819,N_1007,N_495);
nor U1820 (N_1820,N_674,N_919);
or U1821 (N_1821,N_1075,N_1374);
nand U1822 (N_1822,N_885,N_895);
and U1823 (N_1823,N_668,N_1193);
xnor U1824 (N_1824,N_1203,N_245);
nand U1825 (N_1825,N_269,N_1002);
nor U1826 (N_1826,N_910,N_1027);
nor U1827 (N_1827,N_622,N_716);
nor U1828 (N_1828,N_7,N_657);
nand U1829 (N_1829,N_944,N_309);
or U1830 (N_1830,N_706,N_326);
or U1831 (N_1831,N_249,N_1142);
and U1832 (N_1832,N_201,N_44);
xnor U1833 (N_1833,N_145,N_794);
xnor U1834 (N_1834,N_335,N_901);
nand U1835 (N_1835,N_1442,N_1430);
xnor U1836 (N_1836,N_1196,N_595);
and U1837 (N_1837,N_429,N_1330);
or U1838 (N_1838,N_566,N_340);
or U1839 (N_1839,N_1387,N_425);
nor U1840 (N_1840,N_603,N_1473);
or U1841 (N_1841,N_0,N_496);
and U1842 (N_1842,N_517,N_233);
or U1843 (N_1843,N_1356,N_215);
nor U1844 (N_1844,N_205,N_641);
nand U1845 (N_1845,N_42,N_1447);
and U1846 (N_1846,N_1347,N_422);
or U1847 (N_1847,N_492,N_381);
and U1848 (N_1848,N_733,N_257);
nand U1849 (N_1849,N_1216,N_712);
nor U1850 (N_1850,N_1238,N_621);
and U1851 (N_1851,N_151,N_598);
and U1852 (N_1852,N_917,N_1263);
nand U1853 (N_1853,N_1462,N_1083);
nor U1854 (N_1854,N_159,N_489);
nand U1855 (N_1855,N_106,N_1403);
or U1856 (N_1856,N_1215,N_479);
nand U1857 (N_1857,N_632,N_588);
or U1858 (N_1858,N_194,N_1161);
nor U1859 (N_1859,N_490,N_1373);
and U1860 (N_1860,N_1389,N_1477);
nor U1861 (N_1861,N_299,N_1186);
nor U1862 (N_1862,N_314,N_1175);
or U1863 (N_1863,N_182,N_761);
nor U1864 (N_1864,N_1393,N_1017);
nand U1865 (N_1865,N_206,N_1404);
or U1866 (N_1866,N_78,N_164);
nand U1867 (N_1867,N_584,N_856);
or U1868 (N_1868,N_740,N_65);
nor U1869 (N_1869,N_1350,N_957);
xnor U1870 (N_1870,N_923,N_751);
nor U1871 (N_1871,N_274,N_704);
or U1872 (N_1872,N_1408,N_1117);
and U1873 (N_1873,N_1268,N_689);
nand U1874 (N_1874,N_318,N_1231);
and U1875 (N_1875,N_681,N_54);
nand U1876 (N_1876,N_345,N_659);
and U1877 (N_1877,N_93,N_4);
or U1878 (N_1878,N_1489,N_1490);
and U1879 (N_1879,N_376,N_147);
xor U1880 (N_1880,N_1375,N_327);
nor U1881 (N_1881,N_713,N_577);
and U1882 (N_1882,N_993,N_1422);
nand U1883 (N_1883,N_179,N_1118);
or U1884 (N_1884,N_432,N_579);
xor U1885 (N_1885,N_391,N_1125);
or U1886 (N_1886,N_952,N_760);
xnor U1887 (N_1887,N_958,N_829);
nand U1888 (N_1888,N_1001,N_1152);
xor U1889 (N_1889,N_682,N_169);
or U1890 (N_1890,N_820,N_1495);
nor U1891 (N_1891,N_553,N_15);
xor U1892 (N_1892,N_983,N_639);
xnor U1893 (N_1893,N_39,N_1320);
nand U1894 (N_1894,N_1328,N_754);
nor U1895 (N_1895,N_37,N_1044);
and U1896 (N_1896,N_612,N_73);
nand U1897 (N_1897,N_241,N_246);
xor U1898 (N_1898,N_787,N_423);
nor U1899 (N_1899,N_317,N_1306);
nand U1900 (N_1900,N_571,N_146);
and U1901 (N_1901,N_998,N_301);
or U1902 (N_1902,N_1228,N_1034);
and U1903 (N_1903,N_1466,N_1278);
and U1904 (N_1904,N_332,N_1438);
xor U1905 (N_1905,N_1019,N_778);
and U1906 (N_1906,N_398,N_1381);
nand U1907 (N_1907,N_300,N_1322);
or U1908 (N_1908,N_1361,N_353);
and U1909 (N_1909,N_263,N_546);
and U1910 (N_1910,N_707,N_724);
nand U1911 (N_1911,N_886,N_729);
and U1912 (N_1912,N_721,N_774);
nand U1913 (N_1913,N_150,N_252);
nand U1914 (N_1914,N_853,N_1424);
xnor U1915 (N_1915,N_116,N_784);
nand U1916 (N_1916,N_158,N_1073);
nand U1917 (N_1917,N_530,N_798);
and U1918 (N_1918,N_540,N_1289);
xnor U1919 (N_1919,N_554,N_1498);
and U1920 (N_1920,N_400,N_949);
xor U1921 (N_1921,N_1090,N_940);
and U1922 (N_1922,N_392,N_251);
or U1923 (N_1923,N_572,N_334);
nor U1924 (N_1924,N_1281,N_288);
or U1925 (N_1925,N_1030,N_242);
xor U1926 (N_1926,N_1250,N_458);
nand U1927 (N_1927,N_1059,N_656);
nor U1928 (N_1928,N_826,N_819);
or U1929 (N_1929,N_1200,N_538);
nor U1930 (N_1930,N_222,N_38);
and U1931 (N_1931,N_877,N_533);
or U1932 (N_1932,N_905,N_769);
or U1933 (N_1933,N_590,N_524);
nor U1934 (N_1934,N_11,N_74);
and U1935 (N_1935,N_302,N_683);
xor U1936 (N_1936,N_591,N_1070);
nand U1937 (N_1937,N_1344,N_746);
and U1938 (N_1938,N_685,N_446);
xnor U1939 (N_1939,N_995,N_732);
and U1940 (N_1940,N_1470,N_1217);
xnor U1941 (N_1941,N_114,N_1411);
and U1942 (N_1942,N_884,N_351);
and U1943 (N_1943,N_282,N_259);
or U1944 (N_1944,N_1246,N_154);
and U1945 (N_1945,N_1262,N_371);
xnor U1946 (N_1946,N_1264,N_806);
or U1947 (N_1947,N_1094,N_292);
nand U1948 (N_1948,N_1317,N_360);
xnor U1949 (N_1949,N_272,N_532);
nand U1950 (N_1950,N_928,N_386);
nand U1951 (N_1951,N_127,N_323);
and U1952 (N_1952,N_480,N_834);
nand U1953 (N_1953,N_968,N_1310);
and U1954 (N_1954,N_27,N_475);
and U1955 (N_1955,N_1209,N_136);
and U1956 (N_1956,N_815,N_1042);
or U1957 (N_1957,N_1224,N_1406);
and U1958 (N_1958,N_473,N_188);
and U1959 (N_1959,N_266,N_709);
nand U1960 (N_1960,N_1149,N_755);
and U1961 (N_1961,N_315,N_1294);
nand U1962 (N_1962,N_1208,N_177);
xor U1963 (N_1963,N_1391,N_228);
or U1964 (N_1964,N_80,N_1334);
or U1965 (N_1965,N_1095,N_453);
and U1966 (N_1966,N_161,N_662);
and U1967 (N_1967,N_1287,N_53);
and U1968 (N_1968,N_130,N_209);
xnor U1969 (N_1969,N_3,N_131);
xnor U1970 (N_1970,N_1428,N_550);
and U1971 (N_1971,N_1120,N_469);
and U1972 (N_1972,N_644,N_643);
and U1973 (N_1973,N_267,N_1052);
or U1974 (N_1974,N_757,N_1021);
xor U1975 (N_1975,N_468,N_1130);
or U1976 (N_1976,N_543,N_846);
xnor U1977 (N_1977,N_366,N_470);
and U1978 (N_1978,N_946,N_839);
nor U1979 (N_1979,N_920,N_1180);
nor U1980 (N_1980,N_312,N_965);
nor U1981 (N_1981,N_976,N_1198);
nand U1982 (N_1982,N_1032,N_1072);
xnor U1983 (N_1983,N_822,N_1058);
or U1984 (N_1984,N_854,N_1220);
nor U1985 (N_1985,N_1272,N_752);
nand U1986 (N_1986,N_1296,N_1036);
xnor U1987 (N_1987,N_1227,N_1167);
and U1988 (N_1988,N_115,N_397);
xnor U1989 (N_1989,N_1182,N_964);
xor U1990 (N_1990,N_440,N_87);
and U1991 (N_1991,N_433,N_950);
nand U1992 (N_1992,N_770,N_356);
xor U1993 (N_1993,N_1420,N_1401);
or U1994 (N_1994,N_1325,N_549);
xor U1995 (N_1995,N_1313,N_1299);
nor U1996 (N_1996,N_1443,N_227);
nand U1997 (N_1997,N_939,N_1105);
and U1998 (N_1998,N_555,N_25);
nor U1999 (N_1999,N_1365,N_1109);
nor U2000 (N_2000,N_1218,N_336);
nor U2001 (N_2001,N_1499,N_1260);
nand U2002 (N_2002,N_261,N_199);
or U2003 (N_2003,N_1006,N_651);
or U2004 (N_2004,N_875,N_384);
nor U2005 (N_2005,N_420,N_804);
or U2006 (N_2006,N_1368,N_294);
nand U2007 (N_2007,N_1331,N_221);
nand U2008 (N_2008,N_395,N_673);
or U2009 (N_2009,N_1446,N_556);
and U2010 (N_2010,N_1279,N_989);
nand U2011 (N_2011,N_516,N_101);
and U2012 (N_2012,N_933,N_1158);
or U2013 (N_2013,N_1031,N_833);
and U2014 (N_2014,N_1115,N_1230);
or U2015 (N_2015,N_518,N_1103);
nand U2016 (N_2016,N_649,N_625);
xor U2017 (N_2017,N_32,N_890);
and U2018 (N_2018,N_389,N_842);
nor U2019 (N_2019,N_1364,N_1357);
or U2020 (N_2020,N_110,N_1188);
nor U2021 (N_2021,N_1267,N_405);
and U2022 (N_2022,N_1,N_1283);
nand U2023 (N_2023,N_16,N_722);
xor U2024 (N_2024,N_237,N_932);
nand U2025 (N_2025,N_1288,N_640);
xnor U2026 (N_2026,N_975,N_1354);
and U2027 (N_2027,N_67,N_994);
xnor U2028 (N_2028,N_747,N_304);
nor U2029 (N_2029,N_1318,N_868);
nand U2030 (N_2030,N_108,N_521);
nand U2031 (N_2031,N_739,N_235);
and U2032 (N_2032,N_491,N_1483);
xnor U2033 (N_2033,N_831,N_499);
or U2034 (N_2034,N_1222,N_1205);
xnor U2035 (N_2035,N_1257,N_665);
xor U2036 (N_2036,N_174,N_666);
nand U2037 (N_2037,N_559,N_414);
and U2038 (N_2038,N_1273,N_1295);
nand U2039 (N_2039,N_1270,N_1363);
xor U2040 (N_2040,N_1061,N_124);
xnor U2041 (N_2041,N_1303,N_1385);
xnor U2042 (N_2042,N_773,N_1081);
nor U2043 (N_2043,N_807,N_927);
or U2044 (N_2044,N_574,N_1397);
nor U2045 (N_2045,N_504,N_1210);
nor U2046 (N_2046,N_870,N_1418);
nor U2047 (N_2047,N_477,N_1359);
xnor U2048 (N_2048,N_493,N_879);
xnor U2049 (N_2049,N_1362,N_736);
or U2050 (N_2050,N_766,N_935);
nand U2051 (N_2051,N_217,N_984);
nand U2052 (N_2052,N_1229,N_66);
xnor U2053 (N_2053,N_956,N_541);
and U2054 (N_2054,N_1011,N_1050);
nand U2055 (N_2055,N_671,N_382);
or U2056 (N_2056,N_348,N_121);
xor U2057 (N_2057,N_412,N_610);
and U2058 (N_2058,N_1388,N_105);
and U2059 (N_2059,N_34,N_1174);
nand U2060 (N_2060,N_576,N_1412);
or U2061 (N_2061,N_1345,N_280);
xor U2062 (N_2062,N_436,N_830);
nor U2063 (N_2063,N_1219,N_814);
and U2064 (N_2064,N_1133,N_1247);
nand U2065 (N_2065,N_1358,N_642);
or U2066 (N_2066,N_764,N_1197);
and U2067 (N_2067,N_126,N_789);
xor U2068 (N_2068,N_1340,N_393);
xnor U2069 (N_2069,N_783,N_255);
nor U2070 (N_2070,N_88,N_797);
or U2071 (N_2071,N_380,N_139);
nand U2072 (N_2072,N_86,N_1286);
or U2073 (N_2073,N_187,N_85);
nand U2074 (N_2074,N_1020,N_411);
xnor U2075 (N_2075,N_363,N_782);
nor U2076 (N_2076,N_1145,N_1214);
nand U2077 (N_2077,N_803,N_1392);
nand U2078 (N_2078,N_796,N_599);
xor U2079 (N_2079,N_1102,N_1156);
xnor U2080 (N_2080,N_749,N_1134);
nand U2081 (N_2081,N_1326,N_289);
nor U2082 (N_2082,N_1008,N_602);
and U2083 (N_2083,N_122,N_1168);
and U2084 (N_2084,N_502,N_77);
or U2085 (N_2085,N_586,N_2);
and U2086 (N_2086,N_980,N_560);
nand U2087 (N_2087,N_1419,N_522);
and U2088 (N_2088,N_460,N_1112);
nor U2089 (N_2089,N_1141,N_934);
or U2090 (N_2090,N_1367,N_1382);
nand U2091 (N_2091,N_1324,N_378);
nand U2092 (N_2092,N_985,N_1464);
and U2093 (N_2093,N_476,N_203);
nand U2094 (N_2094,N_451,N_930);
nand U2095 (N_2095,N_51,N_585);
and U2096 (N_2096,N_670,N_667);
nand U2097 (N_2097,N_997,N_370);
nor U2098 (N_2098,N_129,N_982);
nand U2099 (N_2099,N_1166,N_865);
nor U2100 (N_2100,N_362,N_1029);
xor U2101 (N_2101,N_581,N_776);
xor U2102 (N_2102,N_900,N_931);
and U2103 (N_2103,N_1415,N_687);
and U2104 (N_2104,N_1431,N_1126);
xor U2105 (N_2105,N_485,N_991);
and U2106 (N_2106,N_1086,N_247);
nand U2107 (N_2107,N_626,N_186);
xnor U2108 (N_2108,N_449,N_911);
or U2109 (N_2109,N_1423,N_416);
and U2110 (N_2110,N_162,N_6);
xnor U2111 (N_2111,N_758,N_1355);
and U2112 (N_2112,N_352,N_390);
nand U2113 (N_2113,N_570,N_1491);
nand U2114 (N_2114,N_24,N_190);
xor U2115 (N_2115,N_791,N_1348);
or U2116 (N_2116,N_1435,N_1277);
and U2117 (N_2117,N_872,N_510);
xor U2118 (N_2118,N_254,N_26);
nand U2119 (N_2119,N_183,N_426);
nand U2120 (N_2120,N_1131,N_1343);
nor U2121 (N_2121,N_421,N_811);
or U2122 (N_2122,N_825,N_536);
xnor U2123 (N_2123,N_620,N_781);
nor U2124 (N_2124,N_1335,N_1338);
nand U2125 (N_2125,N_1323,N_653);
xnor U2126 (N_2126,N_1053,N_1337);
xor U2127 (N_2127,N_611,N_567);
xnor U2128 (N_2128,N_523,N_202);
and U2129 (N_2129,N_467,N_1060);
nor U2130 (N_2130,N_1282,N_793);
nor U2131 (N_2131,N_1057,N_1457);
and U2132 (N_2132,N_852,N_529);
nor U2133 (N_2133,N_184,N_878);
and U2134 (N_2134,N_866,N_22);
nor U2135 (N_2135,N_899,N_763);
nor U2136 (N_2136,N_153,N_1394);
nand U2137 (N_2137,N_542,N_359);
nor U2138 (N_2138,N_1297,N_457);
nor U2139 (N_2139,N_977,N_936);
or U2140 (N_2140,N_113,N_1383);
xor U2141 (N_2141,N_311,N_1253);
and U2142 (N_2142,N_1259,N_564);
or U2143 (N_2143,N_208,N_45);
or U2144 (N_2144,N_893,N_971);
or U2145 (N_2145,N_1266,N_686);
xnor U2146 (N_2146,N_307,N_593);
nor U2147 (N_2147,N_355,N_1305);
xor U2148 (N_2148,N_609,N_786);
or U2149 (N_2149,N_200,N_1097);
and U2150 (N_2150,N_265,N_597);
xnor U2151 (N_2151,N_503,N_802);
nand U2152 (N_2152,N_212,N_36);
nand U2153 (N_2153,N_809,N_232);
and U2154 (N_2154,N_1451,N_1026);
xnor U2155 (N_2155,N_1437,N_1212);
xor U2156 (N_2156,N_592,N_970);
nand U2157 (N_2157,N_103,N_1290);
xnor U2158 (N_2158,N_229,N_1448);
nand U2159 (N_2159,N_1292,N_1065);
nand U2160 (N_2160,N_1496,N_43);
xor U2161 (N_2161,N_527,N_1041);
and U2162 (N_2162,N_1479,N_873);
nor U2163 (N_2163,N_76,N_960);
and U2164 (N_2164,N_1106,N_1372);
xnor U2165 (N_2165,N_1121,N_663);
or U2166 (N_2166,N_634,N_688);
nand U2167 (N_2167,N_535,N_1481);
and U2168 (N_2168,N_1450,N_281);
and U2169 (N_2169,N_23,N_111);
nor U2170 (N_2170,N_347,N_874);
or U2171 (N_2171,N_723,N_1091);
xnor U2172 (N_2172,N_762,N_1204);
nor U2173 (N_2173,N_1468,N_1319);
or U2174 (N_2174,N_1179,N_1114);
xor U2175 (N_2175,N_913,N_1089);
xor U2176 (N_2176,N_439,N_961);
nand U2177 (N_2177,N_275,N_1425);
and U2178 (N_2178,N_1159,N_1150);
or U2179 (N_2179,N_341,N_291);
xnor U2180 (N_2180,N_428,N_515);
nor U2181 (N_2181,N_777,N_1494);
and U2182 (N_2182,N_1370,N_990);
or U2183 (N_2183,N_520,N_824);
or U2184 (N_2184,N_310,N_474);
nor U2185 (N_2185,N_72,N_1146);
nand U2186 (N_2186,N_916,N_117);
and U2187 (N_2187,N_1160,N_655);
xor U2188 (N_2188,N_431,N_1254);
or U2189 (N_2189,N_195,N_144);
nor U2190 (N_2190,N_861,N_357);
xor U2191 (N_2191,N_1243,N_1056);
or U2192 (N_2192,N_684,N_775);
or U2193 (N_2193,N_58,N_1433);
and U2194 (N_2194,N_648,N_772);
xnor U2195 (N_2195,N_926,N_48);
nor U2196 (N_2196,N_531,N_1405);
and U2197 (N_2197,N_1242,N_1051);
nand U2198 (N_2198,N_915,N_583);
nand U2199 (N_2199,N_1184,N_537);
xor U2200 (N_2200,N_1327,N_180);
xnor U2201 (N_2201,N_1071,N_143);
and U2202 (N_2202,N_1055,N_461);
and U2203 (N_2203,N_1353,N_1245);
xnor U2204 (N_2204,N_987,N_1078);
xor U2205 (N_2205,N_862,N_1225);
nand U2206 (N_2206,N_1195,N_552);
nor U2207 (N_2207,N_637,N_672);
and U2208 (N_2208,N_881,N_633);
nand U2209 (N_2209,N_344,N_316);
nand U2210 (N_2210,N_1252,N_908);
nand U2211 (N_2211,N_21,N_456);
xor U2212 (N_2212,N_224,N_996);
xnor U2213 (N_2213,N_1235,N_142);
or U2214 (N_2214,N_832,N_271);
nand U2215 (N_2215,N_624,N_1110);
and U2216 (N_2216,N_273,N_379);
or U2217 (N_2217,N_717,N_629);
nand U2218 (N_2218,N_1025,N_466);
xor U2219 (N_2219,N_896,N_1233);
nand U2220 (N_2220,N_173,N_1321);
nor U2221 (N_2221,N_661,N_324);
or U2222 (N_2222,N_277,N_1376);
nand U2223 (N_2223,N_506,N_452);
nand U2224 (N_2224,N_463,N_279);
or U2225 (N_2225,N_248,N_869);
and U2226 (N_2226,N_83,N_1366);
xor U2227 (N_2227,N_1111,N_97);
xor U2228 (N_2228,N_1234,N_902);
nand U2229 (N_2229,N_1377,N_614);
or U2230 (N_2230,N_415,N_500);
xnor U2231 (N_2231,N_1469,N_1421);
and U2232 (N_2232,N_992,N_364);
and U2233 (N_2233,N_303,N_459);
and U2234 (N_2234,N_253,N_512);
or U2235 (N_2235,N_1079,N_678);
nand U2236 (N_2236,N_1207,N_320);
xor U2237 (N_2237,N_863,N_735);
nor U2238 (N_2238,N_1280,N_498);
nand U2239 (N_2239,N_293,N_907);
xor U2240 (N_2240,N_638,N_1172);
or U2241 (N_2241,N_418,N_816);
and U2242 (N_2242,N_270,N_855);
or U2243 (N_2243,N_95,N_1023);
nor U2244 (N_2244,N_1439,N_330);
or U2245 (N_2245,N_396,N_1178);
nor U2246 (N_2246,N_464,N_20);
and U2247 (N_2247,N_966,N_125);
xor U2248 (N_2248,N_981,N_711);
nor U2249 (N_2249,N_694,N_513);
nor U2250 (N_2250,N_754,N_673);
nand U2251 (N_2251,N_996,N_169);
nor U2252 (N_2252,N_964,N_952);
and U2253 (N_2253,N_1402,N_660);
or U2254 (N_2254,N_262,N_692);
xor U2255 (N_2255,N_1277,N_690);
and U2256 (N_2256,N_1316,N_1224);
or U2257 (N_2257,N_649,N_354);
or U2258 (N_2258,N_602,N_1193);
and U2259 (N_2259,N_681,N_843);
nand U2260 (N_2260,N_62,N_1198);
xnor U2261 (N_2261,N_1336,N_261);
nor U2262 (N_2262,N_566,N_519);
xnor U2263 (N_2263,N_1021,N_369);
nor U2264 (N_2264,N_1023,N_846);
nand U2265 (N_2265,N_805,N_729);
nand U2266 (N_2266,N_843,N_545);
nor U2267 (N_2267,N_1258,N_340);
and U2268 (N_2268,N_701,N_897);
or U2269 (N_2269,N_1424,N_389);
or U2270 (N_2270,N_434,N_715);
xor U2271 (N_2271,N_896,N_1372);
nor U2272 (N_2272,N_61,N_283);
and U2273 (N_2273,N_689,N_193);
or U2274 (N_2274,N_1084,N_75);
xnor U2275 (N_2275,N_729,N_1311);
nand U2276 (N_2276,N_556,N_376);
xor U2277 (N_2277,N_127,N_574);
nor U2278 (N_2278,N_679,N_158);
nand U2279 (N_2279,N_269,N_984);
nand U2280 (N_2280,N_1476,N_1408);
xor U2281 (N_2281,N_1337,N_1036);
nand U2282 (N_2282,N_511,N_243);
nand U2283 (N_2283,N_1492,N_657);
xor U2284 (N_2284,N_268,N_1483);
and U2285 (N_2285,N_1281,N_815);
nor U2286 (N_2286,N_369,N_886);
and U2287 (N_2287,N_577,N_1398);
nand U2288 (N_2288,N_709,N_776);
and U2289 (N_2289,N_96,N_1072);
nor U2290 (N_2290,N_1028,N_202);
and U2291 (N_2291,N_1083,N_39);
or U2292 (N_2292,N_799,N_645);
nand U2293 (N_2293,N_1046,N_637);
and U2294 (N_2294,N_1379,N_776);
xor U2295 (N_2295,N_1315,N_459);
xor U2296 (N_2296,N_978,N_672);
nor U2297 (N_2297,N_875,N_270);
and U2298 (N_2298,N_20,N_657);
nor U2299 (N_2299,N_675,N_351);
xor U2300 (N_2300,N_640,N_629);
nor U2301 (N_2301,N_806,N_1076);
or U2302 (N_2302,N_578,N_67);
nor U2303 (N_2303,N_1445,N_1118);
and U2304 (N_2304,N_1072,N_250);
nand U2305 (N_2305,N_1361,N_46);
xnor U2306 (N_2306,N_728,N_1497);
or U2307 (N_2307,N_1446,N_741);
nor U2308 (N_2308,N_1234,N_1268);
nand U2309 (N_2309,N_1188,N_554);
xor U2310 (N_2310,N_152,N_474);
and U2311 (N_2311,N_1083,N_1125);
xnor U2312 (N_2312,N_312,N_1146);
nand U2313 (N_2313,N_955,N_979);
or U2314 (N_2314,N_162,N_251);
and U2315 (N_2315,N_414,N_340);
and U2316 (N_2316,N_1363,N_1154);
and U2317 (N_2317,N_69,N_1132);
xnor U2318 (N_2318,N_841,N_919);
and U2319 (N_2319,N_307,N_697);
and U2320 (N_2320,N_1435,N_1043);
xnor U2321 (N_2321,N_804,N_1475);
or U2322 (N_2322,N_445,N_938);
or U2323 (N_2323,N_257,N_695);
and U2324 (N_2324,N_278,N_364);
nand U2325 (N_2325,N_1065,N_155);
or U2326 (N_2326,N_79,N_1151);
xnor U2327 (N_2327,N_826,N_216);
xnor U2328 (N_2328,N_173,N_1159);
nor U2329 (N_2329,N_720,N_771);
xnor U2330 (N_2330,N_117,N_1349);
nand U2331 (N_2331,N_1356,N_1379);
xnor U2332 (N_2332,N_530,N_323);
nor U2333 (N_2333,N_734,N_1338);
or U2334 (N_2334,N_312,N_1285);
or U2335 (N_2335,N_623,N_1104);
and U2336 (N_2336,N_1137,N_309);
and U2337 (N_2337,N_226,N_1094);
nand U2338 (N_2338,N_687,N_571);
xor U2339 (N_2339,N_1181,N_709);
nor U2340 (N_2340,N_1074,N_1484);
and U2341 (N_2341,N_484,N_1111);
xor U2342 (N_2342,N_1019,N_489);
nand U2343 (N_2343,N_786,N_207);
or U2344 (N_2344,N_714,N_987);
nand U2345 (N_2345,N_871,N_1096);
nand U2346 (N_2346,N_1455,N_657);
xnor U2347 (N_2347,N_1354,N_414);
nand U2348 (N_2348,N_601,N_915);
and U2349 (N_2349,N_1374,N_19);
xnor U2350 (N_2350,N_691,N_19);
nor U2351 (N_2351,N_190,N_396);
or U2352 (N_2352,N_1106,N_3);
and U2353 (N_2353,N_1188,N_501);
xnor U2354 (N_2354,N_226,N_1338);
nor U2355 (N_2355,N_785,N_737);
and U2356 (N_2356,N_1081,N_326);
or U2357 (N_2357,N_1427,N_33);
nand U2358 (N_2358,N_1491,N_510);
nor U2359 (N_2359,N_860,N_457);
or U2360 (N_2360,N_643,N_401);
or U2361 (N_2361,N_335,N_615);
and U2362 (N_2362,N_666,N_432);
xor U2363 (N_2363,N_112,N_71);
nor U2364 (N_2364,N_734,N_1347);
xor U2365 (N_2365,N_832,N_798);
and U2366 (N_2366,N_605,N_1020);
nand U2367 (N_2367,N_862,N_1250);
nor U2368 (N_2368,N_808,N_331);
or U2369 (N_2369,N_95,N_938);
xnor U2370 (N_2370,N_859,N_226);
and U2371 (N_2371,N_597,N_44);
nor U2372 (N_2372,N_389,N_908);
or U2373 (N_2373,N_1382,N_813);
nor U2374 (N_2374,N_547,N_1247);
nand U2375 (N_2375,N_1392,N_610);
nor U2376 (N_2376,N_983,N_1319);
and U2377 (N_2377,N_261,N_1064);
nor U2378 (N_2378,N_1294,N_870);
or U2379 (N_2379,N_551,N_491);
nand U2380 (N_2380,N_107,N_1355);
and U2381 (N_2381,N_1058,N_515);
nand U2382 (N_2382,N_1411,N_1185);
xnor U2383 (N_2383,N_241,N_387);
nor U2384 (N_2384,N_901,N_962);
nand U2385 (N_2385,N_906,N_318);
xor U2386 (N_2386,N_102,N_532);
or U2387 (N_2387,N_1017,N_685);
or U2388 (N_2388,N_126,N_662);
xor U2389 (N_2389,N_687,N_948);
and U2390 (N_2390,N_186,N_191);
or U2391 (N_2391,N_204,N_255);
or U2392 (N_2392,N_631,N_862);
xor U2393 (N_2393,N_929,N_685);
xnor U2394 (N_2394,N_1130,N_653);
nor U2395 (N_2395,N_403,N_1105);
or U2396 (N_2396,N_1149,N_233);
or U2397 (N_2397,N_1033,N_1032);
and U2398 (N_2398,N_21,N_202);
nor U2399 (N_2399,N_88,N_1007);
or U2400 (N_2400,N_194,N_586);
or U2401 (N_2401,N_638,N_1128);
and U2402 (N_2402,N_771,N_658);
or U2403 (N_2403,N_216,N_676);
nor U2404 (N_2404,N_1326,N_11);
or U2405 (N_2405,N_1245,N_1040);
xor U2406 (N_2406,N_1253,N_593);
nor U2407 (N_2407,N_1201,N_1102);
or U2408 (N_2408,N_673,N_369);
nor U2409 (N_2409,N_592,N_719);
nand U2410 (N_2410,N_901,N_1434);
xnor U2411 (N_2411,N_90,N_1008);
xnor U2412 (N_2412,N_1020,N_1375);
nand U2413 (N_2413,N_570,N_1478);
nor U2414 (N_2414,N_457,N_651);
nor U2415 (N_2415,N_1001,N_510);
nand U2416 (N_2416,N_1032,N_1096);
or U2417 (N_2417,N_1149,N_592);
nor U2418 (N_2418,N_673,N_1111);
nand U2419 (N_2419,N_939,N_1380);
xnor U2420 (N_2420,N_13,N_251);
nor U2421 (N_2421,N_964,N_1404);
nor U2422 (N_2422,N_161,N_243);
xnor U2423 (N_2423,N_36,N_513);
nand U2424 (N_2424,N_1149,N_112);
and U2425 (N_2425,N_496,N_455);
or U2426 (N_2426,N_238,N_1050);
nand U2427 (N_2427,N_491,N_1038);
and U2428 (N_2428,N_400,N_178);
nor U2429 (N_2429,N_373,N_446);
nor U2430 (N_2430,N_77,N_1078);
or U2431 (N_2431,N_1292,N_1425);
or U2432 (N_2432,N_1485,N_774);
xor U2433 (N_2433,N_162,N_781);
xor U2434 (N_2434,N_765,N_1021);
nor U2435 (N_2435,N_1229,N_1432);
xor U2436 (N_2436,N_1395,N_824);
and U2437 (N_2437,N_721,N_913);
nand U2438 (N_2438,N_15,N_42);
or U2439 (N_2439,N_378,N_1416);
nor U2440 (N_2440,N_1249,N_1245);
and U2441 (N_2441,N_1189,N_258);
xnor U2442 (N_2442,N_1420,N_668);
and U2443 (N_2443,N_1187,N_330);
and U2444 (N_2444,N_475,N_1296);
xnor U2445 (N_2445,N_1271,N_1216);
and U2446 (N_2446,N_1068,N_1102);
nor U2447 (N_2447,N_1375,N_735);
nand U2448 (N_2448,N_1282,N_61);
nor U2449 (N_2449,N_1374,N_866);
nor U2450 (N_2450,N_513,N_1427);
nor U2451 (N_2451,N_476,N_678);
xor U2452 (N_2452,N_1457,N_910);
xor U2453 (N_2453,N_898,N_1157);
nand U2454 (N_2454,N_172,N_1138);
nand U2455 (N_2455,N_808,N_502);
and U2456 (N_2456,N_868,N_591);
and U2457 (N_2457,N_877,N_695);
xor U2458 (N_2458,N_369,N_256);
or U2459 (N_2459,N_1306,N_1240);
and U2460 (N_2460,N_688,N_1217);
or U2461 (N_2461,N_1046,N_683);
xnor U2462 (N_2462,N_481,N_793);
nor U2463 (N_2463,N_9,N_556);
and U2464 (N_2464,N_925,N_812);
xnor U2465 (N_2465,N_540,N_180);
xor U2466 (N_2466,N_1306,N_257);
or U2467 (N_2467,N_863,N_1119);
nand U2468 (N_2468,N_759,N_856);
nand U2469 (N_2469,N_630,N_20);
xnor U2470 (N_2470,N_1097,N_1169);
nor U2471 (N_2471,N_878,N_1228);
nand U2472 (N_2472,N_1283,N_1424);
or U2473 (N_2473,N_154,N_565);
and U2474 (N_2474,N_902,N_151);
or U2475 (N_2475,N_732,N_1184);
nand U2476 (N_2476,N_1448,N_1491);
or U2477 (N_2477,N_1386,N_569);
and U2478 (N_2478,N_1391,N_118);
and U2479 (N_2479,N_999,N_1072);
nand U2480 (N_2480,N_1307,N_602);
or U2481 (N_2481,N_811,N_329);
nand U2482 (N_2482,N_820,N_761);
or U2483 (N_2483,N_1016,N_1386);
xnor U2484 (N_2484,N_587,N_350);
xor U2485 (N_2485,N_1284,N_1083);
and U2486 (N_2486,N_380,N_773);
nand U2487 (N_2487,N_792,N_19);
xor U2488 (N_2488,N_384,N_80);
or U2489 (N_2489,N_699,N_564);
and U2490 (N_2490,N_527,N_718);
xor U2491 (N_2491,N_1311,N_145);
or U2492 (N_2492,N_832,N_1240);
nor U2493 (N_2493,N_529,N_842);
and U2494 (N_2494,N_1316,N_1116);
nor U2495 (N_2495,N_710,N_228);
nor U2496 (N_2496,N_660,N_602);
or U2497 (N_2497,N_1093,N_606);
or U2498 (N_2498,N_1197,N_685);
or U2499 (N_2499,N_1112,N_1450);
nand U2500 (N_2500,N_908,N_646);
xor U2501 (N_2501,N_971,N_720);
nor U2502 (N_2502,N_796,N_514);
xor U2503 (N_2503,N_257,N_131);
or U2504 (N_2504,N_586,N_255);
or U2505 (N_2505,N_431,N_471);
nor U2506 (N_2506,N_810,N_433);
nand U2507 (N_2507,N_141,N_443);
nor U2508 (N_2508,N_260,N_1499);
xnor U2509 (N_2509,N_967,N_810);
xor U2510 (N_2510,N_1436,N_582);
nand U2511 (N_2511,N_667,N_1124);
xor U2512 (N_2512,N_1089,N_938);
nor U2513 (N_2513,N_268,N_1075);
or U2514 (N_2514,N_653,N_900);
xor U2515 (N_2515,N_511,N_245);
or U2516 (N_2516,N_508,N_693);
and U2517 (N_2517,N_212,N_181);
xnor U2518 (N_2518,N_55,N_1202);
and U2519 (N_2519,N_459,N_126);
and U2520 (N_2520,N_818,N_1344);
nor U2521 (N_2521,N_916,N_938);
nand U2522 (N_2522,N_502,N_1055);
and U2523 (N_2523,N_100,N_1417);
nand U2524 (N_2524,N_421,N_584);
nand U2525 (N_2525,N_1129,N_1403);
and U2526 (N_2526,N_341,N_188);
or U2527 (N_2527,N_174,N_1052);
and U2528 (N_2528,N_939,N_1324);
nor U2529 (N_2529,N_339,N_1165);
xnor U2530 (N_2530,N_420,N_1369);
xnor U2531 (N_2531,N_1362,N_383);
or U2532 (N_2532,N_1068,N_767);
nor U2533 (N_2533,N_467,N_217);
and U2534 (N_2534,N_1192,N_1223);
or U2535 (N_2535,N_1021,N_232);
nand U2536 (N_2536,N_1494,N_706);
nand U2537 (N_2537,N_481,N_1289);
nor U2538 (N_2538,N_1404,N_1332);
and U2539 (N_2539,N_895,N_667);
and U2540 (N_2540,N_809,N_1016);
and U2541 (N_2541,N_947,N_1301);
nor U2542 (N_2542,N_359,N_472);
or U2543 (N_2543,N_1018,N_252);
nor U2544 (N_2544,N_1228,N_360);
or U2545 (N_2545,N_914,N_1443);
or U2546 (N_2546,N_679,N_12);
nor U2547 (N_2547,N_1469,N_982);
xor U2548 (N_2548,N_774,N_1452);
nand U2549 (N_2549,N_1273,N_1075);
xnor U2550 (N_2550,N_932,N_91);
or U2551 (N_2551,N_448,N_841);
nand U2552 (N_2552,N_558,N_938);
xnor U2553 (N_2553,N_1221,N_218);
and U2554 (N_2554,N_1300,N_1128);
xor U2555 (N_2555,N_603,N_1239);
and U2556 (N_2556,N_1125,N_400);
or U2557 (N_2557,N_1135,N_270);
or U2558 (N_2558,N_309,N_450);
or U2559 (N_2559,N_438,N_429);
nor U2560 (N_2560,N_549,N_276);
and U2561 (N_2561,N_1153,N_1170);
and U2562 (N_2562,N_1337,N_313);
nor U2563 (N_2563,N_1272,N_959);
and U2564 (N_2564,N_1156,N_1279);
nand U2565 (N_2565,N_589,N_1474);
nand U2566 (N_2566,N_138,N_257);
nand U2567 (N_2567,N_331,N_579);
and U2568 (N_2568,N_543,N_704);
and U2569 (N_2569,N_1393,N_342);
xnor U2570 (N_2570,N_1012,N_440);
xnor U2571 (N_2571,N_638,N_142);
or U2572 (N_2572,N_1325,N_415);
nor U2573 (N_2573,N_1485,N_383);
xnor U2574 (N_2574,N_624,N_1278);
xor U2575 (N_2575,N_794,N_1258);
nor U2576 (N_2576,N_1238,N_299);
nand U2577 (N_2577,N_498,N_981);
and U2578 (N_2578,N_1224,N_1071);
xor U2579 (N_2579,N_1098,N_437);
nand U2580 (N_2580,N_1149,N_1197);
nor U2581 (N_2581,N_1035,N_60);
and U2582 (N_2582,N_517,N_842);
and U2583 (N_2583,N_169,N_1311);
or U2584 (N_2584,N_1303,N_1269);
or U2585 (N_2585,N_861,N_1283);
nor U2586 (N_2586,N_1264,N_560);
xor U2587 (N_2587,N_199,N_1128);
nand U2588 (N_2588,N_31,N_847);
and U2589 (N_2589,N_21,N_628);
xnor U2590 (N_2590,N_481,N_231);
and U2591 (N_2591,N_57,N_724);
nand U2592 (N_2592,N_828,N_265);
or U2593 (N_2593,N_697,N_443);
or U2594 (N_2594,N_1320,N_839);
and U2595 (N_2595,N_1325,N_1216);
xnor U2596 (N_2596,N_7,N_473);
and U2597 (N_2597,N_1035,N_198);
nor U2598 (N_2598,N_1279,N_244);
and U2599 (N_2599,N_1438,N_945);
nor U2600 (N_2600,N_353,N_697);
nand U2601 (N_2601,N_1415,N_822);
xnor U2602 (N_2602,N_207,N_1020);
or U2603 (N_2603,N_567,N_316);
or U2604 (N_2604,N_64,N_177);
or U2605 (N_2605,N_439,N_215);
nor U2606 (N_2606,N_58,N_1163);
xor U2607 (N_2607,N_1467,N_62);
xor U2608 (N_2608,N_417,N_132);
nor U2609 (N_2609,N_634,N_553);
or U2610 (N_2610,N_313,N_1241);
nor U2611 (N_2611,N_504,N_1105);
and U2612 (N_2612,N_1206,N_1446);
xor U2613 (N_2613,N_416,N_1372);
and U2614 (N_2614,N_236,N_1118);
xnor U2615 (N_2615,N_748,N_1126);
or U2616 (N_2616,N_1207,N_1093);
or U2617 (N_2617,N_132,N_1359);
nor U2618 (N_2618,N_1241,N_20);
and U2619 (N_2619,N_1293,N_698);
and U2620 (N_2620,N_870,N_1029);
nand U2621 (N_2621,N_358,N_415);
nand U2622 (N_2622,N_376,N_69);
xnor U2623 (N_2623,N_317,N_829);
nand U2624 (N_2624,N_327,N_551);
nor U2625 (N_2625,N_1379,N_360);
nor U2626 (N_2626,N_104,N_609);
nand U2627 (N_2627,N_806,N_285);
or U2628 (N_2628,N_1386,N_1397);
or U2629 (N_2629,N_867,N_875);
nor U2630 (N_2630,N_439,N_235);
or U2631 (N_2631,N_1242,N_1299);
or U2632 (N_2632,N_38,N_689);
nor U2633 (N_2633,N_626,N_1197);
or U2634 (N_2634,N_116,N_462);
nor U2635 (N_2635,N_859,N_706);
nand U2636 (N_2636,N_1425,N_1020);
xnor U2637 (N_2637,N_1409,N_888);
and U2638 (N_2638,N_960,N_1159);
and U2639 (N_2639,N_790,N_575);
or U2640 (N_2640,N_1213,N_97);
nor U2641 (N_2641,N_1469,N_166);
or U2642 (N_2642,N_617,N_57);
and U2643 (N_2643,N_1353,N_427);
nor U2644 (N_2644,N_96,N_1178);
nand U2645 (N_2645,N_247,N_438);
nor U2646 (N_2646,N_790,N_67);
and U2647 (N_2647,N_1429,N_1290);
nand U2648 (N_2648,N_299,N_375);
or U2649 (N_2649,N_437,N_795);
nor U2650 (N_2650,N_1157,N_328);
xor U2651 (N_2651,N_1030,N_622);
nor U2652 (N_2652,N_939,N_734);
nor U2653 (N_2653,N_1124,N_225);
xnor U2654 (N_2654,N_127,N_513);
and U2655 (N_2655,N_637,N_1402);
nand U2656 (N_2656,N_1011,N_152);
or U2657 (N_2657,N_549,N_1219);
xor U2658 (N_2658,N_1480,N_980);
nor U2659 (N_2659,N_503,N_584);
and U2660 (N_2660,N_952,N_384);
or U2661 (N_2661,N_492,N_851);
or U2662 (N_2662,N_1367,N_527);
and U2663 (N_2663,N_857,N_327);
and U2664 (N_2664,N_896,N_1144);
and U2665 (N_2665,N_705,N_422);
nor U2666 (N_2666,N_1289,N_804);
nand U2667 (N_2667,N_891,N_1481);
xnor U2668 (N_2668,N_1027,N_275);
nand U2669 (N_2669,N_1370,N_478);
nor U2670 (N_2670,N_270,N_8);
nor U2671 (N_2671,N_505,N_978);
xnor U2672 (N_2672,N_306,N_834);
nand U2673 (N_2673,N_387,N_625);
nor U2674 (N_2674,N_422,N_796);
xnor U2675 (N_2675,N_1440,N_358);
nand U2676 (N_2676,N_1,N_848);
nor U2677 (N_2677,N_1268,N_748);
and U2678 (N_2678,N_395,N_1231);
nand U2679 (N_2679,N_1344,N_916);
nand U2680 (N_2680,N_700,N_102);
nor U2681 (N_2681,N_234,N_990);
xnor U2682 (N_2682,N_1279,N_1320);
nand U2683 (N_2683,N_844,N_571);
and U2684 (N_2684,N_839,N_843);
and U2685 (N_2685,N_1021,N_64);
xnor U2686 (N_2686,N_373,N_1450);
nor U2687 (N_2687,N_1346,N_588);
nor U2688 (N_2688,N_151,N_1295);
xor U2689 (N_2689,N_497,N_1400);
xnor U2690 (N_2690,N_506,N_256);
nand U2691 (N_2691,N_1031,N_1046);
nand U2692 (N_2692,N_974,N_1222);
or U2693 (N_2693,N_842,N_967);
or U2694 (N_2694,N_394,N_938);
xor U2695 (N_2695,N_1453,N_889);
nor U2696 (N_2696,N_41,N_582);
or U2697 (N_2697,N_1435,N_1034);
xnor U2698 (N_2698,N_1242,N_43);
xnor U2699 (N_2699,N_799,N_339);
xnor U2700 (N_2700,N_1375,N_1319);
and U2701 (N_2701,N_754,N_104);
or U2702 (N_2702,N_472,N_742);
and U2703 (N_2703,N_1009,N_120);
xnor U2704 (N_2704,N_183,N_620);
xnor U2705 (N_2705,N_887,N_581);
and U2706 (N_2706,N_445,N_943);
and U2707 (N_2707,N_1342,N_1462);
and U2708 (N_2708,N_958,N_1068);
and U2709 (N_2709,N_332,N_922);
or U2710 (N_2710,N_103,N_1407);
xnor U2711 (N_2711,N_1321,N_629);
nor U2712 (N_2712,N_1437,N_1470);
xnor U2713 (N_2713,N_589,N_984);
xnor U2714 (N_2714,N_1155,N_532);
or U2715 (N_2715,N_1163,N_1214);
xor U2716 (N_2716,N_436,N_1317);
nor U2717 (N_2717,N_449,N_704);
or U2718 (N_2718,N_251,N_950);
and U2719 (N_2719,N_1343,N_394);
or U2720 (N_2720,N_1280,N_857);
and U2721 (N_2721,N_507,N_1196);
nor U2722 (N_2722,N_253,N_812);
or U2723 (N_2723,N_962,N_1093);
nor U2724 (N_2724,N_1379,N_1334);
or U2725 (N_2725,N_1002,N_720);
xor U2726 (N_2726,N_591,N_299);
nor U2727 (N_2727,N_559,N_753);
or U2728 (N_2728,N_316,N_253);
nor U2729 (N_2729,N_442,N_1190);
nor U2730 (N_2730,N_1129,N_335);
xor U2731 (N_2731,N_1368,N_1213);
or U2732 (N_2732,N_709,N_676);
nor U2733 (N_2733,N_1376,N_979);
and U2734 (N_2734,N_736,N_1209);
nor U2735 (N_2735,N_204,N_817);
nor U2736 (N_2736,N_1303,N_354);
xor U2737 (N_2737,N_639,N_958);
xor U2738 (N_2738,N_452,N_1083);
or U2739 (N_2739,N_256,N_426);
nor U2740 (N_2740,N_1360,N_188);
or U2741 (N_2741,N_400,N_660);
and U2742 (N_2742,N_982,N_673);
nor U2743 (N_2743,N_1299,N_993);
xor U2744 (N_2744,N_32,N_1341);
or U2745 (N_2745,N_1205,N_573);
nor U2746 (N_2746,N_1134,N_262);
nand U2747 (N_2747,N_323,N_1078);
xor U2748 (N_2748,N_387,N_285);
and U2749 (N_2749,N_534,N_1101);
nor U2750 (N_2750,N_921,N_917);
nor U2751 (N_2751,N_802,N_1347);
xor U2752 (N_2752,N_1116,N_269);
or U2753 (N_2753,N_1074,N_1227);
nor U2754 (N_2754,N_1446,N_1468);
xnor U2755 (N_2755,N_1052,N_853);
xor U2756 (N_2756,N_1215,N_1028);
nor U2757 (N_2757,N_1053,N_716);
xor U2758 (N_2758,N_1247,N_1383);
and U2759 (N_2759,N_714,N_54);
or U2760 (N_2760,N_14,N_1027);
nor U2761 (N_2761,N_433,N_1126);
or U2762 (N_2762,N_1126,N_968);
nand U2763 (N_2763,N_944,N_801);
and U2764 (N_2764,N_449,N_627);
and U2765 (N_2765,N_536,N_1371);
xor U2766 (N_2766,N_998,N_68);
or U2767 (N_2767,N_28,N_1350);
and U2768 (N_2768,N_1006,N_721);
and U2769 (N_2769,N_1415,N_904);
xor U2770 (N_2770,N_1187,N_167);
or U2771 (N_2771,N_820,N_999);
nand U2772 (N_2772,N_518,N_679);
xor U2773 (N_2773,N_121,N_409);
nand U2774 (N_2774,N_38,N_1128);
nand U2775 (N_2775,N_668,N_981);
nand U2776 (N_2776,N_1182,N_434);
and U2777 (N_2777,N_1088,N_468);
nand U2778 (N_2778,N_211,N_1143);
xor U2779 (N_2779,N_1332,N_1238);
and U2780 (N_2780,N_1385,N_1081);
nand U2781 (N_2781,N_145,N_1139);
nor U2782 (N_2782,N_1185,N_1032);
nand U2783 (N_2783,N_307,N_1047);
nand U2784 (N_2784,N_338,N_674);
nand U2785 (N_2785,N_853,N_867);
and U2786 (N_2786,N_1362,N_973);
nor U2787 (N_2787,N_517,N_1363);
and U2788 (N_2788,N_520,N_199);
or U2789 (N_2789,N_1444,N_582);
and U2790 (N_2790,N_91,N_149);
and U2791 (N_2791,N_648,N_490);
or U2792 (N_2792,N_1392,N_989);
nor U2793 (N_2793,N_1332,N_611);
nor U2794 (N_2794,N_359,N_1195);
nor U2795 (N_2795,N_1308,N_339);
or U2796 (N_2796,N_657,N_525);
or U2797 (N_2797,N_373,N_816);
nor U2798 (N_2798,N_680,N_564);
and U2799 (N_2799,N_854,N_1123);
nand U2800 (N_2800,N_443,N_1351);
and U2801 (N_2801,N_940,N_827);
xnor U2802 (N_2802,N_1338,N_514);
or U2803 (N_2803,N_1470,N_948);
or U2804 (N_2804,N_332,N_1106);
and U2805 (N_2805,N_944,N_601);
nand U2806 (N_2806,N_231,N_143);
xor U2807 (N_2807,N_1159,N_292);
and U2808 (N_2808,N_889,N_23);
nor U2809 (N_2809,N_439,N_643);
nor U2810 (N_2810,N_847,N_1481);
xor U2811 (N_2811,N_1372,N_324);
nand U2812 (N_2812,N_169,N_1353);
and U2813 (N_2813,N_1155,N_823);
xnor U2814 (N_2814,N_788,N_1377);
nor U2815 (N_2815,N_87,N_469);
nor U2816 (N_2816,N_250,N_934);
or U2817 (N_2817,N_651,N_154);
nor U2818 (N_2818,N_1204,N_91);
nor U2819 (N_2819,N_192,N_1397);
or U2820 (N_2820,N_379,N_508);
xnor U2821 (N_2821,N_582,N_378);
and U2822 (N_2822,N_1202,N_368);
nor U2823 (N_2823,N_614,N_896);
nand U2824 (N_2824,N_497,N_518);
nor U2825 (N_2825,N_1001,N_17);
xor U2826 (N_2826,N_951,N_1469);
nor U2827 (N_2827,N_1170,N_1489);
nand U2828 (N_2828,N_179,N_538);
nand U2829 (N_2829,N_500,N_305);
or U2830 (N_2830,N_494,N_303);
nor U2831 (N_2831,N_976,N_884);
nor U2832 (N_2832,N_965,N_756);
nand U2833 (N_2833,N_33,N_827);
or U2834 (N_2834,N_1313,N_397);
nand U2835 (N_2835,N_647,N_825);
nand U2836 (N_2836,N_1323,N_563);
and U2837 (N_2837,N_1339,N_355);
nand U2838 (N_2838,N_95,N_310);
or U2839 (N_2839,N_1287,N_7);
nand U2840 (N_2840,N_1210,N_775);
nand U2841 (N_2841,N_225,N_111);
and U2842 (N_2842,N_1043,N_1173);
or U2843 (N_2843,N_1480,N_992);
and U2844 (N_2844,N_1441,N_943);
nand U2845 (N_2845,N_186,N_774);
nor U2846 (N_2846,N_640,N_1304);
nand U2847 (N_2847,N_431,N_109);
and U2848 (N_2848,N_290,N_16);
or U2849 (N_2849,N_829,N_387);
xor U2850 (N_2850,N_1033,N_846);
and U2851 (N_2851,N_1114,N_599);
xnor U2852 (N_2852,N_544,N_1347);
nor U2853 (N_2853,N_383,N_1276);
or U2854 (N_2854,N_376,N_928);
and U2855 (N_2855,N_711,N_356);
nor U2856 (N_2856,N_375,N_568);
and U2857 (N_2857,N_671,N_975);
xor U2858 (N_2858,N_1441,N_676);
or U2859 (N_2859,N_120,N_40);
xnor U2860 (N_2860,N_389,N_886);
nor U2861 (N_2861,N_1038,N_968);
nor U2862 (N_2862,N_789,N_1225);
nor U2863 (N_2863,N_109,N_538);
or U2864 (N_2864,N_1046,N_205);
nor U2865 (N_2865,N_1092,N_673);
or U2866 (N_2866,N_905,N_27);
nand U2867 (N_2867,N_37,N_913);
and U2868 (N_2868,N_843,N_1290);
xnor U2869 (N_2869,N_222,N_148);
or U2870 (N_2870,N_1367,N_1498);
xnor U2871 (N_2871,N_883,N_327);
and U2872 (N_2872,N_713,N_933);
nor U2873 (N_2873,N_581,N_289);
nand U2874 (N_2874,N_611,N_1429);
xnor U2875 (N_2875,N_882,N_1231);
nand U2876 (N_2876,N_80,N_1250);
and U2877 (N_2877,N_594,N_833);
nand U2878 (N_2878,N_996,N_1353);
nand U2879 (N_2879,N_1300,N_607);
nand U2880 (N_2880,N_1495,N_628);
nand U2881 (N_2881,N_922,N_1117);
nor U2882 (N_2882,N_1057,N_643);
xnor U2883 (N_2883,N_758,N_423);
nor U2884 (N_2884,N_1220,N_1031);
xnor U2885 (N_2885,N_847,N_1285);
or U2886 (N_2886,N_852,N_1110);
xnor U2887 (N_2887,N_822,N_468);
or U2888 (N_2888,N_512,N_1383);
xor U2889 (N_2889,N_101,N_1431);
xnor U2890 (N_2890,N_907,N_1269);
nor U2891 (N_2891,N_1102,N_95);
nand U2892 (N_2892,N_279,N_373);
xnor U2893 (N_2893,N_878,N_1443);
and U2894 (N_2894,N_689,N_331);
nor U2895 (N_2895,N_335,N_953);
and U2896 (N_2896,N_501,N_896);
nand U2897 (N_2897,N_1100,N_992);
xnor U2898 (N_2898,N_1177,N_672);
nor U2899 (N_2899,N_1081,N_317);
or U2900 (N_2900,N_350,N_335);
or U2901 (N_2901,N_135,N_60);
and U2902 (N_2902,N_1252,N_524);
or U2903 (N_2903,N_1015,N_1014);
nand U2904 (N_2904,N_1301,N_1227);
and U2905 (N_2905,N_933,N_835);
nor U2906 (N_2906,N_125,N_1490);
or U2907 (N_2907,N_631,N_915);
xnor U2908 (N_2908,N_868,N_1272);
and U2909 (N_2909,N_1345,N_903);
or U2910 (N_2910,N_1058,N_953);
nor U2911 (N_2911,N_248,N_985);
nor U2912 (N_2912,N_572,N_594);
xnor U2913 (N_2913,N_1354,N_570);
nand U2914 (N_2914,N_141,N_208);
nand U2915 (N_2915,N_499,N_1361);
or U2916 (N_2916,N_537,N_542);
xnor U2917 (N_2917,N_1002,N_319);
or U2918 (N_2918,N_1003,N_528);
xor U2919 (N_2919,N_1192,N_1268);
xnor U2920 (N_2920,N_546,N_456);
xnor U2921 (N_2921,N_652,N_879);
nor U2922 (N_2922,N_440,N_41);
xor U2923 (N_2923,N_901,N_424);
nand U2924 (N_2924,N_276,N_832);
or U2925 (N_2925,N_251,N_149);
nand U2926 (N_2926,N_155,N_534);
xnor U2927 (N_2927,N_789,N_918);
or U2928 (N_2928,N_1131,N_859);
or U2929 (N_2929,N_410,N_814);
nand U2930 (N_2930,N_1181,N_292);
or U2931 (N_2931,N_14,N_172);
xnor U2932 (N_2932,N_344,N_49);
or U2933 (N_2933,N_978,N_336);
nand U2934 (N_2934,N_1342,N_161);
and U2935 (N_2935,N_702,N_377);
nor U2936 (N_2936,N_251,N_1077);
xor U2937 (N_2937,N_384,N_714);
xor U2938 (N_2938,N_480,N_965);
nor U2939 (N_2939,N_772,N_1212);
nor U2940 (N_2940,N_899,N_1231);
nand U2941 (N_2941,N_1479,N_1062);
and U2942 (N_2942,N_1395,N_1440);
nand U2943 (N_2943,N_459,N_174);
or U2944 (N_2944,N_819,N_1143);
xor U2945 (N_2945,N_338,N_1309);
nand U2946 (N_2946,N_1235,N_1243);
xor U2947 (N_2947,N_1268,N_1117);
nor U2948 (N_2948,N_503,N_590);
or U2949 (N_2949,N_749,N_952);
nor U2950 (N_2950,N_1360,N_1147);
and U2951 (N_2951,N_302,N_801);
nor U2952 (N_2952,N_334,N_297);
xor U2953 (N_2953,N_1268,N_1175);
nand U2954 (N_2954,N_1418,N_402);
nor U2955 (N_2955,N_1473,N_850);
xor U2956 (N_2956,N_394,N_468);
xnor U2957 (N_2957,N_801,N_781);
xnor U2958 (N_2958,N_489,N_889);
xor U2959 (N_2959,N_1195,N_1091);
xor U2960 (N_2960,N_813,N_793);
xor U2961 (N_2961,N_59,N_62);
xnor U2962 (N_2962,N_602,N_634);
xnor U2963 (N_2963,N_566,N_1335);
nand U2964 (N_2964,N_1460,N_338);
nor U2965 (N_2965,N_461,N_460);
or U2966 (N_2966,N_997,N_54);
nand U2967 (N_2967,N_9,N_695);
or U2968 (N_2968,N_889,N_1324);
and U2969 (N_2969,N_1446,N_1412);
nor U2970 (N_2970,N_969,N_852);
and U2971 (N_2971,N_589,N_1357);
nand U2972 (N_2972,N_166,N_1038);
xor U2973 (N_2973,N_1078,N_219);
nand U2974 (N_2974,N_634,N_723);
xnor U2975 (N_2975,N_1117,N_355);
nand U2976 (N_2976,N_576,N_1325);
or U2977 (N_2977,N_645,N_511);
xor U2978 (N_2978,N_605,N_216);
and U2979 (N_2979,N_587,N_37);
and U2980 (N_2980,N_1047,N_309);
xor U2981 (N_2981,N_697,N_1312);
nor U2982 (N_2982,N_713,N_641);
or U2983 (N_2983,N_1012,N_157);
and U2984 (N_2984,N_24,N_874);
nor U2985 (N_2985,N_1031,N_1394);
nand U2986 (N_2986,N_35,N_351);
or U2987 (N_2987,N_1182,N_144);
or U2988 (N_2988,N_12,N_1289);
nand U2989 (N_2989,N_1007,N_1205);
and U2990 (N_2990,N_585,N_503);
xnor U2991 (N_2991,N_891,N_713);
nor U2992 (N_2992,N_372,N_659);
nor U2993 (N_2993,N_501,N_1453);
nor U2994 (N_2994,N_801,N_1221);
or U2995 (N_2995,N_154,N_155);
and U2996 (N_2996,N_1195,N_611);
and U2997 (N_2997,N_1113,N_1293);
or U2998 (N_2998,N_1352,N_342);
or U2999 (N_2999,N_192,N_865);
or U3000 (N_3000,N_2646,N_2050);
or U3001 (N_3001,N_2099,N_2910);
xor U3002 (N_3002,N_1686,N_2361);
nor U3003 (N_3003,N_1550,N_2253);
or U3004 (N_3004,N_1590,N_2865);
or U3005 (N_3005,N_1616,N_2024);
and U3006 (N_3006,N_1776,N_1558);
and U3007 (N_3007,N_1755,N_1775);
nor U3008 (N_3008,N_2570,N_1933);
xor U3009 (N_3009,N_2180,N_2236);
nor U3010 (N_3010,N_2125,N_1709);
and U3011 (N_3011,N_1780,N_2883);
or U3012 (N_3012,N_1834,N_2887);
xnor U3013 (N_3013,N_1760,N_1994);
and U3014 (N_3014,N_2440,N_2963);
and U3015 (N_3015,N_2154,N_2296);
and U3016 (N_3016,N_2218,N_2721);
nand U3017 (N_3017,N_2697,N_2826);
nor U3018 (N_3018,N_2785,N_2936);
nand U3019 (N_3019,N_2012,N_1670);
or U3020 (N_3020,N_2397,N_2542);
nand U3021 (N_3021,N_2411,N_1870);
and U3022 (N_3022,N_2060,N_2039);
nor U3023 (N_3023,N_2607,N_1844);
or U3024 (N_3024,N_1715,N_1826);
nand U3025 (N_3025,N_2392,N_2942);
nor U3026 (N_3026,N_2699,N_1869);
nand U3027 (N_3027,N_1599,N_2226);
nand U3028 (N_3028,N_2745,N_2834);
xor U3029 (N_3029,N_1552,N_2352);
nand U3030 (N_3030,N_2275,N_1716);
and U3031 (N_3031,N_1608,N_2045);
nand U3032 (N_3032,N_1671,N_1965);
nor U3033 (N_3033,N_2813,N_2464);
xnor U3034 (N_3034,N_2533,N_1692);
nand U3035 (N_3035,N_2284,N_1816);
xor U3036 (N_3036,N_1668,N_1974);
nor U3037 (N_3037,N_2162,N_2308);
xnor U3038 (N_3038,N_2021,N_1510);
nor U3039 (N_3039,N_2119,N_2508);
or U3040 (N_3040,N_2825,N_2652);
and U3041 (N_3041,N_2729,N_1751);
and U3042 (N_3042,N_1701,N_1582);
nor U3043 (N_3043,N_1549,N_2685);
nand U3044 (N_3044,N_2769,N_2002);
and U3045 (N_3045,N_1707,N_2069);
and U3046 (N_3046,N_2600,N_2334);
xnor U3047 (N_3047,N_1644,N_1996);
xor U3048 (N_3048,N_2493,N_2297);
or U3049 (N_3049,N_2810,N_2344);
xnor U3050 (N_3050,N_1587,N_2617);
xnor U3051 (N_3051,N_2313,N_2495);
nor U3052 (N_3052,N_2071,N_2609);
or U3053 (N_3053,N_2841,N_1792);
or U3054 (N_3054,N_2677,N_2790);
nor U3055 (N_3055,N_2486,N_2023);
nand U3056 (N_3056,N_1922,N_2482);
or U3057 (N_3057,N_1883,N_2453);
and U3058 (N_3058,N_2294,N_2968);
and U3059 (N_3059,N_2139,N_2648);
and U3060 (N_3060,N_1832,N_2580);
xnor U3061 (N_3061,N_1607,N_2624);
or U3062 (N_3062,N_1837,N_2514);
or U3063 (N_3063,N_2110,N_2232);
nand U3064 (N_3064,N_2639,N_1509);
or U3065 (N_3065,N_2003,N_2475);
and U3066 (N_3066,N_1738,N_2895);
nand U3067 (N_3067,N_1949,N_2808);
or U3068 (N_3068,N_2571,N_1626);
nand U3069 (N_3069,N_2080,N_2563);
nand U3070 (N_3070,N_2282,N_2207);
and U3071 (N_3071,N_1808,N_1989);
nand U3072 (N_3072,N_2916,N_1725);
or U3073 (N_3073,N_2890,N_2703);
nor U3074 (N_3074,N_2714,N_2529);
nor U3075 (N_3075,N_2142,N_2485);
nor U3076 (N_3076,N_2368,N_2788);
nor U3077 (N_3077,N_2324,N_2972);
or U3078 (N_3078,N_2527,N_1782);
nor U3079 (N_3079,N_2688,N_2447);
xnor U3080 (N_3080,N_1501,N_2731);
xnor U3081 (N_3081,N_2399,N_2102);
nand U3082 (N_3082,N_2047,N_1546);
or U3083 (N_3083,N_2927,N_1636);
xor U3084 (N_3084,N_1873,N_2779);
nand U3085 (N_3085,N_1554,N_1547);
and U3086 (N_3086,N_2784,N_2032);
xnor U3087 (N_3087,N_1802,N_2698);
or U3088 (N_3088,N_2242,N_2847);
nand U3089 (N_3089,N_2468,N_1769);
nor U3090 (N_3090,N_1931,N_2262);
and U3091 (N_3091,N_1524,N_1929);
or U3092 (N_3092,N_1932,N_2494);
and U3093 (N_3093,N_2857,N_2492);
xor U3094 (N_3094,N_2436,N_1847);
or U3095 (N_3095,N_2764,N_2064);
xnor U3096 (N_3096,N_1589,N_2220);
nand U3097 (N_3097,N_2097,N_2510);
xor U3098 (N_3098,N_1807,N_2231);
xnor U3099 (N_3099,N_2554,N_2862);
nand U3100 (N_3100,N_2588,N_1528);
nand U3101 (N_3101,N_1655,N_1814);
or U3102 (N_3102,N_2552,N_1525);
and U3103 (N_3103,N_2035,N_2766);
xor U3104 (N_3104,N_2637,N_2960);
nor U3105 (N_3105,N_1817,N_2430);
nand U3106 (N_3106,N_2298,N_1777);
xnor U3107 (N_3107,N_1878,N_2051);
nand U3108 (N_3108,N_2418,N_2442);
nand U3109 (N_3109,N_2901,N_1720);
nand U3110 (N_3110,N_1864,N_2500);
xor U3111 (N_3111,N_2013,N_2780);
nor U3112 (N_3112,N_1646,N_2011);
nand U3113 (N_3113,N_2028,N_1905);
nor U3114 (N_3114,N_1940,N_1544);
or U3115 (N_3115,N_1950,N_2992);
xor U3116 (N_3116,N_1819,N_2844);
nor U3117 (N_3117,N_2522,N_2363);
and U3118 (N_3118,N_1879,N_2777);
nor U3119 (N_3119,N_2305,N_2196);
nor U3120 (N_3120,N_1737,N_2595);
and U3121 (N_3121,N_2015,N_2541);
nand U3122 (N_3122,N_1963,N_1514);
nor U3123 (N_3123,N_1747,N_1604);
nor U3124 (N_3124,N_2722,N_1714);
and U3125 (N_3125,N_1856,N_2423);
and U3126 (N_3126,N_1627,N_1866);
or U3127 (N_3127,N_1954,N_1827);
or U3128 (N_3128,N_2439,N_2585);
xnor U3129 (N_3129,N_2340,N_1538);
nand U3130 (N_3130,N_2031,N_1799);
xnor U3131 (N_3131,N_2962,N_2668);
or U3132 (N_3132,N_1673,N_1763);
or U3133 (N_3133,N_1831,N_2837);
and U3134 (N_3134,N_2311,N_2036);
or U3135 (N_3135,N_2062,N_2303);
or U3136 (N_3136,N_2172,N_1825);
nand U3137 (N_3137,N_1730,N_1642);
and U3138 (N_3138,N_2353,N_2728);
nor U3139 (N_3139,N_2866,N_2077);
or U3140 (N_3140,N_2871,N_1535);
or U3141 (N_3141,N_1679,N_2185);
nor U3142 (N_3142,N_2767,N_2512);
nand U3143 (N_3143,N_2855,N_2118);
nand U3144 (N_3144,N_2754,N_2638);
or U3145 (N_3145,N_1838,N_2647);
nor U3146 (N_3146,N_2557,N_1973);
xor U3147 (N_3147,N_2758,N_2641);
nand U3148 (N_3148,N_2854,N_1860);
or U3149 (N_3149,N_2513,N_1995);
and U3150 (N_3150,N_1648,N_1762);
and U3151 (N_3151,N_2177,N_2944);
nor U3152 (N_3152,N_2759,N_2695);
nor U3153 (N_3153,N_1906,N_2234);
nand U3154 (N_3154,N_1829,N_2285);
nand U3155 (N_3155,N_2355,N_2058);
nor U3156 (N_3156,N_2987,N_2038);
nor U3157 (N_3157,N_1784,N_1536);
or U3158 (N_3158,N_1678,N_2259);
nor U3159 (N_3159,N_1993,N_1764);
or U3160 (N_3160,N_1888,N_2613);
nand U3161 (N_3161,N_1533,N_2875);
xnor U3162 (N_3162,N_2587,N_2105);
xor U3163 (N_3163,N_2822,N_2371);
nand U3164 (N_3164,N_2248,N_2249);
nor U3165 (N_3165,N_2765,N_1664);
and U3166 (N_3166,N_2933,N_2615);
and U3167 (N_3167,N_2267,N_1676);
or U3168 (N_3168,N_1958,N_2351);
and U3169 (N_3169,N_1821,N_2596);
and U3170 (N_3170,N_2863,N_2655);
xor U3171 (N_3171,N_1895,N_2190);
nor U3172 (N_3172,N_2319,N_2280);
or U3173 (N_3173,N_1809,N_2385);
xnor U3174 (N_3174,N_2906,N_1836);
nand U3175 (N_3175,N_1884,N_2073);
nor U3176 (N_3176,N_2739,N_2343);
nand U3177 (N_3177,N_2331,N_2330);
and U3178 (N_3178,N_1592,N_2461);
or U3179 (N_3179,N_2264,N_2473);
xor U3180 (N_3180,N_1946,N_2061);
and U3181 (N_3181,N_1850,N_1962);
or U3182 (N_3182,N_2454,N_2400);
xnor U3183 (N_3183,N_2969,N_1767);
or U3184 (N_3184,N_2551,N_2044);
or U3185 (N_3185,N_2422,N_2431);
or U3186 (N_3186,N_2066,N_2445);
nand U3187 (N_3187,N_2830,N_2052);
and U3188 (N_3188,N_1822,N_1881);
or U3189 (N_3189,N_1904,N_1619);
nor U3190 (N_3190,N_2457,N_2559);
and U3191 (N_3191,N_2009,N_2792);
xnor U3192 (N_3192,N_2221,N_1859);
xnor U3193 (N_3193,N_2832,N_2082);
nor U3194 (N_3194,N_2281,N_1991);
xnor U3195 (N_3195,N_2326,N_2618);
xnor U3196 (N_3196,N_2836,N_2268);
nor U3197 (N_3197,N_2575,N_2138);
and U3198 (N_3198,N_1794,N_1861);
nand U3199 (N_3199,N_2113,N_2474);
nor U3200 (N_3200,N_2446,N_1611);
nand U3201 (N_3201,N_2374,N_1740);
nand U3202 (N_3202,N_2931,N_2437);
nor U3203 (N_3203,N_1721,N_1718);
xnor U3204 (N_3204,N_1894,N_2572);
nor U3205 (N_3205,N_2902,N_2567);
nand U3206 (N_3206,N_1727,N_2643);
nand U3207 (N_3207,N_1943,N_1935);
and U3208 (N_3208,N_1773,N_2880);
or U3209 (N_3209,N_2383,N_2460);
nor U3210 (N_3210,N_2318,N_2347);
nand U3211 (N_3211,N_1577,N_2074);
nor U3212 (N_3212,N_1635,N_1517);
xnor U3213 (N_3213,N_1539,N_1951);
nor U3214 (N_3214,N_1801,N_2915);
nor U3215 (N_3215,N_2574,N_2977);
and U3216 (N_3216,N_1778,N_2908);
nor U3217 (N_3217,N_2250,N_2255);
xor U3218 (N_3218,N_1818,N_2273);
nor U3219 (N_3219,N_2743,N_1529);
xor U3220 (N_3220,N_2922,N_2310);
and U3221 (N_3221,N_1613,N_1977);
nor U3222 (N_3222,N_2578,N_2982);
xnor U3223 (N_3223,N_2725,N_2433);
nand U3224 (N_3224,N_1862,N_1803);
xor U3225 (N_3225,N_2970,N_2175);
nor U3226 (N_3226,N_2621,N_2342);
nand U3227 (N_3227,N_1992,N_1909);
or U3228 (N_3228,N_2389,N_2372);
xnor U3229 (N_3229,N_2043,N_2091);
and U3230 (N_3230,N_2599,N_1796);
nand U3231 (N_3231,N_2472,N_1659);
nor U3232 (N_3232,N_2881,N_2965);
nor U3233 (N_3233,N_1982,N_1921);
or U3234 (N_3234,N_1891,N_1979);
xnor U3235 (N_3235,N_2322,N_2543);
or U3236 (N_3236,N_2116,N_1581);
nand U3237 (N_3237,N_1724,N_2734);
nand U3238 (N_3238,N_2919,N_2499);
nand U3239 (N_3239,N_2809,N_2868);
and U3240 (N_3240,N_1824,N_2186);
nor U3241 (N_3241,N_2197,N_2669);
and U3242 (N_3242,N_2478,N_2896);
nand U3243 (N_3243,N_1938,N_2067);
nand U3244 (N_3244,N_1926,N_1649);
nor U3245 (N_3245,N_2840,N_2148);
or U3246 (N_3246,N_2266,N_2993);
nand U3247 (N_3247,N_2791,N_2664);
or U3248 (N_3248,N_2793,N_1503);
or U3249 (N_3249,N_2424,N_1662);
xnor U3250 (N_3250,N_1735,N_1658);
or U3251 (N_3251,N_2651,N_2042);
and U3252 (N_3252,N_1543,N_2634);
and U3253 (N_3253,N_1537,N_2054);
nor U3254 (N_3254,N_2321,N_1561);
nand U3255 (N_3255,N_2667,N_2631);
and U3256 (N_3256,N_2124,N_2851);
or U3257 (N_3257,N_1706,N_1936);
xnor U3258 (N_3258,N_2362,N_2103);
or U3259 (N_3259,N_2348,N_2828);
or U3260 (N_3260,N_2366,N_2341);
nor U3261 (N_3261,N_1585,N_1609);
or U3262 (N_3262,N_2496,N_1615);
nand U3263 (N_3263,N_2787,N_2597);
and U3264 (N_3264,N_2553,N_2209);
and U3265 (N_3265,N_1956,N_2727);
and U3266 (N_3266,N_2975,N_1512);
and U3267 (N_3267,N_2246,N_1752);
nor U3268 (N_3268,N_1896,N_2923);
nand U3269 (N_3269,N_1942,N_2309);
or U3270 (N_3270,N_2605,N_2573);
nor U3271 (N_3271,N_2451,N_2945);
and U3272 (N_3272,N_1748,N_1882);
nor U3273 (N_3273,N_1653,N_2241);
xnor U3274 (N_3274,N_1971,N_1563);
or U3275 (N_3275,N_2462,N_2428);
or U3276 (N_3276,N_2131,N_2084);
and U3277 (N_3277,N_1813,N_1877);
and U3278 (N_3278,N_1759,N_2092);
nor U3279 (N_3279,N_2692,N_2215);
and U3280 (N_3280,N_1540,N_1574);
or U3281 (N_3281,N_2320,N_1672);
xor U3282 (N_3282,N_1560,N_2415);
xor U3283 (N_3283,N_2818,N_1843);
xnor U3284 (N_3284,N_1772,N_2789);
or U3285 (N_3285,N_2506,N_2258);
and U3286 (N_3286,N_2978,N_2771);
xor U3287 (N_3287,N_2879,N_2252);
nand U3288 (N_3288,N_2187,N_1907);
nor U3289 (N_3289,N_2225,N_1781);
or U3290 (N_3290,N_1732,N_1976);
and U3291 (N_3291,N_1887,N_2477);
or U3292 (N_3292,N_1736,N_1923);
or U3293 (N_3293,N_2864,N_2191);
and U3294 (N_3294,N_2738,N_2452);
xor U3295 (N_3295,N_2804,N_1559);
or U3296 (N_3296,N_2659,N_2206);
nor U3297 (N_3297,N_1790,N_2921);
xnor U3298 (N_3298,N_1912,N_1702);
and U3299 (N_3299,N_2598,N_2239);
xor U3300 (N_3300,N_1614,N_2536);
nand U3301 (N_3301,N_2996,N_1705);
and U3302 (N_3302,N_2360,N_2194);
or U3303 (N_3303,N_2085,N_2546);
nand U3304 (N_3304,N_2746,N_1591);
and U3305 (N_3305,N_2858,N_2345);
nand U3306 (N_3306,N_2426,N_2523);
and U3307 (N_3307,N_1680,N_2670);
or U3308 (N_3308,N_2888,N_2886);
or U3309 (N_3309,N_1774,N_2229);
and U3310 (N_3310,N_2420,N_2682);
xnor U3311 (N_3311,N_2316,N_2405);
and U3312 (N_3312,N_2748,N_2020);
and U3313 (N_3313,N_2136,N_2704);
or U3314 (N_3314,N_1745,N_2724);
or U3315 (N_3315,N_2271,N_1798);
nor U3316 (N_3316,N_1791,N_2635);
and U3317 (N_3317,N_2408,N_2716);
and U3318 (N_3318,N_2932,N_2409);
or U3319 (N_3319,N_1975,N_2870);
or U3320 (N_3320,N_1545,N_2539);
xor U3321 (N_3321,N_2315,N_2336);
or U3322 (N_3322,N_2713,N_2601);
and U3323 (N_3323,N_2957,N_2000);
and U3324 (N_3324,N_2129,N_2776);
nand U3325 (N_3325,N_2693,N_2778);
xor U3326 (N_3326,N_2441,N_2630);
and U3327 (N_3327,N_2954,N_2247);
or U3328 (N_3328,N_2096,N_1930);
nor U3329 (N_3329,N_2534,N_2629);
or U3330 (N_3330,N_2853,N_1955);
nor U3331 (N_3331,N_1917,N_2897);
xor U3332 (N_3332,N_2498,N_2737);
nor U3333 (N_3333,N_2158,N_2072);
nand U3334 (N_3334,N_2885,N_1959);
xor U3335 (N_3335,N_1779,N_2939);
xor U3336 (N_3336,N_1569,N_1594);
or U3337 (N_3337,N_1961,N_2106);
and U3338 (N_3338,N_2007,N_2350);
and U3339 (N_3339,N_1666,N_2237);
and U3340 (N_3340,N_2757,N_1576);
and U3341 (N_3341,N_2645,N_2762);
and U3342 (N_3342,N_1557,N_2481);
xnor U3343 (N_3343,N_2217,N_2414);
or U3344 (N_3344,N_2093,N_1750);
nor U3345 (N_3345,N_2604,N_1507);
nor U3346 (N_3346,N_2427,N_2589);
or U3347 (N_3347,N_2839,N_1984);
or U3348 (N_3348,N_1967,N_1661);
xnor U3349 (N_3349,N_1997,N_2544);
nor U3350 (N_3350,N_1712,N_2056);
and U3351 (N_3351,N_1722,N_2590);
nor U3352 (N_3352,N_2376,N_2277);
and U3353 (N_3353,N_2676,N_1522);
nand U3354 (N_3354,N_2100,N_2112);
xor U3355 (N_3355,N_1812,N_2562);
and U3356 (N_3356,N_2549,N_2917);
nand U3357 (N_3357,N_2182,N_2201);
and U3358 (N_3358,N_2204,N_1553);
nand U3359 (N_3359,N_1830,N_2377);
nand U3360 (N_3360,N_1645,N_1597);
nand U3361 (N_3361,N_2794,N_1562);
nand U3362 (N_3362,N_2999,N_1669);
nand U3363 (N_3363,N_2973,N_2168);
nor U3364 (N_3364,N_2504,N_2517);
nand U3365 (N_3365,N_2869,N_2798);
nor U3366 (N_3366,N_2658,N_2959);
nand U3367 (N_3367,N_1939,N_2990);
nor U3368 (N_3368,N_2114,N_1690);
nand U3369 (N_3369,N_2022,N_1863);
and U3370 (N_3370,N_2260,N_2898);
nand U3371 (N_3371,N_2849,N_1889);
nor U3372 (N_3372,N_2299,N_1811);
xor U3373 (N_3373,N_2251,N_2988);
nor U3374 (N_3374,N_1806,N_2735);
or U3375 (N_3375,N_2934,N_2720);
and U3376 (N_3376,N_2878,N_1743);
nand U3377 (N_3377,N_2270,N_2519);
or U3378 (N_3378,N_2511,N_2329);
and U3379 (N_3379,N_2620,N_1835);
nor U3380 (N_3380,N_2711,N_2833);
or U3381 (N_3381,N_1665,N_1704);
nor U3382 (N_3382,N_2566,N_2911);
nand U3383 (N_3383,N_1875,N_2966);
xnor U3384 (N_3384,N_2068,N_2742);
nand U3385 (N_3385,N_2665,N_2821);
xnor U3386 (N_3386,N_2198,N_2359);
and U3387 (N_3387,N_1710,N_1765);
xnor U3388 (N_3388,N_2608,N_2163);
nor U3389 (N_3389,N_2402,N_2169);
nor U3390 (N_3390,N_2663,N_2123);
xor U3391 (N_3391,N_2986,N_1853);
nand U3392 (N_3392,N_1739,N_2594);
and U3393 (N_3393,N_2079,N_2816);
nor U3394 (N_3394,N_1601,N_2393);
nor U3395 (N_3395,N_2490,N_2732);
and U3396 (N_3396,N_2419,N_2971);
or U3397 (N_3397,N_1744,N_2983);
xor U3398 (N_3398,N_1903,N_2041);
nor U3399 (N_3399,N_2435,N_1911);
nand U3400 (N_3400,N_1952,N_2707);
xnor U3401 (N_3401,N_2955,N_2967);
or U3402 (N_3402,N_2679,N_2365);
or U3403 (N_3403,N_2744,N_2122);
or U3404 (N_3404,N_2081,N_2223);
nand U3405 (N_3405,N_2606,N_2354);
or U3406 (N_3406,N_2033,N_2448);
nor U3407 (N_3407,N_2337,N_2900);
and U3408 (N_3408,N_2558,N_2874);
nor U3409 (N_3409,N_2238,N_1849);
xor U3410 (N_3410,N_2287,N_2132);
xnor U3411 (N_3411,N_2314,N_2749);
or U3412 (N_3412,N_1643,N_2382);
and U3413 (N_3413,N_2302,N_2412);
nand U3414 (N_3414,N_2117,N_2384);
and U3415 (N_3415,N_2660,N_2583);
and U3416 (N_3416,N_2650,N_2128);
nand U3417 (N_3417,N_1788,N_2130);
or U3418 (N_3418,N_1603,N_2565);
nand U3419 (N_3419,N_2991,N_1969);
xnor U3420 (N_3420,N_2947,N_1600);
or U3421 (N_3421,N_2135,N_2741);
xor U3422 (N_3422,N_2867,N_2214);
nor U3423 (N_3423,N_1728,N_2421);
and U3424 (N_3424,N_2661,N_2057);
nor U3425 (N_3425,N_2843,N_1519);
xor U3426 (N_3426,N_2257,N_1840);
nand U3427 (N_3427,N_1502,N_1937);
nand U3428 (N_3428,N_1913,N_2904);
or U3429 (N_3429,N_2432,N_2796);
nor U3430 (N_3430,N_2569,N_1868);
and U3431 (N_3431,N_2407,N_2811);
nor U3432 (N_3432,N_2304,N_2859);
nand U3433 (N_3433,N_2127,N_2367);
nor U3434 (N_3434,N_2882,N_2642);
and U3435 (N_3435,N_2610,N_1757);
xnor U3436 (N_3436,N_1511,N_2357);
nor U3437 (N_3437,N_1674,N_2622);
and U3438 (N_3438,N_2687,N_2375);
nor U3439 (N_3439,N_2040,N_2381);
nand U3440 (N_3440,N_1518,N_1846);
or U3441 (N_3441,N_1695,N_2120);
and U3442 (N_3442,N_2459,N_2480);
xnor U3443 (N_3443,N_2937,N_2403);
nor U3444 (N_3444,N_2396,N_2157);
nand U3445 (N_3445,N_1981,N_2404);
xnor U3446 (N_3446,N_2913,N_2998);
nor U3447 (N_3447,N_2438,N_2306);
nor U3448 (N_3448,N_2391,N_1857);
or U3449 (N_3449,N_1711,N_2487);
nand U3450 (N_3450,N_1625,N_2518);
or U3451 (N_3451,N_1852,N_1948);
nand U3452 (N_3452,N_2774,N_2943);
and U3453 (N_3453,N_2216,N_1928);
nand U3454 (N_3454,N_1500,N_2626);
nand U3455 (N_3455,N_1606,N_1681);
xor U3456 (N_3456,N_2899,N_2520);
xor U3457 (N_3457,N_1786,N_1854);
nor U3458 (N_3458,N_2455,N_2877);
or U3459 (N_3459,N_2672,N_1630);
xor U3460 (N_3460,N_2395,N_1631);
nor U3461 (N_3461,N_2004,N_2592);
xnor U3462 (N_3462,N_2290,N_2233);
or U3463 (N_3463,N_2133,N_2701);
nor U3464 (N_3464,N_2628,N_2410);
or U3465 (N_3465,N_1628,N_2696);
nand U3466 (N_3466,N_1970,N_2170);
or U3467 (N_3467,N_1598,N_1842);
or U3468 (N_3468,N_2561,N_1684);
nand U3469 (N_3469,N_1770,N_2540);
xnor U3470 (N_3470,N_1697,N_2550);
or U3471 (N_3471,N_2509,N_2263);
and U3472 (N_3472,N_2770,N_2662);
nor U3473 (N_3473,N_1687,N_2640);
nor U3474 (N_3474,N_2049,N_2443);
nand U3475 (N_3475,N_2300,N_1910);
nor U3476 (N_3476,N_2497,N_2488);
or U3477 (N_3477,N_1551,N_1916);
or U3478 (N_3478,N_2413,N_2261);
and U3479 (N_3479,N_2434,N_2807);
or U3480 (N_3480,N_1855,N_2333);
nand U3481 (N_3481,N_2274,N_2958);
xor U3482 (N_3482,N_1960,N_1573);
nand U3483 (N_3483,N_1914,N_2961);
and U3484 (N_3484,N_1516,N_1805);
nand U3485 (N_3485,N_2952,N_2802);
and U3486 (N_3486,N_2046,N_2861);
and U3487 (N_3487,N_2245,N_2483);
xnor U3488 (N_3488,N_1761,N_2356);
and U3489 (N_3489,N_2017,N_1513);
or U3490 (N_3490,N_1699,N_2700);
nand U3491 (N_3491,N_1667,N_2165);
or U3492 (N_3492,N_2532,N_2107);
nand U3493 (N_3493,N_2213,N_2465);
nor U3494 (N_3494,N_1640,N_1571);
xor U3495 (N_3495,N_2680,N_2219);
xor U3496 (N_3496,N_2401,N_2476);
xnor U3497 (N_3497,N_2515,N_1564);
xor U3498 (N_3498,N_2346,N_1898);
xor U3499 (N_3499,N_2730,N_1622);
nand U3500 (N_3500,N_2829,N_1980);
xnor U3501 (N_3501,N_2386,N_2719);
nor U3502 (N_3502,N_2016,N_1602);
nand U3503 (N_3503,N_1638,N_2289);
nand U3504 (N_3504,N_2681,N_2456);
nor U3505 (N_3505,N_2027,N_1941);
nor U3506 (N_3506,N_2094,N_2674);
nor U3507 (N_3507,N_2694,N_2755);
and U3508 (N_3508,N_2286,N_1944);
nand U3509 (N_3509,N_2147,N_2702);
nand U3510 (N_3510,N_2503,N_2912);
nand U3511 (N_3511,N_2243,N_2984);
nand U3512 (N_3512,N_2756,N_2269);
nor U3513 (N_3513,N_2526,N_2235);
nor U3514 (N_3514,N_2941,N_2666);
xnor U3515 (N_3515,N_2555,N_1957);
and U3516 (N_3516,N_2926,N_1633);
xor U3517 (N_3517,N_2212,N_2379);
xor U3518 (N_3518,N_1945,N_2835);
nor U3519 (N_3519,N_2614,N_1565);
nor U3520 (N_3520,N_2466,N_2394);
nand U3521 (N_3521,N_1890,N_2918);
or U3522 (N_3522,N_2812,N_2625);
nand U3523 (N_3523,N_1696,N_2953);
nor U3524 (N_3524,N_2083,N_2390);
or U3525 (N_3525,N_2956,N_2889);
nand U3526 (N_3526,N_2852,N_2200);
and U3527 (N_3527,N_2718,N_1689);
xor U3528 (N_3528,N_2801,N_2160);
and U3529 (N_3529,N_1874,N_2188);
nand U3530 (N_3530,N_1708,N_1677);
nand U3531 (N_3531,N_2884,N_1508);
nand U3532 (N_3532,N_1897,N_1754);
xor U3533 (N_3533,N_1783,N_2995);
nand U3534 (N_3534,N_2683,N_2164);
or U3535 (N_3535,N_2782,N_1848);
nand U3536 (N_3536,N_1693,N_1919);
nand U3537 (N_3537,N_2388,N_2623);
or U3538 (N_3538,N_1650,N_1839);
and U3539 (N_3539,N_2781,N_2994);
or U3540 (N_3540,N_2586,N_1685);
nor U3541 (N_3541,N_2053,N_2149);
and U3542 (N_3542,N_1797,N_2034);
xor U3543 (N_3543,N_2203,N_2929);
xnor U3544 (N_3544,N_2750,N_1541);
xor U3545 (N_3545,N_2332,N_1556);
or U3546 (N_3546,N_2584,N_2140);
xnor U3547 (N_3547,N_2531,N_2325);
nor U3548 (N_3548,N_1629,N_1584);
nand U3549 (N_3549,N_1618,N_2705);
nand U3550 (N_3550,N_2181,N_2008);
and U3551 (N_3551,N_2805,N_2930);
or U3552 (N_3552,N_1893,N_1876);
xnor U3553 (N_3553,N_2548,N_1731);
or U3554 (N_3554,N_2005,N_2845);
nor U3555 (N_3555,N_2086,N_2063);
or U3556 (N_3556,N_1785,N_2449);
nand U3557 (N_3557,N_2338,N_1985);
xor U3558 (N_3558,N_2894,N_1531);
and U3559 (N_3559,N_1700,N_1742);
xor U3560 (N_3560,N_2940,N_2581);
nor U3561 (N_3561,N_2167,N_2178);
and U3562 (N_3562,N_2272,N_2150);
xor U3563 (N_3563,N_1694,N_1660);
nand U3564 (N_3564,N_2842,N_1885);
or U3565 (N_3565,N_2006,N_2717);
or U3566 (N_3566,N_2951,N_1851);
nand U3567 (N_3567,N_1793,N_1947);
or U3568 (N_3568,N_2974,N_1927);
xnor U3569 (N_3569,N_2803,N_2278);
nor U3570 (N_3570,N_2657,N_1998);
nand U3571 (N_3571,N_1620,N_1523);
or U3572 (N_3572,N_1924,N_1872);
nor U3573 (N_3573,N_1520,N_2860);
nand U3574 (N_3574,N_2636,N_2141);
nor U3575 (N_3575,N_1717,N_2048);
nand U3576 (N_3576,N_2059,N_1583);
and U3577 (N_3577,N_2317,N_1768);
nor U3578 (N_3578,N_2616,N_2768);
xnor U3579 (N_3579,N_2291,N_2763);
and U3580 (N_3580,N_2265,N_1908);
or U3581 (N_3581,N_1621,N_1566);
nand U3582 (N_3582,N_2450,N_2823);
nand U3583 (N_3583,N_2577,N_2846);
nor U3584 (N_3584,N_2469,N_1688);
xor U3585 (N_3585,N_1624,N_2964);
nor U3586 (N_3586,N_1845,N_2087);
or U3587 (N_3587,N_2786,N_2675);
and U3588 (N_3588,N_2528,N_1787);
or U3589 (N_3589,N_2029,N_1515);
or U3590 (N_3590,N_2949,N_2144);
nand U3591 (N_3591,N_1505,N_1918);
and U3592 (N_3592,N_2684,N_1983);
and U3593 (N_3593,N_2817,N_1530);
xor U3594 (N_3594,N_2070,N_1828);
or U3595 (N_3595,N_2985,N_1641);
or U3596 (N_3596,N_2710,N_2938);
xnor U3597 (N_3597,N_1804,N_1637);
xnor U3598 (N_3598,N_1766,N_1915);
xor U3599 (N_3599,N_2560,N_2980);
and U3600 (N_3600,N_1880,N_2644);
and U3601 (N_3601,N_1758,N_2195);
or U3602 (N_3602,N_1972,N_2507);
or U3603 (N_3603,N_2920,N_2850);
nand U3604 (N_3604,N_2406,N_2612);
xor U3605 (N_3605,N_1596,N_2156);
or U3606 (N_3606,N_1656,N_2535);
xor U3607 (N_3607,N_1586,N_1858);
xnor U3608 (N_3608,N_2525,N_2205);
nand U3609 (N_3609,N_2783,N_1900);
nand U3610 (N_3610,N_1734,N_2712);
nand U3611 (N_3611,N_2387,N_2501);
and U3612 (N_3612,N_1899,N_1865);
nor U3613 (N_3613,N_2121,N_2820);
nor U3614 (N_3614,N_2292,N_2706);
and U3615 (N_3615,N_2184,N_2095);
xor U3616 (N_3616,N_2254,N_2115);
nand U3617 (N_3617,N_2339,N_2173);
xor U3618 (N_3618,N_2760,N_2166);
nand U3619 (N_3619,N_2736,N_1567);
nor U3620 (N_3620,N_2815,N_2417);
or U3621 (N_3621,N_1733,N_2369);
or U3622 (N_3622,N_2814,N_2591);
nand U3623 (N_3623,N_2307,N_1746);
xnor U3624 (N_3624,N_1555,N_2295);
nand U3625 (N_3625,N_1987,N_2089);
and U3626 (N_3626,N_2370,N_2715);
and U3627 (N_3627,N_1867,N_2143);
nor U3628 (N_3628,N_2671,N_2981);
xnor U3629 (N_3629,N_2111,N_1988);
or U3630 (N_3630,N_2155,N_2827);
and U3631 (N_3631,N_1756,N_2976);
or U3632 (N_3632,N_2690,N_2627);
nor U3633 (N_3633,N_2799,N_2380);
nand U3634 (N_3634,N_2176,N_1612);
and U3635 (N_3635,N_2925,N_1871);
xor U3636 (N_3636,N_2924,N_2364);
and U3637 (N_3637,N_2101,N_2358);
or U3638 (N_3638,N_2152,N_2078);
or U3639 (N_3639,N_2775,N_1610);
xor U3640 (N_3640,N_1703,N_2109);
or U3641 (N_3641,N_2171,N_2819);
xnor U3642 (N_3642,N_1588,N_2090);
nand U3643 (N_3643,N_1651,N_1886);
nand U3644 (N_3644,N_2579,N_2547);
xor U3645 (N_3645,N_2293,N_2323);
or U3646 (N_3646,N_1713,N_2484);
nand U3647 (N_3647,N_2416,N_1820);
xor U3648 (N_3648,N_1691,N_2025);
and U3649 (N_3649,N_2603,N_2489);
nand U3650 (N_3650,N_2458,N_2723);
xor U3651 (N_3651,N_1570,N_2240);
xnor U3652 (N_3652,N_2654,N_2378);
nand U3653 (N_3653,N_2467,N_2751);
nor U3654 (N_3654,N_2076,N_2444);
nand U3655 (N_3655,N_2279,N_1534);
xnor U3656 (N_3656,N_2088,N_2151);
or U3657 (N_3657,N_2752,N_2576);
or U3658 (N_3658,N_2530,N_1953);
nand U3659 (N_3659,N_2673,N_1925);
nand U3660 (N_3660,N_2075,N_1632);
or U3661 (N_3661,N_2726,N_2491);
nand U3662 (N_3662,N_2208,N_2611);
or U3663 (N_3663,N_2772,N_2104);
nand U3664 (N_3664,N_1568,N_2055);
xor U3665 (N_3665,N_1749,N_2524);
nand U3666 (N_3666,N_2199,N_1795);
and U3667 (N_3667,N_1892,N_2892);
or U3668 (N_3668,N_2202,N_1506);
and U3669 (N_3669,N_2146,N_2256);
or U3670 (N_3670,N_2708,N_2905);
or U3671 (N_3671,N_2903,N_2893);
or U3672 (N_3672,N_2222,N_2733);
xnor U3673 (N_3673,N_1741,N_2856);
xor U3674 (N_3674,N_1964,N_1966);
or U3675 (N_3675,N_2907,N_2283);
xor U3676 (N_3676,N_2686,N_2373);
or U3677 (N_3677,N_1647,N_2137);
nand U3678 (N_3678,N_1999,N_2161);
and U3679 (N_3679,N_2516,N_2824);
nand U3680 (N_3680,N_2463,N_1934);
and U3681 (N_3681,N_2545,N_2179);
xnor U3682 (N_3682,N_2989,N_1521);
xnor U3683 (N_3683,N_2521,N_2872);
nor U3684 (N_3684,N_1698,N_1968);
nor U3685 (N_3685,N_2026,N_2619);
nand U3686 (N_3686,N_2753,N_2997);
and U3687 (N_3687,N_2010,N_2134);
xnor U3688 (N_3688,N_1719,N_2747);
and U3689 (N_3689,N_2797,N_2806);
and U3690 (N_3690,N_1548,N_2398);
xnor U3691 (N_3691,N_2312,N_1593);
xnor U3692 (N_3692,N_2228,N_2564);
or U3693 (N_3693,N_2653,N_1978);
and U3694 (N_3694,N_1990,N_2505);
nor U3695 (N_3695,N_2538,N_1654);
xor U3696 (N_3696,N_2795,N_2210);
and U3697 (N_3697,N_2537,N_1823);
nor U3698 (N_3698,N_1579,N_2602);
xnor U3699 (N_3699,N_2909,N_1800);
and U3700 (N_3700,N_1532,N_2145);
or U3701 (N_3701,N_2174,N_1815);
and U3702 (N_3702,N_1542,N_2230);
nand U3703 (N_3703,N_2740,N_2335);
or U3704 (N_3704,N_1920,N_2471);
nand U3705 (N_3705,N_2014,N_2979);
xor U3706 (N_3706,N_1617,N_1675);
and U3707 (N_3707,N_1833,N_2328);
nor U3708 (N_3708,N_2678,N_2001);
and U3709 (N_3709,N_2876,N_2192);
or U3710 (N_3710,N_2709,N_1526);
nand U3711 (N_3711,N_2425,N_1723);
xnor U3712 (N_3712,N_1595,N_2244);
nand U3713 (N_3713,N_1634,N_2950);
nand U3714 (N_3714,N_1527,N_2873);
and U3715 (N_3715,N_2183,N_2193);
nand U3716 (N_3716,N_1639,N_2914);
nand U3717 (N_3717,N_2556,N_2470);
nand U3718 (N_3718,N_2327,N_1771);
nand U3719 (N_3719,N_2632,N_1657);
xor U3720 (N_3720,N_2037,N_1753);
nor U3721 (N_3721,N_2276,N_2189);
and U3722 (N_3722,N_2935,N_2429);
nor U3723 (N_3723,N_2018,N_2211);
and U3724 (N_3724,N_1605,N_2030);
and U3725 (N_3725,N_1841,N_2946);
nand U3726 (N_3726,N_2568,N_2349);
xor U3727 (N_3727,N_2065,N_2761);
xnor U3728 (N_3728,N_1901,N_2153);
nor U3729 (N_3729,N_2689,N_2691);
xnor U3730 (N_3730,N_1789,N_1572);
and U3731 (N_3731,N_2773,N_2633);
nor U3732 (N_3732,N_2224,N_1986);
and U3733 (N_3733,N_2479,N_2800);
nor U3734 (N_3734,N_1810,N_2582);
nor U3735 (N_3735,N_2948,N_2502);
and U3736 (N_3736,N_2649,N_2227);
nand U3737 (N_3737,N_1682,N_1683);
and U3738 (N_3738,N_2288,N_1726);
nand U3739 (N_3739,N_2593,N_1580);
nand U3740 (N_3740,N_2928,N_2019);
nand U3741 (N_3741,N_2159,N_2848);
and U3742 (N_3742,N_1729,N_2891);
nand U3743 (N_3743,N_2831,N_2301);
or U3744 (N_3744,N_2656,N_1652);
nand U3745 (N_3745,N_2108,N_1663);
and U3746 (N_3746,N_2838,N_1504);
or U3747 (N_3747,N_1623,N_2126);
nand U3748 (N_3748,N_1575,N_1902);
xnor U3749 (N_3749,N_1578,N_2098);
xnor U3750 (N_3750,N_1895,N_2294);
or U3751 (N_3751,N_2707,N_2460);
or U3752 (N_3752,N_2919,N_1551);
xnor U3753 (N_3753,N_2776,N_2769);
xor U3754 (N_3754,N_2603,N_2679);
nand U3755 (N_3755,N_2263,N_2623);
xor U3756 (N_3756,N_2879,N_2667);
xor U3757 (N_3757,N_2991,N_1728);
xor U3758 (N_3758,N_1516,N_2420);
nor U3759 (N_3759,N_1597,N_2324);
or U3760 (N_3760,N_1696,N_2568);
nor U3761 (N_3761,N_2372,N_2471);
or U3762 (N_3762,N_1716,N_1516);
or U3763 (N_3763,N_2283,N_1725);
or U3764 (N_3764,N_2713,N_2611);
xnor U3765 (N_3765,N_2560,N_2989);
xor U3766 (N_3766,N_1751,N_2520);
or U3767 (N_3767,N_1811,N_1578);
nor U3768 (N_3768,N_2602,N_2980);
nor U3769 (N_3769,N_2231,N_2348);
nor U3770 (N_3770,N_1617,N_1668);
xnor U3771 (N_3771,N_1575,N_2266);
or U3772 (N_3772,N_2861,N_1835);
nor U3773 (N_3773,N_1669,N_2496);
xnor U3774 (N_3774,N_2139,N_2058);
nand U3775 (N_3775,N_1856,N_1868);
xnor U3776 (N_3776,N_2062,N_2836);
and U3777 (N_3777,N_1792,N_2092);
or U3778 (N_3778,N_1934,N_2477);
nand U3779 (N_3779,N_2791,N_2798);
xor U3780 (N_3780,N_2484,N_2281);
xnor U3781 (N_3781,N_1861,N_2743);
nor U3782 (N_3782,N_2058,N_2913);
nor U3783 (N_3783,N_2822,N_2463);
and U3784 (N_3784,N_1662,N_2337);
nand U3785 (N_3785,N_1835,N_2139);
and U3786 (N_3786,N_2160,N_1880);
nor U3787 (N_3787,N_2899,N_2741);
nor U3788 (N_3788,N_2853,N_2249);
nor U3789 (N_3789,N_1669,N_2988);
or U3790 (N_3790,N_1535,N_1637);
and U3791 (N_3791,N_2692,N_2339);
or U3792 (N_3792,N_2130,N_1948);
nand U3793 (N_3793,N_1693,N_2563);
and U3794 (N_3794,N_2940,N_2865);
nor U3795 (N_3795,N_2849,N_2243);
nand U3796 (N_3796,N_1980,N_2790);
nand U3797 (N_3797,N_2530,N_2579);
nand U3798 (N_3798,N_2813,N_2156);
xor U3799 (N_3799,N_1954,N_2189);
nand U3800 (N_3800,N_2121,N_1828);
and U3801 (N_3801,N_2169,N_2520);
nor U3802 (N_3802,N_2405,N_2629);
nand U3803 (N_3803,N_2592,N_1561);
xor U3804 (N_3804,N_2800,N_1681);
or U3805 (N_3805,N_2610,N_1813);
nand U3806 (N_3806,N_2509,N_2403);
nand U3807 (N_3807,N_2377,N_1982);
xnor U3808 (N_3808,N_2724,N_2054);
nor U3809 (N_3809,N_2519,N_2748);
and U3810 (N_3810,N_2381,N_2749);
nand U3811 (N_3811,N_2450,N_1656);
and U3812 (N_3812,N_2918,N_2427);
or U3813 (N_3813,N_1710,N_1750);
xor U3814 (N_3814,N_1680,N_2839);
and U3815 (N_3815,N_2818,N_2978);
nand U3816 (N_3816,N_1996,N_2109);
and U3817 (N_3817,N_1820,N_2494);
or U3818 (N_3818,N_2483,N_2326);
nor U3819 (N_3819,N_2031,N_2227);
nand U3820 (N_3820,N_1962,N_2671);
xor U3821 (N_3821,N_2764,N_1502);
or U3822 (N_3822,N_1716,N_2224);
nor U3823 (N_3823,N_1720,N_1556);
nand U3824 (N_3824,N_1751,N_2249);
and U3825 (N_3825,N_1843,N_1513);
xor U3826 (N_3826,N_2954,N_2592);
xor U3827 (N_3827,N_1532,N_2188);
nand U3828 (N_3828,N_1791,N_2312);
and U3829 (N_3829,N_2638,N_2364);
nor U3830 (N_3830,N_1885,N_2031);
xor U3831 (N_3831,N_1714,N_2537);
or U3832 (N_3832,N_1791,N_1598);
or U3833 (N_3833,N_2789,N_2884);
or U3834 (N_3834,N_2733,N_2252);
nor U3835 (N_3835,N_2524,N_1625);
and U3836 (N_3836,N_1864,N_1996);
xnor U3837 (N_3837,N_1662,N_1858);
and U3838 (N_3838,N_2415,N_1785);
and U3839 (N_3839,N_2206,N_2897);
and U3840 (N_3840,N_2371,N_1701);
xor U3841 (N_3841,N_2388,N_2386);
or U3842 (N_3842,N_2174,N_1764);
nor U3843 (N_3843,N_1632,N_2719);
xnor U3844 (N_3844,N_2151,N_2467);
xor U3845 (N_3845,N_2618,N_2885);
and U3846 (N_3846,N_2577,N_2924);
or U3847 (N_3847,N_2202,N_1698);
xor U3848 (N_3848,N_2244,N_2893);
and U3849 (N_3849,N_1620,N_2826);
nand U3850 (N_3850,N_2991,N_2836);
nor U3851 (N_3851,N_2969,N_2807);
nor U3852 (N_3852,N_2239,N_2141);
xor U3853 (N_3853,N_2682,N_1536);
nor U3854 (N_3854,N_2723,N_1852);
or U3855 (N_3855,N_1753,N_1530);
nand U3856 (N_3856,N_2930,N_2252);
nand U3857 (N_3857,N_2277,N_2534);
nor U3858 (N_3858,N_2642,N_2189);
xor U3859 (N_3859,N_1531,N_2149);
or U3860 (N_3860,N_1545,N_1802);
and U3861 (N_3861,N_1556,N_2962);
and U3862 (N_3862,N_2315,N_2033);
nand U3863 (N_3863,N_2299,N_1816);
nor U3864 (N_3864,N_2464,N_1745);
nand U3865 (N_3865,N_2306,N_2657);
nor U3866 (N_3866,N_2932,N_2876);
nor U3867 (N_3867,N_1961,N_2336);
and U3868 (N_3868,N_2109,N_2292);
or U3869 (N_3869,N_1813,N_1730);
xor U3870 (N_3870,N_1771,N_2998);
xnor U3871 (N_3871,N_2780,N_2414);
nor U3872 (N_3872,N_1912,N_1772);
and U3873 (N_3873,N_2466,N_2191);
or U3874 (N_3874,N_2394,N_2487);
and U3875 (N_3875,N_1537,N_2839);
nand U3876 (N_3876,N_2482,N_1701);
and U3877 (N_3877,N_2741,N_2554);
or U3878 (N_3878,N_2175,N_2476);
xnor U3879 (N_3879,N_1696,N_2033);
or U3880 (N_3880,N_1722,N_2895);
nor U3881 (N_3881,N_2247,N_2834);
or U3882 (N_3882,N_1738,N_1530);
and U3883 (N_3883,N_2902,N_1754);
xor U3884 (N_3884,N_2836,N_2667);
nor U3885 (N_3885,N_2967,N_2589);
and U3886 (N_3886,N_1732,N_2896);
nor U3887 (N_3887,N_2156,N_1619);
xnor U3888 (N_3888,N_1946,N_1756);
nor U3889 (N_3889,N_2157,N_2801);
nand U3890 (N_3890,N_1665,N_1505);
nor U3891 (N_3891,N_2017,N_1862);
or U3892 (N_3892,N_2844,N_2002);
nor U3893 (N_3893,N_1837,N_2701);
xnor U3894 (N_3894,N_1620,N_2642);
xnor U3895 (N_3895,N_2930,N_1719);
or U3896 (N_3896,N_2726,N_2083);
nand U3897 (N_3897,N_2158,N_1552);
nand U3898 (N_3898,N_2944,N_2787);
or U3899 (N_3899,N_2582,N_1559);
nor U3900 (N_3900,N_2708,N_2529);
or U3901 (N_3901,N_2611,N_1698);
xor U3902 (N_3902,N_2688,N_2384);
nand U3903 (N_3903,N_1868,N_2319);
nor U3904 (N_3904,N_2291,N_1749);
nand U3905 (N_3905,N_2383,N_1517);
and U3906 (N_3906,N_2133,N_2850);
xor U3907 (N_3907,N_2007,N_2722);
and U3908 (N_3908,N_2947,N_2891);
xor U3909 (N_3909,N_1579,N_1627);
nor U3910 (N_3910,N_2312,N_2710);
or U3911 (N_3911,N_1750,N_2344);
or U3912 (N_3912,N_1789,N_1972);
and U3913 (N_3913,N_2023,N_2523);
nor U3914 (N_3914,N_1865,N_2437);
and U3915 (N_3915,N_1964,N_1711);
and U3916 (N_3916,N_2246,N_2679);
nand U3917 (N_3917,N_1889,N_2741);
and U3918 (N_3918,N_2760,N_1771);
nor U3919 (N_3919,N_2002,N_2469);
and U3920 (N_3920,N_2734,N_1946);
or U3921 (N_3921,N_1734,N_1663);
xnor U3922 (N_3922,N_1820,N_2038);
nand U3923 (N_3923,N_2734,N_2781);
or U3924 (N_3924,N_2298,N_2617);
xor U3925 (N_3925,N_1991,N_1846);
and U3926 (N_3926,N_1891,N_2167);
or U3927 (N_3927,N_2437,N_1721);
or U3928 (N_3928,N_1659,N_1661);
or U3929 (N_3929,N_1523,N_2995);
nand U3930 (N_3930,N_2492,N_2168);
nand U3931 (N_3931,N_2087,N_1850);
and U3932 (N_3932,N_1981,N_2589);
nor U3933 (N_3933,N_2381,N_2088);
xor U3934 (N_3934,N_2721,N_2189);
or U3935 (N_3935,N_1538,N_1790);
nand U3936 (N_3936,N_2088,N_2686);
nand U3937 (N_3937,N_1930,N_2604);
nand U3938 (N_3938,N_2828,N_1668);
and U3939 (N_3939,N_2531,N_2406);
nor U3940 (N_3940,N_2754,N_2865);
nor U3941 (N_3941,N_1785,N_2571);
or U3942 (N_3942,N_2549,N_2071);
or U3943 (N_3943,N_2796,N_2553);
xnor U3944 (N_3944,N_2587,N_2905);
nor U3945 (N_3945,N_2708,N_1597);
and U3946 (N_3946,N_2245,N_2201);
or U3947 (N_3947,N_2676,N_1885);
nor U3948 (N_3948,N_2172,N_2059);
xor U3949 (N_3949,N_2028,N_2449);
nor U3950 (N_3950,N_2248,N_2932);
and U3951 (N_3951,N_1549,N_2009);
or U3952 (N_3952,N_2187,N_1672);
nand U3953 (N_3953,N_2086,N_2575);
and U3954 (N_3954,N_1504,N_1900);
nor U3955 (N_3955,N_2392,N_2717);
and U3956 (N_3956,N_2358,N_2087);
or U3957 (N_3957,N_1543,N_1717);
or U3958 (N_3958,N_2125,N_2398);
nand U3959 (N_3959,N_1979,N_2187);
or U3960 (N_3960,N_2084,N_2622);
nor U3961 (N_3961,N_2231,N_2497);
or U3962 (N_3962,N_2533,N_2312);
or U3963 (N_3963,N_2893,N_1916);
xor U3964 (N_3964,N_1766,N_1805);
and U3965 (N_3965,N_2692,N_2146);
or U3966 (N_3966,N_2985,N_1774);
nor U3967 (N_3967,N_2203,N_1637);
xnor U3968 (N_3968,N_2880,N_2943);
xnor U3969 (N_3969,N_1568,N_2124);
or U3970 (N_3970,N_2383,N_2841);
and U3971 (N_3971,N_2792,N_2761);
nor U3972 (N_3972,N_2717,N_2590);
and U3973 (N_3973,N_1837,N_2267);
nand U3974 (N_3974,N_2577,N_1916);
nand U3975 (N_3975,N_2659,N_2664);
nor U3976 (N_3976,N_1961,N_2963);
xnor U3977 (N_3977,N_2189,N_2928);
nand U3978 (N_3978,N_2334,N_1727);
or U3979 (N_3979,N_2275,N_2625);
and U3980 (N_3980,N_2208,N_1832);
nand U3981 (N_3981,N_2654,N_1821);
nand U3982 (N_3982,N_2056,N_1503);
or U3983 (N_3983,N_1612,N_2915);
and U3984 (N_3984,N_2575,N_1652);
xnor U3985 (N_3985,N_2050,N_2942);
xnor U3986 (N_3986,N_1957,N_2296);
nor U3987 (N_3987,N_2843,N_2876);
and U3988 (N_3988,N_2731,N_2636);
or U3989 (N_3989,N_1587,N_2210);
and U3990 (N_3990,N_2956,N_2765);
or U3991 (N_3991,N_2287,N_2682);
or U3992 (N_3992,N_1705,N_2186);
and U3993 (N_3993,N_1908,N_2268);
nand U3994 (N_3994,N_2491,N_1805);
and U3995 (N_3995,N_2254,N_1627);
and U3996 (N_3996,N_1800,N_2486);
nor U3997 (N_3997,N_2633,N_1788);
nand U3998 (N_3998,N_2230,N_2995);
nor U3999 (N_3999,N_2256,N_2519);
nand U4000 (N_4000,N_1770,N_2714);
and U4001 (N_4001,N_2837,N_1622);
xor U4002 (N_4002,N_2954,N_2938);
and U4003 (N_4003,N_2553,N_2613);
nand U4004 (N_4004,N_1865,N_2501);
nand U4005 (N_4005,N_2404,N_2211);
or U4006 (N_4006,N_1799,N_1977);
and U4007 (N_4007,N_2062,N_2225);
and U4008 (N_4008,N_2172,N_1658);
and U4009 (N_4009,N_2466,N_2685);
or U4010 (N_4010,N_1993,N_2464);
nor U4011 (N_4011,N_2722,N_2460);
or U4012 (N_4012,N_2958,N_2983);
or U4013 (N_4013,N_2043,N_2634);
and U4014 (N_4014,N_1881,N_2405);
and U4015 (N_4015,N_2526,N_2514);
nor U4016 (N_4016,N_1508,N_2702);
nand U4017 (N_4017,N_1723,N_2891);
nor U4018 (N_4018,N_1985,N_1932);
nor U4019 (N_4019,N_2734,N_2617);
nand U4020 (N_4020,N_2934,N_2009);
nor U4021 (N_4021,N_1901,N_2254);
nand U4022 (N_4022,N_2407,N_1579);
nor U4023 (N_4023,N_2014,N_1580);
or U4024 (N_4024,N_2313,N_2460);
nor U4025 (N_4025,N_1516,N_2502);
nor U4026 (N_4026,N_1697,N_2099);
xor U4027 (N_4027,N_1660,N_2452);
or U4028 (N_4028,N_2426,N_2503);
nor U4029 (N_4029,N_2505,N_2131);
nand U4030 (N_4030,N_2139,N_2746);
nand U4031 (N_4031,N_1960,N_2583);
nand U4032 (N_4032,N_2473,N_2613);
nand U4033 (N_4033,N_2458,N_2447);
or U4034 (N_4034,N_1752,N_2970);
or U4035 (N_4035,N_2546,N_1865);
xnor U4036 (N_4036,N_1968,N_2022);
nand U4037 (N_4037,N_1878,N_2781);
nor U4038 (N_4038,N_2393,N_1580);
nor U4039 (N_4039,N_2892,N_1808);
xor U4040 (N_4040,N_2867,N_2083);
xnor U4041 (N_4041,N_2336,N_2933);
nor U4042 (N_4042,N_2994,N_2155);
nor U4043 (N_4043,N_1930,N_2925);
nor U4044 (N_4044,N_2336,N_2324);
xnor U4045 (N_4045,N_1791,N_2731);
and U4046 (N_4046,N_1698,N_2816);
nor U4047 (N_4047,N_2999,N_1514);
or U4048 (N_4048,N_2598,N_2960);
nand U4049 (N_4049,N_2827,N_2784);
or U4050 (N_4050,N_1646,N_2896);
nand U4051 (N_4051,N_2946,N_1984);
nor U4052 (N_4052,N_2435,N_2630);
and U4053 (N_4053,N_1835,N_2879);
nor U4054 (N_4054,N_1892,N_2027);
xnor U4055 (N_4055,N_2156,N_1610);
or U4056 (N_4056,N_2679,N_2983);
and U4057 (N_4057,N_1796,N_2932);
nor U4058 (N_4058,N_1592,N_2297);
and U4059 (N_4059,N_1783,N_2330);
xor U4060 (N_4060,N_2692,N_2329);
nor U4061 (N_4061,N_2696,N_2821);
xor U4062 (N_4062,N_1724,N_1727);
xor U4063 (N_4063,N_1936,N_2953);
and U4064 (N_4064,N_2003,N_1555);
xnor U4065 (N_4065,N_2386,N_2156);
nor U4066 (N_4066,N_2021,N_1645);
nor U4067 (N_4067,N_2444,N_2598);
xnor U4068 (N_4068,N_2358,N_1716);
nor U4069 (N_4069,N_2222,N_2411);
nand U4070 (N_4070,N_2484,N_1839);
nor U4071 (N_4071,N_2777,N_2701);
nand U4072 (N_4072,N_2792,N_2402);
nor U4073 (N_4073,N_2734,N_1890);
or U4074 (N_4074,N_1644,N_2832);
nand U4075 (N_4075,N_1591,N_2959);
or U4076 (N_4076,N_2055,N_1869);
nor U4077 (N_4077,N_2639,N_2225);
or U4078 (N_4078,N_2645,N_2051);
nor U4079 (N_4079,N_2213,N_1785);
and U4080 (N_4080,N_2770,N_2650);
nand U4081 (N_4081,N_2092,N_2441);
and U4082 (N_4082,N_2822,N_2211);
nor U4083 (N_4083,N_2457,N_2224);
xor U4084 (N_4084,N_2643,N_1896);
nand U4085 (N_4085,N_1605,N_1937);
nor U4086 (N_4086,N_1932,N_2669);
nor U4087 (N_4087,N_2637,N_2401);
xor U4088 (N_4088,N_2961,N_2241);
xor U4089 (N_4089,N_2784,N_2040);
or U4090 (N_4090,N_2099,N_1584);
xnor U4091 (N_4091,N_1658,N_1914);
nor U4092 (N_4092,N_1827,N_2737);
and U4093 (N_4093,N_2987,N_2834);
or U4094 (N_4094,N_2809,N_2929);
nor U4095 (N_4095,N_2132,N_2395);
and U4096 (N_4096,N_2640,N_1534);
and U4097 (N_4097,N_2881,N_1559);
or U4098 (N_4098,N_2864,N_1806);
nor U4099 (N_4099,N_1652,N_2639);
or U4100 (N_4100,N_1796,N_2279);
or U4101 (N_4101,N_2103,N_2871);
or U4102 (N_4102,N_1634,N_1694);
xnor U4103 (N_4103,N_2990,N_2664);
nand U4104 (N_4104,N_1872,N_2736);
and U4105 (N_4105,N_1547,N_2776);
nand U4106 (N_4106,N_2523,N_2013);
and U4107 (N_4107,N_2528,N_2420);
xor U4108 (N_4108,N_2312,N_2908);
xor U4109 (N_4109,N_2200,N_2456);
xnor U4110 (N_4110,N_2593,N_2494);
nor U4111 (N_4111,N_1771,N_2027);
or U4112 (N_4112,N_2851,N_1751);
or U4113 (N_4113,N_1651,N_2813);
or U4114 (N_4114,N_2472,N_2167);
xnor U4115 (N_4115,N_2321,N_1949);
nand U4116 (N_4116,N_2992,N_2914);
xor U4117 (N_4117,N_2742,N_2168);
and U4118 (N_4118,N_2801,N_1585);
xnor U4119 (N_4119,N_2810,N_2795);
nor U4120 (N_4120,N_1708,N_2470);
nor U4121 (N_4121,N_2444,N_2211);
nand U4122 (N_4122,N_2519,N_2917);
nand U4123 (N_4123,N_2935,N_2679);
nand U4124 (N_4124,N_2740,N_2663);
and U4125 (N_4125,N_2219,N_2134);
nand U4126 (N_4126,N_1792,N_1796);
or U4127 (N_4127,N_2888,N_2432);
or U4128 (N_4128,N_2897,N_2156);
and U4129 (N_4129,N_2860,N_1688);
nor U4130 (N_4130,N_2369,N_2965);
nor U4131 (N_4131,N_1659,N_2557);
nand U4132 (N_4132,N_2365,N_1831);
or U4133 (N_4133,N_1665,N_2497);
or U4134 (N_4134,N_2912,N_2947);
nand U4135 (N_4135,N_1571,N_2906);
or U4136 (N_4136,N_2382,N_2719);
xor U4137 (N_4137,N_2645,N_2971);
and U4138 (N_4138,N_1850,N_2217);
nand U4139 (N_4139,N_1785,N_2841);
and U4140 (N_4140,N_1627,N_2884);
and U4141 (N_4141,N_2532,N_2337);
nor U4142 (N_4142,N_2036,N_1682);
nor U4143 (N_4143,N_2429,N_2668);
nor U4144 (N_4144,N_2984,N_2609);
nor U4145 (N_4145,N_2762,N_1846);
nand U4146 (N_4146,N_1624,N_2579);
or U4147 (N_4147,N_2316,N_1609);
xor U4148 (N_4148,N_2338,N_2404);
xor U4149 (N_4149,N_1599,N_2353);
or U4150 (N_4150,N_2419,N_1536);
nor U4151 (N_4151,N_2590,N_1927);
nor U4152 (N_4152,N_2656,N_1625);
xnor U4153 (N_4153,N_2961,N_2944);
and U4154 (N_4154,N_2831,N_2333);
nand U4155 (N_4155,N_2785,N_2218);
nor U4156 (N_4156,N_2158,N_2337);
nor U4157 (N_4157,N_1727,N_2655);
and U4158 (N_4158,N_2975,N_1776);
xnor U4159 (N_4159,N_1821,N_2135);
xor U4160 (N_4160,N_2131,N_1975);
or U4161 (N_4161,N_1683,N_2710);
or U4162 (N_4162,N_2774,N_1619);
xnor U4163 (N_4163,N_2144,N_2781);
xnor U4164 (N_4164,N_2285,N_2060);
or U4165 (N_4165,N_2195,N_1665);
nor U4166 (N_4166,N_2693,N_1682);
or U4167 (N_4167,N_1937,N_2486);
and U4168 (N_4168,N_2260,N_1624);
or U4169 (N_4169,N_1639,N_2468);
or U4170 (N_4170,N_2839,N_1787);
nand U4171 (N_4171,N_2851,N_2489);
and U4172 (N_4172,N_2756,N_2065);
nand U4173 (N_4173,N_2438,N_2354);
or U4174 (N_4174,N_2641,N_2413);
nor U4175 (N_4175,N_2596,N_2176);
nor U4176 (N_4176,N_1797,N_2391);
or U4177 (N_4177,N_2763,N_2015);
or U4178 (N_4178,N_2480,N_1865);
nor U4179 (N_4179,N_2852,N_1870);
or U4180 (N_4180,N_1522,N_2035);
xnor U4181 (N_4181,N_2327,N_2488);
xor U4182 (N_4182,N_1913,N_2057);
and U4183 (N_4183,N_2498,N_2410);
nand U4184 (N_4184,N_2564,N_2014);
and U4185 (N_4185,N_1652,N_2584);
and U4186 (N_4186,N_2852,N_2243);
nor U4187 (N_4187,N_1713,N_2840);
nor U4188 (N_4188,N_1584,N_2596);
or U4189 (N_4189,N_2350,N_2314);
or U4190 (N_4190,N_2899,N_1843);
xor U4191 (N_4191,N_2166,N_2240);
nand U4192 (N_4192,N_1704,N_2418);
xor U4193 (N_4193,N_2381,N_2492);
and U4194 (N_4194,N_1869,N_2842);
xnor U4195 (N_4195,N_2328,N_2839);
and U4196 (N_4196,N_1540,N_2072);
nor U4197 (N_4197,N_2035,N_2891);
and U4198 (N_4198,N_2400,N_1574);
nand U4199 (N_4199,N_2056,N_1587);
nand U4200 (N_4200,N_2591,N_2473);
xnor U4201 (N_4201,N_2848,N_2455);
nand U4202 (N_4202,N_2652,N_2274);
and U4203 (N_4203,N_1686,N_1774);
xnor U4204 (N_4204,N_2239,N_1634);
or U4205 (N_4205,N_2083,N_1647);
nor U4206 (N_4206,N_2175,N_2559);
xnor U4207 (N_4207,N_2259,N_2616);
and U4208 (N_4208,N_1739,N_2631);
xnor U4209 (N_4209,N_1512,N_1950);
or U4210 (N_4210,N_2272,N_2517);
or U4211 (N_4211,N_1882,N_2042);
xnor U4212 (N_4212,N_2787,N_2000);
nor U4213 (N_4213,N_1879,N_2950);
nor U4214 (N_4214,N_2774,N_1809);
nand U4215 (N_4215,N_2973,N_2378);
nand U4216 (N_4216,N_2526,N_2793);
nor U4217 (N_4217,N_2770,N_1778);
nor U4218 (N_4218,N_1746,N_2717);
or U4219 (N_4219,N_1942,N_2072);
nor U4220 (N_4220,N_2309,N_2541);
nor U4221 (N_4221,N_2718,N_1697);
nand U4222 (N_4222,N_1620,N_1530);
nand U4223 (N_4223,N_2392,N_2218);
and U4224 (N_4224,N_2237,N_2279);
or U4225 (N_4225,N_2885,N_2690);
or U4226 (N_4226,N_1611,N_2941);
and U4227 (N_4227,N_1894,N_2302);
and U4228 (N_4228,N_2208,N_2188);
or U4229 (N_4229,N_2783,N_2346);
xor U4230 (N_4230,N_2613,N_2045);
or U4231 (N_4231,N_1816,N_2156);
or U4232 (N_4232,N_2550,N_1956);
xnor U4233 (N_4233,N_2914,N_2305);
nor U4234 (N_4234,N_1680,N_1963);
or U4235 (N_4235,N_2375,N_1695);
nand U4236 (N_4236,N_1607,N_1667);
and U4237 (N_4237,N_2079,N_2556);
or U4238 (N_4238,N_2540,N_2887);
or U4239 (N_4239,N_1983,N_2183);
and U4240 (N_4240,N_2745,N_1711);
or U4241 (N_4241,N_1638,N_2934);
xor U4242 (N_4242,N_2225,N_1801);
nand U4243 (N_4243,N_2575,N_1613);
xor U4244 (N_4244,N_2746,N_1820);
nor U4245 (N_4245,N_1644,N_2064);
and U4246 (N_4246,N_1620,N_1725);
nand U4247 (N_4247,N_2902,N_2403);
nand U4248 (N_4248,N_1583,N_2216);
and U4249 (N_4249,N_2951,N_2394);
and U4250 (N_4250,N_1716,N_2545);
nand U4251 (N_4251,N_2940,N_1583);
nor U4252 (N_4252,N_2926,N_2305);
or U4253 (N_4253,N_2555,N_1999);
or U4254 (N_4254,N_1892,N_2816);
and U4255 (N_4255,N_2277,N_1661);
or U4256 (N_4256,N_2273,N_2622);
and U4257 (N_4257,N_1921,N_1845);
nor U4258 (N_4258,N_1685,N_2287);
or U4259 (N_4259,N_1958,N_2678);
and U4260 (N_4260,N_2191,N_1830);
and U4261 (N_4261,N_2294,N_1568);
nor U4262 (N_4262,N_2132,N_2804);
and U4263 (N_4263,N_1609,N_2257);
and U4264 (N_4264,N_2922,N_2189);
nand U4265 (N_4265,N_2715,N_2047);
nand U4266 (N_4266,N_2681,N_2191);
and U4267 (N_4267,N_1587,N_1556);
nor U4268 (N_4268,N_2675,N_1649);
nand U4269 (N_4269,N_2664,N_2909);
or U4270 (N_4270,N_2841,N_1794);
nand U4271 (N_4271,N_2731,N_2549);
nand U4272 (N_4272,N_1685,N_2083);
or U4273 (N_4273,N_1795,N_2058);
xor U4274 (N_4274,N_2846,N_2573);
nand U4275 (N_4275,N_2068,N_1951);
nor U4276 (N_4276,N_2874,N_2673);
nor U4277 (N_4277,N_1667,N_2417);
xnor U4278 (N_4278,N_2265,N_2433);
and U4279 (N_4279,N_2079,N_2719);
and U4280 (N_4280,N_1800,N_2830);
xnor U4281 (N_4281,N_1691,N_2808);
nor U4282 (N_4282,N_2902,N_2125);
nand U4283 (N_4283,N_1924,N_2072);
nor U4284 (N_4284,N_2386,N_1776);
or U4285 (N_4285,N_2795,N_2792);
or U4286 (N_4286,N_2720,N_2889);
and U4287 (N_4287,N_1839,N_2374);
and U4288 (N_4288,N_2307,N_1727);
or U4289 (N_4289,N_2030,N_1641);
or U4290 (N_4290,N_1713,N_2825);
or U4291 (N_4291,N_1824,N_2211);
xor U4292 (N_4292,N_2458,N_1971);
or U4293 (N_4293,N_2620,N_1724);
xor U4294 (N_4294,N_2961,N_1505);
nand U4295 (N_4295,N_2463,N_2819);
or U4296 (N_4296,N_2836,N_2005);
xor U4297 (N_4297,N_1651,N_2891);
nor U4298 (N_4298,N_2853,N_2951);
nand U4299 (N_4299,N_2725,N_1880);
nor U4300 (N_4300,N_2994,N_2561);
nor U4301 (N_4301,N_1521,N_1927);
nand U4302 (N_4302,N_2267,N_2487);
nand U4303 (N_4303,N_2054,N_2767);
nor U4304 (N_4304,N_2698,N_2715);
or U4305 (N_4305,N_2447,N_2731);
or U4306 (N_4306,N_2850,N_2910);
or U4307 (N_4307,N_2528,N_2384);
nand U4308 (N_4308,N_1767,N_2301);
nor U4309 (N_4309,N_1668,N_2767);
or U4310 (N_4310,N_2377,N_1973);
xor U4311 (N_4311,N_2804,N_1545);
and U4312 (N_4312,N_1708,N_2956);
xor U4313 (N_4313,N_2707,N_1925);
nor U4314 (N_4314,N_2782,N_1611);
xor U4315 (N_4315,N_2597,N_2071);
xor U4316 (N_4316,N_2700,N_1700);
nand U4317 (N_4317,N_1580,N_2249);
and U4318 (N_4318,N_2919,N_1566);
xor U4319 (N_4319,N_2905,N_2866);
nor U4320 (N_4320,N_2490,N_2411);
and U4321 (N_4321,N_1889,N_2179);
nand U4322 (N_4322,N_2253,N_2274);
xor U4323 (N_4323,N_1794,N_2383);
nor U4324 (N_4324,N_2642,N_2296);
nor U4325 (N_4325,N_2497,N_2752);
or U4326 (N_4326,N_2208,N_2916);
xor U4327 (N_4327,N_2440,N_1900);
nand U4328 (N_4328,N_1815,N_2300);
nand U4329 (N_4329,N_2019,N_2695);
nor U4330 (N_4330,N_1963,N_1796);
or U4331 (N_4331,N_2280,N_2684);
or U4332 (N_4332,N_2932,N_1527);
nor U4333 (N_4333,N_1800,N_2820);
nor U4334 (N_4334,N_2186,N_1938);
or U4335 (N_4335,N_2886,N_2910);
xor U4336 (N_4336,N_2724,N_2454);
nand U4337 (N_4337,N_2488,N_2912);
nor U4338 (N_4338,N_2027,N_2130);
nand U4339 (N_4339,N_1596,N_2495);
xnor U4340 (N_4340,N_2722,N_1566);
xnor U4341 (N_4341,N_1761,N_2151);
or U4342 (N_4342,N_2174,N_1970);
or U4343 (N_4343,N_1615,N_2752);
and U4344 (N_4344,N_1710,N_1535);
and U4345 (N_4345,N_1790,N_1763);
and U4346 (N_4346,N_2161,N_2197);
or U4347 (N_4347,N_2951,N_2442);
xnor U4348 (N_4348,N_2487,N_2988);
or U4349 (N_4349,N_2485,N_2420);
and U4350 (N_4350,N_1690,N_2858);
nand U4351 (N_4351,N_1549,N_2031);
or U4352 (N_4352,N_2910,N_1549);
and U4353 (N_4353,N_2640,N_2920);
xnor U4354 (N_4354,N_2216,N_2885);
or U4355 (N_4355,N_2687,N_2506);
and U4356 (N_4356,N_2572,N_2148);
nor U4357 (N_4357,N_2745,N_2852);
xnor U4358 (N_4358,N_1962,N_1740);
nor U4359 (N_4359,N_2832,N_2424);
nor U4360 (N_4360,N_1767,N_2164);
nand U4361 (N_4361,N_2855,N_2884);
xor U4362 (N_4362,N_2192,N_2500);
nor U4363 (N_4363,N_1680,N_2437);
or U4364 (N_4364,N_2496,N_1982);
or U4365 (N_4365,N_1528,N_2475);
xnor U4366 (N_4366,N_2065,N_2538);
nor U4367 (N_4367,N_2109,N_2729);
and U4368 (N_4368,N_2691,N_2510);
or U4369 (N_4369,N_2545,N_2601);
nand U4370 (N_4370,N_2807,N_1518);
or U4371 (N_4371,N_1566,N_2353);
nand U4372 (N_4372,N_2251,N_2849);
nor U4373 (N_4373,N_1527,N_1946);
or U4374 (N_4374,N_2719,N_2822);
or U4375 (N_4375,N_2771,N_1505);
and U4376 (N_4376,N_1733,N_1509);
and U4377 (N_4377,N_2749,N_2012);
and U4378 (N_4378,N_1663,N_2230);
xnor U4379 (N_4379,N_1506,N_1937);
nand U4380 (N_4380,N_2416,N_2712);
xnor U4381 (N_4381,N_2455,N_2123);
xnor U4382 (N_4382,N_1527,N_2911);
nand U4383 (N_4383,N_2692,N_2828);
nand U4384 (N_4384,N_2209,N_1514);
nand U4385 (N_4385,N_2738,N_2779);
xnor U4386 (N_4386,N_2605,N_2691);
and U4387 (N_4387,N_2788,N_2567);
nor U4388 (N_4388,N_2415,N_1881);
nand U4389 (N_4389,N_2598,N_1760);
xor U4390 (N_4390,N_2943,N_2379);
nand U4391 (N_4391,N_2199,N_2372);
xor U4392 (N_4392,N_1924,N_2550);
and U4393 (N_4393,N_2242,N_2795);
nor U4394 (N_4394,N_2397,N_2850);
xor U4395 (N_4395,N_1667,N_1501);
nand U4396 (N_4396,N_1791,N_1759);
nor U4397 (N_4397,N_2700,N_2557);
xor U4398 (N_4398,N_2056,N_2874);
and U4399 (N_4399,N_2815,N_2719);
and U4400 (N_4400,N_2638,N_2206);
nor U4401 (N_4401,N_2779,N_2439);
or U4402 (N_4402,N_2559,N_2978);
or U4403 (N_4403,N_2069,N_2904);
xor U4404 (N_4404,N_2380,N_2082);
nor U4405 (N_4405,N_2334,N_2964);
nand U4406 (N_4406,N_1581,N_2926);
nor U4407 (N_4407,N_2418,N_2732);
or U4408 (N_4408,N_2049,N_2852);
xor U4409 (N_4409,N_2696,N_2187);
nor U4410 (N_4410,N_1931,N_1754);
or U4411 (N_4411,N_1760,N_2401);
nand U4412 (N_4412,N_2909,N_2679);
and U4413 (N_4413,N_2041,N_2878);
and U4414 (N_4414,N_2843,N_2977);
xor U4415 (N_4415,N_2235,N_1962);
and U4416 (N_4416,N_2329,N_2317);
and U4417 (N_4417,N_2919,N_1611);
xor U4418 (N_4418,N_2785,N_1583);
nor U4419 (N_4419,N_1515,N_2416);
xor U4420 (N_4420,N_1585,N_1850);
xnor U4421 (N_4421,N_2770,N_2677);
nand U4422 (N_4422,N_2393,N_2095);
or U4423 (N_4423,N_1692,N_2464);
or U4424 (N_4424,N_1621,N_1504);
nor U4425 (N_4425,N_2720,N_2611);
nor U4426 (N_4426,N_2901,N_2259);
nor U4427 (N_4427,N_2129,N_1814);
or U4428 (N_4428,N_2414,N_2427);
nand U4429 (N_4429,N_1636,N_2219);
nor U4430 (N_4430,N_2612,N_1617);
nor U4431 (N_4431,N_2598,N_1538);
nand U4432 (N_4432,N_2874,N_2219);
nand U4433 (N_4433,N_2636,N_2875);
nand U4434 (N_4434,N_2066,N_1699);
nand U4435 (N_4435,N_2335,N_2799);
nand U4436 (N_4436,N_1540,N_2629);
or U4437 (N_4437,N_2853,N_2392);
xor U4438 (N_4438,N_2838,N_1964);
nor U4439 (N_4439,N_2963,N_2139);
and U4440 (N_4440,N_2675,N_2522);
nor U4441 (N_4441,N_2693,N_2443);
nand U4442 (N_4442,N_2318,N_1581);
nand U4443 (N_4443,N_1890,N_2078);
and U4444 (N_4444,N_2816,N_2688);
or U4445 (N_4445,N_1753,N_2271);
nand U4446 (N_4446,N_2570,N_2683);
or U4447 (N_4447,N_2727,N_2690);
or U4448 (N_4448,N_2909,N_1658);
or U4449 (N_4449,N_2255,N_2260);
nand U4450 (N_4450,N_2020,N_1537);
nor U4451 (N_4451,N_1691,N_2163);
nor U4452 (N_4452,N_1750,N_2555);
xor U4453 (N_4453,N_2552,N_2557);
and U4454 (N_4454,N_2615,N_2829);
nor U4455 (N_4455,N_2012,N_2441);
and U4456 (N_4456,N_1736,N_2170);
xor U4457 (N_4457,N_2982,N_2234);
xnor U4458 (N_4458,N_1817,N_2665);
or U4459 (N_4459,N_2206,N_1670);
nor U4460 (N_4460,N_2549,N_2421);
nor U4461 (N_4461,N_2741,N_2232);
nor U4462 (N_4462,N_1970,N_1737);
nand U4463 (N_4463,N_2138,N_2470);
xor U4464 (N_4464,N_1587,N_2734);
and U4465 (N_4465,N_1777,N_2448);
nand U4466 (N_4466,N_2558,N_2834);
xor U4467 (N_4467,N_1768,N_2557);
and U4468 (N_4468,N_2562,N_2697);
nand U4469 (N_4469,N_2478,N_2458);
or U4470 (N_4470,N_2527,N_2913);
xnor U4471 (N_4471,N_1700,N_2228);
xnor U4472 (N_4472,N_1932,N_2264);
xnor U4473 (N_4473,N_2249,N_2477);
nor U4474 (N_4474,N_2710,N_2815);
nand U4475 (N_4475,N_2231,N_2903);
and U4476 (N_4476,N_2031,N_2546);
and U4477 (N_4477,N_1862,N_2787);
xnor U4478 (N_4478,N_2089,N_2758);
and U4479 (N_4479,N_2280,N_2974);
xnor U4480 (N_4480,N_2549,N_2677);
or U4481 (N_4481,N_2146,N_1998);
and U4482 (N_4482,N_2199,N_2561);
xnor U4483 (N_4483,N_2178,N_2895);
and U4484 (N_4484,N_2571,N_1791);
nand U4485 (N_4485,N_1553,N_1819);
or U4486 (N_4486,N_2377,N_1778);
or U4487 (N_4487,N_1914,N_2253);
xnor U4488 (N_4488,N_1908,N_2604);
nor U4489 (N_4489,N_2337,N_1854);
and U4490 (N_4490,N_1852,N_2073);
nor U4491 (N_4491,N_2438,N_2168);
and U4492 (N_4492,N_1843,N_2328);
xor U4493 (N_4493,N_1641,N_1747);
xnor U4494 (N_4494,N_1529,N_2834);
nand U4495 (N_4495,N_2126,N_2740);
and U4496 (N_4496,N_2027,N_1774);
and U4497 (N_4497,N_1652,N_2295);
or U4498 (N_4498,N_1600,N_2190);
or U4499 (N_4499,N_1870,N_2115);
xnor U4500 (N_4500,N_3184,N_3275);
or U4501 (N_4501,N_3539,N_4301);
and U4502 (N_4502,N_4459,N_3796);
nand U4503 (N_4503,N_3047,N_4270);
nand U4504 (N_4504,N_3654,N_4348);
or U4505 (N_4505,N_3686,N_3610);
nor U4506 (N_4506,N_3671,N_4223);
or U4507 (N_4507,N_4236,N_4052);
and U4508 (N_4508,N_4087,N_3802);
or U4509 (N_4509,N_3567,N_3831);
nand U4510 (N_4510,N_4033,N_3912);
nand U4511 (N_4511,N_4152,N_4228);
nor U4512 (N_4512,N_3987,N_4094);
and U4513 (N_4513,N_3724,N_3417);
and U4514 (N_4514,N_4031,N_3112);
and U4515 (N_4515,N_3027,N_3624);
xnor U4516 (N_4516,N_3630,N_3670);
xor U4517 (N_4517,N_3335,N_3969);
or U4518 (N_4518,N_4313,N_3012);
or U4519 (N_4519,N_3921,N_4201);
or U4520 (N_4520,N_3465,N_3240);
xnor U4521 (N_4521,N_3328,N_3255);
or U4522 (N_4522,N_4012,N_3496);
nor U4523 (N_4523,N_4063,N_3820);
xor U4524 (N_4524,N_3367,N_3786);
or U4525 (N_4525,N_3464,N_3138);
xnor U4526 (N_4526,N_4465,N_3487);
and U4527 (N_4527,N_3731,N_4409);
nor U4528 (N_4528,N_3763,N_4159);
xnor U4529 (N_4529,N_3396,N_3205);
or U4530 (N_4530,N_3893,N_4478);
and U4531 (N_4531,N_3570,N_3156);
nor U4532 (N_4532,N_4410,N_3973);
and U4533 (N_4533,N_3833,N_3766);
nor U4534 (N_4534,N_4456,N_4375);
nor U4535 (N_4535,N_4073,N_4104);
nor U4536 (N_4536,N_3208,N_4383);
xnor U4537 (N_4537,N_4119,N_3433);
or U4538 (N_4538,N_3025,N_3767);
or U4539 (N_4539,N_4428,N_4083);
xnor U4540 (N_4540,N_4058,N_4071);
or U4541 (N_4541,N_4432,N_3867);
and U4542 (N_4542,N_3728,N_4371);
and U4543 (N_4543,N_3805,N_4394);
or U4544 (N_4544,N_3952,N_4424);
xnor U4545 (N_4545,N_3814,N_3979);
or U4546 (N_4546,N_3383,N_4075);
nor U4547 (N_4547,N_3596,N_3504);
nand U4548 (N_4548,N_4145,N_3946);
nor U4549 (N_4549,N_4006,N_3750);
and U4550 (N_4550,N_3536,N_3482);
xnor U4551 (N_4551,N_3378,N_3297);
nand U4552 (N_4552,N_4492,N_3589);
nor U4553 (N_4553,N_4361,N_4476);
or U4554 (N_4554,N_3155,N_3273);
and U4555 (N_4555,N_3350,N_3173);
xor U4556 (N_4556,N_3058,N_4008);
and U4557 (N_4557,N_4067,N_3498);
and U4558 (N_4558,N_3687,N_3294);
or U4559 (N_4559,N_4368,N_3712);
xor U4560 (N_4560,N_3250,N_3582);
nand U4561 (N_4561,N_4376,N_3352);
nor U4562 (N_4562,N_3719,N_4105);
nor U4563 (N_4563,N_3140,N_4421);
nand U4564 (N_4564,N_3020,N_3197);
and U4565 (N_4565,N_3795,N_4319);
and U4566 (N_4566,N_4032,N_3700);
and U4567 (N_4567,N_4382,N_4156);
nand U4568 (N_4568,N_3109,N_3660);
nor U4569 (N_4569,N_3698,N_3067);
nor U4570 (N_4570,N_3530,N_3999);
xor U4571 (N_4571,N_4374,N_3743);
and U4572 (N_4572,N_3800,N_4059);
or U4573 (N_4573,N_3607,N_3543);
and U4574 (N_4574,N_4487,N_3819);
or U4575 (N_4575,N_4475,N_4252);
nand U4576 (N_4576,N_4442,N_3931);
nor U4577 (N_4577,N_3132,N_3391);
nor U4578 (N_4578,N_4339,N_3550);
and U4579 (N_4579,N_3571,N_3829);
nand U4580 (N_4580,N_3420,N_3333);
nor U4581 (N_4581,N_4282,N_3705);
nand U4582 (N_4582,N_3723,N_4286);
nand U4583 (N_4583,N_4360,N_3316);
and U4584 (N_4584,N_3545,N_3072);
nor U4585 (N_4585,N_3726,N_3429);
nor U4586 (N_4586,N_4149,N_4296);
or U4587 (N_4587,N_4316,N_4412);
nand U4588 (N_4588,N_4262,N_4081);
or U4589 (N_4589,N_4212,N_3972);
and U4590 (N_4590,N_4235,N_3659);
nor U4591 (N_4591,N_3157,N_4054);
nand U4592 (N_4592,N_3692,N_4472);
nor U4593 (N_4593,N_4308,N_3890);
and U4594 (N_4594,N_4100,N_4060);
xor U4595 (N_4595,N_3699,N_3754);
nand U4596 (N_4596,N_3597,N_3643);
xor U4597 (N_4597,N_3110,N_3234);
or U4598 (N_4598,N_3438,N_4147);
or U4599 (N_4599,N_3503,N_3292);
xnor U4600 (N_4600,N_3770,N_4381);
xor U4601 (N_4601,N_3259,N_4309);
xor U4602 (N_4602,N_3392,N_3886);
and U4603 (N_4603,N_3863,N_3963);
xnor U4604 (N_4604,N_4333,N_3206);
nor U4605 (N_4605,N_4474,N_3095);
xor U4606 (N_4606,N_3682,N_4085);
or U4607 (N_4607,N_3116,N_4039);
xnor U4608 (N_4608,N_3303,N_3314);
or U4609 (N_4609,N_3559,N_4258);
or U4610 (N_4610,N_3439,N_3163);
and U4611 (N_4611,N_3454,N_3213);
nand U4612 (N_4612,N_3377,N_3771);
nor U4613 (N_4613,N_3204,N_4129);
and U4614 (N_4614,N_3787,N_4022);
or U4615 (N_4615,N_3450,N_4118);
nor U4616 (N_4616,N_3148,N_3744);
xnor U4617 (N_4617,N_4070,N_3913);
nand U4618 (N_4618,N_3821,N_4407);
and U4619 (N_4619,N_3343,N_3996);
nand U4620 (N_4620,N_3798,N_3203);
or U4621 (N_4621,N_3887,N_3480);
nor U4622 (N_4622,N_3431,N_3909);
or U4623 (N_4623,N_4469,N_3511);
and U4624 (N_4624,N_3007,N_3287);
or U4625 (N_4625,N_3778,N_4198);
xnor U4626 (N_4626,N_4323,N_4109);
and U4627 (N_4627,N_3388,N_3428);
and U4628 (N_4628,N_3371,N_3956);
xor U4629 (N_4629,N_3120,N_3579);
or U4630 (N_4630,N_4254,N_4398);
nor U4631 (N_4631,N_3422,N_3218);
xnor U4632 (N_4632,N_3971,N_4385);
xor U4633 (N_4633,N_3151,N_3855);
nor U4634 (N_4634,N_4193,N_4345);
nor U4635 (N_4635,N_4351,N_3907);
or U4636 (N_4636,N_3677,N_3456);
and U4637 (N_4637,N_3419,N_3604);
or U4638 (N_4638,N_4227,N_3021);
nand U4639 (N_4639,N_3953,N_3525);
nand U4640 (N_4640,N_3935,N_3612);
nand U4641 (N_4641,N_3175,N_3172);
xor U4642 (N_4642,N_4233,N_4391);
and U4643 (N_4643,N_3179,N_4215);
nor U4644 (N_4644,N_3748,N_3244);
nor U4645 (N_4645,N_3812,N_3074);
or U4646 (N_4646,N_3801,N_3930);
and U4647 (N_4647,N_3181,N_3858);
nor U4648 (N_4648,N_4176,N_3683);
nand U4649 (N_4649,N_4422,N_3541);
xnor U4650 (N_4650,N_3409,N_4166);
or U4651 (N_4651,N_3411,N_3590);
nor U4652 (N_4652,N_3370,N_4415);
nor U4653 (N_4653,N_3390,N_3103);
nand U4654 (N_4654,N_3653,N_3257);
or U4655 (N_4655,N_3331,N_4413);
xnor U4656 (N_4656,N_4234,N_4148);
nor U4657 (N_4657,N_3752,N_3057);
nand U4658 (N_4658,N_4402,N_3762);
and U4659 (N_4659,N_4435,N_4139);
or U4660 (N_4660,N_4030,N_4390);
xor U4661 (N_4661,N_3540,N_3611);
and U4662 (N_4662,N_3978,N_4480);
xnor U4663 (N_4663,N_4414,N_3060);
or U4664 (N_4664,N_4199,N_4138);
nor U4665 (N_4665,N_3413,N_3399);
and U4666 (N_4666,N_3625,N_4396);
nand U4667 (N_4667,N_3566,N_4047);
nand U4668 (N_4668,N_3920,N_4246);
xnor U4669 (N_4669,N_3828,N_3130);
nor U4670 (N_4670,N_4276,N_4483);
and U4671 (N_4671,N_4167,N_3527);
and U4672 (N_4672,N_3967,N_3284);
nand U4673 (N_4673,N_3874,N_3158);
nand U4674 (N_4674,N_4259,N_4009);
xor U4675 (N_4675,N_3005,N_3400);
nand U4676 (N_4676,N_3210,N_3934);
nor U4677 (N_4677,N_3453,N_3282);
or U4678 (N_4678,N_3732,N_3782);
nand U4679 (N_4679,N_3188,N_3080);
xor U4680 (N_4680,N_3279,N_3299);
nand U4681 (N_4681,N_3729,N_4099);
or U4682 (N_4682,N_4453,N_3246);
nor U4683 (N_4683,N_3477,N_3542);
xor U4684 (N_4684,N_4317,N_4134);
or U4685 (N_4685,N_4369,N_3494);
and U4686 (N_4686,N_3165,N_3461);
nand U4687 (N_4687,N_3779,N_3772);
xnor U4688 (N_4688,N_3514,N_3278);
nand U4689 (N_4689,N_4489,N_4338);
and U4690 (N_4690,N_4384,N_4464);
nand U4691 (N_4691,N_3789,N_3848);
and U4692 (N_4692,N_4454,N_3323);
nor U4693 (N_4693,N_3850,N_4165);
xnor U4694 (N_4694,N_3622,N_3270);
or U4695 (N_4695,N_3024,N_3212);
nor U4696 (N_4696,N_3746,N_3510);
xnor U4697 (N_4697,N_3895,N_4436);
nor U4698 (N_4698,N_4380,N_3271);
and U4699 (N_4699,N_3359,N_3076);
and U4700 (N_4700,N_3416,N_3311);
xnor U4701 (N_4701,N_3619,N_4352);
and U4702 (N_4702,N_3827,N_4204);
nor U4703 (N_4703,N_3055,N_3455);
and U4704 (N_4704,N_4173,N_3864);
and U4705 (N_4705,N_3577,N_3406);
nor U4706 (N_4706,N_3680,N_3003);
nand U4707 (N_4707,N_4493,N_4297);
nand U4708 (N_4708,N_3938,N_4216);
xnor U4709 (N_4709,N_3618,N_3531);
and U4710 (N_4710,N_3127,N_3118);
and U4711 (N_4711,N_3555,N_4448);
and U4712 (N_4712,N_4355,N_3783);
xnor U4713 (N_4713,N_3927,N_3190);
nand U4714 (N_4714,N_4091,N_3853);
and U4715 (N_4715,N_3737,N_3169);
or U4716 (N_4716,N_4076,N_3932);
xor U4717 (N_4717,N_4238,N_3241);
nor U4718 (N_4718,N_4046,N_3681);
xor U4719 (N_4719,N_3500,N_4359);
nand U4720 (N_4720,N_3449,N_3166);
and U4721 (N_4721,N_3004,N_4268);
nor U4722 (N_4722,N_3117,N_4265);
nand U4723 (N_4723,N_3811,N_4066);
xor U4724 (N_4724,N_3337,N_4036);
or U4725 (N_4725,N_3568,N_4337);
nand U4726 (N_4726,N_3048,N_4177);
xor U4727 (N_4727,N_4210,N_3088);
nor U4728 (N_4728,N_4473,N_4458);
nor U4729 (N_4729,N_3185,N_3149);
and U4730 (N_4730,N_4219,N_3096);
xnor U4731 (N_4731,N_3049,N_4019);
and U4732 (N_4732,N_3839,N_4499);
xor U4733 (N_4733,N_3039,N_3101);
nor U4734 (N_4734,N_4090,N_3070);
nand U4735 (N_4735,N_3685,N_3532);
xor U4736 (N_4736,N_3896,N_3189);
xor U4737 (N_4737,N_4000,N_3492);
and U4738 (N_4738,N_3115,N_3790);
or U4739 (N_4739,N_4184,N_3276);
nand U4740 (N_4740,N_4328,N_4164);
or U4741 (N_4741,N_3954,N_4379);
nand U4742 (N_4742,N_4445,N_3629);
and U4743 (N_4743,N_4275,N_3672);
and U4744 (N_4744,N_3903,N_4055);
nor U4745 (N_4745,N_3083,N_3517);
or U4746 (N_4746,N_4170,N_3984);
xnor U4747 (N_4747,N_4029,N_3402);
xnor U4748 (N_4748,N_4449,N_3462);
nand U4749 (N_4749,N_4364,N_4327);
xor U4750 (N_4750,N_4441,N_4273);
nor U4751 (N_4751,N_4174,N_3209);
nand U4752 (N_4752,N_4482,N_3376);
nor U4753 (N_4753,N_3145,N_3214);
nand U4754 (N_4754,N_3232,N_3332);
or U4755 (N_4755,N_4050,N_4124);
nor U4756 (N_4756,N_3836,N_3178);
and U4757 (N_4757,N_3037,N_3602);
nor U4758 (N_4758,N_3929,N_3837);
and U4759 (N_4759,N_3283,N_3452);
nand U4760 (N_4760,N_3147,N_3764);
nand U4761 (N_4761,N_3300,N_3298);
and U4762 (N_4762,N_3369,N_3735);
and U4763 (N_4763,N_3489,N_3817);
and U4764 (N_4764,N_3947,N_3872);
xor U4765 (N_4765,N_3475,N_4315);
nor U4766 (N_4766,N_3387,N_3198);
or U4767 (N_4767,N_3544,N_4336);
nor U4768 (N_4768,N_4195,N_3810);
nor U4769 (N_4769,N_3640,N_3583);
xnor U4770 (N_4770,N_3033,N_3964);
or U4771 (N_4771,N_3761,N_4292);
or U4772 (N_4772,N_3220,N_4111);
xor U4773 (N_4773,N_3014,N_4200);
or U4774 (N_4774,N_4408,N_3182);
nand U4775 (N_4775,N_3034,N_4146);
xor U4776 (N_4776,N_4365,N_3031);
or U4777 (N_4777,N_4477,N_3857);
nand U4778 (N_4778,N_3689,N_3881);
nand U4779 (N_4779,N_3106,N_3776);
nor U4780 (N_4780,N_4330,N_3026);
nor U4781 (N_4781,N_3704,N_3030);
or U4782 (N_4782,N_4217,N_3720);
nor U4783 (N_4783,N_3981,N_3702);
and U4784 (N_4784,N_4334,N_4358);
xnor U4785 (N_4785,N_3261,N_4284);
nor U4786 (N_4786,N_4205,N_3321);
nor U4787 (N_4787,N_3153,N_4023);
and U4788 (N_4788,N_4051,N_3094);
and U4789 (N_4789,N_3207,N_3628);
nor U4790 (N_4790,N_3635,N_4021);
nor U4791 (N_4791,N_4117,N_3623);
or U4792 (N_4792,N_3366,N_3840);
and U4793 (N_4793,N_4057,N_3144);
and U4794 (N_4794,N_3880,N_3111);
or U4795 (N_4795,N_4326,N_3301);
nor U4796 (N_4796,N_3585,N_3940);
and U4797 (N_4797,N_3223,N_3888);
xnor U4798 (N_4798,N_3372,N_3141);
and U4799 (N_4799,N_4405,N_3788);
and U4800 (N_4800,N_4303,N_3708);
nand U4801 (N_4801,N_4224,N_3838);
nor U4802 (N_4802,N_4411,N_4321);
nor U4803 (N_4803,N_3760,N_3528);
xnor U4804 (N_4804,N_3028,N_3363);
nand U4805 (N_4805,N_3632,N_3807);
nand U4806 (N_4806,N_4191,N_3050);
nor U4807 (N_4807,N_3576,N_4079);
xnor U4808 (N_4808,N_4494,N_3382);
nor U4809 (N_4809,N_3286,N_3329);
xor U4810 (N_4810,N_3526,N_3092);
nor U4811 (N_4811,N_4242,N_3041);
or U4812 (N_4812,N_3081,N_3499);
nor U4813 (N_4813,N_4372,N_4426);
xnor U4814 (N_4814,N_4261,N_4125);
and U4815 (N_4815,N_4271,N_3040);
or U4816 (N_4816,N_4264,N_3822);
nor U4817 (N_4817,N_4347,N_3272);
and U4818 (N_4818,N_3557,N_4169);
xnor U4819 (N_4819,N_3397,N_3443);
nand U4820 (N_4820,N_4007,N_4013);
nand U4821 (N_4821,N_3408,N_4089);
nor U4822 (N_4822,N_3649,N_3187);
or U4823 (N_4823,N_3038,N_3884);
nand U4824 (N_4824,N_4386,N_4190);
nor U4825 (N_4825,N_4225,N_3970);
or U4826 (N_4826,N_3753,N_3345);
or U4827 (N_4827,N_4130,N_3052);
xnor U4828 (N_4828,N_4495,N_3315);
nor U4829 (N_4829,N_3725,N_4295);
xnor U4830 (N_4830,N_4042,N_4437);
and U4831 (N_4831,N_4197,N_4484);
and U4832 (N_4832,N_4263,N_3373);
or U4833 (N_4833,N_3520,N_4462);
nor U4834 (N_4834,N_4209,N_3260);
xnor U4835 (N_4835,N_3082,N_4053);
nor U4836 (N_4836,N_3230,N_3191);
nand U4837 (N_4837,N_4028,N_3957);
nor U4838 (N_4838,N_3871,N_3554);
and U4839 (N_4839,N_3922,N_3474);
xor U4840 (N_4840,N_3469,N_3936);
and U4841 (N_4841,N_3523,N_3615);
nor U4842 (N_4842,N_3642,N_3457);
nor U4843 (N_4843,N_3077,N_3824);
xnor U4844 (N_4844,N_3944,N_3695);
or U4845 (N_4845,N_3137,N_3663);
xor U4846 (N_4846,N_3951,N_4102);
nor U4847 (N_4847,N_3393,N_3305);
nand U4848 (N_4848,N_3253,N_3662);
xnor U4849 (N_4849,N_3852,N_4074);
nand U4850 (N_4850,N_4488,N_3134);
nand U4851 (N_4851,N_3780,N_4287);
nor U4852 (N_4852,N_4202,N_4274);
and U4853 (N_4853,N_3358,N_3718);
nand U4854 (N_4854,N_4269,N_3224);
xnor U4855 (N_4855,N_4377,N_4430);
and U4856 (N_4856,N_3269,N_3707);
xnor U4857 (N_4857,N_3084,N_3044);
xor U4858 (N_4858,N_3078,N_3458);
nand U4859 (N_4859,N_4324,N_3295);
nor U4860 (N_4860,N_3473,N_3606);
nor U4861 (N_4861,N_3104,N_3693);
nor U4862 (N_4862,N_3017,N_4243);
nand U4863 (N_4863,N_3879,N_4481);
and U4864 (N_4864,N_4003,N_3302);
nand U4865 (N_4865,N_4043,N_3832);
and U4866 (N_4866,N_4257,N_3497);
nor U4867 (N_4867,N_3274,N_3066);
xnor U4868 (N_4868,N_4266,N_3759);
or U4869 (N_4869,N_3883,N_3318);
nand U4870 (N_4870,N_3751,N_3524);
nand U4871 (N_4871,N_3124,N_3834);
nor U4872 (N_4872,N_4451,N_3404);
xnor U4873 (N_4873,N_3126,N_3785);
and U4874 (N_4874,N_3451,N_3757);
xor U4875 (N_4875,N_3340,N_3285);
or U4876 (N_4876,N_4196,N_4444);
and U4877 (N_4877,N_3123,N_3136);
xnor U4878 (N_4878,N_4239,N_3809);
or U4879 (N_4879,N_3937,N_3551);
or U4880 (N_4880,N_3355,N_3637);
nor U4881 (N_4881,N_4256,N_3564);
xor U4882 (N_4882,N_4367,N_4010);
nor U4883 (N_4883,N_4232,N_3009);
nor U4884 (N_4884,N_3774,N_4230);
nor U4885 (N_4885,N_3289,N_3657);
nand U4886 (N_4886,N_3434,N_4226);
nand U4887 (N_4887,N_3414,N_4439);
nand U4888 (N_4888,N_3010,N_4137);
and U4889 (N_4889,N_4357,N_3985);
and U4890 (N_4890,N_3773,N_3011);
or U4891 (N_4891,N_3418,N_3755);
nor U4892 (N_4892,N_3900,N_4127);
xor U4893 (N_4893,N_4392,N_4342);
nor U4894 (N_4894,N_3977,N_4331);
and U4895 (N_4895,N_3029,N_4106);
and U4896 (N_4896,N_4300,N_4373);
nor U4897 (N_4897,N_4214,N_3509);
and U4898 (N_4898,N_3694,N_3873);
nand U4899 (N_4899,N_4406,N_3068);
xnor U4900 (N_4900,N_3199,N_3484);
and U4901 (N_4901,N_3267,N_4440);
or U4902 (N_4902,N_4045,N_3865);
nand U4903 (N_4903,N_3733,N_4128);
nand U4904 (N_4904,N_3616,N_3717);
nor U4905 (N_4905,N_3098,N_3472);
and U4906 (N_4906,N_4179,N_4332);
xor U4907 (N_4907,N_4400,N_4175);
nor U4908 (N_4908,N_3845,N_3395);
nand U4909 (N_4909,N_3405,N_3375);
or U4910 (N_4910,N_3656,N_4329);
and U4911 (N_4911,N_3679,N_3226);
nand U4912 (N_4912,N_4311,N_3263);
and U4913 (N_4913,N_3097,N_4140);
xnor U4914 (N_4914,N_3231,N_3859);
xor U4915 (N_4915,N_3160,N_3575);
or U4916 (N_4916,N_3633,N_3219);
nor U4917 (N_4917,N_3334,N_3558);
and U4918 (N_4918,N_3018,N_4093);
xor U4919 (N_4919,N_4416,N_3064);
or U4920 (N_4920,N_3515,N_3955);
nor U4921 (N_4921,N_3129,N_4240);
or U4922 (N_4922,N_3741,N_4387);
nor U4923 (N_4923,N_3193,N_4291);
or U4924 (N_4924,N_3983,N_4095);
or U4925 (N_4925,N_3806,N_3892);
and U4926 (N_4926,N_4289,N_4491);
or U4927 (N_4927,N_3114,N_3982);
xnor U4928 (N_4928,N_3631,N_3221);
nor U4929 (N_4929,N_3991,N_4418);
xnor U4930 (N_4930,N_4136,N_3194);
xor U4931 (N_4931,N_3349,N_3646);
or U4932 (N_4932,N_3235,N_3825);
nor U4933 (N_4933,N_3006,N_3361);
or U4934 (N_4934,N_4035,N_3360);
xnor U4935 (N_4935,N_3412,N_4429);
or U4936 (N_4936,N_3522,N_3595);
xor U4937 (N_4937,N_3113,N_3146);
and U4938 (N_4938,N_3792,N_3180);
xor U4939 (N_4939,N_3425,N_4143);
nor U4940 (N_4940,N_3594,N_3684);
nand U4941 (N_4941,N_3364,N_3046);
nand U4942 (N_4942,N_4131,N_4363);
xor U4943 (N_4943,N_3093,N_3356);
xor U4944 (N_4944,N_3620,N_3799);
and U4945 (N_4945,N_3256,N_3065);
xnor U4946 (N_4946,N_3164,N_3714);
nand U4947 (N_4947,N_3877,N_3674);
xnor U4948 (N_4948,N_3901,N_3239);
or U4949 (N_4949,N_3304,N_3357);
xnor U4950 (N_4950,N_4158,N_3354);
xor U4951 (N_4951,N_3990,N_3466);
nor U4952 (N_4952,N_4061,N_3994);
or U4953 (N_4953,N_3745,N_3756);
nor U4954 (N_4954,N_4103,N_4120);
nor U4955 (N_4955,N_4142,N_3013);
xor U4956 (N_4956,N_4157,N_3324);
nor U4957 (N_4957,N_3252,N_4279);
nand U4958 (N_4958,N_3061,N_3085);
nor U4959 (N_4959,N_4293,N_4027);
and U4960 (N_4960,N_3775,N_4314);
and U4961 (N_4961,N_4404,N_4126);
and U4962 (N_4962,N_4171,N_4248);
nor U4963 (N_4963,N_3995,N_4306);
xnor U4964 (N_4964,N_3605,N_3430);
nor U4965 (N_4965,N_3059,N_4155);
xor U4966 (N_4966,N_3980,N_3535);
nor U4967 (N_4967,N_4307,N_3918);
nor U4968 (N_4968,N_3507,N_3960);
xor U4969 (N_4969,N_4221,N_3808);
nand U4970 (N_4970,N_3993,N_3661);
xnor U4971 (N_4971,N_3997,N_3587);
and U4972 (N_4972,N_3665,N_3841);
and U4973 (N_4973,N_4302,N_4471);
and U4974 (N_4974,N_3308,N_3572);
nand U4975 (N_4975,N_4457,N_4450);
and U4976 (N_4976,N_3537,N_4281);
or U4977 (N_4977,N_4389,N_3368);
or U4978 (N_4978,N_4343,N_3854);
nand U4979 (N_4979,N_3490,N_3974);
or U4980 (N_4980,N_3293,N_4037);
and U4981 (N_4981,N_3481,N_4267);
or U4982 (N_4982,N_3254,N_3362);
or U4983 (N_4983,N_3423,N_3251);
or U4984 (N_4984,N_4080,N_3910);
and U4985 (N_4985,N_3945,N_3794);
nand U4986 (N_4986,N_3709,N_3229);
xor U4987 (N_4987,N_3502,N_4260);
nor U4988 (N_4988,N_4399,N_3432);
and U4989 (N_4989,N_3015,N_3100);
or U4990 (N_4990,N_4419,N_3992);
nor U4991 (N_4991,N_3885,N_3784);
and U4992 (N_4992,N_3053,N_3245);
nor U4993 (N_4993,N_3573,N_4108);
or U4994 (N_4994,N_3398,N_3296);
nor U4995 (N_4995,N_4431,N_4305);
nor U4996 (N_4996,N_4020,N_3548);
nor U4997 (N_4997,N_4101,N_3948);
nor U4998 (N_4998,N_4132,N_3675);
or U4999 (N_4999,N_3483,N_4041);
or U5000 (N_5000,N_3152,N_4247);
nor U5001 (N_5001,N_3508,N_3281);
nand U5002 (N_5002,N_3247,N_3634);
nor U5003 (N_5003,N_4272,N_3898);
xor U5004 (N_5004,N_3569,N_3942);
or U5005 (N_5005,N_3804,N_4133);
nor U5006 (N_5006,N_3108,N_4335);
nand U5007 (N_5007,N_3478,N_3581);
nor U5008 (N_5008,N_3338,N_3176);
nand U5009 (N_5009,N_3512,N_3168);
nor U5010 (N_5010,N_4461,N_4341);
xor U5011 (N_5011,N_4350,N_3348);
nand U5012 (N_5012,N_3008,N_4486);
xor U5013 (N_5013,N_3336,N_3739);
xnor U5014 (N_5014,N_3317,N_3962);
or U5015 (N_5015,N_3379,N_3501);
nand U5016 (N_5016,N_3636,N_4397);
xnor U5017 (N_5017,N_3721,N_3621);
or U5018 (N_5018,N_4084,N_3866);
or U5019 (N_5019,N_3552,N_3847);
and U5020 (N_5020,N_4092,N_3002);
or U5021 (N_5021,N_4062,N_3959);
nand U5022 (N_5022,N_3310,N_3915);
xor U5023 (N_5023,N_3035,N_4098);
and U5024 (N_5024,N_3715,N_3706);
or U5025 (N_5025,N_4192,N_4077);
and U5026 (N_5026,N_3747,N_3016);
and U5027 (N_5027,N_3869,N_3609);
or U5028 (N_5028,N_3561,N_3351);
nor U5029 (N_5029,N_4016,N_3186);
and U5030 (N_5030,N_4245,N_4356);
xor U5031 (N_5031,N_3818,N_3891);
or U5032 (N_5032,N_3902,N_3468);
xor U5033 (N_5033,N_4048,N_4163);
or U5034 (N_5034,N_3089,N_4255);
nand U5035 (N_5035,N_3380,N_3105);
and U5036 (N_5036,N_3534,N_3765);
nor U5037 (N_5037,N_4014,N_4049);
nand U5038 (N_5038,N_3381,N_4011);
nor U5039 (N_5039,N_3546,N_4185);
or U5040 (N_5040,N_3403,N_3830);
nor U5041 (N_5041,N_3326,N_4443);
or U5042 (N_5042,N_4299,N_3793);
and U5043 (N_5043,N_3436,N_3736);
nand U5044 (N_5044,N_3950,N_3236);
xnor U5045 (N_5045,N_3758,N_3174);
xnor U5046 (N_5046,N_4064,N_3521);
and U5047 (N_5047,N_3442,N_3086);
nand U5048 (N_5048,N_3407,N_3262);
nor U5049 (N_5049,N_3919,N_3876);
nand U5050 (N_5050,N_3075,N_4114);
and U5051 (N_5051,N_3740,N_3580);
nor U5052 (N_5052,N_4122,N_3645);
or U5053 (N_5053,N_4393,N_4304);
or U5054 (N_5054,N_4318,N_3238);
nor U5055 (N_5055,N_4467,N_4290);
nor U5056 (N_5056,N_3676,N_3102);
nor U5057 (N_5057,N_3131,N_3939);
xnor U5058 (N_5058,N_3467,N_4353);
and U5059 (N_5059,N_3926,N_3655);
or U5060 (N_5060,N_3603,N_3513);
xor U5061 (N_5061,N_3791,N_4161);
or U5062 (N_5062,N_3599,N_4496);
nand U5063 (N_5063,N_4107,N_3878);
nand U5064 (N_5064,N_4229,N_3069);
or U5065 (N_5065,N_3968,N_3965);
nor U5066 (N_5066,N_4320,N_3344);
or U5067 (N_5067,N_4460,N_3617);
xor U5068 (N_5068,N_4249,N_3091);
and U5069 (N_5069,N_4244,N_4188);
xor U5070 (N_5070,N_3384,N_4497);
nor U5071 (N_5071,N_4490,N_3325);
nand U5072 (N_5072,N_3823,N_3374);
nor U5073 (N_5073,N_3815,N_4349);
nor U5074 (N_5074,N_4470,N_3925);
and U5075 (N_5075,N_3079,N_4237);
nor U5076 (N_5076,N_3036,N_3668);
xnor U5077 (N_5077,N_3651,N_3386);
or U5078 (N_5078,N_4001,N_3738);
nor U5079 (N_5079,N_3444,N_4040);
and U5080 (N_5080,N_3322,N_3128);
nor U5081 (N_5081,N_3908,N_4088);
nand U5082 (N_5082,N_3280,N_3192);
nand U5083 (N_5083,N_3437,N_3201);
nor U5084 (N_5084,N_3183,N_3211);
xnor U5085 (N_5085,N_3249,N_3073);
and U5086 (N_5086,N_4154,N_4121);
xor U5087 (N_5087,N_3584,N_4213);
nor U5088 (N_5088,N_3243,N_3549);
xor U5089 (N_5089,N_4446,N_4231);
or U5090 (N_5090,N_3588,N_3917);
or U5091 (N_5091,N_4082,N_3734);
nor U5092 (N_5092,N_4211,N_4346);
xnor U5093 (N_5093,N_3330,N_3479);
nand U5094 (N_5094,N_4024,N_4141);
xor U5095 (N_5095,N_4251,N_3862);
or U5096 (N_5096,N_4025,N_3288);
or U5097 (N_5097,N_3200,N_3894);
or U5098 (N_5098,N_3486,N_3150);
or U5099 (N_5099,N_3673,N_3056);
nand U5100 (N_5100,N_3440,N_3904);
xor U5101 (N_5101,N_4065,N_3664);
nand U5102 (N_5102,N_3488,N_3309);
and U5103 (N_5103,N_4403,N_3849);
nand U5104 (N_5104,N_3519,N_3162);
nand U5105 (N_5105,N_4044,N_4485);
nand U5106 (N_5106,N_4002,N_3342);
or U5107 (N_5107,N_3424,N_3578);
or U5108 (N_5108,N_4112,N_4378);
or U5109 (N_5109,N_3600,N_4447);
or U5110 (N_5110,N_3691,N_4423);
nor U5111 (N_5111,N_3320,N_4115);
nor U5112 (N_5112,N_3813,N_3562);
nor U5113 (N_5113,N_3266,N_4144);
nor U5114 (N_5114,N_3518,N_3923);
xnor U5115 (N_5115,N_3051,N_3045);
or U5116 (N_5116,N_3032,N_3797);
or U5117 (N_5117,N_4250,N_4135);
nor U5118 (N_5118,N_3638,N_4096);
nand U5119 (N_5119,N_4253,N_3319);
nand U5120 (N_5120,N_3727,N_3062);
xor U5121 (N_5121,N_3856,N_3716);
nor U5122 (N_5122,N_3882,N_3769);
xor U5123 (N_5123,N_4160,N_4479);
nand U5124 (N_5124,N_3217,N_3626);
nor U5125 (N_5125,N_3000,N_3491);
nor U5126 (N_5126,N_3989,N_3421);
or U5127 (N_5127,N_3843,N_3516);
or U5128 (N_5128,N_4388,N_3242);
and U5129 (N_5129,N_3592,N_4178);
nor U5130 (N_5130,N_3690,N_3389);
and U5131 (N_5131,N_3170,N_3547);
xor U5132 (N_5132,N_3697,N_3107);
nand U5133 (N_5133,N_3928,N_3023);
or U5134 (N_5134,N_3264,N_3327);
and U5135 (N_5135,N_4312,N_3063);
nor U5136 (N_5136,N_4433,N_3860);
or U5137 (N_5137,N_3353,N_3961);
nand U5138 (N_5138,N_3851,N_3042);
and U5139 (N_5139,N_4370,N_3870);
nor U5140 (N_5140,N_4434,N_4463);
nor U5141 (N_5141,N_4116,N_3291);
xor U5142 (N_5142,N_4026,N_3171);
nand U5143 (N_5143,N_3133,N_3385);
nand U5144 (N_5144,N_3506,N_3658);
xor U5145 (N_5145,N_3538,N_4034);
or U5146 (N_5146,N_4086,N_3598);
nand U5147 (N_5147,N_4452,N_3401);
nor U5148 (N_5148,N_3485,N_4194);
nand U5149 (N_5149,N_4207,N_3447);
nor U5150 (N_5150,N_3943,N_3143);
nand U5151 (N_5151,N_3196,N_3043);
or U5152 (N_5152,N_3905,N_4283);
nand U5153 (N_5153,N_4005,N_3307);
or U5154 (N_5154,N_3446,N_4017);
and U5155 (N_5155,N_3933,N_3730);
nand U5156 (N_5156,N_4153,N_4222);
nor U5157 (N_5157,N_4123,N_3139);
xnor U5158 (N_5158,N_3493,N_4466);
nand U5159 (N_5159,N_4172,N_3875);
nand U5160 (N_5160,N_3435,N_3711);
nand U5161 (N_5161,N_3914,N_3441);
or U5162 (N_5162,N_3722,N_3842);
and U5163 (N_5163,N_3975,N_4354);
or U5164 (N_5164,N_4180,N_3119);
nand U5165 (N_5165,N_3614,N_3001);
xor U5166 (N_5166,N_3265,N_3533);
or U5167 (N_5167,N_3608,N_4018);
xor U5168 (N_5168,N_3346,N_3290);
and U5169 (N_5169,N_4110,N_3868);
and U5170 (N_5170,N_4417,N_4278);
and U5171 (N_5171,N_3966,N_4206);
and U5172 (N_5172,N_3470,N_3341);
nand U5173 (N_5173,N_3574,N_3650);
nand U5174 (N_5174,N_3816,N_3019);
nand U5175 (N_5175,N_4427,N_3142);
or U5176 (N_5176,N_3861,N_3347);
or U5177 (N_5177,N_3495,N_3459);
nand U5178 (N_5178,N_3090,N_4069);
or U5179 (N_5179,N_4183,N_3415);
and U5180 (N_5180,N_4162,N_4186);
or U5181 (N_5181,N_3121,N_4277);
nand U5182 (N_5182,N_3460,N_3505);
and U5183 (N_5183,N_3696,N_3826);
or U5184 (N_5184,N_3087,N_3613);
nor U5185 (N_5185,N_3906,N_3777);
nand U5186 (N_5186,N_3529,N_4072);
nand U5187 (N_5187,N_4366,N_4189);
nand U5188 (N_5188,N_3445,N_4298);
nor U5189 (N_5189,N_3202,N_4113);
nor U5190 (N_5190,N_3916,N_4097);
or U5191 (N_5191,N_4078,N_4280);
nand U5192 (N_5192,N_3553,N_3678);
nand U5193 (N_5193,N_3277,N_3394);
xnor U5194 (N_5194,N_4150,N_3749);
nand U5195 (N_5195,N_3135,N_4038);
xor U5196 (N_5196,N_4322,N_4220);
nor U5197 (N_5197,N_3591,N_3846);
nor U5198 (N_5198,N_3195,N_4498);
xnor U5199 (N_5199,N_3648,N_3216);
nor U5200 (N_5200,N_4340,N_3988);
nor U5201 (N_5201,N_3365,N_3713);
nand U5202 (N_5202,N_3768,N_3237);
nor U5203 (N_5203,N_3803,N_4068);
xor U5204 (N_5204,N_3958,N_3781);
xnor U5205 (N_5205,N_3122,N_3099);
nor U5206 (N_5206,N_4151,N_3161);
or U5207 (N_5207,N_3647,N_3844);
xnor U5208 (N_5208,N_3601,N_3426);
nand U5209 (N_5209,N_3227,N_4004);
xnor U5210 (N_5210,N_4182,N_3125);
nand U5211 (N_5211,N_4455,N_4288);
xnor U5212 (N_5212,N_3560,N_3054);
xor U5213 (N_5213,N_3897,N_4468);
and U5214 (N_5214,N_4181,N_3742);
and U5215 (N_5215,N_4015,N_3911);
and U5216 (N_5216,N_3652,N_3701);
and U5217 (N_5217,N_3565,N_3228);
nand U5218 (N_5218,N_3644,N_3949);
or U5219 (N_5219,N_3639,N_4218);
or U5220 (N_5220,N_3312,N_3159);
nor U5221 (N_5221,N_4056,N_3899);
xor U5222 (N_5222,N_3258,N_3248);
xnor U5223 (N_5223,N_3710,N_3022);
nor U5224 (N_5224,N_3339,N_4401);
and U5225 (N_5225,N_4168,N_3666);
or U5226 (N_5226,N_3222,N_3586);
xor U5227 (N_5227,N_3463,N_3986);
and U5228 (N_5228,N_3313,N_4285);
nand U5229 (N_5229,N_4362,N_3448);
nand U5230 (N_5230,N_3215,N_3593);
xnor U5231 (N_5231,N_4325,N_3177);
or U5232 (N_5232,N_3306,N_3071);
nand U5233 (N_5233,N_3268,N_3225);
nor U5234 (N_5234,N_4310,N_3410);
xnor U5235 (N_5235,N_4420,N_3471);
nand U5236 (N_5236,N_4187,N_3627);
nand U5237 (N_5237,N_3167,N_3703);
nand U5238 (N_5238,N_3476,N_3688);
nand U5239 (N_5239,N_4395,N_4203);
nand U5240 (N_5240,N_3154,N_3233);
and U5241 (N_5241,N_3669,N_3889);
nor U5242 (N_5242,N_4208,N_4241);
xor U5243 (N_5243,N_3998,N_3556);
or U5244 (N_5244,N_3667,N_3835);
xnor U5245 (N_5245,N_4438,N_3427);
or U5246 (N_5246,N_4294,N_3641);
xnor U5247 (N_5247,N_3924,N_3941);
or U5248 (N_5248,N_4425,N_4344);
and U5249 (N_5249,N_3563,N_3976);
xnor U5250 (N_5250,N_3732,N_3470);
nand U5251 (N_5251,N_3726,N_4126);
and U5252 (N_5252,N_4356,N_4003);
nor U5253 (N_5253,N_3351,N_3352);
and U5254 (N_5254,N_4012,N_3284);
or U5255 (N_5255,N_3896,N_3776);
xor U5256 (N_5256,N_3663,N_3604);
nand U5257 (N_5257,N_4218,N_3282);
xor U5258 (N_5258,N_4063,N_3065);
or U5259 (N_5259,N_4475,N_3202);
and U5260 (N_5260,N_3966,N_4132);
and U5261 (N_5261,N_3873,N_3129);
or U5262 (N_5262,N_3515,N_3335);
or U5263 (N_5263,N_3921,N_3942);
nand U5264 (N_5264,N_3366,N_4440);
nand U5265 (N_5265,N_3164,N_3812);
nor U5266 (N_5266,N_3570,N_3906);
xnor U5267 (N_5267,N_3078,N_3531);
xnor U5268 (N_5268,N_4108,N_3955);
or U5269 (N_5269,N_4377,N_3098);
nand U5270 (N_5270,N_4074,N_3686);
and U5271 (N_5271,N_3510,N_3819);
nor U5272 (N_5272,N_3658,N_4003);
xnor U5273 (N_5273,N_3551,N_4387);
xnor U5274 (N_5274,N_3408,N_4025);
nor U5275 (N_5275,N_4373,N_3455);
nor U5276 (N_5276,N_3702,N_3828);
nor U5277 (N_5277,N_4338,N_3898);
nor U5278 (N_5278,N_3432,N_3827);
xor U5279 (N_5279,N_3386,N_4332);
xnor U5280 (N_5280,N_4406,N_4284);
nor U5281 (N_5281,N_4120,N_3883);
and U5282 (N_5282,N_4029,N_4371);
xnor U5283 (N_5283,N_3323,N_3633);
xor U5284 (N_5284,N_4412,N_3899);
xor U5285 (N_5285,N_3444,N_4157);
nor U5286 (N_5286,N_3921,N_4308);
nand U5287 (N_5287,N_4455,N_4210);
nand U5288 (N_5288,N_3026,N_4423);
nor U5289 (N_5289,N_4012,N_4431);
nor U5290 (N_5290,N_3083,N_3178);
xor U5291 (N_5291,N_3932,N_3490);
xor U5292 (N_5292,N_3561,N_3596);
xnor U5293 (N_5293,N_3603,N_3236);
nor U5294 (N_5294,N_4054,N_3746);
nand U5295 (N_5295,N_3969,N_4409);
nand U5296 (N_5296,N_4416,N_3749);
nand U5297 (N_5297,N_4381,N_4383);
nand U5298 (N_5298,N_3961,N_3903);
nand U5299 (N_5299,N_3661,N_3049);
nor U5300 (N_5300,N_4235,N_4209);
xnor U5301 (N_5301,N_3131,N_3246);
xor U5302 (N_5302,N_3674,N_3929);
nand U5303 (N_5303,N_3812,N_4177);
and U5304 (N_5304,N_3262,N_4363);
or U5305 (N_5305,N_3216,N_3241);
nand U5306 (N_5306,N_4253,N_3540);
and U5307 (N_5307,N_4147,N_3930);
or U5308 (N_5308,N_3619,N_4087);
or U5309 (N_5309,N_3350,N_3106);
xor U5310 (N_5310,N_3181,N_3104);
and U5311 (N_5311,N_3512,N_3560);
nand U5312 (N_5312,N_4407,N_4410);
or U5313 (N_5313,N_3716,N_3761);
and U5314 (N_5314,N_4366,N_3662);
nand U5315 (N_5315,N_3421,N_3191);
xor U5316 (N_5316,N_3087,N_3242);
xnor U5317 (N_5317,N_3040,N_3886);
nor U5318 (N_5318,N_3819,N_4204);
xor U5319 (N_5319,N_3245,N_3232);
or U5320 (N_5320,N_3753,N_4334);
nor U5321 (N_5321,N_3193,N_3170);
nor U5322 (N_5322,N_3059,N_3979);
xnor U5323 (N_5323,N_4213,N_4234);
or U5324 (N_5324,N_4301,N_4292);
or U5325 (N_5325,N_3342,N_3529);
and U5326 (N_5326,N_4234,N_3267);
or U5327 (N_5327,N_3326,N_3241);
xnor U5328 (N_5328,N_3286,N_3112);
and U5329 (N_5329,N_3192,N_3625);
or U5330 (N_5330,N_3318,N_3354);
nor U5331 (N_5331,N_4290,N_3914);
and U5332 (N_5332,N_3228,N_3722);
nor U5333 (N_5333,N_3150,N_3124);
and U5334 (N_5334,N_3661,N_3110);
xor U5335 (N_5335,N_3322,N_3875);
nand U5336 (N_5336,N_4017,N_3465);
and U5337 (N_5337,N_3445,N_4367);
xnor U5338 (N_5338,N_4277,N_3694);
or U5339 (N_5339,N_3230,N_4251);
nor U5340 (N_5340,N_3138,N_4333);
or U5341 (N_5341,N_3205,N_3186);
xnor U5342 (N_5342,N_3519,N_3632);
and U5343 (N_5343,N_3125,N_4395);
and U5344 (N_5344,N_3678,N_3641);
and U5345 (N_5345,N_4174,N_4378);
xnor U5346 (N_5346,N_3896,N_3528);
nand U5347 (N_5347,N_3638,N_3600);
nand U5348 (N_5348,N_3428,N_3187);
and U5349 (N_5349,N_3661,N_3480);
nand U5350 (N_5350,N_4134,N_4149);
and U5351 (N_5351,N_3487,N_3543);
xor U5352 (N_5352,N_3913,N_3910);
xor U5353 (N_5353,N_3849,N_3967);
or U5354 (N_5354,N_4317,N_3645);
nand U5355 (N_5355,N_4492,N_4040);
and U5356 (N_5356,N_3038,N_3550);
or U5357 (N_5357,N_4342,N_3995);
and U5358 (N_5358,N_4224,N_3749);
xnor U5359 (N_5359,N_3183,N_3056);
nand U5360 (N_5360,N_3348,N_3795);
xor U5361 (N_5361,N_3816,N_3538);
xor U5362 (N_5362,N_3993,N_4183);
nor U5363 (N_5363,N_3938,N_3320);
and U5364 (N_5364,N_3017,N_3377);
nand U5365 (N_5365,N_4372,N_3995);
nand U5366 (N_5366,N_3581,N_3469);
and U5367 (N_5367,N_3077,N_3931);
nor U5368 (N_5368,N_4162,N_3591);
xnor U5369 (N_5369,N_3924,N_4431);
xnor U5370 (N_5370,N_3996,N_3966);
nor U5371 (N_5371,N_4284,N_4064);
xor U5372 (N_5372,N_3245,N_4489);
xnor U5373 (N_5373,N_4284,N_4466);
or U5374 (N_5374,N_4200,N_3887);
or U5375 (N_5375,N_3498,N_4401);
nand U5376 (N_5376,N_4077,N_4239);
xor U5377 (N_5377,N_3904,N_3381);
or U5378 (N_5378,N_3921,N_4027);
xnor U5379 (N_5379,N_4121,N_4493);
or U5380 (N_5380,N_4075,N_3634);
nor U5381 (N_5381,N_3120,N_3819);
nor U5382 (N_5382,N_4035,N_3291);
and U5383 (N_5383,N_3764,N_3679);
xor U5384 (N_5384,N_3117,N_4222);
nand U5385 (N_5385,N_4094,N_3917);
or U5386 (N_5386,N_3818,N_3193);
nor U5387 (N_5387,N_3862,N_3902);
and U5388 (N_5388,N_4405,N_4318);
or U5389 (N_5389,N_4337,N_3092);
xnor U5390 (N_5390,N_3758,N_3666);
nand U5391 (N_5391,N_3232,N_4087);
nor U5392 (N_5392,N_4101,N_3901);
and U5393 (N_5393,N_3889,N_3834);
nand U5394 (N_5394,N_4417,N_3094);
nor U5395 (N_5395,N_3689,N_4346);
or U5396 (N_5396,N_3420,N_3323);
and U5397 (N_5397,N_3501,N_3639);
and U5398 (N_5398,N_4175,N_4354);
and U5399 (N_5399,N_3233,N_4405);
nor U5400 (N_5400,N_4300,N_4350);
or U5401 (N_5401,N_4341,N_3773);
and U5402 (N_5402,N_3186,N_4270);
and U5403 (N_5403,N_4227,N_3799);
or U5404 (N_5404,N_3092,N_3127);
nor U5405 (N_5405,N_4035,N_3174);
nand U5406 (N_5406,N_3758,N_3154);
nand U5407 (N_5407,N_3425,N_3173);
nand U5408 (N_5408,N_3409,N_3912);
nor U5409 (N_5409,N_3654,N_3797);
xor U5410 (N_5410,N_4482,N_3586);
nor U5411 (N_5411,N_3841,N_3182);
nor U5412 (N_5412,N_3149,N_4443);
and U5413 (N_5413,N_4277,N_3411);
nor U5414 (N_5414,N_3385,N_3475);
nand U5415 (N_5415,N_4416,N_4314);
nand U5416 (N_5416,N_3379,N_3834);
or U5417 (N_5417,N_3824,N_3712);
xor U5418 (N_5418,N_4273,N_3050);
nand U5419 (N_5419,N_3071,N_4087);
or U5420 (N_5420,N_4496,N_3965);
nor U5421 (N_5421,N_3121,N_3257);
xnor U5422 (N_5422,N_4470,N_3384);
nand U5423 (N_5423,N_3390,N_4121);
and U5424 (N_5424,N_4033,N_3804);
and U5425 (N_5425,N_4086,N_3157);
and U5426 (N_5426,N_3910,N_3570);
or U5427 (N_5427,N_3279,N_3571);
nand U5428 (N_5428,N_3134,N_4130);
xnor U5429 (N_5429,N_3192,N_3349);
or U5430 (N_5430,N_3118,N_4012);
nor U5431 (N_5431,N_3917,N_3472);
and U5432 (N_5432,N_3297,N_3420);
nor U5433 (N_5433,N_3577,N_4079);
nand U5434 (N_5434,N_4366,N_3523);
and U5435 (N_5435,N_3061,N_4319);
nand U5436 (N_5436,N_3610,N_3887);
nor U5437 (N_5437,N_3932,N_3737);
nand U5438 (N_5438,N_3302,N_3057);
or U5439 (N_5439,N_3981,N_3154);
and U5440 (N_5440,N_3289,N_3632);
nor U5441 (N_5441,N_3888,N_4232);
nand U5442 (N_5442,N_3761,N_3546);
and U5443 (N_5443,N_4362,N_3609);
nand U5444 (N_5444,N_4371,N_3894);
nand U5445 (N_5445,N_4098,N_3705);
nand U5446 (N_5446,N_4230,N_3154);
xnor U5447 (N_5447,N_4371,N_4495);
or U5448 (N_5448,N_4367,N_4217);
nand U5449 (N_5449,N_3025,N_3597);
nand U5450 (N_5450,N_3500,N_4198);
or U5451 (N_5451,N_4374,N_4298);
or U5452 (N_5452,N_4173,N_3354);
nor U5453 (N_5453,N_4350,N_3219);
or U5454 (N_5454,N_4185,N_4201);
and U5455 (N_5455,N_3370,N_3780);
xnor U5456 (N_5456,N_3949,N_3602);
and U5457 (N_5457,N_3273,N_4147);
nand U5458 (N_5458,N_4044,N_4352);
or U5459 (N_5459,N_3121,N_3322);
or U5460 (N_5460,N_4081,N_3671);
xnor U5461 (N_5461,N_3679,N_3315);
or U5462 (N_5462,N_3238,N_3902);
nor U5463 (N_5463,N_3552,N_3244);
or U5464 (N_5464,N_3096,N_4484);
nor U5465 (N_5465,N_4344,N_4244);
nand U5466 (N_5466,N_3344,N_4267);
xor U5467 (N_5467,N_3975,N_3490);
and U5468 (N_5468,N_4045,N_3997);
xor U5469 (N_5469,N_3855,N_3757);
and U5470 (N_5470,N_3301,N_4088);
xor U5471 (N_5471,N_3052,N_3994);
nor U5472 (N_5472,N_3825,N_3584);
or U5473 (N_5473,N_4374,N_3270);
nand U5474 (N_5474,N_3318,N_4409);
nand U5475 (N_5475,N_3863,N_3288);
or U5476 (N_5476,N_4415,N_4324);
nor U5477 (N_5477,N_4499,N_3037);
and U5478 (N_5478,N_3580,N_4078);
xor U5479 (N_5479,N_4423,N_4292);
xnor U5480 (N_5480,N_3137,N_3006);
nor U5481 (N_5481,N_3550,N_4222);
and U5482 (N_5482,N_3639,N_4123);
and U5483 (N_5483,N_3413,N_3805);
nand U5484 (N_5484,N_4228,N_3158);
nand U5485 (N_5485,N_3702,N_3198);
and U5486 (N_5486,N_3833,N_3775);
nand U5487 (N_5487,N_3850,N_4440);
nor U5488 (N_5488,N_4169,N_3122);
nor U5489 (N_5489,N_4114,N_4322);
and U5490 (N_5490,N_3470,N_4082);
nand U5491 (N_5491,N_4123,N_3280);
nor U5492 (N_5492,N_3668,N_4336);
or U5493 (N_5493,N_3701,N_3014);
nor U5494 (N_5494,N_3851,N_3292);
nand U5495 (N_5495,N_3715,N_4180);
and U5496 (N_5496,N_4498,N_3796);
nor U5497 (N_5497,N_4328,N_3946);
nor U5498 (N_5498,N_3456,N_4187);
and U5499 (N_5499,N_4199,N_3880);
nor U5500 (N_5500,N_3416,N_3911);
xor U5501 (N_5501,N_3264,N_3107);
and U5502 (N_5502,N_3414,N_4393);
and U5503 (N_5503,N_3436,N_4469);
nor U5504 (N_5504,N_3607,N_3661);
and U5505 (N_5505,N_4361,N_3168);
and U5506 (N_5506,N_4092,N_3362);
or U5507 (N_5507,N_3788,N_3981);
xnor U5508 (N_5508,N_3306,N_3923);
and U5509 (N_5509,N_4233,N_4020);
and U5510 (N_5510,N_3990,N_4436);
or U5511 (N_5511,N_3741,N_3931);
nor U5512 (N_5512,N_3226,N_4029);
or U5513 (N_5513,N_4212,N_3865);
xnor U5514 (N_5514,N_4279,N_3954);
nand U5515 (N_5515,N_3507,N_4214);
nor U5516 (N_5516,N_4378,N_3363);
xor U5517 (N_5517,N_3159,N_3748);
xnor U5518 (N_5518,N_3111,N_3729);
nand U5519 (N_5519,N_3731,N_3225);
or U5520 (N_5520,N_4242,N_3893);
or U5521 (N_5521,N_4148,N_4226);
and U5522 (N_5522,N_4129,N_3328);
nor U5523 (N_5523,N_4142,N_3412);
xor U5524 (N_5524,N_4134,N_3801);
xor U5525 (N_5525,N_3187,N_3434);
xnor U5526 (N_5526,N_3994,N_3959);
nor U5527 (N_5527,N_4410,N_4031);
xnor U5528 (N_5528,N_3227,N_3441);
nor U5529 (N_5529,N_4408,N_3163);
and U5530 (N_5530,N_3409,N_3408);
xnor U5531 (N_5531,N_3372,N_3253);
or U5532 (N_5532,N_3678,N_3510);
and U5533 (N_5533,N_4044,N_4270);
nor U5534 (N_5534,N_3095,N_4306);
and U5535 (N_5535,N_4184,N_3833);
or U5536 (N_5536,N_4046,N_3012);
nor U5537 (N_5537,N_4188,N_3432);
xor U5538 (N_5538,N_3827,N_4211);
nor U5539 (N_5539,N_3749,N_4482);
nand U5540 (N_5540,N_4168,N_4082);
and U5541 (N_5541,N_4004,N_3334);
xnor U5542 (N_5542,N_3596,N_4457);
nor U5543 (N_5543,N_3031,N_4340);
xnor U5544 (N_5544,N_3560,N_4006);
and U5545 (N_5545,N_3768,N_3954);
nor U5546 (N_5546,N_3568,N_4242);
and U5547 (N_5547,N_3643,N_3527);
and U5548 (N_5548,N_4315,N_3545);
xnor U5549 (N_5549,N_3334,N_3619);
and U5550 (N_5550,N_3570,N_3344);
nor U5551 (N_5551,N_4296,N_3714);
and U5552 (N_5552,N_3123,N_4366);
nand U5553 (N_5553,N_3364,N_3613);
or U5554 (N_5554,N_3317,N_3607);
or U5555 (N_5555,N_3980,N_4264);
xnor U5556 (N_5556,N_3526,N_3976);
nor U5557 (N_5557,N_4372,N_3442);
or U5558 (N_5558,N_4099,N_4231);
xnor U5559 (N_5559,N_4033,N_3648);
nand U5560 (N_5560,N_4298,N_4079);
and U5561 (N_5561,N_3580,N_3547);
or U5562 (N_5562,N_3934,N_4076);
nor U5563 (N_5563,N_3742,N_3943);
nor U5564 (N_5564,N_3679,N_3891);
and U5565 (N_5565,N_3766,N_3615);
or U5566 (N_5566,N_3663,N_4373);
and U5567 (N_5567,N_3686,N_3262);
and U5568 (N_5568,N_3332,N_3856);
and U5569 (N_5569,N_4419,N_3472);
xnor U5570 (N_5570,N_4106,N_3279);
and U5571 (N_5571,N_3394,N_3447);
nand U5572 (N_5572,N_3353,N_4484);
or U5573 (N_5573,N_3694,N_3070);
nor U5574 (N_5574,N_3492,N_3560);
nand U5575 (N_5575,N_3605,N_3753);
nand U5576 (N_5576,N_4183,N_3087);
nand U5577 (N_5577,N_4480,N_4309);
or U5578 (N_5578,N_3298,N_3527);
nor U5579 (N_5579,N_4365,N_3766);
or U5580 (N_5580,N_4424,N_4386);
xnor U5581 (N_5581,N_3139,N_4233);
nor U5582 (N_5582,N_3186,N_3730);
and U5583 (N_5583,N_4151,N_4118);
xnor U5584 (N_5584,N_3479,N_3854);
nor U5585 (N_5585,N_3330,N_4472);
nor U5586 (N_5586,N_4413,N_3597);
nand U5587 (N_5587,N_4280,N_3004);
xor U5588 (N_5588,N_3528,N_4464);
nand U5589 (N_5589,N_3500,N_3016);
or U5590 (N_5590,N_4087,N_3613);
nor U5591 (N_5591,N_3323,N_4389);
nand U5592 (N_5592,N_3751,N_4350);
xor U5593 (N_5593,N_3562,N_3844);
and U5594 (N_5594,N_4185,N_4480);
and U5595 (N_5595,N_4164,N_4206);
or U5596 (N_5596,N_3705,N_3093);
xnor U5597 (N_5597,N_4287,N_4227);
or U5598 (N_5598,N_3634,N_3306);
xor U5599 (N_5599,N_3300,N_3475);
nor U5600 (N_5600,N_3040,N_4181);
xor U5601 (N_5601,N_3947,N_3442);
nand U5602 (N_5602,N_4345,N_4274);
xnor U5603 (N_5603,N_3175,N_4142);
nor U5604 (N_5604,N_4086,N_4208);
xnor U5605 (N_5605,N_4338,N_3261);
or U5606 (N_5606,N_3358,N_3308);
nor U5607 (N_5607,N_3178,N_3401);
nand U5608 (N_5608,N_4318,N_3536);
or U5609 (N_5609,N_3810,N_3456);
nor U5610 (N_5610,N_3574,N_3381);
nand U5611 (N_5611,N_3078,N_3685);
or U5612 (N_5612,N_4276,N_3506);
or U5613 (N_5613,N_3588,N_4434);
nand U5614 (N_5614,N_3777,N_3928);
or U5615 (N_5615,N_4301,N_3190);
or U5616 (N_5616,N_3336,N_3729);
nor U5617 (N_5617,N_4436,N_3347);
and U5618 (N_5618,N_3082,N_3941);
nor U5619 (N_5619,N_4234,N_3743);
and U5620 (N_5620,N_4014,N_3903);
nand U5621 (N_5621,N_3942,N_4434);
or U5622 (N_5622,N_4281,N_3624);
and U5623 (N_5623,N_3060,N_3143);
nand U5624 (N_5624,N_3842,N_3941);
nor U5625 (N_5625,N_3323,N_3088);
nor U5626 (N_5626,N_3580,N_4130);
nand U5627 (N_5627,N_3262,N_4044);
nor U5628 (N_5628,N_3546,N_3291);
nor U5629 (N_5629,N_3705,N_4368);
and U5630 (N_5630,N_4403,N_3996);
and U5631 (N_5631,N_3179,N_3978);
nand U5632 (N_5632,N_3720,N_3055);
xor U5633 (N_5633,N_3760,N_3605);
nor U5634 (N_5634,N_3075,N_3122);
or U5635 (N_5635,N_3741,N_4269);
and U5636 (N_5636,N_3214,N_3139);
nand U5637 (N_5637,N_4390,N_3235);
nand U5638 (N_5638,N_3320,N_3501);
or U5639 (N_5639,N_3580,N_4312);
or U5640 (N_5640,N_3682,N_3441);
and U5641 (N_5641,N_3674,N_3822);
or U5642 (N_5642,N_4282,N_3106);
or U5643 (N_5643,N_4327,N_3232);
nand U5644 (N_5644,N_3831,N_3360);
xor U5645 (N_5645,N_4099,N_4212);
nand U5646 (N_5646,N_3881,N_3542);
nand U5647 (N_5647,N_4150,N_3464);
nor U5648 (N_5648,N_3152,N_3876);
nor U5649 (N_5649,N_3694,N_3390);
or U5650 (N_5650,N_3979,N_4298);
nand U5651 (N_5651,N_3400,N_3139);
nand U5652 (N_5652,N_3696,N_4361);
or U5653 (N_5653,N_3290,N_3264);
nor U5654 (N_5654,N_4278,N_4075);
nand U5655 (N_5655,N_3879,N_3982);
nand U5656 (N_5656,N_3210,N_3967);
nor U5657 (N_5657,N_3491,N_3084);
and U5658 (N_5658,N_3293,N_3101);
xor U5659 (N_5659,N_3171,N_3592);
and U5660 (N_5660,N_3877,N_3123);
or U5661 (N_5661,N_4150,N_3764);
nor U5662 (N_5662,N_3722,N_4102);
or U5663 (N_5663,N_3506,N_3618);
nor U5664 (N_5664,N_3938,N_4479);
and U5665 (N_5665,N_3296,N_3466);
xor U5666 (N_5666,N_4027,N_3922);
and U5667 (N_5667,N_3709,N_3947);
and U5668 (N_5668,N_3596,N_4381);
or U5669 (N_5669,N_3017,N_4137);
xor U5670 (N_5670,N_3389,N_4439);
and U5671 (N_5671,N_3554,N_4207);
nand U5672 (N_5672,N_4258,N_4295);
or U5673 (N_5673,N_4236,N_3155);
xor U5674 (N_5674,N_3957,N_4355);
nand U5675 (N_5675,N_3167,N_3444);
and U5676 (N_5676,N_3589,N_4395);
and U5677 (N_5677,N_3103,N_3781);
nor U5678 (N_5678,N_3377,N_3174);
and U5679 (N_5679,N_3149,N_3352);
and U5680 (N_5680,N_3072,N_3499);
nor U5681 (N_5681,N_3379,N_3325);
nand U5682 (N_5682,N_3453,N_4178);
nand U5683 (N_5683,N_3594,N_3464);
xnor U5684 (N_5684,N_4365,N_4220);
and U5685 (N_5685,N_4015,N_4181);
or U5686 (N_5686,N_3049,N_4087);
xnor U5687 (N_5687,N_4376,N_3691);
xnor U5688 (N_5688,N_3911,N_4420);
nor U5689 (N_5689,N_3961,N_3987);
or U5690 (N_5690,N_3995,N_3424);
nand U5691 (N_5691,N_3527,N_3394);
xor U5692 (N_5692,N_4230,N_3537);
or U5693 (N_5693,N_3275,N_4493);
and U5694 (N_5694,N_4449,N_3322);
xnor U5695 (N_5695,N_3598,N_3072);
xnor U5696 (N_5696,N_3908,N_3631);
nand U5697 (N_5697,N_3213,N_3498);
nand U5698 (N_5698,N_3679,N_4189);
xnor U5699 (N_5699,N_3589,N_3216);
nor U5700 (N_5700,N_3058,N_3831);
nor U5701 (N_5701,N_3156,N_4441);
xor U5702 (N_5702,N_3061,N_4161);
nand U5703 (N_5703,N_4287,N_4382);
or U5704 (N_5704,N_3586,N_3508);
or U5705 (N_5705,N_3450,N_4322);
nand U5706 (N_5706,N_4130,N_3000);
and U5707 (N_5707,N_4080,N_3202);
or U5708 (N_5708,N_3478,N_4097);
xor U5709 (N_5709,N_4434,N_3955);
or U5710 (N_5710,N_3282,N_4194);
xnor U5711 (N_5711,N_3667,N_4440);
nor U5712 (N_5712,N_3018,N_3780);
nor U5713 (N_5713,N_3559,N_3633);
nor U5714 (N_5714,N_3985,N_3970);
or U5715 (N_5715,N_3608,N_3016);
nand U5716 (N_5716,N_3276,N_4491);
and U5717 (N_5717,N_4140,N_4218);
nand U5718 (N_5718,N_3546,N_3677);
nand U5719 (N_5719,N_4162,N_3702);
nor U5720 (N_5720,N_3087,N_3647);
and U5721 (N_5721,N_4347,N_4042);
xor U5722 (N_5722,N_3822,N_3099);
nor U5723 (N_5723,N_3446,N_4047);
nor U5724 (N_5724,N_3647,N_4082);
nor U5725 (N_5725,N_3031,N_3645);
nand U5726 (N_5726,N_3564,N_4029);
nor U5727 (N_5727,N_4371,N_3150);
xor U5728 (N_5728,N_3828,N_4271);
xnor U5729 (N_5729,N_3230,N_3716);
xor U5730 (N_5730,N_3506,N_3753);
xor U5731 (N_5731,N_3098,N_3086);
or U5732 (N_5732,N_4417,N_4267);
and U5733 (N_5733,N_4488,N_3101);
and U5734 (N_5734,N_3611,N_3887);
nand U5735 (N_5735,N_3086,N_3344);
and U5736 (N_5736,N_3643,N_3310);
nor U5737 (N_5737,N_3567,N_3605);
nand U5738 (N_5738,N_3806,N_3717);
xnor U5739 (N_5739,N_4209,N_3015);
or U5740 (N_5740,N_4061,N_4023);
nor U5741 (N_5741,N_3172,N_3132);
xnor U5742 (N_5742,N_4124,N_3016);
nand U5743 (N_5743,N_3224,N_3811);
and U5744 (N_5744,N_3789,N_3572);
and U5745 (N_5745,N_3013,N_3664);
xnor U5746 (N_5746,N_3289,N_3128);
xor U5747 (N_5747,N_3661,N_3782);
or U5748 (N_5748,N_4169,N_3777);
xor U5749 (N_5749,N_3167,N_4115);
xor U5750 (N_5750,N_4195,N_4303);
or U5751 (N_5751,N_3661,N_4094);
or U5752 (N_5752,N_4054,N_3765);
xnor U5753 (N_5753,N_3453,N_3708);
nor U5754 (N_5754,N_3590,N_3198);
nor U5755 (N_5755,N_4168,N_3306);
nand U5756 (N_5756,N_4267,N_3672);
nand U5757 (N_5757,N_3298,N_3519);
nand U5758 (N_5758,N_3985,N_3789);
and U5759 (N_5759,N_3342,N_3578);
xnor U5760 (N_5760,N_4444,N_4309);
or U5761 (N_5761,N_3138,N_3249);
or U5762 (N_5762,N_3687,N_3549);
and U5763 (N_5763,N_4122,N_3191);
and U5764 (N_5764,N_4137,N_3456);
xnor U5765 (N_5765,N_4366,N_3655);
nor U5766 (N_5766,N_3794,N_4153);
and U5767 (N_5767,N_3970,N_4218);
xnor U5768 (N_5768,N_3846,N_3961);
nand U5769 (N_5769,N_3909,N_3451);
or U5770 (N_5770,N_3123,N_3451);
or U5771 (N_5771,N_3352,N_4475);
and U5772 (N_5772,N_3971,N_3014);
xor U5773 (N_5773,N_3106,N_4249);
and U5774 (N_5774,N_4208,N_4053);
nor U5775 (N_5775,N_4128,N_3981);
and U5776 (N_5776,N_3147,N_3547);
or U5777 (N_5777,N_3371,N_3278);
and U5778 (N_5778,N_3003,N_3178);
xnor U5779 (N_5779,N_4024,N_3602);
and U5780 (N_5780,N_3380,N_3096);
xnor U5781 (N_5781,N_4214,N_3168);
or U5782 (N_5782,N_3878,N_4094);
nor U5783 (N_5783,N_3117,N_4474);
xor U5784 (N_5784,N_3648,N_3407);
or U5785 (N_5785,N_3415,N_4176);
or U5786 (N_5786,N_3166,N_4467);
nand U5787 (N_5787,N_3086,N_3718);
nor U5788 (N_5788,N_3424,N_4345);
nand U5789 (N_5789,N_3815,N_3951);
nor U5790 (N_5790,N_3734,N_3080);
and U5791 (N_5791,N_3264,N_3349);
nand U5792 (N_5792,N_3895,N_3803);
nand U5793 (N_5793,N_4264,N_4338);
xor U5794 (N_5794,N_3174,N_3281);
nor U5795 (N_5795,N_3432,N_3833);
or U5796 (N_5796,N_3681,N_3148);
xnor U5797 (N_5797,N_3337,N_3518);
xnor U5798 (N_5798,N_3102,N_4394);
nor U5799 (N_5799,N_3445,N_3578);
xnor U5800 (N_5800,N_3283,N_3617);
nor U5801 (N_5801,N_3501,N_3293);
or U5802 (N_5802,N_4021,N_3630);
and U5803 (N_5803,N_4305,N_4188);
nand U5804 (N_5804,N_3387,N_3861);
nand U5805 (N_5805,N_4255,N_4156);
nand U5806 (N_5806,N_4236,N_4350);
and U5807 (N_5807,N_3524,N_3248);
or U5808 (N_5808,N_3015,N_3503);
xnor U5809 (N_5809,N_4200,N_4096);
nand U5810 (N_5810,N_4116,N_4139);
nor U5811 (N_5811,N_3857,N_3317);
nor U5812 (N_5812,N_4270,N_3834);
nor U5813 (N_5813,N_4267,N_4189);
or U5814 (N_5814,N_3959,N_3330);
xor U5815 (N_5815,N_4391,N_3430);
xor U5816 (N_5816,N_3483,N_3918);
xor U5817 (N_5817,N_3477,N_3769);
nand U5818 (N_5818,N_4042,N_3317);
xor U5819 (N_5819,N_4185,N_3776);
xor U5820 (N_5820,N_4482,N_4389);
or U5821 (N_5821,N_3180,N_4178);
xor U5822 (N_5822,N_3689,N_4246);
nor U5823 (N_5823,N_4047,N_3821);
and U5824 (N_5824,N_4190,N_4415);
or U5825 (N_5825,N_3438,N_4419);
xor U5826 (N_5826,N_4074,N_4262);
and U5827 (N_5827,N_3246,N_3124);
nor U5828 (N_5828,N_3276,N_4243);
nand U5829 (N_5829,N_3708,N_3785);
nand U5830 (N_5830,N_4096,N_3136);
xor U5831 (N_5831,N_3856,N_3641);
xor U5832 (N_5832,N_4362,N_3807);
and U5833 (N_5833,N_4428,N_4075);
xnor U5834 (N_5834,N_3159,N_3377);
or U5835 (N_5835,N_3250,N_3443);
nand U5836 (N_5836,N_4105,N_4402);
nor U5837 (N_5837,N_3965,N_3385);
xnor U5838 (N_5838,N_4193,N_3211);
nand U5839 (N_5839,N_3814,N_3913);
and U5840 (N_5840,N_3725,N_3251);
and U5841 (N_5841,N_4001,N_4404);
xor U5842 (N_5842,N_4287,N_4309);
and U5843 (N_5843,N_3703,N_3080);
nor U5844 (N_5844,N_4258,N_4058);
and U5845 (N_5845,N_3158,N_3622);
nand U5846 (N_5846,N_4031,N_3461);
xor U5847 (N_5847,N_3599,N_3584);
and U5848 (N_5848,N_3303,N_3632);
nor U5849 (N_5849,N_4206,N_4186);
nor U5850 (N_5850,N_3633,N_3562);
xor U5851 (N_5851,N_4222,N_4191);
nand U5852 (N_5852,N_3335,N_4021);
nand U5853 (N_5853,N_4321,N_3968);
and U5854 (N_5854,N_3780,N_4309);
and U5855 (N_5855,N_4268,N_4472);
nor U5856 (N_5856,N_4051,N_3766);
xor U5857 (N_5857,N_3212,N_3679);
nand U5858 (N_5858,N_4153,N_4260);
nor U5859 (N_5859,N_4138,N_3394);
nor U5860 (N_5860,N_3305,N_4177);
or U5861 (N_5861,N_3750,N_3575);
xnor U5862 (N_5862,N_4018,N_3417);
and U5863 (N_5863,N_4382,N_4200);
or U5864 (N_5864,N_3730,N_3902);
nor U5865 (N_5865,N_4015,N_3188);
nor U5866 (N_5866,N_3084,N_3779);
and U5867 (N_5867,N_4156,N_4170);
nor U5868 (N_5868,N_3052,N_3277);
nand U5869 (N_5869,N_3875,N_4120);
and U5870 (N_5870,N_3972,N_3190);
nand U5871 (N_5871,N_3755,N_4173);
xnor U5872 (N_5872,N_4078,N_3355);
and U5873 (N_5873,N_4332,N_4222);
xor U5874 (N_5874,N_3815,N_3226);
or U5875 (N_5875,N_3895,N_3038);
or U5876 (N_5876,N_3711,N_3834);
and U5877 (N_5877,N_3689,N_3692);
xnor U5878 (N_5878,N_4120,N_3629);
nand U5879 (N_5879,N_3979,N_4106);
nor U5880 (N_5880,N_3084,N_3514);
or U5881 (N_5881,N_3511,N_3395);
or U5882 (N_5882,N_3578,N_3736);
and U5883 (N_5883,N_3897,N_3793);
xnor U5884 (N_5884,N_4429,N_3262);
nand U5885 (N_5885,N_3908,N_3248);
or U5886 (N_5886,N_3969,N_3138);
or U5887 (N_5887,N_3841,N_4095);
nand U5888 (N_5888,N_4375,N_3111);
nor U5889 (N_5889,N_3930,N_3567);
or U5890 (N_5890,N_3641,N_4210);
nand U5891 (N_5891,N_4367,N_3557);
and U5892 (N_5892,N_4449,N_3882);
xnor U5893 (N_5893,N_3062,N_4337);
and U5894 (N_5894,N_3539,N_3732);
xor U5895 (N_5895,N_3568,N_3548);
nor U5896 (N_5896,N_4226,N_3048);
nand U5897 (N_5897,N_3399,N_3203);
xor U5898 (N_5898,N_3813,N_4382);
and U5899 (N_5899,N_3472,N_4276);
xnor U5900 (N_5900,N_3593,N_4025);
nand U5901 (N_5901,N_4381,N_3758);
and U5902 (N_5902,N_3164,N_3282);
or U5903 (N_5903,N_3677,N_3932);
and U5904 (N_5904,N_3996,N_3563);
or U5905 (N_5905,N_3186,N_4352);
nor U5906 (N_5906,N_4098,N_3254);
nand U5907 (N_5907,N_3875,N_3281);
nor U5908 (N_5908,N_4268,N_4346);
nor U5909 (N_5909,N_3993,N_3969);
xor U5910 (N_5910,N_3934,N_4183);
nand U5911 (N_5911,N_4125,N_3675);
nor U5912 (N_5912,N_4050,N_3602);
xnor U5913 (N_5913,N_3621,N_3531);
or U5914 (N_5914,N_4175,N_3948);
nor U5915 (N_5915,N_4453,N_3498);
or U5916 (N_5916,N_4250,N_3267);
and U5917 (N_5917,N_4339,N_4025);
and U5918 (N_5918,N_3800,N_3227);
nand U5919 (N_5919,N_4308,N_3421);
xor U5920 (N_5920,N_3688,N_4050);
nor U5921 (N_5921,N_3265,N_3928);
or U5922 (N_5922,N_3519,N_4068);
or U5923 (N_5923,N_3702,N_4374);
or U5924 (N_5924,N_4128,N_3484);
xor U5925 (N_5925,N_3936,N_3176);
nand U5926 (N_5926,N_3449,N_4320);
nand U5927 (N_5927,N_3323,N_3346);
or U5928 (N_5928,N_3107,N_4094);
and U5929 (N_5929,N_4135,N_4313);
and U5930 (N_5930,N_4118,N_4337);
or U5931 (N_5931,N_4262,N_3354);
xor U5932 (N_5932,N_3947,N_3528);
and U5933 (N_5933,N_4329,N_4254);
nand U5934 (N_5934,N_3598,N_3975);
nand U5935 (N_5935,N_3479,N_3488);
xnor U5936 (N_5936,N_3180,N_3807);
xor U5937 (N_5937,N_3639,N_3876);
or U5938 (N_5938,N_3978,N_3505);
nand U5939 (N_5939,N_4246,N_3027);
or U5940 (N_5940,N_3145,N_3161);
nand U5941 (N_5941,N_4460,N_3074);
and U5942 (N_5942,N_4415,N_3397);
and U5943 (N_5943,N_3823,N_3049);
nand U5944 (N_5944,N_3162,N_3397);
or U5945 (N_5945,N_3828,N_4043);
nand U5946 (N_5946,N_3633,N_3195);
xor U5947 (N_5947,N_3766,N_3438);
nand U5948 (N_5948,N_4274,N_3873);
nand U5949 (N_5949,N_3907,N_3123);
xnor U5950 (N_5950,N_4202,N_3413);
nand U5951 (N_5951,N_3130,N_3359);
xor U5952 (N_5952,N_3268,N_4161);
nand U5953 (N_5953,N_3995,N_3604);
xor U5954 (N_5954,N_3907,N_3672);
and U5955 (N_5955,N_3487,N_3177);
and U5956 (N_5956,N_3685,N_3766);
or U5957 (N_5957,N_3993,N_4143);
and U5958 (N_5958,N_3724,N_4431);
nor U5959 (N_5959,N_3102,N_4349);
nand U5960 (N_5960,N_3268,N_3822);
nor U5961 (N_5961,N_3789,N_3606);
and U5962 (N_5962,N_4055,N_3563);
nand U5963 (N_5963,N_4140,N_4397);
and U5964 (N_5964,N_3839,N_4339);
or U5965 (N_5965,N_3748,N_3389);
nor U5966 (N_5966,N_4316,N_4327);
nand U5967 (N_5967,N_3414,N_3380);
nor U5968 (N_5968,N_3184,N_3083);
or U5969 (N_5969,N_3695,N_3530);
or U5970 (N_5970,N_3747,N_3992);
nor U5971 (N_5971,N_3969,N_4104);
xor U5972 (N_5972,N_4391,N_4377);
xor U5973 (N_5973,N_3757,N_4350);
nand U5974 (N_5974,N_3848,N_3169);
and U5975 (N_5975,N_4128,N_3678);
nor U5976 (N_5976,N_4188,N_3519);
xnor U5977 (N_5977,N_4275,N_3464);
xnor U5978 (N_5978,N_3182,N_4362);
and U5979 (N_5979,N_3499,N_3597);
or U5980 (N_5980,N_3815,N_4230);
and U5981 (N_5981,N_4122,N_3033);
xor U5982 (N_5982,N_3618,N_3963);
xnor U5983 (N_5983,N_3565,N_4231);
xnor U5984 (N_5984,N_4133,N_3034);
xnor U5985 (N_5985,N_3578,N_3371);
or U5986 (N_5986,N_4240,N_4224);
or U5987 (N_5987,N_4074,N_3368);
and U5988 (N_5988,N_3056,N_3639);
nand U5989 (N_5989,N_3049,N_4289);
nand U5990 (N_5990,N_3643,N_3751);
nand U5991 (N_5991,N_4427,N_3251);
nor U5992 (N_5992,N_4136,N_4045);
xor U5993 (N_5993,N_3844,N_3334);
and U5994 (N_5994,N_3318,N_3189);
or U5995 (N_5995,N_4217,N_3288);
nor U5996 (N_5996,N_4497,N_3407);
and U5997 (N_5997,N_3925,N_4265);
xnor U5998 (N_5998,N_3039,N_3333);
nor U5999 (N_5999,N_3784,N_3975);
xnor U6000 (N_6000,N_5136,N_4621);
or U6001 (N_6001,N_5916,N_5227);
or U6002 (N_6002,N_5103,N_5390);
and U6003 (N_6003,N_5025,N_4967);
nand U6004 (N_6004,N_5127,N_5878);
or U6005 (N_6005,N_4701,N_5310);
xor U6006 (N_6006,N_5991,N_4812);
and U6007 (N_6007,N_4911,N_5496);
or U6008 (N_6008,N_4732,N_5909);
nor U6009 (N_6009,N_5929,N_5652);
and U6010 (N_6010,N_5234,N_4814);
xnor U6011 (N_6011,N_4971,N_5764);
and U6012 (N_6012,N_5529,N_4596);
xor U6013 (N_6013,N_4841,N_5282);
and U6014 (N_6014,N_5182,N_4548);
nor U6015 (N_6015,N_4510,N_5226);
xor U6016 (N_6016,N_5613,N_5321);
nand U6017 (N_6017,N_5618,N_5525);
nor U6018 (N_6018,N_5352,N_5159);
nor U6019 (N_6019,N_4585,N_5459);
or U6020 (N_6020,N_5960,N_5461);
nand U6021 (N_6021,N_5924,N_4933);
xor U6022 (N_6022,N_5172,N_5162);
and U6023 (N_6023,N_4941,N_5768);
or U6024 (N_6024,N_4910,N_5434);
xnor U6025 (N_6025,N_4724,N_5617);
nand U6026 (N_6026,N_5179,N_5245);
nand U6027 (N_6027,N_4833,N_4736);
and U6028 (N_6028,N_4803,N_4968);
nor U6029 (N_6029,N_5847,N_5448);
xor U6030 (N_6030,N_4892,N_5432);
and U6031 (N_6031,N_5668,N_5985);
or U6032 (N_6032,N_4709,N_4593);
or U6033 (N_6033,N_4738,N_5389);
nand U6034 (N_6034,N_4895,N_5413);
and U6035 (N_6035,N_5160,N_5262);
nor U6036 (N_6036,N_5287,N_5299);
xnor U6037 (N_6037,N_5317,N_5216);
nor U6038 (N_6038,N_4850,N_5962);
xor U6039 (N_6039,N_5697,N_5951);
or U6040 (N_6040,N_5957,N_5830);
xnor U6041 (N_6041,N_4780,N_5372);
nor U6042 (N_6042,N_5480,N_4748);
or U6043 (N_6043,N_4974,N_4707);
nand U6044 (N_6044,N_5938,N_4770);
nand U6045 (N_6045,N_5253,N_5666);
xor U6046 (N_6046,N_5431,N_5521);
nor U6047 (N_6047,N_5414,N_5647);
or U6048 (N_6048,N_5126,N_5501);
xnor U6049 (N_6049,N_5988,N_5391);
nor U6050 (N_6050,N_4702,N_4582);
xor U6051 (N_6051,N_4898,N_4900);
nor U6052 (N_6052,N_5333,N_5087);
xnor U6053 (N_6053,N_5983,N_5889);
nor U6054 (N_6054,N_5005,N_4614);
xnor U6055 (N_6055,N_5114,N_5782);
or U6056 (N_6056,N_5573,N_4986);
or U6057 (N_6057,N_5642,N_5270);
nand U6058 (N_6058,N_5438,N_5837);
xnor U6059 (N_6059,N_4790,N_5732);
nand U6060 (N_6060,N_4729,N_4792);
nand U6061 (N_6061,N_5140,N_5718);
nor U6062 (N_6062,N_4944,N_4563);
and U6063 (N_6063,N_5853,N_5588);
or U6064 (N_6064,N_4540,N_4718);
xor U6065 (N_6065,N_4549,N_5393);
and U6066 (N_6066,N_4849,N_4672);
nand U6067 (N_6067,N_5865,N_5061);
nor U6068 (N_6068,N_5238,N_5728);
xor U6069 (N_6069,N_4581,N_5691);
and U6070 (N_6070,N_5706,N_4637);
or U6071 (N_6071,N_5619,N_5116);
nor U6072 (N_6072,N_5898,N_5774);
xor U6073 (N_6073,N_5311,N_5382);
nand U6074 (N_6074,N_5300,N_5215);
and U6075 (N_6075,N_4514,N_4584);
and U6076 (N_6076,N_4861,N_4807);
and U6077 (N_6077,N_5113,N_5156);
nor U6078 (N_6078,N_5828,N_5435);
nand U6079 (N_6079,N_4851,N_5819);
nor U6080 (N_6080,N_5007,N_5301);
and U6081 (N_6081,N_5604,N_5540);
nand U6082 (N_6082,N_4991,N_4662);
or U6083 (N_6083,N_5967,N_5703);
and U6084 (N_6084,N_4950,N_4570);
xor U6085 (N_6085,N_4726,N_4889);
nor U6086 (N_6086,N_5293,N_5132);
xnor U6087 (N_6087,N_5692,N_5682);
or U6088 (N_6088,N_5646,N_4739);
or U6089 (N_6089,N_5055,N_4901);
xnor U6090 (N_6090,N_4524,N_5188);
or U6091 (N_6091,N_4737,N_5135);
nor U6092 (N_6092,N_5404,N_5729);
or U6093 (N_6093,N_5771,N_4800);
nor U6094 (N_6094,N_5532,N_5765);
nor U6095 (N_6095,N_5142,N_5048);
nor U6096 (N_6096,N_5073,N_5769);
or U6097 (N_6097,N_5096,N_4823);
xor U6098 (N_6098,N_5026,N_5277);
xnor U6099 (N_6099,N_5396,N_5399);
and U6100 (N_6100,N_5328,N_5705);
and U6101 (N_6101,N_4806,N_4537);
nor U6102 (N_6102,N_4542,N_4754);
and U6103 (N_6103,N_5043,N_5428);
or U6104 (N_6104,N_5552,N_5206);
nand U6105 (N_6105,N_4762,N_4728);
nand U6106 (N_6106,N_5046,N_5454);
or U6107 (N_6107,N_5338,N_5809);
nand U6108 (N_6108,N_4560,N_5515);
and U6109 (N_6109,N_5437,N_5063);
nand U6110 (N_6110,N_5637,N_5775);
or U6111 (N_6111,N_5921,N_5392);
nand U6112 (N_6112,N_5799,N_4873);
and U6113 (N_6113,N_5421,N_4503);
nand U6114 (N_6114,N_5365,N_5856);
nor U6115 (N_6115,N_5696,N_5358);
xnor U6116 (N_6116,N_5419,N_5485);
and U6117 (N_6117,N_5152,N_4569);
and U6118 (N_6118,N_5394,N_5109);
nand U6119 (N_6119,N_4880,N_4978);
nand U6120 (N_6120,N_5258,N_5122);
nand U6121 (N_6121,N_4932,N_5045);
nor U6122 (N_6122,N_5385,N_5327);
and U6123 (N_6123,N_4845,N_5336);
and U6124 (N_6124,N_5292,N_5143);
nand U6125 (N_6125,N_5289,N_5543);
xnor U6126 (N_6126,N_5032,N_4970);
xor U6127 (N_6127,N_5850,N_5213);
nor U6128 (N_6128,N_4568,N_5012);
xor U6129 (N_6129,N_4700,N_4506);
or U6130 (N_6130,N_5963,N_4985);
nor U6131 (N_6131,N_4987,N_4964);
and U6132 (N_6132,N_5244,N_5243);
and U6133 (N_6133,N_4763,N_5915);
xor U6134 (N_6134,N_5731,N_4714);
nor U6135 (N_6135,N_4886,N_5084);
or U6136 (N_6136,N_4599,N_5675);
nor U6137 (N_6137,N_5357,N_5319);
and U6138 (N_6138,N_5019,N_5631);
and U6139 (N_6139,N_5773,N_5939);
nor U6140 (N_6140,N_5551,N_5651);
nor U6141 (N_6141,N_4559,N_5458);
xnor U6142 (N_6142,N_5037,N_5209);
and U6143 (N_6143,N_4558,N_5316);
nand U6144 (N_6144,N_5247,N_5934);
or U6145 (N_6145,N_5513,N_5484);
or U6146 (N_6146,N_5449,N_5595);
and U6147 (N_6147,N_5306,N_4578);
and U6148 (N_6148,N_5498,N_4867);
xor U6149 (N_6149,N_5836,N_4580);
xnor U6150 (N_6150,N_5408,N_5488);
xor U6151 (N_6151,N_4645,N_5749);
xor U6152 (N_6152,N_5469,N_5423);
nand U6153 (N_6153,N_5854,N_4517);
or U6154 (N_6154,N_5883,N_5153);
nand U6155 (N_6155,N_5895,N_5362);
nor U6156 (N_6156,N_5871,N_4694);
nand U6157 (N_6157,N_4550,N_5777);
nor U6158 (N_6158,N_4853,N_4866);
nand U6159 (N_6159,N_5332,N_4627);
xor U6160 (N_6160,N_5817,N_5489);
xnor U6161 (N_6161,N_5430,N_4538);
nor U6162 (N_6162,N_5471,N_4544);
nor U6163 (N_6163,N_5189,N_5776);
nand U6164 (N_6164,N_4612,N_5455);
nor U6165 (N_6165,N_5487,N_4766);
xor U6166 (N_6166,N_5383,N_5843);
or U6167 (N_6167,N_5173,N_4565);
nand U6168 (N_6168,N_5516,N_5091);
xor U6169 (N_6169,N_5767,N_5246);
and U6170 (N_6170,N_4904,N_4797);
or U6171 (N_6171,N_5526,N_4528);
xor U6172 (N_6172,N_5584,N_5254);
nand U6173 (N_6173,N_5908,N_4505);
or U6174 (N_6174,N_5196,N_4830);
xor U6175 (N_6175,N_5914,N_4894);
nand U6176 (N_6176,N_4551,N_5740);
nor U6177 (N_6177,N_5470,N_5344);
xnor U6178 (N_6178,N_5267,N_5639);
xnor U6179 (N_6179,N_5948,N_5147);
or U6180 (N_6180,N_5861,N_5881);
nand U6181 (N_6181,N_4740,N_5743);
nand U6182 (N_6182,N_5761,N_5686);
and U6183 (N_6183,N_5266,N_5466);
and U6184 (N_6184,N_5356,N_4990);
nand U6185 (N_6185,N_5904,N_5912);
and U6186 (N_6186,N_4647,N_5574);
nor U6187 (N_6187,N_5190,N_4864);
xor U6188 (N_6188,N_5279,N_5309);
nand U6189 (N_6189,N_5911,N_5330);
xnor U6190 (N_6190,N_4798,N_4523);
and U6191 (N_6191,N_5973,N_5214);
and U6192 (N_6192,N_4883,N_5659);
and U6193 (N_6193,N_5022,N_4522);
xor U6194 (N_6194,N_5814,N_5553);
xor U6195 (N_6195,N_5753,N_4843);
or U6196 (N_6196,N_5987,N_5313);
and U6197 (N_6197,N_5260,N_5715);
nor U6198 (N_6198,N_5542,N_4888);
and U6199 (N_6199,N_4715,N_5677);
nor U6200 (N_6200,N_4896,N_4882);
and U6201 (N_6201,N_5971,N_4553);
nand U6202 (N_6202,N_5994,N_4682);
and U6203 (N_6203,N_5822,N_5069);
and U6204 (N_6204,N_4855,N_5401);
or U6205 (N_6205,N_5165,N_4785);
and U6206 (N_6206,N_5020,N_5681);
and U6207 (N_6207,N_5980,N_5474);
and U6208 (N_6208,N_5242,N_5802);
and U6209 (N_6209,N_5680,N_5068);
nand U6210 (N_6210,N_5101,N_4781);
or U6211 (N_6211,N_4905,N_4848);
nand U6212 (N_6212,N_4652,N_5925);
xnor U6213 (N_6213,N_4535,N_5024);
xnor U6214 (N_6214,N_5636,N_5578);
and U6215 (N_6215,N_4623,N_5033);
or U6216 (N_6216,N_5086,N_4742);
nor U6217 (N_6217,N_5166,N_5996);
xor U6218 (N_6218,N_5472,N_5566);
xor U6219 (N_6219,N_4995,N_4897);
or U6220 (N_6220,N_5931,N_5150);
nor U6221 (N_6221,N_5905,N_5935);
and U6222 (N_6222,N_5842,N_5755);
nand U6223 (N_6223,N_4717,N_5679);
nand U6224 (N_6224,N_5285,N_5972);
nor U6225 (N_6225,N_5491,N_5427);
nor U6226 (N_6226,N_5808,N_5855);
nor U6227 (N_6227,N_5082,N_5936);
and U6228 (N_6228,N_5707,N_5118);
and U6229 (N_6229,N_5593,N_5123);
and U6230 (N_6230,N_4519,N_4829);
and U6231 (N_6231,N_5120,N_5514);
or U6232 (N_6232,N_5756,N_5548);
nand U6233 (N_6233,N_4981,N_4712);
and U6234 (N_6234,N_4509,N_4607);
xnor U6235 (N_6235,N_5323,N_4909);
xnor U6236 (N_6236,N_4872,N_5483);
or U6237 (N_6237,N_4928,N_4711);
nand U6238 (N_6238,N_5504,N_5575);
xnor U6239 (N_6239,N_5351,N_4828);
nor U6240 (N_6240,N_4821,N_5104);
and U6241 (N_6241,N_5239,N_5256);
nand U6242 (N_6242,N_5608,N_4959);
and U6243 (N_6243,N_5088,N_5900);
xnor U6244 (N_6244,N_4648,N_5687);
nor U6245 (N_6245,N_4634,N_5410);
nor U6246 (N_6246,N_4720,N_5602);
nor U6247 (N_6247,N_4816,N_5549);
or U6248 (N_6248,N_5121,N_5630);
and U6249 (N_6249,N_4692,N_4907);
xor U6250 (N_6250,N_4969,N_5700);
or U6251 (N_6251,N_5559,N_4778);
xor U6252 (N_6252,N_4500,N_4541);
and U6253 (N_6253,N_5056,N_5535);
nor U6254 (N_6254,N_4539,N_5500);
nand U6255 (N_6255,N_5318,N_5094);
xor U6256 (N_6256,N_5479,N_5337);
nand U6257 (N_6257,N_4604,N_5719);
nand U6258 (N_6258,N_5654,N_4730);
nand U6259 (N_6259,N_5062,N_5028);
xnor U6260 (N_6260,N_5537,N_4638);
xor U6261 (N_6261,N_4917,N_5265);
nand U6262 (N_6262,N_5629,N_5149);
or U6263 (N_6263,N_4681,N_5615);
nor U6264 (N_6264,N_5952,N_5065);
and U6265 (N_6265,N_4779,N_5494);
and U6266 (N_6266,N_5374,N_5272);
nor U6267 (N_6267,N_5252,N_4617);
nor U6268 (N_6268,N_5841,N_5581);
xnor U6269 (N_6269,N_4914,N_5997);
xnor U6270 (N_6270,N_4751,N_4804);
xnor U6271 (N_6271,N_4605,N_4719);
or U6272 (N_6272,N_5294,N_4608);
nor U6273 (N_6273,N_5597,N_4639);
or U6274 (N_6274,N_5864,N_5560);
or U6275 (N_6275,N_4773,N_5711);
nand U6276 (N_6276,N_5493,N_5436);
or U6277 (N_6277,N_5119,N_4994);
nand U6278 (N_6278,N_5857,N_5168);
or U6279 (N_6279,N_5801,N_5286);
and U6280 (N_6280,N_5250,N_4508);
xor U6281 (N_6281,N_5251,N_5187);
and U6282 (N_6282,N_5353,N_4590);
nor U6283 (N_6283,N_5240,N_4939);
nor U6284 (N_6284,N_5657,N_5606);
nand U6285 (N_6285,N_4699,N_4735);
nand U6286 (N_6286,N_4965,N_5704);
nor U6287 (N_6287,N_5770,N_5018);
or U6288 (N_6288,N_5497,N_5860);
xor U6289 (N_6289,N_5913,N_5820);
xor U6290 (N_6290,N_5102,N_4511);
nand U6291 (N_6291,N_4741,N_4870);
xnor U6292 (N_6292,N_5892,N_5499);
or U6293 (N_6293,N_5989,N_5906);
and U6294 (N_6294,N_5229,N_5425);
nor U6295 (N_6295,N_5610,N_5027);
xor U6296 (N_6296,N_5161,N_5066);
nor U6297 (N_6297,N_5378,N_5439);
and U6298 (N_6298,N_5009,N_5098);
or U6299 (N_6299,N_5381,N_4518);
xnor U6300 (N_6300,N_5348,N_4920);
nor U6301 (N_6301,N_4862,N_5053);
or U6302 (N_6302,N_5546,N_5124);
nor U6303 (N_6303,N_5507,N_5180);
and U6304 (N_6304,N_4598,N_5750);
nand U6305 (N_6305,N_5057,N_5844);
nor U6306 (N_6306,N_4961,N_5922);
and U6307 (N_6307,N_4597,N_5223);
or U6308 (N_6308,N_5561,N_5274);
nor U6309 (N_6309,N_5360,N_4564);
and U6310 (N_6310,N_5674,N_5442);
nand U6311 (N_6311,N_5418,N_4592);
and U6312 (N_6312,N_5685,N_4743);
xor U6313 (N_6313,N_5510,N_5611);
or U6314 (N_6314,N_5954,N_5601);
or U6315 (N_6315,N_4931,N_5283);
nor U6316 (N_6316,N_5205,N_4858);
or U6317 (N_6317,N_5752,N_5517);
or U6318 (N_6318,N_5000,N_4938);
nor U6319 (N_6319,N_5052,N_5614);
or U6320 (N_6320,N_4611,N_4536);
xor U6321 (N_6321,N_5926,N_4817);
or U6322 (N_6322,N_5653,N_5523);
nor U6323 (N_6323,N_4591,N_5664);
nand U6324 (N_6324,N_4982,N_5363);
or U6325 (N_6325,N_5355,N_4633);
and U6326 (N_6326,N_4529,N_5937);
nor U6327 (N_6327,N_4556,N_4688);
nand U6328 (N_6328,N_5380,N_4769);
xnor U6329 (N_6329,N_4955,N_5417);
nand U6330 (N_6330,N_5231,N_4587);
nand U6331 (N_6331,N_5805,N_5185);
nand U6332 (N_6332,N_5656,N_5138);
or U6333 (N_6333,N_5141,N_5708);
and U6334 (N_6334,N_4573,N_5530);
nor U6335 (N_6335,N_5722,N_5100);
and U6336 (N_6336,N_4574,N_4943);
and U6337 (N_6337,N_5456,N_5476);
and U6338 (N_6338,N_5903,N_5004);
nor U6339 (N_6339,N_5021,N_5999);
nor U6340 (N_6340,N_5093,N_5139);
nor U6341 (N_6341,N_5424,N_5804);
xnor U6342 (N_6342,N_4670,N_4975);
xor U6343 (N_6343,N_4846,N_5859);
xnor U6344 (N_6344,N_4879,N_5402);
or U6345 (N_6345,N_5475,N_4912);
nand U6346 (N_6346,N_4847,N_5993);
nor U6347 (N_6347,N_4836,N_4577);
nand U6348 (N_6348,N_4813,N_5545);
xor U6349 (N_6349,N_5145,N_4903);
nor U6350 (N_6350,N_4502,N_5465);
and U6351 (N_6351,N_4989,N_4727);
nor U6352 (N_6352,N_4919,N_5605);
or U6353 (N_6353,N_4767,N_4760);
nand U6354 (N_6354,N_5563,N_5727);
nor U6355 (N_6355,N_5930,N_5186);
xnor U6356 (N_6356,N_5482,N_5040);
or U6357 (N_6357,N_4650,N_5111);
nand U6358 (N_6358,N_5942,N_5232);
or U6359 (N_6359,N_5961,N_5622);
or U6360 (N_6360,N_4752,N_5237);
nor U6361 (N_6361,N_4992,N_4875);
nor U6362 (N_6362,N_4703,N_5468);
xor U6363 (N_6363,N_5342,N_5081);
and U6364 (N_6364,N_5144,N_5320);
xnor U6365 (N_6365,N_5016,N_4902);
nor U6366 (N_6366,N_5958,N_4856);
and U6367 (N_6367,N_5580,N_5170);
xnor U6368 (N_6368,N_5036,N_5133);
nor U6369 (N_6369,N_5716,N_5868);
nand U6370 (N_6370,N_4945,N_4572);
nand U6371 (N_6371,N_4734,N_5899);
nand U6372 (N_6372,N_5589,N_5444);
nand U6373 (N_6373,N_5834,N_4929);
xnor U6374 (N_6374,N_4554,N_4776);
or U6375 (N_6375,N_5284,N_4721);
nor U6376 (N_6376,N_4948,N_4906);
or U6377 (N_6377,N_4656,N_4979);
nor U6378 (N_6378,N_4787,N_4690);
and U6379 (N_6379,N_5840,N_5273);
or U6380 (N_6380,N_4531,N_5945);
or U6381 (N_6381,N_5008,N_5167);
or U6382 (N_6382,N_4876,N_5193);
nor U6383 (N_6383,N_5210,N_5203);
or U6384 (N_6384,N_4628,N_5815);
and U6385 (N_6385,N_5789,N_5778);
and U6386 (N_6386,N_4571,N_5695);
nand U6387 (N_6387,N_5154,N_4857);
and U6388 (N_6388,N_5964,N_5195);
nor U6389 (N_6389,N_5790,N_5090);
or U6390 (N_6390,N_5812,N_5616);
xor U6391 (N_6391,N_5249,N_5528);
or U6392 (N_6392,N_4784,N_5029);
nand U6393 (N_6393,N_5339,N_5041);
nand U6394 (N_6394,N_4723,N_5953);
nor U6395 (N_6395,N_5271,N_4606);
xnor U6396 (N_6396,N_4746,N_5896);
or U6397 (N_6397,N_5975,N_5085);
xor U6398 (N_6398,N_4801,N_5059);
nand U6399 (N_6399,N_5816,N_5222);
nand U6400 (N_6400,N_5742,N_4795);
or U6401 (N_6401,N_5092,N_4827);
xor U6402 (N_6402,N_4868,N_5699);
or U6403 (N_6403,N_4893,N_5257);
nor U6404 (N_6404,N_5174,N_5839);
nor U6405 (N_6405,N_5017,N_5502);
nor U6406 (N_6406,N_4545,N_5280);
nor U6407 (N_6407,N_5956,N_5712);
nand U6408 (N_6408,N_5295,N_5876);
nand U6409 (N_6409,N_4957,N_5891);
and U6410 (N_6410,N_4844,N_5303);
or U6411 (N_6411,N_4689,N_4641);
and U6412 (N_6412,N_5624,N_5198);
nand U6413 (N_6413,N_5709,N_4818);
and U6414 (N_6414,N_5694,N_5569);
nand U6415 (N_6415,N_5796,N_5733);
or U6416 (N_6416,N_5006,N_4675);
or U6417 (N_6417,N_5851,N_5288);
and U6418 (N_6418,N_4666,N_5632);
nand U6419 (N_6419,N_5640,N_5050);
or U6420 (N_6420,N_4678,N_5869);
or U6421 (N_6421,N_4834,N_5981);
nor U6422 (N_6422,N_4820,N_5723);
xnor U6423 (N_6423,N_4695,N_4659);
nand U6424 (N_6424,N_5191,N_5315);
or U6425 (N_6425,N_5970,N_5838);
nor U6426 (N_6426,N_5995,N_5178);
nand U6427 (N_6427,N_4824,N_5011);
or U6428 (N_6428,N_5058,N_4504);
xor U6429 (N_6429,N_5757,N_5885);
xnor U6430 (N_6430,N_4501,N_5870);
nor U6431 (N_6431,N_5806,N_4869);
nor U6432 (N_6432,N_4533,N_5369);
nand U6433 (N_6433,N_5524,N_5599);
xnor U6434 (N_6434,N_5984,N_5658);
nor U6435 (N_6435,N_5562,N_5304);
nand U6436 (N_6436,N_5933,N_4629);
nor U6437 (N_6437,N_5717,N_4973);
xor U6438 (N_6438,N_4777,N_5398);
and U6439 (N_6439,N_5415,N_5541);
nand U6440 (N_6440,N_5477,N_4977);
nand U6441 (N_6441,N_5690,N_4934);
or U6442 (N_6442,N_4937,N_4758);
nand U6443 (N_6443,N_5807,N_4774);
and U6444 (N_6444,N_5835,N_5698);
nand U6445 (N_6445,N_4704,N_4984);
nand U6446 (N_6446,N_5181,N_4878);
or U6447 (N_6447,N_5151,N_5641);
nand U6448 (N_6448,N_5786,N_5326);
nor U6449 (N_6449,N_5623,N_5076);
nand U6450 (N_6450,N_5781,N_5832);
or U6451 (N_6451,N_5276,N_4786);
xnor U6452 (N_6452,N_5446,N_4636);
and U6453 (N_6453,N_5117,N_4713);
nor U6454 (N_6454,N_4755,N_5341);
and U6455 (N_6455,N_5329,N_4842);
xor U6456 (N_6456,N_5522,N_5660);
or U6457 (N_6457,N_5405,N_4860);
and U6458 (N_6458,N_5979,N_4586);
xor U6459 (N_6459,N_5726,N_5671);
nand U6460 (N_6460,N_5130,N_4775);
nor U6461 (N_6461,N_4854,N_5131);
nand U6462 (N_6462,N_5002,N_5831);
or U6463 (N_6463,N_5741,N_4999);
xor U6464 (N_6464,N_5001,N_5334);
nand U6465 (N_6465,N_5940,N_5386);
or U6466 (N_6466,N_5099,N_5955);
and U6467 (N_6467,N_5112,N_5462);
nor U6468 (N_6468,N_5079,N_5095);
xor U6469 (N_6469,N_5787,N_5297);
nor U6470 (N_6470,N_4791,N_5531);
and U6471 (N_6471,N_5872,N_4543);
nor U6472 (N_6472,N_4783,N_5772);
and U6473 (N_6473,N_5571,N_4525);
and U6474 (N_6474,N_5207,N_5965);
nor U6475 (N_6475,N_5074,N_5388);
nor U6476 (N_6476,N_4625,N_4983);
and U6477 (N_6477,N_5966,N_5793);
xor U6478 (N_6478,N_5758,N_5212);
nor U6479 (N_6479,N_5263,N_5290);
nor U6480 (N_6480,N_5661,N_5201);
xnor U6481 (N_6481,N_5441,N_5492);
xor U6482 (N_6482,N_4789,N_5946);
and U6483 (N_6483,N_5557,N_4935);
or U6484 (N_6484,N_5060,N_5928);
and U6485 (N_6485,N_4810,N_5576);
nor U6486 (N_6486,N_5089,N_5670);
nand U6487 (N_6487,N_5014,N_4683);
xnor U6488 (N_6488,N_5917,N_5902);
nand U6489 (N_6489,N_4826,N_5447);
nor U6490 (N_6490,N_5416,N_5108);
and U6491 (N_6491,N_5678,N_5202);
xnor U6492 (N_6492,N_5509,N_5071);
and U6493 (N_6493,N_5810,N_5042);
nand U6494 (N_6494,N_5490,N_5555);
or U6495 (N_6495,N_4722,N_5982);
xnor U6496 (N_6496,N_4676,N_4840);
nor U6497 (N_6497,N_4993,N_4516);
and U6498 (N_6498,N_5950,N_5230);
nor U6499 (N_6499,N_4603,N_5407);
xor U6500 (N_6500,N_4725,N_5473);
and U6501 (N_6501,N_5146,N_5565);
and U6502 (N_6502,N_4588,N_5554);
nand U6503 (N_6503,N_5354,N_5795);
nor U6504 (N_6504,N_4616,N_5072);
or U6505 (N_6505,N_5791,N_5433);
or U6506 (N_6506,N_4673,N_5325);
and U6507 (N_6507,N_4745,N_5440);
xor U6508 (N_6508,N_5371,N_5880);
nand U6509 (N_6509,N_5078,N_4815);
nand U6510 (N_6510,N_5739,N_5628);
or U6511 (N_6511,N_4561,N_4532);
nand U6512 (N_6512,N_5314,N_5780);
nand U6513 (N_6513,N_5976,N_5598);
xor U6514 (N_6514,N_5255,N_5335);
nand U6515 (N_6515,N_4805,N_4927);
nand U6516 (N_6516,N_5751,N_5224);
nor U6517 (N_6517,N_4874,N_4940);
nor U6518 (N_6518,N_5638,N_5669);
nand U6519 (N_6519,N_4921,N_5766);
xor U6520 (N_6520,N_5067,N_4680);
or U6521 (N_6521,N_5564,N_5594);
nand U6522 (N_6522,N_4696,N_5422);
nor U6523 (N_6523,N_5376,N_5648);
nand U6524 (N_6524,N_4749,N_5218);
or U6525 (N_6525,N_5225,N_5745);
or U6526 (N_6526,N_4881,N_4915);
nand U6527 (N_6527,N_5403,N_5077);
or U6528 (N_6528,N_4534,N_5655);
nor U6529 (N_6529,N_4997,N_5762);
and U6530 (N_6530,N_5901,N_5625);
xnor U6531 (N_6531,N_5920,N_4972);
xnor U6532 (N_6532,N_4575,N_5083);
nor U6533 (N_6533,N_4685,N_5759);
nor U6534 (N_6534,N_5049,N_4884);
or U6535 (N_6535,N_5824,N_5848);
nand U6536 (N_6536,N_4552,N_5397);
and U6537 (N_6537,N_5361,N_5281);
and U6538 (N_6538,N_4674,N_5296);
and U6539 (N_6539,N_5721,N_5520);
xor U6540 (N_6540,N_4546,N_5533);
or U6541 (N_6541,N_5643,N_5877);
nand U6542 (N_6542,N_4899,N_4958);
or U6543 (N_6543,N_5370,N_5710);
and U6544 (N_6544,N_5291,N_5137);
xnor U6545 (N_6545,N_5148,N_5959);
and U6546 (N_6546,N_5607,N_5794);
nand U6547 (N_6547,N_5867,N_4630);
xnor U6548 (N_6548,N_5888,N_5411);
and U6549 (N_6549,N_4677,N_4952);
xnor U6550 (N_6550,N_5744,N_5667);
and U6551 (N_6551,N_4747,N_5672);
nand U6552 (N_6552,N_5969,N_4796);
nand U6553 (N_6553,N_4618,N_5467);
and U6554 (N_6554,N_5737,N_4622);
nand U6555 (N_6555,N_5663,N_4753);
nor U6556 (N_6556,N_4926,N_5241);
nor U6557 (N_6557,N_5821,N_5199);
nor U6558 (N_6558,N_5259,N_5725);
xor U6559 (N_6559,N_5884,N_4530);
or U6560 (N_6560,N_4936,N_5720);
nor U6561 (N_6561,N_4930,N_4520);
xnor U6562 (N_6562,N_5811,N_4687);
and U6563 (N_6563,N_5798,N_5034);
xnor U6564 (N_6564,N_4835,N_5713);
and U6565 (N_6565,N_4589,N_5512);
nor U6566 (N_6566,N_5412,N_5044);
and U6567 (N_6567,N_5633,N_5689);
or U6568 (N_6568,N_5075,N_5184);
and U6569 (N_6569,N_5890,N_5823);
xor U6570 (N_6570,N_5379,N_5550);
or U6571 (N_6571,N_4594,N_4764);
xor U6572 (N_6572,N_4942,N_4632);
nand U6573 (N_6573,N_5347,N_4839);
or U6574 (N_6574,N_4665,N_5115);
nor U6575 (N_6575,N_4863,N_5734);
and U6576 (N_6576,N_5849,N_4643);
and U6577 (N_6577,N_5164,N_5579);
nor U6578 (N_6578,N_4859,N_5627);
or U6579 (N_6579,N_5208,N_5219);
or U6580 (N_6580,N_4976,N_5927);
or U6581 (N_6581,N_5346,N_5264);
nand U6582 (N_6582,N_5887,N_5463);
nand U6583 (N_6583,N_4567,N_4809);
and U6584 (N_6584,N_4655,N_5192);
and U6585 (N_6585,N_5714,N_5367);
and U6586 (N_6586,N_5384,N_5577);
nand U6587 (N_6587,N_4887,N_4610);
and U6588 (N_6588,N_5833,N_5373);
nand U6589 (N_6589,N_4664,N_5974);
xnor U6590 (N_6590,N_5665,N_5070);
and U6591 (N_6591,N_5107,N_5506);
nor U6592 (N_6592,N_5846,N_4819);
and U6593 (N_6593,N_5220,N_5724);
or U6594 (N_6594,N_4646,N_5177);
nand U6595 (N_6595,N_5275,N_5503);
nor U6596 (N_6596,N_4925,N_4808);
or U6597 (N_6597,N_4731,N_4877);
or U6598 (N_6598,N_4691,N_4507);
nor U6599 (N_6599,N_5375,N_4947);
nand U6600 (N_6600,N_4733,N_5409);
and U6601 (N_6601,N_5228,N_4890);
and U6602 (N_6602,N_5730,N_4838);
nor U6603 (N_6603,N_5591,N_5583);
or U6604 (N_6604,N_5511,N_4684);
nand U6605 (N_6605,N_5612,N_5157);
nor U6606 (N_6606,N_5097,N_5478);
xor U6607 (N_6607,N_5155,N_5785);
nor U6608 (N_6608,N_5986,N_4602);
nor U6609 (N_6609,N_4706,N_5582);
nand U6610 (N_6610,N_5204,N_5932);
nand U6611 (N_6611,N_4660,N_5539);
and U6612 (N_6612,N_5702,N_4642);
nand U6613 (N_6613,N_5600,N_5803);
or U6614 (N_6614,N_5845,N_5236);
xor U6615 (N_6615,N_5194,N_5110);
xnor U6616 (N_6616,N_5827,N_4802);
and U6617 (N_6617,N_4963,N_5527);
nor U6618 (N_6618,N_4710,N_4793);
xor U6619 (N_6619,N_5457,N_4954);
and U6620 (N_6620,N_4698,N_5923);
nor U6621 (N_6621,N_4988,N_5596);
nor U6622 (N_6622,N_4799,N_5308);
xnor U6623 (N_6623,N_5278,N_5943);
nor U6624 (N_6624,N_5163,N_4512);
nand U6625 (N_6625,N_5990,N_5866);
or U6626 (N_6626,N_5039,N_5746);
and U6627 (N_6627,N_5736,N_4547);
or U6628 (N_6628,N_4668,N_4600);
xor U6629 (N_6629,N_5125,N_4953);
and U6630 (N_6630,N_4998,N_4772);
nand U6631 (N_6631,N_4667,N_5343);
nor U6632 (N_6632,N_5377,N_4996);
nand U6633 (N_6633,N_4918,N_5518);
or U6634 (N_6634,N_5106,N_5387);
nor U6635 (N_6635,N_5587,N_5592);
xor U6636 (N_6636,N_4576,N_4651);
or U6637 (N_6637,N_5673,N_4671);
xnor U6638 (N_6638,N_5556,N_5968);
or U6639 (N_6639,N_4771,N_5464);
xnor U6640 (N_6640,N_5261,N_5893);
or U6641 (N_6641,N_4613,N_5248);
and U6642 (N_6642,N_4708,N_5105);
xnor U6643 (N_6643,N_4566,N_5738);
or U6644 (N_6644,N_4653,N_5302);
xor U6645 (N_6645,N_5626,N_5534);
and U6646 (N_6646,N_5800,N_5064);
or U6647 (N_6647,N_4649,N_5395);
or U6648 (N_6648,N_5620,N_4946);
xor U6649 (N_6649,N_5128,N_5788);
or U6650 (N_6650,N_5349,N_5858);
and U6651 (N_6651,N_5873,N_4750);
xnor U6652 (N_6652,N_5031,N_5030);
xnor U6653 (N_6653,N_5350,N_5013);
and U6654 (N_6654,N_5919,N_5211);
nand U6655 (N_6655,N_5233,N_4794);
and U6656 (N_6656,N_5221,N_5015);
nand U6657 (N_6657,N_4885,N_5312);
nor U6658 (N_6658,N_4825,N_4757);
or U6659 (N_6659,N_4635,N_4624);
and U6660 (N_6660,N_5038,N_5634);
nand U6661 (N_6661,N_4716,N_5894);
or U6662 (N_6662,N_4923,N_5688);
and U6663 (N_6663,N_5693,N_4759);
xor U6664 (N_6664,N_5676,N_5235);
and U6665 (N_6665,N_5538,N_4640);
or U6666 (N_6666,N_4609,N_5324);
xnor U6667 (N_6667,N_4601,N_5486);
nand U6668 (N_6668,N_5217,N_5683);
xnor U6669 (N_6669,N_5536,N_5818);
nor U6670 (N_6670,N_5169,N_4908);
nor U6671 (N_6671,N_5570,N_5450);
nor U6672 (N_6672,N_5197,N_4615);
nor U6673 (N_6673,N_5748,N_5763);
xnor U6674 (N_6674,N_5586,N_4913);
xnor U6675 (N_6675,N_4527,N_5400);
or U6676 (N_6676,N_4822,N_5609);
or U6677 (N_6677,N_5829,N_5949);
and U6678 (N_6678,N_5568,N_4557);
nand U6679 (N_6679,N_5645,N_5897);
xor U6680 (N_6680,N_5590,N_4595);
xnor U6681 (N_6681,N_5875,N_5519);
and U6682 (N_6682,N_5558,N_5429);
and U6683 (N_6683,N_4620,N_4761);
or U6684 (N_6684,N_5547,N_5992);
or U6685 (N_6685,N_4661,N_5340);
nor U6686 (N_6686,N_5003,N_5176);
or U6687 (N_6687,N_5662,N_4679);
or U6688 (N_6688,N_5035,N_4644);
nand U6689 (N_6689,N_5650,N_5879);
nor U6690 (N_6690,N_4811,N_5307);
or U6691 (N_6691,N_5451,N_5886);
xnor U6692 (N_6692,N_4631,N_5874);
and U6693 (N_6693,N_5947,N_5941);
xor U6694 (N_6694,N_5701,N_5345);
xor U6695 (N_6695,N_5825,N_4956);
nand U6696 (N_6696,N_5910,N_4515);
and U6697 (N_6697,N_4871,N_4788);
or U6698 (N_6698,N_5644,N_5452);
xnor U6699 (N_6699,N_4583,N_5754);
or U6700 (N_6700,N_5200,N_5366);
xnor U6701 (N_6701,N_5426,N_4765);
nand U6702 (N_6702,N_5779,N_5649);
nor U6703 (N_6703,N_5420,N_5508);
and U6704 (N_6704,N_5882,N_5453);
and U6705 (N_6705,N_5918,N_5998);
or U6706 (N_6706,N_5826,N_4744);
or U6707 (N_6707,N_5364,N_4922);
nand U6708 (N_6708,N_5572,N_4837);
nor U6709 (N_6709,N_5359,N_4619);
nor U6710 (N_6710,N_5080,N_5760);
xor U6711 (N_6711,N_4705,N_5813);
nor U6712 (N_6712,N_5784,N_4697);
nand U6713 (N_6713,N_5907,N_4521);
xor U6714 (N_6714,N_5129,N_4960);
nor U6715 (N_6715,N_4980,N_5862);
and U6716 (N_6716,N_4782,N_4924);
and U6717 (N_6717,N_4669,N_5171);
and U6718 (N_6718,N_4756,N_4693);
or U6719 (N_6719,N_4949,N_5944);
nand U6720 (N_6720,N_5621,N_5268);
nor U6721 (N_6721,N_4951,N_5635);
nor U6722 (N_6722,N_4891,N_5368);
nand U6723 (N_6723,N_5406,N_5445);
or U6724 (N_6724,N_4916,N_5183);
nor U6725 (N_6725,N_5792,N_4663);
and U6726 (N_6726,N_5322,N_4579);
or U6727 (N_6727,N_5505,N_4852);
and U6728 (N_6728,N_5544,N_4654);
or U6729 (N_6729,N_4526,N_5443);
nor U6730 (N_6730,N_5158,N_4626);
nor U6731 (N_6731,N_5603,N_4555);
or U6732 (N_6732,N_5269,N_4962);
or U6733 (N_6733,N_5797,N_4831);
nor U6734 (N_6734,N_5863,N_5047);
and U6735 (N_6735,N_5054,N_5010);
and U6736 (N_6736,N_5735,N_5175);
or U6737 (N_6737,N_5495,N_5978);
or U6738 (N_6738,N_5298,N_4686);
xor U6739 (N_6739,N_5585,N_5134);
nor U6740 (N_6740,N_5747,N_4657);
xor U6741 (N_6741,N_4562,N_5051);
nand U6742 (N_6742,N_5783,N_4513);
nand U6743 (N_6743,N_5460,N_4832);
nor U6744 (N_6744,N_5331,N_4658);
or U6745 (N_6745,N_5684,N_4966);
or U6746 (N_6746,N_4865,N_5481);
and U6747 (N_6747,N_5977,N_5852);
or U6748 (N_6748,N_4768,N_5567);
nor U6749 (N_6749,N_5023,N_5305);
and U6750 (N_6750,N_5969,N_5772);
xor U6751 (N_6751,N_5832,N_5658);
and U6752 (N_6752,N_5900,N_4639);
xor U6753 (N_6753,N_4957,N_5544);
and U6754 (N_6754,N_4561,N_5474);
xnor U6755 (N_6755,N_5046,N_4937);
or U6756 (N_6756,N_4621,N_4912);
and U6757 (N_6757,N_5793,N_4873);
nor U6758 (N_6758,N_5558,N_4624);
and U6759 (N_6759,N_4750,N_5653);
and U6760 (N_6760,N_5352,N_5255);
xor U6761 (N_6761,N_4909,N_4785);
nor U6762 (N_6762,N_5329,N_5099);
or U6763 (N_6763,N_5893,N_5500);
nor U6764 (N_6764,N_5611,N_4675);
nor U6765 (N_6765,N_4652,N_4759);
or U6766 (N_6766,N_5448,N_5097);
nand U6767 (N_6767,N_5132,N_5331);
nor U6768 (N_6768,N_4801,N_5964);
nand U6769 (N_6769,N_5143,N_4656);
and U6770 (N_6770,N_5149,N_5665);
xor U6771 (N_6771,N_4574,N_5270);
nor U6772 (N_6772,N_4799,N_4815);
and U6773 (N_6773,N_5105,N_5277);
nor U6774 (N_6774,N_5187,N_4603);
nand U6775 (N_6775,N_4929,N_4722);
nand U6776 (N_6776,N_4716,N_4966);
xnor U6777 (N_6777,N_5263,N_5059);
or U6778 (N_6778,N_4667,N_5714);
nand U6779 (N_6779,N_5899,N_4784);
xor U6780 (N_6780,N_4797,N_5880);
nand U6781 (N_6781,N_5488,N_5331);
xor U6782 (N_6782,N_5492,N_4800);
nand U6783 (N_6783,N_5643,N_5958);
nor U6784 (N_6784,N_5622,N_4822);
or U6785 (N_6785,N_5977,N_5342);
or U6786 (N_6786,N_5675,N_5762);
or U6787 (N_6787,N_4518,N_5467);
nor U6788 (N_6788,N_5781,N_5675);
nand U6789 (N_6789,N_5265,N_4505);
nor U6790 (N_6790,N_5421,N_4523);
nand U6791 (N_6791,N_5590,N_4644);
xnor U6792 (N_6792,N_5432,N_5311);
and U6793 (N_6793,N_5908,N_5805);
nor U6794 (N_6794,N_5910,N_5592);
xnor U6795 (N_6795,N_5557,N_4707);
xnor U6796 (N_6796,N_4830,N_5183);
nor U6797 (N_6797,N_4876,N_5316);
and U6798 (N_6798,N_5692,N_4930);
nor U6799 (N_6799,N_5240,N_5096);
nor U6800 (N_6800,N_5383,N_5830);
and U6801 (N_6801,N_5584,N_5518);
nand U6802 (N_6802,N_4965,N_4767);
nor U6803 (N_6803,N_5937,N_5610);
and U6804 (N_6804,N_4673,N_5106);
and U6805 (N_6805,N_5665,N_5886);
or U6806 (N_6806,N_5938,N_5196);
or U6807 (N_6807,N_5964,N_5776);
nor U6808 (N_6808,N_5501,N_4789);
nand U6809 (N_6809,N_5532,N_5813);
or U6810 (N_6810,N_5920,N_5403);
nand U6811 (N_6811,N_4961,N_4594);
and U6812 (N_6812,N_5673,N_5556);
and U6813 (N_6813,N_5311,N_5970);
xor U6814 (N_6814,N_4943,N_4572);
nand U6815 (N_6815,N_5226,N_5046);
or U6816 (N_6816,N_5734,N_4749);
nor U6817 (N_6817,N_5714,N_4892);
xnor U6818 (N_6818,N_5738,N_4764);
nand U6819 (N_6819,N_4898,N_4871);
nor U6820 (N_6820,N_5630,N_4778);
nor U6821 (N_6821,N_4834,N_5075);
nand U6822 (N_6822,N_4681,N_5664);
xnor U6823 (N_6823,N_4552,N_5391);
xor U6824 (N_6824,N_5274,N_5336);
and U6825 (N_6825,N_5491,N_4877);
nor U6826 (N_6826,N_4655,N_5296);
nand U6827 (N_6827,N_4729,N_4859);
xnor U6828 (N_6828,N_5558,N_5939);
nor U6829 (N_6829,N_5301,N_4573);
xnor U6830 (N_6830,N_4779,N_4751);
nor U6831 (N_6831,N_5560,N_4540);
or U6832 (N_6832,N_4701,N_5016);
nor U6833 (N_6833,N_4806,N_4783);
nand U6834 (N_6834,N_5100,N_4929);
and U6835 (N_6835,N_4539,N_5095);
and U6836 (N_6836,N_5791,N_5364);
or U6837 (N_6837,N_5276,N_5267);
xor U6838 (N_6838,N_5917,N_5048);
or U6839 (N_6839,N_5670,N_5986);
nor U6840 (N_6840,N_5987,N_5406);
xnor U6841 (N_6841,N_5324,N_5857);
and U6842 (N_6842,N_4987,N_5416);
xnor U6843 (N_6843,N_4666,N_5485);
xnor U6844 (N_6844,N_5920,N_5076);
nor U6845 (N_6845,N_5785,N_5512);
and U6846 (N_6846,N_4881,N_4739);
nand U6847 (N_6847,N_5325,N_4873);
or U6848 (N_6848,N_5991,N_4945);
xor U6849 (N_6849,N_4909,N_5086);
or U6850 (N_6850,N_4873,N_5216);
or U6851 (N_6851,N_4626,N_5314);
nor U6852 (N_6852,N_5343,N_4746);
or U6853 (N_6853,N_4677,N_4894);
nor U6854 (N_6854,N_4775,N_4695);
nand U6855 (N_6855,N_5736,N_5806);
nor U6856 (N_6856,N_5282,N_5523);
or U6857 (N_6857,N_5417,N_5033);
or U6858 (N_6858,N_5332,N_5567);
nor U6859 (N_6859,N_5838,N_5939);
xnor U6860 (N_6860,N_5189,N_5448);
or U6861 (N_6861,N_4664,N_5681);
and U6862 (N_6862,N_4959,N_5368);
or U6863 (N_6863,N_5296,N_4820);
xor U6864 (N_6864,N_4575,N_4846);
xnor U6865 (N_6865,N_5197,N_5587);
nor U6866 (N_6866,N_4611,N_5436);
nand U6867 (N_6867,N_5142,N_4985);
and U6868 (N_6868,N_5752,N_4613);
nor U6869 (N_6869,N_5808,N_5275);
nor U6870 (N_6870,N_5768,N_5797);
nand U6871 (N_6871,N_5299,N_4872);
nor U6872 (N_6872,N_5913,N_4578);
xnor U6873 (N_6873,N_5486,N_5964);
nor U6874 (N_6874,N_4822,N_5527);
or U6875 (N_6875,N_5542,N_4805);
and U6876 (N_6876,N_5155,N_4701);
nand U6877 (N_6877,N_5711,N_5332);
nor U6878 (N_6878,N_4793,N_5218);
xnor U6879 (N_6879,N_4994,N_5707);
or U6880 (N_6880,N_4659,N_5248);
xnor U6881 (N_6881,N_5745,N_5090);
xor U6882 (N_6882,N_4645,N_5346);
nand U6883 (N_6883,N_5978,N_5479);
or U6884 (N_6884,N_5952,N_5146);
xnor U6885 (N_6885,N_5019,N_4969);
and U6886 (N_6886,N_5789,N_4503);
nand U6887 (N_6887,N_4945,N_4941);
or U6888 (N_6888,N_5869,N_5123);
and U6889 (N_6889,N_5566,N_5514);
xor U6890 (N_6890,N_5734,N_5355);
and U6891 (N_6891,N_4919,N_5009);
or U6892 (N_6892,N_5620,N_4781);
and U6893 (N_6893,N_5607,N_5498);
xnor U6894 (N_6894,N_5373,N_5059);
nor U6895 (N_6895,N_5066,N_5022);
xor U6896 (N_6896,N_5495,N_4835);
and U6897 (N_6897,N_5093,N_5408);
and U6898 (N_6898,N_5178,N_5392);
nand U6899 (N_6899,N_4786,N_5814);
xor U6900 (N_6900,N_5604,N_4563);
or U6901 (N_6901,N_5577,N_5556);
or U6902 (N_6902,N_5772,N_5824);
and U6903 (N_6903,N_4553,N_4515);
nor U6904 (N_6904,N_5032,N_5989);
nand U6905 (N_6905,N_4556,N_4872);
xnor U6906 (N_6906,N_5244,N_4658);
xnor U6907 (N_6907,N_4777,N_4708);
and U6908 (N_6908,N_4614,N_4720);
nand U6909 (N_6909,N_4949,N_5633);
xor U6910 (N_6910,N_5553,N_5208);
or U6911 (N_6911,N_4757,N_5175);
nor U6912 (N_6912,N_5803,N_5739);
or U6913 (N_6913,N_5546,N_5002);
and U6914 (N_6914,N_4779,N_5159);
nor U6915 (N_6915,N_4500,N_5723);
nor U6916 (N_6916,N_5511,N_4664);
nand U6917 (N_6917,N_5258,N_4877);
and U6918 (N_6918,N_4571,N_5323);
and U6919 (N_6919,N_5679,N_4910);
nor U6920 (N_6920,N_5052,N_5968);
and U6921 (N_6921,N_4605,N_4601);
nand U6922 (N_6922,N_5571,N_4936);
nand U6923 (N_6923,N_5999,N_5982);
nor U6924 (N_6924,N_5188,N_5893);
xnor U6925 (N_6925,N_5787,N_4553);
nand U6926 (N_6926,N_4902,N_5756);
and U6927 (N_6927,N_5727,N_5652);
and U6928 (N_6928,N_5141,N_5466);
or U6929 (N_6929,N_5505,N_4962);
or U6930 (N_6930,N_5677,N_5151);
and U6931 (N_6931,N_5951,N_5675);
and U6932 (N_6932,N_5572,N_5692);
xor U6933 (N_6933,N_5919,N_5504);
xnor U6934 (N_6934,N_5312,N_5098);
or U6935 (N_6935,N_4573,N_5208);
nand U6936 (N_6936,N_5080,N_4934);
nand U6937 (N_6937,N_5744,N_5211);
xnor U6938 (N_6938,N_5350,N_5653);
and U6939 (N_6939,N_5563,N_4849);
and U6940 (N_6940,N_5420,N_5626);
nand U6941 (N_6941,N_5556,N_5700);
or U6942 (N_6942,N_5381,N_4723);
or U6943 (N_6943,N_4877,N_5148);
nor U6944 (N_6944,N_5757,N_4634);
xnor U6945 (N_6945,N_5714,N_4835);
nor U6946 (N_6946,N_5792,N_4676);
xor U6947 (N_6947,N_5116,N_5520);
and U6948 (N_6948,N_5833,N_5477);
and U6949 (N_6949,N_5898,N_4638);
and U6950 (N_6950,N_5316,N_5118);
or U6951 (N_6951,N_5634,N_5270);
nand U6952 (N_6952,N_4831,N_5051);
or U6953 (N_6953,N_5712,N_5313);
or U6954 (N_6954,N_5073,N_5427);
xnor U6955 (N_6955,N_4748,N_5009);
nand U6956 (N_6956,N_5606,N_4501);
nor U6957 (N_6957,N_5607,N_4971);
nand U6958 (N_6958,N_5361,N_4918);
xor U6959 (N_6959,N_4957,N_4998);
nor U6960 (N_6960,N_5299,N_4512);
xnor U6961 (N_6961,N_5551,N_5654);
nor U6962 (N_6962,N_5125,N_4503);
xnor U6963 (N_6963,N_4890,N_5369);
nor U6964 (N_6964,N_5858,N_5941);
or U6965 (N_6965,N_5732,N_5252);
nor U6966 (N_6966,N_4763,N_5578);
and U6967 (N_6967,N_5131,N_4963);
xnor U6968 (N_6968,N_5417,N_4866);
nor U6969 (N_6969,N_5948,N_5412);
or U6970 (N_6970,N_4573,N_5654);
xnor U6971 (N_6971,N_4795,N_4678);
xor U6972 (N_6972,N_4529,N_5176);
nor U6973 (N_6973,N_4580,N_4911);
and U6974 (N_6974,N_5035,N_5518);
xor U6975 (N_6975,N_5988,N_5563);
xor U6976 (N_6976,N_4915,N_5357);
or U6977 (N_6977,N_5098,N_5336);
nor U6978 (N_6978,N_4590,N_5649);
nor U6979 (N_6979,N_5596,N_5486);
or U6980 (N_6980,N_4883,N_5467);
nand U6981 (N_6981,N_5591,N_5522);
xnor U6982 (N_6982,N_5466,N_4669);
or U6983 (N_6983,N_5074,N_5097);
xor U6984 (N_6984,N_4698,N_5860);
nand U6985 (N_6985,N_4821,N_5489);
nand U6986 (N_6986,N_5001,N_4621);
or U6987 (N_6987,N_5426,N_5730);
nand U6988 (N_6988,N_5914,N_5491);
and U6989 (N_6989,N_5727,N_5379);
nand U6990 (N_6990,N_4845,N_4505);
or U6991 (N_6991,N_4707,N_4699);
xnor U6992 (N_6992,N_4599,N_5756);
or U6993 (N_6993,N_5433,N_4566);
and U6994 (N_6994,N_5038,N_5426);
and U6995 (N_6995,N_4520,N_4686);
xnor U6996 (N_6996,N_5374,N_4719);
nor U6997 (N_6997,N_5973,N_5180);
nor U6998 (N_6998,N_5728,N_5955);
and U6999 (N_6999,N_5348,N_4582);
nand U7000 (N_7000,N_5701,N_5487);
or U7001 (N_7001,N_5350,N_4691);
nor U7002 (N_7002,N_5284,N_4895);
nand U7003 (N_7003,N_5010,N_5521);
and U7004 (N_7004,N_5061,N_5824);
and U7005 (N_7005,N_5955,N_5960);
and U7006 (N_7006,N_5958,N_5288);
xor U7007 (N_7007,N_5727,N_4737);
xnor U7008 (N_7008,N_4535,N_5515);
nand U7009 (N_7009,N_4752,N_5301);
and U7010 (N_7010,N_4800,N_5736);
nand U7011 (N_7011,N_5789,N_5494);
or U7012 (N_7012,N_4894,N_4853);
and U7013 (N_7013,N_4598,N_4698);
and U7014 (N_7014,N_4923,N_4697);
xor U7015 (N_7015,N_4844,N_4867);
nor U7016 (N_7016,N_5760,N_5146);
xor U7017 (N_7017,N_5627,N_4850);
nand U7018 (N_7018,N_5077,N_4775);
or U7019 (N_7019,N_5117,N_5307);
nand U7020 (N_7020,N_4939,N_5401);
or U7021 (N_7021,N_5501,N_4515);
and U7022 (N_7022,N_5677,N_5810);
nor U7023 (N_7023,N_5538,N_5106);
xor U7024 (N_7024,N_4741,N_4586);
and U7025 (N_7025,N_5785,N_4722);
and U7026 (N_7026,N_5738,N_5314);
nor U7027 (N_7027,N_5465,N_5173);
and U7028 (N_7028,N_5872,N_5863);
and U7029 (N_7029,N_5391,N_5581);
and U7030 (N_7030,N_4875,N_5213);
or U7031 (N_7031,N_4959,N_5227);
nor U7032 (N_7032,N_4916,N_4501);
nand U7033 (N_7033,N_5715,N_5799);
nand U7034 (N_7034,N_5868,N_4545);
xor U7035 (N_7035,N_4952,N_5064);
or U7036 (N_7036,N_4826,N_5535);
xor U7037 (N_7037,N_5706,N_4942);
xor U7038 (N_7038,N_4556,N_4640);
nand U7039 (N_7039,N_5183,N_5425);
xor U7040 (N_7040,N_5421,N_5868);
or U7041 (N_7041,N_5747,N_4637);
and U7042 (N_7042,N_4995,N_5943);
nor U7043 (N_7043,N_5499,N_5856);
or U7044 (N_7044,N_4749,N_4748);
xnor U7045 (N_7045,N_5086,N_5119);
or U7046 (N_7046,N_5530,N_5471);
xor U7047 (N_7047,N_5908,N_5616);
nand U7048 (N_7048,N_5087,N_5533);
nor U7049 (N_7049,N_5177,N_5189);
nand U7050 (N_7050,N_5715,N_4920);
and U7051 (N_7051,N_5193,N_5650);
or U7052 (N_7052,N_5230,N_4602);
xnor U7053 (N_7053,N_5613,N_5165);
nand U7054 (N_7054,N_4915,N_5479);
nand U7055 (N_7055,N_4843,N_5296);
nor U7056 (N_7056,N_5337,N_5478);
and U7057 (N_7057,N_4904,N_5045);
or U7058 (N_7058,N_4574,N_5052);
xor U7059 (N_7059,N_5914,N_5721);
and U7060 (N_7060,N_5639,N_4690);
and U7061 (N_7061,N_5103,N_4730);
and U7062 (N_7062,N_5880,N_5698);
nor U7063 (N_7063,N_5558,N_5336);
and U7064 (N_7064,N_4979,N_4574);
xor U7065 (N_7065,N_5545,N_5029);
nor U7066 (N_7066,N_5809,N_5522);
xor U7067 (N_7067,N_5257,N_5600);
nand U7068 (N_7068,N_5502,N_5259);
or U7069 (N_7069,N_5558,N_4641);
nand U7070 (N_7070,N_5531,N_4516);
and U7071 (N_7071,N_5516,N_5230);
nand U7072 (N_7072,N_5213,N_5432);
nand U7073 (N_7073,N_5022,N_5794);
nand U7074 (N_7074,N_5144,N_5250);
xor U7075 (N_7075,N_4503,N_5972);
and U7076 (N_7076,N_5010,N_5277);
and U7077 (N_7077,N_5192,N_5405);
nand U7078 (N_7078,N_4551,N_5838);
and U7079 (N_7079,N_5566,N_5540);
nor U7080 (N_7080,N_5973,N_5446);
nor U7081 (N_7081,N_5270,N_4962);
and U7082 (N_7082,N_5287,N_5259);
nand U7083 (N_7083,N_5922,N_4949);
nor U7084 (N_7084,N_5645,N_5409);
or U7085 (N_7085,N_5067,N_5903);
or U7086 (N_7086,N_5255,N_5775);
nand U7087 (N_7087,N_4828,N_5875);
xnor U7088 (N_7088,N_5210,N_5209);
nand U7089 (N_7089,N_4881,N_5969);
nor U7090 (N_7090,N_5875,N_5931);
or U7091 (N_7091,N_4883,N_5021);
or U7092 (N_7092,N_5540,N_5965);
nand U7093 (N_7093,N_5878,N_5378);
nor U7094 (N_7094,N_4828,N_5262);
nand U7095 (N_7095,N_5867,N_5271);
nand U7096 (N_7096,N_5897,N_4719);
or U7097 (N_7097,N_5688,N_5609);
nand U7098 (N_7098,N_4643,N_5749);
xnor U7099 (N_7099,N_4602,N_5001);
nand U7100 (N_7100,N_4577,N_5532);
xnor U7101 (N_7101,N_5498,N_5936);
xor U7102 (N_7102,N_5098,N_5170);
nor U7103 (N_7103,N_5520,N_4667);
xnor U7104 (N_7104,N_5270,N_4585);
or U7105 (N_7105,N_5603,N_4888);
xor U7106 (N_7106,N_5306,N_4671);
and U7107 (N_7107,N_4716,N_5461);
and U7108 (N_7108,N_4849,N_4704);
nand U7109 (N_7109,N_5696,N_4990);
nand U7110 (N_7110,N_4896,N_5846);
xnor U7111 (N_7111,N_4731,N_5779);
nor U7112 (N_7112,N_5268,N_4613);
nand U7113 (N_7113,N_5910,N_5395);
xnor U7114 (N_7114,N_5321,N_5994);
xnor U7115 (N_7115,N_5269,N_5894);
xnor U7116 (N_7116,N_5609,N_5361);
xnor U7117 (N_7117,N_4846,N_4567);
and U7118 (N_7118,N_4907,N_5828);
nor U7119 (N_7119,N_4850,N_5068);
and U7120 (N_7120,N_5511,N_4709);
nor U7121 (N_7121,N_4894,N_5378);
nor U7122 (N_7122,N_5269,N_4880);
xnor U7123 (N_7123,N_4750,N_5603);
nand U7124 (N_7124,N_4971,N_5949);
nor U7125 (N_7125,N_4953,N_5241);
or U7126 (N_7126,N_5335,N_4778);
xor U7127 (N_7127,N_5121,N_4817);
xnor U7128 (N_7128,N_5423,N_4830);
nor U7129 (N_7129,N_5332,N_5480);
xnor U7130 (N_7130,N_5375,N_5208);
or U7131 (N_7131,N_5799,N_5348);
and U7132 (N_7132,N_5041,N_5026);
and U7133 (N_7133,N_4936,N_4807);
xnor U7134 (N_7134,N_5015,N_5500);
nand U7135 (N_7135,N_4638,N_5857);
and U7136 (N_7136,N_4947,N_5863);
and U7137 (N_7137,N_5619,N_4704);
and U7138 (N_7138,N_5017,N_5482);
nand U7139 (N_7139,N_5520,N_5955);
xor U7140 (N_7140,N_4683,N_5648);
nand U7141 (N_7141,N_5480,N_4696);
nor U7142 (N_7142,N_4750,N_5270);
nand U7143 (N_7143,N_4982,N_5754);
and U7144 (N_7144,N_4854,N_5733);
nor U7145 (N_7145,N_4667,N_5988);
or U7146 (N_7146,N_5291,N_4731);
and U7147 (N_7147,N_5822,N_4881);
nor U7148 (N_7148,N_5276,N_5205);
and U7149 (N_7149,N_5008,N_4605);
nand U7150 (N_7150,N_5673,N_5535);
nor U7151 (N_7151,N_4985,N_5352);
nor U7152 (N_7152,N_5965,N_5416);
nor U7153 (N_7153,N_5077,N_5569);
or U7154 (N_7154,N_4542,N_5335);
nor U7155 (N_7155,N_5519,N_5554);
xor U7156 (N_7156,N_5432,N_4575);
nor U7157 (N_7157,N_4513,N_5449);
or U7158 (N_7158,N_4656,N_5641);
nand U7159 (N_7159,N_4594,N_5005);
and U7160 (N_7160,N_5688,N_4766);
and U7161 (N_7161,N_4732,N_5158);
xor U7162 (N_7162,N_5709,N_5447);
or U7163 (N_7163,N_5752,N_5280);
xnor U7164 (N_7164,N_5155,N_5363);
or U7165 (N_7165,N_4862,N_4504);
and U7166 (N_7166,N_5645,N_5943);
or U7167 (N_7167,N_5923,N_5656);
nand U7168 (N_7168,N_5598,N_5047);
or U7169 (N_7169,N_4526,N_5257);
or U7170 (N_7170,N_5304,N_4575);
or U7171 (N_7171,N_5473,N_5780);
nand U7172 (N_7172,N_5665,N_5112);
nor U7173 (N_7173,N_5789,N_5908);
or U7174 (N_7174,N_5333,N_5523);
nor U7175 (N_7175,N_4592,N_5763);
nor U7176 (N_7176,N_5288,N_5959);
xnor U7177 (N_7177,N_4725,N_5403);
and U7178 (N_7178,N_5905,N_5082);
xor U7179 (N_7179,N_4847,N_4988);
xor U7180 (N_7180,N_4849,N_5502);
nor U7181 (N_7181,N_5464,N_5747);
and U7182 (N_7182,N_4563,N_5330);
or U7183 (N_7183,N_4600,N_4669);
or U7184 (N_7184,N_5376,N_4819);
nand U7185 (N_7185,N_5034,N_4972);
and U7186 (N_7186,N_4747,N_5727);
or U7187 (N_7187,N_4837,N_5018);
and U7188 (N_7188,N_5401,N_4605);
nor U7189 (N_7189,N_5240,N_5824);
nand U7190 (N_7190,N_4755,N_5854);
or U7191 (N_7191,N_4973,N_5572);
or U7192 (N_7192,N_5389,N_5756);
nor U7193 (N_7193,N_5758,N_5683);
and U7194 (N_7194,N_4977,N_4856);
xor U7195 (N_7195,N_5416,N_5076);
nor U7196 (N_7196,N_4800,N_5733);
nand U7197 (N_7197,N_5578,N_4536);
nand U7198 (N_7198,N_5197,N_5109);
nand U7199 (N_7199,N_5718,N_4999);
xnor U7200 (N_7200,N_4891,N_5177);
nor U7201 (N_7201,N_5846,N_4669);
xor U7202 (N_7202,N_4653,N_4799);
xnor U7203 (N_7203,N_4680,N_4627);
nand U7204 (N_7204,N_5196,N_5551);
or U7205 (N_7205,N_4586,N_5290);
xor U7206 (N_7206,N_5669,N_5198);
or U7207 (N_7207,N_4541,N_5649);
or U7208 (N_7208,N_4874,N_5585);
and U7209 (N_7209,N_4989,N_5317);
xor U7210 (N_7210,N_5058,N_5479);
nor U7211 (N_7211,N_5856,N_4845);
xor U7212 (N_7212,N_5853,N_5898);
xor U7213 (N_7213,N_4882,N_5911);
xnor U7214 (N_7214,N_5907,N_5241);
xnor U7215 (N_7215,N_4717,N_5619);
xnor U7216 (N_7216,N_5716,N_4677);
nand U7217 (N_7217,N_4985,N_4531);
xnor U7218 (N_7218,N_5802,N_5673);
nor U7219 (N_7219,N_5017,N_4581);
or U7220 (N_7220,N_4989,N_5468);
nand U7221 (N_7221,N_5954,N_5054);
nor U7222 (N_7222,N_5320,N_4622);
and U7223 (N_7223,N_5093,N_5430);
and U7224 (N_7224,N_5598,N_5403);
xor U7225 (N_7225,N_5188,N_4617);
and U7226 (N_7226,N_5212,N_4991);
or U7227 (N_7227,N_5201,N_5927);
and U7228 (N_7228,N_5808,N_4552);
and U7229 (N_7229,N_4934,N_5836);
nor U7230 (N_7230,N_5504,N_4614);
xor U7231 (N_7231,N_5232,N_4680);
or U7232 (N_7232,N_5259,N_5423);
xor U7233 (N_7233,N_5906,N_5736);
xnor U7234 (N_7234,N_5446,N_4552);
and U7235 (N_7235,N_5289,N_5978);
or U7236 (N_7236,N_5206,N_5669);
and U7237 (N_7237,N_5103,N_5555);
nor U7238 (N_7238,N_4584,N_4907);
or U7239 (N_7239,N_4765,N_5390);
and U7240 (N_7240,N_5772,N_4568);
nor U7241 (N_7241,N_4674,N_5259);
nand U7242 (N_7242,N_4994,N_5956);
and U7243 (N_7243,N_4557,N_4963);
xnor U7244 (N_7244,N_4613,N_5762);
or U7245 (N_7245,N_5281,N_5772);
and U7246 (N_7246,N_5896,N_5497);
or U7247 (N_7247,N_4719,N_4723);
nand U7248 (N_7248,N_5204,N_4721);
or U7249 (N_7249,N_4927,N_5611);
nand U7250 (N_7250,N_5978,N_5268);
or U7251 (N_7251,N_5545,N_5997);
nor U7252 (N_7252,N_4657,N_4832);
and U7253 (N_7253,N_4668,N_5029);
nand U7254 (N_7254,N_5361,N_5555);
xnor U7255 (N_7255,N_5891,N_5846);
nor U7256 (N_7256,N_4745,N_5443);
xnor U7257 (N_7257,N_4936,N_5439);
and U7258 (N_7258,N_5275,N_5814);
and U7259 (N_7259,N_4630,N_5518);
or U7260 (N_7260,N_4554,N_4501);
xnor U7261 (N_7261,N_5411,N_5487);
or U7262 (N_7262,N_5678,N_4552);
xnor U7263 (N_7263,N_5361,N_4741);
and U7264 (N_7264,N_5833,N_4919);
and U7265 (N_7265,N_5504,N_5507);
and U7266 (N_7266,N_4684,N_4590);
or U7267 (N_7267,N_5421,N_5005);
or U7268 (N_7268,N_4644,N_4967);
nand U7269 (N_7269,N_4713,N_5996);
xnor U7270 (N_7270,N_5248,N_5417);
nor U7271 (N_7271,N_4712,N_5448);
xnor U7272 (N_7272,N_4727,N_5797);
xor U7273 (N_7273,N_5617,N_5864);
and U7274 (N_7274,N_5694,N_5787);
xnor U7275 (N_7275,N_4705,N_5247);
or U7276 (N_7276,N_4995,N_4557);
nand U7277 (N_7277,N_4691,N_5388);
nand U7278 (N_7278,N_5143,N_5693);
nor U7279 (N_7279,N_5032,N_5169);
and U7280 (N_7280,N_4702,N_4876);
nor U7281 (N_7281,N_5558,N_5400);
nand U7282 (N_7282,N_4927,N_5342);
or U7283 (N_7283,N_4888,N_5243);
or U7284 (N_7284,N_5718,N_5103);
and U7285 (N_7285,N_5287,N_5342);
and U7286 (N_7286,N_5972,N_5961);
nor U7287 (N_7287,N_5235,N_4956);
nor U7288 (N_7288,N_4664,N_4813);
and U7289 (N_7289,N_4638,N_4867);
nor U7290 (N_7290,N_5111,N_5452);
nor U7291 (N_7291,N_5880,N_5884);
or U7292 (N_7292,N_4761,N_5170);
nor U7293 (N_7293,N_5641,N_5934);
and U7294 (N_7294,N_4661,N_4810);
or U7295 (N_7295,N_4598,N_4643);
nand U7296 (N_7296,N_5700,N_5838);
and U7297 (N_7297,N_5104,N_5876);
xnor U7298 (N_7298,N_5947,N_5027);
xnor U7299 (N_7299,N_4536,N_4711);
nand U7300 (N_7300,N_4912,N_5638);
nor U7301 (N_7301,N_4883,N_4688);
nand U7302 (N_7302,N_5053,N_4933);
and U7303 (N_7303,N_5420,N_5173);
nand U7304 (N_7304,N_4578,N_5138);
nor U7305 (N_7305,N_5491,N_5988);
nor U7306 (N_7306,N_5796,N_4756);
nor U7307 (N_7307,N_4828,N_5851);
nand U7308 (N_7308,N_4692,N_5164);
and U7309 (N_7309,N_4960,N_5866);
nor U7310 (N_7310,N_5471,N_5154);
xnor U7311 (N_7311,N_5580,N_5985);
or U7312 (N_7312,N_5792,N_4576);
or U7313 (N_7313,N_5947,N_5117);
nor U7314 (N_7314,N_4745,N_5618);
nor U7315 (N_7315,N_5163,N_5645);
or U7316 (N_7316,N_4555,N_5127);
or U7317 (N_7317,N_5091,N_4838);
or U7318 (N_7318,N_4586,N_4887);
nand U7319 (N_7319,N_5817,N_5782);
nor U7320 (N_7320,N_5589,N_5447);
or U7321 (N_7321,N_5641,N_4913);
or U7322 (N_7322,N_4626,N_5766);
nor U7323 (N_7323,N_4612,N_4546);
xor U7324 (N_7324,N_4860,N_5631);
nand U7325 (N_7325,N_5022,N_5897);
nor U7326 (N_7326,N_5060,N_5613);
or U7327 (N_7327,N_5847,N_4828);
xnor U7328 (N_7328,N_5051,N_5840);
nor U7329 (N_7329,N_4731,N_5090);
nand U7330 (N_7330,N_5701,N_4805);
nor U7331 (N_7331,N_4721,N_5509);
or U7332 (N_7332,N_5805,N_4925);
or U7333 (N_7333,N_5353,N_4884);
xor U7334 (N_7334,N_5234,N_4719);
xnor U7335 (N_7335,N_5319,N_5856);
nor U7336 (N_7336,N_4740,N_4784);
nor U7337 (N_7337,N_5355,N_5938);
xnor U7338 (N_7338,N_5401,N_5164);
nor U7339 (N_7339,N_5812,N_4587);
nor U7340 (N_7340,N_5246,N_4692);
xor U7341 (N_7341,N_5124,N_5337);
nor U7342 (N_7342,N_5289,N_5328);
nand U7343 (N_7343,N_5702,N_5889);
nand U7344 (N_7344,N_5286,N_5614);
xnor U7345 (N_7345,N_5295,N_5284);
or U7346 (N_7346,N_4863,N_4855);
or U7347 (N_7347,N_5945,N_5593);
or U7348 (N_7348,N_5290,N_5306);
and U7349 (N_7349,N_5407,N_5902);
or U7350 (N_7350,N_5104,N_5220);
and U7351 (N_7351,N_5583,N_5910);
or U7352 (N_7352,N_5662,N_5434);
nand U7353 (N_7353,N_5967,N_4722);
or U7354 (N_7354,N_5184,N_4833);
xnor U7355 (N_7355,N_5395,N_5317);
and U7356 (N_7356,N_5520,N_4726);
nand U7357 (N_7357,N_5897,N_5245);
and U7358 (N_7358,N_5922,N_4588);
nor U7359 (N_7359,N_5681,N_5532);
xor U7360 (N_7360,N_4537,N_5900);
nand U7361 (N_7361,N_4804,N_4522);
and U7362 (N_7362,N_5927,N_5764);
nand U7363 (N_7363,N_4702,N_4661);
nand U7364 (N_7364,N_4789,N_5172);
xnor U7365 (N_7365,N_5733,N_5985);
nand U7366 (N_7366,N_5150,N_5810);
nor U7367 (N_7367,N_4548,N_4580);
xnor U7368 (N_7368,N_5623,N_4646);
or U7369 (N_7369,N_5322,N_5152);
or U7370 (N_7370,N_5362,N_4841);
nand U7371 (N_7371,N_5578,N_4741);
nor U7372 (N_7372,N_4821,N_5711);
or U7373 (N_7373,N_5803,N_4517);
and U7374 (N_7374,N_5535,N_5976);
or U7375 (N_7375,N_5502,N_4683);
and U7376 (N_7376,N_4570,N_5997);
nor U7377 (N_7377,N_5115,N_5095);
nand U7378 (N_7378,N_5042,N_4595);
xnor U7379 (N_7379,N_4606,N_5700);
nand U7380 (N_7380,N_5115,N_5369);
nand U7381 (N_7381,N_4650,N_4525);
xnor U7382 (N_7382,N_4998,N_5975);
xnor U7383 (N_7383,N_5479,N_5231);
nor U7384 (N_7384,N_5349,N_5041);
or U7385 (N_7385,N_5313,N_5890);
nand U7386 (N_7386,N_5773,N_5928);
nor U7387 (N_7387,N_5666,N_5388);
or U7388 (N_7388,N_5795,N_5278);
xnor U7389 (N_7389,N_5581,N_4728);
xnor U7390 (N_7390,N_5899,N_5480);
xnor U7391 (N_7391,N_5641,N_4508);
or U7392 (N_7392,N_5821,N_5266);
and U7393 (N_7393,N_5605,N_4527);
nand U7394 (N_7394,N_5644,N_5335);
and U7395 (N_7395,N_5368,N_5431);
or U7396 (N_7396,N_4993,N_5721);
xor U7397 (N_7397,N_5773,N_5221);
and U7398 (N_7398,N_4956,N_5488);
xor U7399 (N_7399,N_5048,N_4510);
or U7400 (N_7400,N_5657,N_5816);
xnor U7401 (N_7401,N_4722,N_5304);
xnor U7402 (N_7402,N_5367,N_4537);
xnor U7403 (N_7403,N_4500,N_4668);
and U7404 (N_7404,N_4874,N_5661);
nor U7405 (N_7405,N_5983,N_4891);
xnor U7406 (N_7406,N_4962,N_5484);
nand U7407 (N_7407,N_5418,N_5397);
or U7408 (N_7408,N_5771,N_5838);
or U7409 (N_7409,N_5036,N_5886);
nand U7410 (N_7410,N_4664,N_5629);
or U7411 (N_7411,N_5598,N_5771);
or U7412 (N_7412,N_4855,N_4847);
xor U7413 (N_7413,N_4574,N_5421);
nor U7414 (N_7414,N_5450,N_4590);
nand U7415 (N_7415,N_4587,N_4973);
nor U7416 (N_7416,N_4597,N_4842);
xnor U7417 (N_7417,N_5486,N_5522);
nand U7418 (N_7418,N_5483,N_4525);
nor U7419 (N_7419,N_4715,N_5201);
xnor U7420 (N_7420,N_4838,N_5318);
xor U7421 (N_7421,N_4778,N_4723);
or U7422 (N_7422,N_5049,N_5527);
nor U7423 (N_7423,N_4823,N_5624);
and U7424 (N_7424,N_4675,N_5628);
nand U7425 (N_7425,N_5543,N_4927);
nor U7426 (N_7426,N_5144,N_4738);
nor U7427 (N_7427,N_5858,N_4602);
or U7428 (N_7428,N_5487,N_5433);
nand U7429 (N_7429,N_5768,N_5071);
or U7430 (N_7430,N_4823,N_4961);
and U7431 (N_7431,N_5108,N_4868);
xnor U7432 (N_7432,N_5549,N_5976);
nand U7433 (N_7433,N_5868,N_5377);
and U7434 (N_7434,N_4548,N_5608);
xnor U7435 (N_7435,N_4818,N_5416);
xnor U7436 (N_7436,N_4641,N_5040);
nand U7437 (N_7437,N_5978,N_4930);
and U7438 (N_7438,N_5024,N_4846);
nor U7439 (N_7439,N_4999,N_5519);
xor U7440 (N_7440,N_5529,N_5854);
xnor U7441 (N_7441,N_5876,N_4575);
nor U7442 (N_7442,N_4783,N_5340);
xor U7443 (N_7443,N_5086,N_5730);
nand U7444 (N_7444,N_5633,N_5743);
nor U7445 (N_7445,N_5296,N_4898);
or U7446 (N_7446,N_5785,N_5563);
nand U7447 (N_7447,N_4749,N_4804);
xnor U7448 (N_7448,N_4711,N_5788);
or U7449 (N_7449,N_4801,N_4788);
or U7450 (N_7450,N_5953,N_5410);
or U7451 (N_7451,N_5302,N_5580);
and U7452 (N_7452,N_5581,N_4798);
nand U7453 (N_7453,N_4947,N_5743);
nand U7454 (N_7454,N_4729,N_4518);
and U7455 (N_7455,N_4693,N_4615);
and U7456 (N_7456,N_5621,N_5646);
nand U7457 (N_7457,N_5055,N_4792);
or U7458 (N_7458,N_5276,N_5182);
and U7459 (N_7459,N_5328,N_5014);
nor U7460 (N_7460,N_5657,N_5652);
nand U7461 (N_7461,N_5357,N_5883);
xnor U7462 (N_7462,N_5960,N_5771);
nor U7463 (N_7463,N_4535,N_5719);
xnor U7464 (N_7464,N_5605,N_4999);
xor U7465 (N_7465,N_5441,N_5370);
or U7466 (N_7466,N_5435,N_4718);
nand U7467 (N_7467,N_5687,N_4819);
or U7468 (N_7468,N_5649,N_5856);
or U7469 (N_7469,N_4510,N_5948);
and U7470 (N_7470,N_4931,N_5490);
nand U7471 (N_7471,N_5601,N_5921);
and U7472 (N_7472,N_5985,N_5494);
xnor U7473 (N_7473,N_5418,N_5196);
nor U7474 (N_7474,N_5331,N_5854);
nand U7475 (N_7475,N_4706,N_5381);
nor U7476 (N_7476,N_4847,N_5326);
or U7477 (N_7477,N_4625,N_4722);
nand U7478 (N_7478,N_4932,N_4609);
and U7479 (N_7479,N_5882,N_5908);
nand U7480 (N_7480,N_4708,N_5127);
nand U7481 (N_7481,N_5196,N_5098);
xor U7482 (N_7482,N_5781,N_5804);
and U7483 (N_7483,N_5977,N_5590);
nand U7484 (N_7484,N_5474,N_4834);
and U7485 (N_7485,N_5872,N_5188);
xor U7486 (N_7486,N_4825,N_4519);
nand U7487 (N_7487,N_4880,N_4601);
and U7488 (N_7488,N_5535,N_5934);
xor U7489 (N_7489,N_5994,N_5449);
and U7490 (N_7490,N_4866,N_4982);
nor U7491 (N_7491,N_4618,N_4891);
xor U7492 (N_7492,N_5897,N_4722);
or U7493 (N_7493,N_5396,N_5158);
and U7494 (N_7494,N_4908,N_5362);
nand U7495 (N_7495,N_5385,N_5989);
and U7496 (N_7496,N_5826,N_5525);
xor U7497 (N_7497,N_5448,N_5145);
nand U7498 (N_7498,N_5000,N_4928);
nor U7499 (N_7499,N_4850,N_5858);
or U7500 (N_7500,N_7054,N_6064);
nor U7501 (N_7501,N_7316,N_6834);
xnor U7502 (N_7502,N_7340,N_7288);
or U7503 (N_7503,N_6151,N_6517);
nand U7504 (N_7504,N_6004,N_6667);
nor U7505 (N_7505,N_6784,N_6943);
nor U7506 (N_7506,N_6208,N_6286);
nand U7507 (N_7507,N_7448,N_6692);
nor U7508 (N_7508,N_7167,N_6913);
or U7509 (N_7509,N_6197,N_6966);
xnor U7510 (N_7510,N_7387,N_6069);
and U7511 (N_7511,N_7335,N_6079);
xor U7512 (N_7512,N_6068,N_7375);
and U7513 (N_7513,N_7108,N_7256);
xor U7514 (N_7514,N_6283,N_7091);
nand U7515 (N_7515,N_6923,N_6013);
or U7516 (N_7516,N_6685,N_6892);
xnor U7517 (N_7517,N_6594,N_6108);
and U7518 (N_7518,N_7456,N_6718);
nor U7519 (N_7519,N_6047,N_6840);
or U7520 (N_7520,N_6462,N_7084);
nand U7521 (N_7521,N_6878,N_6478);
and U7522 (N_7522,N_6743,N_6691);
xnor U7523 (N_7523,N_6779,N_6360);
nor U7524 (N_7524,N_6401,N_7396);
nor U7525 (N_7525,N_6346,N_6394);
or U7526 (N_7526,N_6119,N_7028);
nor U7527 (N_7527,N_7063,N_7174);
nand U7528 (N_7528,N_6760,N_7219);
nand U7529 (N_7529,N_7402,N_7373);
nor U7530 (N_7530,N_6989,N_6166);
or U7531 (N_7531,N_7092,N_6547);
and U7532 (N_7532,N_7045,N_6831);
nand U7533 (N_7533,N_7380,N_7474);
nand U7534 (N_7534,N_7309,N_6527);
nor U7535 (N_7535,N_6549,N_7307);
or U7536 (N_7536,N_7194,N_6332);
or U7537 (N_7537,N_6537,N_6931);
nor U7538 (N_7538,N_6277,N_6359);
xnor U7539 (N_7539,N_7445,N_6444);
nor U7540 (N_7540,N_7107,N_6920);
xor U7541 (N_7541,N_6625,N_6599);
xor U7542 (N_7542,N_7218,N_6681);
and U7543 (N_7543,N_6876,N_6765);
and U7544 (N_7544,N_7186,N_6485);
and U7545 (N_7545,N_6821,N_6545);
nand U7546 (N_7546,N_6341,N_6597);
and U7547 (N_7547,N_6149,N_6621);
xnor U7548 (N_7548,N_6045,N_6483);
nand U7549 (N_7549,N_7144,N_7357);
xnor U7550 (N_7550,N_6558,N_6721);
and U7551 (N_7551,N_7492,N_6933);
nor U7552 (N_7552,N_6790,N_6805);
nand U7553 (N_7553,N_6023,N_7113);
xnor U7554 (N_7554,N_6622,N_6315);
nand U7555 (N_7555,N_6711,N_7188);
and U7556 (N_7556,N_6000,N_6115);
xor U7557 (N_7557,N_7130,N_7459);
or U7558 (N_7558,N_6551,N_6266);
nand U7559 (N_7559,N_6781,N_6252);
and U7560 (N_7560,N_6029,N_7145);
nand U7561 (N_7561,N_6814,N_6163);
xnor U7562 (N_7562,N_6010,N_7290);
nand U7563 (N_7563,N_7035,N_7246);
and U7564 (N_7564,N_6526,N_6435);
or U7565 (N_7565,N_7417,N_6355);
xor U7566 (N_7566,N_7230,N_6492);
and U7567 (N_7567,N_7315,N_6875);
xnor U7568 (N_7568,N_6240,N_7351);
nand U7569 (N_7569,N_7029,N_6367);
nand U7570 (N_7570,N_6124,N_6123);
xnor U7571 (N_7571,N_7025,N_6279);
and U7572 (N_7572,N_6179,N_6488);
nand U7573 (N_7573,N_7381,N_6648);
or U7574 (N_7574,N_6481,N_6349);
or U7575 (N_7575,N_7329,N_7434);
xor U7576 (N_7576,N_6363,N_6410);
nor U7577 (N_7577,N_6906,N_7319);
and U7578 (N_7578,N_7300,N_7242);
nand U7579 (N_7579,N_7070,N_7446);
and U7580 (N_7580,N_7318,N_6869);
or U7581 (N_7581,N_6027,N_6505);
or U7582 (N_7582,N_6979,N_6147);
or U7583 (N_7583,N_6601,N_7040);
or U7584 (N_7584,N_6881,N_6736);
or U7585 (N_7585,N_7111,N_6969);
nand U7586 (N_7586,N_6998,N_6055);
xnor U7587 (N_7587,N_7237,N_6666);
xor U7588 (N_7588,N_7075,N_6433);
nand U7589 (N_7589,N_7385,N_6173);
and U7590 (N_7590,N_6323,N_6523);
and U7591 (N_7591,N_7039,N_6971);
xnor U7592 (N_7592,N_7293,N_6900);
or U7593 (N_7593,N_7216,N_6705);
or U7594 (N_7594,N_7151,N_6375);
or U7595 (N_7595,N_7060,N_6986);
nor U7596 (N_7596,N_6507,N_6334);
and U7597 (N_7597,N_7030,N_6562);
nor U7598 (N_7598,N_7048,N_6511);
nor U7599 (N_7599,N_6466,N_6644);
or U7600 (N_7600,N_7409,N_6372);
or U7601 (N_7601,N_6141,N_6019);
nand U7602 (N_7602,N_7401,N_6182);
nand U7603 (N_7603,N_6387,N_6703);
nand U7604 (N_7604,N_7490,N_7245);
or U7605 (N_7605,N_6215,N_6871);
nand U7606 (N_7606,N_7481,N_7143);
xor U7607 (N_7607,N_6585,N_7200);
and U7608 (N_7608,N_7422,N_7004);
nor U7609 (N_7609,N_6991,N_6615);
xor U7610 (N_7610,N_7299,N_7050);
nand U7611 (N_7611,N_6139,N_6500);
and U7612 (N_7612,N_6620,N_7198);
and U7613 (N_7613,N_7139,N_7163);
xor U7614 (N_7614,N_7394,N_6235);
nor U7615 (N_7615,N_6456,N_7160);
xnor U7616 (N_7616,N_6860,N_6231);
nand U7617 (N_7617,N_7213,N_7240);
xor U7618 (N_7618,N_6428,N_7430);
nand U7619 (N_7619,N_6476,N_6455);
nand U7620 (N_7620,N_6312,N_6114);
xnor U7621 (N_7621,N_6745,N_7243);
xnor U7622 (N_7622,N_6651,N_6659);
xnor U7623 (N_7623,N_6270,N_7125);
or U7624 (N_7624,N_6710,N_7444);
or U7625 (N_7625,N_6160,N_6035);
nand U7626 (N_7626,N_6824,N_6448);
nor U7627 (N_7627,N_6238,N_7023);
and U7628 (N_7628,N_6624,N_6596);
or U7629 (N_7629,N_7321,N_6144);
or U7630 (N_7630,N_7497,N_6351);
and U7631 (N_7631,N_6501,N_6944);
nand U7632 (N_7632,N_6614,N_7159);
and U7633 (N_7633,N_6598,N_6934);
and U7634 (N_7634,N_6085,N_6409);
xnor U7635 (N_7635,N_7291,N_6643);
xor U7636 (N_7636,N_6928,N_7332);
and U7637 (N_7637,N_7486,N_6259);
nand U7638 (N_7638,N_6138,N_7333);
nor U7639 (N_7639,N_6749,N_6439);
xnor U7640 (N_7640,N_6411,N_6084);
nor U7641 (N_7641,N_6185,N_6515);
xnor U7642 (N_7642,N_6532,N_6525);
nand U7643 (N_7643,N_6368,N_6136);
xor U7644 (N_7644,N_6658,N_6070);
and U7645 (N_7645,N_6239,N_6497);
and U7646 (N_7646,N_6992,N_7372);
and U7647 (N_7647,N_6775,N_6699);
xnor U7648 (N_7648,N_7146,N_6945);
or U7649 (N_7649,N_6832,N_6377);
xnor U7650 (N_7650,N_7005,N_6091);
xnor U7651 (N_7651,N_6129,N_7418);
or U7652 (N_7652,N_6168,N_7353);
xnor U7653 (N_7653,N_6778,N_6678);
xnor U7654 (N_7654,N_6234,N_6285);
or U7655 (N_7655,N_6042,N_7432);
nor U7656 (N_7656,N_6586,N_6113);
nand U7657 (N_7657,N_6970,N_6227);
or U7658 (N_7658,N_6740,N_6726);
nor U7659 (N_7659,N_7308,N_6797);
nand U7660 (N_7660,N_6610,N_6403);
or U7661 (N_7661,N_7260,N_6461);
nor U7662 (N_7662,N_6954,N_6521);
or U7663 (N_7663,N_6443,N_7026);
xnor U7664 (N_7664,N_6415,N_6157);
xor U7665 (N_7665,N_6962,N_6660);
nand U7666 (N_7666,N_6929,N_6072);
nor U7667 (N_7667,N_6078,N_6026);
and U7668 (N_7668,N_6490,N_6339);
xnor U7669 (N_7669,N_6327,N_7475);
and U7670 (N_7670,N_6576,N_6959);
or U7671 (N_7671,N_7449,N_6416);
and U7672 (N_7672,N_6390,N_6417);
and U7673 (N_7673,N_6309,N_6608);
xnor U7674 (N_7674,N_6353,N_6216);
or U7675 (N_7675,N_6406,N_7201);
nor U7676 (N_7676,N_6189,N_6039);
nand U7677 (N_7677,N_6638,N_6534);
and U7678 (N_7678,N_6287,N_7082);
and U7679 (N_7679,N_7129,N_7354);
or U7680 (N_7680,N_7367,N_6720);
nor U7681 (N_7681,N_6102,N_6661);
or U7682 (N_7682,N_6373,N_7002);
or U7683 (N_7683,N_6841,N_7410);
nor U7684 (N_7684,N_7020,N_6117);
xnor U7685 (N_7685,N_7262,N_6898);
nand U7686 (N_7686,N_6708,N_6634);
and U7687 (N_7687,N_6901,N_6260);
nand U7688 (N_7688,N_6542,N_7115);
nor U7689 (N_7689,N_6434,N_6310);
nand U7690 (N_7690,N_6299,N_6639);
nor U7691 (N_7691,N_6391,N_6686);
nand U7692 (N_7692,N_7133,N_6024);
nand U7693 (N_7693,N_7093,N_7205);
or U7694 (N_7694,N_6487,N_6696);
nand U7695 (N_7695,N_6999,N_7429);
xnor U7696 (N_7696,N_6771,N_6879);
xnor U7697 (N_7697,N_6171,N_6762);
and U7698 (N_7698,N_6975,N_6008);
xor U7699 (N_7699,N_6093,N_6005);
xor U7700 (N_7700,N_6963,N_7254);
nor U7701 (N_7701,N_7470,N_7202);
xor U7702 (N_7702,N_6473,N_7124);
nand U7703 (N_7703,N_6425,N_7136);
nand U7704 (N_7704,N_6172,N_6396);
nand U7705 (N_7705,N_6637,N_6071);
and U7706 (N_7706,N_7206,N_6167);
xor U7707 (N_7707,N_6715,N_6449);
nor U7708 (N_7708,N_6857,N_6995);
nor U7709 (N_7709,N_6431,N_6746);
and U7710 (N_7710,N_6393,N_7066);
and U7711 (N_7711,N_7140,N_6541);
nor U7712 (N_7712,N_6578,N_7441);
and U7713 (N_7713,N_6100,N_6539);
nor U7714 (N_7714,N_6560,N_7489);
xor U7715 (N_7715,N_7261,N_7487);
nor U7716 (N_7716,N_6910,N_7494);
nor U7717 (N_7717,N_7350,N_7000);
or U7718 (N_7718,N_6727,N_6628);
nor U7719 (N_7719,N_6827,N_6502);
nand U7720 (N_7720,N_6981,N_6801);
xnor U7721 (N_7721,N_6424,N_7480);
nor U7722 (N_7722,N_6499,N_6003);
nand U7723 (N_7723,N_7165,N_6457);
nand U7724 (N_7724,N_7241,N_6633);
nor U7725 (N_7725,N_6063,N_6818);
xnor U7726 (N_7726,N_7024,N_6052);
xnor U7727 (N_7727,N_7021,N_7119);
nor U7728 (N_7728,N_6577,N_7484);
nor U7729 (N_7729,N_7104,N_7226);
nor U7730 (N_7730,N_6122,N_6858);
nand U7731 (N_7731,N_6847,N_7064);
nor U7732 (N_7732,N_6595,N_6641);
nand U7733 (N_7733,N_6739,N_6925);
nor U7734 (N_7734,N_7478,N_6036);
or U7735 (N_7735,N_6237,N_6571);
nor U7736 (N_7736,N_7452,N_6861);
and U7737 (N_7737,N_6965,N_6081);
nor U7738 (N_7738,N_6961,N_6978);
nand U7739 (N_7739,N_6421,N_7098);
and U7740 (N_7740,N_6859,N_6230);
and U7741 (N_7741,N_7044,N_7031);
or U7742 (N_7742,N_7471,N_6125);
and U7743 (N_7743,N_7339,N_6581);
nand U7744 (N_7744,N_7062,N_6932);
nor U7745 (N_7745,N_6697,N_6565);
xor U7746 (N_7746,N_7424,N_6130);
or U7747 (N_7747,N_6572,N_6937);
and U7748 (N_7748,N_6698,N_7152);
and U7749 (N_7749,N_6265,N_6987);
or U7750 (N_7750,N_6912,N_6960);
or U7751 (N_7751,N_6343,N_6142);
nor U7752 (N_7752,N_7110,N_6682);
or U7753 (N_7753,N_7466,N_6664);
or U7754 (N_7754,N_7232,N_6430);
nor U7755 (N_7755,N_6616,N_6973);
xor U7756 (N_7756,N_7345,N_6848);
xnor U7757 (N_7757,N_6494,N_6398);
or U7758 (N_7758,N_6675,N_6447);
nor U7759 (N_7759,N_6942,N_6303);
or U7760 (N_7760,N_7341,N_7343);
or U7761 (N_7761,N_6330,N_6754);
and U7762 (N_7762,N_6313,N_6025);
nand U7763 (N_7763,N_7181,N_6165);
and U7764 (N_7764,N_6076,N_6935);
nand U7765 (N_7765,N_7297,N_6800);
nor U7766 (N_7766,N_6470,N_6017);
xor U7767 (N_7767,N_6742,N_7313);
nand U7768 (N_7768,N_6241,N_7137);
nor U7769 (N_7769,N_6738,N_6325);
nand U7770 (N_7770,N_6938,N_6217);
xnor U7771 (N_7771,N_6164,N_6210);
and U7772 (N_7772,N_6947,N_6837);
xor U7773 (N_7773,N_7338,N_7118);
and U7774 (N_7774,N_6680,N_7266);
or U7775 (N_7775,N_6802,N_6657);
and U7776 (N_7776,N_7461,N_6649);
xor U7777 (N_7777,N_7094,N_7013);
and U7778 (N_7778,N_6066,N_7427);
nand U7779 (N_7779,N_7052,N_6361);
or U7780 (N_7780,N_7056,N_7325);
nand U7781 (N_7781,N_7042,N_6438);
nand U7782 (N_7782,N_6324,N_7252);
and U7783 (N_7783,N_6101,N_7349);
and U7784 (N_7784,N_7102,N_6154);
nor U7785 (N_7785,N_7249,N_7172);
or U7786 (N_7786,N_6573,N_6250);
nand U7787 (N_7787,N_7276,N_6020);
nor U7788 (N_7788,N_7404,N_7154);
nand U7789 (N_7789,N_6441,N_6750);
nand U7790 (N_7790,N_6180,N_6980);
nor U7791 (N_7791,N_6903,N_7083);
or U7792 (N_7792,N_6865,N_7057);
xor U7793 (N_7793,N_6451,N_7199);
xnor U7794 (N_7794,N_6902,N_6090);
xor U7795 (N_7795,N_6253,N_6899);
or U7796 (N_7796,N_6034,N_6564);
and U7797 (N_7797,N_6278,N_7175);
nor U7798 (N_7798,N_7184,N_7499);
nand U7799 (N_7799,N_6924,N_6673);
and U7800 (N_7800,N_6789,N_6040);
nand U7801 (N_7801,N_7458,N_6550);
and U7802 (N_7802,N_6529,N_6491);
xnor U7803 (N_7803,N_7298,N_6722);
and U7804 (N_7804,N_6972,N_6022);
xor U7805 (N_7805,N_7037,N_7248);
and U7806 (N_7806,N_6612,N_7149);
or U7807 (N_7807,N_6508,N_6689);
and U7808 (N_7808,N_6314,N_7009);
and U7809 (N_7809,N_6716,N_6719);
or U7810 (N_7810,N_6246,N_6380);
nor U7811 (N_7811,N_6856,N_6940);
nor U7812 (N_7812,N_7334,N_7450);
nor U7813 (N_7813,N_6833,N_7324);
or U7814 (N_7814,N_6242,N_6099);
nor U7815 (N_7815,N_6553,N_7431);
and U7816 (N_7816,N_7155,N_6582);
nor U7817 (N_7817,N_6060,N_7120);
nor U7818 (N_7818,N_6559,N_7421);
xor U7819 (N_7819,N_6748,N_7126);
nand U7820 (N_7820,N_7277,N_6904);
nand U7821 (N_7821,N_7271,N_6674);
nand U7822 (N_7822,N_7142,N_6062);
nand U7823 (N_7823,N_7428,N_7073);
xor U7824 (N_7824,N_6484,N_6662);
nand U7825 (N_7825,N_7089,N_7437);
and U7826 (N_7826,N_6528,N_6463);
nor U7827 (N_7827,N_6602,N_7258);
nor U7828 (N_7828,N_6994,N_7166);
nor U7829 (N_7829,N_6454,N_6606);
xor U7830 (N_7830,N_6863,N_7247);
or U7831 (N_7831,N_6844,N_7229);
or U7832 (N_7832,N_6236,N_6429);
nand U7833 (N_7833,N_6561,N_6838);
nor U7834 (N_7834,N_6317,N_6244);
and U7835 (N_7835,N_6836,N_6877);
and U7836 (N_7836,N_6195,N_7074);
or U7837 (N_7837,N_6474,N_6756);
and U7838 (N_7838,N_7103,N_7231);
and U7839 (N_7839,N_6701,N_7457);
nand U7840 (N_7840,N_6759,N_7388);
or U7841 (N_7841,N_6348,N_6524);
xor U7842 (N_7842,N_7420,N_6530);
nor U7843 (N_7843,N_6974,N_6894);
and U7844 (N_7844,N_6379,N_6829);
xor U7845 (N_7845,N_6326,N_6137);
xor U7846 (N_7846,N_6150,N_6870);
nand U7847 (N_7847,N_6471,N_7150);
xnor U7848 (N_7848,N_6049,N_6964);
xnor U7849 (N_7849,N_6446,N_7378);
or U7850 (N_7850,N_6842,N_7001);
xnor U7851 (N_7851,N_6132,N_6272);
nor U7852 (N_7852,N_6819,N_7365);
nor U7853 (N_7853,N_7384,N_7036);
nand U7854 (N_7854,N_6798,N_6053);
nor U7855 (N_7855,N_7304,N_6785);
or U7856 (N_7856,N_6825,N_7192);
nor U7857 (N_7857,N_7018,N_6219);
nor U7858 (N_7858,N_6282,N_6522);
and U7859 (N_7859,N_6795,N_6952);
nor U7860 (N_7860,N_7389,N_7439);
nor U7861 (N_7861,N_6713,N_6128);
and U7862 (N_7862,N_6854,N_6489);
nor U7863 (N_7863,N_6714,N_7121);
nor U7864 (N_7864,N_7485,N_6768);
nor U7865 (N_7865,N_6290,N_6477);
and U7866 (N_7866,N_6732,N_6201);
nor U7867 (N_7867,N_6245,N_6866);
nand U7868 (N_7868,N_7171,N_6028);
and U7869 (N_7869,N_6755,N_7051);
nand U7870 (N_7870,N_6362,N_7465);
xor U7871 (N_7871,N_6843,N_7253);
and U7872 (N_7872,N_6335,N_6226);
nand U7873 (N_7873,N_6757,N_7209);
nor U7874 (N_7874,N_7215,N_6222);
nand U7875 (N_7875,N_6298,N_7462);
nor U7876 (N_7876,N_6399,N_6887);
and U7877 (N_7877,N_6255,N_6918);
xnor U7878 (N_7878,N_6822,N_6958);
nand U7879 (N_7879,N_6583,N_7285);
nand U7880 (N_7880,N_7287,N_6949);
and U7881 (N_7881,N_6855,N_7483);
or U7882 (N_7882,N_6437,N_6450);
xnor U7883 (N_7883,N_7268,N_6280);
and U7884 (N_7884,N_6381,N_7019);
xor U7885 (N_7885,N_6220,N_7027);
or U7886 (N_7886,N_6709,N_7033);
nor U7887 (N_7887,N_6030,N_6120);
or U7888 (N_7888,N_7105,N_6806);
nor U7889 (N_7889,N_7408,N_7482);
and U7890 (N_7890,N_6690,N_7058);
xnor U7891 (N_7891,N_7468,N_6557);
xnor U7892 (N_7892,N_6460,N_6915);
nor U7893 (N_7893,N_6930,N_6533);
or U7894 (N_7894,N_7046,N_6518);
nand U7895 (N_7895,N_6316,N_7411);
nor U7896 (N_7896,N_6955,N_6849);
xor U7897 (N_7897,N_6385,N_6103);
or U7898 (N_7898,N_6654,N_7006);
xor U7899 (N_7899,N_6546,N_7012);
nand U7900 (N_7900,N_6402,N_7182);
nor U7901 (N_7901,N_7068,N_6872);
or U7902 (N_7902,N_6880,N_7179);
nand U7903 (N_7903,N_7127,N_7195);
nor U7904 (N_7904,N_7363,N_7162);
xnor U7905 (N_7905,N_7210,N_6774);
or U7906 (N_7906,N_6811,N_7217);
or U7907 (N_7907,N_7158,N_6788);
and U7908 (N_7908,N_6535,N_6472);
and U7909 (N_7909,N_6306,N_6273);
nor U7910 (N_7910,N_7259,N_7336);
xnor U7911 (N_7911,N_6555,N_6569);
and U7912 (N_7912,N_6092,N_7273);
and U7913 (N_7913,N_6383,N_6570);
and U7914 (N_7914,N_6397,N_6342);
xor U7915 (N_7915,N_6358,N_6687);
nand U7916 (N_7916,N_6941,N_7392);
nor U7917 (N_7917,N_6605,N_6480);
and U7918 (N_7918,N_6655,N_7153);
and U7919 (N_7919,N_7295,N_7269);
nand U7920 (N_7920,N_6556,N_6693);
xor U7921 (N_7921,N_7301,N_6772);
xnor U7922 (N_7922,N_7374,N_7122);
nand U7923 (N_7923,N_6207,N_6767);
or U7924 (N_7924,N_7358,N_6835);
or U7925 (N_7925,N_6823,N_6243);
and U7926 (N_7926,N_6683,N_6328);
nor U7927 (N_7927,N_7250,N_6589);
xnor U7928 (N_7928,N_6753,N_6552);
xor U7929 (N_7929,N_6187,N_7203);
and U7930 (N_7930,N_7224,N_7306);
and U7931 (N_7931,N_6810,N_6050);
or U7932 (N_7932,N_6203,N_7379);
xnor U7933 (N_7933,N_6131,N_6400);
and U7934 (N_7934,N_6412,N_7283);
nor U7935 (N_7935,N_7447,N_6882);
xnor U7936 (N_7936,N_6311,N_6468);
nor U7937 (N_7937,N_7370,N_7320);
and U7938 (N_7938,N_7178,N_7397);
nand U7939 (N_7939,N_6262,N_7348);
or U7940 (N_7940,N_6769,N_6777);
nand U7941 (N_7941,N_7138,N_6868);
xor U7942 (N_7942,N_6213,N_7112);
nand U7943 (N_7943,N_7106,N_6850);
xnor U7944 (N_7944,N_7225,N_6194);
or U7945 (N_7945,N_6015,N_6540);
and U7946 (N_7946,N_6791,N_7355);
nor U7947 (N_7947,N_6224,N_6631);
or U7948 (N_7948,N_6065,N_7011);
and U7949 (N_7949,N_6724,N_7323);
or U7950 (N_7950,N_6786,N_6618);
xnor U7951 (N_7951,N_6057,N_7041);
nor U7952 (N_7952,N_6075,N_7239);
xor U7953 (N_7953,N_6747,N_7101);
nand U7954 (N_7954,N_6922,N_6807);
nand U7955 (N_7955,N_7085,N_7128);
xnor U7956 (N_7956,N_6269,N_6169);
xnor U7957 (N_7957,N_7227,N_6640);
xnor U7958 (N_7958,N_7204,N_6820);
and U7959 (N_7959,N_6688,N_6983);
nand U7960 (N_7960,N_6404,N_6504);
nor U7961 (N_7961,N_6907,N_6885);
xor U7962 (N_7962,N_6080,N_6110);
and U7963 (N_7963,N_6896,N_6735);
nand U7964 (N_7964,N_6436,N_6751);
xor U7965 (N_7965,N_6803,N_6459);
xor U7966 (N_7966,N_6184,N_6074);
nand U7967 (N_7967,N_6734,N_6408);
nand U7968 (N_7968,N_6354,N_7134);
and U7969 (N_7969,N_7177,N_6737);
nand U7970 (N_7970,N_7327,N_6853);
or U7971 (N_7971,N_7087,N_6544);
and U7972 (N_7972,N_6851,N_7117);
nand U7973 (N_7973,N_6752,N_6482);
and U7974 (N_7974,N_6432,N_6916);
xor U7975 (N_7975,N_6388,N_7311);
and U7976 (N_7976,N_6109,N_7148);
or U7977 (N_7977,N_6178,N_6225);
or U7978 (N_7978,N_6274,N_7435);
xor U7979 (N_7979,N_6469,N_7141);
xnor U7980 (N_7980,N_6982,N_6427);
and U7981 (N_7981,N_7359,N_6096);
or U7982 (N_7982,N_7047,N_7495);
xor U7983 (N_7983,N_7185,N_6506);
or U7984 (N_7984,N_6407,N_6389);
xor U7985 (N_7985,N_6374,N_7438);
nor U7986 (N_7986,N_6744,N_6190);
nor U7987 (N_7987,N_6232,N_6672);
and U7988 (N_7988,N_6567,N_6414);
and U7989 (N_7989,N_7472,N_6116);
xnor U7990 (N_7990,N_6914,N_6318);
xor U7991 (N_7991,N_6148,N_6619);
xnor U7992 (N_7992,N_6319,N_7097);
and U7993 (N_7993,N_6809,N_6088);
nand U7994 (N_7994,N_7322,N_6543);
nand U7995 (N_7995,N_6095,N_6956);
or U7996 (N_7996,N_6369,N_7086);
nor U7997 (N_7997,N_6548,N_7377);
nor U7998 (N_7998,N_7053,N_7281);
xor U7999 (N_7999,N_6112,N_6665);
xor U8000 (N_8000,N_7114,N_6939);
and U8001 (N_8001,N_6647,N_6909);
or U8002 (N_8002,N_7017,N_6761);
xnor U8003 (N_8003,N_6635,N_6006);
nor U8004 (N_8004,N_6725,N_6264);
nor U8005 (N_8005,N_6950,N_7196);
and U8006 (N_8006,N_6308,N_6204);
nand U8007 (N_8007,N_6617,N_6083);
nand U8008 (N_8008,N_7015,N_6127);
xor U8009 (N_8009,N_7236,N_6782);
and U8010 (N_8010,N_6636,N_7352);
nor U8011 (N_8011,N_7233,N_6568);
or U8012 (N_8012,N_6193,N_7368);
xor U8013 (N_8013,N_6632,N_6340);
or U8014 (N_8014,N_7069,N_7426);
nor U8015 (N_8015,N_7081,N_7034);
or U8016 (N_8016,N_6174,N_7289);
or U8017 (N_8017,N_6927,N_6498);
and U8018 (N_8018,N_6267,N_6300);
nor U8019 (N_8019,N_6712,N_6007);
nor U8020 (N_8020,N_7223,N_6365);
nand U8021 (N_8021,N_6175,N_7493);
or U8022 (N_8022,N_6134,N_6170);
and U8023 (N_8023,N_6356,N_6817);
nor U8024 (N_8024,N_7065,N_7270);
nand U8025 (N_8025,N_6717,N_6580);
xor U8026 (N_8026,N_6845,N_6370);
and U8027 (N_8027,N_6307,N_6256);
or U8028 (N_8028,N_6413,N_6741);
nand U8029 (N_8029,N_6650,N_6209);
xor U8030 (N_8030,N_6073,N_6794);
nor U8031 (N_8031,N_6733,N_7376);
nor U8032 (N_8032,N_7328,N_6067);
and U8033 (N_8033,N_6105,N_6087);
xor U8034 (N_8034,N_6921,N_6611);
nand U8035 (N_8035,N_6516,N_7010);
and U8036 (N_8036,N_6161,N_6350);
nor U8037 (N_8037,N_7257,N_6574);
nand U8038 (N_8038,N_7049,N_6158);
nand U8039 (N_8039,N_6320,N_6593);
and U8040 (N_8040,N_6247,N_6082);
nand U8041 (N_8041,N_6812,N_6357);
nor U8042 (N_8042,N_6422,N_6271);
or U8043 (N_8043,N_6382,N_6936);
or U8044 (N_8044,N_7220,N_6893);
or U8045 (N_8045,N_6249,N_6951);
or U8046 (N_8046,N_6384,N_6452);
and U8047 (N_8047,N_6155,N_6192);
and U8048 (N_8048,N_7425,N_6419);
and U8049 (N_8049,N_6584,N_7067);
nor U8050 (N_8050,N_6159,N_7292);
or U8051 (N_8051,N_6152,N_7235);
and U8052 (N_8052,N_7415,N_7395);
nand U8053 (N_8053,N_6458,N_7043);
nor U8054 (N_8054,N_7423,N_6135);
nand U8055 (N_8055,N_7014,N_7071);
nor U8056 (N_8056,N_6206,N_6301);
xnor U8057 (N_8057,N_6405,N_6669);
xor U8058 (N_8058,N_6104,N_6867);
or U8059 (N_8059,N_7274,N_7022);
and U8060 (N_8060,N_7080,N_6826);
nor U8061 (N_8061,N_6813,N_6985);
nor U8062 (N_8062,N_6347,N_7265);
nor U8063 (N_8063,N_6630,N_7302);
nor U8064 (N_8064,N_6467,N_7440);
and U8065 (N_8065,N_6496,N_7488);
and U8066 (N_8066,N_6094,N_6156);
xnor U8067 (N_8067,N_6107,N_6176);
or U8068 (N_8068,N_7362,N_6294);
xnor U8069 (N_8069,N_6371,N_7059);
and U8070 (N_8070,N_6291,N_7190);
and U8071 (N_8071,N_7208,N_7310);
nor U8072 (N_8072,N_6297,N_7016);
xor U8073 (N_8073,N_6445,N_6627);
or U8074 (N_8074,N_6984,N_6479);
nor U8075 (N_8075,N_6322,N_7109);
and U8076 (N_8076,N_7442,N_6889);
nand U8077 (N_8077,N_7294,N_7364);
nor U8078 (N_8078,N_7371,N_6591);
xnor U8079 (N_8079,N_7038,N_7399);
nand U8080 (N_8080,N_6111,N_6228);
nor U8081 (N_8081,N_6033,N_6289);
or U8082 (N_8082,N_6338,N_6663);
and U8083 (N_8083,N_6623,N_6670);
nand U8084 (N_8084,N_7096,N_6002);
xnor U8085 (N_8085,N_6873,N_7100);
xor U8086 (N_8086,N_6191,N_6223);
xnor U8087 (N_8087,N_6146,N_7454);
or U8088 (N_8088,N_7383,N_6976);
or U8089 (N_8089,N_7400,N_7346);
and U8090 (N_8090,N_7406,N_7282);
and U8091 (N_8091,N_6926,N_6776);
nand U8092 (N_8092,N_7267,N_6538);
nor U8093 (N_8093,N_7275,N_7366);
and U8094 (N_8094,N_6783,N_6758);
nand U8095 (N_8095,N_6153,N_7286);
or U8096 (N_8096,N_7331,N_6183);
and U8097 (N_8097,N_6442,N_6799);
or U8098 (N_8098,N_6531,N_6626);
nor U8099 (N_8099,N_7116,N_6058);
nand U8100 (N_8100,N_6607,N_7079);
and U8101 (N_8101,N_6764,N_6031);
nand U8102 (N_8102,N_6423,N_6305);
and U8103 (N_8103,N_6337,N_6656);
or U8104 (N_8104,N_6588,N_6514);
nand U8105 (N_8105,N_6808,N_6609);
xnor U8106 (N_8106,N_7061,N_7491);
nand U8107 (N_8107,N_6766,N_6679);
nand U8108 (N_8108,N_7244,N_7284);
nor U8109 (N_8109,N_7419,N_6600);
nand U8110 (N_8110,N_7099,N_6186);
and U8111 (N_8111,N_7391,N_6864);
xor U8112 (N_8112,N_7222,N_6694);
and U8113 (N_8113,N_6495,N_6205);
xnor U8114 (N_8114,N_6464,N_6329);
and U8115 (N_8115,N_7342,N_6018);
and U8116 (N_8116,N_6276,N_6001);
nor U8117 (N_8117,N_6603,N_6919);
and U8118 (N_8118,N_6592,N_6792);
and U8119 (N_8119,N_6118,N_7464);
or U8120 (N_8120,N_6646,N_6671);
nand U8121 (N_8121,N_6181,N_6804);
xor U8122 (N_8122,N_6199,N_7238);
and U8123 (N_8123,N_6012,N_7207);
and U8124 (N_8124,N_7296,N_6575);
and U8125 (N_8125,N_7095,N_7436);
or U8126 (N_8126,N_6331,N_6106);
nand U8127 (N_8127,N_7164,N_6846);
or U8128 (N_8128,N_6061,N_6214);
xnor U8129 (N_8129,N_6728,N_7168);
or U8130 (N_8130,N_7279,N_6200);
or U8131 (N_8131,N_7403,N_7312);
or U8132 (N_8132,N_7479,N_6566);
nand U8133 (N_8133,N_6773,N_6378);
xnor U8134 (N_8134,N_6486,N_6037);
nand U8135 (N_8135,N_6133,N_6059);
and U8136 (N_8136,N_7003,N_6536);
nand U8137 (N_8137,N_6212,N_7135);
or U8138 (N_8138,N_6296,N_6780);
or U8139 (N_8139,N_7212,N_7131);
nor U8140 (N_8140,N_7330,N_6706);
nor U8141 (N_8141,N_7180,N_6392);
nand U8142 (N_8142,N_6288,N_6263);
or U8143 (N_8143,N_7390,N_6051);
or U8144 (N_8144,N_6874,N_6086);
nand U8145 (N_8145,N_6321,N_6221);
and U8146 (N_8146,N_7477,N_7090);
xor U8147 (N_8147,N_6275,N_6908);
nand U8148 (N_8148,N_6077,N_6891);
xor U8149 (N_8149,N_6590,N_6702);
nand U8150 (N_8150,N_6828,N_7088);
nor U8151 (N_8151,N_7473,N_7156);
nor U8152 (N_8152,N_7214,N_6304);
nor U8153 (N_8153,N_6044,N_6977);
nand U8154 (N_8154,N_6440,N_6009);
nand U8155 (N_8155,N_7416,N_7280);
or U8156 (N_8156,N_6890,N_7303);
nor U8157 (N_8157,N_6770,N_6883);
or U8158 (N_8158,N_6032,N_6089);
nor U8159 (N_8159,N_7078,N_7455);
nor U8160 (N_8160,N_6917,N_6613);
and U8161 (N_8161,N_7077,N_6731);
and U8162 (N_8162,N_6642,N_6519);
nor U8163 (N_8163,N_6520,N_7317);
xor U8164 (N_8164,N_6229,N_6704);
xnor U8165 (N_8165,N_7147,N_7443);
or U8166 (N_8166,N_6376,N_6302);
nor U8167 (N_8167,N_6014,N_6587);
and U8168 (N_8168,N_6295,N_7412);
and U8169 (N_8169,N_7032,N_7451);
nand U8170 (N_8170,N_6420,N_7453);
and U8171 (N_8171,N_6554,N_6258);
nand U8172 (N_8172,N_7193,N_6344);
or U8173 (N_8173,N_6793,N_6426);
xnor U8174 (N_8174,N_7251,N_7413);
or U8175 (N_8175,N_6996,N_6254);
and U8176 (N_8176,N_6905,N_7264);
nand U8177 (N_8177,N_6695,N_7460);
nor U8178 (N_8178,N_6503,N_6677);
xor U8179 (N_8179,N_6862,N_6948);
or U8180 (N_8180,N_6386,N_6126);
or U8181 (N_8181,N_6188,N_6395);
nand U8182 (N_8182,N_6011,N_7344);
and U8183 (N_8183,N_7191,N_7123);
nand U8184 (N_8184,N_6988,N_6493);
nand U8185 (N_8185,N_7467,N_7255);
nor U8186 (N_8186,N_7469,N_7405);
xor U8187 (N_8187,N_6098,N_6196);
xor U8188 (N_8188,N_6140,N_6563);
nor U8189 (N_8189,N_6465,N_6579);
nor U8190 (N_8190,N_7356,N_6418);
or U8191 (N_8191,N_7211,N_6993);
nor U8192 (N_8192,N_7360,N_6261);
xor U8193 (N_8193,N_7393,N_6763);
xor U8194 (N_8194,N_6211,N_6729);
nor U8195 (N_8195,N_6796,N_7498);
xor U8196 (N_8196,N_6281,N_6897);
nor U8197 (N_8197,N_6946,N_7170);
nor U8198 (N_8198,N_6967,N_7463);
and U8199 (N_8199,N_6048,N_6162);
nor U8200 (N_8200,N_7278,N_6097);
or U8201 (N_8201,N_7221,N_6645);
nor U8202 (N_8202,N_6653,N_6723);
nor U8203 (N_8203,N_7414,N_6839);
nand U8204 (N_8204,N_6352,N_6512);
xnor U8205 (N_8205,N_7369,N_6041);
and U8206 (N_8206,N_6911,N_6852);
nor U8207 (N_8207,N_7008,N_6202);
xnor U8208 (N_8208,N_6038,N_6676);
or U8209 (N_8209,N_6046,N_7132);
nor U8210 (N_8210,N_7007,N_7176);
xnor U8211 (N_8211,N_6054,N_6684);
nor U8212 (N_8212,N_7326,N_6895);
and U8213 (N_8213,N_6043,N_7072);
and U8214 (N_8214,N_6284,N_7347);
nand U8215 (N_8215,N_6143,N_7337);
or U8216 (N_8216,N_7234,N_7433);
or U8217 (N_8217,N_6513,N_6251);
nand U8218 (N_8218,N_6453,N_6629);
nand U8219 (N_8219,N_6364,N_6366);
nor U8220 (N_8220,N_6787,N_6145);
nand U8221 (N_8221,N_6668,N_6888);
nand U8222 (N_8222,N_6177,N_7076);
or U8223 (N_8223,N_6509,N_6016);
or U8224 (N_8224,N_7398,N_7305);
xor U8225 (N_8225,N_7055,N_6957);
and U8226 (N_8226,N_6121,N_6233);
xor U8227 (N_8227,N_7272,N_6604);
or U8228 (N_8228,N_7496,N_7197);
nand U8229 (N_8229,N_6816,N_7169);
xnor U8230 (N_8230,N_6968,N_6700);
nand U8231 (N_8231,N_6884,N_7228);
nand U8232 (N_8232,N_7386,N_7361);
nand U8233 (N_8233,N_6730,N_7187);
nor U8234 (N_8234,N_6815,N_7161);
or U8235 (N_8235,N_7382,N_6707);
xnor U8236 (N_8236,N_6990,N_7263);
xor U8237 (N_8237,N_7476,N_7173);
nor U8238 (N_8238,N_7157,N_6248);
nor U8239 (N_8239,N_6830,N_6886);
xor U8240 (N_8240,N_7189,N_6953);
and U8241 (N_8241,N_6292,N_6345);
xor U8242 (N_8242,N_6056,N_6293);
or U8243 (N_8243,N_6021,N_6268);
or U8244 (N_8244,N_6198,N_6652);
nand U8245 (N_8245,N_7314,N_6333);
nand U8246 (N_8246,N_6336,N_7183);
xnor U8247 (N_8247,N_6475,N_6997);
nand U8248 (N_8248,N_7407,N_6510);
nor U8249 (N_8249,N_6257,N_6218);
nand U8250 (N_8250,N_6700,N_7207);
xnor U8251 (N_8251,N_6867,N_7094);
nand U8252 (N_8252,N_6681,N_6478);
or U8253 (N_8253,N_6883,N_6258);
xnor U8254 (N_8254,N_6500,N_6444);
nor U8255 (N_8255,N_6949,N_6380);
or U8256 (N_8256,N_7499,N_6234);
and U8257 (N_8257,N_7356,N_6719);
or U8258 (N_8258,N_6805,N_6574);
nor U8259 (N_8259,N_6178,N_6858);
nand U8260 (N_8260,N_6659,N_6048);
or U8261 (N_8261,N_7075,N_7206);
and U8262 (N_8262,N_7068,N_6410);
nor U8263 (N_8263,N_6453,N_7446);
nand U8264 (N_8264,N_6402,N_7331);
nand U8265 (N_8265,N_6250,N_7145);
or U8266 (N_8266,N_7368,N_7039);
nand U8267 (N_8267,N_6925,N_7057);
xor U8268 (N_8268,N_6417,N_6643);
and U8269 (N_8269,N_6239,N_7446);
xor U8270 (N_8270,N_6055,N_6857);
nand U8271 (N_8271,N_6421,N_6657);
and U8272 (N_8272,N_7496,N_7027);
xor U8273 (N_8273,N_6938,N_6889);
and U8274 (N_8274,N_7397,N_7066);
xnor U8275 (N_8275,N_6624,N_7459);
or U8276 (N_8276,N_6851,N_7381);
nand U8277 (N_8277,N_7053,N_6112);
nor U8278 (N_8278,N_6768,N_6266);
and U8279 (N_8279,N_6676,N_6486);
nor U8280 (N_8280,N_7192,N_7062);
or U8281 (N_8281,N_6541,N_6429);
or U8282 (N_8282,N_6365,N_6893);
nand U8283 (N_8283,N_7422,N_7419);
and U8284 (N_8284,N_7417,N_6148);
or U8285 (N_8285,N_6261,N_7225);
xor U8286 (N_8286,N_7424,N_6488);
xnor U8287 (N_8287,N_6741,N_7346);
xor U8288 (N_8288,N_6539,N_6623);
or U8289 (N_8289,N_6268,N_6868);
nand U8290 (N_8290,N_6355,N_6421);
and U8291 (N_8291,N_6988,N_6333);
nor U8292 (N_8292,N_7438,N_6968);
and U8293 (N_8293,N_7279,N_6758);
nor U8294 (N_8294,N_7182,N_6215);
nand U8295 (N_8295,N_7013,N_6271);
and U8296 (N_8296,N_7306,N_7443);
and U8297 (N_8297,N_7497,N_6988);
xnor U8298 (N_8298,N_7427,N_7357);
and U8299 (N_8299,N_7331,N_7114);
nor U8300 (N_8300,N_6525,N_6530);
or U8301 (N_8301,N_6921,N_6377);
nor U8302 (N_8302,N_6956,N_6982);
nor U8303 (N_8303,N_6066,N_7405);
xnor U8304 (N_8304,N_6104,N_7473);
nand U8305 (N_8305,N_6675,N_6649);
nor U8306 (N_8306,N_7331,N_7209);
or U8307 (N_8307,N_6145,N_7019);
or U8308 (N_8308,N_6661,N_6386);
nor U8309 (N_8309,N_6687,N_7261);
and U8310 (N_8310,N_6764,N_6780);
nor U8311 (N_8311,N_6377,N_6968);
nor U8312 (N_8312,N_7422,N_7073);
and U8313 (N_8313,N_7220,N_6184);
nand U8314 (N_8314,N_7175,N_6560);
nor U8315 (N_8315,N_7361,N_6744);
and U8316 (N_8316,N_6235,N_7174);
xnor U8317 (N_8317,N_6701,N_7196);
xor U8318 (N_8318,N_6245,N_6023);
xnor U8319 (N_8319,N_7355,N_7246);
xnor U8320 (N_8320,N_6293,N_6259);
nor U8321 (N_8321,N_6489,N_6634);
nor U8322 (N_8322,N_6974,N_6191);
xnor U8323 (N_8323,N_6235,N_6043);
or U8324 (N_8324,N_6624,N_7213);
nor U8325 (N_8325,N_7392,N_7176);
or U8326 (N_8326,N_6980,N_6987);
and U8327 (N_8327,N_7241,N_7353);
nor U8328 (N_8328,N_6635,N_6617);
nor U8329 (N_8329,N_6270,N_6332);
xnor U8330 (N_8330,N_6791,N_6327);
xor U8331 (N_8331,N_7275,N_6210);
nor U8332 (N_8332,N_7351,N_6759);
nand U8333 (N_8333,N_6169,N_6080);
nand U8334 (N_8334,N_7164,N_6651);
and U8335 (N_8335,N_6897,N_6711);
xor U8336 (N_8336,N_6943,N_7052);
xor U8337 (N_8337,N_7077,N_6629);
or U8338 (N_8338,N_6787,N_6901);
and U8339 (N_8339,N_7021,N_7102);
nor U8340 (N_8340,N_6713,N_6995);
or U8341 (N_8341,N_6362,N_6853);
nand U8342 (N_8342,N_7372,N_6925);
nand U8343 (N_8343,N_6696,N_6106);
nand U8344 (N_8344,N_7023,N_6815);
or U8345 (N_8345,N_6639,N_6414);
nand U8346 (N_8346,N_6768,N_6843);
or U8347 (N_8347,N_6112,N_6279);
or U8348 (N_8348,N_6406,N_6883);
nor U8349 (N_8349,N_7098,N_6414);
and U8350 (N_8350,N_6179,N_6061);
nor U8351 (N_8351,N_6071,N_6983);
and U8352 (N_8352,N_7414,N_6914);
and U8353 (N_8353,N_6214,N_6265);
xor U8354 (N_8354,N_6697,N_6891);
nor U8355 (N_8355,N_6608,N_7482);
nand U8356 (N_8356,N_6985,N_6946);
nor U8357 (N_8357,N_6209,N_6995);
or U8358 (N_8358,N_6271,N_6738);
and U8359 (N_8359,N_6710,N_6731);
or U8360 (N_8360,N_7305,N_6802);
xnor U8361 (N_8361,N_6987,N_6163);
nand U8362 (N_8362,N_6151,N_7382);
nor U8363 (N_8363,N_6582,N_6494);
or U8364 (N_8364,N_7083,N_6579);
nor U8365 (N_8365,N_6812,N_6887);
xnor U8366 (N_8366,N_6856,N_6314);
nand U8367 (N_8367,N_6957,N_7394);
nor U8368 (N_8368,N_6859,N_7137);
nand U8369 (N_8369,N_7043,N_6107);
and U8370 (N_8370,N_7190,N_7331);
or U8371 (N_8371,N_6328,N_6931);
nor U8372 (N_8372,N_6002,N_7338);
nor U8373 (N_8373,N_6926,N_7263);
or U8374 (N_8374,N_6389,N_6199);
xor U8375 (N_8375,N_7471,N_6455);
or U8376 (N_8376,N_7219,N_6902);
nand U8377 (N_8377,N_7297,N_7011);
or U8378 (N_8378,N_7330,N_6633);
nor U8379 (N_8379,N_6644,N_6395);
nor U8380 (N_8380,N_7003,N_6363);
or U8381 (N_8381,N_6948,N_6502);
or U8382 (N_8382,N_6447,N_7017);
and U8383 (N_8383,N_6427,N_6529);
xnor U8384 (N_8384,N_7492,N_7472);
xor U8385 (N_8385,N_6456,N_7431);
or U8386 (N_8386,N_7010,N_6408);
xnor U8387 (N_8387,N_6732,N_7078);
or U8388 (N_8388,N_7147,N_6489);
xnor U8389 (N_8389,N_6272,N_6878);
xnor U8390 (N_8390,N_6810,N_7326);
xor U8391 (N_8391,N_7319,N_6846);
xor U8392 (N_8392,N_6592,N_6240);
nor U8393 (N_8393,N_7096,N_6701);
nand U8394 (N_8394,N_7174,N_7468);
nand U8395 (N_8395,N_6895,N_6688);
or U8396 (N_8396,N_6282,N_6217);
xor U8397 (N_8397,N_6665,N_6926);
nand U8398 (N_8398,N_6804,N_6737);
and U8399 (N_8399,N_6589,N_6766);
and U8400 (N_8400,N_6652,N_7040);
xnor U8401 (N_8401,N_7488,N_6164);
and U8402 (N_8402,N_7130,N_7495);
and U8403 (N_8403,N_7167,N_6010);
nor U8404 (N_8404,N_6135,N_7021);
xor U8405 (N_8405,N_6818,N_7496);
nand U8406 (N_8406,N_6574,N_7478);
and U8407 (N_8407,N_7345,N_6386);
or U8408 (N_8408,N_6855,N_7012);
xor U8409 (N_8409,N_6877,N_6691);
xnor U8410 (N_8410,N_6836,N_7119);
and U8411 (N_8411,N_7223,N_7182);
or U8412 (N_8412,N_7031,N_7431);
and U8413 (N_8413,N_7478,N_7445);
nor U8414 (N_8414,N_6761,N_6058);
nor U8415 (N_8415,N_6528,N_6583);
nand U8416 (N_8416,N_6827,N_6266);
nor U8417 (N_8417,N_7440,N_7081);
and U8418 (N_8418,N_6632,N_6065);
nand U8419 (N_8419,N_6711,N_6109);
or U8420 (N_8420,N_6565,N_6668);
or U8421 (N_8421,N_7454,N_6440);
and U8422 (N_8422,N_6078,N_7092);
nand U8423 (N_8423,N_7489,N_6613);
and U8424 (N_8424,N_6634,N_6079);
or U8425 (N_8425,N_6163,N_6182);
or U8426 (N_8426,N_6083,N_6498);
nand U8427 (N_8427,N_6577,N_7063);
and U8428 (N_8428,N_6782,N_7258);
xor U8429 (N_8429,N_7334,N_6981);
and U8430 (N_8430,N_7348,N_6160);
nand U8431 (N_8431,N_6892,N_6174);
xor U8432 (N_8432,N_6538,N_7065);
xor U8433 (N_8433,N_6436,N_6738);
nor U8434 (N_8434,N_6683,N_6348);
nor U8435 (N_8435,N_7024,N_6502);
nor U8436 (N_8436,N_7123,N_7422);
nor U8437 (N_8437,N_6673,N_7250);
or U8438 (N_8438,N_7019,N_6374);
or U8439 (N_8439,N_7168,N_7203);
and U8440 (N_8440,N_6641,N_6985);
nand U8441 (N_8441,N_6167,N_6348);
nand U8442 (N_8442,N_7485,N_7026);
nor U8443 (N_8443,N_6173,N_6549);
and U8444 (N_8444,N_6226,N_6026);
and U8445 (N_8445,N_6269,N_6190);
xnor U8446 (N_8446,N_7185,N_6642);
and U8447 (N_8447,N_6348,N_7399);
nor U8448 (N_8448,N_6933,N_6632);
and U8449 (N_8449,N_6080,N_6543);
nand U8450 (N_8450,N_7001,N_7143);
xnor U8451 (N_8451,N_6222,N_6043);
nor U8452 (N_8452,N_6376,N_6642);
and U8453 (N_8453,N_7055,N_6248);
nor U8454 (N_8454,N_7434,N_7441);
and U8455 (N_8455,N_6747,N_6633);
nor U8456 (N_8456,N_7014,N_7383);
xor U8457 (N_8457,N_6763,N_7465);
and U8458 (N_8458,N_6211,N_6988);
and U8459 (N_8459,N_6450,N_6890);
nand U8460 (N_8460,N_7191,N_6223);
nor U8461 (N_8461,N_6389,N_6157);
nor U8462 (N_8462,N_6318,N_6043);
xor U8463 (N_8463,N_6463,N_6396);
nand U8464 (N_8464,N_6614,N_7291);
nand U8465 (N_8465,N_6433,N_6753);
and U8466 (N_8466,N_7309,N_6991);
xor U8467 (N_8467,N_6806,N_6575);
xnor U8468 (N_8468,N_7000,N_6917);
xor U8469 (N_8469,N_7316,N_7406);
and U8470 (N_8470,N_6392,N_6466);
and U8471 (N_8471,N_6520,N_7122);
xnor U8472 (N_8472,N_7239,N_6273);
and U8473 (N_8473,N_7445,N_6705);
and U8474 (N_8474,N_7390,N_7027);
nand U8475 (N_8475,N_6269,N_7031);
and U8476 (N_8476,N_7264,N_6576);
nor U8477 (N_8477,N_6621,N_7430);
nor U8478 (N_8478,N_6111,N_6095);
nor U8479 (N_8479,N_7410,N_6637);
and U8480 (N_8480,N_7131,N_6441);
nor U8481 (N_8481,N_6254,N_6311);
xnor U8482 (N_8482,N_6872,N_6370);
xor U8483 (N_8483,N_6817,N_7153);
nor U8484 (N_8484,N_6393,N_6646);
or U8485 (N_8485,N_6103,N_7365);
xnor U8486 (N_8486,N_7354,N_6671);
or U8487 (N_8487,N_7279,N_6008);
and U8488 (N_8488,N_6078,N_7282);
or U8489 (N_8489,N_6003,N_6282);
xnor U8490 (N_8490,N_7256,N_6278);
and U8491 (N_8491,N_6350,N_6698);
and U8492 (N_8492,N_6562,N_7012);
or U8493 (N_8493,N_6791,N_6493);
xor U8494 (N_8494,N_7489,N_6079);
nand U8495 (N_8495,N_6398,N_6253);
or U8496 (N_8496,N_6795,N_7410);
and U8497 (N_8497,N_6198,N_6335);
nor U8498 (N_8498,N_6916,N_7148);
or U8499 (N_8499,N_7335,N_6343);
nand U8500 (N_8500,N_7305,N_6701);
nand U8501 (N_8501,N_6188,N_6316);
and U8502 (N_8502,N_6900,N_7147);
xor U8503 (N_8503,N_6718,N_7049);
nor U8504 (N_8504,N_7327,N_6946);
nand U8505 (N_8505,N_7028,N_6043);
and U8506 (N_8506,N_7071,N_7486);
and U8507 (N_8507,N_6822,N_6379);
xnor U8508 (N_8508,N_6490,N_6558);
and U8509 (N_8509,N_6257,N_6490);
or U8510 (N_8510,N_6432,N_6403);
and U8511 (N_8511,N_6608,N_6386);
and U8512 (N_8512,N_6775,N_6782);
nand U8513 (N_8513,N_6514,N_7381);
or U8514 (N_8514,N_6390,N_6608);
xnor U8515 (N_8515,N_6015,N_6690);
and U8516 (N_8516,N_7008,N_6233);
nand U8517 (N_8517,N_7237,N_6842);
nor U8518 (N_8518,N_6815,N_6742);
xor U8519 (N_8519,N_6109,N_6423);
or U8520 (N_8520,N_7365,N_6616);
nand U8521 (N_8521,N_6888,N_7106);
nand U8522 (N_8522,N_7032,N_6950);
nand U8523 (N_8523,N_7191,N_7284);
xor U8524 (N_8524,N_6013,N_6918);
nand U8525 (N_8525,N_6635,N_6948);
or U8526 (N_8526,N_6157,N_6584);
nand U8527 (N_8527,N_6800,N_6878);
nand U8528 (N_8528,N_6024,N_6565);
nor U8529 (N_8529,N_6075,N_6461);
xor U8530 (N_8530,N_6833,N_6622);
xor U8531 (N_8531,N_7213,N_6982);
nand U8532 (N_8532,N_6040,N_7309);
or U8533 (N_8533,N_6333,N_6562);
and U8534 (N_8534,N_6547,N_7230);
nor U8535 (N_8535,N_6583,N_6340);
or U8536 (N_8536,N_7280,N_6990);
and U8537 (N_8537,N_6198,N_7011);
xnor U8538 (N_8538,N_7473,N_6841);
and U8539 (N_8539,N_6899,N_6953);
nand U8540 (N_8540,N_6722,N_6924);
nand U8541 (N_8541,N_7418,N_7195);
nor U8542 (N_8542,N_6827,N_6805);
or U8543 (N_8543,N_6729,N_7310);
or U8544 (N_8544,N_6343,N_6349);
xnor U8545 (N_8545,N_6351,N_6850);
nand U8546 (N_8546,N_7089,N_6595);
and U8547 (N_8547,N_6884,N_6506);
and U8548 (N_8548,N_6684,N_7020);
xnor U8549 (N_8549,N_6768,N_7441);
nor U8550 (N_8550,N_7263,N_6220);
nand U8551 (N_8551,N_6354,N_6122);
or U8552 (N_8552,N_6716,N_7247);
nor U8553 (N_8553,N_6578,N_7140);
nor U8554 (N_8554,N_6131,N_6704);
and U8555 (N_8555,N_6889,N_7294);
and U8556 (N_8556,N_7342,N_6527);
nor U8557 (N_8557,N_6337,N_7406);
and U8558 (N_8558,N_7096,N_6138);
or U8559 (N_8559,N_6441,N_6613);
xor U8560 (N_8560,N_6514,N_7459);
or U8561 (N_8561,N_7311,N_6137);
and U8562 (N_8562,N_6674,N_7473);
xor U8563 (N_8563,N_7179,N_7284);
or U8564 (N_8564,N_6719,N_7395);
and U8565 (N_8565,N_7346,N_6225);
and U8566 (N_8566,N_7341,N_6986);
or U8567 (N_8567,N_7302,N_6220);
and U8568 (N_8568,N_6017,N_6757);
nor U8569 (N_8569,N_6570,N_7181);
xnor U8570 (N_8570,N_6339,N_6954);
xnor U8571 (N_8571,N_6250,N_7213);
nand U8572 (N_8572,N_7036,N_6296);
and U8573 (N_8573,N_6881,N_7496);
nand U8574 (N_8574,N_7057,N_7399);
and U8575 (N_8575,N_7478,N_6201);
xnor U8576 (N_8576,N_6944,N_7477);
xnor U8577 (N_8577,N_7300,N_7099);
nand U8578 (N_8578,N_7496,N_7452);
or U8579 (N_8579,N_7108,N_7328);
and U8580 (N_8580,N_7005,N_6075);
xor U8581 (N_8581,N_7045,N_7303);
nor U8582 (N_8582,N_6719,N_6063);
and U8583 (N_8583,N_7152,N_6464);
xor U8584 (N_8584,N_7401,N_6690);
nor U8585 (N_8585,N_6547,N_6725);
nor U8586 (N_8586,N_6500,N_7415);
nor U8587 (N_8587,N_6403,N_6035);
xnor U8588 (N_8588,N_7321,N_6052);
xor U8589 (N_8589,N_6752,N_6316);
nand U8590 (N_8590,N_6172,N_7344);
or U8591 (N_8591,N_6402,N_6416);
or U8592 (N_8592,N_6491,N_6999);
nor U8593 (N_8593,N_7315,N_7358);
nand U8594 (N_8594,N_6357,N_7370);
xnor U8595 (N_8595,N_7005,N_7173);
nand U8596 (N_8596,N_6055,N_6475);
nor U8597 (N_8597,N_6052,N_6061);
nor U8598 (N_8598,N_6513,N_6485);
and U8599 (N_8599,N_6377,N_6651);
nand U8600 (N_8600,N_6058,N_6609);
nor U8601 (N_8601,N_7307,N_6987);
or U8602 (N_8602,N_6585,N_6269);
nand U8603 (N_8603,N_6858,N_7397);
nand U8604 (N_8604,N_6723,N_6899);
nand U8605 (N_8605,N_7464,N_7468);
nor U8606 (N_8606,N_7036,N_6673);
nand U8607 (N_8607,N_6528,N_6883);
xor U8608 (N_8608,N_6978,N_6579);
nand U8609 (N_8609,N_7449,N_6833);
and U8610 (N_8610,N_6692,N_7147);
nor U8611 (N_8611,N_6337,N_6016);
and U8612 (N_8612,N_7119,N_6135);
and U8613 (N_8613,N_6919,N_6426);
or U8614 (N_8614,N_7045,N_6891);
or U8615 (N_8615,N_6915,N_6051);
or U8616 (N_8616,N_7020,N_6697);
nor U8617 (N_8617,N_7161,N_6542);
and U8618 (N_8618,N_6219,N_6447);
nand U8619 (N_8619,N_6057,N_7195);
and U8620 (N_8620,N_6187,N_6359);
and U8621 (N_8621,N_6176,N_6904);
nand U8622 (N_8622,N_7053,N_6986);
nor U8623 (N_8623,N_6328,N_6593);
xnor U8624 (N_8624,N_7061,N_6388);
nand U8625 (N_8625,N_6336,N_7143);
nor U8626 (N_8626,N_6790,N_6514);
xor U8627 (N_8627,N_7376,N_6427);
or U8628 (N_8628,N_6583,N_6568);
nand U8629 (N_8629,N_7236,N_6195);
nor U8630 (N_8630,N_6606,N_7033);
and U8631 (N_8631,N_6181,N_6071);
nor U8632 (N_8632,N_7007,N_6660);
or U8633 (N_8633,N_7490,N_7456);
xor U8634 (N_8634,N_6531,N_6013);
xor U8635 (N_8635,N_7053,N_6153);
and U8636 (N_8636,N_6538,N_7138);
or U8637 (N_8637,N_6881,N_6232);
nor U8638 (N_8638,N_7028,N_7090);
nand U8639 (N_8639,N_7213,N_6654);
xnor U8640 (N_8640,N_6424,N_6809);
and U8641 (N_8641,N_7494,N_7061);
xnor U8642 (N_8642,N_7080,N_6589);
nand U8643 (N_8643,N_6951,N_7126);
nor U8644 (N_8644,N_6615,N_6418);
or U8645 (N_8645,N_6236,N_6802);
nor U8646 (N_8646,N_6885,N_7402);
nor U8647 (N_8647,N_6802,N_6374);
nand U8648 (N_8648,N_6318,N_7485);
nand U8649 (N_8649,N_6725,N_6645);
and U8650 (N_8650,N_6857,N_7457);
and U8651 (N_8651,N_7152,N_6982);
or U8652 (N_8652,N_7203,N_6421);
nand U8653 (N_8653,N_7001,N_6460);
xnor U8654 (N_8654,N_7285,N_6991);
nor U8655 (N_8655,N_7166,N_7378);
nand U8656 (N_8656,N_6365,N_7489);
or U8657 (N_8657,N_7133,N_6557);
nor U8658 (N_8658,N_6065,N_6472);
xnor U8659 (N_8659,N_7170,N_7019);
and U8660 (N_8660,N_7287,N_7179);
nor U8661 (N_8661,N_6359,N_6205);
nand U8662 (N_8662,N_6048,N_7006);
and U8663 (N_8663,N_6936,N_6394);
or U8664 (N_8664,N_6481,N_6559);
or U8665 (N_8665,N_6532,N_6884);
xnor U8666 (N_8666,N_6653,N_6262);
or U8667 (N_8667,N_6726,N_6613);
and U8668 (N_8668,N_7181,N_6521);
and U8669 (N_8669,N_6386,N_6527);
or U8670 (N_8670,N_6458,N_6622);
or U8671 (N_8671,N_7005,N_6748);
xor U8672 (N_8672,N_6361,N_6441);
xor U8673 (N_8673,N_6242,N_7083);
nand U8674 (N_8674,N_6517,N_7390);
and U8675 (N_8675,N_7498,N_6701);
xnor U8676 (N_8676,N_6835,N_7346);
nor U8677 (N_8677,N_6901,N_6938);
xor U8678 (N_8678,N_6490,N_7242);
or U8679 (N_8679,N_6410,N_6388);
and U8680 (N_8680,N_6893,N_6089);
or U8681 (N_8681,N_6969,N_6385);
and U8682 (N_8682,N_7471,N_6361);
nor U8683 (N_8683,N_6325,N_7355);
or U8684 (N_8684,N_6038,N_6978);
or U8685 (N_8685,N_6807,N_6382);
and U8686 (N_8686,N_6471,N_6084);
and U8687 (N_8687,N_7461,N_6415);
or U8688 (N_8688,N_6135,N_7370);
nand U8689 (N_8689,N_6887,N_6546);
xnor U8690 (N_8690,N_6430,N_7190);
xor U8691 (N_8691,N_6865,N_6978);
or U8692 (N_8692,N_6158,N_6224);
nand U8693 (N_8693,N_6198,N_6667);
nand U8694 (N_8694,N_7325,N_6960);
xnor U8695 (N_8695,N_7409,N_6957);
nand U8696 (N_8696,N_6645,N_6583);
and U8697 (N_8697,N_6343,N_6173);
nand U8698 (N_8698,N_6440,N_7130);
nand U8699 (N_8699,N_6382,N_7452);
nor U8700 (N_8700,N_7095,N_6934);
or U8701 (N_8701,N_7341,N_6319);
and U8702 (N_8702,N_7483,N_7311);
nor U8703 (N_8703,N_6932,N_6546);
nor U8704 (N_8704,N_7143,N_6497);
xor U8705 (N_8705,N_6496,N_6833);
nand U8706 (N_8706,N_6504,N_6986);
and U8707 (N_8707,N_6260,N_6316);
or U8708 (N_8708,N_6682,N_7287);
or U8709 (N_8709,N_6571,N_6103);
and U8710 (N_8710,N_6421,N_6381);
nand U8711 (N_8711,N_7064,N_6188);
xor U8712 (N_8712,N_6851,N_6835);
and U8713 (N_8713,N_6619,N_7132);
xnor U8714 (N_8714,N_6911,N_7372);
nor U8715 (N_8715,N_6407,N_6888);
nor U8716 (N_8716,N_6618,N_6411);
nor U8717 (N_8717,N_6158,N_6531);
and U8718 (N_8718,N_6831,N_6334);
and U8719 (N_8719,N_7268,N_6921);
nand U8720 (N_8720,N_6868,N_6098);
nand U8721 (N_8721,N_7247,N_6935);
xnor U8722 (N_8722,N_6866,N_6315);
nand U8723 (N_8723,N_6632,N_6373);
or U8724 (N_8724,N_6789,N_6020);
nand U8725 (N_8725,N_6217,N_6375);
nor U8726 (N_8726,N_7495,N_6401);
nand U8727 (N_8727,N_6329,N_7445);
nor U8728 (N_8728,N_6897,N_6581);
and U8729 (N_8729,N_7135,N_6890);
or U8730 (N_8730,N_6512,N_7259);
or U8731 (N_8731,N_7058,N_6688);
and U8732 (N_8732,N_7118,N_6413);
nand U8733 (N_8733,N_6606,N_6030);
xnor U8734 (N_8734,N_7041,N_7491);
nand U8735 (N_8735,N_6154,N_6239);
nor U8736 (N_8736,N_7484,N_7320);
nand U8737 (N_8737,N_7149,N_7061);
nor U8738 (N_8738,N_7446,N_7361);
nor U8739 (N_8739,N_7283,N_6875);
nand U8740 (N_8740,N_7125,N_6408);
or U8741 (N_8741,N_6938,N_6120);
nand U8742 (N_8742,N_7310,N_6164);
and U8743 (N_8743,N_6060,N_6290);
and U8744 (N_8744,N_7185,N_6049);
nor U8745 (N_8745,N_7003,N_6342);
xor U8746 (N_8746,N_7257,N_6500);
and U8747 (N_8747,N_6781,N_7125);
or U8748 (N_8748,N_6102,N_6278);
or U8749 (N_8749,N_7100,N_6783);
nor U8750 (N_8750,N_6416,N_6031);
nand U8751 (N_8751,N_6572,N_6308);
nand U8752 (N_8752,N_6872,N_6493);
xor U8753 (N_8753,N_6726,N_7046);
nand U8754 (N_8754,N_6825,N_7286);
nand U8755 (N_8755,N_6217,N_6120);
or U8756 (N_8756,N_6009,N_6362);
nor U8757 (N_8757,N_6758,N_6322);
xor U8758 (N_8758,N_6461,N_6070);
nand U8759 (N_8759,N_6072,N_6194);
or U8760 (N_8760,N_7008,N_6201);
xnor U8761 (N_8761,N_6186,N_6729);
nor U8762 (N_8762,N_6397,N_7173);
nand U8763 (N_8763,N_6123,N_6561);
xor U8764 (N_8764,N_7128,N_6736);
xnor U8765 (N_8765,N_7353,N_6338);
nand U8766 (N_8766,N_6842,N_6002);
nand U8767 (N_8767,N_6487,N_7129);
nand U8768 (N_8768,N_6239,N_6845);
nor U8769 (N_8769,N_6328,N_6974);
and U8770 (N_8770,N_6695,N_7344);
and U8771 (N_8771,N_6041,N_6760);
nand U8772 (N_8772,N_7140,N_6935);
nand U8773 (N_8773,N_6549,N_6612);
xor U8774 (N_8774,N_6583,N_7064);
and U8775 (N_8775,N_6802,N_6847);
xor U8776 (N_8776,N_6603,N_6436);
xnor U8777 (N_8777,N_7335,N_6877);
nor U8778 (N_8778,N_6561,N_7321);
or U8779 (N_8779,N_6693,N_6105);
nor U8780 (N_8780,N_6064,N_6696);
and U8781 (N_8781,N_7137,N_6324);
nor U8782 (N_8782,N_6621,N_7394);
nand U8783 (N_8783,N_6356,N_7466);
and U8784 (N_8784,N_7305,N_6883);
nand U8785 (N_8785,N_7072,N_6983);
nand U8786 (N_8786,N_6097,N_6019);
nor U8787 (N_8787,N_6237,N_6890);
or U8788 (N_8788,N_7412,N_7469);
and U8789 (N_8789,N_6781,N_6589);
xor U8790 (N_8790,N_6672,N_7127);
or U8791 (N_8791,N_7310,N_7023);
xnor U8792 (N_8792,N_6225,N_7345);
nand U8793 (N_8793,N_7448,N_7003);
xnor U8794 (N_8794,N_7413,N_6863);
xnor U8795 (N_8795,N_6187,N_6412);
or U8796 (N_8796,N_6506,N_6981);
nor U8797 (N_8797,N_6471,N_7386);
xnor U8798 (N_8798,N_7014,N_6346);
nor U8799 (N_8799,N_6780,N_6432);
or U8800 (N_8800,N_6198,N_6457);
nor U8801 (N_8801,N_6157,N_7166);
nand U8802 (N_8802,N_6783,N_6557);
nor U8803 (N_8803,N_7461,N_6778);
xnor U8804 (N_8804,N_6989,N_6933);
nor U8805 (N_8805,N_7326,N_7034);
xor U8806 (N_8806,N_6262,N_6635);
and U8807 (N_8807,N_6939,N_6041);
xnor U8808 (N_8808,N_6008,N_6697);
and U8809 (N_8809,N_6009,N_6980);
nand U8810 (N_8810,N_6287,N_7245);
or U8811 (N_8811,N_7364,N_7395);
nor U8812 (N_8812,N_7293,N_6912);
nor U8813 (N_8813,N_7328,N_6200);
or U8814 (N_8814,N_7222,N_6231);
and U8815 (N_8815,N_7000,N_7315);
nand U8816 (N_8816,N_7025,N_6070);
and U8817 (N_8817,N_6322,N_6267);
nor U8818 (N_8818,N_6691,N_6160);
or U8819 (N_8819,N_7244,N_6237);
nand U8820 (N_8820,N_6228,N_6305);
or U8821 (N_8821,N_6200,N_6920);
and U8822 (N_8822,N_7424,N_7000);
xor U8823 (N_8823,N_7031,N_6774);
xnor U8824 (N_8824,N_6372,N_6839);
or U8825 (N_8825,N_7386,N_7100);
nor U8826 (N_8826,N_6684,N_6283);
and U8827 (N_8827,N_6119,N_7253);
nand U8828 (N_8828,N_7179,N_7426);
or U8829 (N_8829,N_6272,N_6258);
xnor U8830 (N_8830,N_7212,N_6761);
xor U8831 (N_8831,N_7048,N_7070);
nand U8832 (N_8832,N_6426,N_7390);
nor U8833 (N_8833,N_6546,N_6857);
xor U8834 (N_8834,N_6470,N_6368);
or U8835 (N_8835,N_6440,N_7253);
nor U8836 (N_8836,N_7096,N_6798);
nand U8837 (N_8837,N_6399,N_6390);
nor U8838 (N_8838,N_6248,N_7197);
or U8839 (N_8839,N_6271,N_7041);
or U8840 (N_8840,N_6371,N_7334);
or U8841 (N_8841,N_6256,N_6457);
and U8842 (N_8842,N_6757,N_6916);
and U8843 (N_8843,N_6823,N_7405);
nor U8844 (N_8844,N_6697,N_6103);
nor U8845 (N_8845,N_6676,N_6320);
nor U8846 (N_8846,N_7472,N_6983);
nor U8847 (N_8847,N_7352,N_7136);
nand U8848 (N_8848,N_6634,N_6987);
and U8849 (N_8849,N_6786,N_6757);
or U8850 (N_8850,N_6233,N_7465);
xnor U8851 (N_8851,N_6425,N_6307);
nand U8852 (N_8852,N_6818,N_6542);
xor U8853 (N_8853,N_6796,N_7107);
or U8854 (N_8854,N_6057,N_7083);
xnor U8855 (N_8855,N_6225,N_6364);
nand U8856 (N_8856,N_6003,N_7365);
xor U8857 (N_8857,N_6108,N_7311);
or U8858 (N_8858,N_6018,N_7406);
and U8859 (N_8859,N_7105,N_6371);
nand U8860 (N_8860,N_7023,N_6265);
nand U8861 (N_8861,N_6711,N_6695);
xnor U8862 (N_8862,N_6405,N_7444);
nand U8863 (N_8863,N_6022,N_6453);
nand U8864 (N_8864,N_6518,N_7071);
nand U8865 (N_8865,N_7258,N_6550);
nand U8866 (N_8866,N_6201,N_6914);
nand U8867 (N_8867,N_7081,N_6515);
xor U8868 (N_8868,N_6632,N_6488);
nor U8869 (N_8869,N_6174,N_6226);
xor U8870 (N_8870,N_6590,N_7253);
and U8871 (N_8871,N_6585,N_6865);
xnor U8872 (N_8872,N_7081,N_7451);
or U8873 (N_8873,N_6659,N_6194);
xor U8874 (N_8874,N_7425,N_6062);
and U8875 (N_8875,N_7364,N_6402);
or U8876 (N_8876,N_7201,N_6501);
nand U8877 (N_8877,N_6121,N_6969);
nor U8878 (N_8878,N_6056,N_6011);
and U8879 (N_8879,N_7115,N_6635);
or U8880 (N_8880,N_6763,N_6548);
and U8881 (N_8881,N_7212,N_7400);
nor U8882 (N_8882,N_6201,N_6447);
nor U8883 (N_8883,N_6704,N_7470);
or U8884 (N_8884,N_6302,N_6733);
xnor U8885 (N_8885,N_7271,N_6114);
or U8886 (N_8886,N_6186,N_7021);
nand U8887 (N_8887,N_6649,N_7477);
or U8888 (N_8888,N_7042,N_7161);
nand U8889 (N_8889,N_7000,N_7094);
or U8890 (N_8890,N_6521,N_6935);
or U8891 (N_8891,N_6310,N_7424);
or U8892 (N_8892,N_7238,N_7306);
nor U8893 (N_8893,N_7068,N_6770);
xnor U8894 (N_8894,N_6157,N_7085);
or U8895 (N_8895,N_6377,N_6867);
or U8896 (N_8896,N_6719,N_7049);
and U8897 (N_8897,N_6167,N_6021);
nor U8898 (N_8898,N_6296,N_6536);
nand U8899 (N_8899,N_6519,N_7287);
xnor U8900 (N_8900,N_7055,N_7204);
nand U8901 (N_8901,N_7349,N_7100);
nor U8902 (N_8902,N_6464,N_6826);
nand U8903 (N_8903,N_6861,N_6047);
and U8904 (N_8904,N_7059,N_7377);
or U8905 (N_8905,N_6752,N_7296);
and U8906 (N_8906,N_6848,N_6602);
nand U8907 (N_8907,N_6427,N_6623);
nand U8908 (N_8908,N_7490,N_6791);
nor U8909 (N_8909,N_6416,N_7306);
or U8910 (N_8910,N_7000,N_6253);
or U8911 (N_8911,N_6550,N_6602);
and U8912 (N_8912,N_7248,N_6447);
nand U8913 (N_8913,N_6204,N_6386);
and U8914 (N_8914,N_7401,N_6646);
or U8915 (N_8915,N_7120,N_7134);
or U8916 (N_8916,N_7201,N_6732);
or U8917 (N_8917,N_6606,N_6116);
nand U8918 (N_8918,N_6186,N_6877);
xnor U8919 (N_8919,N_6796,N_7162);
nor U8920 (N_8920,N_6065,N_7115);
nor U8921 (N_8921,N_6117,N_7355);
nand U8922 (N_8922,N_6156,N_6123);
nand U8923 (N_8923,N_6924,N_7197);
nor U8924 (N_8924,N_7266,N_6353);
or U8925 (N_8925,N_6124,N_6218);
nand U8926 (N_8926,N_6142,N_7262);
or U8927 (N_8927,N_7326,N_7104);
xnor U8928 (N_8928,N_6344,N_7443);
and U8929 (N_8929,N_6304,N_7302);
or U8930 (N_8930,N_6673,N_6389);
xor U8931 (N_8931,N_6511,N_6162);
and U8932 (N_8932,N_6216,N_6060);
and U8933 (N_8933,N_7156,N_7494);
and U8934 (N_8934,N_6059,N_6596);
nand U8935 (N_8935,N_6304,N_6818);
xor U8936 (N_8936,N_6478,N_6243);
nand U8937 (N_8937,N_7007,N_6580);
nor U8938 (N_8938,N_6821,N_7472);
xnor U8939 (N_8939,N_7025,N_6137);
or U8940 (N_8940,N_6194,N_7382);
nand U8941 (N_8941,N_7392,N_6377);
xnor U8942 (N_8942,N_6500,N_6383);
nand U8943 (N_8943,N_6871,N_7455);
xor U8944 (N_8944,N_6008,N_7148);
xor U8945 (N_8945,N_6208,N_6307);
nand U8946 (N_8946,N_7012,N_6518);
nor U8947 (N_8947,N_6719,N_7191);
xnor U8948 (N_8948,N_6460,N_7280);
and U8949 (N_8949,N_6695,N_7392);
and U8950 (N_8950,N_6555,N_6621);
and U8951 (N_8951,N_6702,N_6005);
nand U8952 (N_8952,N_7020,N_6633);
and U8953 (N_8953,N_6737,N_6211);
xnor U8954 (N_8954,N_7080,N_7293);
nor U8955 (N_8955,N_7220,N_7029);
xnor U8956 (N_8956,N_7456,N_6059);
and U8957 (N_8957,N_6652,N_6408);
nand U8958 (N_8958,N_7424,N_7204);
or U8959 (N_8959,N_6340,N_7041);
nor U8960 (N_8960,N_6277,N_7109);
nor U8961 (N_8961,N_7105,N_7110);
nand U8962 (N_8962,N_6734,N_7154);
nor U8963 (N_8963,N_6186,N_6234);
or U8964 (N_8964,N_6233,N_6064);
xor U8965 (N_8965,N_7211,N_6022);
nand U8966 (N_8966,N_7373,N_6473);
nor U8967 (N_8967,N_6080,N_7293);
or U8968 (N_8968,N_6880,N_7227);
or U8969 (N_8969,N_6884,N_7104);
or U8970 (N_8970,N_6023,N_6779);
xor U8971 (N_8971,N_6013,N_6846);
and U8972 (N_8972,N_7223,N_7162);
and U8973 (N_8973,N_7169,N_6482);
nand U8974 (N_8974,N_6041,N_6837);
nor U8975 (N_8975,N_6586,N_7491);
nor U8976 (N_8976,N_6234,N_7428);
nor U8977 (N_8977,N_6006,N_6259);
nand U8978 (N_8978,N_7285,N_6295);
xnor U8979 (N_8979,N_6293,N_7250);
or U8980 (N_8980,N_6460,N_6079);
nor U8981 (N_8981,N_6341,N_6773);
nor U8982 (N_8982,N_6601,N_6967);
xnor U8983 (N_8983,N_6414,N_6129);
or U8984 (N_8984,N_7267,N_7024);
nor U8985 (N_8985,N_6213,N_7152);
or U8986 (N_8986,N_6275,N_6523);
nand U8987 (N_8987,N_6759,N_6032);
nand U8988 (N_8988,N_7089,N_6558);
nor U8989 (N_8989,N_7046,N_6794);
nor U8990 (N_8990,N_7025,N_7320);
or U8991 (N_8991,N_6938,N_6065);
nand U8992 (N_8992,N_6693,N_7402);
xor U8993 (N_8993,N_6650,N_6198);
nor U8994 (N_8994,N_6191,N_6235);
nand U8995 (N_8995,N_7387,N_7331);
xor U8996 (N_8996,N_7321,N_6143);
xor U8997 (N_8997,N_7065,N_6799);
or U8998 (N_8998,N_6577,N_6788);
or U8999 (N_8999,N_7024,N_6314);
nand U9000 (N_9000,N_8721,N_8060);
xnor U9001 (N_9001,N_8379,N_8324);
and U9002 (N_9002,N_7740,N_8053);
nor U9003 (N_9003,N_7515,N_8040);
xnor U9004 (N_9004,N_7888,N_8454);
nand U9005 (N_9005,N_7542,N_8984);
nand U9006 (N_9006,N_8108,N_7937);
and U9007 (N_9007,N_8847,N_8240);
xnor U9008 (N_9008,N_8153,N_8348);
xor U9009 (N_9009,N_8321,N_8876);
xnor U9010 (N_9010,N_8026,N_8238);
or U9011 (N_9011,N_8794,N_8043);
and U9012 (N_9012,N_8411,N_8129);
or U9013 (N_9013,N_7609,N_8436);
nor U9014 (N_9014,N_7640,N_8112);
nor U9015 (N_9015,N_8715,N_8091);
and U9016 (N_9016,N_8466,N_8550);
nor U9017 (N_9017,N_8219,N_7772);
and U9018 (N_9018,N_8848,N_8490);
nand U9019 (N_9019,N_7842,N_7755);
xor U9020 (N_9020,N_7719,N_8966);
and U9021 (N_9021,N_8271,N_8549);
and U9022 (N_9022,N_7853,N_8662);
nor U9023 (N_9023,N_7865,N_8429);
and U9024 (N_9024,N_7819,N_8789);
nand U9025 (N_9025,N_8113,N_8941);
nor U9026 (N_9026,N_7926,N_7899);
or U9027 (N_9027,N_8004,N_8872);
nand U9028 (N_9028,N_8650,N_8840);
or U9029 (N_9029,N_8774,N_8824);
and U9030 (N_9030,N_7827,N_7783);
xor U9031 (N_9031,N_7681,N_8335);
nor U9032 (N_9032,N_8388,N_8798);
nand U9033 (N_9033,N_8455,N_8187);
and U9034 (N_9034,N_7934,N_8277);
xor U9035 (N_9035,N_8709,N_8139);
xnor U9036 (N_9036,N_8969,N_8297);
nor U9037 (N_9037,N_7919,N_8780);
xor U9038 (N_9038,N_8904,N_8703);
nor U9039 (N_9039,N_8796,N_7737);
nand U9040 (N_9040,N_7773,N_8110);
and U9041 (N_9041,N_8536,N_7929);
nor U9042 (N_9042,N_7803,N_7547);
nor U9043 (N_9043,N_8916,N_8667);
nand U9044 (N_9044,N_8276,N_7968);
xor U9045 (N_9045,N_8836,N_8548);
and U9046 (N_9046,N_8125,N_7675);
or U9047 (N_9047,N_8989,N_8396);
nand U9048 (N_9048,N_7702,N_7788);
nand U9049 (N_9049,N_8417,N_8172);
or U9050 (N_9050,N_8878,N_8671);
nand U9051 (N_9051,N_8222,N_8855);
or U9052 (N_9052,N_8821,N_8502);
or U9053 (N_9053,N_7916,N_7875);
and U9054 (N_9054,N_8543,N_8033);
or U9055 (N_9055,N_8259,N_8556);
xor U9056 (N_9056,N_7859,N_8733);
nand U9057 (N_9057,N_8516,N_8022);
or U9058 (N_9058,N_7513,N_8460);
xor U9059 (N_9059,N_8024,N_7603);
nand U9060 (N_9060,N_8037,N_8408);
nor U9061 (N_9061,N_8511,N_8001);
nand U9062 (N_9062,N_8771,N_8599);
nand U9063 (N_9063,N_7543,N_7502);
or U9064 (N_9064,N_8155,N_8235);
nor U9065 (N_9065,N_7801,N_8608);
and U9066 (N_9066,N_7684,N_8575);
and U9067 (N_9067,N_8160,N_7596);
xnor U9068 (N_9068,N_8860,N_7594);
xnor U9069 (N_9069,N_7568,N_8227);
nand U9070 (N_9070,N_8712,N_8293);
or U9071 (N_9071,N_7832,N_8882);
xor U9072 (N_9072,N_8370,N_8631);
and U9073 (N_9073,N_7687,N_8369);
or U9074 (N_9074,N_7703,N_8143);
nor U9075 (N_9075,N_8165,N_8098);
xor U9076 (N_9076,N_8717,N_7650);
and U9077 (N_9077,N_7501,N_8419);
and U9078 (N_9078,N_8497,N_7860);
xnor U9079 (N_9079,N_7733,N_8641);
xor U9080 (N_9080,N_8327,N_8784);
nor U9081 (N_9081,N_8507,N_7995);
or U9082 (N_9082,N_8623,N_8723);
and U9083 (N_9083,N_8152,N_7619);
xnor U9084 (N_9084,N_8158,N_8869);
nand U9085 (N_9085,N_8530,N_8011);
xnor U9086 (N_9086,N_8965,N_7845);
nand U9087 (N_9087,N_8504,N_7994);
nand U9088 (N_9088,N_8072,N_8978);
nand U9089 (N_9089,N_8206,N_8194);
and U9090 (N_9090,N_8842,N_8047);
or U9091 (N_9091,N_8131,N_8318);
and U9092 (N_9092,N_8215,N_8216);
nor U9093 (N_9093,N_7572,N_7894);
xnor U9094 (N_9094,N_7586,N_8565);
nand U9095 (N_9095,N_8724,N_7563);
and U9096 (N_9096,N_8957,N_8613);
xnor U9097 (N_9097,N_8870,N_7953);
or U9098 (N_9098,N_8330,N_7711);
xnor U9099 (N_9099,N_8791,N_7779);
xor U9100 (N_9100,N_8517,N_7727);
xnor U9101 (N_9101,N_8693,N_7777);
nand U9102 (N_9102,N_7752,N_8603);
nand U9103 (N_9103,N_8677,N_8170);
or U9104 (N_9104,N_7597,N_7565);
or U9105 (N_9105,N_7508,N_8479);
and U9106 (N_9106,N_8820,N_8000);
xor U9107 (N_9107,N_8220,N_7536);
or U9108 (N_9108,N_8336,N_8583);
xnor U9109 (N_9109,N_8175,N_8415);
nor U9110 (N_9110,N_8493,N_7993);
or U9111 (N_9111,N_8880,N_7790);
and U9112 (N_9112,N_7530,N_8384);
nor U9113 (N_9113,N_8156,N_7570);
or U9114 (N_9114,N_8101,N_8624);
and U9115 (N_9115,N_8768,N_8298);
xor U9116 (N_9116,N_7511,N_8439);
and U9117 (N_9117,N_8078,N_8185);
nand U9118 (N_9118,N_8616,N_8264);
nor U9119 (N_9119,N_7722,N_8779);
and U9120 (N_9120,N_7524,N_7754);
nor U9121 (N_9121,N_7954,N_8280);
and U9122 (N_9122,N_7841,N_7961);
or U9123 (N_9123,N_7900,N_7742);
or U9124 (N_9124,N_8403,N_8023);
xnor U9125 (N_9125,N_8105,N_8376);
and U9126 (N_9126,N_7504,N_8122);
or U9127 (N_9127,N_8312,N_8056);
xnor U9128 (N_9128,N_8405,N_8900);
and U9129 (N_9129,N_8955,N_7784);
nand U9130 (N_9130,N_8992,N_8529);
and U9131 (N_9131,N_8469,N_8601);
and U9132 (N_9132,N_7720,N_8050);
xor U9133 (N_9133,N_7962,N_8862);
nand U9134 (N_9134,N_8115,N_7991);
nor U9135 (N_9135,N_7880,N_8804);
nand U9136 (N_9136,N_8982,N_8289);
xnor U9137 (N_9137,N_8036,N_7904);
and U9138 (N_9138,N_8811,N_8903);
and U9139 (N_9139,N_8308,N_7840);
nand U9140 (N_9140,N_8873,N_8964);
xor U9141 (N_9141,N_8427,N_7906);
nor U9142 (N_9142,N_8250,N_8267);
nand U9143 (N_9143,N_7761,N_8672);
or U9144 (N_9144,N_8897,N_7966);
nor U9145 (N_9145,N_7930,N_7855);
and U9146 (N_9146,N_7553,N_8935);
xor U9147 (N_9147,N_7573,N_7802);
nand U9148 (N_9148,N_7863,N_8385);
and U9149 (N_9149,N_8232,N_7647);
or U9150 (N_9150,N_8448,N_7712);
xor U9151 (N_9151,N_8985,N_8559);
nor U9152 (N_9152,N_8598,N_8892);
xnor U9153 (N_9153,N_7695,N_8462);
nand U9154 (N_9154,N_8760,N_7615);
and U9155 (N_9155,N_7918,N_8148);
nand U9156 (N_9156,N_8274,N_8169);
xnor U9157 (N_9157,N_8594,N_8674);
and U9158 (N_9158,N_7861,N_7560);
xnor U9159 (N_9159,N_8857,N_8372);
or U9160 (N_9160,N_8781,N_8423);
or U9161 (N_9161,N_8934,N_7963);
or U9162 (N_9162,N_7938,N_8576);
and U9163 (N_9163,N_7598,N_8525);
nor U9164 (N_9164,N_7810,N_8640);
xor U9165 (N_9165,N_7555,N_8795);
xor U9166 (N_9166,N_7756,N_8118);
nand U9167 (N_9167,N_8828,N_8633);
or U9168 (N_9168,N_7591,N_7662);
or U9169 (N_9169,N_8629,N_7868);
or U9170 (N_9170,N_8407,N_8426);
xnor U9171 (N_9171,N_8952,N_8763);
or U9172 (N_9172,N_8881,N_8015);
nor U9173 (N_9173,N_8099,N_8726);
and U9174 (N_9174,N_8279,N_7655);
nor U9175 (N_9175,N_7723,N_8109);
xnor U9176 (N_9176,N_7716,N_8266);
nor U9177 (N_9177,N_8545,N_7884);
xor U9178 (N_9178,N_8573,N_8496);
xnor U9179 (N_9179,N_8694,N_7750);
nor U9180 (N_9180,N_8681,N_8838);
nor U9181 (N_9181,N_7920,N_7585);
xor U9182 (N_9182,N_8885,N_8670);
xor U9183 (N_9183,N_7799,N_7935);
nor U9184 (N_9184,N_7562,N_7521);
and U9185 (N_9185,N_8807,N_8644);
or U9186 (N_9186,N_8132,N_7660);
or U9187 (N_9187,N_8533,N_7520);
nor U9188 (N_9188,N_8494,N_8485);
xor U9189 (N_9189,N_8766,N_8213);
nand U9190 (N_9190,N_7985,N_8449);
xor U9191 (N_9191,N_7793,N_8765);
nor U9192 (N_9192,N_8962,N_8665);
xor U9193 (N_9193,N_7569,N_8104);
or U9194 (N_9194,N_8702,N_8815);
and U9195 (N_9195,N_8371,N_7898);
and U9196 (N_9196,N_8199,N_8930);
or U9197 (N_9197,N_8571,N_8532);
and U9198 (N_9198,N_8524,N_7529);
nor U9199 (N_9199,N_8928,N_7850);
and U9200 (N_9200,N_8970,N_8566);
nand U9201 (N_9201,N_8755,N_8757);
nor U9202 (N_9202,N_7951,N_7658);
and U9203 (N_9203,N_8720,N_8664);
nand U9204 (N_9204,N_7984,N_8179);
or U9205 (N_9205,N_8141,N_8697);
xnor U9206 (N_9206,N_8446,N_7554);
nand U9207 (N_9207,N_8166,N_8950);
nand U9208 (N_9208,N_8711,N_7804);
and U9209 (N_9209,N_7694,N_8741);
or U9210 (N_9210,N_7725,N_7765);
or U9211 (N_9211,N_8863,N_8729);
nand U9212 (N_9212,N_7541,N_8996);
nor U9213 (N_9213,N_8183,N_7908);
and U9214 (N_9214,N_8188,N_8938);
nor U9215 (N_9215,N_8508,N_8925);
xnor U9216 (N_9216,N_8328,N_8245);
and U9217 (N_9217,N_8971,N_7879);
or U9218 (N_9218,N_8444,N_8406);
xor U9219 (N_9219,N_8021,N_8300);
or U9220 (N_9220,N_7972,N_8803);
and U9221 (N_9221,N_7751,N_8636);
xor U9222 (N_9222,N_8753,N_8059);
nand U9223 (N_9223,N_8147,N_8258);
or U9224 (N_9224,N_7843,N_7897);
nor U9225 (N_9225,N_8871,N_8822);
nand U9226 (N_9226,N_7539,N_7673);
and U9227 (N_9227,N_8182,N_8651);
nor U9228 (N_9228,N_8542,N_8630);
nor U9229 (N_9229,N_8195,N_8749);
xnor U9230 (N_9230,N_7924,N_8716);
and U9231 (N_9231,N_7786,N_7805);
xor U9232 (N_9232,N_7815,N_8646);
and U9233 (N_9233,N_8745,N_8910);
and U9234 (N_9234,N_8572,N_8354);
nand U9235 (N_9235,N_8018,N_8177);
nand U9236 (N_9236,N_8577,N_8946);
nor U9237 (N_9237,N_8899,N_8332);
and U9238 (N_9238,N_8605,N_8410);
nand U9239 (N_9239,N_7651,N_8117);
nand U9240 (N_9240,N_8073,N_8120);
xnor U9241 (N_9241,N_7714,N_7915);
xnor U9242 (N_9242,N_7856,N_7693);
xnor U9243 (N_9243,N_7905,N_7821);
and U9244 (N_9244,N_8083,N_8786);
and U9245 (N_9245,N_7545,N_7854);
and U9246 (N_9246,N_7818,N_8189);
or U9247 (N_9247,N_8048,N_8625);
and U9248 (N_9248,N_8588,N_8400);
and U9249 (N_9249,N_8349,N_8224);
nor U9250 (N_9250,N_8116,N_7644);
and U9251 (N_9251,N_8919,N_8019);
or U9252 (N_9252,N_7600,N_8911);
nand U9253 (N_9253,N_8775,N_8247);
and U9254 (N_9254,N_8392,N_8311);
and U9255 (N_9255,N_7576,N_7578);
nand U9256 (N_9256,N_7923,N_7577);
or U9257 (N_9257,N_8002,N_7724);
and U9258 (N_9258,N_7680,N_7770);
or U9259 (N_9259,N_8688,N_8350);
nand U9260 (N_9260,N_7566,N_7838);
xnor U9261 (N_9261,N_7623,N_8812);
nand U9262 (N_9262,N_7606,N_7958);
or U9263 (N_9263,N_8301,N_8802);
nand U9264 (N_9264,N_7528,N_8528);
nand U9265 (N_9265,N_7811,N_8197);
and U9266 (N_9266,N_7901,N_7654);
nand U9267 (N_9267,N_8713,N_7736);
and U9268 (N_9268,N_8217,N_7957);
or U9269 (N_9269,N_7977,N_8339);
or U9270 (N_9270,N_8364,N_7574);
nand U9271 (N_9271,N_8655,N_7685);
nor U9272 (N_9272,N_8866,N_7895);
nand U9273 (N_9273,N_8212,N_8157);
or U9274 (N_9274,N_8676,N_8642);
and U9275 (N_9275,N_8178,N_8431);
nand U9276 (N_9276,N_8558,N_8102);
xor U9277 (N_9277,N_8657,N_7708);
and U9278 (N_9278,N_8069,N_8684);
xnor U9279 (N_9279,N_8704,N_8894);
nor U9280 (N_9280,N_8959,N_8200);
nor U9281 (N_9281,N_8695,N_7605);
and U9282 (N_9282,N_8025,N_8639);
xnor U9283 (N_9283,N_7726,N_8805);
nor U9284 (N_9284,N_7653,N_8288);
xnor U9285 (N_9285,N_8149,N_8028);
nand U9286 (N_9286,N_8397,N_7835);
nor U9287 (N_9287,N_7652,N_7933);
nor U9288 (N_9288,N_8521,N_8399);
xor U9289 (N_9289,N_8334,N_8579);
and U9290 (N_9290,N_8128,N_8981);
xor U9291 (N_9291,N_7999,N_8389);
xnor U9292 (N_9292,N_7877,N_8648);
nand U9293 (N_9293,N_8007,N_8788);
and U9294 (N_9294,N_8140,N_7974);
or U9295 (N_9295,N_8617,N_8658);
or U9296 (N_9296,N_8722,N_8081);
nor U9297 (N_9297,N_8159,N_7707);
nor U9298 (N_9298,N_7557,N_8951);
nor U9299 (N_9299,N_7500,N_8858);
xnor U9300 (N_9300,N_7638,N_8303);
or U9301 (N_9301,N_7980,N_7834);
nand U9302 (N_9302,N_8831,N_7769);
or U9303 (N_9303,N_8647,N_8555);
or U9304 (N_9304,N_8225,N_7925);
xnor U9305 (N_9305,N_8680,N_8489);
and U9306 (N_9306,N_8706,N_7833);
xnor U9307 (N_9307,N_8719,N_8936);
and U9308 (N_9308,N_8239,N_8103);
or U9309 (N_9309,N_8922,N_7849);
nor U9310 (N_9310,N_8174,N_7981);
xnor U9311 (N_9311,N_7886,N_7851);
xnor U9312 (N_9312,N_7857,N_7914);
xor U9313 (N_9313,N_8307,N_7829);
xor U9314 (N_9314,N_8202,N_8736);
or U9315 (N_9315,N_8070,N_7505);
or U9316 (N_9316,N_8510,N_8750);
xnor U9317 (N_9317,N_8086,N_8123);
or U9318 (N_9318,N_7706,N_7697);
nand U9319 (N_9319,N_7814,N_7731);
and U9320 (N_9320,N_8544,N_7670);
nand U9321 (N_9321,N_8320,N_7969);
xnor U9322 (N_9322,N_7964,N_7575);
or U9323 (N_9323,N_8375,N_7602);
nor U9324 (N_9324,N_8012,N_8394);
and U9325 (N_9325,N_8747,N_8531);
and U9326 (N_9326,N_8045,N_8926);
and U9327 (N_9327,N_8538,N_8698);
xor U9328 (N_9328,N_8778,N_8452);
nand U9329 (N_9329,N_8701,N_8346);
xnor U9330 (N_9330,N_7721,N_8825);
and U9331 (N_9331,N_8690,N_7683);
xnor U9332 (N_9332,N_7696,N_8600);
and U9333 (N_9333,N_7639,N_8292);
xnor U9334 (N_9334,N_7518,N_8854);
or U9335 (N_9335,N_8231,N_8470);
nor U9336 (N_9336,N_8203,N_7584);
nand U9337 (N_9337,N_8668,N_8323);
and U9338 (N_9338,N_7688,N_8888);
nand U9339 (N_9339,N_8834,N_8967);
and U9340 (N_9340,N_7910,N_8409);
and U9341 (N_9341,N_7948,N_8357);
nor U9342 (N_9342,N_8835,N_8127);
xnor U9343 (N_9343,N_8972,N_8163);
nor U9344 (N_9344,N_8638,N_8268);
nor U9345 (N_9345,N_8005,N_7635);
or U9346 (N_9346,N_8929,N_8696);
or U9347 (N_9347,N_8463,N_7789);
and U9348 (N_9348,N_8087,N_7656);
xnor U9349 (N_9349,N_7763,N_7766);
xor U9350 (N_9350,N_7713,N_8945);
or U9351 (N_9351,N_7955,N_8198);
xnor U9352 (N_9352,N_8275,N_8746);
nand U9353 (N_9353,N_8171,N_8180);
nor U9354 (N_9354,N_7912,N_8666);
nand U9355 (N_9355,N_8373,N_7676);
nand U9356 (N_9356,N_8865,N_8265);
xnor U9357 (N_9357,N_8580,N_7758);
xor U9358 (N_9358,N_8253,N_8014);
or U9359 (N_9359,N_7990,N_7588);
nor U9360 (N_9360,N_7873,N_7881);
or U9361 (N_9361,N_8682,N_8578);
xor U9362 (N_9362,N_8679,N_8793);
nor U9363 (N_9363,N_8433,N_8874);
and U9364 (N_9364,N_7891,N_7913);
or U9365 (N_9365,N_8061,N_7844);
xor U9366 (N_9366,N_8027,N_8707);
xnor U9367 (N_9367,N_7593,N_7589);
nand U9368 (N_9368,N_8382,N_8907);
and U9369 (N_9369,N_8252,N_8973);
nor U9370 (N_9370,N_8917,N_8269);
xnor U9371 (N_9371,N_8546,N_8420);
or U9372 (N_9372,N_7649,N_7625);
and U9373 (N_9373,N_8818,N_8823);
and U9374 (N_9374,N_8810,N_8193);
and U9375 (N_9375,N_7823,N_8582);
or U9376 (N_9376,N_8136,N_8075);
or U9377 (N_9377,N_7978,N_7571);
and U9378 (N_9378,N_7590,N_8509);
or U9379 (N_9379,N_8886,N_8480);
nand U9380 (N_9380,N_8445,N_8121);
nand U9381 (N_9381,N_8909,N_8475);
or U9382 (N_9382,N_7988,N_8859);
xor U9383 (N_9383,N_7669,N_8345);
or U9384 (N_9384,N_8034,N_8309);
and U9385 (N_9385,N_8322,N_7604);
nand U9386 (N_9386,N_7728,N_8527);
or U9387 (N_9387,N_8491,N_8994);
xnor U9388 (N_9388,N_8961,N_8233);
xnor U9389 (N_9389,N_8205,N_8678);
nand U9390 (N_9390,N_8285,N_8111);
and U9391 (N_9391,N_7889,N_7852);
xor U9392 (N_9392,N_8209,N_8352);
nor U9393 (N_9393,N_8464,N_8782);
and U9394 (N_9394,N_8473,N_8949);
xnor U9395 (N_9395,N_7883,N_8414);
nand U9396 (N_9396,N_7667,N_8797);
or U9397 (N_9397,N_8776,N_8808);
or U9398 (N_9398,N_7893,N_8079);
nor U9399 (N_9399,N_8792,N_8759);
xor U9400 (N_9400,N_8705,N_8564);
and U9401 (N_9401,N_8853,N_7764);
xnor U9402 (N_9402,N_7816,N_7748);
and U9403 (N_9403,N_7734,N_8817);
or U9404 (N_9404,N_7581,N_8619);
xnor U9405 (N_9405,N_8421,N_8609);
xor U9406 (N_9406,N_8317,N_7872);
or U9407 (N_9407,N_8898,N_8124);
nor U9408 (N_9408,N_8777,N_8150);
nor U9409 (N_9409,N_8621,N_7794);
or U9410 (N_9410,N_7858,N_8628);
nor U9411 (N_9411,N_8673,N_8767);
and U9412 (N_9412,N_7780,N_8241);
nor U9413 (N_9413,N_7689,N_7847);
and U9414 (N_9414,N_8041,N_8740);
or U9415 (N_9415,N_8783,N_8077);
xor U9416 (N_9416,N_8515,N_7741);
and U9417 (N_9417,N_8761,N_8923);
and U9418 (N_9418,N_8669,N_8020);
nor U9419 (N_9419,N_7885,N_7642);
nand U9420 (N_9420,N_7611,N_8895);
nor U9421 (N_9421,N_7607,N_8236);
xor U9422 (N_9422,N_8088,N_7665);
and U9423 (N_9423,N_7986,N_8687);
xnor U9424 (N_9424,N_7771,N_7787);
nand U9425 (N_9425,N_7613,N_8095);
or U9426 (N_9426,N_7965,N_8367);
nand U9427 (N_9427,N_7837,N_7546);
nor U9428 (N_9428,N_8262,N_8341);
xnor U9429 (N_9429,N_8013,N_8735);
xor U9430 (N_9430,N_8381,N_8844);
nor U9431 (N_9431,N_7882,N_8319);
nand U9432 (N_9432,N_7551,N_8246);
xnor U9433 (N_9433,N_8570,N_8365);
or U9434 (N_9434,N_8074,N_8204);
nor U9435 (N_9435,N_8362,N_7830);
and U9436 (N_9436,N_8856,N_8329);
xor U9437 (N_9437,N_8523,N_8467);
xor U9438 (N_9438,N_8082,N_7747);
and U9439 (N_9439,N_7595,N_8432);
nand U9440 (N_9440,N_8734,N_8913);
nor U9441 (N_9441,N_7645,N_8833);
xor U9442 (N_9442,N_8830,N_8956);
nor U9443 (N_9443,N_7550,N_8539);
xor U9444 (N_9444,N_8044,N_8282);
and U9445 (N_9445,N_8085,N_7798);
nand U9446 (N_9446,N_7629,N_8416);
or U9447 (N_9447,N_8347,N_8868);
nor U9448 (N_9448,N_7776,N_8879);
or U9449 (N_9449,N_7682,N_7759);
and U9450 (N_9450,N_7632,N_7775);
and U9451 (N_9451,N_8526,N_8867);
or U9452 (N_9452,N_8809,N_8988);
nor U9453 (N_9453,N_7732,N_8584);
nand U9454 (N_9454,N_8049,N_7839);
nand U9455 (N_9455,N_7580,N_7970);
nand U9456 (N_9456,N_8211,N_7657);
or U9457 (N_9457,N_7952,N_8114);
or U9458 (N_9458,N_8813,N_7946);
xor U9459 (N_9459,N_8832,N_8901);
and U9460 (N_9460,N_8162,N_7690);
nand U9461 (N_9461,N_8977,N_7992);
and U9462 (N_9462,N_7987,N_7630);
and U9463 (N_9463,N_7917,N_8649);
nand U9464 (N_9464,N_8154,N_8402);
nor U9465 (N_9465,N_7812,N_8652);
nand U9466 (N_9466,N_8428,N_8850);
xor U9467 (N_9467,N_7809,N_8864);
and U9468 (N_9468,N_8585,N_8656);
or U9469 (N_9469,N_8762,N_7514);
xnor U9470 (N_9470,N_7622,N_8645);
nand U9471 (N_9471,N_8441,N_8632);
and U9472 (N_9472,N_8424,N_8412);
and U9473 (N_9473,N_7532,N_7892);
nor U9474 (N_9474,N_8875,N_8980);
or U9475 (N_9475,N_7537,N_8819);
xor U9476 (N_9476,N_7579,N_8270);
xor U9477 (N_9477,N_8986,N_8884);
or U9478 (N_9478,N_8990,N_8430);
or U9479 (N_9479,N_8386,N_8210);
or U9480 (N_9480,N_8451,N_7778);
or U9481 (N_9481,N_8541,N_8912);
nor U9482 (N_9482,N_8134,N_8361);
nand U9483 (N_9483,N_7648,N_7526);
or U9484 (N_9484,N_8229,N_7762);
nor U9485 (N_9485,N_8918,N_8046);
and U9486 (N_9486,N_8016,N_7887);
xnor U9487 (N_9487,N_8520,N_8482);
nand U9488 (N_9488,N_8168,N_7975);
or U9489 (N_9489,N_7561,N_8943);
nand U9490 (N_9490,N_7668,N_7729);
xnor U9491 (N_9491,N_7909,N_7943);
xnor U9492 (N_9492,N_8921,N_8067);
xnor U9493 (N_9493,N_7902,N_7691);
and U9494 (N_9494,N_8413,N_7808);
nor U9495 (N_9495,N_8751,N_8841);
nor U9496 (N_9496,N_7890,N_7587);
or U9497 (N_9497,N_7768,N_8093);
nand U9498 (N_9498,N_8896,N_8581);
xnor U9499 (N_9499,N_7674,N_8999);
xnor U9500 (N_9500,N_7846,N_7939);
nor U9501 (N_9501,N_8255,N_8487);
and U9502 (N_9502,N_7807,N_8457);
nor U9503 (N_9503,N_7621,N_8756);
or U9504 (N_9504,N_8979,N_8477);
or U9505 (N_9505,N_8806,N_7704);
xor U9506 (N_9506,N_8574,N_7749);
and U9507 (N_9507,N_8974,N_7633);
nand U9508 (N_9508,N_8290,N_8042);
nor U9509 (N_9509,N_8196,N_8186);
nor U9510 (N_9510,N_8390,N_7636);
xor U9511 (N_9511,N_8338,N_8281);
and U9512 (N_9512,N_8754,N_8718);
xnor U9513 (N_9513,N_7896,N_8100);
nor U9514 (N_9514,N_8221,N_8495);
nand U9515 (N_9515,N_8010,N_8484);
nor U9516 (N_9516,N_7945,N_7610);
and U9517 (N_9517,N_7628,N_8344);
xor U9518 (N_9518,N_8234,N_7624);
and U9519 (N_9519,N_7718,N_8244);
or U9520 (N_9520,N_8360,N_8620);
nand U9521 (N_9521,N_7634,N_8622);
nor U9522 (N_9522,N_8286,N_7864);
xor U9523 (N_9523,N_8450,N_8260);
and U9524 (N_9524,N_8039,N_8054);
and U9525 (N_9525,N_7612,N_8291);
and U9526 (N_9526,N_8191,N_8228);
nand U9527 (N_9527,N_7549,N_7618);
xor U9528 (N_9528,N_8438,N_8201);
or U9529 (N_9529,N_7525,N_8237);
nor U9530 (N_9530,N_8092,N_8660);
or U9531 (N_9531,N_8256,N_7976);
nor U9532 (N_9532,N_7944,N_7614);
and U9533 (N_9533,N_8587,N_8590);
or U9534 (N_9534,N_8960,N_8133);
or U9535 (N_9535,N_8947,N_8058);
and U9536 (N_9536,N_7949,N_8223);
xor U9537 (N_9537,N_8135,N_8353);
xnor U9538 (N_9538,N_8906,N_8637);
or U9539 (N_9539,N_8519,N_8401);
xnor U9540 (N_9540,N_8553,N_7538);
nand U9541 (N_9541,N_7767,N_7941);
xnor U9542 (N_9542,N_8192,N_7982);
xor U9543 (N_9543,N_7608,N_8889);
nor U9544 (N_9544,N_8604,N_7757);
nor U9545 (N_9545,N_8066,N_7931);
or U9546 (N_9546,N_8326,N_8106);
or U9547 (N_9547,N_8614,N_8356);
nand U9548 (N_9548,N_8313,N_8483);
or U9549 (N_9549,N_8785,N_8852);
nand U9550 (N_9550,N_8063,N_8068);
nor U9551 (N_9551,N_8249,N_8968);
xnor U9552 (N_9552,N_7903,N_7874);
nor U9553 (N_9553,N_8440,N_7583);
nor U9554 (N_9554,N_8514,N_8331);
nand U9555 (N_9555,N_7738,N_8983);
xor U9556 (N_9556,N_8727,N_8486);
and U9557 (N_9557,N_8843,N_8342);
nand U9558 (N_9558,N_8764,N_8643);
nor U9559 (N_9559,N_7950,N_8456);
xnor U9560 (N_9560,N_8096,N_8954);
or U9561 (N_9561,N_8355,N_8474);
nand U9562 (N_9562,N_8461,N_8130);
nor U9563 (N_9563,N_8800,N_8366);
nand U9564 (N_9564,N_7743,N_8686);
xor U9565 (N_9565,N_8710,N_8927);
nand U9566 (N_9566,N_7567,N_7921);
or U9567 (N_9567,N_8499,N_8948);
or U9568 (N_9568,N_8453,N_8437);
and U9569 (N_9569,N_8107,N_8908);
nand U9570 (N_9570,N_8963,N_7971);
or U9571 (N_9571,N_8752,N_8743);
nor U9572 (N_9572,N_7782,N_8031);
or U9573 (N_9573,N_8562,N_7671);
xnor U9574 (N_9574,N_8931,N_8932);
nand U9575 (N_9575,N_7730,N_7552);
xnor U9576 (N_9576,N_7517,N_7556);
or U9577 (N_9577,N_8518,N_8465);
nor U9578 (N_9578,N_8940,N_8374);
nor U9579 (N_9579,N_8708,N_8663);
or U9580 (N_9580,N_8691,N_7663);
nor U9581 (N_9581,N_8052,N_8030);
nor U9582 (N_9582,N_8845,N_8084);
or U9583 (N_9583,N_8167,N_8772);
and U9584 (N_9584,N_8310,N_8062);
xnor U9585 (N_9585,N_8097,N_8017);
or U9586 (N_9586,N_8161,N_8595);
or U9587 (N_9587,N_7997,N_7641);
nand U9588 (N_9588,N_8283,N_8554);
nand U9589 (N_9589,N_8714,N_8243);
xnor U9590 (N_9590,N_8893,N_8877);
and U9591 (N_9591,N_8611,N_7753);
xnor U9592 (N_9592,N_8325,N_8032);
nand U9593 (N_9593,N_8551,N_8801);
or U9594 (N_9594,N_8602,N_8368);
and U9595 (N_9595,N_7661,N_7989);
or U9596 (N_9596,N_7973,N_7817);
or U9597 (N_9597,N_8003,N_8552);
or U9598 (N_9598,N_8905,N_7535);
or U9599 (N_9599,N_8009,N_7631);
and U9600 (N_9600,N_8887,N_8038);
nor U9601 (N_9601,N_7800,N_8398);
and U9602 (N_9602,N_8387,N_8476);
or U9603 (N_9603,N_7940,N_8447);
xnor U9604 (N_9604,N_8993,N_8257);
xor U9605 (N_9605,N_8890,N_8635);
nand U9606 (N_9606,N_8654,N_7544);
xor U9607 (N_9607,N_7878,N_8659);
xnor U9608 (N_9608,N_8471,N_8391);
nand U9609 (N_9609,N_8254,N_7672);
nand U9610 (N_9610,N_7745,N_8569);
xor U9611 (N_9611,N_7831,N_8591);
and U9612 (N_9612,N_7922,N_7744);
xor U9613 (N_9613,N_7548,N_8425);
and U9614 (N_9614,N_8535,N_7659);
nand U9615 (N_9615,N_7717,N_8799);
and U9616 (N_9616,N_8333,N_7715);
nor U9617 (N_9617,N_8627,N_8567);
nor U9618 (N_9618,N_8442,N_7698);
xnor U9619 (N_9619,N_8942,N_8610);
and U9620 (N_9620,N_8488,N_7705);
and U9621 (N_9621,N_8218,N_8997);
nor U9622 (N_9622,N_7699,N_8506);
or U9623 (N_9623,N_7592,N_8589);
nor U9624 (N_9624,N_7996,N_7826);
and U9625 (N_9625,N_8468,N_8145);
xor U9626 (N_9626,N_7983,N_8730);
and U9627 (N_9627,N_8146,N_8849);
nand U9628 (N_9628,N_8748,N_7825);
xnor U9629 (N_9629,N_8586,N_7820);
nor U9630 (N_9630,N_8343,N_8975);
nor U9631 (N_9631,N_7700,N_8699);
nor U9632 (N_9632,N_7527,N_7796);
xnor U9633 (N_9633,N_7813,N_7503);
nor U9634 (N_9634,N_8915,N_7867);
nand U9635 (N_9635,N_8299,N_7534);
nor U9636 (N_9636,N_8090,N_8758);
or U9637 (N_9637,N_8278,N_8164);
or U9638 (N_9638,N_7792,N_8790);
nand U9639 (N_9639,N_8359,N_8839);
and U9640 (N_9640,N_8296,N_8958);
xor U9641 (N_9641,N_8534,N_8287);
nor U9642 (N_9642,N_7523,N_8505);
nand U9643 (N_9643,N_8055,N_7519);
xnor U9644 (N_9644,N_8190,N_7866);
nor U9645 (N_9645,N_7907,N_8363);
nor U9646 (N_9646,N_8126,N_8404);
and U9647 (N_9647,N_8176,N_8902);
or U9648 (N_9648,N_8592,N_7739);
and U9649 (N_9649,N_8478,N_8207);
nor U9650 (N_9650,N_8597,N_7509);
and U9651 (N_9651,N_8065,N_8057);
and U9652 (N_9652,N_7791,N_8184);
and U9653 (N_9653,N_8006,N_7871);
xnor U9654 (N_9654,N_8076,N_8472);
nand U9655 (N_9655,N_7760,N_7998);
nor U9656 (N_9656,N_8737,N_7911);
xor U9657 (N_9657,N_8492,N_8337);
or U9658 (N_9658,N_7797,N_7936);
and U9659 (N_9659,N_7620,N_8302);
xor U9660 (N_9660,N_7522,N_8606);
xnor U9661 (N_9661,N_8512,N_8144);
nand U9662 (N_9662,N_8089,N_8503);
xor U9663 (N_9663,N_8443,N_8242);
or U9664 (N_9664,N_8920,N_7806);
nand U9665 (N_9665,N_8976,N_8612);
and U9666 (N_9666,N_7876,N_8029);
and U9667 (N_9667,N_7862,N_8883);
xor U9668 (N_9668,N_8284,N_8991);
nand U9669 (N_9669,N_8683,N_8251);
nand U9670 (N_9670,N_7558,N_8596);
xor U9671 (N_9671,N_8501,N_8728);
nand U9672 (N_9672,N_8138,N_8263);
xor U9673 (N_9673,N_7785,N_7942);
or U9674 (N_9674,N_8939,N_7795);
nor U9675 (N_9675,N_8891,N_8700);
or U9676 (N_9676,N_8725,N_7848);
xor U9677 (N_9677,N_8305,N_8458);
xnor U9678 (N_9678,N_7869,N_8769);
xor U9679 (N_9679,N_8739,N_8933);
nand U9680 (N_9680,N_8314,N_7627);
xnor U9681 (N_9681,N_8661,N_8626);
nand U9682 (N_9682,N_8422,N_7746);
xnor U9683 (N_9683,N_7678,N_7956);
nor U9684 (N_9684,N_7686,N_8261);
nor U9685 (N_9685,N_7960,N_8846);
xor U9686 (N_9686,N_8816,N_8731);
nand U9687 (N_9687,N_7822,N_8732);
nor U9688 (N_9688,N_8851,N_7599);
nor U9689 (N_9689,N_7870,N_7947);
xor U9690 (N_9690,N_8094,N_8226);
nand U9691 (N_9691,N_8080,N_8208);
nor U9692 (N_9692,N_7516,N_7828);
and U9693 (N_9693,N_8738,N_8607);
or U9694 (N_9694,N_8615,N_8557);
and U9695 (N_9695,N_8151,N_8814);
nand U9696 (N_9696,N_8273,N_7616);
nand U9697 (N_9697,N_8787,N_8837);
nor U9698 (N_9698,N_7564,N_7531);
nand U9699 (N_9699,N_8142,N_7664);
xnor U9700 (N_9700,N_7506,N_7836);
or U9701 (N_9701,N_8634,N_7559);
nor U9702 (N_9702,N_7679,N_8435);
xor U9703 (N_9703,N_8944,N_8540);
or U9704 (N_9704,N_8563,N_7959);
or U9705 (N_9705,N_8008,N_8924);
and U9706 (N_9706,N_8937,N_8380);
nand U9707 (N_9707,N_8248,N_8692);
or U9708 (N_9708,N_7643,N_8744);
and U9709 (N_9709,N_8119,N_7824);
xnor U9710 (N_9710,N_8522,N_7774);
xnor U9711 (N_9711,N_7927,N_8304);
or U9712 (N_9712,N_8537,N_7533);
nor U9713 (N_9713,N_8561,N_8742);
nand U9714 (N_9714,N_7928,N_8035);
or U9715 (N_9715,N_7692,N_8618);
xnor U9716 (N_9716,N_8214,N_8071);
nor U9717 (N_9717,N_8315,N_8064);
and U9718 (N_9718,N_8773,N_8137);
and U9719 (N_9719,N_7626,N_8861);
nand U9720 (N_9720,N_8051,N_8995);
xor U9721 (N_9721,N_8827,N_8459);
nand U9722 (N_9722,N_7709,N_7979);
and U9723 (N_9723,N_8272,N_7646);
xnor U9724 (N_9724,N_8316,N_8230);
nor U9725 (N_9725,N_8481,N_8340);
nor U9726 (N_9726,N_8685,N_8560);
and U9727 (N_9727,N_7540,N_7512);
nor U9728 (N_9728,N_7582,N_8351);
or U9729 (N_9729,N_8295,N_8500);
xnor U9730 (N_9730,N_8513,N_7617);
xnor U9731 (N_9731,N_8418,N_8498);
and U9732 (N_9732,N_7637,N_7735);
and U9733 (N_9733,N_8358,N_7932);
and U9734 (N_9734,N_7510,N_8393);
xnor U9735 (N_9735,N_7710,N_7666);
nor U9736 (N_9736,N_8547,N_8383);
nor U9737 (N_9737,N_7967,N_8829);
nor U9738 (N_9738,N_8434,N_8987);
xnor U9739 (N_9739,N_8998,N_8568);
and U9740 (N_9740,N_8689,N_8395);
or U9741 (N_9741,N_8378,N_7507);
and U9742 (N_9742,N_8953,N_8294);
nand U9743 (N_9743,N_8593,N_8826);
or U9744 (N_9744,N_8914,N_7677);
nor U9745 (N_9745,N_8675,N_8306);
or U9746 (N_9746,N_7701,N_7781);
nand U9747 (N_9747,N_8377,N_8173);
xor U9748 (N_9748,N_8653,N_8770);
nand U9749 (N_9749,N_7601,N_8181);
nand U9750 (N_9750,N_7678,N_7973);
or U9751 (N_9751,N_7591,N_8627);
nor U9752 (N_9752,N_8053,N_7718);
nand U9753 (N_9753,N_7797,N_7905);
xnor U9754 (N_9754,N_8395,N_8318);
nand U9755 (N_9755,N_8635,N_8286);
nand U9756 (N_9756,N_8773,N_8513);
or U9757 (N_9757,N_8450,N_7712);
nor U9758 (N_9758,N_8673,N_7867);
nor U9759 (N_9759,N_7847,N_8741);
xnor U9760 (N_9760,N_7860,N_8263);
or U9761 (N_9761,N_7883,N_7995);
and U9762 (N_9762,N_8343,N_8780);
nor U9763 (N_9763,N_7977,N_7637);
or U9764 (N_9764,N_8884,N_8308);
nor U9765 (N_9765,N_8262,N_7878);
nor U9766 (N_9766,N_8056,N_7662);
nand U9767 (N_9767,N_7909,N_7502);
nand U9768 (N_9768,N_7853,N_7767);
nand U9769 (N_9769,N_8559,N_8253);
or U9770 (N_9770,N_8272,N_8486);
or U9771 (N_9771,N_7547,N_7939);
nand U9772 (N_9772,N_8466,N_8097);
and U9773 (N_9773,N_8083,N_7668);
nand U9774 (N_9774,N_7543,N_8601);
nand U9775 (N_9775,N_8775,N_8823);
or U9776 (N_9776,N_8309,N_8567);
nand U9777 (N_9777,N_8571,N_7723);
or U9778 (N_9778,N_7611,N_8962);
or U9779 (N_9779,N_7575,N_8801);
xnor U9780 (N_9780,N_8727,N_8315);
nand U9781 (N_9781,N_7836,N_8667);
nand U9782 (N_9782,N_7766,N_8081);
nor U9783 (N_9783,N_7659,N_7958);
nor U9784 (N_9784,N_7525,N_8376);
and U9785 (N_9785,N_7953,N_8230);
and U9786 (N_9786,N_8253,N_8255);
and U9787 (N_9787,N_8242,N_8440);
xor U9788 (N_9788,N_7823,N_8967);
or U9789 (N_9789,N_8437,N_8853);
or U9790 (N_9790,N_8572,N_8048);
nand U9791 (N_9791,N_8117,N_8361);
xor U9792 (N_9792,N_8914,N_7882);
xor U9793 (N_9793,N_8009,N_7879);
nand U9794 (N_9794,N_7788,N_8154);
or U9795 (N_9795,N_7653,N_8342);
or U9796 (N_9796,N_8929,N_7718);
or U9797 (N_9797,N_8448,N_7980);
xor U9798 (N_9798,N_7852,N_8107);
nand U9799 (N_9799,N_8188,N_7688);
nor U9800 (N_9800,N_7676,N_8728);
xnor U9801 (N_9801,N_7753,N_8208);
xor U9802 (N_9802,N_8674,N_8008);
nor U9803 (N_9803,N_7639,N_7565);
nand U9804 (N_9804,N_7935,N_7676);
and U9805 (N_9805,N_7894,N_8454);
nor U9806 (N_9806,N_8508,N_8781);
or U9807 (N_9807,N_8030,N_7738);
or U9808 (N_9808,N_8986,N_8724);
nor U9809 (N_9809,N_8906,N_8652);
or U9810 (N_9810,N_7916,N_8431);
and U9811 (N_9811,N_8865,N_8906);
or U9812 (N_9812,N_8562,N_8845);
or U9813 (N_9813,N_8782,N_7520);
nand U9814 (N_9814,N_8370,N_8181);
or U9815 (N_9815,N_8575,N_7800);
or U9816 (N_9816,N_8485,N_7902);
and U9817 (N_9817,N_8466,N_8288);
or U9818 (N_9818,N_7682,N_8919);
xor U9819 (N_9819,N_8273,N_7860);
nor U9820 (N_9820,N_8313,N_8449);
xnor U9821 (N_9821,N_8430,N_7727);
or U9822 (N_9822,N_7796,N_8606);
nand U9823 (N_9823,N_8800,N_7564);
or U9824 (N_9824,N_8274,N_8254);
and U9825 (N_9825,N_8009,N_7601);
and U9826 (N_9826,N_8913,N_8671);
nor U9827 (N_9827,N_8713,N_8777);
nand U9828 (N_9828,N_8904,N_7960);
and U9829 (N_9829,N_8349,N_8320);
nor U9830 (N_9830,N_7572,N_8207);
xnor U9831 (N_9831,N_8260,N_8116);
or U9832 (N_9832,N_8030,N_7693);
and U9833 (N_9833,N_7598,N_8046);
nand U9834 (N_9834,N_7605,N_8348);
nor U9835 (N_9835,N_8122,N_8403);
xor U9836 (N_9836,N_7538,N_7993);
or U9837 (N_9837,N_7954,N_7881);
or U9838 (N_9838,N_7899,N_7923);
nand U9839 (N_9839,N_7933,N_7999);
xor U9840 (N_9840,N_8640,N_8511);
or U9841 (N_9841,N_8218,N_8388);
nand U9842 (N_9842,N_7772,N_7533);
xor U9843 (N_9843,N_7752,N_8216);
and U9844 (N_9844,N_8337,N_8919);
and U9845 (N_9845,N_8372,N_8898);
or U9846 (N_9846,N_8313,N_7610);
nor U9847 (N_9847,N_8915,N_8334);
and U9848 (N_9848,N_7581,N_7838);
nand U9849 (N_9849,N_8905,N_8676);
or U9850 (N_9850,N_8746,N_7557);
or U9851 (N_9851,N_8408,N_7665);
xnor U9852 (N_9852,N_8352,N_8194);
or U9853 (N_9853,N_8919,N_7916);
and U9854 (N_9854,N_8022,N_8646);
nor U9855 (N_9855,N_8616,N_7505);
nand U9856 (N_9856,N_8860,N_8682);
nand U9857 (N_9857,N_8411,N_8637);
or U9858 (N_9858,N_8831,N_8555);
nor U9859 (N_9859,N_8789,N_8822);
nor U9860 (N_9860,N_7524,N_7833);
or U9861 (N_9861,N_8666,N_7831);
or U9862 (N_9862,N_8030,N_8109);
nor U9863 (N_9863,N_7838,N_8874);
or U9864 (N_9864,N_8110,N_8497);
nand U9865 (N_9865,N_8941,N_8995);
nor U9866 (N_9866,N_8289,N_8467);
nor U9867 (N_9867,N_7556,N_7914);
or U9868 (N_9868,N_8430,N_8528);
nor U9869 (N_9869,N_7517,N_8693);
nand U9870 (N_9870,N_8999,N_8312);
xor U9871 (N_9871,N_8891,N_8626);
and U9872 (N_9872,N_7507,N_7524);
and U9873 (N_9873,N_8923,N_8828);
xor U9874 (N_9874,N_8968,N_7906);
and U9875 (N_9875,N_7887,N_8705);
nor U9876 (N_9876,N_8784,N_8287);
and U9877 (N_9877,N_7526,N_8026);
nor U9878 (N_9878,N_8599,N_7825);
and U9879 (N_9879,N_7999,N_8646);
nand U9880 (N_9880,N_8082,N_8243);
nand U9881 (N_9881,N_8879,N_8582);
xor U9882 (N_9882,N_7692,N_8843);
or U9883 (N_9883,N_8131,N_7680);
and U9884 (N_9884,N_8410,N_7696);
nand U9885 (N_9885,N_7755,N_7570);
or U9886 (N_9886,N_7699,N_7913);
and U9887 (N_9887,N_8697,N_8307);
or U9888 (N_9888,N_7864,N_8775);
nand U9889 (N_9889,N_8848,N_8717);
nand U9890 (N_9890,N_8122,N_8845);
nor U9891 (N_9891,N_8534,N_8028);
xor U9892 (N_9892,N_8277,N_7842);
nor U9893 (N_9893,N_8829,N_8005);
and U9894 (N_9894,N_8150,N_8238);
nand U9895 (N_9895,N_8463,N_7696);
xnor U9896 (N_9896,N_8576,N_7500);
and U9897 (N_9897,N_8298,N_8147);
or U9898 (N_9898,N_8982,N_8189);
and U9899 (N_9899,N_8281,N_8019);
nor U9900 (N_9900,N_7762,N_7742);
nor U9901 (N_9901,N_7534,N_8243);
nor U9902 (N_9902,N_8785,N_7990);
or U9903 (N_9903,N_8445,N_8205);
or U9904 (N_9904,N_8797,N_8885);
or U9905 (N_9905,N_7932,N_7738);
and U9906 (N_9906,N_8425,N_8120);
xnor U9907 (N_9907,N_8983,N_7981);
nand U9908 (N_9908,N_7975,N_8857);
nor U9909 (N_9909,N_8136,N_8058);
nor U9910 (N_9910,N_7990,N_7814);
nor U9911 (N_9911,N_7647,N_8533);
xor U9912 (N_9912,N_8118,N_8346);
nor U9913 (N_9913,N_8289,N_8126);
nand U9914 (N_9914,N_8690,N_8371);
nand U9915 (N_9915,N_8227,N_8684);
xnor U9916 (N_9916,N_7997,N_7853);
xnor U9917 (N_9917,N_7808,N_8544);
nor U9918 (N_9918,N_7748,N_7519);
xnor U9919 (N_9919,N_7732,N_8914);
and U9920 (N_9920,N_8739,N_8730);
and U9921 (N_9921,N_8540,N_8547);
xor U9922 (N_9922,N_7688,N_8102);
nand U9923 (N_9923,N_8159,N_8767);
nand U9924 (N_9924,N_7751,N_8378);
nand U9925 (N_9925,N_8483,N_8969);
nor U9926 (N_9926,N_8120,N_8096);
or U9927 (N_9927,N_8229,N_8419);
and U9928 (N_9928,N_8888,N_8123);
or U9929 (N_9929,N_8798,N_7527);
or U9930 (N_9930,N_8020,N_8256);
xor U9931 (N_9931,N_8490,N_8244);
nor U9932 (N_9932,N_8365,N_8876);
nor U9933 (N_9933,N_8942,N_7681);
nor U9934 (N_9934,N_8858,N_8530);
nand U9935 (N_9935,N_8019,N_7519);
and U9936 (N_9936,N_8912,N_8038);
xor U9937 (N_9937,N_7771,N_8972);
nor U9938 (N_9938,N_8652,N_8045);
nand U9939 (N_9939,N_8476,N_8846);
and U9940 (N_9940,N_7763,N_7743);
nand U9941 (N_9941,N_7503,N_8059);
and U9942 (N_9942,N_7791,N_7661);
xnor U9943 (N_9943,N_8480,N_8809);
nor U9944 (N_9944,N_7974,N_8316);
nor U9945 (N_9945,N_8201,N_7944);
nand U9946 (N_9946,N_8925,N_8966);
nand U9947 (N_9947,N_7821,N_7779);
xor U9948 (N_9948,N_8382,N_8281);
or U9949 (N_9949,N_7654,N_8018);
xor U9950 (N_9950,N_7802,N_7907);
or U9951 (N_9951,N_8748,N_8511);
nor U9952 (N_9952,N_7907,N_8397);
and U9953 (N_9953,N_8517,N_8507);
nand U9954 (N_9954,N_8427,N_8054);
xnor U9955 (N_9955,N_7769,N_7801);
and U9956 (N_9956,N_8215,N_8258);
nor U9957 (N_9957,N_8080,N_8026);
nand U9958 (N_9958,N_8582,N_7777);
xnor U9959 (N_9959,N_8752,N_8454);
xor U9960 (N_9960,N_8700,N_8031);
or U9961 (N_9961,N_7677,N_8261);
and U9962 (N_9962,N_7805,N_8824);
and U9963 (N_9963,N_8711,N_8413);
nand U9964 (N_9964,N_8218,N_8342);
and U9965 (N_9965,N_8884,N_8879);
nand U9966 (N_9966,N_7891,N_8575);
and U9967 (N_9967,N_8193,N_8671);
xnor U9968 (N_9968,N_7747,N_7895);
and U9969 (N_9969,N_7508,N_7959);
xor U9970 (N_9970,N_7589,N_7955);
and U9971 (N_9971,N_8796,N_8394);
and U9972 (N_9972,N_8258,N_8893);
xnor U9973 (N_9973,N_7951,N_8466);
nand U9974 (N_9974,N_8889,N_8691);
nor U9975 (N_9975,N_8174,N_8478);
or U9976 (N_9976,N_8517,N_7671);
nor U9977 (N_9977,N_8406,N_8577);
nand U9978 (N_9978,N_8657,N_7848);
xor U9979 (N_9979,N_8227,N_8574);
and U9980 (N_9980,N_8565,N_8681);
and U9981 (N_9981,N_7883,N_7981);
nand U9982 (N_9982,N_7950,N_8200);
or U9983 (N_9983,N_7719,N_7553);
xor U9984 (N_9984,N_8269,N_7608);
xnor U9985 (N_9985,N_7783,N_7861);
nor U9986 (N_9986,N_8841,N_8772);
xor U9987 (N_9987,N_8776,N_8858);
nand U9988 (N_9988,N_7608,N_8023);
nor U9989 (N_9989,N_8367,N_7629);
nand U9990 (N_9990,N_8615,N_8581);
nor U9991 (N_9991,N_7574,N_7983);
xor U9992 (N_9992,N_8315,N_8780);
or U9993 (N_9993,N_7703,N_7999);
nand U9994 (N_9994,N_7929,N_7520);
xnor U9995 (N_9995,N_8923,N_7621);
xnor U9996 (N_9996,N_8404,N_7676);
nor U9997 (N_9997,N_8423,N_7640);
or U9998 (N_9998,N_8116,N_8312);
or U9999 (N_9999,N_8358,N_7714);
or U10000 (N_10000,N_8177,N_8058);
and U10001 (N_10001,N_7820,N_7970);
or U10002 (N_10002,N_7651,N_8864);
xnor U10003 (N_10003,N_7794,N_7923);
and U10004 (N_10004,N_8229,N_7929);
or U10005 (N_10005,N_8787,N_8139);
nand U10006 (N_10006,N_7802,N_8923);
and U10007 (N_10007,N_7842,N_8215);
and U10008 (N_10008,N_8890,N_8277);
or U10009 (N_10009,N_7673,N_8927);
and U10010 (N_10010,N_8637,N_7684);
nand U10011 (N_10011,N_8636,N_8684);
nor U10012 (N_10012,N_7570,N_8548);
nor U10013 (N_10013,N_7579,N_8873);
nor U10014 (N_10014,N_8435,N_8044);
xor U10015 (N_10015,N_8228,N_8162);
xnor U10016 (N_10016,N_7755,N_8411);
and U10017 (N_10017,N_8976,N_7620);
nor U10018 (N_10018,N_7876,N_7576);
or U10019 (N_10019,N_7725,N_8263);
nor U10020 (N_10020,N_8681,N_7968);
and U10021 (N_10021,N_8868,N_7895);
or U10022 (N_10022,N_8153,N_8325);
nor U10023 (N_10023,N_8555,N_7779);
or U10024 (N_10024,N_7738,N_8066);
and U10025 (N_10025,N_8444,N_7616);
nand U10026 (N_10026,N_8013,N_8258);
or U10027 (N_10027,N_7697,N_7702);
xnor U10028 (N_10028,N_8309,N_8087);
or U10029 (N_10029,N_8192,N_8905);
nor U10030 (N_10030,N_7594,N_8573);
or U10031 (N_10031,N_8252,N_8931);
nand U10032 (N_10032,N_8089,N_8259);
nand U10033 (N_10033,N_8400,N_8161);
nor U10034 (N_10034,N_8590,N_8206);
nand U10035 (N_10035,N_8509,N_8284);
or U10036 (N_10036,N_7538,N_8500);
and U10037 (N_10037,N_7999,N_8073);
nor U10038 (N_10038,N_8255,N_8532);
or U10039 (N_10039,N_8785,N_7641);
xnor U10040 (N_10040,N_8960,N_8772);
and U10041 (N_10041,N_8633,N_8196);
nor U10042 (N_10042,N_8047,N_8991);
nand U10043 (N_10043,N_8337,N_8921);
and U10044 (N_10044,N_7836,N_7585);
nor U10045 (N_10045,N_8702,N_7688);
nor U10046 (N_10046,N_7836,N_8542);
xnor U10047 (N_10047,N_8850,N_8033);
and U10048 (N_10048,N_8845,N_7767);
and U10049 (N_10049,N_8064,N_7913);
nand U10050 (N_10050,N_8339,N_8027);
nand U10051 (N_10051,N_8639,N_8853);
nand U10052 (N_10052,N_7875,N_7879);
nor U10053 (N_10053,N_8488,N_8168);
and U10054 (N_10054,N_8817,N_8159);
or U10055 (N_10055,N_8517,N_8927);
xor U10056 (N_10056,N_8235,N_8469);
or U10057 (N_10057,N_8778,N_7658);
xor U10058 (N_10058,N_7693,N_8572);
nor U10059 (N_10059,N_8479,N_8612);
or U10060 (N_10060,N_7691,N_8112);
nand U10061 (N_10061,N_8555,N_8808);
xnor U10062 (N_10062,N_8706,N_8003);
or U10063 (N_10063,N_8996,N_8465);
or U10064 (N_10064,N_8575,N_8312);
and U10065 (N_10065,N_7604,N_7550);
nor U10066 (N_10066,N_7745,N_8494);
and U10067 (N_10067,N_7970,N_8189);
and U10068 (N_10068,N_8980,N_8888);
nand U10069 (N_10069,N_8705,N_7922);
xor U10070 (N_10070,N_8973,N_8199);
nand U10071 (N_10071,N_8387,N_7749);
xor U10072 (N_10072,N_7513,N_8504);
xor U10073 (N_10073,N_8100,N_8987);
nor U10074 (N_10074,N_8614,N_8281);
nand U10075 (N_10075,N_8540,N_8299);
nor U10076 (N_10076,N_8692,N_8618);
xnor U10077 (N_10077,N_8292,N_8780);
and U10078 (N_10078,N_7687,N_8298);
or U10079 (N_10079,N_8611,N_8704);
or U10080 (N_10080,N_8819,N_7787);
nor U10081 (N_10081,N_8049,N_8447);
or U10082 (N_10082,N_8391,N_8276);
nor U10083 (N_10083,N_8375,N_7814);
and U10084 (N_10084,N_7630,N_8674);
nor U10085 (N_10085,N_8967,N_7892);
or U10086 (N_10086,N_7606,N_7862);
nor U10087 (N_10087,N_7756,N_8439);
nand U10088 (N_10088,N_8530,N_8020);
nor U10089 (N_10089,N_8377,N_7963);
and U10090 (N_10090,N_8407,N_8999);
nor U10091 (N_10091,N_8491,N_7970);
xor U10092 (N_10092,N_8484,N_8407);
nor U10093 (N_10093,N_7960,N_7639);
nor U10094 (N_10094,N_8231,N_7785);
xor U10095 (N_10095,N_8927,N_7967);
or U10096 (N_10096,N_7765,N_8901);
or U10097 (N_10097,N_8246,N_7941);
and U10098 (N_10098,N_8216,N_8582);
nor U10099 (N_10099,N_8886,N_8105);
and U10100 (N_10100,N_8705,N_8233);
and U10101 (N_10101,N_7792,N_7852);
xor U10102 (N_10102,N_8196,N_7714);
xor U10103 (N_10103,N_8970,N_8388);
nor U10104 (N_10104,N_7701,N_8794);
nor U10105 (N_10105,N_8119,N_8080);
and U10106 (N_10106,N_7794,N_7720);
xnor U10107 (N_10107,N_7952,N_8482);
xnor U10108 (N_10108,N_7843,N_7728);
nand U10109 (N_10109,N_8936,N_7859);
and U10110 (N_10110,N_7585,N_8365);
nor U10111 (N_10111,N_8678,N_7523);
xnor U10112 (N_10112,N_8719,N_7608);
nor U10113 (N_10113,N_7944,N_7939);
or U10114 (N_10114,N_8684,N_8863);
xor U10115 (N_10115,N_8648,N_8383);
or U10116 (N_10116,N_8004,N_8215);
or U10117 (N_10117,N_8677,N_7864);
xnor U10118 (N_10118,N_7694,N_7541);
xor U10119 (N_10119,N_8979,N_8097);
nand U10120 (N_10120,N_8027,N_7956);
or U10121 (N_10121,N_8861,N_8743);
nor U10122 (N_10122,N_8752,N_7919);
nor U10123 (N_10123,N_8890,N_8219);
nand U10124 (N_10124,N_8667,N_8746);
xnor U10125 (N_10125,N_7521,N_8429);
xor U10126 (N_10126,N_8353,N_8697);
nand U10127 (N_10127,N_8269,N_8419);
nor U10128 (N_10128,N_7934,N_8482);
or U10129 (N_10129,N_7527,N_7913);
nand U10130 (N_10130,N_8473,N_7910);
xor U10131 (N_10131,N_7525,N_7873);
or U10132 (N_10132,N_7600,N_7599);
xor U10133 (N_10133,N_8886,N_8239);
nor U10134 (N_10134,N_8695,N_7970);
or U10135 (N_10135,N_7617,N_8206);
nand U10136 (N_10136,N_8070,N_7898);
xor U10137 (N_10137,N_8686,N_7868);
xor U10138 (N_10138,N_7619,N_8789);
nor U10139 (N_10139,N_8423,N_8549);
xor U10140 (N_10140,N_8618,N_8569);
xor U10141 (N_10141,N_8665,N_8037);
or U10142 (N_10142,N_7601,N_8590);
nand U10143 (N_10143,N_8415,N_8512);
or U10144 (N_10144,N_8156,N_7869);
nor U10145 (N_10145,N_8633,N_8934);
nor U10146 (N_10146,N_7562,N_8373);
nor U10147 (N_10147,N_8943,N_8809);
or U10148 (N_10148,N_8059,N_7530);
nor U10149 (N_10149,N_8209,N_7625);
or U10150 (N_10150,N_7984,N_8840);
or U10151 (N_10151,N_7657,N_7824);
xor U10152 (N_10152,N_7955,N_7525);
nor U10153 (N_10153,N_7874,N_7576);
nand U10154 (N_10154,N_8137,N_8651);
or U10155 (N_10155,N_8535,N_7649);
or U10156 (N_10156,N_7605,N_8168);
and U10157 (N_10157,N_7508,N_7595);
nor U10158 (N_10158,N_7622,N_8606);
and U10159 (N_10159,N_8681,N_7691);
nor U10160 (N_10160,N_8925,N_8432);
xor U10161 (N_10161,N_8654,N_8414);
xnor U10162 (N_10162,N_8233,N_8607);
or U10163 (N_10163,N_7503,N_8384);
or U10164 (N_10164,N_8830,N_7897);
nor U10165 (N_10165,N_8700,N_8481);
nand U10166 (N_10166,N_8151,N_7957);
and U10167 (N_10167,N_8540,N_7622);
and U10168 (N_10168,N_8270,N_8499);
and U10169 (N_10169,N_8645,N_8430);
and U10170 (N_10170,N_7586,N_7657);
nor U10171 (N_10171,N_7883,N_8085);
xor U10172 (N_10172,N_8754,N_8890);
and U10173 (N_10173,N_8033,N_8350);
nand U10174 (N_10174,N_8795,N_8082);
or U10175 (N_10175,N_8002,N_8085);
nor U10176 (N_10176,N_8928,N_7612);
or U10177 (N_10177,N_7634,N_7707);
or U10178 (N_10178,N_8387,N_7770);
nor U10179 (N_10179,N_7733,N_8654);
or U10180 (N_10180,N_8253,N_8307);
xnor U10181 (N_10181,N_8987,N_8931);
and U10182 (N_10182,N_8705,N_8403);
nand U10183 (N_10183,N_8881,N_8800);
nand U10184 (N_10184,N_8816,N_8971);
and U10185 (N_10185,N_7766,N_7843);
nor U10186 (N_10186,N_7796,N_7755);
or U10187 (N_10187,N_7953,N_8609);
xor U10188 (N_10188,N_8775,N_8528);
nand U10189 (N_10189,N_8059,N_8748);
and U10190 (N_10190,N_8552,N_8454);
xnor U10191 (N_10191,N_8048,N_8593);
nand U10192 (N_10192,N_8078,N_7904);
or U10193 (N_10193,N_8607,N_8919);
or U10194 (N_10194,N_8118,N_8782);
nand U10195 (N_10195,N_7959,N_8035);
nor U10196 (N_10196,N_7966,N_7558);
nand U10197 (N_10197,N_8237,N_8854);
nand U10198 (N_10198,N_8637,N_8152);
nor U10199 (N_10199,N_8567,N_8644);
or U10200 (N_10200,N_8283,N_8110);
or U10201 (N_10201,N_8959,N_8873);
or U10202 (N_10202,N_8001,N_8488);
xnor U10203 (N_10203,N_7569,N_8657);
nor U10204 (N_10204,N_7924,N_8852);
nand U10205 (N_10205,N_8425,N_8539);
nand U10206 (N_10206,N_8229,N_7687);
and U10207 (N_10207,N_8300,N_8069);
nand U10208 (N_10208,N_8407,N_8986);
or U10209 (N_10209,N_7891,N_7994);
nand U10210 (N_10210,N_8939,N_7962);
nand U10211 (N_10211,N_7905,N_8142);
or U10212 (N_10212,N_8610,N_8928);
or U10213 (N_10213,N_7979,N_8865);
nor U10214 (N_10214,N_8621,N_8087);
xor U10215 (N_10215,N_8012,N_7656);
and U10216 (N_10216,N_8524,N_8377);
xnor U10217 (N_10217,N_8667,N_7864);
nor U10218 (N_10218,N_8770,N_7894);
and U10219 (N_10219,N_7635,N_8929);
and U10220 (N_10220,N_8112,N_8132);
and U10221 (N_10221,N_8457,N_7581);
and U10222 (N_10222,N_8426,N_7552);
nand U10223 (N_10223,N_8793,N_7977);
and U10224 (N_10224,N_8754,N_7770);
and U10225 (N_10225,N_7822,N_8251);
or U10226 (N_10226,N_8290,N_7988);
or U10227 (N_10227,N_8483,N_8801);
xor U10228 (N_10228,N_8758,N_8348);
xor U10229 (N_10229,N_8232,N_8841);
nor U10230 (N_10230,N_8252,N_8211);
xor U10231 (N_10231,N_8191,N_8696);
or U10232 (N_10232,N_8273,N_7938);
xor U10233 (N_10233,N_7895,N_7598);
nand U10234 (N_10234,N_7904,N_7954);
or U10235 (N_10235,N_7986,N_8933);
nor U10236 (N_10236,N_8454,N_7996);
nand U10237 (N_10237,N_8234,N_8072);
and U10238 (N_10238,N_8453,N_8132);
xnor U10239 (N_10239,N_8582,N_7762);
xor U10240 (N_10240,N_7661,N_8111);
or U10241 (N_10241,N_8354,N_8738);
and U10242 (N_10242,N_7537,N_7927);
nand U10243 (N_10243,N_8835,N_7873);
nor U10244 (N_10244,N_7554,N_8551);
and U10245 (N_10245,N_8013,N_8885);
and U10246 (N_10246,N_8247,N_8201);
or U10247 (N_10247,N_7513,N_7673);
nand U10248 (N_10248,N_7547,N_7720);
xnor U10249 (N_10249,N_7908,N_8987);
nand U10250 (N_10250,N_7996,N_8240);
nor U10251 (N_10251,N_8364,N_7648);
nor U10252 (N_10252,N_8729,N_7833);
and U10253 (N_10253,N_8334,N_8353);
nor U10254 (N_10254,N_8261,N_8791);
xnor U10255 (N_10255,N_7939,N_8829);
or U10256 (N_10256,N_7695,N_7665);
xor U10257 (N_10257,N_8134,N_8826);
or U10258 (N_10258,N_8503,N_8839);
and U10259 (N_10259,N_8614,N_8629);
or U10260 (N_10260,N_7623,N_8604);
nand U10261 (N_10261,N_8455,N_8208);
nand U10262 (N_10262,N_8797,N_7572);
and U10263 (N_10263,N_8971,N_8151);
xor U10264 (N_10264,N_7801,N_7638);
nand U10265 (N_10265,N_8761,N_8336);
xnor U10266 (N_10266,N_7683,N_8997);
or U10267 (N_10267,N_8084,N_8069);
xnor U10268 (N_10268,N_7873,N_8945);
xor U10269 (N_10269,N_8553,N_8938);
and U10270 (N_10270,N_7825,N_7916);
or U10271 (N_10271,N_8673,N_8208);
or U10272 (N_10272,N_7822,N_8852);
and U10273 (N_10273,N_7601,N_8082);
and U10274 (N_10274,N_7941,N_7971);
and U10275 (N_10275,N_8436,N_8724);
or U10276 (N_10276,N_8733,N_8224);
and U10277 (N_10277,N_8225,N_8217);
or U10278 (N_10278,N_7772,N_8631);
xor U10279 (N_10279,N_8421,N_8999);
and U10280 (N_10280,N_8404,N_8807);
nor U10281 (N_10281,N_7622,N_8605);
or U10282 (N_10282,N_7552,N_7860);
nor U10283 (N_10283,N_7908,N_7524);
nor U10284 (N_10284,N_7610,N_7788);
nand U10285 (N_10285,N_7896,N_8819);
and U10286 (N_10286,N_7671,N_8990);
nand U10287 (N_10287,N_7917,N_8890);
xnor U10288 (N_10288,N_8383,N_8754);
or U10289 (N_10289,N_8833,N_8955);
nor U10290 (N_10290,N_8933,N_7653);
nand U10291 (N_10291,N_8693,N_8091);
nor U10292 (N_10292,N_8466,N_8678);
xnor U10293 (N_10293,N_7515,N_8557);
xnor U10294 (N_10294,N_8859,N_8225);
or U10295 (N_10295,N_7591,N_8386);
or U10296 (N_10296,N_8480,N_8192);
xnor U10297 (N_10297,N_8661,N_8405);
nor U10298 (N_10298,N_7546,N_8749);
nor U10299 (N_10299,N_8810,N_8405);
nor U10300 (N_10300,N_7575,N_7948);
nor U10301 (N_10301,N_7715,N_7674);
or U10302 (N_10302,N_8561,N_8418);
xnor U10303 (N_10303,N_7532,N_8356);
or U10304 (N_10304,N_7546,N_8111);
nand U10305 (N_10305,N_8473,N_8476);
and U10306 (N_10306,N_8329,N_8440);
or U10307 (N_10307,N_8111,N_8892);
nand U10308 (N_10308,N_8963,N_8101);
and U10309 (N_10309,N_8390,N_8513);
xnor U10310 (N_10310,N_7634,N_8563);
or U10311 (N_10311,N_7657,N_7621);
nor U10312 (N_10312,N_7802,N_8741);
nand U10313 (N_10313,N_7533,N_8045);
xor U10314 (N_10314,N_8091,N_8737);
or U10315 (N_10315,N_8413,N_8488);
nor U10316 (N_10316,N_7626,N_8978);
nand U10317 (N_10317,N_8658,N_8279);
nor U10318 (N_10318,N_8916,N_8284);
or U10319 (N_10319,N_7667,N_8083);
nand U10320 (N_10320,N_7987,N_7691);
nor U10321 (N_10321,N_8888,N_7764);
and U10322 (N_10322,N_8987,N_7643);
or U10323 (N_10323,N_7537,N_7943);
or U10324 (N_10324,N_8766,N_8674);
and U10325 (N_10325,N_7656,N_8443);
nand U10326 (N_10326,N_8297,N_8161);
or U10327 (N_10327,N_8121,N_8663);
xnor U10328 (N_10328,N_8622,N_8383);
xor U10329 (N_10329,N_7632,N_7619);
xor U10330 (N_10330,N_7847,N_7556);
or U10331 (N_10331,N_8465,N_8067);
or U10332 (N_10332,N_7630,N_8019);
nand U10333 (N_10333,N_8968,N_8138);
nand U10334 (N_10334,N_8076,N_8116);
xnor U10335 (N_10335,N_7879,N_8860);
xnor U10336 (N_10336,N_8480,N_8635);
or U10337 (N_10337,N_8129,N_8573);
xnor U10338 (N_10338,N_8613,N_8170);
nand U10339 (N_10339,N_7514,N_8692);
and U10340 (N_10340,N_7787,N_8323);
xnor U10341 (N_10341,N_8103,N_8335);
or U10342 (N_10342,N_7678,N_8232);
and U10343 (N_10343,N_7640,N_7541);
nor U10344 (N_10344,N_8289,N_8986);
and U10345 (N_10345,N_7874,N_8029);
xor U10346 (N_10346,N_8978,N_7973);
xnor U10347 (N_10347,N_7849,N_8556);
or U10348 (N_10348,N_8434,N_8324);
and U10349 (N_10349,N_8449,N_7575);
xor U10350 (N_10350,N_8849,N_8108);
or U10351 (N_10351,N_7868,N_7709);
xor U10352 (N_10352,N_7666,N_8404);
nand U10353 (N_10353,N_8607,N_7710);
nor U10354 (N_10354,N_7594,N_8910);
or U10355 (N_10355,N_8115,N_7892);
nor U10356 (N_10356,N_8893,N_8419);
xnor U10357 (N_10357,N_8445,N_8929);
nand U10358 (N_10358,N_7803,N_8543);
nand U10359 (N_10359,N_7780,N_8979);
xor U10360 (N_10360,N_7641,N_8076);
and U10361 (N_10361,N_8639,N_8466);
nor U10362 (N_10362,N_8004,N_8354);
and U10363 (N_10363,N_8666,N_8254);
xor U10364 (N_10364,N_7507,N_8301);
nand U10365 (N_10365,N_7555,N_8590);
nor U10366 (N_10366,N_7826,N_8037);
nand U10367 (N_10367,N_8106,N_8472);
and U10368 (N_10368,N_8083,N_8779);
xor U10369 (N_10369,N_7736,N_7650);
nand U10370 (N_10370,N_8417,N_8501);
and U10371 (N_10371,N_8722,N_8813);
nand U10372 (N_10372,N_8408,N_8124);
and U10373 (N_10373,N_8504,N_8903);
nand U10374 (N_10374,N_8161,N_8917);
xor U10375 (N_10375,N_7648,N_7690);
or U10376 (N_10376,N_8804,N_7993);
or U10377 (N_10377,N_8374,N_7643);
and U10378 (N_10378,N_8991,N_7842);
nor U10379 (N_10379,N_7867,N_8979);
and U10380 (N_10380,N_7647,N_8467);
xnor U10381 (N_10381,N_8949,N_7889);
nand U10382 (N_10382,N_8661,N_8176);
xor U10383 (N_10383,N_7928,N_8554);
and U10384 (N_10384,N_7918,N_8011);
or U10385 (N_10385,N_7661,N_7776);
or U10386 (N_10386,N_8187,N_8201);
nand U10387 (N_10387,N_8881,N_8743);
and U10388 (N_10388,N_8209,N_7612);
nor U10389 (N_10389,N_7623,N_8943);
or U10390 (N_10390,N_8601,N_8754);
nand U10391 (N_10391,N_7951,N_8812);
xor U10392 (N_10392,N_7675,N_7963);
or U10393 (N_10393,N_8094,N_8460);
xor U10394 (N_10394,N_8539,N_8249);
nor U10395 (N_10395,N_7504,N_8622);
nor U10396 (N_10396,N_8534,N_8087);
or U10397 (N_10397,N_7526,N_8498);
nor U10398 (N_10398,N_8739,N_7559);
nor U10399 (N_10399,N_8953,N_7912);
or U10400 (N_10400,N_8275,N_8377);
or U10401 (N_10401,N_7913,N_7928);
and U10402 (N_10402,N_8003,N_8372);
xnor U10403 (N_10403,N_7823,N_7767);
nand U10404 (N_10404,N_7724,N_8493);
or U10405 (N_10405,N_8701,N_7739);
or U10406 (N_10406,N_8542,N_8316);
nand U10407 (N_10407,N_8056,N_7862);
xnor U10408 (N_10408,N_8642,N_8558);
or U10409 (N_10409,N_7734,N_7736);
xnor U10410 (N_10410,N_8298,N_7741);
nand U10411 (N_10411,N_7712,N_8756);
or U10412 (N_10412,N_8129,N_8471);
xor U10413 (N_10413,N_8746,N_8026);
nand U10414 (N_10414,N_8565,N_8573);
nor U10415 (N_10415,N_8271,N_8734);
xnor U10416 (N_10416,N_8222,N_8001);
or U10417 (N_10417,N_7852,N_7747);
or U10418 (N_10418,N_8582,N_8329);
nand U10419 (N_10419,N_7660,N_8971);
nor U10420 (N_10420,N_8819,N_7817);
xor U10421 (N_10421,N_8586,N_8247);
or U10422 (N_10422,N_8886,N_8257);
nand U10423 (N_10423,N_7811,N_8608);
and U10424 (N_10424,N_8978,N_8288);
or U10425 (N_10425,N_8814,N_8857);
nor U10426 (N_10426,N_8406,N_8086);
and U10427 (N_10427,N_8468,N_8172);
nand U10428 (N_10428,N_7662,N_7936);
xor U10429 (N_10429,N_8151,N_7636);
nand U10430 (N_10430,N_8057,N_7842);
or U10431 (N_10431,N_8363,N_7929);
xor U10432 (N_10432,N_8443,N_8452);
nor U10433 (N_10433,N_8355,N_8508);
or U10434 (N_10434,N_7994,N_8267);
or U10435 (N_10435,N_7613,N_8136);
and U10436 (N_10436,N_8064,N_8430);
nand U10437 (N_10437,N_8040,N_8760);
and U10438 (N_10438,N_8888,N_7773);
or U10439 (N_10439,N_8527,N_8024);
nand U10440 (N_10440,N_7917,N_7745);
xnor U10441 (N_10441,N_8312,N_8016);
and U10442 (N_10442,N_8175,N_8002);
or U10443 (N_10443,N_7856,N_8780);
xor U10444 (N_10444,N_7630,N_8435);
nor U10445 (N_10445,N_7579,N_8585);
xor U10446 (N_10446,N_7847,N_8926);
xnor U10447 (N_10447,N_8365,N_8805);
nor U10448 (N_10448,N_8452,N_8973);
nand U10449 (N_10449,N_8047,N_8653);
nand U10450 (N_10450,N_8566,N_7919);
and U10451 (N_10451,N_7522,N_8091);
or U10452 (N_10452,N_8335,N_8949);
or U10453 (N_10453,N_8938,N_8308);
xnor U10454 (N_10454,N_8112,N_7824);
nand U10455 (N_10455,N_8896,N_8839);
xor U10456 (N_10456,N_8661,N_8958);
and U10457 (N_10457,N_8636,N_7736);
and U10458 (N_10458,N_8776,N_7802);
nor U10459 (N_10459,N_8644,N_8828);
nor U10460 (N_10460,N_8028,N_8977);
or U10461 (N_10461,N_8663,N_8335);
xor U10462 (N_10462,N_8600,N_8452);
nor U10463 (N_10463,N_8853,N_8892);
and U10464 (N_10464,N_7808,N_7671);
nand U10465 (N_10465,N_8774,N_8692);
nand U10466 (N_10466,N_8944,N_8100);
or U10467 (N_10467,N_8902,N_7715);
or U10468 (N_10468,N_8261,N_8374);
or U10469 (N_10469,N_8026,N_8535);
nor U10470 (N_10470,N_8271,N_7614);
xnor U10471 (N_10471,N_7602,N_8611);
or U10472 (N_10472,N_7750,N_8154);
nand U10473 (N_10473,N_8741,N_8465);
and U10474 (N_10474,N_7691,N_8547);
nor U10475 (N_10475,N_8641,N_7967);
nor U10476 (N_10476,N_7865,N_8354);
nand U10477 (N_10477,N_8065,N_8255);
nand U10478 (N_10478,N_7598,N_7896);
nand U10479 (N_10479,N_8908,N_8756);
nand U10480 (N_10480,N_8155,N_8994);
nand U10481 (N_10481,N_8000,N_7512);
or U10482 (N_10482,N_8948,N_7953);
or U10483 (N_10483,N_8624,N_8182);
nor U10484 (N_10484,N_7726,N_8121);
and U10485 (N_10485,N_7571,N_8168);
and U10486 (N_10486,N_8842,N_8315);
or U10487 (N_10487,N_8637,N_8394);
nand U10488 (N_10488,N_8374,N_8945);
or U10489 (N_10489,N_8020,N_8813);
nor U10490 (N_10490,N_7582,N_8829);
xor U10491 (N_10491,N_8381,N_8905);
nor U10492 (N_10492,N_8729,N_7858);
or U10493 (N_10493,N_8630,N_8473);
xor U10494 (N_10494,N_8994,N_8406);
xor U10495 (N_10495,N_7980,N_8401);
nor U10496 (N_10496,N_8222,N_8676);
and U10497 (N_10497,N_7996,N_8174);
or U10498 (N_10498,N_8800,N_8192);
nor U10499 (N_10499,N_8181,N_8420);
and U10500 (N_10500,N_10049,N_9878);
nor U10501 (N_10501,N_9501,N_10156);
xor U10502 (N_10502,N_10448,N_9844);
or U10503 (N_10503,N_9447,N_9240);
and U10504 (N_10504,N_9037,N_10416);
and U10505 (N_10505,N_9009,N_10423);
and U10506 (N_10506,N_10101,N_9884);
nor U10507 (N_10507,N_9904,N_9534);
xnor U10508 (N_10508,N_10118,N_9306);
and U10509 (N_10509,N_10075,N_9492);
and U10510 (N_10510,N_9111,N_9473);
xor U10511 (N_10511,N_10497,N_9033);
nand U10512 (N_10512,N_9368,N_9161);
and U10513 (N_10513,N_9462,N_9711);
nand U10514 (N_10514,N_10474,N_9935);
or U10515 (N_10515,N_10026,N_9087);
and U10516 (N_10516,N_9493,N_9923);
xnor U10517 (N_10517,N_9200,N_9331);
xor U10518 (N_10518,N_10360,N_9661);
nand U10519 (N_10519,N_9470,N_10337);
or U10520 (N_10520,N_10232,N_9336);
xor U10521 (N_10521,N_10123,N_9750);
xor U10522 (N_10522,N_9848,N_9619);
nor U10523 (N_10523,N_9321,N_10334);
nor U10524 (N_10524,N_9029,N_9951);
nor U10525 (N_10525,N_10256,N_9660);
nand U10526 (N_10526,N_10287,N_10457);
or U10527 (N_10527,N_9245,N_9141);
nand U10528 (N_10528,N_9633,N_9516);
nor U10529 (N_10529,N_9254,N_9498);
nand U10530 (N_10530,N_10456,N_9965);
nand U10531 (N_10531,N_9605,N_10144);
xor U10532 (N_10532,N_9128,N_9603);
xor U10533 (N_10533,N_9337,N_9713);
xor U10534 (N_10534,N_9068,N_10235);
xnor U10535 (N_10535,N_10175,N_10453);
nand U10536 (N_10536,N_9913,N_9433);
nor U10537 (N_10537,N_9806,N_10335);
or U10538 (N_10538,N_9397,N_9294);
nand U10539 (N_10539,N_10293,N_9872);
nand U10540 (N_10540,N_9512,N_9461);
nand U10541 (N_10541,N_9517,N_9518);
nor U10542 (N_10542,N_10259,N_9443);
xor U10543 (N_10543,N_9456,N_9197);
nand U10544 (N_10544,N_9561,N_9837);
and U10545 (N_10545,N_9757,N_10260);
nand U10546 (N_10546,N_9258,N_10310);
xnor U10547 (N_10547,N_10447,N_10097);
nand U10548 (N_10548,N_10429,N_9706);
nor U10549 (N_10549,N_9278,N_10017);
nor U10550 (N_10550,N_9914,N_10289);
xor U10551 (N_10551,N_9975,N_9910);
nand U10552 (N_10552,N_9808,N_9487);
or U10553 (N_10553,N_10234,N_10299);
or U10554 (N_10554,N_9595,N_9001);
and U10555 (N_10555,N_9234,N_9202);
or U10556 (N_10556,N_10014,N_9530);
xor U10557 (N_10557,N_9880,N_9210);
or U10558 (N_10558,N_9007,N_10090);
nand U10559 (N_10559,N_10094,N_9869);
or U10560 (N_10560,N_9101,N_10476);
or U10561 (N_10561,N_9268,N_9537);
and U10562 (N_10562,N_9286,N_10152);
nor U10563 (N_10563,N_9908,N_9296);
nor U10564 (N_10564,N_9526,N_9751);
xnor U10565 (N_10565,N_10327,N_9421);
nand U10566 (N_10566,N_10063,N_10137);
nand U10567 (N_10567,N_9395,N_10394);
nand U10568 (N_10568,N_10043,N_9220);
xor U10569 (N_10569,N_10353,N_10300);
and U10570 (N_10570,N_9986,N_9227);
nand U10571 (N_10571,N_10011,N_9825);
xnor U10572 (N_10572,N_9628,N_9264);
nand U10573 (N_10573,N_9369,N_10395);
nand U10574 (N_10574,N_10076,N_9155);
and U10575 (N_10575,N_9702,N_9484);
xnor U10576 (N_10576,N_9957,N_9683);
or U10577 (N_10577,N_9795,N_10182);
or U10578 (N_10578,N_9644,N_10323);
or U10579 (N_10579,N_10404,N_10085);
and U10580 (N_10580,N_9119,N_9066);
xor U10581 (N_10581,N_9123,N_10460);
or U10582 (N_10582,N_9873,N_9819);
nand U10583 (N_10583,N_9906,N_9250);
nand U10584 (N_10584,N_9246,N_9838);
nor U10585 (N_10585,N_10467,N_9899);
and U10586 (N_10586,N_10045,N_9973);
nand U10587 (N_10587,N_9055,N_9002);
and U10588 (N_10588,N_9723,N_9771);
nor U10589 (N_10589,N_9737,N_9247);
nor U10590 (N_10590,N_10158,N_9292);
nand U10591 (N_10591,N_10082,N_9849);
xor U10592 (N_10592,N_10095,N_9366);
and U10593 (N_10593,N_9347,N_10122);
xnor U10594 (N_10594,N_10445,N_10272);
nor U10595 (N_10595,N_9499,N_9449);
nand U10596 (N_10596,N_9866,N_9617);
and U10597 (N_10597,N_10393,N_9677);
xnor U10598 (N_10598,N_9569,N_9021);
xnor U10599 (N_10599,N_9828,N_9401);
xor U10600 (N_10600,N_9544,N_10473);
xnor U10601 (N_10601,N_9558,N_9062);
xnor U10602 (N_10602,N_9172,N_9414);
or U10603 (N_10603,N_9792,N_10107);
or U10604 (N_10604,N_10325,N_10146);
xnor U10605 (N_10605,N_9483,N_9094);
nand U10606 (N_10606,N_9931,N_9375);
xor U10607 (N_10607,N_9998,N_9404);
or U10608 (N_10608,N_10336,N_10074);
xor U10609 (N_10609,N_9417,N_9394);
and U10610 (N_10610,N_10003,N_9237);
and U10611 (N_10611,N_9497,N_9471);
nand U10612 (N_10612,N_10406,N_9173);
xor U10613 (N_10613,N_9511,N_9427);
xor U10614 (N_10614,N_9047,N_9129);
nor U10615 (N_10615,N_9672,N_9898);
and U10616 (N_10616,N_9276,N_10153);
nor U10617 (N_10617,N_9658,N_10266);
xor U10618 (N_10618,N_9359,N_10060);
nand U10619 (N_10619,N_9142,N_9620);
or U10620 (N_10620,N_10389,N_10160);
xor U10621 (N_10621,N_9460,N_10405);
xnor U10622 (N_10622,N_9508,N_9540);
or U10623 (N_10623,N_9810,N_10058);
and U10624 (N_10624,N_10297,N_10145);
and U10625 (N_10625,N_9715,N_9136);
xnor U10626 (N_10626,N_9550,N_9139);
xor U10627 (N_10627,N_9106,N_9695);
and U10628 (N_10628,N_9663,N_10113);
nand U10629 (N_10629,N_9831,N_9432);
and U10630 (N_10630,N_10485,N_10154);
and U10631 (N_10631,N_9145,N_10044);
and U10632 (N_10632,N_9153,N_9410);
nor U10633 (N_10633,N_9862,N_9624);
nor U10634 (N_10634,N_9575,N_9478);
xnor U10635 (N_10635,N_9870,N_9938);
nand U10636 (N_10636,N_10440,N_9284);
nor U10637 (N_10637,N_9398,N_9285);
nor U10638 (N_10638,N_10414,N_9939);
xnor U10639 (N_10639,N_10126,N_9360);
and U10640 (N_10640,N_10274,N_9669);
xor U10641 (N_10641,N_10252,N_9385);
nand U10642 (N_10642,N_9097,N_9084);
and U10643 (N_10643,N_9670,N_9339);
nand U10644 (N_10644,N_10087,N_9112);
xnor U10645 (N_10645,N_10285,N_9753);
nand U10646 (N_10646,N_9598,N_9697);
xor U10647 (N_10647,N_9547,N_9266);
and U10648 (N_10648,N_9754,N_10243);
or U10649 (N_10649,N_9437,N_9448);
nor U10650 (N_10650,N_9177,N_9010);
and U10651 (N_10651,N_10140,N_9761);
or U10652 (N_10652,N_9978,N_10210);
and U10653 (N_10653,N_9747,N_9921);
nand U10654 (N_10654,N_9272,N_10065);
xor U10655 (N_10655,N_10373,N_9459);
nor U10656 (N_10656,N_9131,N_9157);
and U10657 (N_10657,N_10073,N_10403);
xnor U10658 (N_10658,N_9515,N_9358);
and U10659 (N_10659,N_9728,N_9779);
xor U10660 (N_10660,N_9566,N_9950);
nand U10661 (N_10661,N_9730,N_9820);
xor U10662 (N_10662,N_9580,N_10315);
and U10663 (N_10663,N_10007,N_10171);
or U10664 (N_10664,N_9122,N_10281);
nand U10665 (N_10665,N_10498,N_10039);
and U10666 (N_10666,N_9583,N_9428);
and U10667 (N_10667,N_9228,N_10368);
and U10668 (N_10668,N_10472,N_9996);
and U10669 (N_10669,N_9548,N_9942);
nand U10670 (N_10670,N_9796,N_9961);
nand U10671 (N_10671,N_9564,N_9623);
nand U10672 (N_10672,N_10419,N_9915);
or U10673 (N_10673,N_9574,N_10383);
nor U10674 (N_10674,N_9774,N_9287);
xnor U10675 (N_10675,N_10169,N_10173);
nand U10676 (N_10676,N_10214,N_10271);
and U10677 (N_10677,N_9496,N_9152);
nand U10678 (N_10678,N_9940,N_9926);
or U10679 (N_10679,N_10374,N_9570);
xnor U10680 (N_10680,N_10277,N_9643);
xnor U10681 (N_10681,N_9219,N_10278);
or U10682 (N_10682,N_10016,N_9242);
or U10683 (N_10683,N_10211,N_10181);
nor U10684 (N_10684,N_10046,N_10320);
nor U10685 (N_10685,N_9997,N_9768);
or U10686 (N_10686,N_9992,N_9507);
xnor U10687 (N_10687,N_10066,N_9045);
xor U10688 (N_10688,N_10301,N_9291);
nand U10689 (N_10689,N_9041,N_9626);
and U10690 (N_10690,N_9650,N_9146);
and U10691 (N_10691,N_10262,N_9221);
nand U10692 (N_10692,N_9143,N_9503);
and U10693 (N_10693,N_9834,N_10163);
nand U10694 (N_10694,N_9922,N_9308);
and U10695 (N_10695,N_9412,N_9743);
nor U10696 (N_10696,N_10290,N_9042);
xor U10697 (N_10697,N_10324,N_9093);
nand U10698 (N_10698,N_10298,N_9257);
xnor U10699 (N_10699,N_9364,N_10209);
nand U10700 (N_10700,N_9634,N_9968);
and U10701 (N_10701,N_9019,N_9393);
xor U10702 (N_10702,N_9351,N_9678);
nand U10703 (N_10703,N_9400,N_9107);
and U10704 (N_10704,N_9759,N_9164);
nor U10705 (N_10705,N_9431,N_9630);
nand U10706 (N_10706,N_10319,N_9165);
xor U10707 (N_10707,N_10139,N_9439);
and U10708 (N_10708,N_9453,N_9857);
nand U10709 (N_10709,N_10254,N_9399);
and U10710 (N_10710,N_10286,N_10420);
nand U10711 (N_10711,N_9912,N_9746);
xor U10712 (N_10712,N_9475,N_9151);
nand U10713 (N_10713,N_10151,N_9271);
nor U10714 (N_10714,N_9382,N_9253);
nand U10715 (N_10715,N_9874,N_10331);
nand U10716 (N_10716,N_9451,N_9436);
and U10717 (N_10717,N_9786,N_9841);
xor U10718 (N_10718,N_9827,N_10443);
nand U10719 (N_10719,N_10031,N_9091);
nor U10720 (N_10720,N_10080,N_9749);
and U10721 (N_10721,N_10109,N_9689);
xnor U10722 (N_10722,N_9947,N_10461);
or U10723 (N_10723,N_9147,N_9944);
nand U10724 (N_10724,N_9435,N_9373);
nand U10725 (N_10725,N_9556,N_10358);
nor U10726 (N_10726,N_9936,N_9799);
and U10727 (N_10727,N_9323,N_10023);
and U10728 (N_10728,N_10413,N_9290);
nor U10729 (N_10729,N_9303,N_10083);
nand U10730 (N_10730,N_9764,N_9752);
nand U10731 (N_10731,N_9787,N_9557);
xnor U10732 (N_10732,N_10350,N_9946);
xor U10733 (N_10733,N_10032,N_9724);
nand U10734 (N_10734,N_9704,N_9543);
nand U10735 (N_10735,N_9571,N_9735);
nand U10736 (N_10736,N_9046,N_9967);
nand U10737 (N_10737,N_9896,N_10417);
nand U10738 (N_10738,N_10370,N_9847);
or U10739 (N_10739,N_10048,N_10427);
and U10740 (N_10740,N_9283,N_9627);
xnor U10741 (N_10741,N_9408,N_10333);
xor U10742 (N_10742,N_9158,N_9314);
xnor U10743 (N_10743,N_10422,N_9481);
nor U10744 (N_10744,N_9260,N_9017);
nor U10745 (N_10745,N_9117,N_9618);
nor U10746 (N_10746,N_10435,N_9334);
nand U10747 (N_10747,N_9244,N_9765);
xnor U10748 (N_10748,N_9241,N_10084);
nand U10749 (N_10749,N_9892,N_10008);
or U10750 (N_10750,N_9629,N_9554);
and U10751 (N_10751,N_9674,N_9034);
and U10752 (N_10752,N_9440,N_9324);
or U10753 (N_10753,N_9977,N_10069);
nor U10754 (N_10754,N_9013,N_9175);
nor U10755 (N_10755,N_9805,N_10465);
and U10756 (N_10756,N_10332,N_10451);
or U10757 (N_10757,N_9927,N_9252);
xnor U10758 (N_10758,N_9355,N_9745);
nand U10759 (N_10759,N_10437,N_9816);
or U10760 (N_10760,N_9519,N_9609);
and U10761 (N_10761,N_9450,N_9654);
or U10762 (N_10762,N_9154,N_9160);
nor U10763 (N_10763,N_10072,N_9316);
xor U10764 (N_10764,N_9269,N_10407);
nor U10765 (N_10765,N_10219,N_9933);
nand U10766 (N_10766,N_9708,N_9277);
or U10767 (N_10767,N_9879,N_9971);
and U10768 (N_10768,N_10105,N_10352);
and U10769 (N_10769,N_10067,N_10459);
xor U10770 (N_10770,N_10167,N_9187);
or U10771 (N_10771,N_10041,N_10313);
and U10772 (N_10772,N_9807,N_9549);
xor U10773 (N_10773,N_9059,N_10086);
or U10774 (N_10774,N_10196,N_10365);
nand U10775 (N_10775,N_10280,N_9419);
and U10776 (N_10776,N_9299,N_9030);
nor U10777 (N_10777,N_10304,N_9125);
and U10778 (N_10778,N_9482,N_9109);
or U10779 (N_10779,N_9022,N_10050);
xnor U10780 (N_10780,N_9144,N_9201);
or U10781 (N_10781,N_9063,N_10180);
or U10782 (N_10782,N_10070,N_9486);
xor U10783 (N_10783,N_10489,N_9166);
xor U10784 (N_10784,N_9867,N_9632);
nand U10785 (N_10785,N_10390,N_10054);
xnor U10786 (N_10786,N_10379,N_9803);
xor U10787 (N_10787,N_9226,N_9053);
nor U10788 (N_10788,N_9189,N_10159);
xor U10789 (N_10789,N_9858,N_10378);
or U10790 (N_10790,N_10446,N_10077);
nand U10791 (N_10791,N_10364,N_9929);
or U10792 (N_10792,N_9409,N_10255);
xnor U10793 (N_10793,N_10356,N_9963);
xnor U10794 (N_10794,N_9918,N_9315);
xor U10795 (N_10795,N_10469,N_9687);
xor U10796 (N_10796,N_10068,N_9261);
xnor U10797 (N_10797,N_10279,N_9829);
xnor U10798 (N_10798,N_9008,N_10096);
and U10799 (N_10799,N_10000,N_9777);
nand U10800 (N_10800,N_9020,N_9667);
and U10801 (N_10801,N_9374,N_9104);
and U10802 (N_10802,N_9073,N_10071);
and U10803 (N_10803,N_10265,N_10454);
or U10804 (N_10804,N_10291,N_9529);
xnor U10805 (N_10805,N_9920,N_9089);
nand U10806 (N_10806,N_9864,N_10369);
and U10807 (N_10807,N_9686,N_10436);
xor U10808 (N_10808,N_9523,N_10288);
and U10809 (N_10809,N_9585,N_9536);
nand U10810 (N_10810,N_9811,N_9108);
xor U10811 (N_10811,N_10317,N_9974);
and U10812 (N_10812,N_9607,N_9930);
xor U10813 (N_10813,N_10006,N_9891);
and U10814 (N_10814,N_10246,N_10191);
nand U10815 (N_10815,N_10098,N_10468);
and U10816 (N_10816,N_9466,N_9680);
xnor U10817 (N_10817,N_9895,N_9733);
xor U10818 (N_10818,N_9190,N_9835);
nor U10819 (N_10819,N_10387,N_10021);
xor U10820 (N_10820,N_9179,N_10455);
or U10821 (N_10821,N_9541,N_9991);
xnor U10822 (N_10822,N_10491,N_10239);
xnor U10823 (N_10823,N_9812,N_9772);
xor U10824 (N_10824,N_9140,N_9781);
or U10825 (N_10825,N_9953,N_10248);
xor U10826 (N_10826,N_10092,N_9070);
xor U10827 (N_10827,N_10292,N_10062);
or U10828 (N_10828,N_10268,N_9510);
nor U10829 (N_10829,N_9163,N_9325);
nor U10830 (N_10830,N_9591,N_9911);
nand U10831 (N_10831,N_9600,N_10177);
or U10832 (N_10832,N_9881,N_10036);
nand U10833 (N_10833,N_9340,N_9238);
xor U10834 (N_10834,N_9608,N_9668);
nor U10835 (N_10835,N_9304,N_10375);
xor U10836 (N_10836,N_10424,N_9211);
xnor U10837 (N_10837,N_9185,N_10164);
nand U10838 (N_10838,N_9442,N_10061);
nor U10839 (N_10839,N_10012,N_10481);
or U10840 (N_10840,N_10380,N_9701);
and U10841 (N_10841,N_9300,N_9684);
and U10842 (N_10842,N_10345,N_9673);
xor U10843 (N_10843,N_9124,N_9649);
and U10844 (N_10844,N_9945,N_9763);
or U10845 (N_10845,N_9937,N_9958);
xnor U10846 (N_10846,N_9365,N_9602);
nand U10847 (N_10847,N_9876,N_9824);
or U10848 (N_10848,N_9567,N_10376);
and U10849 (N_10849,N_10463,N_9345);
or U10850 (N_10850,N_9424,N_10149);
nand U10851 (N_10851,N_9578,N_9514);
nand U10852 (N_10852,N_10240,N_9601);
and U10853 (N_10853,N_9954,N_10306);
and U10854 (N_10854,N_10157,N_10480);
and U10855 (N_10855,N_10125,N_10218);
nand U10856 (N_10856,N_10212,N_9215);
nor U10857 (N_10857,N_9061,N_9096);
nor U10858 (N_10858,N_10458,N_9114);
nand U10859 (N_10859,N_10314,N_10493);
or U10860 (N_10860,N_10206,N_9208);
or U10861 (N_10861,N_10487,N_10193);
or U10862 (N_10862,N_9330,N_9472);
nand U10863 (N_10863,N_9760,N_10386);
nor U10864 (N_10864,N_9413,N_9741);
and U10865 (N_10865,N_9983,N_9818);
or U10866 (N_10866,N_10190,N_9302);
or U10867 (N_10867,N_9348,N_9714);
nand U10868 (N_10868,N_10222,N_10110);
nor U10869 (N_10869,N_9092,N_10432);
xnor U10870 (N_10870,N_9229,N_10203);
or U10871 (N_10871,N_9357,N_9889);
or U10872 (N_10872,N_9665,N_10185);
xnor U10873 (N_10873,N_10261,N_9979);
nor U10874 (N_10874,N_10247,N_10385);
xor U10875 (N_10875,N_10479,N_9137);
or U10876 (N_10876,N_9298,N_9318);
and U10877 (N_10877,N_9727,N_10019);
or U10878 (N_10878,N_9069,N_9295);
and U10879 (N_10879,N_10205,N_9794);
nand U10880 (N_10880,N_9095,N_9744);
nand U10881 (N_10881,N_9637,N_9722);
xnor U10882 (N_10882,N_10047,N_9297);
or U10883 (N_10883,N_10344,N_9110);
nand U10884 (N_10884,N_10148,N_9716);
xnor U10885 (N_10885,N_9115,N_9489);
or U10886 (N_10886,N_9804,N_9490);
xor U10887 (N_10887,N_9793,N_9116);
or U10888 (N_10888,N_9026,N_9885);
nand U10889 (N_10889,N_10001,N_9445);
xor U10890 (N_10890,N_10131,N_9662);
xor U10891 (N_10891,N_9363,N_9981);
or U10892 (N_10892,N_10347,N_9988);
xor U10893 (N_10893,N_10362,N_9987);
and U10894 (N_10894,N_10172,N_10035);
or U10895 (N_10895,N_10184,N_10127);
nand U10896 (N_10896,N_10270,N_9192);
nor U10897 (N_10897,N_10229,N_9532);
xor U10898 (N_10898,N_9495,N_9589);
nor U10899 (N_10899,N_9132,N_9383);
nand U10900 (N_10900,N_10161,N_10197);
nand U10901 (N_10901,N_9748,N_10138);
nand U10902 (N_10902,N_9188,N_9802);
and U10903 (N_10903,N_9265,N_9313);
and U10904 (N_10904,N_9797,N_9823);
or U10905 (N_10905,N_9040,N_10377);
or U10906 (N_10906,N_9681,N_9186);
nor U10907 (N_10907,N_9718,N_10466);
and U10908 (N_10908,N_10482,N_9354);
nor U10909 (N_10909,N_9434,N_10117);
nor U10910 (N_10910,N_10115,N_10116);
and U10911 (N_10911,N_10400,N_9048);
nor U10912 (N_10912,N_9388,N_10147);
and U10913 (N_10913,N_10484,N_10475);
xnor U10914 (N_10914,N_10307,N_10015);
nor U10915 (N_10915,N_9280,N_9994);
nand U10916 (N_10916,N_9615,N_9352);
nand U10917 (N_10917,N_10119,N_10078);
nand U10918 (N_10918,N_9016,N_9893);
nor U10919 (N_10919,N_10490,N_9328);
or U10920 (N_10920,N_9477,N_9319);
or U10921 (N_10921,N_9180,N_10309);
nand U10922 (N_10922,N_10284,N_9648);
nand U10923 (N_10923,N_10189,N_10183);
and U10924 (N_10924,N_10464,N_9830);
xor U10925 (N_10925,N_10442,N_10056);
or U10926 (N_10926,N_10020,N_9076);
nand U10927 (N_10927,N_9756,N_9080);
nor U10928 (N_10928,N_10305,N_10471);
and U10929 (N_10929,N_10207,N_9102);
nand U10930 (N_10930,N_9350,N_9389);
or U10931 (N_10931,N_9120,N_9218);
nand U10932 (N_10932,N_9039,N_9288);
xnor U10933 (N_10933,N_10186,N_9584);
nor U10934 (N_10934,N_9506,N_10418);
or U10935 (N_10935,N_9446,N_9568);
or U10936 (N_10936,N_9642,N_10081);
xor U10937 (N_10937,N_9692,N_9441);
or U10938 (N_10938,N_9025,N_9865);
or U10939 (N_10939,N_9613,N_9035);
or U10940 (N_10940,N_9731,N_10361);
xor U10941 (N_10941,N_9652,N_9457);
and U10942 (N_10942,N_9058,N_9989);
or U10943 (N_10943,N_10228,N_10408);
nand U10944 (N_10944,N_9943,N_9758);
xnor U10945 (N_10945,N_10253,N_10022);
xor U10946 (N_10946,N_9023,N_9966);
nand U10947 (N_10947,N_9871,N_9176);
xnor U10948 (N_10948,N_9616,N_10302);
or U10949 (N_10949,N_10318,N_10341);
nor U10950 (N_10950,N_10141,N_9635);
nor U10951 (N_10951,N_10402,N_9332);
nand U10952 (N_10952,N_9338,N_9289);
xnor U10953 (N_10953,N_10059,N_10415);
nand U10954 (N_10954,N_10295,N_9156);
and U10955 (N_10955,N_9552,N_9485);
and U10956 (N_10956,N_9479,N_9209);
nand U10957 (N_10957,N_9995,N_9740);
nand U10958 (N_10958,N_9962,N_9028);
and U10959 (N_10959,N_9535,N_9312);
or U10960 (N_10960,N_10339,N_9604);
nand U10961 (N_10961,N_10296,N_9705);
nor U10962 (N_10962,N_9367,N_9928);
nand U10963 (N_10963,N_9463,N_9729);
or U10964 (N_10964,N_9814,N_10208);
nor U10965 (N_10965,N_9640,N_9868);
xnor U10966 (N_10966,N_10216,N_10162);
and U10967 (N_10967,N_10276,N_9082);
nor U10968 (N_10968,N_9262,N_9387);
xnor U10969 (N_10969,N_10321,N_9588);
and U10970 (N_10970,N_9577,N_9327);
nand U10971 (N_10971,N_9888,N_9167);
nor U10972 (N_10972,N_10294,N_9842);
nand U10973 (N_10973,N_9239,N_9719);
and U10974 (N_10974,N_10150,N_9625);
and U10975 (N_10975,N_9148,N_9183);
xor U10976 (N_10976,N_9390,N_9085);
xor U10977 (N_10977,N_10037,N_9392);
or U10978 (N_10978,N_9322,N_9491);
or U10979 (N_10979,N_10030,N_10124);
and U10980 (N_10980,N_9181,N_9833);
nor U10981 (N_10981,N_9659,N_10338);
xnor U10982 (N_10982,N_10194,N_10174);
nor U10983 (N_10983,N_10308,N_10439);
or U10984 (N_10984,N_9476,N_10411);
xor U10985 (N_10985,N_10462,N_9249);
nor U10986 (N_10986,N_9370,N_10004);
xnor U10987 (N_10987,N_10340,N_9948);
xor U10988 (N_10988,N_10371,N_9438);
xnor U10989 (N_10989,N_10382,N_10367);
nor U10990 (N_10990,N_9356,N_9972);
nand U10991 (N_10991,N_10057,N_10053);
and U10992 (N_10992,N_10396,N_9088);
or U10993 (N_10993,N_9853,N_9311);
or U10994 (N_10994,N_9320,N_10135);
xnor U10995 (N_10995,N_9243,N_10267);
or U10996 (N_10996,N_9118,N_9418);
xnor U10997 (N_10997,N_9317,N_10034);
or U10998 (N_10998,N_10275,N_9361);
or U10999 (N_10999,N_9054,N_10195);
nor U11000 (N_11000,N_9699,N_9664);
and U11001 (N_11001,N_10486,N_9329);
or U11002 (N_11002,N_9279,N_9402);
xor U11003 (N_11003,N_9700,N_9480);
nor U11004 (N_11004,N_9901,N_9984);
xnor U11005 (N_11005,N_10391,N_10244);
or U11006 (N_11006,N_9646,N_9206);
nand U11007 (N_11007,N_10496,N_9416);
or U11008 (N_11008,N_9454,N_9582);
nand U11009 (N_11009,N_9196,N_9647);
or U11010 (N_11010,N_9698,N_9083);
or U11011 (N_11011,N_9344,N_9964);
nor U11012 (N_11012,N_10238,N_9909);
xor U11013 (N_11013,N_10355,N_9883);
or U11014 (N_11014,N_9839,N_9105);
or U11015 (N_11015,N_9378,N_10166);
xnor U11016 (N_11016,N_9732,N_9133);
nand U11017 (N_11017,N_9845,N_10249);
nand U11018 (N_11018,N_9012,N_9126);
nor U11019 (N_11019,N_10093,N_10002);
and U11020 (N_11020,N_10410,N_9075);
nand U11021 (N_11021,N_10282,N_10328);
and U11022 (N_11022,N_10111,N_10351);
or U11023 (N_11023,N_9043,N_10384);
xor U11024 (N_11024,N_10263,N_9504);
or U11025 (N_11025,N_9565,N_9099);
and U11026 (N_11026,N_9381,N_9500);
and U11027 (N_11027,N_10354,N_10311);
xnor U11028 (N_11028,N_9710,N_9403);
and U11029 (N_11029,N_10114,N_10392);
or U11030 (N_11030,N_10326,N_10102);
nor U11031 (N_11031,N_10492,N_9924);
or U11032 (N_11032,N_9693,N_9212);
nand U11033 (N_11033,N_9800,N_9738);
or U11034 (N_11034,N_10100,N_9612);
and U11035 (N_11035,N_9721,N_9422);
and U11036 (N_11036,N_9293,N_9970);
and U11037 (N_11037,N_10033,N_9840);
and U11038 (N_11038,N_10129,N_10176);
xor U11039 (N_11039,N_9855,N_9191);
or U11040 (N_11040,N_9464,N_9343);
or U11041 (N_11041,N_9657,N_9690);
or U11042 (N_11042,N_10434,N_9709);
xnor U11043 (N_11043,N_9011,N_9533);
xor U11044 (N_11044,N_9606,N_10024);
and U11045 (N_11045,N_10303,N_10038);
nor U11046 (N_11046,N_10227,N_10200);
nor U11047 (N_11047,N_9694,N_9003);
nand U11048 (N_11048,N_9232,N_9138);
nor U11049 (N_11049,N_9259,N_9856);
and U11050 (N_11050,N_9121,N_10204);
or U11051 (N_11051,N_10433,N_9169);
nor U11052 (N_11052,N_9377,N_10231);
nand U11053 (N_11053,N_9307,N_9980);
nand U11054 (N_11054,N_9894,N_9900);
or U11055 (N_11055,N_9579,N_9391);
and U11056 (N_11056,N_9521,N_9813);
or U11057 (N_11057,N_9420,N_9000);
nor U11058 (N_11058,N_9224,N_10201);
xnor U11059 (N_11059,N_9406,N_10132);
or U11060 (N_11060,N_9776,N_9005);
or U11061 (N_11061,N_9767,N_9773);
xor U11062 (N_11062,N_9952,N_10236);
xor U11063 (N_11063,N_9815,N_9203);
and U11064 (N_11064,N_9217,N_10258);
xor U11065 (N_11065,N_9386,N_9572);
nor U11066 (N_11066,N_10088,N_9233);
xor U11067 (N_11067,N_9782,N_9353);
xor U11068 (N_11068,N_9852,N_10343);
nand U11069 (N_11069,N_9326,N_10198);
nand U11070 (N_11070,N_9999,N_9941);
and U11071 (N_11071,N_9522,N_9982);
and U11072 (N_11072,N_9090,N_9528);
nor U11073 (N_11073,N_10438,N_9969);
and U11074 (N_11074,N_9594,N_9411);
and U11075 (N_11075,N_9726,N_9494);
and U11076 (N_11076,N_9551,N_10494);
and U11077 (N_11077,N_9778,N_9596);
nand U11078 (N_11078,N_10128,N_9100);
or U11079 (N_11079,N_10136,N_10426);
nand U11080 (N_11080,N_9655,N_9052);
nand U11081 (N_11081,N_10441,N_9426);
nand U11082 (N_11082,N_9273,N_9843);
nand U11083 (N_11083,N_9060,N_9465);
nor U11084 (N_11084,N_9875,N_9919);
nand U11085 (N_11085,N_9956,N_9809);
and U11086 (N_11086,N_9127,N_9538);
nand U11087 (N_11087,N_10091,N_10168);
and U11088 (N_11088,N_9072,N_9555);
nand U11089 (N_11089,N_10220,N_10027);
and U11090 (N_11090,N_9251,N_9882);
nor U11091 (N_11091,N_9525,N_9791);
xor U11092 (N_11092,N_10316,N_9455);
or U11093 (N_11093,N_9335,N_9452);
or U11094 (N_11094,N_10366,N_10192);
xnor U11095 (N_11095,N_9645,N_9785);
xnor U11096 (N_11096,N_10170,N_9006);
nor U11097 (N_11097,N_9917,N_10241);
xor U11098 (N_11098,N_9934,N_9194);
or U11099 (N_11099,N_9639,N_9204);
nand U11100 (N_11100,N_10452,N_9907);
nand U11101 (N_11101,N_9079,N_9651);
nand U11102 (N_11102,N_10421,N_9641);
and U11103 (N_11103,N_9309,N_10143);
nor U11104 (N_11104,N_10251,N_9581);
xor U11105 (N_11105,N_9783,N_10042);
nor U11106 (N_11106,N_9790,N_9916);
nand U11107 (N_11107,N_10202,N_9734);
nand U11108 (N_11108,N_9762,N_10401);
nand U11109 (N_11109,N_9717,N_9405);
and U11110 (N_11110,N_10425,N_9990);
nand U11111 (N_11111,N_9223,N_10359);
nand U11112 (N_11112,N_10230,N_9231);
nand U11113 (N_11113,N_9149,N_10449);
nand U11114 (N_11114,N_9230,N_9134);
or U11115 (N_11115,N_10273,N_9178);
or U11116 (N_11116,N_10470,N_9836);
nand U11117 (N_11117,N_10217,N_10499);
nor U11118 (N_11118,N_9766,N_10226);
or U11119 (N_11119,N_10106,N_9064);
nor U11120 (N_11120,N_9396,N_10346);
nor U11121 (N_11121,N_10018,N_9769);
nand U11122 (N_11122,N_9362,N_9597);
or U11123 (N_11123,N_10283,N_9505);
xor U11124 (N_11124,N_10223,N_10478);
nor U11125 (N_11125,N_10103,N_9184);
nand U11126 (N_11126,N_9576,N_9859);
or U11127 (N_11127,N_9542,N_9044);
nor U11128 (N_11128,N_9425,N_9056);
nor U11129 (N_11129,N_10187,N_9955);
or U11130 (N_11130,N_9676,N_9621);
or U11131 (N_11131,N_10250,N_9174);
xnor U11132 (N_11132,N_10025,N_9074);
or U11133 (N_11133,N_9346,N_9553);
nor U11134 (N_11134,N_9671,N_10409);
or U11135 (N_11135,N_10224,N_10178);
nand U11136 (N_11136,N_9103,N_10079);
or U11137 (N_11137,N_10450,N_9707);
nor U11138 (N_11138,N_9255,N_10155);
nand U11139 (N_11139,N_9205,N_9004);
nor U11140 (N_11140,N_9712,N_10040);
or U11141 (N_11141,N_10188,N_10215);
xnor U11142 (N_11142,N_9788,N_10388);
xnor U11143 (N_11143,N_9902,N_10329);
nor U11144 (N_11144,N_9301,N_9216);
nand U11145 (N_11145,N_10055,N_10483);
or U11146 (N_11146,N_9474,N_9488);
xnor U11147 (N_11147,N_9696,N_9275);
xor U11148 (N_11148,N_9036,N_9691);
xor U11149 (N_11149,N_10312,N_9851);
and U11150 (N_11150,N_9038,N_10225);
xor U11151 (N_11151,N_9599,N_10120);
nor U11152 (N_11152,N_10104,N_9586);
and U11153 (N_11153,N_9531,N_9592);
nand U11154 (N_11154,N_9078,N_9235);
or U11155 (N_11155,N_9817,N_9614);
or U11156 (N_11156,N_9371,N_9198);
and U11157 (N_11157,N_9631,N_9587);
and U11158 (N_11158,N_10430,N_9985);
and U11159 (N_11159,N_9267,N_9086);
and U11160 (N_11160,N_9057,N_9380);
nand U11161 (N_11161,N_9636,N_9832);
nor U11162 (N_11162,N_10179,N_9031);
xnor U11163 (N_11163,N_9458,N_10348);
and U11164 (N_11164,N_9376,N_9349);
xnor U11165 (N_11165,N_9468,N_10269);
nor U11166 (N_11166,N_10381,N_9770);
nor U11167 (N_11167,N_10213,N_9736);
nand U11168 (N_11168,N_9801,N_9342);
nand U11169 (N_11169,N_9653,N_10005);
nand U11170 (N_11170,N_10349,N_9520);
nor U11171 (N_11171,N_9854,N_9850);
nand U11172 (N_11172,N_10398,N_9236);
nand U11173 (N_11173,N_9077,N_9049);
or U11174 (N_11174,N_10089,N_10357);
nand U11175 (N_11175,N_9524,N_10029);
and U11176 (N_11176,N_9281,N_9282);
xnor U11177 (N_11177,N_9135,N_9014);
nor U11178 (N_11178,N_9423,N_10495);
xnor U11179 (N_11179,N_10330,N_9222);
xnor U11180 (N_11180,N_10428,N_9469);
xor U11181 (N_11181,N_9467,N_10064);
xor U11182 (N_11182,N_9993,N_9846);
xor U11183 (N_11183,N_9780,N_9826);
or U11184 (N_11184,N_9513,N_9949);
xnor U11185 (N_11185,N_9113,N_9213);
and U11186 (N_11186,N_9860,N_9755);
xnor U11187 (N_11187,N_9071,N_10245);
and U11188 (N_11188,N_9798,N_10412);
xnor U11189 (N_11189,N_9720,N_9685);
nor U11190 (N_11190,N_10477,N_9263);
or U11191 (N_11191,N_9573,N_9861);
and U11192 (N_11192,N_9195,N_9675);
and U11193 (N_11193,N_9150,N_9877);
nor U11194 (N_11194,N_9546,N_10397);
or U11195 (N_11195,N_10051,N_9274);
or U11196 (N_11196,N_10028,N_9539);
nor U11197 (N_11197,N_10444,N_10130);
or U11198 (N_11198,N_10142,N_9333);
nor U11199 (N_11199,N_9903,N_9018);
nand U11200 (N_11200,N_9430,N_9682);
and U11201 (N_11201,N_9725,N_10342);
or U11202 (N_11202,N_10108,N_9890);
nand U11203 (N_11203,N_9784,N_9822);
nand U11204 (N_11204,N_9065,N_10322);
nand U11205 (N_11205,N_10133,N_9562);
or U11206 (N_11206,N_9341,N_9638);
nor U11207 (N_11207,N_9429,N_9656);
xor U11208 (N_11208,N_9863,N_9563);
xnor U11209 (N_11209,N_10112,N_9024);
xnor U11210 (N_11210,N_9162,N_9593);
and U11211 (N_11211,N_9821,N_9527);
and U11212 (N_11212,N_9739,N_9081);
or U11213 (N_11213,N_10013,N_9905);
and U11214 (N_11214,N_10052,N_9372);
nand U11215 (N_11215,N_9742,N_9193);
nor U11216 (N_11216,N_9015,N_9171);
xor U11217 (N_11217,N_9976,N_10010);
nor U11218 (N_11218,N_9182,N_9067);
nand U11219 (N_11219,N_9225,N_10165);
nor U11220 (N_11220,N_10134,N_9159);
nor U11221 (N_11221,N_9775,N_9098);
nor U11222 (N_11222,N_9959,N_10242);
nand U11223 (N_11223,N_9032,N_10009);
and U11224 (N_11224,N_9886,N_10237);
xor U11225 (N_11225,N_9688,N_9199);
and U11226 (N_11226,N_10233,N_9679);
and U11227 (N_11227,N_9407,N_9666);
and U11228 (N_11228,N_9248,N_9170);
nand U11229 (N_11229,N_9703,N_9207);
xor U11230 (N_11230,N_9559,N_9560);
nand U11231 (N_11231,N_9887,N_10363);
or U11232 (N_11232,N_9925,N_9051);
and U11233 (N_11233,N_9590,N_9502);
nand U11234 (N_11234,N_10488,N_9168);
xor U11235 (N_11235,N_9789,N_9130);
nor U11236 (N_11236,N_9050,N_9897);
xor U11237 (N_11237,N_9545,N_9932);
or U11238 (N_11238,N_9622,N_9310);
xnor U11239 (N_11239,N_9444,N_10221);
nand U11240 (N_11240,N_9256,N_9214);
nand U11241 (N_11241,N_9270,N_10264);
and U11242 (N_11242,N_9610,N_9305);
nor U11243 (N_11243,N_10121,N_9027);
nor U11244 (N_11244,N_10372,N_10399);
or U11245 (N_11245,N_9379,N_9509);
xnor U11246 (N_11246,N_9415,N_9611);
or U11247 (N_11247,N_10257,N_10199);
nand U11248 (N_11248,N_10099,N_10431);
nor U11249 (N_11249,N_9384,N_9960);
xnor U11250 (N_11250,N_10017,N_9247);
nand U11251 (N_11251,N_9038,N_10203);
xnor U11252 (N_11252,N_9729,N_9000);
and U11253 (N_11253,N_9438,N_9884);
and U11254 (N_11254,N_9971,N_9301);
xor U11255 (N_11255,N_10224,N_10204);
nor U11256 (N_11256,N_9005,N_9462);
xor U11257 (N_11257,N_9839,N_9250);
nor U11258 (N_11258,N_9244,N_10365);
or U11259 (N_11259,N_9854,N_10369);
or U11260 (N_11260,N_9166,N_9148);
nor U11261 (N_11261,N_9841,N_9035);
nand U11262 (N_11262,N_9134,N_9828);
and U11263 (N_11263,N_9936,N_10021);
xnor U11264 (N_11264,N_9072,N_9529);
xor U11265 (N_11265,N_9462,N_10042);
or U11266 (N_11266,N_9986,N_9234);
and U11267 (N_11267,N_9876,N_9748);
or U11268 (N_11268,N_10094,N_10227);
nor U11269 (N_11269,N_9800,N_9868);
and U11270 (N_11270,N_9781,N_10093);
nand U11271 (N_11271,N_9185,N_9648);
nor U11272 (N_11272,N_9833,N_9665);
nor U11273 (N_11273,N_10394,N_9402);
and U11274 (N_11274,N_9661,N_10250);
nor U11275 (N_11275,N_9855,N_10379);
or U11276 (N_11276,N_10428,N_9406);
nand U11277 (N_11277,N_9907,N_10241);
nand U11278 (N_11278,N_10098,N_9433);
nand U11279 (N_11279,N_9048,N_10241);
nor U11280 (N_11280,N_9618,N_9272);
nand U11281 (N_11281,N_9758,N_10053);
xnor U11282 (N_11282,N_9282,N_9519);
and U11283 (N_11283,N_10033,N_9005);
xnor U11284 (N_11284,N_9476,N_9621);
or U11285 (N_11285,N_10002,N_9612);
xnor U11286 (N_11286,N_9262,N_9319);
or U11287 (N_11287,N_9522,N_9132);
nand U11288 (N_11288,N_10131,N_10416);
xnor U11289 (N_11289,N_9145,N_9127);
or U11290 (N_11290,N_9596,N_9801);
nand U11291 (N_11291,N_10167,N_10227);
nor U11292 (N_11292,N_9566,N_9410);
xor U11293 (N_11293,N_10016,N_10187);
and U11294 (N_11294,N_9256,N_9224);
or U11295 (N_11295,N_9531,N_10488);
or U11296 (N_11296,N_9701,N_9577);
or U11297 (N_11297,N_9485,N_9166);
and U11298 (N_11298,N_9060,N_9023);
or U11299 (N_11299,N_9537,N_9030);
xnor U11300 (N_11300,N_9281,N_9473);
xor U11301 (N_11301,N_9288,N_10261);
xor U11302 (N_11302,N_10107,N_10312);
and U11303 (N_11303,N_9931,N_10315);
nand U11304 (N_11304,N_10464,N_9970);
nand U11305 (N_11305,N_9017,N_10038);
nor U11306 (N_11306,N_9840,N_9839);
nor U11307 (N_11307,N_10343,N_9129);
or U11308 (N_11308,N_9366,N_10447);
nand U11309 (N_11309,N_9838,N_10208);
nand U11310 (N_11310,N_9585,N_9581);
and U11311 (N_11311,N_9547,N_9869);
and U11312 (N_11312,N_9473,N_9165);
xor U11313 (N_11313,N_9487,N_9811);
or U11314 (N_11314,N_9396,N_9259);
and U11315 (N_11315,N_9702,N_9317);
nand U11316 (N_11316,N_10138,N_10294);
or U11317 (N_11317,N_10304,N_9877);
or U11318 (N_11318,N_9842,N_9359);
xor U11319 (N_11319,N_9393,N_10263);
nand U11320 (N_11320,N_9155,N_9017);
nor U11321 (N_11321,N_10393,N_10283);
nor U11322 (N_11322,N_10481,N_9934);
or U11323 (N_11323,N_9908,N_10486);
xor U11324 (N_11324,N_9015,N_10173);
or U11325 (N_11325,N_9888,N_9602);
xnor U11326 (N_11326,N_9287,N_9172);
nand U11327 (N_11327,N_9920,N_10263);
and U11328 (N_11328,N_9753,N_9805);
or U11329 (N_11329,N_9844,N_9006);
or U11330 (N_11330,N_9375,N_9503);
or U11331 (N_11331,N_9327,N_9606);
or U11332 (N_11332,N_10109,N_10215);
or U11333 (N_11333,N_10024,N_9238);
nand U11334 (N_11334,N_9189,N_10134);
and U11335 (N_11335,N_10230,N_10413);
nand U11336 (N_11336,N_9524,N_9832);
or U11337 (N_11337,N_10172,N_9755);
and U11338 (N_11338,N_9912,N_9657);
nand U11339 (N_11339,N_9774,N_9275);
or U11340 (N_11340,N_10435,N_9126);
nand U11341 (N_11341,N_9298,N_10202);
nand U11342 (N_11342,N_9795,N_9105);
and U11343 (N_11343,N_9068,N_9405);
nor U11344 (N_11344,N_9062,N_9728);
nand U11345 (N_11345,N_10246,N_9503);
nand U11346 (N_11346,N_10065,N_9770);
nand U11347 (N_11347,N_10213,N_10468);
or U11348 (N_11348,N_10429,N_9113);
xor U11349 (N_11349,N_9671,N_9871);
nand U11350 (N_11350,N_9900,N_9609);
nor U11351 (N_11351,N_9464,N_10165);
and U11352 (N_11352,N_9629,N_9358);
nand U11353 (N_11353,N_9779,N_9218);
nand U11354 (N_11354,N_9777,N_9702);
and U11355 (N_11355,N_9574,N_9069);
and U11356 (N_11356,N_9746,N_9530);
nor U11357 (N_11357,N_10247,N_9778);
nand U11358 (N_11358,N_9318,N_10073);
and U11359 (N_11359,N_10346,N_9803);
and U11360 (N_11360,N_10268,N_9995);
nor U11361 (N_11361,N_9192,N_9590);
nor U11362 (N_11362,N_10014,N_9219);
xor U11363 (N_11363,N_10222,N_9253);
nor U11364 (N_11364,N_10336,N_10361);
xnor U11365 (N_11365,N_9185,N_9199);
xor U11366 (N_11366,N_9495,N_10085);
xnor U11367 (N_11367,N_10257,N_10104);
xor U11368 (N_11368,N_9090,N_10394);
and U11369 (N_11369,N_9819,N_9082);
and U11370 (N_11370,N_9465,N_10180);
or U11371 (N_11371,N_9125,N_10145);
and U11372 (N_11372,N_10040,N_9546);
xor U11373 (N_11373,N_9375,N_9451);
xnor U11374 (N_11374,N_9927,N_9183);
nand U11375 (N_11375,N_10492,N_9007);
xor U11376 (N_11376,N_10242,N_9777);
or U11377 (N_11377,N_9647,N_9600);
or U11378 (N_11378,N_10286,N_9832);
or U11379 (N_11379,N_9241,N_9892);
xnor U11380 (N_11380,N_9773,N_10102);
xor U11381 (N_11381,N_10271,N_9036);
xor U11382 (N_11382,N_10316,N_10271);
or U11383 (N_11383,N_9278,N_9220);
or U11384 (N_11384,N_9267,N_9948);
nor U11385 (N_11385,N_10499,N_9254);
and U11386 (N_11386,N_9109,N_9770);
or U11387 (N_11387,N_10454,N_10118);
and U11388 (N_11388,N_9035,N_9547);
nand U11389 (N_11389,N_10096,N_9065);
and U11390 (N_11390,N_9247,N_9934);
xor U11391 (N_11391,N_9420,N_9940);
nor U11392 (N_11392,N_10457,N_10296);
or U11393 (N_11393,N_10273,N_9274);
nand U11394 (N_11394,N_9940,N_10457);
or U11395 (N_11395,N_9517,N_9882);
xnor U11396 (N_11396,N_9374,N_10332);
and U11397 (N_11397,N_9092,N_10243);
nand U11398 (N_11398,N_10450,N_9559);
and U11399 (N_11399,N_10156,N_9504);
and U11400 (N_11400,N_9747,N_9599);
nand U11401 (N_11401,N_10337,N_9737);
nand U11402 (N_11402,N_10440,N_10481);
xor U11403 (N_11403,N_10022,N_9968);
and U11404 (N_11404,N_9641,N_9325);
nand U11405 (N_11405,N_10153,N_9305);
nor U11406 (N_11406,N_10331,N_10243);
nor U11407 (N_11407,N_10256,N_9478);
or U11408 (N_11408,N_9977,N_9166);
nand U11409 (N_11409,N_10347,N_10202);
or U11410 (N_11410,N_10356,N_9126);
and U11411 (N_11411,N_10203,N_9117);
and U11412 (N_11412,N_10367,N_9108);
nor U11413 (N_11413,N_9834,N_9078);
nor U11414 (N_11414,N_9809,N_9444);
xnor U11415 (N_11415,N_9382,N_9363);
and U11416 (N_11416,N_10143,N_9078);
xnor U11417 (N_11417,N_9736,N_10438);
or U11418 (N_11418,N_10023,N_9073);
or U11419 (N_11419,N_9953,N_10075);
and U11420 (N_11420,N_9115,N_10484);
nor U11421 (N_11421,N_9237,N_10001);
nor U11422 (N_11422,N_10404,N_10252);
nand U11423 (N_11423,N_10171,N_9525);
xnor U11424 (N_11424,N_10498,N_10328);
and U11425 (N_11425,N_9107,N_10459);
nor U11426 (N_11426,N_9898,N_10249);
nor U11427 (N_11427,N_10357,N_10381);
and U11428 (N_11428,N_9749,N_10352);
nor U11429 (N_11429,N_9674,N_9284);
nor U11430 (N_11430,N_9159,N_9044);
or U11431 (N_11431,N_9882,N_9338);
nand U11432 (N_11432,N_9097,N_9364);
nand U11433 (N_11433,N_9926,N_9870);
and U11434 (N_11434,N_9391,N_9373);
or U11435 (N_11435,N_9988,N_10163);
nor U11436 (N_11436,N_10307,N_10348);
and U11437 (N_11437,N_9778,N_9677);
nor U11438 (N_11438,N_10498,N_10117);
and U11439 (N_11439,N_9764,N_9366);
nand U11440 (N_11440,N_9166,N_9312);
or U11441 (N_11441,N_9825,N_9065);
or U11442 (N_11442,N_9644,N_9170);
and U11443 (N_11443,N_9253,N_10306);
nand U11444 (N_11444,N_10116,N_9672);
nor U11445 (N_11445,N_9631,N_9974);
nand U11446 (N_11446,N_10007,N_9861);
or U11447 (N_11447,N_10104,N_9842);
and U11448 (N_11448,N_9060,N_9330);
nand U11449 (N_11449,N_9148,N_10158);
or U11450 (N_11450,N_10409,N_9858);
nor U11451 (N_11451,N_10428,N_10300);
or U11452 (N_11452,N_9828,N_9868);
nand U11453 (N_11453,N_10201,N_10339);
nand U11454 (N_11454,N_10256,N_10286);
nand U11455 (N_11455,N_9191,N_9145);
or U11456 (N_11456,N_9380,N_9761);
and U11457 (N_11457,N_10127,N_9553);
or U11458 (N_11458,N_9674,N_9925);
nor U11459 (N_11459,N_9676,N_9388);
xnor U11460 (N_11460,N_10081,N_9266);
nand U11461 (N_11461,N_9085,N_10470);
nor U11462 (N_11462,N_10224,N_9344);
and U11463 (N_11463,N_9834,N_10122);
nand U11464 (N_11464,N_10409,N_10077);
nand U11465 (N_11465,N_9338,N_9931);
xnor U11466 (N_11466,N_9792,N_10227);
or U11467 (N_11467,N_10274,N_10332);
nor U11468 (N_11468,N_10143,N_10351);
nand U11469 (N_11469,N_9451,N_10038);
nor U11470 (N_11470,N_9531,N_9905);
and U11471 (N_11471,N_10459,N_9907);
nand U11472 (N_11472,N_9179,N_10115);
xor U11473 (N_11473,N_9716,N_10356);
xnor U11474 (N_11474,N_10309,N_9099);
or U11475 (N_11475,N_10305,N_9889);
nand U11476 (N_11476,N_9660,N_10138);
nand U11477 (N_11477,N_10373,N_9167);
or U11478 (N_11478,N_9495,N_10425);
xnor U11479 (N_11479,N_10263,N_9266);
xnor U11480 (N_11480,N_9338,N_9621);
xor U11481 (N_11481,N_10179,N_10351);
nand U11482 (N_11482,N_9811,N_10320);
and U11483 (N_11483,N_10322,N_10372);
or U11484 (N_11484,N_10171,N_9003);
nand U11485 (N_11485,N_9834,N_10457);
nand U11486 (N_11486,N_9996,N_9801);
nand U11487 (N_11487,N_9316,N_9235);
and U11488 (N_11488,N_9631,N_10053);
and U11489 (N_11489,N_9816,N_10459);
nor U11490 (N_11490,N_10187,N_9616);
xor U11491 (N_11491,N_9914,N_9297);
nand U11492 (N_11492,N_9034,N_9096);
nand U11493 (N_11493,N_9648,N_10092);
nor U11494 (N_11494,N_9294,N_9504);
nand U11495 (N_11495,N_10459,N_9376);
xor U11496 (N_11496,N_9082,N_10010);
and U11497 (N_11497,N_9083,N_9959);
xnor U11498 (N_11498,N_9689,N_9580);
nand U11499 (N_11499,N_9799,N_9490);
xnor U11500 (N_11500,N_9587,N_10476);
nand U11501 (N_11501,N_9578,N_10119);
and U11502 (N_11502,N_9850,N_10051);
or U11503 (N_11503,N_9560,N_9127);
and U11504 (N_11504,N_9812,N_9074);
xor U11505 (N_11505,N_9199,N_9968);
and U11506 (N_11506,N_9920,N_9204);
and U11507 (N_11507,N_9018,N_9473);
nand U11508 (N_11508,N_9892,N_9470);
or U11509 (N_11509,N_10444,N_10020);
xor U11510 (N_11510,N_10386,N_10104);
and U11511 (N_11511,N_10126,N_9409);
or U11512 (N_11512,N_9395,N_9886);
or U11513 (N_11513,N_9689,N_10200);
xor U11514 (N_11514,N_9413,N_9629);
and U11515 (N_11515,N_9120,N_9979);
nor U11516 (N_11516,N_9246,N_10261);
xnor U11517 (N_11517,N_10035,N_9323);
nor U11518 (N_11518,N_9354,N_9904);
or U11519 (N_11519,N_10301,N_9723);
nand U11520 (N_11520,N_9769,N_9479);
or U11521 (N_11521,N_10133,N_9813);
nor U11522 (N_11522,N_9807,N_9137);
nand U11523 (N_11523,N_10024,N_10478);
and U11524 (N_11524,N_10458,N_9948);
and U11525 (N_11525,N_10105,N_9810);
xnor U11526 (N_11526,N_9947,N_9112);
and U11527 (N_11527,N_9877,N_10414);
or U11528 (N_11528,N_10135,N_9886);
nand U11529 (N_11529,N_10039,N_9830);
or U11530 (N_11530,N_9024,N_9553);
xnor U11531 (N_11531,N_9347,N_10094);
xor U11532 (N_11532,N_10102,N_10377);
or U11533 (N_11533,N_9976,N_9864);
and U11534 (N_11534,N_9488,N_9622);
and U11535 (N_11535,N_9522,N_9394);
nand U11536 (N_11536,N_9920,N_10499);
nand U11537 (N_11537,N_10180,N_9695);
nand U11538 (N_11538,N_9279,N_10176);
or U11539 (N_11539,N_10442,N_9737);
nor U11540 (N_11540,N_10078,N_9105);
and U11541 (N_11541,N_9389,N_10445);
xnor U11542 (N_11542,N_9421,N_9978);
nor U11543 (N_11543,N_9823,N_9879);
nor U11544 (N_11544,N_10250,N_9641);
xor U11545 (N_11545,N_10351,N_9340);
and U11546 (N_11546,N_9921,N_9930);
nand U11547 (N_11547,N_10427,N_9389);
or U11548 (N_11548,N_10134,N_9209);
and U11549 (N_11549,N_9566,N_9880);
nor U11550 (N_11550,N_9732,N_9892);
and U11551 (N_11551,N_9700,N_9497);
nor U11552 (N_11552,N_10263,N_10445);
nand U11553 (N_11553,N_9494,N_10303);
and U11554 (N_11554,N_10336,N_10266);
and U11555 (N_11555,N_9632,N_9559);
or U11556 (N_11556,N_9161,N_10388);
xnor U11557 (N_11557,N_9217,N_10169);
and U11558 (N_11558,N_9756,N_10400);
nor U11559 (N_11559,N_10080,N_9887);
xnor U11560 (N_11560,N_9893,N_9128);
nand U11561 (N_11561,N_9966,N_9288);
and U11562 (N_11562,N_10350,N_10125);
and U11563 (N_11563,N_10384,N_10026);
nand U11564 (N_11564,N_10104,N_10441);
nand U11565 (N_11565,N_9596,N_9873);
or U11566 (N_11566,N_9396,N_9075);
or U11567 (N_11567,N_10224,N_10098);
nand U11568 (N_11568,N_10427,N_9917);
xnor U11569 (N_11569,N_9571,N_10006);
xor U11570 (N_11570,N_9317,N_9713);
nor U11571 (N_11571,N_10264,N_10053);
and U11572 (N_11572,N_9021,N_9237);
nor U11573 (N_11573,N_10425,N_9911);
and U11574 (N_11574,N_9621,N_9163);
nor U11575 (N_11575,N_9917,N_9519);
nand U11576 (N_11576,N_9463,N_9948);
xor U11577 (N_11577,N_10319,N_9326);
nand U11578 (N_11578,N_10153,N_9889);
nor U11579 (N_11579,N_9439,N_9349);
or U11580 (N_11580,N_10314,N_10492);
nor U11581 (N_11581,N_9024,N_10209);
nor U11582 (N_11582,N_9892,N_9716);
nand U11583 (N_11583,N_9169,N_10125);
xnor U11584 (N_11584,N_9894,N_10237);
or U11585 (N_11585,N_9304,N_9992);
nand U11586 (N_11586,N_10227,N_9312);
and U11587 (N_11587,N_10422,N_10124);
or U11588 (N_11588,N_10142,N_9504);
or U11589 (N_11589,N_9677,N_9422);
or U11590 (N_11590,N_9089,N_10335);
nand U11591 (N_11591,N_10102,N_9351);
xor U11592 (N_11592,N_9194,N_9277);
nor U11593 (N_11593,N_10438,N_9416);
or U11594 (N_11594,N_10314,N_9958);
and U11595 (N_11595,N_9382,N_10466);
xor U11596 (N_11596,N_9786,N_9440);
xor U11597 (N_11597,N_9677,N_9456);
xnor U11598 (N_11598,N_9539,N_9220);
nand U11599 (N_11599,N_9271,N_10272);
or U11600 (N_11600,N_9715,N_10001);
and U11601 (N_11601,N_9736,N_10065);
nor U11602 (N_11602,N_9230,N_9275);
xor U11603 (N_11603,N_9283,N_9212);
and U11604 (N_11604,N_10240,N_9935);
and U11605 (N_11605,N_9003,N_9474);
xnor U11606 (N_11606,N_10310,N_9996);
and U11607 (N_11607,N_9932,N_9429);
or U11608 (N_11608,N_9683,N_10139);
nand U11609 (N_11609,N_10203,N_9889);
and U11610 (N_11610,N_9073,N_9430);
and U11611 (N_11611,N_9519,N_9033);
nor U11612 (N_11612,N_10273,N_9075);
nor U11613 (N_11613,N_9827,N_9564);
or U11614 (N_11614,N_9994,N_9039);
xnor U11615 (N_11615,N_9271,N_9305);
nand U11616 (N_11616,N_10137,N_10035);
and U11617 (N_11617,N_10077,N_9646);
xnor U11618 (N_11618,N_10465,N_9465);
xnor U11619 (N_11619,N_9172,N_9171);
or U11620 (N_11620,N_9224,N_9798);
nor U11621 (N_11621,N_9335,N_10100);
xor U11622 (N_11622,N_9148,N_10144);
or U11623 (N_11623,N_9804,N_9835);
nand U11624 (N_11624,N_10156,N_9629);
or U11625 (N_11625,N_9157,N_10145);
xor U11626 (N_11626,N_9942,N_10271);
and U11627 (N_11627,N_9592,N_9706);
or U11628 (N_11628,N_10042,N_10115);
and U11629 (N_11629,N_9924,N_9782);
nor U11630 (N_11630,N_10185,N_9254);
nand U11631 (N_11631,N_9978,N_9086);
and U11632 (N_11632,N_9208,N_9458);
nand U11633 (N_11633,N_10215,N_9817);
or U11634 (N_11634,N_10044,N_9642);
nand U11635 (N_11635,N_9392,N_10186);
and U11636 (N_11636,N_10216,N_9492);
nor U11637 (N_11637,N_9904,N_9554);
nand U11638 (N_11638,N_9443,N_10120);
and U11639 (N_11639,N_9826,N_10353);
xor U11640 (N_11640,N_9901,N_9401);
nand U11641 (N_11641,N_9623,N_9600);
xnor U11642 (N_11642,N_9827,N_9957);
or U11643 (N_11643,N_9302,N_10316);
and U11644 (N_11644,N_9116,N_10455);
or U11645 (N_11645,N_9798,N_10053);
and U11646 (N_11646,N_9383,N_9039);
or U11647 (N_11647,N_9406,N_9216);
and U11648 (N_11648,N_10407,N_9108);
and U11649 (N_11649,N_9680,N_9139);
nand U11650 (N_11650,N_9853,N_9419);
and U11651 (N_11651,N_10445,N_10479);
xor U11652 (N_11652,N_9732,N_10284);
nor U11653 (N_11653,N_9961,N_9789);
nor U11654 (N_11654,N_9706,N_9764);
nand U11655 (N_11655,N_9332,N_9177);
nor U11656 (N_11656,N_9331,N_9499);
and U11657 (N_11657,N_10021,N_9645);
nor U11658 (N_11658,N_10146,N_9392);
or U11659 (N_11659,N_9826,N_9917);
and U11660 (N_11660,N_9885,N_10065);
nand U11661 (N_11661,N_9819,N_9017);
xnor U11662 (N_11662,N_9028,N_9140);
and U11663 (N_11663,N_9153,N_9854);
xor U11664 (N_11664,N_10116,N_10026);
and U11665 (N_11665,N_9807,N_9567);
and U11666 (N_11666,N_9136,N_9127);
nand U11667 (N_11667,N_10189,N_10118);
and U11668 (N_11668,N_10292,N_10318);
and U11669 (N_11669,N_9297,N_10445);
xnor U11670 (N_11670,N_9021,N_10209);
and U11671 (N_11671,N_9749,N_9152);
xnor U11672 (N_11672,N_10143,N_10114);
nor U11673 (N_11673,N_9040,N_9980);
and U11674 (N_11674,N_9524,N_10204);
and U11675 (N_11675,N_9763,N_10247);
nand U11676 (N_11676,N_9213,N_9966);
xnor U11677 (N_11677,N_9846,N_9415);
xor U11678 (N_11678,N_9599,N_10483);
xnor U11679 (N_11679,N_9325,N_9229);
nor U11680 (N_11680,N_9813,N_10472);
and U11681 (N_11681,N_9029,N_9766);
xor U11682 (N_11682,N_9113,N_10010);
xor U11683 (N_11683,N_10063,N_9241);
and U11684 (N_11684,N_9010,N_10463);
nand U11685 (N_11685,N_9994,N_9145);
xnor U11686 (N_11686,N_9908,N_9726);
nor U11687 (N_11687,N_9094,N_9007);
xor U11688 (N_11688,N_9810,N_10012);
or U11689 (N_11689,N_9320,N_9239);
or U11690 (N_11690,N_9634,N_9047);
xnor U11691 (N_11691,N_9262,N_10347);
xnor U11692 (N_11692,N_10402,N_10147);
and U11693 (N_11693,N_9228,N_9520);
nor U11694 (N_11694,N_9594,N_9665);
nor U11695 (N_11695,N_9841,N_9080);
xnor U11696 (N_11696,N_9536,N_9825);
nand U11697 (N_11697,N_10080,N_10245);
and U11698 (N_11698,N_9442,N_10170);
and U11699 (N_11699,N_9692,N_10184);
xor U11700 (N_11700,N_9450,N_9773);
nand U11701 (N_11701,N_10262,N_9478);
and U11702 (N_11702,N_9167,N_9247);
nor U11703 (N_11703,N_9393,N_9745);
nor U11704 (N_11704,N_9879,N_9620);
or U11705 (N_11705,N_9723,N_9857);
xor U11706 (N_11706,N_10279,N_9582);
xor U11707 (N_11707,N_10452,N_9218);
nor U11708 (N_11708,N_9939,N_9924);
and U11709 (N_11709,N_10387,N_9085);
nor U11710 (N_11710,N_9380,N_9265);
xnor U11711 (N_11711,N_9108,N_9935);
xnor U11712 (N_11712,N_10406,N_10060);
nand U11713 (N_11713,N_9000,N_9573);
and U11714 (N_11714,N_9565,N_9661);
xor U11715 (N_11715,N_9477,N_10240);
or U11716 (N_11716,N_9166,N_9935);
nand U11717 (N_11717,N_10311,N_9061);
or U11718 (N_11718,N_9843,N_10150);
xor U11719 (N_11719,N_9279,N_9099);
nand U11720 (N_11720,N_10180,N_9789);
nand U11721 (N_11721,N_9288,N_9715);
and U11722 (N_11722,N_9720,N_10057);
nand U11723 (N_11723,N_10106,N_9557);
or U11724 (N_11724,N_9327,N_10378);
xnor U11725 (N_11725,N_9064,N_9090);
nor U11726 (N_11726,N_10484,N_9857);
and U11727 (N_11727,N_9018,N_9869);
xor U11728 (N_11728,N_10326,N_9482);
nor U11729 (N_11729,N_9225,N_9826);
nor U11730 (N_11730,N_10088,N_10234);
xor U11731 (N_11731,N_9124,N_9114);
nand U11732 (N_11732,N_10497,N_10013);
xnor U11733 (N_11733,N_10420,N_9015);
nor U11734 (N_11734,N_9112,N_10333);
and U11735 (N_11735,N_9387,N_9995);
xor U11736 (N_11736,N_9422,N_10266);
xor U11737 (N_11737,N_9270,N_9568);
nor U11738 (N_11738,N_9085,N_9922);
nor U11739 (N_11739,N_9638,N_9867);
xor U11740 (N_11740,N_9255,N_9298);
nand U11741 (N_11741,N_10274,N_10154);
and U11742 (N_11742,N_9411,N_10401);
or U11743 (N_11743,N_9685,N_10465);
or U11744 (N_11744,N_9340,N_10136);
nor U11745 (N_11745,N_9000,N_9597);
nand U11746 (N_11746,N_10046,N_10476);
nand U11747 (N_11747,N_9990,N_9903);
nand U11748 (N_11748,N_10235,N_9163);
or U11749 (N_11749,N_9790,N_9053);
xnor U11750 (N_11750,N_9929,N_9968);
xor U11751 (N_11751,N_9353,N_9584);
or U11752 (N_11752,N_10356,N_10324);
or U11753 (N_11753,N_10376,N_10137);
nor U11754 (N_11754,N_9460,N_9021);
xor U11755 (N_11755,N_10265,N_9144);
nor U11756 (N_11756,N_10032,N_9035);
nor U11757 (N_11757,N_9720,N_9035);
xnor U11758 (N_11758,N_9557,N_10085);
nor U11759 (N_11759,N_9777,N_9497);
and U11760 (N_11760,N_10220,N_9661);
nor U11761 (N_11761,N_10125,N_9618);
or U11762 (N_11762,N_9763,N_10161);
xor U11763 (N_11763,N_9579,N_9092);
xor U11764 (N_11764,N_9598,N_9585);
xnor U11765 (N_11765,N_9396,N_9250);
nand U11766 (N_11766,N_10052,N_10131);
nor U11767 (N_11767,N_9272,N_10310);
nor U11768 (N_11768,N_10449,N_10065);
nand U11769 (N_11769,N_10331,N_9814);
or U11770 (N_11770,N_9838,N_9407);
xor U11771 (N_11771,N_9341,N_9657);
and U11772 (N_11772,N_9886,N_9493);
and U11773 (N_11773,N_9973,N_10410);
nand U11774 (N_11774,N_10442,N_10255);
xnor U11775 (N_11775,N_10419,N_10278);
nand U11776 (N_11776,N_10248,N_9707);
and U11777 (N_11777,N_9192,N_9385);
xor U11778 (N_11778,N_9268,N_9053);
and U11779 (N_11779,N_9937,N_9579);
nand U11780 (N_11780,N_9788,N_9292);
and U11781 (N_11781,N_10164,N_9585);
xnor U11782 (N_11782,N_9842,N_10386);
nor U11783 (N_11783,N_10211,N_9906);
nor U11784 (N_11784,N_9851,N_9767);
xnor U11785 (N_11785,N_9885,N_9247);
nand U11786 (N_11786,N_9920,N_9243);
or U11787 (N_11787,N_9535,N_10158);
and U11788 (N_11788,N_10165,N_9293);
and U11789 (N_11789,N_9010,N_9220);
nand U11790 (N_11790,N_9778,N_10408);
nor U11791 (N_11791,N_9455,N_9612);
nor U11792 (N_11792,N_10228,N_10222);
nand U11793 (N_11793,N_10176,N_9317);
nor U11794 (N_11794,N_9467,N_10039);
nor U11795 (N_11795,N_9565,N_9256);
xor U11796 (N_11796,N_10221,N_10041);
nand U11797 (N_11797,N_9107,N_10425);
xnor U11798 (N_11798,N_9244,N_9850);
nor U11799 (N_11799,N_9735,N_9850);
xnor U11800 (N_11800,N_9286,N_10036);
or U11801 (N_11801,N_9328,N_9380);
xnor U11802 (N_11802,N_10238,N_9464);
nor U11803 (N_11803,N_10298,N_9355);
or U11804 (N_11804,N_9532,N_9069);
or U11805 (N_11805,N_9488,N_9764);
or U11806 (N_11806,N_10411,N_10463);
nand U11807 (N_11807,N_10240,N_9109);
xor U11808 (N_11808,N_9683,N_10311);
nand U11809 (N_11809,N_10350,N_9682);
or U11810 (N_11810,N_9973,N_10372);
and U11811 (N_11811,N_10069,N_10361);
xnor U11812 (N_11812,N_9741,N_10100);
or U11813 (N_11813,N_9137,N_9368);
and U11814 (N_11814,N_9765,N_9743);
and U11815 (N_11815,N_9820,N_9896);
and U11816 (N_11816,N_9296,N_9166);
and U11817 (N_11817,N_9728,N_10451);
nand U11818 (N_11818,N_10250,N_10001);
xnor U11819 (N_11819,N_10469,N_10087);
xnor U11820 (N_11820,N_9276,N_9543);
or U11821 (N_11821,N_10177,N_10080);
xor U11822 (N_11822,N_10487,N_9250);
or U11823 (N_11823,N_9172,N_9016);
or U11824 (N_11824,N_9138,N_9197);
nand U11825 (N_11825,N_9722,N_9898);
and U11826 (N_11826,N_10421,N_9776);
or U11827 (N_11827,N_10041,N_10134);
nor U11828 (N_11828,N_10121,N_9498);
xor U11829 (N_11829,N_10018,N_9036);
xnor U11830 (N_11830,N_10214,N_9014);
and U11831 (N_11831,N_10111,N_9464);
xnor U11832 (N_11832,N_9184,N_9798);
xor U11833 (N_11833,N_9149,N_10316);
xnor U11834 (N_11834,N_9841,N_9952);
or U11835 (N_11835,N_9341,N_10038);
or U11836 (N_11836,N_9193,N_10429);
and U11837 (N_11837,N_9902,N_9610);
and U11838 (N_11838,N_10421,N_9019);
and U11839 (N_11839,N_10373,N_9744);
nor U11840 (N_11840,N_10041,N_10448);
xnor U11841 (N_11841,N_9485,N_9146);
or U11842 (N_11842,N_9458,N_10112);
and U11843 (N_11843,N_10038,N_9434);
and U11844 (N_11844,N_9324,N_10154);
and U11845 (N_11845,N_9237,N_9088);
and U11846 (N_11846,N_10208,N_9853);
nor U11847 (N_11847,N_9156,N_10389);
or U11848 (N_11848,N_9605,N_10159);
nand U11849 (N_11849,N_9364,N_9435);
nand U11850 (N_11850,N_9970,N_9819);
nand U11851 (N_11851,N_9602,N_10064);
or U11852 (N_11852,N_10455,N_9468);
xnor U11853 (N_11853,N_9224,N_10292);
and U11854 (N_11854,N_10314,N_10089);
nand U11855 (N_11855,N_10019,N_10207);
and U11856 (N_11856,N_10186,N_10285);
nor U11857 (N_11857,N_10364,N_10279);
xnor U11858 (N_11858,N_9208,N_10327);
or U11859 (N_11859,N_9043,N_10293);
and U11860 (N_11860,N_9711,N_10008);
nand U11861 (N_11861,N_9400,N_9780);
nand U11862 (N_11862,N_9395,N_9374);
xnor U11863 (N_11863,N_9031,N_10448);
or U11864 (N_11864,N_10335,N_9401);
or U11865 (N_11865,N_9058,N_9041);
xor U11866 (N_11866,N_9558,N_9237);
nor U11867 (N_11867,N_9340,N_9126);
or U11868 (N_11868,N_9849,N_9964);
xor U11869 (N_11869,N_9019,N_9631);
nand U11870 (N_11870,N_10027,N_10392);
and U11871 (N_11871,N_10388,N_9711);
nand U11872 (N_11872,N_9833,N_9126);
and U11873 (N_11873,N_9958,N_10142);
and U11874 (N_11874,N_9341,N_9031);
nor U11875 (N_11875,N_9069,N_9691);
and U11876 (N_11876,N_9016,N_9547);
and U11877 (N_11877,N_10307,N_10220);
or U11878 (N_11878,N_9729,N_10122);
nor U11879 (N_11879,N_10075,N_9969);
and U11880 (N_11880,N_9156,N_10131);
xor U11881 (N_11881,N_9322,N_9676);
nor U11882 (N_11882,N_9917,N_10322);
xnor U11883 (N_11883,N_9327,N_9654);
and U11884 (N_11884,N_9339,N_9945);
nand U11885 (N_11885,N_9865,N_10179);
or U11886 (N_11886,N_9276,N_9928);
nor U11887 (N_11887,N_9842,N_9505);
or U11888 (N_11888,N_9734,N_9832);
or U11889 (N_11889,N_9773,N_10022);
or U11890 (N_11890,N_9276,N_9236);
and U11891 (N_11891,N_9103,N_9171);
nor U11892 (N_11892,N_10465,N_9132);
nor U11893 (N_11893,N_10404,N_9351);
or U11894 (N_11894,N_9404,N_9846);
and U11895 (N_11895,N_9808,N_10396);
or U11896 (N_11896,N_10136,N_10435);
nand U11897 (N_11897,N_10014,N_9156);
nor U11898 (N_11898,N_9672,N_9859);
nor U11899 (N_11899,N_9208,N_9575);
or U11900 (N_11900,N_10362,N_10016);
nand U11901 (N_11901,N_9204,N_10224);
or U11902 (N_11902,N_10490,N_10224);
nand U11903 (N_11903,N_9665,N_9376);
and U11904 (N_11904,N_10407,N_10329);
nor U11905 (N_11905,N_9931,N_9857);
or U11906 (N_11906,N_9819,N_9187);
nand U11907 (N_11907,N_9832,N_9313);
and U11908 (N_11908,N_9411,N_9559);
nor U11909 (N_11909,N_9821,N_9239);
nor U11910 (N_11910,N_9728,N_9230);
nor U11911 (N_11911,N_9014,N_9765);
or U11912 (N_11912,N_9720,N_9946);
nand U11913 (N_11913,N_10116,N_9473);
and U11914 (N_11914,N_10376,N_9345);
and U11915 (N_11915,N_9101,N_9057);
nand U11916 (N_11916,N_9039,N_10426);
or U11917 (N_11917,N_9616,N_10179);
nand U11918 (N_11918,N_9373,N_9843);
nand U11919 (N_11919,N_9123,N_9512);
and U11920 (N_11920,N_10380,N_9365);
and U11921 (N_11921,N_9577,N_10426);
nand U11922 (N_11922,N_9014,N_9717);
xor U11923 (N_11923,N_10133,N_10222);
and U11924 (N_11924,N_10392,N_9782);
xor U11925 (N_11925,N_10399,N_10355);
xnor U11926 (N_11926,N_9217,N_9025);
nand U11927 (N_11927,N_10241,N_9899);
and U11928 (N_11928,N_9941,N_10277);
nand U11929 (N_11929,N_9033,N_9002);
or U11930 (N_11930,N_9666,N_9037);
xor U11931 (N_11931,N_9664,N_9563);
nand U11932 (N_11932,N_10383,N_9615);
xor U11933 (N_11933,N_9254,N_9992);
nand U11934 (N_11934,N_10251,N_9689);
and U11935 (N_11935,N_10362,N_10035);
or U11936 (N_11936,N_10463,N_9232);
xnor U11937 (N_11937,N_10233,N_9637);
or U11938 (N_11938,N_9417,N_10354);
and U11939 (N_11939,N_10153,N_9389);
or U11940 (N_11940,N_10338,N_10399);
nor U11941 (N_11941,N_9003,N_9055);
xor U11942 (N_11942,N_9543,N_9962);
and U11943 (N_11943,N_10331,N_9050);
xnor U11944 (N_11944,N_10286,N_9968);
xor U11945 (N_11945,N_10008,N_9311);
or U11946 (N_11946,N_9236,N_9721);
xor U11947 (N_11947,N_9732,N_10346);
and U11948 (N_11948,N_9801,N_9474);
xnor U11949 (N_11949,N_9312,N_10285);
xor U11950 (N_11950,N_10243,N_9076);
or U11951 (N_11951,N_9606,N_9126);
and U11952 (N_11952,N_10216,N_9045);
nor U11953 (N_11953,N_9791,N_9056);
nor U11954 (N_11954,N_10411,N_9881);
nor U11955 (N_11955,N_9379,N_9425);
xor U11956 (N_11956,N_10091,N_9319);
xnor U11957 (N_11957,N_10313,N_10101);
and U11958 (N_11958,N_9190,N_9436);
and U11959 (N_11959,N_10196,N_9104);
and U11960 (N_11960,N_9437,N_10413);
xnor U11961 (N_11961,N_10203,N_9806);
and U11962 (N_11962,N_10078,N_9173);
and U11963 (N_11963,N_9950,N_9655);
xor U11964 (N_11964,N_9348,N_10019);
and U11965 (N_11965,N_10240,N_10378);
nor U11966 (N_11966,N_9495,N_10168);
nor U11967 (N_11967,N_9762,N_9152);
and U11968 (N_11968,N_9896,N_9166);
nor U11969 (N_11969,N_9437,N_10313);
xnor U11970 (N_11970,N_9292,N_9279);
xor U11971 (N_11971,N_9939,N_9888);
nand U11972 (N_11972,N_9658,N_9439);
or U11973 (N_11973,N_10340,N_10175);
and U11974 (N_11974,N_10179,N_10068);
xnor U11975 (N_11975,N_9959,N_9002);
nand U11976 (N_11976,N_10122,N_9599);
nand U11977 (N_11977,N_9004,N_9916);
and U11978 (N_11978,N_9790,N_10317);
nand U11979 (N_11979,N_9116,N_9505);
and U11980 (N_11980,N_10118,N_9674);
and U11981 (N_11981,N_9526,N_9035);
xnor U11982 (N_11982,N_9682,N_10220);
xor U11983 (N_11983,N_10416,N_9282);
nor U11984 (N_11984,N_10380,N_9330);
nor U11985 (N_11985,N_10416,N_10232);
nor U11986 (N_11986,N_9754,N_9742);
and U11987 (N_11987,N_10185,N_10390);
and U11988 (N_11988,N_9204,N_10099);
nor U11989 (N_11989,N_9882,N_10474);
nor U11990 (N_11990,N_9452,N_9339);
nor U11991 (N_11991,N_9467,N_10272);
xor U11992 (N_11992,N_10428,N_9366);
xor U11993 (N_11993,N_10208,N_10269);
xnor U11994 (N_11994,N_10137,N_9374);
nand U11995 (N_11995,N_9785,N_9955);
xor U11996 (N_11996,N_9619,N_9796);
nand U11997 (N_11997,N_9985,N_9548);
nor U11998 (N_11998,N_9901,N_10267);
and U11999 (N_11999,N_9563,N_9427);
and U12000 (N_12000,N_11697,N_10637);
xor U12001 (N_12001,N_11074,N_11396);
nand U12002 (N_12002,N_10501,N_11889);
or U12003 (N_12003,N_11938,N_10709);
nor U12004 (N_12004,N_11923,N_11212);
xor U12005 (N_12005,N_11080,N_11975);
nand U12006 (N_12006,N_10574,N_11307);
nand U12007 (N_12007,N_10808,N_11281);
nand U12008 (N_12008,N_11497,N_11877);
nand U12009 (N_12009,N_11252,N_11266);
nor U12010 (N_12010,N_11053,N_10803);
or U12011 (N_12011,N_10911,N_11827);
and U12012 (N_12012,N_11452,N_11614);
nor U12013 (N_12013,N_11814,N_10851);
xnor U12014 (N_12014,N_10938,N_10664);
xnor U12015 (N_12015,N_11406,N_11190);
or U12016 (N_12016,N_11071,N_10845);
and U12017 (N_12017,N_11665,N_11952);
and U12018 (N_12018,N_11059,N_10799);
nor U12019 (N_12019,N_10502,N_11234);
and U12020 (N_12020,N_11024,N_10602);
nor U12021 (N_12021,N_11692,N_11533);
nor U12022 (N_12022,N_11134,N_11639);
xor U12023 (N_12023,N_11850,N_11137);
and U12024 (N_12024,N_11143,N_10548);
or U12025 (N_12025,N_11591,N_10721);
and U12026 (N_12026,N_10766,N_10886);
and U12027 (N_12027,N_11379,N_10974);
xor U12028 (N_12028,N_11010,N_10545);
xor U12029 (N_12029,N_11690,N_10941);
nor U12030 (N_12030,N_11806,N_10642);
and U12031 (N_12031,N_11846,N_10961);
and U12032 (N_12032,N_11186,N_10777);
nor U12033 (N_12033,N_10983,N_10913);
nor U12034 (N_12034,N_10718,N_11739);
nor U12035 (N_12035,N_10677,N_10739);
or U12036 (N_12036,N_10633,N_10921);
or U12037 (N_12037,N_11661,N_11681);
nand U12038 (N_12038,N_11094,N_11855);
xor U12039 (N_12039,N_10990,N_11476);
nand U12040 (N_12040,N_11364,N_11226);
and U12041 (N_12041,N_10853,N_10940);
or U12042 (N_12042,N_11713,N_10842);
or U12043 (N_12043,N_10559,N_10641);
nand U12044 (N_12044,N_10686,N_10942);
or U12045 (N_12045,N_10634,N_11368);
xor U12046 (N_12046,N_11544,N_10922);
nor U12047 (N_12047,N_11289,N_11482);
nand U12048 (N_12048,N_10763,N_11757);
nand U12049 (N_12049,N_11508,N_10948);
or U12050 (N_12050,N_11909,N_11637);
xor U12051 (N_12051,N_11068,N_11869);
nor U12052 (N_12052,N_11560,N_11572);
nor U12053 (N_12053,N_11890,N_11898);
xnor U12054 (N_12054,N_11417,N_11125);
and U12055 (N_12055,N_10771,N_11478);
xor U12056 (N_12056,N_10910,N_11404);
nor U12057 (N_12057,N_11357,N_11087);
nor U12058 (N_12058,N_11781,N_10820);
nand U12059 (N_12059,N_11891,N_10705);
nor U12060 (N_12060,N_11774,N_11049);
and U12061 (N_12061,N_10752,N_10958);
or U12062 (N_12062,N_10629,N_11982);
or U12063 (N_12063,N_11044,N_11703);
and U12064 (N_12064,N_11521,N_11162);
or U12065 (N_12065,N_10540,N_10659);
xor U12066 (N_12066,N_10571,N_11054);
nand U12067 (N_12067,N_11386,N_11410);
xnor U12068 (N_12068,N_11383,N_10749);
nor U12069 (N_12069,N_11444,N_10952);
and U12070 (N_12070,N_11997,N_10750);
xor U12071 (N_12071,N_11841,N_11423);
nor U12072 (N_12072,N_10861,N_11193);
or U12073 (N_12073,N_10617,N_11579);
or U12074 (N_12074,N_10618,N_11012);
and U12075 (N_12075,N_11389,N_11920);
or U12076 (N_12076,N_11902,N_11412);
and U12077 (N_12077,N_11426,N_11667);
or U12078 (N_12078,N_11886,N_11896);
and U12079 (N_12079,N_11025,N_10555);
xnor U12080 (N_12080,N_11937,N_11787);
nor U12081 (N_12081,N_10524,N_10957);
xnor U12082 (N_12082,N_10514,N_11786);
or U12083 (N_12083,N_11565,N_10673);
xnor U12084 (N_12084,N_11441,N_11953);
nand U12085 (N_12085,N_10909,N_11677);
nor U12086 (N_12086,N_10863,N_11834);
nand U12087 (N_12087,N_10950,N_11618);
and U12088 (N_12088,N_11339,N_11790);
xor U12089 (N_12089,N_10830,N_10920);
nand U12090 (N_12090,N_11202,N_11459);
nor U12091 (N_12091,N_11915,N_11675);
xor U12092 (N_12092,N_11797,N_11282);
nand U12093 (N_12093,N_10773,N_11951);
and U12094 (N_12094,N_10534,N_11195);
nand U12095 (N_12095,N_10811,N_11216);
nand U12096 (N_12096,N_10683,N_11325);
nor U12097 (N_12097,N_11931,N_11556);
and U12098 (N_12098,N_10769,N_11935);
or U12099 (N_12099,N_11306,N_10562);
xnor U12100 (N_12100,N_11130,N_10969);
and U12101 (N_12101,N_10793,N_11220);
nand U12102 (N_12102,N_11812,N_11326);
xor U12103 (N_12103,N_10531,N_10724);
nand U12104 (N_12104,N_11696,N_11369);
nor U12105 (N_12105,N_11061,N_11669);
and U12106 (N_12106,N_11308,N_11081);
or U12107 (N_12107,N_10813,N_11484);
and U12108 (N_12108,N_11050,N_10682);
nor U12109 (N_12109,N_10954,N_10521);
or U12110 (N_12110,N_11399,N_11318);
and U12111 (N_12111,N_11084,N_10719);
nor U12112 (N_12112,N_11332,N_11553);
and U12113 (N_12113,N_11615,N_11187);
xnor U12114 (N_12114,N_11721,N_11179);
and U12115 (N_12115,N_11783,N_11447);
and U12116 (N_12116,N_11972,N_11392);
and U12117 (N_12117,N_11241,N_10575);
xnor U12118 (N_12118,N_10668,N_11780);
xor U12119 (N_12119,N_11973,N_10876);
or U12120 (N_12120,N_10888,N_11839);
and U12121 (N_12121,N_10966,N_11321);
xnor U12122 (N_12122,N_11005,N_11062);
nand U12123 (N_12123,N_11494,N_11117);
nor U12124 (N_12124,N_11983,N_11227);
nor U12125 (N_12125,N_10850,N_10947);
or U12126 (N_12126,N_11448,N_11501);
or U12127 (N_12127,N_11057,N_11424);
nor U12128 (N_12128,N_11726,N_11156);
xor U12129 (N_12129,N_11142,N_11279);
and U12130 (N_12130,N_11322,N_11122);
xor U12131 (N_12131,N_11990,N_11330);
and U12132 (N_12132,N_11633,N_11178);
and U12133 (N_12133,N_10512,N_11925);
and U12134 (N_12134,N_10836,N_11225);
or U12135 (N_12135,N_11722,N_11414);
or U12136 (N_12136,N_10585,N_11901);
nor U12137 (N_12137,N_10840,N_11916);
xor U12138 (N_12138,N_11425,N_11033);
nor U12139 (N_12139,N_11845,N_11040);
xnor U12140 (N_12140,N_10572,N_11286);
and U12141 (N_12141,N_11168,N_11837);
nand U12142 (N_12142,N_10993,N_10879);
nor U12143 (N_12143,N_11601,N_11177);
or U12144 (N_12144,N_11408,N_11163);
and U12145 (N_12145,N_10680,N_11014);
or U12146 (N_12146,N_11471,N_11802);
xor U12147 (N_12147,N_11658,N_11748);
or U12148 (N_12148,N_10848,N_11950);
and U12149 (N_12149,N_11235,N_11535);
and U12150 (N_12150,N_10784,N_11984);
xnor U12151 (N_12151,N_11843,N_11347);
or U12152 (N_12152,N_10726,N_11752);
nand U12153 (N_12153,N_11345,N_11201);
nor U12154 (N_12154,N_10511,N_11641);
and U12155 (N_12155,N_11016,N_11131);
xor U12156 (N_12156,N_10797,N_11929);
and U12157 (N_12157,N_11430,N_11320);
nor U12158 (N_12158,N_11934,N_11680);
and U12159 (N_12159,N_10608,N_10939);
nand U12160 (N_12160,N_11564,N_11968);
nand U12161 (N_12161,N_11099,N_11547);
or U12162 (N_12162,N_11336,N_11007);
nand U12163 (N_12163,N_11461,N_10729);
and U12164 (N_12164,N_11363,N_11283);
nor U12165 (N_12165,N_11815,N_11582);
nor U12166 (N_12166,N_11836,N_10734);
nand U12167 (N_12167,N_10662,N_11340);
nand U12168 (N_12168,N_10785,N_11872);
nand U12169 (N_12169,N_10589,N_11686);
xor U12170 (N_12170,N_10880,N_10755);
or U12171 (N_12171,N_10866,N_11782);
nor U12172 (N_12172,N_11362,N_11958);
nor U12173 (N_12173,N_11903,N_11470);
or U12174 (N_12174,N_11096,N_11894);
and U12175 (N_12175,N_11867,N_11769);
nor U12176 (N_12176,N_11715,N_11491);
nand U12177 (N_12177,N_11173,N_10651);
xor U12178 (N_12178,N_10944,N_11439);
nand U12179 (N_12179,N_11807,N_10706);
xor U12180 (N_12180,N_10544,N_10523);
nand U12181 (N_12181,N_11954,N_11718);
nor U12182 (N_12182,N_11302,N_10537);
and U12183 (N_12183,N_11558,N_11645);
nor U12184 (N_12184,N_10834,N_10529);
or U12185 (N_12185,N_10945,N_11371);
and U12186 (N_12186,N_11421,N_11671);
xor U12187 (N_12187,N_11003,N_10566);
or U12188 (N_12188,N_11924,N_11531);
and U12189 (N_12189,N_11128,N_11454);
or U12190 (N_12190,N_11192,N_10871);
or U12191 (N_12191,N_11828,N_11204);
or U12192 (N_12192,N_11239,N_11659);
or U12193 (N_12193,N_11039,N_11303);
nand U12194 (N_12194,N_10991,N_11875);
nor U12195 (N_12195,N_10713,N_11811);
or U12196 (N_12196,N_11546,N_10758);
and U12197 (N_12197,N_11309,N_10774);
or U12198 (N_12198,N_11545,N_10963);
or U12199 (N_12199,N_10789,N_11067);
xor U12200 (N_12200,N_11754,N_11211);
or U12201 (N_12201,N_11413,N_10747);
or U12202 (N_12202,N_11324,N_10710);
nand U12203 (N_12203,N_11581,N_11589);
or U12204 (N_12204,N_11691,N_11354);
or U12205 (N_12205,N_11189,N_11758);
xor U12206 (N_12206,N_10688,N_11575);
nand U12207 (N_12207,N_11188,N_11858);
and U12208 (N_12208,N_10924,N_11970);
or U12209 (N_12209,N_11648,N_11027);
and U12210 (N_12210,N_11292,N_11394);
or U12211 (N_12211,N_10778,N_11549);
xnor U12212 (N_12212,N_10505,N_11947);
and U12213 (N_12213,N_11609,N_10959);
nor U12214 (N_12214,N_10744,N_11056);
and U12215 (N_12215,N_11767,N_11191);
and U12216 (N_12216,N_10646,N_10996);
nor U12217 (N_12217,N_10893,N_10628);
xnor U12218 (N_12218,N_11268,N_11611);
xnor U12219 (N_12219,N_11310,N_11817);
nand U12220 (N_12220,N_11020,N_11616);
or U12221 (N_12221,N_10875,N_11230);
nand U12222 (N_12222,N_11112,N_11569);
nand U12223 (N_12223,N_10670,N_11416);
nand U12224 (N_12224,N_10666,N_11486);
nor U12225 (N_12225,N_11047,N_11538);
nor U12226 (N_12226,N_10835,N_11231);
xor U12227 (N_12227,N_10615,N_11693);
nand U12228 (N_12228,N_10819,N_11500);
and U12229 (N_12229,N_11119,N_10802);
or U12230 (N_12230,N_10895,N_11826);
or U12231 (N_12231,N_11247,N_10564);
nor U12232 (N_12232,N_11750,N_11479);
nand U12233 (N_12233,N_11120,N_10852);
or U12234 (N_12234,N_10552,N_11017);
nor U12235 (N_12235,N_11495,N_11945);
and U12236 (N_12236,N_10827,N_11510);
and U12237 (N_12237,N_11794,N_10591);
or U12238 (N_12238,N_10611,N_10931);
and U12239 (N_12239,N_11160,N_10607);
or U12240 (N_12240,N_11291,N_11833);
and U12241 (N_12241,N_11069,N_10975);
and U12242 (N_12242,N_11514,N_11385);
and U12243 (N_12243,N_11219,N_11037);
nor U12244 (N_12244,N_11621,N_11801);
or U12245 (N_12245,N_11906,N_11316);
nand U12246 (N_12246,N_11208,N_10989);
and U12247 (N_12247,N_10728,N_10902);
nor U12248 (N_12248,N_11182,N_10560);
or U12249 (N_12249,N_11388,N_11270);
nand U12250 (N_12250,N_11458,N_10885);
or U12251 (N_12251,N_11695,N_10672);
xnor U12252 (N_12252,N_11210,N_11624);
xor U12253 (N_12253,N_10513,N_11157);
or U12254 (N_12254,N_10603,N_11612);
nor U12255 (N_12255,N_11493,N_11004);
xor U12256 (N_12256,N_11070,N_11907);
nand U12257 (N_12257,N_11809,N_11778);
nand U12258 (N_12258,N_10970,N_11356);
nand U12259 (N_12259,N_11274,N_11029);
xor U12260 (N_12260,N_11380,N_11248);
nor U12261 (N_12261,N_10814,N_11825);
xnor U12262 (N_12262,N_11232,N_10576);
or U12263 (N_12263,N_11735,N_11199);
or U12264 (N_12264,N_11810,N_11684);
and U12265 (N_12265,N_10600,N_11224);
nand U12266 (N_12266,N_11298,N_11963);
nand U12267 (N_12267,N_10711,N_11602);
or U12268 (N_12268,N_11606,N_10985);
and U12269 (N_12269,N_10551,N_11725);
nand U12270 (N_12270,N_10693,N_11573);
nor U12271 (N_12271,N_11859,N_11060);
and U12272 (N_12272,N_11028,N_11164);
or U12273 (N_12273,N_11150,N_11881);
and U12274 (N_12274,N_11578,N_11803);
xnor U12275 (N_12275,N_10647,N_11873);
xnor U12276 (N_12276,N_10855,N_11346);
nor U12277 (N_12277,N_11851,N_11467);
nand U12278 (N_12278,N_10700,N_11652);
and U12279 (N_12279,N_10509,N_11251);
xor U12280 (N_12280,N_10932,N_11646);
or U12281 (N_12281,N_11422,N_11245);
and U12282 (N_12282,N_11237,N_11759);
nand U12283 (N_12283,N_10971,N_10864);
and U12284 (N_12284,N_10503,N_10767);
xnor U12285 (N_12285,N_10896,N_11969);
xnor U12286 (N_12286,N_11456,N_11397);
or U12287 (N_12287,N_11683,N_10674);
nor U12288 (N_12288,N_10554,N_11361);
or U12289 (N_12289,N_11058,N_10815);
and U12290 (N_12290,N_10809,N_10746);
or U12291 (N_12291,N_11136,N_11995);
xnor U12292 (N_12292,N_10689,N_11939);
and U12293 (N_12293,N_11473,N_10725);
nand U12294 (N_12294,N_10708,N_11745);
and U12295 (N_12295,N_11240,N_11640);
nand U12296 (N_12296,N_10905,N_11642);
and U12297 (N_12297,N_11770,N_10772);
or U12298 (N_12298,N_11688,N_11311);
nor U12299 (N_12299,N_11496,N_11355);
or U12300 (N_12300,N_11663,N_11480);
or U12301 (N_12301,N_10581,N_11910);
nor U12302 (N_12302,N_11876,N_11152);
nand U12303 (N_12303,N_10919,N_11359);
nand U12304 (N_12304,N_11174,N_11411);
or U12305 (N_12305,N_11580,N_10696);
and U12306 (N_12306,N_11527,N_11490);
or U12307 (N_12307,N_11751,N_11552);
and U12308 (N_12308,N_11250,N_11315);
nor U12309 (N_12309,N_11800,N_11360);
xor U12310 (N_12310,N_11576,N_11358);
nor U12311 (N_12311,N_11747,N_10597);
nand U12312 (N_12312,N_11451,N_11035);
nand U12313 (N_12313,N_11222,N_11073);
xor U12314 (N_12314,N_11734,N_11146);
and U12315 (N_12315,N_11246,N_11185);
and U12316 (N_12316,N_10923,N_11290);
xor U12317 (N_12317,N_11960,N_11124);
and U12318 (N_12318,N_10640,N_11197);
or U12319 (N_12319,N_11905,N_10526);
nand U12320 (N_12320,N_11716,N_11926);
nor U12321 (N_12321,N_10854,N_11804);
or U12322 (N_12322,N_10847,N_10660);
or U12323 (N_12323,N_10517,N_11526);
or U12324 (N_12324,N_10669,N_11349);
nor U12325 (N_12325,N_11986,N_10928);
or U12326 (N_12326,N_10882,N_10818);
xnor U12327 (N_12327,N_10997,N_10570);
xor U12328 (N_12328,N_11568,N_11957);
nand U12329 (N_12329,N_11849,N_11223);
nand U12330 (N_12330,N_11707,N_10624);
or U12331 (N_12331,N_10578,N_11460);
or U12332 (N_12332,N_11104,N_11001);
xor U12333 (N_12333,N_11936,N_11052);
xnor U12334 (N_12334,N_10507,N_11636);
and U12335 (N_12335,N_11737,N_10656);
nor U12336 (N_12336,N_11305,N_10881);
or U12337 (N_12337,N_10687,N_10759);
or U12338 (N_12338,N_10745,N_10891);
or U12339 (N_12339,N_11114,N_11978);
xnor U12340 (N_12340,N_11741,N_11089);
or U12341 (N_12341,N_10704,N_10829);
or U12342 (N_12342,N_11314,N_11273);
nor U12343 (N_12343,N_11730,N_11530);
xor U12344 (N_12344,N_11518,N_10590);
nand U12345 (N_12345,N_10592,N_10884);
nand U12346 (N_12346,N_11329,N_10730);
nor U12347 (N_12347,N_11650,N_10565);
or U12348 (N_12348,N_11698,N_11874);
or U12349 (N_12349,N_11838,N_11353);
and U12350 (N_12350,N_11766,N_11561);
and U12351 (N_12351,N_11861,N_10506);
xor U12352 (N_12352,N_11238,N_10968);
and U12353 (N_12353,N_11265,N_10794);
nor U12354 (N_12354,N_10638,N_11487);
xor U12355 (N_12355,N_11045,N_11749);
nand U12356 (N_12356,N_11832,N_10619);
nand U12357 (N_12357,N_10798,N_11632);
and U12358 (N_12358,N_11599,N_10796);
nand U12359 (N_12359,N_10860,N_11788);
xor U12360 (N_12360,N_11228,N_11440);
and U12361 (N_12361,N_10841,N_10723);
xnor U12362 (N_12362,N_11154,N_10890);
nand U12363 (N_12363,N_10953,N_10609);
or U12364 (N_12364,N_11313,N_10768);
nand U12365 (N_12365,N_11180,N_10580);
or U12366 (N_12366,N_11704,N_10962);
or U12367 (N_12367,N_10987,N_11450);
nor U12368 (N_12368,N_11327,N_10695);
and U12369 (N_12369,N_11477,N_11532);
nor U12370 (N_12370,N_11824,N_11543);
or U12371 (N_12371,N_11701,N_11086);
nor U12372 (N_12372,N_10714,N_11337);
or U12373 (N_12373,N_11799,N_11622);
nor U12374 (N_12374,N_10518,N_11036);
or U12375 (N_12375,N_11438,N_10692);
or U12376 (N_12376,N_11000,N_11333);
nand U12377 (N_12377,N_11091,N_10762);
nand U12378 (N_12378,N_10956,N_11654);
nor U12379 (N_12379,N_11145,N_10753);
and U12380 (N_12380,N_10912,N_11147);
nand U12381 (N_12381,N_10889,N_11673);
and U12382 (N_12382,N_10735,N_11537);
xnor U12383 (N_12383,N_10779,N_10907);
nand U12384 (N_12384,N_11194,N_10584);
or U12385 (N_12385,N_10527,N_11293);
nor U12386 (N_12386,N_11868,N_11261);
xnor U12387 (N_12387,N_10828,N_11466);
or U12388 (N_12388,N_11856,N_10715);
xor U12389 (N_12389,N_11419,N_10716);
and U12390 (N_12390,N_11348,N_10694);
xnor U12391 (N_12391,N_11285,N_10553);
or U12392 (N_12392,N_11917,N_11229);
and U12393 (N_12393,N_10675,N_11334);
or U12394 (N_12394,N_10832,N_11196);
nand U12395 (N_12395,N_11634,N_11221);
xor U12396 (N_12396,N_11013,N_11709);
or U12397 (N_12397,N_11746,N_10900);
nand U12398 (N_12398,N_11719,N_10804);
nor U12399 (N_12399,N_11338,N_11702);
nor U12400 (N_12400,N_10620,N_11301);
nor U12401 (N_12401,N_11262,N_11300);
and U12402 (N_12402,N_11375,N_11277);
xor U12403 (N_12403,N_10622,N_11511);
xnor U12404 (N_12404,N_11175,N_10515);
or U12405 (N_12405,N_10982,N_11083);
nor U12406 (N_12406,N_11512,N_11708);
nand U12407 (N_12407,N_11630,N_11139);
and U12408 (N_12408,N_11598,N_11026);
nand U12409 (N_12409,N_11525,N_11078);
nand U12410 (N_12410,N_10776,N_10795);
or U12411 (N_12411,N_10904,N_10906);
xnor U12412 (N_12412,N_11762,N_10568);
and U12413 (N_12413,N_11434,N_11835);
nor U12414 (N_12414,N_11551,N_11006);
and U12415 (N_12415,N_10612,N_10760);
and U12416 (N_12416,N_11135,N_11200);
xor U12417 (N_12417,N_11792,N_11823);
nand U12418 (N_12418,N_10859,N_11031);
and U12419 (N_12419,N_11455,N_11100);
nand U12420 (N_12420,N_11276,N_11443);
xor U12421 (N_12421,N_11259,N_11209);
nor U12422 (N_12422,N_11149,N_10510);
and U12423 (N_12423,N_10599,N_10899);
or U12424 (N_12424,N_11299,N_11366);
nand U12425 (N_12425,N_11866,N_11672);
xor U12426 (N_12426,N_11966,N_11092);
xor U12427 (N_12427,N_11249,N_11930);
nand U12428 (N_12428,N_10781,N_11727);
or U12429 (N_12429,N_11773,N_10800);
and U12430 (N_12430,N_11133,N_11822);
or U12431 (N_12431,N_11030,N_11761);
xnor U12432 (N_12432,N_11623,N_11974);
or U12433 (N_12433,N_11167,N_11244);
or U12434 (N_12434,N_11205,N_11166);
or U12435 (N_12435,N_11795,N_10582);
nor U12436 (N_12436,N_10538,N_11269);
and U12437 (N_12437,N_11918,N_11021);
nor U12438 (N_12438,N_11217,N_11097);
nand U12439 (N_12439,N_11048,N_11015);
nor U12440 (N_12440,N_11002,N_10598);
nor U12441 (N_12441,N_11432,N_11882);
or U12442 (N_12442,N_11429,N_11522);
and U12443 (N_12443,N_11402,N_11400);
xor U12444 (N_12444,N_11852,N_11848);
nand U12445 (N_12445,N_11678,N_11644);
and U12446 (N_12446,N_11011,N_11942);
xor U12447 (N_12447,N_11880,N_10650);
nor U12448 (N_12448,N_10702,N_11481);
xnor U12449 (N_12449,N_10678,N_10791);
xor U12450 (N_12450,N_11075,N_11342);
nor U12451 (N_12451,N_11956,N_11018);
or U12452 (N_12452,N_10536,N_10869);
nor U12453 (N_12453,N_10894,N_11445);
nand U12454 (N_12454,N_11888,N_11853);
or U12455 (N_12455,N_10636,N_11720);
nor U12456 (N_12456,N_11607,N_11959);
or U12457 (N_12457,N_11263,N_11887);
nor U12458 (N_12458,N_11541,N_11732);
and U12459 (N_12459,N_10533,N_10874);
nor U12460 (N_12460,N_10837,N_10539);
xnor U12461 (N_12461,N_10901,N_11008);
nor U12462 (N_12462,N_11415,N_11108);
or U12463 (N_12463,N_10976,N_10935);
nor U12464 (N_12464,N_10583,N_11506);
nand U12465 (N_12465,N_10878,N_11520);
or U12466 (N_12466,N_10712,N_11908);
nand U12467 (N_12467,N_10626,N_11555);
and U12468 (N_12468,N_11631,N_10782);
nand U12469 (N_12469,N_11105,N_11294);
nor U12470 (N_12470,N_11666,N_10632);
xnor U12471 (N_12471,N_11516,N_10504);
nand U12472 (N_12472,N_11367,N_10535);
or U12473 (N_12473,N_11585,N_11577);
xnor U12474 (N_12474,N_11829,N_11148);
nor U12475 (N_12475,N_10732,N_10816);
xnor U12476 (N_12476,N_10917,N_10934);
xor U12477 (N_12477,N_11784,N_11176);
nand U12478 (N_12478,N_11158,N_10817);
and U12479 (N_12479,N_10978,N_11275);
or U12480 (N_12480,N_10787,N_11593);
and U12481 (N_12481,N_11857,N_10743);
xnor U12482 (N_12482,N_11655,N_11492);
nand U12483 (N_12483,N_10601,N_10955);
and U12484 (N_12484,N_10806,N_10960);
nand U12485 (N_12485,N_11893,N_10541);
and U12486 (N_12486,N_10697,N_11840);
xor U12487 (N_12487,N_11862,N_11647);
nand U12488 (N_12488,N_11777,N_10522);
nand U12489 (N_12489,N_11554,N_11566);
nand U12490 (N_12490,N_10964,N_10707);
nand U12491 (N_12491,N_11079,N_10937);
or U12492 (N_12492,N_11608,N_11382);
nand U12493 (N_12493,N_11098,N_10946);
or U12494 (N_12494,N_11038,N_10929);
and U12495 (N_12495,N_10500,N_11865);
xnor U12496 (N_12496,N_10737,N_11932);
nand U12497 (N_12497,N_11870,N_11662);
and U12498 (N_12498,N_11141,N_11453);
xnor U12499 (N_12499,N_11243,N_10943);
nand U12500 (N_12500,N_11793,N_10530);
or U12501 (N_12501,N_11427,N_11132);
xor U12502 (N_12502,N_11161,N_11433);
or U12503 (N_12503,N_10988,N_11312);
or U12504 (N_12504,N_10972,N_11323);
and U12505 (N_12505,N_11600,N_11449);
or U12506 (N_12506,N_10843,N_11821);
nor U12507 (N_12507,N_11472,N_11335);
nor U12508 (N_12508,N_11879,N_11253);
or U12509 (N_12509,N_10858,N_10655);
nand U12510 (N_12510,N_11387,N_11213);
nand U12511 (N_12511,N_11962,N_10754);
nand U12512 (N_12512,N_11993,N_10933);
or U12513 (N_12513,N_11989,N_11842);
nand U12514 (N_12514,N_11928,N_11922);
nor U12515 (N_12515,N_11948,N_11331);
nor U12516 (N_12516,N_11431,N_11592);
xor U12517 (N_12517,N_10748,N_11465);
xnor U12518 (N_12518,N_11878,N_11921);
nand U12519 (N_12519,N_11446,N_10764);
or U12520 (N_12520,N_10898,N_11604);
xnor U12521 (N_12521,N_10731,N_10916);
or U12522 (N_12522,N_11933,N_10998);
nor U12523 (N_12523,N_10949,N_11297);
nor U12524 (N_12524,N_11032,N_11871);
nor U12525 (N_12525,N_11170,N_11127);
nand U12526 (N_12526,N_11118,N_11528);
or U12527 (N_12527,N_11517,N_11764);
nand U12528 (N_12528,N_11756,N_11489);
and U12529 (N_12529,N_10665,N_11376);
and U12530 (N_12530,N_11390,N_11548);
nor U12531 (N_12531,N_11864,N_10698);
or U12532 (N_12532,N_11207,N_11740);
nor U12533 (N_12533,N_11771,N_11236);
or U12534 (N_12534,N_10586,N_10722);
and U12535 (N_12535,N_11409,N_11628);
nand U12536 (N_12536,N_11328,N_10738);
nor U12537 (N_12537,N_11711,N_11106);
nand U12538 (N_12538,N_11093,N_11557);
and U12539 (N_12539,N_11689,N_11796);
and U12540 (N_12540,N_11463,N_10631);
nor U12541 (N_12541,N_10516,N_11590);
xor U12542 (N_12542,N_11436,N_11381);
or U12543 (N_12543,N_10648,N_11911);
nand U12544 (N_12544,N_11884,N_11485);
nand U12545 (N_12545,N_10546,N_11679);
or U12546 (N_12546,N_11107,N_11949);
xor U12547 (N_12547,N_10685,N_11912);
nor U12548 (N_12548,N_11287,N_10645);
xnor U12549 (N_12549,N_10833,N_11736);
nor U12550 (N_12550,N_11892,N_10561);
or U12551 (N_12551,N_11961,N_11085);
xnor U12552 (N_12552,N_11597,N_11442);
nand U12553 (N_12553,N_11352,N_11171);
or U12554 (N_12554,N_10873,N_10606);
and U12555 (N_12555,N_11126,N_10826);
xor U12556 (N_12556,N_11267,N_11284);
nor U12557 (N_12557,N_10903,N_11763);
xor U12558 (N_12558,N_11116,N_10525);
and U12559 (N_12559,N_11534,N_11077);
or U12560 (N_12560,N_11288,N_10865);
nor U12561 (N_12561,N_11717,N_11258);
and U12562 (N_12562,N_11798,N_11435);
or U12563 (N_12563,N_11964,N_11583);
and U12564 (N_12564,N_11785,N_11055);
nand U12565 (N_12565,N_11140,N_10751);
or U12566 (N_12566,N_11617,N_10643);
nor U12567 (N_12567,N_11296,N_11101);
nand U12568 (N_12568,N_11980,N_11542);
and U12569 (N_12569,N_10740,N_11676);
nor U12570 (N_12570,N_11724,N_11373);
nand U12571 (N_12571,N_10567,N_11588);
nor U12572 (N_12572,N_11041,N_10596);
xnor U12573 (N_12573,N_11418,N_11206);
and U12574 (N_12574,N_10691,N_11513);
or U12575 (N_12575,N_11317,N_10877);
or U12576 (N_12576,N_10756,N_11144);
xor U12577 (N_12577,N_11536,N_11523);
nor U12578 (N_12578,N_11883,N_11789);
and U12579 (N_12579,N_11505,N_10579);
nand U12580 (N_12580,N_11550,N_11981);
and U12581 (N_12581,N_11255,N_11619);
nand U12582 (N_12582,N_11063,N_10918);
nor U12583 (N_12583,N_11562,N_11023);
nor U12584 (N_12584,N_11066,N_11022);
nor U12585 (N_12585,N_11110,N_11627);
xor U12586 (N_12586,N_10805,N_10594);
or U12587 (N_12587,N_11603,N_10825);
nor U12588 (N_12588,N_10528,N_10658);
xor U12589 (N_12589,N_10610,N_10569);
nand U12590 (N_12590,N_10720,N_10936);
or U12591 (N_12591,N_11775,N_11256);
xor U12592 (N_12592,N_10595,N_11529);
or U12593 (N_12593,N_11457,N_10699);
nand U12594 (N_12594,N_10831,N_11395);
nand U12595 (N_12595,N_10926,N_11350);
and U12596 (N_12596,N_10679,N_10547);
and U12597 (N_12597,N_10783,N_11046);
nor U12598 (N_12598,N_10951,N_11319);
or U12599 (N_12599,N_10824,N_11744);
and U12600 (N_12600,N_11813,N_11653);
and U12601 (N_12601,N_10532,N_11499);
xnor U12602 (N_12602,N_10792,N_10573);
nand U12603 (N_12603,N_10979,N_11090);
and U12604 (N_12604,N_10995,N_11899);
xor U12605 (N_12605,N_10870,N_10867);
nor U12606 (N_12606,N_10742,N_11344);
xor U12607 (N_12607,N_11183,N_11109);
and U12608 (N_12608,N_10788,N_11153);
nor U12609 (N_12609,N_10604,N_11051);
xnor U12610 (N_12610,N_11370,N_11009);
or U12611 (N_12611,N_11169,N_11076);
and U12612 (N_12612,N_11420,N_10653);
and U12613 (N_12613,N_10892,N_11805);
xnor U12614 (N_12614,N_11668,N_11694);
and U12615 (N_12615,N_10810,N_11498);
or U12616 (N_12616,N_10786,N_11103);
or U12617 (N_12617,N_10549,N_11584);
nor U12618 (N_12618,N_11914,N_11998);
or U12619 (N_12619,N_10807,N_10872);
nand U12620 (N_12620,N_10856,N_11398);
or U12621 (N_12621,N_11996,N_10908);
nand U12622 (N_12622,N_11816,N_11203);
nand U12623 (N_12623,N_11034,N_11643);
xnor U12624 (N_12624,N_10984,N_11102);
and U12625 (N_12625,N_11768,N_10973);
or U12626 (N_12626,N_10844,N_11927);
xor U12627 (N_12627,N_10508,N_11121);
nand U12628 (N_12628,N_11111,N_11563);
or U12629 (N_12629,N_10994,N_10801);
nor U12630 (N_12630,N_10727,N_11574);
nor U12631 (N_12631,N_11507,N_11743);
nand U12632 (N_12632,N_11264,N_11976);
or U12633 (N_12633,N_11095,N_11991);
nor U12634 (N_12634,N_10977,N_11705);
nor U12635 (N_12635,N_11474,N_10623);
and U12636 (N_12636,N_11660,N_11738);
and U12637 (N_12637,N_11198,N_11437);
xnor U12638 (N_12638,N_10661,N_11731);
nor U12639 (N_12639,N_10986,N_11710);
nor U12640 (N_12640,N_11184,N_10862);
and U12641 (N_12641,N_11765,N_11808);
xor U12642 (N_12642,N_11831,N_11295);
xor U12643 (N_12643,N_11594,N_11714);
or U12644 (N_12644,N_11651,N_10780);
and U12645 (N_12645,N_11895,N_11042);
nand U12646 (N_12646,N_11257,N_11687);
and U12647 (N_12647,N_11987,N_11272);
nor U12648 (N_12648,N_10999,N_11772);
nor U12649 (N_12649,N_11985,N_10701);
or U12650 (N_12650,N_10649,N_11065);
and U12651 (N_12651,N_11625,N_10927);
xor U12652 (N_12652,N_10627,N_11464);
and U12653 (N_12653,N_11155,N_10684);
xnor U12654 (N_12654,N_11115,N_10733);
or U12655 (N_12655,N_10630,N_11753);
and U12656 (N_12656,N_10965,N_11214);
and U12657 (N_12657,N_10822,N_11776);
or U12658 (N_12658,N_11977,N_11254);
xor U12659 (N_12659,N_11699,N_11365);
xor U12660 (N_12660,N_10868,N_11885);
nor U12661 (N_12661,N_11913,N_11941);
and U12662 (N_12662,N_11384,N_11965);
nor U12663 (N_12663,N_10635,N_11728);
xnor U12664 (N_12664,N_11072,N_11586);
nor U12665 (N_12665,N_11165,N_10839);
nor U12666 (N_12666,N_10838,N_11509);
nand U12667 (N_12667,N_10703,N_10563);
xor U12668 (N_12668,N_10639,N_10887);
nor U12669 (N_12669,N_11405,N_11779);
nor U12670 (N_12670,N_10761,N_11088);
nor U12671 (N_12671,N_11610,N_11519);
and U12672 (N_12672,N_10520,N_11407);
xnor U12673 (N_12673,N_11567,N_10992);
nand U12674 (N_12674,N_10897,N_10883);
nor U12675 (N_12675,N_11515,N_11940);
nand U12676 (N_12676,N_11129,N_10925);
nor U12677 (N_12677,N_11700,N_11682);
or U12678 (N_12678,N_11181,N_10652);
nand U12679 (N_12679,N_11844,N_10821);
and U12680 (N_12680,N_11524,N_11596);
xor U12681 (N_12681,N_11919,N_11955);
xnor U12682 (N_12682,N_11830,N_11979);
or U12683 (N_12683,N_10543,N_11502);
nor U12684 (N_12684,N_11123,N_11755);
nand U12685 (N_12685,N_11994,N_10967);
or U12686 (N_12686,N_11897,N_11685);
or U12687 (N_12687,N_10846,N_11629);
nor U12688 (N_12688,N_11271,N_11967);
nor U12689 (N_12689,N_11138,N_11860);
xor U12690 (N_12690,N_10542,N_10614);
nand U12691 (N_12691,N_11587,N_11378);
or U12692 (N_12692,N_10593,N_10587);
and U12693 (N_12693,N_11504,N_11900);
and U12694 (N_12694,N_10981,N_10657);
or U12695 (N_12695,N_11943,N_10625);
and U12696 (N_12696,N_11571,N_11863);
nand U12697 (N_12697,N_11791,N_11151);
nand U12698 (N_12698,N_11483,N_10914);
xor U12699 (N_12699,N_11742,N_11620);
and U12700 (N_12700,N_11341,N_10557);
nor U12701 (N_12701,N_11082,N_11706);
nand U12702 (N_12702,N_11649,N_11712);
xnor U12703 (N_12703,N_11613,N_10676);
and U12704 (N_12704,N_10857,N_11729);
and U12705 (N_12705,N_11723,N_10550);
nand U12706 (N_12706,N_11540,N_11818);
nor U12707 (N_12707,N_10812,N_10980);
or U12708 (N_12708,N_10556,N_11372);
nor U12709 (N_12709,N_11656,N_11233);
or U12710 (N_12710,N_11172,N_11260);
xnor U12711 (N_12711,N_10690,N_10663);
nand U12712 (N_12712,N_11847,N_11638);
xnor U12713 (N_12713,N_10736,N_11539);
and U12714 (N_12714,N_11626,N_10616);
xnor U12715 (N_12715,N_11971,N_10605);
and U12716 (N_12716,N_11670,N_11401);
and U12717 (N_12717,N_10621,N_11043);
xor U12718 (N_12718,N_11664,N_10741);
xor U12719 (N_12719,N_11988,N_10717);
nor U12720 (N_12720,N_10915,N_11113);
or U12721 (N_12721,N_11343,N_11999);
xnor U12722 (N_12722,N_11488,N_11674);
or U12723 (N_12723,N_10775,N_11280);
nor U12724 (N_12724,N_11159,N_11475);
xnor U12725 (N_12725,N_11820,N_10823);
xor U12726 (N_12726,N_11559,N_10681);
or U12727 (N_12727,N_11595,N_11374);
xor U12728 (N_12728,N_10757,N_11733);
nand U12729 (N_12729,N_10930,N_11304);
xor U12730 (N_12730,N_11944,N_10613);
nor U12731 (N_12731,N_11992,N_11351);
xnor U12732 (N_12732,N_11854,N_11635);
nor U12733 (N_12733,N_10577,N_11904);
nor U12734 (N_12734,N_11391,N_11019);
nand U12735 (N_12735,N_11278,N_11468);
and U12736 (N_12736,N_10765,N_11242);
nor U12737 (N_12737,N_11215,N_10667);
or U12738 (N_12738,N_11605,N_10644);
nand U12739 (N_12739,N_10588,N_11819);
and U12740 (N_12740,N_10654,N_11064);
or U12741 (N_12741,N_10790,N_11218);
or U12742 (N_12742,N_10849,N_10558);
xor U12743 (N_12743,N_11760,N_10770);
or U12744 (N_12744,N_11403,N_11393);
and U12745 (N_12745,N_11946,N_11503);
or U12746 (N_12746,N_10671,N_11657);
or U12747 (N_12747,N_11469,N_11377);
xnor U12748 (N_12748,N_10519,N_11570);
nor U12749 (N_12749,N_11428,N_11462);
xor U12750 (N_12750,N_10995,N_11838);
nand U12751 (N_12751,N_11389,N_10869);
nand U12752 (N_12752,N_10853,N_11079);
and U12753 (N_12753,N_10946,N_11664);
nor U12754 (N_12754,N_10843,N_11410);
nand U12755 (N_12755,N_10743,N_11005);
and U12756 (N_12756,N_10797,N_11325);
and U12757 (N_12757,N_11747,N_11380);
and U12758 (N_12758,N_11538,N_11108);
xnor U12759 (N_12759,N_10593,N_11440);
xnor U12760 (N_12760,N_11666,N_11515);
xor U12761 (N_12761,N_10961,N_11117);
xnor U12762 (N_12762,N_10918,N_11664);
or U12763 (N_12763,N_10702,N_11725);
nor U12764 (N_12764,N_10738,N_11498);
nor U12765 (N_12765,N_11786,N_11664);
nand U12766 (N_12766,N_11877,N_11312);
nand U12767 (N_12767,N_11601,N_11192);
or U12768 (N_12768,N_10973,N_10785);
or U12769 (N_12769,N_11071,N_11525);
nand U12770 (N_12770,N_10636,N_11248);
xnor U12771 (N_12771,N_11230,N_10965);
and U12772 (N_12772,N_11730,N_11414);
nand U12773 (N_12773,N_10751,N_11271);
and U12774 (N_12774,N_11598,N_11123);
or U12775 (N_12775,N_11565,N_11259);
and U12776 (N_12776,N_11199,N_10814);
or U12777 (N_12777,N_10983,N_10514);
nand U12778 (N_12778,N_11446,N_10567);
and U12779 (N_12779,N_10995,N_11255);
nor U12780 (N_12780,N_11346,N_11856);
and U12781 (N_12781,N_11283,N_10677);
nor U12782 (N_12782,N_10659,N_11182);
and U12783 (N_12783,N_11736,N_10973);
and U12784 (N_12784,N_10932,N_11268);
nor U12785 (N_12785,N_11195,N_10761);
nand U12786 (N_12786,N_11127,N_10622);
xor U12787 (N_12787,N_10705,N_11981);
nor U12788 (N_12788,N_11923,N_11390);
or U12789 (N_12789,N_10717,N_11595);
and U12790 (N_12790,N_10523,N_11776);
or U12791 (N_12791,N_10958,N_11769);
and U12792 (N_12792,N_11322,N_11353);
nor U12793 (N_12793,N_11522,N_11495);
or U12794 (N_12794,N_11600,N_11410);
nor U12795 (N_12795,N_11140,N_10603);
xnor U12796 (N_12796,N_11059,N_11935);
or U12797 (N_12797,N_11747,N_10957);
nand U12798 (N_12798,N_11912,N_11780);
nand U12799 (N_12799,N_10669,N_11670);
xnor U12800 (N_12800,N_11922,N_10946);
nor U12801 (N_12801,N_10573,N_11829);
xor U12802 (N_12802,N_11172,N_11702);
nor U12803 (N_12803,N_11129,N_11890);
or U12804 (N_12804,N_10980,N_11410);
nor U12805 (N_12805,N_11052,N_11735);
and U12806 (N_12806,N_10915,N_11277);
nand U12807 (N_12807,N_11493,N_11150);
or U12808 (N_12808,N_10619,N_11333);
xnor U12809 (N_12809,N_10884,N_11802);
nor U12810 (N_12810,N_11326,N_11543);
or U12811 (N_12811,N_11994,N_10936);
xor U12812 (N_12812,N_11234,N_11763);
xor U12813 (N_12813,N_11585,N_10573);
nor U12814 (N_12814,N_10639,N_11173);
nor U12815 (N_12815,N_10545,N_11555);
and U12816 (N_12816,N_11928,N_11542);
or U12817 (N_12817,N_11169,N_11103);
xor U12818 (N_12818,N_11072,N_11714);
nor U12819 (N_12819,N_11399,N_10654);
nor U12820 (N_12820,N_11399,N_10676);
and U12821 (N_12821,N_11270,N_11557);
or U12822 (N_12822,N_11903,N_11662);
or U12823 (N_12823,N_11923,N_11321);
nand U12824 (N_12824,N_10681,N_11913);
xor U12825 (N_12825,N_11839,N_11597);
xnor U12826 (N_12826,N_11055,N_11975);
and U12827 (N_12827,N_11620,N_11837);
nor U12828 (N_12828,N_11122,N_10844);
and U12829 (N_12829,N_10712,N_11624);
or U12830 (N_12830,N_10908,N_10587);
nor U12831 (N_12831,N_11860,N_11204);
nor U12832 (N_12832,N_10649,N_10893);
xnor U12833 (N_12833,N_11382,N_11658);
xnor U12834 (N_12834,N_11308,N_11270);
or U12835 (N_12835,N_11297,N_10734);
or U12836 (N_12836,N_11543,N_11587);
or U12837 (N_12837,N_10555,N_10745);
and U12838 (N_12838,N_11857,N_10633);
nor U12839 (N_12839,N_11092,N_11699);
or U12840 (N_12840,N_11095,N_11949);
and U12841 (N_12841,N_10680,N_11208);
xnor U12842 (N_12842,N_10830,N_11368);
nor U12843 (N_12843,N_10615,N_11468);
or U12844 (N_12844,N_11890,N_10830);
or U12845 (N_12845,N_11998,N_10622);
nand U12846 (N_12846,N_11319,N_10737);
nor U12847 (N_12847,N_11990,N_11176);
xor U12848 (N_12848,N_11156,N_10581);
and U12849 (N_12849,N_11110,N_11834);
and U12850 (N_12850,N_10794,N_10788);
or U12851 (N_12851,N_10957,N_11876);
nand U12852 (N_12852,N_11679,N_11254);
or U12853 (N_12853,N_11423,N_11477);
xor U12854 (N_12854,N_11711,N_11685);
xor U12855 (N_12855,N_11059,N_11513);
nand U12856 (N_12856,N_11545,N_10914);
and U12857 (N_12857,N_10839,N_11474);
and U12858 (N_12858,N_11568,N_10793);
xor U12859 (N_12859,N_11735,N_11885);
xnor U12860 (N_12860,N_11808,N_10807);
nand U12861 (N_12861,N_11080,N_10871);
xor U12862 (N_12862,N_10667,N_11790);
and U12863 (N_12863,N_10990,N_10528);
nand U12864 (N_12864,N_11002,N_11613);
xnor U12865 (N_12865,N_11002,N_11395);
xnor U12866 (N_12866,N_11721,N_11659);
xor U12867 (N_12867,N_11066,N_11616);
nor U12868 (N_12868,N_11075,N_11536);
or U12869 (N_12869,N_11802,N_10655);
or U12870 (N_12870,N_11757,N_11358);
and U12871 (N_12871,N_11568,N_10981);
and U12872 (N_12872,N_10532,N_10682);
or U12873 (N_12873,N_11771,N_11046);
or U12874 (N_12874,N_11007,N_10773);
nor U12875 (N_12875,N_11246,N_11702);
and U12876 (N_12876,N_11975,N_11430);
nor U12877 (N_12877,N_11196,N_11408);
nand U12878 (N_12878,N_11175,N_10895);
nand U12879 (N_12879,N_11331,N_10554);
nor U12880 (N_12880,N_11454,N_11448);
or U12881 (N_12881,N_11807,N_11982);
and U12882 (N_12882,N_11366,N_11356);
and U12883 (N_12883,N_11180,N_11273);
nor U12884 (N_12884,N_10935,N_11870);
nand U12885 (N_12885,N_11054,N_11403);
and U12886 (N_12886,N_11821,N_11018);
or U12887 (N_12887,N_10985,N_11696);
nor U12888 (N_12888,N_11767,N_11953);
xor U12889 (N_12889,N_10786,N_11454);
xor U12890 (N_12890,N_11155,N_11214);
and U12891 (N_12891,N_11578,N_11486);
and U12892 (N_12892,N_10525,N_10550);
and U12893 (N_12893,N_10957,N_10940);
or U12894 (N_12894,N_11491,N_11913);
and U12895 (N_12895,N_11988,N_11074);
nor U12896 (N_12896,N_10605,N_11975);
or U12897 (N_12897,N_11694,N_11154);
and U12898 (N_12898,N_11678,N_10810);
nor U12899 (N_12899,N_10649,N_11934);
nor U12900 (N_12900,N_11943,N_11366);
and U12901 (N_12901,N_11128,N_11369);
and U12902 (N_12902,N_11922,N_11051);
and U12903 (N_12903,N_11881,N_11139);
xnor U12904 (N_12904,N_11119,N_11647);
xor U12905 (N_12905,N_11624,N_11154);
and U12906 (N_12906,N_10652,N_11980);
nand U12907 (N_12907,N_10665,N_11475);
xor U12908 (N_12908,N_11583,N_11843);
xnor U12909 (N_12909,N_11573,N_11036);
or U12910 (N_12910,N_10945,N_10665);
nand U12911 (N_12911,N_10807,N_11608);
nand U12912 (N_12912,N_11334,N_10957);
nor U12913 (N_12913,N_11150,N_11280);
and U12914 (N_12914,N_11204,N_11700);
nand U12915 (N_12915,N_11450,N_11047);
or U12916 (N_12916,N_11930,N_10582);
and U12917 (N_12917,N_10715,N_11964);
and U12918 (N_12918,N_11341,N_11488);
xor U12919 (N_12919,N_11710,N_10977);
nor U12920 (N_12920,N_11786,N_10857);
nor U12921 (N_12921,N_11509,N_11397);
nand U12922 (N_12922,N_11116,N_11034);
xor U12923 (N_12923,N_10843,N_11168);
and U12924 (N_12924,N_10538,N_11125);
or U12925 (N_12925,N_10524,N_11198);
xor U12926 (N_12926,N_11390,N_11546);
nand U12927 (N_12927,N_11909,N_10911);
and U12928 (N_12928,N_11686,N_11655);
nor U12929 (N_12929,N_11650,N_11819);
or U12930 (N_12930,N_11148,N_11871);
xor U12931 (N_12931,N_10970,N_10872);
nor U12932 (N_12932,N_10900,N_11728);
nor U12933 (N_12933,N_10926,N_11337);
and U12934 (N_12934,N_11417,N_11862);
and U12935 (N_12935,N_10659,N_11636);
nand U12936 (N_12936,N_10759,N_11037);
xnor U12937 (N_12937,N_11490,N_11079);
xnor U12938 (N_12938,N_11752,N_11824);
or U12939 (N_12939,N_11745,N_11478);
nor U12940 (N_12940,N_11189,N_11696);
xor U12941 (N_12941,N_11042,N_11565);
and U12942 (N_12942,N_11142,N_10596);
nand U12943 (N_12943,N_10913,N_11939);
xnor U12944 (N_12944,N_10740,N_10638);
xnor U12945 (N_12945,N_11780,N_11430);
nor U12946 (N_12946,N_11075,N_11713);
nor U12947 (N_12947,N_10625,N_11161);
nand U12948 (N_12948,N_11290,N_10976);
or U12949 (N_12949,N_10514,N_10513);
or U12950 (N_12950,N_11213,N_10744);
nor U12951 (N_12951,N_11533,N_11820);
or U12952 (N_12952,N_11187,N_10910);
nand U12953 (N_12953,N_10541,N_11348);
xor U12954 (N_12954,N_10951,N_11220);
xnor U12955 (N_12955,N_11769,N_11650);
nand U12956 (N_12956,N_10598,N_11447);
xor U12957 (N_12957,N_11620,N_10769);
nor U12958 (N_12958,N_11300,N_11677);
nor U12959 (N_12959,N_11635,N_10677);
and U12960 (N_12960,N_11315,N_10631);
or U12961 (N_12961,N_11112,N_10840);
or U12962 (N_12962,N_10504,N_11279);
nand U12963 (N_12963,N_11625,N_11447);
and U12964 (N_12964,N_10694,N_11718);
and U12965 (N_12965,N_11344,N_11130);
and U12966 (N_12966,N_11368,N_10944);
nand U12967 (N_12967,N_11835,N_10674);
and U12968 (N_12968,N_11828,N_11244);
and U12969 (N_12969,N_11757,N_10688);
xor U12970 (N_12970,N_10857,N_11783);
xnor U12971 (N_12971,N_11575,N_11008);
nand U12972 (N_12972,N_11037,N_11196);
nor U12973 (N_12973,N_10807,N_10975);
and U12974 (N_12974,N_11278,N_11735);
and U12975 (N_12975,N_10772,N_11368);
nand U12976 (N_12976,N_10735,N_10775);
nor U12977 (N_12977,N_10862,N_11817);
xnor U12978 (N_12978,N_11367,N_10623);
xnor U12979 (N_12979,N_11367,N_11143);
xnor U12980 (N_12980,N_10660,N_11138);
or U12981 (N_12981,N_11414,N_11635);
or U12982 (N_12982,N_11580,N_10889);
xnor U12983 (N_12983,N_11335,N_11559);
nand U12984 (N_12984,N_10552,N_10679);
nor U12985 (N_12985,N_11092,N_11478);
nor U12986 (N_12986,N_11842,N_11715);
nor U12987 (N_12987,N_10852,N_11648);
nand U12988 (N_12988,N_11120,N_11564);
and U12989 (N_12989,N_10981,N_10950);
nand U12990 (N_12990,N_10725,N_11985);
xor U12991 (N_12991,N_11314,N_10510);
nand U12992 (N_12992,N_11686,N_11822);
xnor U12993 (N_12993,N_10741,N_11751);
or U12994 (N_12994,N_11007,N_11735);
nand U12995 (N_12995,N_11846,N_11038);
or U12996 (N_12996,N_11952,N_11639);
nand U12997 (N_12997,N_10618,N_11599);
nor U12998 (N_12998,N_10768,N_10521);
and U12999 (N_12999,N_11284,N_11159);
nand U13000 (N_13000,N_10513,N_11796);
nor U13001 (N_13001,N_11038,N_11218);
and U13002 (N_13002,N_11139,N_11738);
nor U13003 (N_13003,N_11529,N_11312);
nor U13004 (N_13004,N_11254,N_11696);
nand U13005 (N_13005,N_10732,N_10937);
nand U13006 (N_13006,N_11061,N_11738);
xnor U13007 (N_13007,N_10852,N_11373);
or U13008 (N_13008,N_10591,N_10797);
or U13009 (N_13009,N_10557,N_11486);
nand U13010 (N_13010,N_10559,N_10742);
and U13011 (N_13011,N_11062,N_11716);
or U13012 (N_13012,N_11732,N_11866);
xnor U13013 (N_13013,N_10554,N_11639);
and U13014 (N_13014,N_11447,N_11603);
nor U13015 (N_13015,N_11056,N_10791);
xnor U13016 (N_13016,N_11778,N_11740);
nand U13017 (N_13017,N_11155,N_11633);
nand U13018 (N_13018,N_11396,N_10658);
nand U13019 (N_13019,N_10889,N_11610);
xnor U13020 (N_13020,N_11633,N_11531);
nor U13021 (N_13021,N_11742,N_11694);
or U13022 (N_13022,N_10628,N_10682);
nor U13023 (N_13023,N_10887,N_10967);
or U13024 (N_13024,N_11233,N_11983);
nand U13025 (N_13025,N_11447,N_10564);
nand U13026 (N_13026,N_11052,N_11413);
nor U13027 (N_13027,N_11498,N_11858);
xnor U13028 (N_13028,N_11532,N_11415);
nand U13029 (N_13029,N_10540,N_11973);
xnor U13030 (N_13030,N_11537,N_10538);
xor U13031 (N_13031,N_10705,N_11309);
xnor U13032 (N_13032,N_11261,N_11134);
nand U13033 (N_13033,N_11441,N_10656);
or U13034 (N_13034,N_11155,N_11788);
xor U13035 (N_13035,N_11945,N_11591);
nand U13036 (N_13036,N_11954,N_11822);
nand U13037 (N_13037,N_11055,N_10622);
xor U13038 (N_13038,N_11170,N_11611);
or U13039 (N_13039,N_11506,N_10854);
xnor U13040 (N_13040,N_11439,N_11897);
and U13041 (N_13041,N_10789,N_11333);
nand U13042 (N_13042,N_11187,N_11120);
nand U13043 (N_13043,N_11558,N_10715);
nand U13044 (N_13044,N_11370,N_11286);
xnor U13045 (N_13045,N_11339,N_10991);
xor U13046 (N_13046,N_10968,N_11132);
nand U13047 (N_13047,N_11041,N_10573);
nand U13048 (N_13048,N_11937,N_11261);
or U13049 (N_13049,N_10958,N_11210);
or U13050 (N_13050,N_10546,N_10962);
xnor U13051 (N_13051,N_10803,N_10687);
xnor U13052 (N_13052,N_10897,N_11305);
and U13053 (N_13053,N_11853,N_11804);
nand U13054 (N_13054,N_11759,N_10564);
and U13055 (N_13055,N_11579,N_11549);
nand U13056 (N_13056,N_10870,N_10691);
nand U13057 (N_13057,N_10993,N_10557);
xor U13058 (N_13058,N_11748,N_10550);
nand U13059 (N_13059,N_11191,N_11641);
xnor U13060 (N_13060,N_11166,N_11830);
xnor U13061 (N_13061,N_11724,N_11067);
and U13062 (N_13062,N_11853,N_11491);
and U13063 (N_13063,N_10851,N_11792);
and U13064 (N_13064,N_11249,N_11564);
or U13065 (N_13065,N_11032,N_10731);
xor U13066 (N_13066,N_10699,N_11268);
or U13067 (N_13067,N_11385,N_10939);
or U13068 (N_13068,N_11298,N_10648);
nand U13069 (N_13069,N_11741,N_11950);
nand U13070 (N_13070,N_11199,N_10528);
nand U13071 (N_13071,N_11568,N_11032);
nor U13072 (N_13072,N_11918,N_11652);
and U13073 (N_13073,N_11281,N_11493);
nor U13074 (N_13074,N_11312,N_10816);
nand U13075 (N_13075,N_11141,N_11815);
xnor U13076 (N_13076,N_11392,N_11094);
or U13077 (N_13077,N_11422,N_11080);
and U13078 (N_13078,N_10891,N_11561);
nand U13079 (N_13079,N_11231,N_10818);
and U13080 (N_13080,N_11145,N_10739);
xor U13081 (N_13081,N_10735,N_10552);
xnor U13082 (N_13082,N_10865,N_10645);
xor U13083 (N_13083,N_10597,N_11710);
nor U13084 (N_13084,N_11442,N_10988);
nor U13085 (N_13085,N_10835,N_11749);
nor U13086 (N_13086,N_11067,N_11745);
nor U13087 (N_13087,N_11101,N_10700);
xor U13088 (N_13088,N_11579,N_11179);
or U13089 (N_13089,N_11021,N_10995);
nor U13090 (N_13090,N_11585,N_11374);
nor U13091 (N_13091,N_10572,N_11904);
xor U13092 (N_13092,N_10544,N_11768);
nand U13093 (N_13093,N_11520,N_10865);
xnor U13094 (N_13094,N_11803,N_10682);
nor U13095 (N_13095,N_11078,N_11752);
and U13096 (N_13096,N_11680,N_10747);
nand U13097 (N_13097,N_11754,N_11422);
and U13098 (N_13098,N_11206,N_11073);
nor U13099 (N_13099,N_10568,N_11804);
or U13100 (N_13100,N_10704,N_11597);
and U13101 (N_13101,N_11234,N_10715);
nor U13102 (N_13102,N_11350,N_10883);
and U13103 (N_13103,N_11122,N_11120);
and U13104 (N_13104,N_10650,N_10626);
nand U13105 (N_13105,N_11947,N_11093);
nor U13106 (N_13106,N_11212,N_11401);
nand U13107 (N_13107,N_11416,N_11691);
xor U13108 (N_13108,N_10573,N_10654);
or U13109 (N_13109,N_11757,N_11043);
nand U13110 (N_13110,N_11467,N_11339);
and U13111 (N_13111,N_11422,N_11472);
and U13112 (N_13112,N_11939,N_11416);
nor U13113 (N_13113,N_11823,N_11827);
or U13114 (N_13114,N_11987,N_11828);
and U13115 (N_13115,N_10699,N_10961);
nand U13116 (N_13116,N_11335,N_11441);
xor U13117 (N_13117,N_10523,N_11104);
xnor U13118 (N_13118,N_11266,N_11201);
and U13119 (N_13119,N_10968,N_10834);
and U13120 (N_13120,N_10998,N_11430);
and U13121 (N_13121,N_11617,N_10851);
nand U13122 (N_13122,N_10643,N_10839);
and U13123 (N_13123,N_11727,N_11649);
nand U13124 (N_13124,N_11590,N_11852);
nand U13125 (N_13125,N_11426,N_11079);
nor U13126 (N_13126,N_11739,N_10544);
nand U13127 (N_13127,N_11912,N_11240);
or U13128 (N_13128,N_11536,N_11487);
nand U13129 (N_13129,N_11912,N_10852);
nand U13130 (N_13130,N_11600,N_10529);
or U13131 (N_13131,N_11296,N_11905);
nor U13132 (N_13132,N_10842,N_10667);
and U13133 (N_13133,N_10764,N_11189);
nor U13134 (N_13134,N_10618,N_10608);
nand U13135 (N_13135,N_11998,N_11091);
or U13136 (N_13136,N_11146,N_11519);
xor U13137 (N_13137,N_10871,N_11824);
nor U13138 (N_13138,N_11861,N_10991);
and U13139 (N_13139,N_11896,N_11278);
nor U13140 (N_13140,N_11445,N_10501);
nor U13141 (N_13141,N_11138,N_10549);
xnor U13142 (N_13142,N_11585,N_11960);
or U13143 (N_13143,N_11720,N_11166);
and U13144 (N_13144,N_11171,N_11684);
nand U13145 (N_13145,N_11991,N_11886);
xor U13146 (N_13146,N_11352,N_10566);
nand U13147 (N_13147,N_10633,N_10534);
nor U13148 (N_13148,N_11857,N_10541);
or U13149 (N_13149,N_10562,N_10815);
nand U13150 (N_13150,N_10765,N_11919);
or U13151 (N_13151,N_11478,N_11886);
nor U13152 (N_13152,N_11442,N_11016);
nand U13153 (N_13153,N_10879,N_11362);
and U13154 (N_13154,N_10947,N_11745);
nor U13155 (N_13155,N_10862,N_11063);
and U13156 (N_13156,N_10967,N_11897);
or U13157 (N_13157,N_11626,N_11103);
or U13158 (N_13158,N_10539,N_10791);
xnor U13159 (N_13159,N_11151,N_11285);
or U13160 (N_13160,N_11013,N_11271);
and U13161 (N_13161,N_11180,N_10776);
xor U13162 (N_13162,N_11535,N_11084);
nand U13163 (N_13163,N_11881,N_11186);
nand U13164 (N_13164,N_11455,N_11962);
xnor U13165 (N_13165,N_11286,N_11533);
or U13166 (N_13166,N_10511,N_11809);
nand U13167 (N_13167,N_11387,N_10558);
nand U13168 (N_13168,N_11344,N_11037);
nor U13169 (N_13169,N_10840,N_10674);
xor U13170 (N_13170,N_11294,N_11940);
nor U13171 (N_13171,N_11243,N_10651);
nor U13172 (N_13172,N_11748,N_11923);
nor U13173 (N_13173,N_10957,N_11919);
nor U13174 (N_13174,N_11737,N_10623);
nor U13175 (N_13175,N_11895,N_10793);
nand U13176 (N_13176,N_10962,N_11731);
or U13177 (N_13177,N_10923,N_11142);
nand U13178 (N_13178,N_11194,N_11967);
nor U13179 (N_13179,N_10532,N_10701);
nor U13180 (N_13180,N_11399,N_11075);
nand U13181 (N_13181,N_11211,N_10634);
nor U13182 (N_13182,N_11033,N_11288);
and U13183 (N_13183,N_11817,N_11226);
and U13184 (N_13184,N_11308,N_11487);
nor U13185 (N_13185,N_10682,N_10549);
xnor U13186 (N_13186,N_11756,N_11067);
xor U13187 (N_13187,N_11424,N_11510);
or U13188 (N_13188,N_11367,N_10558);
xnor U13189 (N_13189,N_11098,N_10878);
or U13190 (N_13190,N_10897,N_11882);
xnor U13191 (N_13191,N_11616,N_11927);
nor U13192 (N_13192,N_11247,N_11822);
nor U13193 (N_13193,N_11646,N_10544);
and U13194 (N_13194,N_11125,N_10501);
and U13195 (N_13195,N_11337,N_10921);
nand U13196 (N_13196,N_10819,N_10914);
nand U13197 (N_13197,N_11757,N_11521);
nand U13198 (N_13198,N_10992,N_11493);
nand U13199 (N_13199,N_11444,N_11589);
or U13200 (N_13200,N_10680,N_11745);
and U13201 (N_13201,N_11706,N_11989);
xnor U13202 (N_13202,N_10751,N_11516);
and U13203 (N_13203,N_11954,N_10562);
nand U13204 (N_13204,N_11624,N_11382);
xnor U13205 (N_13205,N_11734,N_10684);
and U13206 (N_13206,N_11816,N_11695);
nand U13207 (N_13207,N_10755,N_11932);
xnor U13208 (N_13208,N_11637,N_10782);
xnor U13209 (N_13209,N_11956,N_10915);
xnor U13210 (N_13210,N_10760,N_10704);
or U13211 (N_13211,N_11198,N_11774);
and U13212 (N_13212,N_11739,N_10950);
and U13213 (N_13213,N_11254,N_11922);
or U13214 (N_13214,N_10976,N_11415);
and U13215 (N_13215,N_10783,N_11857);
nor U13216 (N_13216,N_10698,N_10608);
and U13217 (N_13217,N_11759,N_10511);
and U13218 (N_13218,N_11198,N_11459);
and U13219 (N_13219,N_11887,N_11503);
xor U13220 (N_13220,N_11289,N_10884);
or U13221 (N_13221,N_11293,N_11488);
nor U13222 (N_13222,N_11562,N_11641);
and U13223 (N_13223,N_10963,N_11007);
nand U13224 (N_13224,N_11149,N_10626);
nor U13225 (N_13225,N_11343,N_10822);
nor U13226 (N_13226,N_11269,N_10745);
and U13227 (N_13227,N_10573,N_11705);
nor U13228 (N_13228,N_11797,N_11772);
xor U13229 (N_13229,N_11606,N_10932);
and U13230 (N_13230,N_10927,N_10584);
and U13231 (N_13231,N_11139,N_11326);
and U13232 (N_13232,N_10833,N_10718);
and U13233 (N_13233,N_11104,N_10581);
and U13234 (N_13234,N_11470,N_11402);
xor U13235 (N_13235,N_11367,N_10827);
nor U13236 (N_13236,N_11238,N_11854);
or U13237 (N_13237,N_11898,N_11499);
nor U13238 (N_13238,N_10899,N_11461);
and U13239 (N_13239,N_11408,N_11625);
xnor U13240 (N_13240,N_11274,N_10765);
nor U13241 (N_13241,N_10596,N_11878);
or U13242 (N_13242,N_11155,N_10876);
and U13243 (N_13243,N_11284,N_11480);
nand U13244 (N_13244,N_11746,N_10778);
xor U13245 (N_13245,N_11292,N_11881);
and U13246 (N_13246,N_11270,N_10717);
and U13247 (N_13247,N_11116,N_11744);
and U13248 (N_13248,N_11996,N_10765);
nand U13249 (N_13249,N_10787,N_11128);
nand U13250 (N_13250,N_11417,N_11189);
xor U13251 (N_13251,N_10732,N_10961);
or U13252 (N_13252,N_11004,N_11532);
nor U13253 (N_13253,N_11562,N_10572);
or U13254 (N_13254,N_11477,N_10692);
and U13255 (N_13255,N_11223,N_11431);
and U13256 (N_13256,N_11005,N_11361);
or U13257 (N_13257,N_11726,N_11899);
nor U13258 (N_13258,N_10718,N_11860);
and U13259 (N_13259,N_11283,N_10882);
nand U13260 (N_13260,N_11189,N_11884);
nand U13261 (N_13261,N_10834,N_11179);
xor U13262 (N_13262,N_11290,N_11616);
nand U13263 (N_13263,N_11478,N_11182);
and U13264 (N_13264,N_11741,N_11655);
nand U13265 (N_13265,N_10752,N_11280);
nor U13266 (N_13266,N_11118,N_11246);
nor U13267 (N_13267,N_10649,N_11307);
xnor U13268 (N_13268,N_11847,N_11087);
xor U13269 (N_13269,N_11784,N_11266);
xor U13270 (N_13270,N_11607,N_11907);
and U13271 (N_13271,N_11208,N_11016);
xor U13272 (N_13272,N_11890,N_11776);
nand U13273 (N_13273,N_11794,N_10724);
nand U13274 (N_13274,N_11353,N_11055);
nand U13275 (N_13275,N_10711,N_11460);
or U13276 (N_13276,N_10542,N_10628);
and U13277 (N_13277,N_10556,N_11856);
nand U13278 (N_13278,N_11133,N_11012);
xnor U13279 (N_13279,N_11772,N_11439);
or U13280 (N_13280,N_10543,N_10923);
nor U13281 (N_13281,N_11882,N_10529);
and U13282 (N_13282,N_11652,N_11595);
nand U13283 (N_13283,N_11516,N_10943);
and U13284 (N_13284,N_10942,N_11537);
nor U13285 (N_13285,N_10677,N_10627);
and U13286 (N_13286,N_10722,N_11433);
nor U13287 (N_13287,N_11448,N_11344);
xnor U13288 (N_13288,N_11649,N_10509);
and U13289 (N_13289,N_11040,N_10699);
or U13290 (N_13290,N_10674,N_11871);
nand U13291 (N_13291,N_10874,N_11558);
and U13292 (N_13292,N_11455,N_11388);
or U13293 (N_13293,N_11124,N_11313);
and U13294 (N_13294,N_10633,N_10818);
xor U13295 (N_13295,N_10554,N_11735);
and U13296 (N_13296,N_10692,N_11057);
nor U13297 (N_13297,N_11578,N_10531);
and U13298 (N_13298,N_10837,N_11916);
nand U13299 (N_13299,N_11568,N_11493);
and U13300 (N_13300,N_11236,N_11112);
and U13301 (N_13301,N_11643,N_11171);
xor U13302 (N_13302,N_11967,N_11569);
xnor U13303 (N_13303,N_10635,N_11883);
and U13304 (N_13304,N_10519,N_11631);
nand U13305 (N_13305,N_11916,N_10780);
or U13306 (N_13306,N_11318,N_11075);
nand U13307 (N_13307,N_11146,N_11798);
nand U13308 (N_13308,N_11132,N_10566);
or U13309 (N_13309,N_10879,N_11371);
and U13310 (N_13310,N_11664,N_11814);
and U13311 (N_13311,N_10883,N_10722);
xnor U13312 (N_13312,N_10850,N_11841);
nor U13313 (N_13313,N_11697,N_11292);
nand U13314 (N_13314,N_11157,N_10556);
nand U13315 (N_13315,N_10523,N_11513);
nand U13316 (N_13316,N_11115,N_11876);
or U13317 (N_13317,N_10902,N_11385);
nor U13318 (N_13318,N_10573,N_11295);
nand U13319 (N_13319,N_11901,N_11208);
and U13320 (N_13320,N_11472,N_10507);
nand U13321 (N_13321,N_11705,N_10531);
nor U13322 (N_13322,N_11707,N_10762);
or U13323 (N_13323,N_11750,N_11976);
or U13324 (N_13324,N_11870,N_11183);
or U13325 (N_13325,N_10873,N_11616);
or U13326 (N_13326,N_11988,N_11924);
or U13327 (N_13327,N_10667,N_11504);
or U13328 (N_13328,N_11807,N_10784);
xor U13329 (N_13329,N_11589,N_11567);
or U13330 (N_13330,N_11121,N_11020);
or U13331 (N_13331,N_11494,N_11594);
xnor U13332 (N_13332,N_11526,N_11873);
or U13333 (N_13333,N_11929,N_11965);
and U13334 (N_13334,N_11395,N_11303);
xnor U13335 (N_13335,N_10658,N_11368);
or U13336 (N_13336,N_11550,N_11113);
nand U13337 (N_13337,N_11135,N_10939);
nand U13338 (N_13338,N_11857,N_11768);
and U13339 (N_13339,N_11143,N_11665);
xnor U13340 (N_13340,N_11435,N_10557);
nor U13341 (N_13341,N_11666,N_11157);
nand U13342 (N_13342,N_10749,N_11178);
nor U13343 (N_13343,N_10729,N_11975);
or U13344 (N_13344,N_10904,N_10781);
and U13345 (N_13345,N_11302,N_11828);
nor U13346 (N_13346,N_11176,N_11846);
xor U13347 (N_13347,N_11901,N_11669);
xnor U13348 (N_13348,N_11573,N_10819);
nand U13349 (N_13349,N_11507,N_11419);
nor U13350 (N_13350,N_11992,N_10779);
and U13351 (N_13351,N_11165,N_10863);
xor U13352 (N_13352,N_11700,N_11114);
and U13353 (N_13353,N_10673,N_11854);
nor U13354 (N_13354,N_11982,N_11033);
nor U13355 (N_13355,N_11309,N_11151);
nor U13356 (N_13356,N_11460,N_11481);
nand U13357 (N_13357,N_10932,N_11126);
nor U13358 (N_13358,N_11574,N_11549);
xnor U13359 (N_13359,N_11155,N_11956);
nor U13360 (N_13360,N_11341,N_10999);
nand U13361 (N_13361,N_10869,N_10865);
xnor U13362 (N_13362,N_11187,N_11121);
xor U13363 (N_13363,N_11258,N_11415);
nor U13364 (N_13364,N_11943,N_11163);
xor U13365 (N_13365,N_11549,N_10547);
and U13366 (N_13366,N_11271,N_11308);
nand U13367 (N_13367,N_11832,N_11666);
nand U13368 (N_13368,N_11072,N_10753);
nand U13369 (N_13369,N_11095,N_11156);
nor U13370 (N_13370,N_11506,N_11640);
or U13371 (N_13371,N_10595,N_11532);
nor U13372 (N_13372,N_11333,N_10606);
and U13373 (N_13373,N_11930,N_11066);
nand U13374 (N_13374,N_10663,N_10977);
nand U13375 (N_13375,N_11733,N_10508);
and U13376 (N_13376,N_10651,N_11920);
nor U13377 (N_13377,N_10502,N_11221);
nand U13378 (N_13378,N_11378,N_11801);
or U13379 (N_13379,N_11964,N_11742);
and U13380 (N_13380,N_10831,N_11400);
nand U13381 (N_13381,N_11216,N_11281);
nand U13382 (N_13382,N_10723,N_10599);
nor U13383 (N_13383,N_11176,N_10985);
and U13384 (N_13384,N_10818,N_11435);
xor U13385 (N_13385,N_11350,N_11571);
and U13386 (N_13386,N_11802,N_11012);
or U13387 (N_13387,N_10697,N_10783);
xnor U13388 (N_13388,N_10725,N_11156);
and U13389 (N_13389,N_11890,N_10815);
nor U13390 (N_13390,N_10914,N_11012);
xor U13391 (N_13391,N_11810,N_11628);
and U13392 (N_13392,N_10585,N_10832);
and U13393 (N_13393,N_11440,N_11622);
xnor U13394 (N_13394,N_11070,N_11753);
and U13395 (N_13395,N_11369,N_11592);
nor U13396 (N_13396,N_11544,N_11749);
and U13397 (N_13397,N_11658,N_11699);
nand U13398 (N_13398,N_11716,N_10849);
or U13399 (N_13399,N_10671,N_10550);
and U13400 (N_13400,N_11546,N_10960);
and U13401 (N_13401,N_11508,N_11983);
and U13402 (N_13402,N_11495,N_11071);
nand U13403 (N_13403,N_10970,N_11432);
xor U13404 (N_13404,N_11907,N_11727);
and U13405 (N_13405,N_11233,N_11615);
xor U13406 (N_13406,N_10992,N_11065);
and U13407 (N_13407,N_11911,N_10985);
and U13408 (N_13408,N_11791,N_11893);
nor U13409 (N_13409,N_10902,N_11753);
xnor U13410 (N_13410,N_11531,N_10825);
nor U13411 (N_13411,N_10760,N_11399);
xor U13412 (N_13412,N_11697,N_11491);
nor U13413 (N_13413,N_11569,N_11140);
and U13414 (N_13414,N_10707,N_10728);
nand U13415 (N_13415,N_10863,N_11608);
or U13416 (N_13416,N_11758,N_10718);
or U13417 (N_13417,N_11322,N_10631);
and U13418 (N_13418,N_11270,N_11960);
xor U13419 (N_13419,N_11681,N_11565);
xnor U13420 (N_13420,N_10533,N_11925);
nor U13421 (N_13421,N_10550,N_10913);
and U13422 (N_13422,N_11258,N_11734);
nand U13423 (N_13423,N_11672,N_11164);
xor U13424 (N_13424,N_11198,N_10622);
and U13425 (N_13425,N_11270,N_11330);
nand U13426 (N_13426,N_11899,N_11214);
nor U13427 (N_13427,N_10660,N_11531);
xnor U13428 (N_13428,N_11301,N_11648);
xor U13429 (N_13429,N_10997,N_11598);
nand U13430 (N_13430,N_11400,N_10615);
and U13431 (N_13431,N_11279,N_11879);
nor U13432 (N_13432,N_10637,N_11076);
nor U13433 (N_13433,N_11033,N_11164);
and U13434 (N_13434,N_10745,N_11150);
nand U13435 (N_13435,N_11663,N_11519);
or U13436 (N_13436,N_11068,N_10938);
nor U13437 (N_13437,N_11821,N_11732);
and U13438 (N_13438,N_11506,N_10958);
nor U13439 (N_13439,N_11362,N_11814);
nor U13440 (N_13440,N_11131,N_11391);
xnor U13441 (N_13441,N_10953,N_11534);
xnor U13442 (N_13442,N_11964,N_10664);
nor U13443 (N_13443,N_10592,N_11875);
nand U13444 (N_13444,N_10687,N_11817);
and U13445 (N_13445,N_11592,N_11848);
xnor U13446 (N_13446,N_11089,N_10738);
nor U13447 (N_13447,N_10865,N_11275);
nor U13448 (N_13448,N_11826,N_11657);
xor U13449 (N_13449,N_11194,N_11390);
or U13450 (N_13450,N_10884,N_10632);
or U13451 (N_13451,N_11057,N_11926);
nor U13452 (N_13452,N_11503,N_11765);
nor U13453 (N_13453,N_11545,N_11678);
or U13454 (N_13454,N_11707,N_10992);
xnor U13455 (N_13455,N_11636,N_11912);
nor U13456 (N_13456,N_11869,N_10717);
or U13457 (N_13457,N_11717,N_11594);
or U13458 (N_13458,N_11723,N_10839);
and U13459 (N_13459,N_11923,N_11730);
or U13460 (N_13460,N_10887,N_10767);
and U13461 (N_13461,N_11238,N_11147);
and U13462 (N_13462,N_11894,N_10696);
and U13463 (N_13463,N_11601,N_11575);
or U13464 (N_13464,N_11175,N_11244);
or U13465 (N_13465,N_11551,N_11150);
xnor U13466 (N_13466,N_11906,N_11377);
nand U13467 (N_13467,N_11020,N_10765);
xnor U13468 (N_13468,N_11664,N_10659);
or U13469 (N_13469,N_10964,N_10824);
xor U13470 (N_13470,N_10759,N_11085);
nand U13471 (N_13471,N_10517,N_10940);
nand U13472 (N_13472,N_11432,N_10538);
and U13473 (N_13473,N_11001,N_10506);
nand U13474 (N_13474,N_11927,N_10694);
nand U13475 (N_13475,N_10839,N_11230);
or U13476 (N_13476,N_11670,N_11849);
nor U13477 (N_13477,N_11457,N_10793);
nor U13478 (N_13478,N_11484,N_10728);
or U13479 (N_13479,N_11476,N_11101);
xnor U13480 (N_13480,N_11457,N_11033);
nor U13481 (N_13481,N_10768,N_11653);
or U13482 (N_13482,N_11933,N_11983);
xnor U13483 (N_13483,N_11806,N_11763);
nand U13484 (N_13484,N_10649,N_11148);
or U13485 (N_13485,N_11763,N_11392);
nand U13486 (N_13486,N_11215,N_10992);
and U13487 (N_13487,N_11892,N_11226);
nor U13488 (N_13488,N_10940,N_11508);
or U13489 (N_13489,N_11561,N_10770);
and U13490 (N_13490,N_11127,N_11609);
xnor U13491 (N_13491,N_11850,N_11236);
xnor U13492 (N_13492,N_11795,N_11322);
and U13493 (N_13493,N_11826,N_11638);
nand U13494 (N_13494,N_11860,N_11843);
or U13495 (N_13495,N_11100,N_10715);
xnor U13496 (N_13496,N_11511,N_11148);
and U13497 (N_13497,N_11306,N_11597);
nor U13498 (N_13498,N_10884,N_10996);
nor U13499 (N_13499,N_10500,N_11629);
xor U13500 (N_13500,N_12675,N_13208);
or U13501 (N_13501,N_12437,N_13345);
or U13502 (N_13502,N_13029,N_12701);
or U13503 (N_13503,N_12497,N_12456);
and U13504 (N_13504,N_13230,N_12649);
xor U13505 (N_13505,N_12622,N_13490);
and U13506 (N_13506,N_13065,N_12094);
xor U13507 (N_13507,N_13116,N_12699);
or U13508 (N_13508,N_12284,N_12875);
nand U13509 (N_13509,N_12042,N_12218);
or U13510 (N_13510,N_12950,N_12796);
nor U13511 (N_13511,N_12627,N_12471);
and U13512 (N_13512,N_13396,N_12345);
nand U13513 (N_13513,N_12269,N_13172);
nor U13514 (N_13514,N_12494,N_13128);
and U13515 (N_13515,N_12669,N_13434);
nor U13516 (N_13516,N_13046,N_12524);
nand U13517 (N_13517,N_12697,N_13427);
nor U13518 (N_13518,N_12806,N_13071);
xor U13519 (N_13519,N_13151,N_13095);
xor U13520 (N_13520,N_12883,N_13120);
or U13521 (N_13521,N_13248,N_13359);
and U13522 (N_13522,N_12947,N_12886);
xnor U13523 (N_13523,N_13090,N_12346);
nor U13524 (N_13524,N_12526,N_12703);
nor U13525 (N_13525,N_12731,N_12339);
or U13526 (N_13526,N_12532,N_12992);
nand U13527 (N_13527,N_12889,N_12679);
nor U13528 (N_13528,N_12977,N_12991);
or U13529 (N_13529,N_12579,N_13408);
or U13530 (N_13530,N_12152,N_12521);
nand U13531 (N_13531,N_12079,N_12890);
nor U13532 (N_13532,N_12563,N_13253);
or U13533 (N_13533,N_13334,N_12747);
xor U13534 (N_13534,N_13291,N_12088);
nor U13535 (N_13535,N_13107,N_12067);
or U13536 (N_13536,N_13101,N_13482);
nor U13537 (N_13537,N_13064,N_12343);
xor U13538 (N_13538,N_12432,N_13495);
nand U13539 (N_13539,N_12485,N_12593);
and U13540 (N_13540,N_13104,N_13215);
nor U13541 (N_13541,N_13382,N_12382);
nor U13542 (N_13542,N_12828,N_12658);
xor U13543 (N_13543,N_12283,N_13445);
or U13544 (N_13544,N_12785,N_12989);
nand U13545 (N_13545,N_12009,N_12290);
or U13546 (N_13546,N_13013,N_12921);
and U13547 (N_13547,N_12619,N_13349);
nor U13548 (N_13548,N_13370,N_13143);
nor U13549 (N_13549,N_12849,N_12933);
nand U13550 (N_13550,N_13337,N_13368);
and U13551 (N_13551,N_12920,N_12827);
and U13552 (N_13552,N_12842,N_13367);
and U13553 (N_13553,N_13252,N_12516);
and U13554 (N_13554,N_12909,N_12967);
and U13555 (N_13555,N_12755,N_12436);
or U13556 (N_13556,N_12386,N_12234);
nor U13557 (N_13557,N_12771,N_12417);
and U13558 (N_13558,N_12200,N_12207);
nand U13559 (N_13559,N_13493,N_12262);
xnor U13560 (N_13560,N_13134,N_13273);
nor U13561 (N_13561,N_13148,N_12746);
or U13562 (N_13562,N_12765,N_12766);
nand U13563 (N_13563,N_12550,N_12279);
or U13564 (N_13564,N_13147,N_12098);
or U13565 (N_13565,N_12605,N_13006);
nor U13566 (N_13566,N_12617,N_12134);
and U13567 (N_13567,N_12435,N_12880);
nor U13568 (N_13568,N_12916,N_12519);
nand U13569 (N_13569,N_12544,N_13199);
or U13570 (N_13570,N_13381,N_12130);
nor U13571 (N_13571,N_12076,N_12195);
xnor U13572 (N_13572,N_13183,N_12548);
or U13573 (N_13573,N_13470,N_12955);
or U13574 (N_13574,N_13043,N_12392);
nor U13575 (N_13575,N_12214,N_12710);
nor U13576 (N_13576,N_13339,N_13110);
or U13577 (N_13577,N_12807,N_13139);
nor U13578 (N_13578,N_12228,N_12882);
xor U13579 (N_13579,N_12112,N_13330);
or U13580 (N_13580,N_12668,N_12408);
or U13581 (N_13581,N_12155,N_12135);
nand U13582 (N_13582,N_13193,N_12581);
xnor U13583 (N_13583,N_12501,N_13233);
nand U13584 (N_13584,N_12015,N_12705);
or U13585 (N_13585,N_12823,N_12227);
xor U13586 (N_13586,N_12203,N_13210);
nand U13587 (N_13587,N_13177,N_12693);
and U13588 (N_13588,N_12085,N_12483);
nor U13589 (N_13589,N_12154,N_12953);
or U13590 (N_13590,N_12707,N_12175);
nand U13591 (N_13591,N_13073,N_12303);
xnor U13592 (N_13592,N_13093,N_13196);
nor U13593 (N_13593,N_12212,N_12353);
xnor U13594 (N_13594,N_13483,N_13133);
nand U13595 (N_13595,N_12294,N_12420);
and U13596 (N_13596,N_12254,N_12180);
nor U13597 (N_13597,N_12728,N_12601);
xnor U13598 (N_13598,N_12209,N_13258);
nand U13599 (N_13599,N_12610,N_12572);
nor U13600 (N_13600,N_12414,N_12852);
or U13601 (N_13601,N_12413,N_12522);
and U13602 (N_13602,N_12751,N_12691);
nand U13603 (N_13603,N_12841,N_12275);
xor U13604 (N_13604,N_13352,N_12257);
and U13605 (N_13605,N_13220,N_12385);
nor U13606 (N_13606,N_12517,N_12141);
nand U13607 (N_13607,N_13243,N_12231);
nor U13608 (N_13608,N_12598,N_12259);
nor U13609 (N_13609,N_12565,N_12110);
xnor U13610 (N_13610,N_12684,N_13435);
nand U13611 (N_13611,N_12356,N_12282);
nand U13612 (N_13612,N_12726,N_13040);
nand U13613 (N_13613,N_12018,N_13300);
and U13614 (N_13614,N_13092,N_12361);
or U13615 (N_13615,N_12270,N_13262);
nand U13616 (N_13616,N_12850,N_12127);
nor U13617 (N_13617,N_12545,N_13308);
and U13618 (N_13618,N_13010,N_12370);
xnor U13619 (N_13619,N_13179,N_12190);
or U13620 (N_13620,N_13355,N_12367);
nor U13621 (N_13621,N_13226,N_13269);
nand U13622 (N_13622,N_12744,N_13313);
nor U13623 (N_13623,N_13437,N_12578);
and U13624 (N_13624,N_13433,N_12981);
nand U13625 (N_13625,N_12419,N_12586);
nor U13626 (N_13626,N_12451,N_12553);
xor U13627 (N_13627,N_12647,N_13084);
nor U13628 (N_13628,N_12122,N_12253);
nand U13629 (N_13629,N_13447,N_13260);
and U13630 (N_13630,N_12761,N_13096);
and U13631 (N_13631,N_13033,N_12039);
xor U13632 (N_13632,N_12910,N_12655);
nand U13633 (N_13633,N_12201,N_13247);
nor U13634 (N_13634,N_12278,N_12782);
xnor U13635 (N_13635,N_12260,N_12873);
or U13636 (N_13636,N_13327,N_12441);
nor U13637 (N_13637,N_13332,N_13008);
nor U13638 (N_13638,N_12809,N_12969);
nor U13639 (N_13639,N_13238,N_13217);
xnor U13640 (N_13640,N_13000,N_12964);
nor U13641 (N_13641,N_13244,N_12261);
nor U13642 (N_13642,N_13213,N_13072);
xnor U13643 (N_13643,N_13054,N_12461);
nor U13644 (N_13644,N_12005,N_13003);
xor U13645 (N_13645,N_13295,N_13305);
nor U13646 (N_13646,N_13192,N_13232);
and U13647 (N_13647,N_12695,N_13146);
or U13648 (N_13648,N_12006,N_12355);
and U13649 (N_13649,N_12416,N_12080);
nor U13650 (N_13650,N_13201,N_12641);
xor U13651 (N_13651,N_13378,N_12129);
nand U13652 (N_13652,N_12944,N_12439);
or U13653 (N_13653,N_12768,N_13289);
and U13654 (N_13654,N_12819,N_12597);
nand U13655 (N_13655,N_12896,N_12354);
xor U13656 (N_13656,N_12198,N_12443);
nor U13657 (N_13657,N_12963,N_13286);
or U13658 (N_13658,N_12791,N_12558);
nor U13659 (N_13659,N_13162,N_12723);
nor U13660 (N_13660,N_12583,N_12412);
xor U13661 (N_13661,N_12833,N_12786);
or U13662 (N_13662,N_12452,N_12683);
or U13663 (N_13663,N_12325,N_13460);
or U13664 (N_13664,N_12531,N_12749);
nand U13665 (N_13665,N_13156,N_12799);
xnor U13666 (N_13666,N_12378,N_12616);
or U13667 (N_13667,N_12948,N_12090);
xor U13668 (N_13668,N_12245,N_12306);
or U13669 (N_13669,N_12631,N_12041);
xor U13670 (N_13670,N_12255,N_12169);
and U13671 (N_13671,N_13113,N_13492);
nand U13672 (N_13672,N_12859,N_12189);
xnor U13673 (N_13673,N_12584,N_12008);
xor U13674 (N_13674,N_13324,N_12037);
nand U13675 (N_13675,N_12241,N_12341);
xnor U13676 (N_13676,N_12300,N_12700);
or U13677 (N_13677,N_13325,N_13060);
and U13678 (N_13678,N_12727,N_12124);
and U13679 (N_13679,N_12721,N_13121);
or U13680 (N_13680,N_12934,N_12478);
and U13681 (N_13681,N_12863,N_12680);
xor U13682 (N_13682,N_12315,N_12470);
xor U13683 (N_13683,N_12793,N_12176);
or U13684 (N_13684,N_13221,N_12525);
xnor U13685 (N_13685,N_12638,N_12732);
and U13686 (N_13686,N_13207,N_12380);
or U13687 (N_13687,N_12800,N_12252);
xnor U13688 (N_13688,N_13016,N_12011);
or U13689 (N_13689,N_12359,N_12552);
nor U13690 (N_13690,N_12029,N_13271);
xor U13691 (N_13691,N_12895,N_13356);
nand U13692 (N_13692,N_12081,N_12832);
or U13693 (N_13693,N_13028,N_12131);
xnor U13694 (N_13694,N_13266,N_12686);
and U13695 (N_13695,N_13392,N_13170);
xor U13696 (N_13696,N_12139,N_12932);
or U13697 (N_13697,N_13165,N_12074);
or U13698 (N_13698,N_12936,N_12236);
nor U13699 (N_13699,N_12321,N_13117);
or U13700 (N_13700,N_12543,N_13280);
or U13701 (N_13701,N_12116,N_12106);
and U13702 (N_13702,N_12970,N_12220);
xor U13703 (N_13703,N_12159,N_12289);
xnor U13704 (N_13704,N_12855,N_12802);
nand U13705 (N_13705,N_12724,N_12334);
xor U13706 (N_13706,N_12857,N_12708);
nand U13707 (N_13707,N_13395,N_12459);
or U13708 (N_13708,N_13274,N_13077);
xor U13709 (N_13709,N_13469,N_12838);
nor U13710 (N_13710,N_12835,N_12375);
xor U13711 (N_13711,N_12021,N_13276);
nand U13712 (N_13712,N_12312,N_12898);
nor U13713 (N_13713,N_12313,N_13414);
nor U13714 (N_13714,N_12960,N_13144);
xnor U13715 (N_13715,N_12824,N_12671);
nand U13716 (N_13716,N_13188,N_12070);
nand U13717 (N_13717,N_12718,N_12266);
xor U13718 (N_13718,N_12128,N_12528);
xnor U13719 (N_13719,N_12017,N_13239);
xor U13720 (N_13720,N_12337,N_13191);
or U13721 (N_13721,N_12144,N_12538);
nor U13722 (N_13722,N_12784,N_12058);
nor U13723 (N_13723,N_13039,N_13374);
nor U13724 (N_13724,N_13441,N_12285);
and U13725 (N_13725,N_12347,N_12156);
nand U13726 (N_13726,N_12957,N_12892);
or U13727 (N_13727,N_12150,N_12491);
xor U13728 (N_13728,N_12506,N_13049);
or U13729 (N_13729,N_12663,N_13479);
or U13730 (N_13730,N_13254,N_12351);
or U13731 (N_13731,N_13453,N_12427);
nand U13732 (N_13732,N_13058,N_12546);
and U13733 (N_13733,N_12666,N_12625);
or U13734 (N_13734,N_12047,N_12908);
nand U13735 (N_13735,N_12945,N_12946);
nor U13736 (N_13736,N_12462,N_13027);
xor U13737 (N_13737,N_12899,N_12052);
or U13738 (N_13738,N_12000,N_13108);
or U13739 (N_13739,N_12826,N_12320);
nand U13740 (N_13740,N_12066,N_13444);
xnor U13741 (N_13741,N_12783,N_12535);
nand U13742 (N_13742,N_13203,N_12002);
nand U13743 (N_13743,N_12170,N_13467);
and U13744 (N_13744,N_13336,N_13393);
xor U13745 (N_13745,N_12615,N_13042);
or U13746 (N_13746,N_12575,N_12221);
xnor U13747 (N_13747,N_12962,N_12258);
xnor U13748 (N_13748,N_13184,N_13481);
and U13749 (N_13749,N_12089,N_13489);
xnor U13750 (N_13750,N_12770,N_12268);
and U13751 (N_13751,N_12878,N_13038);
nand U13752 (N_13752,N_12696,N_12958);
nand U13753 (N_13753,N_12928,N_12464);
nand U13754 (N_13754,N_13261,N_12556);
and U13755 (N_13755,N_13399,N_12153);
or U13756 (N_13756,N_13420,N_12562);
nand U13757 (N_13757,N_12810,N_12888);
nand U13758 (N_13758,N_12979,N_13487);
or U13759 (N_13759,N_12288,N_13051);
and U13760 (N_13760,N_13080,N_12032);
xnor U13761 (N_13761,N_12287,N_12233);
or U13762 (N_13762,N_12792,N_12376);
nand U13763 (N_13763,N_12816,N_12238);
nor U13764 (N_13764,N_12271,N_12702);
xor U13765 (N_13765,N_12330,N_12489);
nor U13766 (N_13766,N_13229,N_12788);
nor U13767 (N_13767,N_13005,N_12038);
nand U13768 (N_13768,N_12711,N_12426);
nand U13769 (N_13769,N_13100,N_12912);
xor U13770 (N_13770,N_13315,N_12564);
and U13771 (N_13771,N_13440,N_13344);
nand U13772 (N_13772,N_12324,N_12049);
or U13773 (N_13773,N_12603,N_12879);
nand U13774 (N_13774,N_12588,N_12894);
xnor U13775 (N_13775,N_12160,N_12650);
nor U13776 (N_13776,N_13316,N_12537);
xnor U13777 (N_13777,N_12511,N_13214);
nor U13778 (N_13778,N_13034,N_13255);
and U13779 (N_13779,N_13057,N_12352);
nand U13780 (N_13780,N_12273,N_12225);
xnor U13781 (N_13781,N_13087,N_13474);
and U13782 (N_13782,N_12541,N_13137);
nand U13783 (N_13783,N_12274,N_13175);
or U13784 (N_13784,N_13459,N_12309);
and U13785 (N_13785,N_13045,N_13242);
nor U13786 (N_13786,N_12188,N_12196);
nor U13787 (N_13787,N_12513,N_12034);
nand U13788 (N_13788,N_13299,N_13023);
and U13789 (N_13789,N_13485,N_12348);
and U13790 (N_13790,N_13112,N_12120);
nor U13791 (N_13791,N_12014,N_13142);
nand U13792 (N_13792,N_12529,N_13135);
and U13793 (N_13793,N_13462,N_12972);
nand U13794 (N_13794,N_12893,N_12192);
or U13795 (N_13795,N_12372,N_13302);
or U13796 (N_13796,N_12900,N_13007);
nand U13797 (N_13797,N_12256,N_12764);
nand U13798 (N_13798,N_13473,N_12599);
xor U13799 (N_13799,N_12687,N_13081);
or U13800 (N_13800,N_12682,N_13168);
nor U13801 (N_13801,N_12993,N_13197);
and U13802 (N_13802,N_12871,N_12568);
and U13803 (N_13803,N_12971,N_12381);
nand U13804 (N_13804,N_12719,N_13138);
or U13805 (N_13805,N_12499,N_12571);
nor U13806 (N_13806,N_12400,N_13363);
nor U13807 (N_13807,N_13037,N_12713);
or U13808 (N_13808,N_13418,N_12569);
xor U13809 (N_13809,N_12142,N_12740);
and U13810 (N_13810,N_12342,N_13109);
or U13811 (N_13811,N_13155,N_13307);
nand U13812 (N_13812,N_13451,N_13257);
xnor U13813 (N_13813,N_12813,N_12643);
xor U13814 (N_13814,N_12917,N_13259);
and U13815 (N_13815,N_13102,N_12421);
or U13816 (N_13816,N_13141,N_13019);
and U13817 (N_13817,N_12118,N_12481);
nor U13818 (N_13818,N_13311,N_12418);
nand U13819 (N_13819,N_12186,N_12523);
and U13820 (N_13820,N_13303,N_12618);
xnor U13821 (N_13821,N_12798,N_12063);
xnor U13822 (N_13822,N_13486,N_13263);
xnor U13823 (N_13823,N_12398,N_12165);
or U13824 (N_13824,N_12885,N_12316);
xor U13825 (N_13825,N_12554,N_12004);
nor U13826 (N_13826,N_13119,N_13091);
nor U13827 (N_13827,N_12665,N_12405);
and U13828 (N_13828,N_13386,N_13373);
xnor U13829 (N_13829,N_12045,N_13224);
and U13830 (N_13830,N_12639,N_13428);
nand U13831 (N_13831,N_12903,N_12612);
nor U13832 (N_13832,N_12735,N_12265);
and U13833 (N_13833,N_13180,N_12092);
and U13834 (N_13834,N_12407,N_12843);
xnor U13835 (N_13835,N_13237,N_13484);
nor U13836 (N_13836,N_12741,N_13331);
xnor U13837 (N_13837,N_12716,N_12108);
and U13838 (N_13838,N_12121,N_12390);
nor U13839 (N_13839,N_12831,N_12183);
and U13840 (N_13840,N_13338,N_12549);
or U13841 (N_13841,N_13290,N_12656);
or U13842 (N_13842,N_12698,N_12725);
and U13843 (N_13843,N_12357,N_12825);
nor U13844 (N_13844,N_12117,N_12445);
nand U13845 (N_13845,N_12628,N_12263);
or U13846 (N_13846,N_12817,N_12847);
and U13847 (N_13847,N_12344,N_12502);
nor U13848 (N_13848,N_12336,N_13178);
nand U13849 (N_13849,N_12514,N_12976);
or U13850 (N_13850,N_13089,N_12566);
and U13851 (N_13851,N_12844,N_12943);
and U13852 (N_13852,N_12590,N_13014);
nor U13853 (N_13853,N_12866,N_13041);
nor U13854 (N_13854,N_12520,N_12387);
nand U13855 (N_13855,N_12447,N_12988);
or U13856 (N_13856,N_12101,N_12397);
nor U13857 (N_13857,N_12931,N_12064);
nor U13858 (N_13858,N_12775,N_12830);
nand U13859 (N_13859,N_12125,N_13383);
or U13860 (N_13860,N_13153,N_12776);
and U13861 (N_13861,N_12677,N_12480);
nor U13862 (N_13862,N_13472,N_13118);
or U13863 (N_13863,N_12887,N_12404);
xor U13864 (N_13864,N_13353,N_12001);
xnor U13865 (N_13865,N_12918,N_13401);
nor U13866 (N_13866,N_12244,N_12409);
xnor U13867 (N_13867,N_13278,N_12086);
or U13868 (N_13868,N_13205,N_13463);
nor U13869 (N_13869,N_13127,N_12465);
nor U13870 (N_13870,N_12595,N_12384);
xor U13871 (N_13871,N_12422,N_12512);
nand U13872 (N_13872,N_12267,N_12291);
xnor U13873 (N_13873,N_12822,N_13202);
nand U13874 (N_13874,N_13284,N_13129);
or U13875 (N_13875,N_13377,N_12318);
or U13876 (N_13876,N_12580,N_12591);
nand U13877 (N_13877,N_12230,N_12667);
nand U13878 (N_13878,N_13249,N_12795);
and U13879 (N_13879,N_13319,N_13044);
and U13880 (N_13880,N_13075,N_12814);
xor U13881 (N_13881,N_12999,N_12745);
and U13882 (N_13882,N_12363,N_13343);
or U13883 (N_13883,N_12046,N_13412);
nand U13884 (N_13884,N_13328,N_13456);
nand U13885 (N_13885,N_12304,N_13194);
nand U13886 (N_13886,N_12623,N_12206);
nand U13887 (N_13887,N_12335,N_12406);
xnor U13888 (N_13888,N_12652,N_12661);
nor U13889 (N_13889,N_12906,N_13436);
and U13890 (N_13890,N_12013,N_12468);
nand U13891 (N_13891,N_12298,N_12488);
and U13892 (N_13892,N_13068,N_12057);
or U13893 (N_13893,N_12614,N_12323);
or U13894 (N_13894,N_12688,N_12033);
nand U13895 (N_13895,N_12848,N_12854);
nand U13896 (N_13896,N_12737,N_13018);
xor U13897 (N_13897,N_12482,N_12199);
xor U13898 (N_13898,N_12450,N_13391);
or U13899 (N_13899,N_12082,N_13145);
xor U13900 (N_13900,N_12179,N_12808);
and U13901 (N_13901,N_12856,N_12305);
xor U13902 (N_13902,N_13225,N_13407);
nand U13903 (N_13903,N_12508,N_13275);
and U13904 (N_13904,N_12389,N_12840);
xnor U13905 (N_13905,N_12503,N_12358);
xor U13906 (N_13906,N_13466,N_12994);
and U13907 (N_13907,N_12924,N_12927);
xor U13908 (N_13908,N_12901,N_12237);
xor U13909 (N_13909,N_13468,N_12007);
or U13910 (N_13910,N_12243,N_12454);
nand U13911 (N_13911,N_12054,N_12985);
and U13912 (N_13912,N_12954,N_12393);
and U13913 (N_13913,N_12694,N_13372);
or U13914 (N_13914,N_13314,N_12171);
nand U13915 (N_13915,N_12197,N_12959);
xnor U13916 (N_13916,N_12010,N_12410);
nor U13917 (N_13917,N_12941,N_12664);
or U13918 (N_13918,N_13497,N_12922);
nand U13919 (N_13919,N_12487,N_12310);
and U13920 (N_13920,N_12913,N_12191);
nor U13921 (N_13921,N_12217,N_12624);
or U13922 (N_13922,N_13264,N_12987);
nor U13923 (N_13923,N_13322,N_12115);
xor U13924 (N_13924,N_12251,N_13326);
nand U13925 (N_13925,N_13002,N_13052);
or U13926 (N_13926,N_12996,N_12322);
nand U13927 (N_13927,N_12036,N_12103);
nor U13928 (N_13928,N_13158,N_12003);
nor U13929 (N_13929,N_12560,N_12250);
nand U13930 (N_13930,N_12174,N_13149);
xnor U13931 (N_13931,N_13390,N_13169);
nand U13932 (N_13932,N_12479,N_12570);
xnor U13933 (N_13933,N_13020,N_13222);
nand U13934 (N_13934,N_13364,N_13419);
or U13935 (N_13935,N_12084,N_13397);
or U13936 (N_13936,N_13333,N_13425);
and U13937 (N_13937,N_13298,N_12019);
or U13938 (N_13938,N_13021,N_12317);
or U13939 (N_13939,N_13310,N_12223);
nand U13940 (N_13940,N_12507,N_13312);
nand U13941 (N_13941,N_13024,N_12736);
or U13942 (N_13942,N_13360,N_12247);
or U13943 (N_13943,N_13415,N_12219);
nand U13944 (N_13944,N_12096,N_13219);
or U13945 (N_13945,N_12016,N_12242);
or U13946 (N_13946,N_12099,N_13061);
or U13947 (N_13947,N_12690,N_13380);
nand U13948 (N_13948,N_13410,N_13454);
xor U13949 (N_13949,N_12202,N_12653);
nand U13950 (N_13950,N_12442,N_12557);
and U13951 (N_13951,N_12821,N_12048);
or U13952 (N_13952,N_12477,N_13288);
xnor U13953 (N_13953,N_12138,N_13405);
nand U13954 (N_13954,N_12781,N_12148);
or U13955 (N_13955,N_13082,N_12975);
and U13956 (N_13956,N_13228,N_13130);
xor U13957 (N_13957,N_12145,N_12637);
nand U13958 (N_13958,N_12773,N_12423);
and U13959 (N_13959,N_12143,N_12555);
xor U13960 (N_13960,N_12635,N_12277);
and U13961 (N_13961,N_13223,N_13036);
and U13962 (N_13962,N_12163,N_12069);
nand U13963 (N_13963,N_12172,N_12659);
and U13964 (N_13964,N_12026,N_13422);
nand U13965 (N_13965,N_12168,N_12496);
nand U13966 (N_13966,N_13190,N_12573);
or U13967 (N_13967,N_12567,N_12071);
xnor U13968 (N_13968,N_12978,N_12332);
nor U13969 (N_13969,N_12474,N_12877);
or U13970 (N_13970,N_13204,N_12062);
or U13971 (N_13971,N_13017,N_12504);
xor U13972 (N_13972,N_12329,N_13309);
or U13973 (N_13973,N_12640,N_12208);
or U13974 (N_13974,N_12911,N_12072);
and U13975 (N_13975,N_12246,N_12113);
xnor U13976 (N_13976,N_13362,N_13235);
xor U13977 (N_13977,N_12493,N_12391);
nor U13978 (N_13978,N_12527,N_12301);
xor U13979 (N_13979,N_12986,N_12951);
and U13980 (N_13980,N_12040,N_13176);
and U13981 (N_13981,N_13211,N_12308);
xnor U13982 (N_13982,N_12053,N_12073);
nor U13983 (N_13983,N_12399,N_12743);
or U13984 (N_13984,N_12660,N_13423);
or U13985 (N_13985,N_13212,N_12248);
nor U13986 (N_13986,N_12876,N_12606);
or U13987 (N_13987,N_13186,N_12297);
nor U13988 (N_13988,N_12107,N_12956);
nor U13989 (N_13989,N_13056,N_13251);
nor U13990 (N_13990,N_12714,N_13371);
or U13991 (N_13991,N_12974,N_12022);
and U13992 (N_13992,N_12651,N_13004);
nand U13993 (N_13993,N_13458,N_13384);
nor U13994 (N_13994,N_13099,N_13358);
or U13995 (N_13995,N_13402,N_12068);
and U13996 (N_13996,N_13431,N_12379);
or U13997 (N_13997,N_13385,N_12184);
nor U13998 (N_13998,N_12146,N_13069);
or U13999 (N_13999,N_13050,N_13231);
or U14000 (N_14000,N_12777,N_12025);
xor U14001 (N_14001,N_12331,N_13446);
nand U14002 (N_14002,N_13079,N_12167);
nor U14003 (N_14003,N_12604,N_12050);
and U14004 (N_14004,N_13150,N_12868);
nand U14005 (N_14005,N_12440,N_13185);
nor U14006 (N_14006,N_13256,N_12884);
xor U14007 (N_14007,N_12360,N_12292);
nor U14008 (N_14008,N_12706,N_13340);
or U14009 (N_14009,N_12326,N_12539);
or U14010 (N_14010,N_12949,N_12812);
or U14011 (N_14011,N_13160,N_13122);
or U14012 (N_14012,N_13083,N_12938);
nand U14013 (N_14013,N_12561,N_12239);
nor U14014 (N_14014,N_13365,N_12559);
and U14015 (N_14015,N_12164,N_12730);
nor U14016 (N_14016,N_12276,N_12448);
or U14017 (N_14017,N_13471,N_13464);
or U14018 (N_14018,N_13376,N_12870);
nor U14019 (N_14019,N_12055,N_12109);
or U14020 (N_14020,N_12430,N_12805);
or U14021 (N_14021,N_12102,N_13457);
or U14022 (N_14022,N_12907,N_12692);
nand U14023 (N_14023,N_12600,N_13088);
or U14024 (N_14024,N_12780,N_13086);
or U14025 (N_14025,N_12845,N_12678);
nor U14026 (N_14026,N_12028,N_13281);
and U14027 (N_14027,N_12602,N_12327);
and U14028 (N_14028,N_13246,N_13159);
or U14029 (N_14029,N_12264,N_13348);
nor U14030 (N_14030,N_13209,N_13106);
and U14031 (N_14031,N_12869,N_13025);
or U14032 (N_14032,N_12087,N_12645);
nor U14033 (N_14033,N_13318,N_12093);
nand U14034 (N_14034,N_12281,N_12926);
nand U14035 (N_14035,N_13001,N_12712);
xnor U14036 (N_14036,N_12753,N_12672);
or U14037 (N_14037,N_13398,N_12119);
and U14038 (N_14038,N_12997,N_13163);
nand U14039 (N_14039,N_12091,N_13366);
nor U14040 (N_14040,N_13189,N_12193);
nand U14041 (N_14041,N_13424,N_12424);
or U14042 (N_14042,N_12194,N_13394);
or U14043 (N_14043,N_12177,N_12295);
nand U14044 (N_14044,N_12542,N_12388);
xnor U14045 (N_14045,N_12820,N_13452);
xor U14046 (N_14046,N_12044,N_12670);
or U14047 (N_14047,N_12862,N_13066);
nor U14048 (N_14048,N_12804,N_13498);
nor U14049 (N_14049,N_13055,N_13476);
nor U14050 (N_14050,N_12429,N_12314);
xnor U14051 (N_14051,N_13494,N_12829);
and U14052 (N_14052,N_12759,N_13063);
and U14053 (N_14053,N_13283,N_13292);
and U14054 (N_14054,N_13241,N_13167);
nand U14055 (N_14055,N_12673,N_12232);
or U14056 (N_14056,N_12722,N_12942);
and U14057 (N_14057,N_12185,N_12100);
xnor U14058 (N_14058,N_12867,N_12815);
or U14059 (N_14059,N_13268,N_12364);
or U14060 (N_14060,N_12754,N_12463);
xnor U14061 (N_14061,N_12229,N_12366);
nand U14062 (N_14062,N_13346,N_12224);
xor U14063 (N_14063,N_13012,N_13067);
nor U14064 (N_14064,N_12794,N_12097);
nor U14065 (N_14065,N_12715,N_12648);
or U14066 (N_14066,N_12484,N_12173);
nand U14067 (N_14067,N_12787,N_12905);
or U14068 (N_14068,N_12995,N_12940);
xnor U14069 (N_14069,N_12860,N_12574);
or U14070 (N_14070,N_12476,N_13491);
and U14071 (N_14071,N_13448,N_12756);
and U14072 (N_14072,N_12328,N_13022);
and U14073 (N_14073,N_13465,N_13136);
xnor U14074 (N_14074,N_13126,N_13123);
nor U14075 (N_14075,N_13114,N_13455);
xnor U14076 (N_14076,N_12646,N_13438);
nor U14077 (N_14077,N_12767,N_12444);
nand U14078 (N_14078,N_13265,N_13461);
nor U14079 (N_14079,N_13478,N_12056);
or U14080 (N_14080,N_13047,N_13499);
or U14081 (N_14081,N_12757,N_13323);
nand U14082 (N_14082,N_12662,N_13426);
xor U14083 (N_14083,N_12181,N_12839);
and U14084 (N_14084,N_12861,N_13171);
xnor U14085 (N_14085,N_12075,N_13245);
nor U14086 (N_14086,N_12738,N_12151);
and U14087 (N_14087,N_12338,N_13411);
or U14088 (N_14088,N_13161,N_12803);
nor U14089 (N_14089,N_13124,N_12915);
nand U14090 (N_14090,N_13335,N_12473);
xnor U14091 (N_14091,N_12769,N_12874);
xor U14092 (N_14092,N_12158,N_12457);
nand U14093 (N_14093,N_12704,N_13195);
xor U14094 (N_14094,N_12530,N_12340);
and U14095 (N_14095,N_12633,N_12362);
nor U14096 (N_14096,N_13416,N_12161);
nand U14097 (N_14097,N_13206,N_12973);
nand U14098 (N_14098,N_13035,N_13304);
nor U14099 (N_14099,N_12968,N_12914);
xnor U14100 (N_14100,N_13250,N_12709);
or U14101 (N_14101,N_12140,N_12302);
nor U14102 (N_14102,N_12644,N_13187);
or U14103 (N_14103,N_13240,N_12428);
nor U14104 (N_14104,N_12609,N_12834);
nor U14105 (N_14105,N_12187,N_13011);
or U14106 (N_14106,N_13296,N_13430);
and U14107 (N_14107,N_13285,N_13350);
nor U14108 (N_14108,N_12061,N_13293);
or U14109 (N_14109,N_13015,N_12872);
xor U14110 (N_14110,N_12739,N_12434);
nor U14111 (N_14111,N_13070,N_12585);
and U14112 (N_14112,N_12642,N_12373);
xor U14113 (N_14113,N_12060,N_12752);
or U14114 (N_14114,N_12689,N_12453);
and U14115 (N_14115,N_13354,N_13218);
xnor U14116 (N_14116,N_12307,N_12369);
or U14117 (N_14117,N_13413,N_13496);
nand U14118 (N_14118,N_13432,N_12162);
xor U14119 (N_14119,N_12460,N_12495);
xnor U14120 (N_14120,N_12925,N_12433);
nor U14121 (N_14121,N_13389,N_12059);
and U14122 (N_14122,N_13361,N_13227);
xnor U14123 (N_14123,N_13270,N_13320);
or U14124 (N_14124,N_12083,N_12077);
or U14125 (N_14125,N_12582,N_13198);
and U14126 (N_14126,N_12607,N_12438);
or U14127 (N_14127,N_12990,N_12030);
and U14128 (N_14128,N_12216,N_12613);
nor U14129 (N_14129,N_12533,N_12982);
nand U14130 (N_14130,N_12213,N_13449);
or U14131 (N_14131,N_13157,N_12515);
xor U14132 (N_14132,N_12576,N_13031);
or U14133 (N_14133,N_13098,N_12935);
or U14134 (N_14134,N_13103,N_13488);
and U14135 (N_14135,N_12469,N_12980);
nand U14136 (N_14136,N_12864,N_13406);
nor U14137 (N_14137,N_13388,N_13279);
or U14138 (N_14138,N_12717,N_12024);
nor U14139 (N_14139,N_13387,N_13342);
xor U14140 (N_14140,N_12065,N_12365);
nand U14141 (N_14141,N_12235,N_12368);
and U14142 (N_14142,N_13030,N_13076);
nor U14143 (N_14143,N_12371,N_13094);
xnor U14144 (N_14144,N_12750,N_12965);
nand U14145 (N_14145,N_12621,N_12779);
nor U14146 (N_14146,N_13277,N_12758);
nand U14147 (N_14147,N_12939,N_12629);
xor U14148 (N_14148,N_13182,N_12534);
nand U14149 (N_14149,N_12458,N_13125);
and U14150 (N_14150,N_12891,N_13347);
and U14151 (N_14151,N_12126,N_13173);
nor U14152 (N_14152,N_12547,N_12772);
or U14153 (N_14153,N_12760,N_12836);
xor U14154 (N_14154,N_12540,N_12472);
or U14155 (N_14155,N_12240,N_13009);
nor U14156 (N_14156,N_12774,N_12505);
xnor U14157 (N_14157,N_12961,N_12455);
or U14158 (N_14158,N_12681,N_12111);
and U14159 (N_14159,N_13074,N_13294);
nand U14160 (N_14160,N_13097,N_13105);
and U14161 (N_14161,N_12594,N_12937);
xnor U14162 (N_14162,N_12147,N_12396);
or U14163 (N_14163,N_12818,N_12383);
nand U14164 (N_14164,N_12449,N_13272);
nor U14165 (N_14165,N_12846,N_13282);
nand U14166 (N_14166,N_13301,N_13403);
and U14167 (N_14167,N_12431,N_12349);
and U14168 (N_14168,N_13477,N_12475);
and U14169 (N_14169,N_13154,N_12952);
and U14170 (N_14170,N_13131,N_12020);
nand U14171 (N_14171,N_12498,N_12510);
or U14172 (N_14172,N_12636,N_12790);
xnor U14173 (N_14173,N_13351,N_12105);
or U14174 (N_14174,N_12133,N_12865);
nor U14175 (N_14175,N_12998,N_13429);
nor U14176 (N_14176,N_12577,N_13375);
and U14177 (N_14177,N_12486,N_13216);
nand U14178 (N_14178,N_13329,N_12136);
xor U14179 (N_14179,N_12929,N_12132);
nor U14180 (N_14180,N_12904,N_12748);
nor U14181 (N_14181,N_12411,N_12490);
or U14182 (N_14182,N_12210,N_13166);
and U14183 (N_14183,N_12674,N_12676);
or U14184 (N_14184,N_12897,N_13480);
xor U14185 (N_14185,N_12299,N_12446);
nor U14186 (N_14186,N_12966,N_12881);
nor U14187 (N_14187,N_12596,N_12401);
or U14188 (N_14188,N_12509,N_12012);
and U14189 (N_14189,N_13085,N_12211);
nor U14190 (N_14190,N_13032,N_12930);
nand U14191 (N_14191,N_12425,N_13297);
xor U14192 (N_14192,N_13181,N_13442);
or U14193 (N_14193,N_12226,N_13404);
and U14194 (N_14194,N_12630,N_12923);
xnor U14195 (N_14195,N_13078,N_12902);
nor U14196 (N_14196,N_12031,N_12051);
nor U14197 (N_14197,N_13439,N_12333);
nand U14198 (N_14198,N_12632,N_12729);
nor U14199 (N_14199,N_12611,N_12286);
or U14200 (N_14200,N_12592,N_13152);
or U14201 (N_14201,N_12114,N_12634);
nand U14202 (N_14202,N_12023,N_12415);
nor U14203 (N_14203,N_13357,N_12983);
nand U14204 (N_14204,N_13048,N_12394);
nor U14205 (N_14205,N_13443,N_12182);
nor U14206 (N_14206,N_13287,N_12403);
nand U14207 (N_14207,N_12853,N_12395);
and U14208 (N_14208,N_13267,N_12858);
or U14209 (N_14209,N_12492,N_12919);
nand U14210 (N_14210,N_12608,N_13132);
nor U14211 (N_14211,N_12801,N_13200);
xnor U14212 (N_14212,N_12311,N_13421);
nor U14213 (N_14213,N_12377,N_12762);
nor U14214 (N_14214,N_12742,N_12078);
and U14215 (N_14215,N_12763,N_13053);
or U14216 (N_14216,N_12293,N_13417);
nor U14217 (N_14217,N_13059,N_12296);
nor U14218 (N_14218,N_13236,N_13164);
nand U14219 (N_14219,N_13115,N_12215);
and U14220 (N_14220,N_12536,N_12137);
nor U14221 (N_14221,N_12851,N_13409);
nor U14222 (N_14222,N_12149,N_12249);
nor U14223 (N_14223,N_12374,N_12657);
xnor U14224 (N_14224,N_12500,N_12837);
and U14225 (N_14225,N_12734,N_12587);
or U14226 (N_14226,N_12272,N_12027);
nor U14227 (N_14227,N_12104,N_13400);
nand U14228 (N_14228,N_12204,N_13234);
nor U14229 (N_14229,N_12797,N_12095);
nor U14230 (N_14230,N_12811,N_12589);
xor U14231 (N_14231,N_12178,N_12551);
nor U14232 (N_14232,N_13062,N_12402);
nor U14233 (N_14233,N_13317,N_12685);
nor U14234 (N_14234,N_12466,N_13379);
nor U14235 (N_14235,N_12654,N_12222);
xnor U14236 (N_14236,N_13369,N_12350);
or U14237 (N_14237,N_12620,N_13026);
and U14238 (N_14238,N_13321,N_12720);
and U14239 (N_14239,N_13174,N_12035);
nand U14240 (N_14240,N_13450,N_12319);
or U14241 (N_14241,N_13306,N_12518);
xor U14242 (N_14242,N_12984,N_13341);
nand U14243 (N_14243,N_12733,N_12626);
xor U14244 (N_14244,N_12123,N_13475);
or U14245 (N_14245,N_12166,N_13111);
or U14246 (N_14246,N_12778,N_12789);
nand U14247 (N_14247,N_12157,N_12043);
or U14248 (N_14248,N_12467,N_12205);
and U14249 (N_14249,N_13140,N_12280);
xor U14250 (N_14250,N_12299,N_12520);
xnor U14251 (N_14251,N_12102,N_13142);
xor U14252 (N_14252,N_12741,N_12313);
nor U14253 (N_14253,N_12119,N_13105);
nor U14254 (N_14254,N_12997,N_13195);
nor U14255 (N_14255,N_12937,N_13375);
xnor U14256 (N_14256,N_13461,N_12924);
xnor U14257 (N_14257,N_12721,N_12257);
and U14258 (N_14258,N_13148,N_12458);
or U14259 (N_14259,N_12431,N_13256);
nor U14260 (N_14260,N_13195,N_12667);
xnor U14261 (N_14261,N_13490,N_12599);
and U14262 (N_14262,N_12053,N_13403);
xnor U14263 (N_14263,N_12349,N_13054);
nand U14264 (N_14264,N_12618,N_13370);
xor U14265 (N_14265,N_13379,N_13480);
nand U14266 (N_14266,N_12050,N_12399);
or U14267 (N_14267,N_13365,N_12534);
and U14268 (N_14268,N_12793,N_12183);
nand U14269 (N_14269,N_12611,N_13272);
xor U14270 (N_14270,N_13260,N_13474);
and U14271 (N_14271,N_13341,N_13226);
nand U14272 (N_14272,N_12798,N_13042);
and U14273 (N_14273,N_12724,N_12128);
or U14274 (N_14274,N_12721,N_12627);
nand U14275 (N_14275,N_13106,N_13240);
or U14276 (N_14276,N_12922,N_12712);
nor U14277 (N_14277,N_12944,N_12421);
nor U14278 (N_14278,N_12605,N_13021);
xnor U14279 (N_14279,N_13454,N_12641);
nor U14280 (N_14280,N_12360,N_13151);
nor U14281 (N_14281,N_13498,N_12204);
nand U14282 (N_14282,N_12543,N_12288);
nand U14283 (N_14283,N_12919,N_13020);
nand U14284 (N_14284,N_13211,N_13355);
nand U14285 (N_14285,N_12958,N_12309);
nand U14286 (N_14286,N_12978,N_12002);
and U14287 (N_14287,N_13271,N_12854);
nand U14288 (N_14288,N_12914,N_12008);
nor U14289 (N_14289,N_13010,N_12401);
xor U14290 (N_14290,N_12209,N_12204);
nand U14291 (N_14291,N_13412,N_12304);
nand U14292 (N_14292,N_12830,N_13422);
nor U14293 (N_14293,N_13221,N_12278);
nand U14294 (N_14294,N_13232,N_12411);
nor U14295 (N_14295,N_13459,N_12307);
nor U14296 (N_14296,N_12786,N_13040);
xor U14297 (N_14297,N_13315,N_12059);
and U14298 (N_14298,N_12796,N_12311);
nand U14299 (N_14299,N_13085,N_12809);
and U14300 (N_14300,N_12933,N_13135);
nand U14301 (N_14301,N_12087,N_13185);
or U14302 (N_14302,N_12594,N_12373);
xor U14303 (N_14303,N_12612,N_12861);
nor U14304 (N_14304,N_13495,N_13355);
and U14305 (N_14305,N_12583,N_12968);
xor U14306 (N_14306,N_13199,N_12207);
and U14307 (N_14307,N_13436,N_12411);
nand U14308 (N_14308,N_13495,N_12964);
nand U14309 (N_14309,N_13389,N_12568);
or U14310 (N_14310,N_12142,N_13483);
nand U14311 (N_14311,N_12052,N_13281);
nand U14312 (N_14312,N_12643,N_12497);
nand U14313 (N_14313,N_12489,N_13335);
xor U14314 (N_14314,N_13094,N_12569);
xnor U14315 (N_14315,N_12571,N_12848);
nor U14316 (N_14316,N_12780,N_12737);
nor U14317 (N_14317,N_13056,N_12282);
nand U14318 (N_14318,N_13350,N_12763);
xnor U14319 (N_14319,N_12990,N_13061);
and U14320 (N_14320,N_12465,N_12234);
or U14321 (N_14321,N_13046,N_13068);
and U14322 (N_14322,N_12380,N_12909);
nor U14323 (N_14323,N_12168,N_12133);
or U14324 (N_14324,N_12022,N_13474);
or U14325 (N_14325,N_13453,N_12641);
and U14326 (N_14326,N_12582,N_12376);
and U14327 (N_14327,N_12223,N_12081);
xnor U14328 (N_14328,N_13384,N_12820);
nor U14329 (N_14329,N_13128,N_13111);
nor U14330 (N_14330,N_12684,N_12137);
or U14331 (N_14331,N_12154,N_12079);
and U14332 (N_14332,N_13253,N_13301);
nand U14333 (N_14333,N_12424,N_13189);
or U14334 (N_14334,N_12858,N_12934);
xor U14335 (N_14335,N_12097,N_12953);
or U14336 (N_14336,N_12057,N_12794);
nand U14337 (N_14337,N_12430,N_12515);
and U14338 (N_14338,N_13451,N_13142);
nand U14339 (N_14339,N_13120,N_13157);
or U14340 (N_14340,N_12531,N_13278);
and U14341 (N_14341,N_12577,N_13459);
xnor U14342 (N_14342,N_12074,N_12175);
or U14343 (N_14343,N_12415,N_12743);
or U14344 (N_14344,N_12172,N_12565);
nor U14345 (N_14345,N_12493,N_13287);
nand U14346 (N_14346,N_12007,N_12215);
xor U14347 (N_14347,N_12997,N_13452);
and U14348 (N_14348,N_13433,N_13431);
and U14349 (N_14349,N_12859,N_13407);
or U14350 (N_14350,N_12144,N_12314);
or U14351 (N_14351,N_12760,N_12301);
or U14352 (N_14352,N_12781,N_12911);
xor U14353 (N_14353,N_12030,N_12459);
or U14354 (N_14354,N_13213,N_12940);
nand U14355 (N_14355,N_12240,N_12144);
and U14356 (N_14356,N_12216,N_12990);
and U14357 (N_14357,N_12168,N_13080);
and U14358 (N_14358,N_13476,N_13430);
and U14359 (N_14359,N_13443,N_12139);
xnor U14360 (N_14360,N_13481,N_13489);
and U14361 (N_14361,N_12738,N_13077);
nand U14362 (N_14362,N_12595,N_13287);
nor U14363 (N_14363,N_13221,N_12506);
or U14364 (N_14364,N_13197,N_12505);
xnor U14365 (N_14365,N_12048,N_12194);
nand U14366 (N_14366,N_12720,N_13249);
and U14367 (N_14367,N_13416,N_12128);
or U14368 (N_14368,N_12674,N_13128);
nor U14369 (N_14369,N_13465,N_12164);
nor U14370 (N_14370,N_12897,N_13371);
nor U14371 (N_14371,N_12117,N_12222);
nand U14372 (N_14372,N_12424,N_12113);
and U14373 (N_14373,N_13214,N_12524);
nor U14374 (N_14374,N_13377,N_13051);
and U14375 (N_14375,N_12416,N_13488);
xnor U14376 (N_14376,N_13028,N_12732);
xnor U14377 (N_14377,N_12811,N_13402);
or U14378 (N_14378,N_12629,N_12274);
and U14379 (N_14379,N_13258,N_13238);
nand U14380 (N_14380,N_12040,N_13215);
xnor U14381 (N_14381,N_13227,N_12165);
or U14382 (N_14382,N_12799,N_12873);
nor U14383 (N_14383,N_12839,N_13103);
and U14384 (N_14384,N_12949,N_12684);
nand U14385 (N_14385,N_12824,N_12499);
nor U14386 (N_14386,N_12821,N_12603);
xor U14387 (N_14387,N_12734,N_12486);
nand U14388 (N_14388,N_13381,N_12958);
nand U14389 (N_14389,N_12274,N_12440);
nor U14390 (N_14390,N_12510,N_12033);
nor U14391 (N_14391,N_12224,N_12992);
xor U14392 (N_14392,N_13050,N_13405);
or U14393 (N_14393,N_13229,N_12554);
nand U14394 (N_14394,N_12892,N_12540);
nor U14395 (N_14395,N_12711,N_13159);
nor U14396 (N_14396,N_12257,N_12861);
and U14397 (N_14397,N_13183,N_12684);
or U14398 (N_14398,N_13227,N_13116);
nor U14399 (N_14399,N_12316,N_13417);
or U14400 (N_14400,N_13443,N_12515);
or U14401 (N_14401,N_12546,N_13281);
nor U14402 (N_14402,N_13030,N_12484);
nor U14403 (N_14403,N_13100,N_12013);
xor U14404 (N_14404,N_12656,N_12845);
xor U14405 (N_14405,N_12726,N_13067);
and U14406 (N_14406,N_13230,N_12098);
or U14407 (N_14407,N_13178,N_12862);
xor U14408 (N_14408,N_13492,N_12341);
xor U14409 (N_14409,N_12524,N_13203);
and U14410 (N_14410,N_13030,N_12426);
nor U14411 (N_14411,N_13033,N_12189);
nor U14412 (N_14412,N_13022,N_12318);
and U14413 (N_14413,N_13472,N_13168);
nor U14414 (N_14414,N_12678,N_13170);
or U14415 (N_14415,N_12417,N_12223);
nor U14416 (N_14416,N_12799,N_12649);
nor U14417 (N_14417,N_12991,N_13116);
xor U14418 (N_14418,N_13254,N_13045);
xor U14419 (N_14419,N_12362,N_12015);
nor U14420 (N_14420,N_12835,N_13309);
nand U14421 (N_14421,N_13213,N_12451);
xnor U14422 (N_14422,N_13411,N_12961);
and U14423 (N_14423,N_13366,N_12683);
nand U14424 (N_14424,N_12761,N_12128);
xnor U14425 (N_14425,N_12852,N_12599);
xnor U14426 (N_14426,N_13050,N_12072);
nor U14427 (N_14427,N_13454,N_12657);
nand U14428 (N_14428,N_13252,N_13005);
xnor U14429 (N_14429,N_13322,N_13361);
nand U14430 (N_14430,N_12250,N_12350);
nand U14431 (N_14431,N_12074,N_12000);
nor U14432 (N_14432,N_12370,N_13307);
or U14433 (N_14433,N_13131,N_12937);
nand U14434 (N_14434,N_12382,N_13371);
nand U14435 (N_14435,N_12801,N_13311);
nor U14436 (N_14436,N_12165,N_12495);
and U14437 (N_14437,N_13028,N_12709);
and U14438 (N_14438,N_12754,N_12242);
or U14439 (N_14439,N_12417,N_12359);
nand U14440 (N_14440,N_12656,N_12226);
xor U14441 (N_14441,N_13004,N_12018);
nor U14442 (N_14442,N_12430,N_12645);
nand U14443 (N_14443,N_12775,N_13425);
or U14444 (N_14444,N_13037,N_12664);
and U14445 (N_14445,N_13259,N_13214);
nand U14446 (N_14446,N_12587,N_12544);
xnor U14447 (N_14447,N_13126,N_12394);
and U14448 (N_14448,N_12187,N_12373);
or U14449 (N_14449,N_12391,N_13115);
xnor U14450 (N_14450,N_12042,N_12846);
xor U14451 (N_14451,N_12599,N_12992);
nand U14452 (N_14452,N_12980,N_13344);
and U14453 (N_14453,N_12133,N_13237);
and U14454 (N_14454,N_12807,N_12166);
or U14455 (N_14455,N_12587,N_13106);
xnor U14456 (N_14456,N_13388,N_12265);
nor U14457 (N_14457,N_13253,N_12772);
nor U14458 (N_14458,N_12887,N_13064);
or U14459 (N_14459,N_13368,N_12686);
or U14460 (N_14460,N_13486,N_12613);
and U14461 (N_14461,N_12669,N_12124);
nor U14462 (N_14462,N_12822,N_13420);
nor U14463 (N_14463,N_12900,N_12446);
xor U14464 (N_14464,N_12715,N_12110);
xor U14465 (N_14465,N_13346,N_13215);
and U14466 (N_14466,N_13358,N_12020);
and U14467 (N_14467,N_13023,N_12898);
or U14468 (N_14468,N_12740,N_12755);
and U14469 (N_14469,N_12309,N_12770);
or U14470 (N_14470,N_12432,N_12545);
and U14471 (N_14471,N_13446,N_12636);
xnor U14472 (N_14472,N_12978,N_12728);
xnor U14473 (N_14473,N_12634,N_12100);
or U14474 (N_14474,N_13054,N_13200);
nor U14475 (N_14475,N_12459,N_12412);
and U14476 (N_14476,N_13185,N_12724);
xor U14477 (N_14477,N_12761,N_12376);
nand U14478 (N_14478,N_12375,N_12139);
xnor U14479 (N_14479,N_12151,N_12306);
xor U14480 (N_14480,N_13340,N_12198);
or U14481 (N_14481,N_12159,N_13378);
nor U14482 (N_14482,N_12437,N_12523);
nand U14483 (N_14483,N_12163,N_12555);
and U14484 (N_14484,N_13106,N_12832);
nor U14485 (N_14485,N_13250,N_12653);
nand U14486 (N_14486,N_13422,N_12413);
or U14487 (N_14487,N_12685,N_13129);
or U14488 (N_14488,N_12849,N_12493);
nand U14489 (N_14489,N_12662,N_12846);
xnor U14490 (N_14490,N_13352,N_13398);
or U14491 (N_14491,N_12338,N_12987);
or U14492 (N_14492,N_12068,N_13363);
nor U14493 (N_14493,N_12278,N_12186);
xor U14494 (N_14494,N_12700,N_13294);
xor U14495 (N_14495,N_12005,N_12202);
or U14496 (N_14496,N_13311,N_12079);
nor U14497 (N_14497,N_13483,N_12634);
nand U14498 (N_14498,N_13391,N_12889);
nand U14499 (N_14499,N_13038,N_12377);
and U14500 (N_14500,N_12155,N_12975);
nor U14501 (N_14501,N_13093,N_12127);
nor U14502 (N_14502,N_12611,N_12182);
nor U14503 (N_14503,N_13090,N_13412);
and U14504 (N_14504,N_12558,N_12623);
xnor U14505 (N_14505,N_12169,N_13026);
nor U14506 (N_14506,N_12329,N_12796);
nand U14507 (N_14507,N_12889,N_12272);
or U14508 (N_14508,N_12185,N_13085);
or U14509 (N_14509,N_13024,N_13128);
xnor U14510 (N_14510,N_12182,N_12050);
nand U14511 (N_14511,N_13462,N_12921);
xor U14512 (N_14512,N_13181,N_13166);
xor U14513 (N_14513,N_12564,N_13487);
nor U14514 (N_14514,N_12871,N_12194);
xor U14515 (N_14515,N_12845,N_13341);
nor U14516 (N_14516,N_13392,N_12763);
and U14517 (N_14517,N_12913,N_12244);
xor U14518 (N_14518,N_12559,N_12339);
or U14519 (N_14519,N_13169,N_12564);
or U14520 (N_14520,N_12654,N_12954);
nand U14521 (N_14521,N_12656,N_12216);
and U14522 (N_14522,N_12311,N_12920);
and U14523 (N_14523,N_13251,N_12245);
or U14524 (N_14524,N_13170,N_13013);
and U14525 (N_14525,N_12068,N_13242);
nor U14526 (N_14526,N_13416,N_12379);
nand U14527 (N_14527,N_13218,N_12210);
or U14528 (N_14528,N_12021,N_13432);
xnor U14529 (N_14529,N_12449,N_12590);
nor U14530 (N_14530,N_13033,N_13303);
and U14531 (N_14531,N_12838,N_13072);
nand U14532 (N_14532,N_12720,N_12395);
and U14533 (N_14533,N_12965,N_13277);
nor U14534 (N_14534,N_12135,N_13474);
and U14535 (N_14535,N_12100,N_12838);
nor U14536 (N_14536,N_12715,N_12807);
nor U14537 (N_14537,N_12622,N_13394);
xor U14538 (N_14538,N_13364,N_12082);
nor U14539 (N_14539,N_12926,N_12399);
or U14540 (N_14540,N_12789,N_13037);
nor U14541 (N_14541,N_12597,N_12429);
and U14542 (N_14542,N_12951,N_13447);
or U14543 (N_14543,N_13232,N_12509);
and U14544 (N_14544,N_13422,N_12114);
or U14545 (N_14545,N_12287,N_12353);
or U14546 (N_14546,N_12896,N_12542);
and U14547 (N_14547,N_12452,N_12698);
nand U14548 (N_14548,N_12173,N_13059);
xor U14549 (N_14549,N_13120,N_13085);
xnor U14550 (N_14550,N_13382,N_13056);
or U14551 (N_14551,N_13457,N_13317);
nor U14552 (N_14552,N_13302,N_12589);
or U14553 (N_14553,N_12330,N_12542);
xor U14554 (N_14554,N_13057,N_12354);
nand U14555 (N_14555,N_12935,N_13134);
and U14556 (N_14556,N_12737,N_13120);
xor U14557 (N_14557,N_12222,N_13058);
nor U14558 (N_14558,N_12513,N_12181);
xor U14559 (N_14559,N_12604,N_12665);
nand U14560 (N_14560,N_13405,N_13495);
xor U14561 (N_14561,N_12774,N_12367);
xor U14562 (N_14562,N_12312,N_12552);
and U14563 (N_14563,N_13055,N_13182);
xor U14564 (N_14564,N_12346,N_12252);
or U14565 (N_14565,N_12136,N_12981);
nand U14566 (N_14566,N_12086,N_13298);
nand U14567 (N_14567,N_12560,N_12344);
xnor U14568 (N_14568,N_12512,N_12555);
nor U14569 (N_14569,N_13169,N_12113);
and U14570 (N_14570,N_13234,N_13203);
nor U14571 (N_14571,N_12035,N_13448);
nand U14572 (N_14572,N_12944,N_13305);
and U14573 (N_14573,N_12761,N_13154);
xnor U14574 (N_14574,N_12809,N_12484);
and U14575 (N_14575,N_13041,N_13315);
nor U14576 (N_14576,N_12603,N_12392);
nand U14577 (N_14577,N_12505,N_12199);
nand U14578 (N_14578,N_13043,N_12340);
or U14579 (N_14579,N_12296,N_12080);
and U14580 (N_14580,N_12877,N_12073);
nor U14581 (N_14581,N_12356,N_12213);
xnor U14582 (N_14582,N_13341,N_13324);
and U14583 (N_14583,N_12902,N_12420);
or U14584 (N_14584,N_12967,N_12794);
or U14585 (N_14585,N_12138,N_12933);
nand U14586 (N_14586,N_12042,N_12621);
xor U14587 (N_14587,N_12724,N_12841);
and U14588 (N_14588,N_12696,N_12811);
nor U14589 (N_14589,N_12668,N_13267);
or U14590 (N_14590,N_12364,N_12074);
nand U14591 (N_14591,N_12717,N_12971);
and U14592 (N_14592,N_13018,N_12968);
and U14593 (N_14593,N_12445,N_12604);
xnor U14594 (N_14594,N_13112,N_12184);
xor U14595 (N_14595,N_12053,N_12608);
xor U14596 (N_14596,N_12291,N_12414);
nand U14597 (N_14597,N_12075,N_12511);
and U14598 (N_14598,N_12332,N_12526);
or U14599 (N_14599,N_13386,N_13313);
and U14600 (N_14600,N_12363,N_12210);
or U14601 (N_14601,N_12087,N_12545);
nor U14602 (N_14602,N_12516,N_12003);
nand U14603 (N_14603,N_12100,N_12549);
xnor U14604 (N_14604,N_12167,N_13311);
nand U14605 (N_14605,N_12640,N_13105);
or U14606 (N_14606,N_12867,N_12464);
nor U14607 (N_14607,N_12836,N_12925);
nor U14608 (N_14608,N_12545,N_13103);
or U14609 (N_14609,N_12285,N_13460);
xnor U14610 (N_14610,N_13412,N_13037);
or U14611 (N_14611,N_12140,N_12162);
nand U14612 (N_14612,N_12769,N_12812);
xnor U14613 (N_14613,N_13054,N_12972);
and U14614 (N_14614,N_13446,N_12621);
nand U14615 (N_14615,N_12776,N_12407);
nand U14616 (N_14616,N_12771,N_12841);
nand U14617 (N_14617,N_12065,N_12886);
nand U14618 (N_14618,N_13035,N_12625);
or U14619 (N_14619,N_12565,N_13111);
and U14620 (N_14620,N_12402,N_13007);
and U14621 (N_14621,N_12788,N_12941);
xor U14622 (N_14622,N_12909,N_12135);
nand U14623 (N_14623,N_12704,N_12886);
xor U14624 (N_14624,N_12915,N_13088);
nor U14625 (N_14625,N_12767,N_13202);
and U14626 (N_14626,N_13128,N_12238);
xnor U14627 (N_14627,N_13477,N_12876);
xor U14628 (N_14628,N_12695,N_12864);
or U14629 (N_14629,N_13107,N_12292);
or U14630 (N_14630,N_12598,N_13134);
nand U14631 (N_14631,N_12900,N_12667);
or U14632 (N_14632,N_12006,N_12488);
nor U14633 (N_14633,N_13028,N_12185);
nand U14634 (N_14634,N_12555,N_12126);
and U14635 (N_14635,N_12763,N_12968);
nand U14636 (N_14636,N_12227,N_13335);
nand U14637 (N_14637,N_12956,N_12567);
nand U14638 (N_14638,N_12255,N_12191);
nor U14639 (N_14639,N_13333,N_12498);
xor U14640 (N_14640,N_13119,N_12087);
or U14641 (N_14641,N_12859,N_12710);
xor U14642 (N_14642,N_12866,N_12993);
nand U14643 (N_14643,N_12261,N_12173);
and U14644 (N_14644,N_13345,N_12765);
nor U14645 (N_14645,N_13003,N_12670);
or U14646 (N_14646,N_12105,N_13416);
or U14647 (N_14647,N_13068,N_12268);
and U14648 (N_14648,N_12392,N_12080);
nor U14649 (N_14649,N_13292,N_12922);
and U14650 (N_14650,N_12638,N_12789);
nor U14651 (N_14651,N_13400,N_12912);
and U14652 (N_14652,N_13090,N_13261);
xnor U14653 (N_14653,N_13463,N_12417);
or U14654 (N_14654,N_12452,N_12279);
and U14655 (N_14655,N_13306,N_13065);
nor U14656 (N_14656,N_13380,N_13080);
xnor U14657 (N_14657,N_12565,N_12757);
or U14658 (N_14658,N_13313,N_13202);
or U14659 (N_14659,N_13421,N_13122);
xnor U14660 (N_14660,N_12835,N_12093);
or U14661 (N_14661,N_13375,N_12524);
nand U14662 (N_14662,N_12060,N_12986);
and U14663 (N_14663,N_13479,N_13030);
and U14664 (N_14664,N_13148,N_13016);
nand U14665 (N_14665,N_12392,N_12361);
xnor U14666 (N_14666,N_12836,N_12645);
nor U14667 (N_14667,N_12146,N_12912);
and U14668 (N_14668,N_12402,N_12271);
nand U14669 (N_14669,N_12178,N_12646);
xnor U14670 (N_14670,N_13403,N_12291);
xor U14671 (N_14671,N_12505,N_13452);
nand U14672 (N_14672,N_12082,N_12418);
xor U14673 (N_14673,N_12063,N_13223);
nand U14674 (N_14674,N_12314,N_12394);
xor U14675 (N_14675,N_12031,N_12062);
nor U14676 (N_14676,N_12449,N_13053);
and U14677 (N_14677,N_13213,N_13195);
nor U14678 (N_14678,N_12432,N_12539);
and U14679 (N_14679,N_12809,N_12504);
or U14680 (N_14680,N_12548,N_13305);
nand U14681 (N_14681,N_12470,N_12225);
or U14682 (N_14682,N_13352,N_12491);
nand U14683 (N_14683,N_12409,N_12547);
and U14684 (N_14684,N_12653,N_13141);
and U14685 (N_14685,N_12098,N_12481);
nor U14686 (N_14686,N_13159,N_13187);
nor U14687 (N_14687,N_13277,N_12983);
xor U14688 (N_14688,N_13040,N_13327);
nand U14689 (N_14689,N_13171,N_12125);
and U14690 (N_14690,N_13047,N_13251);
nand U14691 (N_14691,N_13094,N_12937);
nor U14692 (N_14692,N_13493,N_13474);
xnor U14693 (N_14693,N_12300,N_12825);
nor U14694 (N_14694,N_13095,N_13492);
xor U14695 (N_14695,N_12796,N_13107);
xnor U14696 (N_14696,N_13144,N_12174);
xnor U14697 (N_14697,N_12848,N_13031);
xor U14698 (N_14698,N_12124,N_12214);
and U14699 (N_14699,N_12433,N_12816);
and U14700 (N_14700,N_13037,N_12823);
or U14701 (N_14701,N_12999,N_12873);
nor U14702 (N_14702,N_12189,N_13105);
xnor U14703 (N_14703,N_13438,N_12278);
xnor U14704 (N_14704,N_13084,N_13287);
or U14705 (N_14705,N_13132,N_12111);
or U14706 (N_14706,N_13011,N_13138);
nor U14707 (N_14707,N_12302,N_13079);
or U14708 (N_14708,N_12470,N_13112);
nand U14709 (N_14709,N_12418,N_12732);
nor U14710 (N_14710,N_13371,N_12052);
and U14711 (N_14711,N_12117,N_12158);
nor U14712 (N_14712,N_13472,N_12285);
nand U14713 (N_14713,N_12579,N_12849);
or U14714 (N_14714,N_12671,N_12300);
or U14715 (N_14715,N_12730,N_12017);
nand U14716 (N_14716,N_12066,N_12462);
and U14717 (N_14717,N_12776,N_12331);
and U14718 (N_14718,N_13339,N_12946);
or U14719 (N_14719,N_12805,N_13413);
nand U14720 (N_14720,N_13379,N_12000);
nor U14721 (N_14721,N_12658,N_13142);
nand U14722 (N_14722,N_12604,N_12816);
nand U14723 (N_14723,N_12821,N_12809);
or U14724 (N_14724,N_12671,N_13011);
xor U14725 (N_14725,N_12867,N_12857);
xnor U14726 (N_14726,N_12791,N_13346);
and U14727 (N_14727,N_12341,N_12103);
nor U14728 (N_14728,N_12682,N_12257);
nor U14729 (N_14729,N_12915,N_12080);
nor U14730 (N_14730,N_13329,N_12467);
or U14731 (N_14731,N_12696,N_12599);
and U14732 (N_14732,N_13429,N_13148);
nor U14733 (N_14733,N_12162,N_13400);
xor U14734 (N_14734,N_12867,N_12729);
xor U14735 (N_14735,N_12749,N_12342);
and U14736 (N_14736,N_13419,N_13160);
xnor U14737 (N_14737,N_12773,N_13250);
and U14738 (N_14738,N_12217,N_12103);
nor U14739 (N_14739,N_12783,N_12216);
nand U14740 (N_14740,N_12424,N_12306);
or U14741 (N_14741,N_12876,N_12172);
xor U14742 (N_14742,N_13237,N_13463);
nand U14743 (N_14743,N_12576,N_13170);
xor U14744 (N_14744,N_12525,N_12556);
xnor U14745 (N_14745,N_12407,N_12456);
nor U14746 (N_14746,N_12798,N_12799);
and U14747 (N_14747,N_13260,N_13039);
and U14748 (N_14748,N_12672,N_12060);
nor U14749 (N_14749,N_12268,N_12169);
nand U14750 (N_14750,N_13444,N_13018);
and U14751 (N_14751,N_12198,N_12654);
or U14752 (N_14752,N_12851,N_12161);
and U14753 (N_14753,N_12583,N_13224);
nor U14754 (N_14754,N_12228,N_13474);
nand U14755 (N_14755,N_13485,N_13324);
nand U14756 (N_14756,N_13198,N_12349);
nor U14757 (N_14757,N_13423,N_13467);
xor U14758 (N_14758,N_12532,N_12939);
xor U14759 (N_14759,N_12101,N_13370);
or U14760 (N_14760,N_12818,N_12640);
nor U14761 (N_14761,N_13099,N_12153);
nand U14762 (N_14762,N_12935,N_13193);
nand U14763 (N_14763,N_13326,N_12805);
nand U14764 (N_14764,N_13083,N_12196);
and U14765 (N_14765,N_13132,N_12777);
nor U14766 (N_14766,N_12390,N_12516);
nand U14767 (N_14767,N_12596,N_13314);
nand U14768 (N_14768,N_12418,N_13145);
nor U14769 (N_14769,N_13014,N_12306);
nor U14770 (N_14770,N_12519,N_12753);
nand U14771 (N_14771,N_12183,N_12947);
nor U14772 (N_14772,N_12550,N_12324);
nand U14773 (N_14773,N_12199,N_12240);
nor U14774 (N_14774,N_12519,N_13380);
nor U14775 (N_14775,N_12319,N_13184);
nor U14776 (N_14776,N_13270,N_12551);
xor U14777 (N_14777,N_12899,N_12752);
or U14778 (N_14778,N_12638,N_12870);
and U14779 (N_14779,N_12470,N_12786);
or U14780 (N_14780,N_13376,N_13286);
and U14781 (N_14781,N_12841,N_13416);
nor U14782 (N_14782,N_12094,N_12271);
xor U14783 (N_14783,N_12440,N_12627);
nand U14784 (N_14784,N_13287,N_12712);
xnor U14785 (N_14785,N_12553,N_12607);
or U14786 (N_14786,N_12809,N_12813);
or U14787 (N_14787,N_13399,N_12208);
or U14788 (N_14788,N_13253,N_12449);
nand U14789 (N_14789,N_13379,N_13132);
or U14790 (N_14790,N_13398,N_13350);
and U14791 (N_14791,N_13223,N_12306);
nand U14792 (N_14792,N_12769,N_12495);
nor U14793 (N_14793,N_12261,N_12986);
and U14794 (N_14794,N_13233,N_13383);
nand U14795 (N_14795,N_12149,N_12355);
nand U14796 (N_14796,N_12725,N_13069);
or U14797 (N_14797,N_12805,N_12675);
nor U14798 (N_14798,N_12157,N_12512);
nand U14799 (N_14799,N_13065,N_12787);
xor U14800 (N_14800,N_12623,N_12648);
nand U14801 (N_14801,N_12125,N_12078);
xor U14802 (N_14802,N_12349,N_12256);
xnor U14803 (N_14803,N_12610,N_12627);
or U14804 (N_14804,N_13246,N_13152);
nand U14805 (N_14805,N_12464,N_13454);
xnor U14806 (N_14806,N_13122,N_12835);
nor U14807 (N_14807,N_13275,N_12449);
xnor U14808 (N_14808,N_12079,N_12896);
and U14809 (N_14809,N_12105,N_12915);
and U14810 (N_14810,N_12027,N_12267);
nand U14811 (N_14811,N_13291,N_12920);
nand U14812 (N_14812,N_12313,N_13428);
nand U14813 (N_14813,N_13413,N_12884);
and U14814 (N_14814,N_12831,N_13494);
or U14815 (N_14815,N_12979,N_12299);
or U14816 (N_14816,N_13373,N_13183);
and U14817 (N_14817,N_13050,N_12025);
xor U14818 (N_14818,N_12728,N_12369);
nand U14819 (N_14819,N_13088,N_12476);
and U14820 (N_14820,N_12010,N_13255);
xnor U14821 (N_14821,N_12832,N_12355);
xor U14822 (N_14822,N_12218,N_13266);
nand U14823 (N_14823,N_12300,N_12413);
xnor U14824 (N_14824,N_12969,N_13468);
and U14825 (N_14825,N_12441,N_12564);
nand U14826 (N_14826,N_13385,N_12342);
nor U14827 (N_14827,N_12531,N_13499);
or U14828 (N_14828,N_12206,N_12522);
xnor U14829 (N_14829,N_13391,N_12934);
or U14830 (N_14830,N_13245,N_12411);
and U14831 (N_14831,N_12687,N_12908);
or U14832 (N_14832,N_13296,N_12396);
nand U14833 (N_14833,N_13364,N_12146);
xor U14834 (N_14834,N_12548,N_12459);
nor U14835 (N_14835,N_12796,N_12290);
and U14836 (N_14836,N_12317,N_12702);
nor U14837 (N_14837,N_13258,N_12968);
and U14838 (N_14838,N_12425,N_12752);
xnor U14839 (N_14839,N_12691,N_12829);
nand U14840 (N_14840,N_12044,N_12326);
nor U14841 (N_14841,N_12572,N_12061);
nand U14842 (N_14842,N_12696,N_12719);
nand U14843 (N_14843,N_12736,N_13354);
nor U14844 (N_14844,N_12504,N_13154);
nor U14845 (N_14845,N_12204,N_13185);
or U14846 (N_14846,N_12184,N_12404);
or U14847 (N_14847,N_13265,N_12309);
and U14848 (N_14848,N_12515,N_12909);
nand U14849 (N_14849,N_13088,N_12860);
or U14850 (N_14850,N_12418,N_13341);
or U14851 (N_14851,N_12839,N_12781);
or U14852 (N_14852,N_13256,N_12824);
nand U14853 (N_14853,N_12112,N_12878);
xnor U14854 (N_14854,N_12903,N_12219);
and U14855 (N_14855,N_12517,N_12410);
or U14856 (N_14856,N_12593,N_12198);
nor U14857 (N_14857,N_13009,N_12711);
and U14858 (N_14858,N_12055,N_13468);
and U14859 (N_14859,N_12825,N_13302);
and U14860 (N_14860,N_12446,N_13320);
and U14861 (N_14861,N_12859,N_13294);
xor U14862 (N_14862,N_12666,N_12179);
and U14863 (N_14863,N_12968,N_13374);
nand U14864 (N_14864,N_13309,N_12826);
xnor U14865 (N_14865,N_12255,N_13276);
or U14866 (N_14866,N_12194,N_13498);
nor U14867 (N_14867,N_12410,N_12262);
nor U14868 (N_14868,N_12009,N_13068);
or U14869 (N_14869,N_12255,N_12573);
or U14870 (N_14870,N_12666,N_12247);
nand U14871 (N_14871,N_12293,N_12573);
or U14872 (N_14872,N_12443,N_13080);
xnor U14873 (N_14873,N_13060,N_13093);
nand U14874 (N_14874,N_13384,N_13147);
nand U14875 (N_14875,N_13276,N_12692);
nand U14876 (N_14876,N_12308,N_13087);
or U14877 (N_14877,N_12704,N_13246);
nor U14878 (N_14878,N_12520,N_12838);
or U14879 (N_14879,N_12313,N_13392);
and U14880 (N_14880,N_13202,N_12602);
and U14881 (N_14881,N_12468,N_12118);
nand U14882 (N_14882,N_12700,N_13433);
nor U14883 (N_14883,N_12560,N_12113);
and U14884 (N_14884,N_12115,N_12034);
nor U14885 (N_14885,N_13383,N_13373);
nand U14886 (N_14886,N_12159,N_13126);
and U14887 (N_14887,N_13189,N_13330);
nor U14888 (N_14888,N_12523,N_13313);
and U14889 (N_14889,N_13374,N_13246);
and U14890 (N_14890,N_12229,N_12864);
xor U14891 (N_14891,N_12208,N_12284);
or U14892 (N_14892,N_12696,N_12175);
xnor U14893 (N_14893,N_12355,N_13370);
nand U14894 (N_14894,N_13440,N_12585);
nand U14895 (N_14895,N_12746,N_12786);
or U14896 (N_14896,N_13479,N_12501);
and U14897 (N_14897,N_13297,N_13035);
xnor U14898 (N_14898,N_12086,N_13331);
nor U14899 (N_14899,N_12337,N_13471);
xnor U14900 (N_14900,N_12035,N_12890);
xnor U14901 (N_14901,N_12536,N_12861);
xnor U14902 (N_14902,N_13324,N_13458);
nand U14903 (N_14903,N_12714,N_12500);
nor U14904 (N_14904,N_12629,N_12158);
xnor U14905 (N_14905,N_13186,N_13192);
xor U14906 (N_14906,N_12025,N_13368);
xor U14907 (N_14907,N_12475,N_12569);
or U14908 (N_14908,N_12470,N_12709);
and U14909 (N_14909,N_12841,N_13404);
nand U14910 (N_14910,N_12557,N_13444);
or U14911 (N_14911,N_12205,N_12670);
nand U14912 (N_14912,N_12981,N_12753);
and U14913 (N_14913,N_13249,N_12176);
nor U14914 (N_14914,N_12597,N_12958);
and U14915 (N_14915,N_12668,N_12386);
nor U14916 (N_14916,N_12091,N_12428);
and U14917 (N_14917,N_13290,N_12122);
and U14918 (N_14918,N_12017,N_12262);
nor U14919 (N_14919,N_12732,N_13253);
or U14920 (N_14920,N_13349,N_13308);
or U14921 (N_14921,N_12982,N_12083);
nand U14922 (N_14922,N_12305,N_12831);
xnor U14923 (N_14923,N_13021,N_13456);
or U14924 (N_14924,N_12292,N_12571);
xor U14925 (N_14925,N_13065,N_12716);
and U14926 (N_14926,N_12775,N_13452);
and U14927 (N_14927,N_12936,N_12235);
nand U14928 (N_14928,N_13003,N_12850);
nand U14929 (N_14929,N_13288,N_13381);
nand U14930 (N_14930,N_12546,N_12140);
nor U14931 (N_14931,N_12595,N_13459);
or U14932 (N_14932,N_13368,N_13076);
nand U14933 (N_14933,N_12142,N_12866);
xor U14934 (N_14934,N_12347,N_12913);
and U14935 (N_14935,N_13485,N_12195);
nand U14936 (N_14936,N_12799,N_12097);
or U14937 (N_14937,N_13455,N_12149);
and U14938 (N_14938,N_12117,N_12811);
and U14939 (N_14939,N_12042,N_12755);
nand U14940 (N_14940,N_13142,N_12666);
xor U14941 (N_14941,N_12830,N_12309);
or U14942 (N_14942,N_12152,N_12853);
xor U14943 (N_14943,N_13299,N_12066);
nand U14944 (N_14944,N_12846,N_13153);
nand U14945 (N_14945,N_12894,N_13485);
xnor U14946 (N_14946,N_13490,N_13012);
nor U14947 (N_14947,N_12603,N_13012);
nand U14948 (N_14948,N_13384,N_12016);
or U14949 (N_14949,N_12461,N_13303);
nor U14950 (N_14950,N_12231,N_12282);
nand U14951 (N_14951,N_12127,N_12023);
or U14952 (N_14952,N_13359,N_12522);
and U14953 (N_14953,N_12674,N_13028);
and U14954 (N_14954,N_13061,N_12775);
or U14955 (N_14955,N_13136,N_13462);
or U14956 (N_14956,N_12024,N_12398);
xnor U14957 (N_14957,N_13466,N_13492);
xnor U14958 (N_14958,N_12341,N_13206);
or U14959 (N_14959,N_12880,N_12542);
nand U14960 (N_14960,N_13402,N_12454);
nand U14961 (N_14961,N_12477,N_12458);
or U14962 (N_14962,N_13322,N_12899);
or U14963 (N_14963,N_13382,N_13218);
and U14964 (N_14964,N_13443,N_13406);
and U14965 (N_14965,N_13111,N_12920);
or U14966 (N_14966,N_13084,N_12490);
or U14967 (N_14967,N_12476,N_12336);
nand U14968 (N_14968,N_13115,N_12550);
nor U14969 (N_14969,N_12987,N_12268);
nor U14970 (N_14970,N_12032,N_12876);
nand U14971 (N_14971,N_12749,N_12946);
nor U14972 (N_14972,N_12936,N_12188);
nor U14973 (N_14973,N_13383,N_12341);
xnor U14974 (N_14974,N_12868,N_12062);
or U14975 (N_14975,N_12250,N_12673);
nor U14976 (N_14976,N_12226,N_13479);
or U14977 (N_14977,N_12977,N_12097);
or U14978 (N_14978,N_12327,N_12733);
and U14979 (N_14979,N_12949,N_12119);
nand U14980 (N_14980,N_13409,N_13146);
nor U14981 (N_14981,N_13428,N_12412);
and U14982 (N_14982,N_13250,N_12993);
or U14983 (N_14983,N_12865,N_12341);
or U14984 (N_14984,N_12466,N_12215);
nor U14985 (N_14985,N_12310,N_12325);
and U14986 (N_14986,N_12811,N_12937);
nand U14987 (N_14987,N_12773,N_12652);
nor U14988 (N_14988,N_12638,N_12044);
and U14989 (N_14989,N_12072,N_13171);
nor U14990 (N_14990,N_13139,N_12764);
xnor U14991 (N_14991,N_13145,N_13292);
xor U14992 (N_14992,N_12481,N_13458);
nor U14993 (N_14993,N_12110,N_13407);
nor U14994 (N_14994,N_12025,N_13148);
xor U14995 (N_14995,N_12302,N_12683);
nand U14996 (N_14996,N_12274,N_12911);
nor U14997 (N_14997,N_12889,N_12474);
or U14998 (N_14998,N_12386,N_12871);
xnor U14999 (N_14999,N_12426,N_12762);
or UO_0 (O_0,N_13725,N_13560);
nand UO_1 (O_1,N_13569,N_13822);
or UO_2 (O_2,N_14260,N_14554);
nand UO_3 (O_3,N_14794,N_14327);
nor UO_4 (O_4,N_13803,N_14171);
or UO_5 (O_5,N_14611,N_14409);
nand UO_6 (O_6,N_14702,N_14205);
nor UO_7 (O_7,N_14383,N_14164);
or UO_8 (O_8,N_14182,N_14743);
or UO_9 (O_9,N_14669,N_14655);
or UO_10 (O_10,N_14757,N_13793);
xnor UO_11 (O_11,N_14213,N_13788);
nand UO_12 (O_12,N_14201,N_13740);
xnor UO_13 (O_13,N_13513,N_14496);
and UO_14 (O_14,N_14696,N_14298);
xor UO_15 (O_15,N_14106,N_14139);
xnor UO_16 (O_16,N_14031,N_13970);
xnor UO_17 (O_17,N_13898,N_14278);
xnor UO_18 (O_18,N_14402,N_14077);
nand UO_19 (O_19,N_14482,N_14452);
and UO_20 (O_20,N_13629,N_13991);
xnor UO_21 (O_21,N_14878,N_14625);
and UO_22 (O_22,N_14271,N_14528);
nand UO_23 (O_23,N_13979,N_14360);
and UO_24 (O_24,N_13829,N_13996);
xor UO_25 (O_25,N_14776,N_14082);
nor UO_26 (O_26,N_13533,N_14939);
nand UO_27 (O_27,N_14958,N_13728);
nor UO_28 (O_28,N_14300,N_14584);
and UO_29 (O_29,N_14886,N_14431);
or UO_30 (O_30,N_13696,N_13734);
and UO_31 (O_31,N_14473,N_14007);
or UO_32 (O_32,N_13971,N_14324);
or UO_33 (O_33,N_13877,N_14196);
xnor UO_34 (O_34,N_14217,N_13630);
nand UO_35 (O_35,N_14718,N_14469);
xnor UO_36 (O_36,N_14839,N_13522);
nor UO_37 (O_37,N_14583,N_14859);
nand UO_38 (O_38,N_13792,N_14172);
and UO_39 (O_39,N_13860,N_14270);
xor UO_40 (O_40,N_13949,N_14912);
nor UO_41 (O_41,N_14115,N_14935);
or UO_42 (O_42,N_14520,N_14050);
or UO_43 (O_43,N_14305,N_13854);
nand UO_44 (O_44,N_14425,N_14013);
nor UO_45 (O_45,N_14899,N_13928);
nand UO_46 (O_46,N_14773,N_14328);
nand UO_47 (O_47,N_14098,N_13907);
and UO_48 (O_48,N_14051,N_14600);
and UO_49 (O_49,N_13779,N_13948);
and UO_50 (O_50,N_13733,N_13889);
nor UO_51 (O_51,N_14665,N_13802);
nor UO_52 (O_52,N_14130,N_14789);
or UO_53 (O_53,N_14489,N_13963);
nor UO_54 (O_54,N_13552,N_13842);
and UO_55 (O_55,N_13591,N_14382);
xor UO_56 (O_56,N_14845,N_14184);
xnor UO_57 (O_57,N_14813,N_13915);
nand UO_58 (O_58,N_13738,N_13605);
nor UO_59 (O_59,N_14786,N_14986);
and UO_60 (O_60,N_13755,N_13878);
nand UO_61 (O_61,N_14540,N_14578);
or UO_62 (O_62,N_14936,N_14323);
nand UO_63 (O_63,N_14998,N_13961);
and UO_64 (O_64,N_13615,N_14762);
or UO_65 (O_65,N_13544,N_13632);
or UO_66 (O_66,N_14165,N_14512);
or UO_67 (O_67,N_13504,N_14390);
and UO_68 (O_68,N_13864,N_13609);
or UO_69 (O_69,N_13910,N_14840);
xor UO_70 (O_70,N_13767,N_14521);
nor UO_71 (O_71,N_14570,N_13776);
nor UO_72 (O_72,N_14101,N_13703);
xnor UO_73 (O_73,N_14945,N_13758);
and UO_74 (O_74,N_13590,N_14189);
or UO_75 (O_75,N_14000,N_14395);
or UO_76 (O_76,N_14946,N_13699);
and UO_77 (O_77,N_14032,N_13697);
nand UO_78 (O_78,N_14659,N_13550);
nand UO_79 (O_79,N_14123,N_14285);
xnor UO_80 (O_80,N_14487,N_13627);
nand UO_81 (O_81,N_14124,N_14349);
xor UO_82 (O_82,N_14310,N_13862);
or UO_83 (O_83,N_13705,N_14564);
nand UO_84 (O_84,N_14286,N_14175);
and UO_85 (O_85,N_14396,N_14351);
or UO_86 (O_86,N_14713,N_14420);
nand UO_87 (O_87,N_13594,N_14519);
nor UO_88 (O_88,N_13821,N_13894);
and UO_89 (O_89,N_13893,N_13818);
or UO_90 (O_90,N_13859,N_14173);
nand UO_91 (O_91,N_14903,N_14118);
or UO_92 (O_92,N_13631,N_13500);
or UO_93 (O_93,N_13678,N_14767);
and UO_94 (O_94,N_13865,N_14345);
and UO_95 (O_95,N_14891,N_14837);
nor UO_96 (O_96,N_13811,N_14072);
xnor UO_97 (O_97,N_14879,N_14457);
and UO_98 (O_98,N_13666,N_14257);
and UO_99 (O_99,N_13518,N_14526);
xnor UO_100 (O_100,N_14251,N_14111);
xnor UO_101 (O_101,N_14577,N_14507);
nand UO_102 (O_102,N_14846,N_14277);
nor UO_103 (O_103,N_14373,N_14368);
xor UO_104 (O_104,N_14694,N_14557);
xnor UO_105 (O_105,N_14188,N_14036);
nand UO_106 (O_106,N_14601,N_14391);
nor UO_107 (O_107,N_13625,N_14092);
or UO_108 (O_108,N_14571,N_14574);
nor UO_109 (O_109,N_13837,N_14437);
nor UO_110 (O_110,N_14445,N_13742);
nand UO_111 (O_111,N_13838,N_13551);
and UO_112 (O_112,N_14350,N_14353);
or UO_113 (O_113,N_14676,N_14261);
and UO_114 (O_114,N_14318,N_14947);
or UO_115 (O_115,N_14765,N_13580);
and UO_116 (O_116,N_14599,N_13538);
and UO_117 (O_117,N_14258,N_14126);
nor UO_118 (O_118,N_13801,N_14864);
nand UO_119 (O_119,N_14099,N_13932);
xor UO_120 (O_120,N_14059,N_14400);
and UO_121 (O_121,N_13724,N_14957);
or UO_122 (O_122,N_13945,N_13817);
nor UO_123 (O_123,N_13529,N_14888);
and UO_124 (O_124,N_14208,N_14569);
nand UO_125 (O_125,N_13735,N_14547);
xor UO_126 (O_126,N_14125,N_14313);
or UO_127 (O_127,N_14828,N_13954);
xnor UO_128 (O_128,N_14340,N_13897);
xor UO_129 (O_129,N_14646,N_14800);
nand UO_130 (O_130,N_14410,N_13964);
and UO_131 (O_131,N_14307,N_14754);
nand UO_132 (O_132,N_13641,N_14472);
and UO_133 (O_133,N_14769,N_14679);
nor UO_134 (O_134,N_14451,N_14668);
and UO_135 (O_135,N_14783,N_14635);
nand UO_136 (O_136,N_13731,N_14596);
nand UO_137 (O_137,N_13923,N_14114);
or UO_138 (O_138,N_14083,N_14008);
xor UO_139 (O_139,N_13691,N_13913);
and UO_140 (O_140,N_14953,N_13503);
nand UO_141 (O_141,N_14359,N_13834);
nand UO_142 (O_142,N_14576,N_14052);
nand UO_143 (O_143,N_13832,N_14833);
and UO_144 (O_144,N_14136,N_14399);
nor UO_145 (O_145,N_14931,N_14242);
xor UO_146 (O_146,N_14781,N_13657);
or UO_147 (O_147,N_14597,N_13583);
nor UO_148 (O_148,N_14023,N_14636);
or UO_149 (O_149,N_14291,N_14621);
xor UO_150 (O_150,N_14219,N_14296);
and UO_151 (O_151,N_14539,N_13671);
and UO_152 (O_152,N_14742,N_13927);
nor UO_153 (O_153,N_14568,N_13649);
or UO_154 (O_154,N_14272,N_14731);
nor UO_155 (O_155,N_13872,N_14394);
nor UO_156 (O_156,N_14216,N_14921);
and UO_157 (O_157,N_14440,N_13925);
xnor UO_158 (O_158,N_13506,N_13637);
nor UO_159 (O_159,N_14110,N_14084);
nor UO_160 (O_160,N_14553,N_14593);
and UO_161 (O_161,N_13798,N_13562);
xnor UO_162 (O_162,N_14075,N_14501);
xnor UO_163 (O_163,N_14483,N_14037);
or UO_164 (O_164,N_13698,N_14458);
and UO_165 (O_165,N_14346,N_13739);
nor UO_166 (O_166,N_14317,N_13748);
xnor UO_167 (O_167,N_14787,N_13828);
and UO_168 (O_168,N_14068,N_13804);
or UO_169 (O_169,N_14901,N_14397);
nand UO_170 (O_170,N_14380,N_14955);
or UO_171 (O_171,N_14645,N_14476);
nand UO_172 (O_172,N_13723,N_14985);
nand UO_173 (O_173,N_14371,N_14211);
nor UO_174 (O_174,N_14705,N_14893);
and UO_175 (O_175,N_14259,N_14478);
xor UO_176 (O_176,N_14950,N_14620);
xor UO_177 (O_177,N_13519,N_13572);
or UO_178 (O_178,N_13726,N_14863);
and UO_179 (O_179,N_13539,N_13711);
or UO_180 (O_180,N_14230,N_14628);
and UO_181 (O_181,N_14143,N_13962);
and UO_182 (O_182,N_14289,N_14269);
nand UO_183 (O_183,N_14653,N_14057);
or UO_184 (O_184,N_14081,N_13730);
nor UO_185 (O_185,N_14943,N_13757);
nand UO_186 (O_186,N_14214,N_14393);
nor UO_187 (O_187,N_14290,N_14322);
and UO_188 (O_188,N_14215,N_14464);
and UO_189 (O_189,N_14502,N_14632);
nand UO_190 (O_190,N_13814,N_14799);
and UO_191 (O_191,N_13589,N_13542);
nor UO_192 (O_192,N_14090,N_14884);
xnor UO_193 (O_193,N_13866,N_14709);
or UO_194 (O_194,N_14352,N_14775);
nor UO_195 (O_195,N_13879,N_14011);
and UO_196 (O_196,N_13940,N_13880);
xnor UO_197 (O_197,N_14369,N_14686);
and UO_198 (O_198,N_14212,N_13887);
or UO_199 (O_199,N_14316,N_14804);
nor UO_200 (O_200,N_14944,N_14825);
and UO_201 (O_201,N_14151,N_13823);
or UO_202 (O_202,N_14657,N_14342);
nand UO_203 (O_203,N_14039,N_14681);
nor UO_204 (O_204,N_14674,N_13869);
or UO_205 (O_205,N_14163,N_14745);
or UO_206 (O_206,N_14224,N_14002);
nand UO_207 (O_207,N_13981,N_14241);
nand UO_208 (O_208,N_14723,N_14329);
or UO_209 (O_209,N_14060,N_14510);
xor UO_210 (O_210,N_14275,N_14306);
nand UO_211 (O_211,N_14087,N_14357);
and UO_212 (O_212,N_14870,N_13772);
nor UO_213 (O_213,N_13520,N_14695);
xor UO_214 (O_214,N_14732,N_14253);
nand UO_215 (O_215,N_14119,N_14406);
or UO_216 (O_216,N_14595,N_14877);
and UO_217 (O_217,N_14479,N_13936);
nand UO_218 (O_218,N_13867,N_14146);
xor UO_219 (O_219,N_14848,N_13848);
or UO_220 (O_220,N_13807,N_13515);
xnor UO_221 (O_221,N_14690,N_13511);
xnor UO_222 (O_222,N_14811,N_14245);
and UO_223 (O_223,N_14439,N_13507);
or UO_224 (O_224,N_14860,N_14546);
nor UO_225 (O_225,N_14838,N_13890);
or UO_226 (O_226,N_13931,N_14281);
xor UO_227 (O_227,N_13824,N_13899);
and UO_228 (O_228,N_14503,N_14375);
xnor UO_229 (O_229,N_13516,N_14630);
nor UO_230 (O_230,N_14456,N_14065);
and UO_231 (O_231,N_13935,N_13623);
nand UO_232 (O_232,N_14384,N_14698);
or UO_233 (O_233,N_13694,N_13980);
nor UO_234 (O_234,N_14887,N_14462);
and UO_235 (O_235,N_13791,N_14268);
nor UO_236 (O_236,N_13617,N_14766);
nor UO_237 (O_237,N_14461,N_14187);
xnor UO_238 (O_238,N_14134,N_14807);
nand UO_239 (O_239,N_14527,N_14552);
nand UO_240 (O_240,N_14062,N_14466);
nor UO_241 (O_241,N_14490,N_13718);
and UO_242 (O_242,N_14429,N_13836);
nand UO_243 (O_243,N_14565,N_14778);
and UO_244 (O_244,N_14774,N_13926);
and UO_245 (O_245,N_14956,N_14532);
and UO_246 (O_246,N_13958,N_14685);
nor UO_247 (O_247,N_14549,N_14193);
nand UO_248 (O_248,N_14256,N_13598);
nand UO_249 (O_249,N_14024,N_14049);
and UO_250 (O_250,N_14430,N_14844);
or UO_251 (O_251,N_14386,N_14021);
xor UO_252 (O_252,N_13786,N_14591);
or UO_253 (O_253,N_14169,N_14894);
and UO_254 (O_254,N_14882,N_14923);
xor UO_255 (O_255,N_14426,N_14561);
nor UO_256 (O_256,N_14204,N_13827);
nand UO_257 (O_257,N_13536,N_14304);
xnor UO_258 (O_258,N_13690,N_14150);
nand UO_259 (O_259,N_14728,N_14895);
nand UO_260 (O_260,N_13669,N_14379);
and UO_261 (O_261,N_14977,N_13687);
or UO_262 (O_262,N_14744,N_14623);
and UO_263 (O_263,N_14548,N_14952);
nand UO_264 (O_264,N_14881,N_13595);
and UO_265 (O_265,N_14474,N_13985);
nand UO_266 (O_266,N_14356,N_14999);
and UO_267 (O_267,N_13933,N_14969);
or UO_268 (O_268,N_13722,N_13847);
nor UO_269 (O_269,N_14274,N_14834);
nand UO_270 (O_270,N_14941,N_14243);
nor UO_271 (O_271,N_14103,N_14581);
and UO_272 (O_272,N_13553,N_13709);
nand UO_273 (O_273,N_14616,N_13689);
nand UO_274 (O_274,N_14792,N_14897);
and UO_275 (O_275,N_13628,N_14129);
xor UO_276 (O_276,N_14029,N_14132);
nor UO_277 (O_277,N_14720,N_13902);
nor UO_278 (O_278,N_13568,N_14917);
nand UO_279 (O_279,N_13712,N_13686);
nor UO_280 (O_280,N_13639,N_14691);
and UO_281 (O_281,N_13976,N_14603);
nor UO_282 (O_282,N_13903,N_14707);
and UO_283 (O_283,N_14942,N_14209);
xor UO_284 (O_284,N_13799,N_14160);
nand UO_285 (O_285,N_14017,N_14613);
and UO_286 (O_286,N_14711,N_14566);
or UO_287 (O_287,N_14314,N_14078);
or UO_288 (O_288,N_14159,N_14876);
or UO_289 (O_289,N_14419,N_14580);
or UO_290 (O_290,N_14378,N_14610);
nand UO_291 (O_291,N_13951,N_14325);
xnor UO_292 (O_292,N_13588,N_14348);
nor UO_293 (O_293,N_13912,N_14053);
and UO_294 (O_294,N_14135,N_13756);
xnor UO_295 (O_295,N_14856,N_13787);
nand UO_296 (O_296,N_14010,N_14167);
or UO_297 (O_297,N_14889,N_14055);
and UO_298 (O_298,N_14333,N_14176);
and UO_299 (O_299,N_14066,N_14207);
nand UO_300 (O_300,N_14477,N_14654);
or UO_301 (O_301,N_14725,N_13762);
nand UO_302 (O_302,N_14093,N_14040);
nor UO_303 (O_303,N_14320,N_14726);
and UO_304 (O_304,N_14658,N_14096);
nor UO_305 (O_305,N_14722,N_13651);
nor UO_306 (O_306,N_14843,N_13874);
nor UO_307 (O_307,N_14928,N_14818);
or UO_308 (O_308,N_14388,N_14988);
nor UO_309 (O_309,N_14377,N_14675);
nor UO_310 (O_310,N_14531,N_14232);
and UO_311 (O_311,N_13921,N_14225);
and UO_312 (O_312,N_14308,N_14220);
and UO_313 (O_313,N_13843,N_14004);
xor UO_314 (O_314,N_13660,N_14047);
nor UO_315 (O_315,N_13541,N_14138);
nand UO_316 (O_316,N_14233,N_14738);
and UO_317 (O_317,N_14868,N_13673);
or UO_318 (O_318,N_14337,N_14663);
and UO_319 (O_319,N_14435,N_13707);
and UO_320 (O_320,N_14244,N_13825);
xnor UO_321 (O_321,N_13797,N_14166);
nor UO_322 (O_322,N_14624,N_14976);
and UO_323 (O_323,N_14045,N_14949);
nand UO_324 (O_324,N_13622,N_14930);
nor UO_325 (O_325,N_14226,N_14575);
or UO_326 (O_326,N_13905,N_13614);
nand UO_327 (O_327,N_14602,N_14609);
nor UO_328 (O_328,N_14934,N_14341);
xnor UO_329 (O_329,N_14044,N_14816);
nor UO_330 (O_330,N_14697,N_14760);
nand UO_331 (O_331,N_14438,N_14805);
nor UO_332 (O_332,N_14128,N_14617);
and UO_333 (O_333,N_14513,N_14442);
or UO_334 (O_334,N_14538,N_14534);
nand UO_335 (O_335,N_13741,N_14853);
nand UO_336 (O_336,N_14319,N_14303);
nor UO_337 (O_337,N_14692,N_14585);
nor UO_338 (O_338,N_14434,N_14819);
nand UO_339 (O_339,N_13620,N_14606);
nor UO_340 (O_340,N_14486,N_13557);
xor UO_341 (O_341,N_13561,N_14417);
or UO_342 (O_342,N_13839,N_14122);
nor UO_343 (O_343,N_13987,N_14687);
nand UO_344 (O_344,N_13886,N_14475);
and UO_345 (O_345,N_13960,N_14142);
xnor UO_346 (O_346,N_13577,N_14265);
nor UO_347 (O_347,N_14033,N_13853);
nor UO_348 (O_348,N_14974,N_14688);
nand UO_349 (O_349,N_14823,N_13806);
nor UO_350 (O_350,N_14407,N_14492);
or UO_351 (O_351,N_13567,N_13876);
nor UO_352 (O_352,N_14117,N_13773);
xnor UO_353 (O_353,N_14835,N_14283);
nand UO_354 (O_354,N_13713,N_14755);
nor UO_355 (O_355,N_13545,N_14642);
nand UO_356 (O_356,N_14749,N_13685);
xnor UO_357 (O_357,N_14467,N_14076);
xor UO_358 (O_358,N_13770,N_14206);
xor UO_359 (O_359,N_14071,N_13548);
nor UO_360 (O_360,N_14504,N_14218);
nand UO_361 (O_361,N_13775,N_14018);
or UO_362 (O_362,N_14362,N_14385);
nand UO_363 (O_363,N_13900,N_14841);
nor UO_364 (O_364,N_14523,N_13579);
xor UO_365 (O_365,N_13992,N_14847);
or UO_366 (O_366,N_14761,N_14682);
or UO_367 (O_367,N_13574,N_13596);
and UO_368 (O_368,N_14174,N_13535);
xor UO_369 (O_369,N_13676,N_13967);
nor UO_370 (O_370,N_14481,N_13861);
nor UO_371 (O_371,N_13835,N_14815);
or UO_372 (O_372,N_14006,N_14292);
nor UO_373 (O_373,N_14598,N_13582);
nand UO_374 (O_374,N_14716,N_14727);
and UO_375 (O_375,N_14647,N_13665);
or UO_376 (O_376,N_13512,N_13700);
nor UO_377 (O_377,N_14756,N_13968);
or UO_378 (O_378,N_14719,N_14276);
xor UO_379 (O_379,N_14180,N_14148);
xor UO_380 (O_380,N_13809,N_13808);
and UO_381 (O_381,N_14963,N_14714);
nand UO_382 (O_382,N_14608,N_13653);
xnor UO_383 (O_383,N_13969,N_14906);
nand UO_384 (O_384,N_14890,N_14444);
nor UO_385 (O_385,N_14951,N_14618);
nor UO_386 (O_386,N_14460,N_14293);
and UO_387 (O_387,N_14508,N_14607);
or UO_388 (O_388,N_13941,N_14104);
or UO_389 (O_389,N_13844,N_14671);
nor UO_390 (O_390,N_14192,N_13959);
nand UO_391 (O_391,N_14109,N_14038);
nand UO_392 (O_392,N_13584,N_14954);
nor UO_393 (O_393,N_13692,N_13729);
or UO_394 (O_394,N_14121,N_13855);
xor UO_395 (O_395,N_14924,N_14493);
xnor UO_396 (O_396,N_13763,N_14043);
and UO_397 (O_397,N_13736,N_14488);
and UO_398 (O_398,N_14423,N_14177);
and UO_399 (O_399,N_14721,N_14237);
nand UO_400 (O_400,N_13558,N_14972);
nand UO_401 (O_401,N_14824,N_13505);
or UO_402 (O_402,N_14905,N_14614);
nand UO_403 (O_403,N_14803,N_14336);
nor UO_404 (O_404,N_14900,N_13634);
xor UO_405 (O_405,N_13523,N_14465);
or UO_406 (O_406,N_14249,N_14374);
and UO_407 (O_407,N_14959,N_13546);
and UO_408 (O_408,N_13904,N_14874);
nor UO_409 (O_409,N_14414,N_13708);
and UO_410 (O_410,N_14842,N_14330);
nor UO_411 (O_411,N_14938,N_14734);
and UO_412 (O_412,N_14195,N_13796);
and UO_413 (O_413,N_14817,N_13895);
and UO_414 (O_414,N_13918,N_14730);
xnor UO_415 (O_415,N_14662,N_14433);
nor UO_416 (O_416,N_14063,N_14515);
xnor UO_417 (O_417,N_13619,N_13587);
xor UO_418 (O_418,N_13565,N_14222);
and UO_419 (O_419,N_14915,N_14338);
or UO_420 (O_420,N_14637,N_14067);
nor UO_421 (O_421,N_13717,N_14471);
nand UO_422 (O_422,N_14470,N_14358);
or UO_423 (O_423,N_14354,N_13576);
xnor UO_424 (O_424,N_14186,N_14459);
nor UO_425 (O_425,N_14364,N_14416);
and UO_426 (O_426,N_13621,N_14693);
and UO_427 (O_427,N_13668,N_13603);
or UO_428 (O_428,N_14592,N_13883);
or UO_429 (O_429,N_14056,N_14074);
nand UO_430 (O_430,N_13785,N_13950);
and UO_431 (O_431,N_13957,N_13974);
or UO_432 (O_432,N_13563,N_14904);
xor UO_433 (O_433,N_14820,N_13765);
or UO_434 (O_434,N_13909,N_13953);
nor UO_435 (O_435,N_14793,N_14048);
and UO_436 (O_436,N_14763,N_14850);
nor UO_437 (O_437,N_14750,N_14061);
xor UO_438 (O_438,N_13986,N_14131);
nand UO_439 (O_439,N_13527,N_14545);
nor UO_440 (O_440,N_13841,N_14643);
nor UO_441 (O_441,N_14558,N_14133);
nand UO_442 (O_442,N_13680,N_14246);
nor UO_443 (O_443,N_14965,N_13911);
nand UO_444 (O_444,N_14594,N_14559);
xor UO_445 (O_445,N_14808,N_13831);
nand UO_446 (O_446,N_14009,N_14740);
and UO_447 (O_447,N_13679,N_13752);
nor UO_448 (O_448,N_13934,N_13988);
nand UO_449 (O_449,N_13661,N_13789);
nand UO_450 (O_450,N_14925,N_14447);
or UO_451 (O_451,N_13531,N_13783);
nor UO_452 (O_452,N_14003,N_14480);
xnor UO_453 (O_453,N_14387,N_13721);
xnor UO_454 (O_454,N_13599,N_14927);
or UO_455 (O_455,N_14372,N_14537);
xnor UO_456 (O_456,N_13664,N_13652);
nor UO_457 (O_457,N_14588,N_14582);
nor UO_458 (O_458,N_14398,N_14499);
xnor UO_459 (O_459,N_14550,N_14535);
nand UO_460 (O_460,N_14780,N_14234);
and UO_461 (O_461,N_14911,N_14401);
xnor UO_462 (O_462,N_14966,N_13704);
nor UO_463 (O_463,N_14996,N_14315);
xor UO_464 (O_464,N_13695,N_13759);
nor UO_465 (O_465,N_13606,N_13849);
nand UO_466 (O_466,N_14405,N_13743);
or UO_467 (O_467,N_14615,N_14343);
and UO_468 (O_468,N_14144,N_13858);
xor UO_469 (O_469,N_14197,N_14147);
or UO_470 (O_470,N_14759,N_14670);
xor UO_471 (O_471,N_13524,N_13999);
nand UO_472 (O_472,N_14962,N_14858);
and UO_473 (O_473,N_14883,N_14748);
nand UO_474 (O_474,N_13677,N_14231);
or UO_475 (O_475,N_14255,N_14376);
xor UO_476 (O_476,N_13501,N_13761);
xnor UO_477 (O_477,N_13607,N_14854);
nor UO_478 (O_478,N_13944,N_14673);
xor UO_479 (O_479,N_14604,N_14105);
nand UO_480 (O_480,N_14677,N_14516);
or UO_481 (O_481,N_14875,N_14700);
nor UO_482 (O_482,N_14411,N_13920);
nand UO_483 (O_483,N_14266,N_14831);
xnor UO_484 (O_484,N_13532,N_14155);
or UO_485 (O_485,N_14543,N_14035);
nor UO_486 (O_486,N_14712,N_14724);
nand UO_487 (O_487,N_14267,N_13947);
or UO_488 (O_488,N_14107,N_13517);
nor UO_489 (O_489,N_14079,N_14530);
nor UO_490 (O_490,N_14961,N_13737);
xnor UO_491 (O_491,N_14454,N_14770);
nand UO_492 (O_492,N_14703,N_14992);
or UO_493 (O_493,N_14273,N_14252);
nand UO_494 (O_494,N_14729,N_13857);
nand UO_495 (O_495,N_14661,N_14542);
nand UO_496 (O_496,N_14086,N_13896);
or UO_497 (O_497,N_14733,N_13509);
nand UO_498 (O_498,N_13593,N_13514);
xnor UO_499 (O_499,N_14975,N_14027);
or UO_500 (O_500,N_13871,N_13845);
xnor UO_501 (O_501,N_13924,N_14240);
nand UO_502 (O_502,N_14484,N_13840);
and UO_503 (O_503,N_14403,N_14170);
nand UO_504 (O_504,N_14990,N_13764);
or UO_505 (O_505,N_13601,N_14415);
nor UO_506 (O_506,N_14857,N_13597);
nand UO_507 (O_507,N_14861,N_14832);
nand UO_508 (O_508,N_14649,N_13820);
nor UO_509 (O_509,N_14015,N_13943);
nand UO_510 (O_510,N_14153,N_14994);
and UO_511 (O_511,N_13647,N_13774);
nor UO_512 (O_512,N_13656,N_14221);
nand UO_513 (O_513,N_14367,N_14287);
xor UO_514 (O_514,N_14809,N_14849);
nand UO_515 (O_515,N_13648,N_14228);
nor UO_516 (O_516,N_14737,N_14964);
and UO_517 (O_517,N_13662,N_13994);
nor UO_518 (O_518,N_14524,N_13990);
or UO_519 (O_519,N_14790,N_13795);
nor UO_520 (O_520,N_13732,N_14463);
nor UO_521 (O_521,N_14495,N_13942);
nor UO_522 (O_522,N_14198,N_13777);
nand UO_523 (O_523,N_14518,N_13908);
nand UO_524 (O_524,N_14455,N_14822);
and UO_525 (O_525,N_13586,N_13502);
nand UO_526 (O_526,N_14190,N_14448);
nor UO_527 (O_527,N_14046,N_14161);
xor UO_528 (O_528,N_14660,N_13884);
nor UO_529 (O_529,N_13901,N_14555);
nor UO_530 (O_530,N_13573,N_13720);
nor UO_531 (O_531,N_14706,N_14651);
nor UO_532 (O_532,N_13667,N_14238);
or UO_533 (O_533,N_14739,N_13833);
or UO_534 (O_534,N_13682,N_14191);
and UO_535 (O_535,N_14979,N_13939);
nor UO_536 (O_536,N_14741,N_14871);
nand UO_537 (O_537,N_14080,N_14937);
xnor UO_538 (O_538,N_13870,N_14453);
and UO_539 (O_539,N_14254,N_14920);
xnor UO_540 (O_540,N_13638,N_14648);
and UO_541 (O_541,N_13972,N_14179);
xor UO_542 (O_542,N_14094,N_14796);
xor UO_543 (O_543,N_14529,N_14710);
and UO_544 (O_544,N_14517,N_14752);
and UO_545 (O_545,N_14666,N_14590);
nand UO_546 (O_546,N_14149,N_14088);
or UO_547 (O_547,N_14626,N_14699);
nand UO_548 (O_548,N_14113,N_14301);
and UO_549 (O_549,N_13782,N_14446);
xnor UO_550 (O_550,N_13701,N_13984);
xnor UO_551 (O_551,N_14366,N_14299);
nor UO_552 (O_552,N_14223,N_14424);
or UO_553 (O_553,N_13640,N_14157);
nand UO_554 (O_554,N_14701,N_14672);
nand UO_555 (O_555,N_14779,N_14041);
nor UO_556 (O_556,N_14069,N_13525);
and UO_557 (O_557,N_14806,N_14468);
and UO_558 (O_558,N_13863,N_14814);
or UO_559 (O_559,N_14573,N_14302);
and UO_560 (O_560,N_13922,N_14797);
and UO_561 (O_561,N_13674,N_14100);
and UO_562 (O_562,N_14933,N_14812);
nor UO_563 (O_563,N_13554,N_14450);
and UO_564 (O_564,N_13683,N_14162);
or UO_565 (O_565,N_13812,N_14639);
and UO_566 (O_566,N_13747,N_14680);
and UO_567 (O_567,N_13604,N_14284);
or UO_568 (O_568,N_13805,N_14443);
and UO_569 (O_569,N_14408,N_14418);
nand UO_570 (O_570,N_13744,N_14782);
xnor UO_571 (O_571,N_14355,N_14562);
nor UO_572 (O_572,N_14137,N_13975);
nand UO_573 (O_573,N_14108,N_14326);
xor UO_574 (O_574,N_14089,N_14427);
nand UO_575 (O_575,N_13693,N_13891);
nor UO_576 (O_576,N_14509,N_14152);
or UO_577 (O_577,N_13559,N_13571);
xor UO_578 (O_578,N_14909,N_13633);
xor UO_579 (O_579,N_14913,N_13534);
or UO_580 (O_580,N_13715,N_14514);
or UO_581 (O_581,N_14332,N_14851);
and UO_582 (O_582,N_14073,N_13714);
nor UO_583 (O_583,N_14960,N_13781);
and UO_584 (O_584,N_14058,N_14541);
nor UO_585 (O_585,N_13989,N_14158);
or UO_586 (O_586,N_13646,N_14629);
nor UO_587 (O_587,N_13766,N_14494);
xnor UO_588 (O_588,N_14982,N_14202);
xnor UO_589 (O_589,N_14926,N_14826);
xor UO_590 (O_590,N_14971,N_13800);
nor UO_591 (O_591,N_13750,N_14309);
or UO_592 (O_592,N_14683,N_14652);
xor UO_593 (O_593,N_14168,N_14987);
and UO_594 (O_594,N_14533,N_14634);
or UO_595 (O_595,N_14363,N_14898);
or UO_596 (O_596,N_13875,N_13616);
xnor UO_597 (O_597,N_13982,N_14500);
and UO_598 (O_598,N_14973,N_13659);
nand UO_599 (O_599,N_14932,N_14758);
or UO_600 (O_600,N_14784,N_13917);
nand UO_601 (O_601,N_13626,N_14746);
nand UO_602 (O_602,N_14589,N_14865);
nor UO_603 (O_603,N_14070,N_14321);
xor UO_604 (O_604,N_14311,N_14019);
xnor UO_605 (O_605,N_14633,N_13508);
nor UO_606 (O_606,N_14827,N_13952);
nor UO_607 (O_607,N_14919,N_14295);
xnor UO_608 (O_608,N_14717,N_13618);
or UO_609 (O_609,N_13643,N_13751);
nor UO_610 (O_610,N_14016,N_14279);
xor UO_611 (O_611,N_13881,N_14312);
nor UO_612 (O_612,N_14830,N_13760);
and UO_613 (O_613,N_13938,N_13727);
nand UO_614 (O_614,N_14948,N_13906);
and UO_615 (O_615,N_13570,N_14736);
xnor UO_616 (O_616,N_13575,N_14872);
nand UO_617 (O_617,N_14210,N_14989);
and UO_618 (O_618,N_14235,N_14156);
nand UO_619 (O_619,N_14587,N_13790);
xnor UO_620 (O_620,N_14412,N_13780);
or UO_621 (O_621,N_13816,N_13644);
xor UO_622 (O_622,N_13611,N_13753);
nor UO_623 (O_623,N_13778,N_14892);
and UO_624 (O_624,N_13675,N_14751);
nand UO_625 (O_625,N_14282,N_14112);
or UO_626 (O_626,N_14525,N_14764);
nand UO_627 (O_627,N_14922,N_14280);
xnor UO_628 (O_628,N_13610,N_13636);
or UO_629 (O_629,N_13530,N_14183);
and UO_630 (O_630,N_14993,N_14014);
nand UO_631 (O_631,N_14236,N_14704);
nand UO_632 (O_632,N_13937,N_13965);
xor UO_633 (O_633,N_14772,N_14001);
nor UO_634 (O_634,N_13655,N_14638);
xnor UO_635 (O_635,N_14127,N_14715);
xnor UO_636 (O_636,N_14030,N_14064);
or UO_637 (O_637,N_13684,N_13526);
and UO_638 (O_638,N_13745,N_14929);
and UO_639 (O_639,N_14768,N_14026);
or UO_640 (O_640,N_14619,N_14567);
nand UO_641 (O_641,N_14239,N_14862);
or UO_642 (O_642,N_13998,N_13566);
or UO_643 (O_643,N_14248,N_14991);
nor UO_644 (O_644,N_14914,N_14511);
nor UO_645 (O_645,N_14498,N_13585);
and UO_646 (O_646,N_14263,N_14970);
or UO_647 (O_647,N_13578,N_14428);
nand UO_648 (O_648,N_14344,N_14650);
xnor UO_649 (O_649,N_13528,N_13672);
and UO_650 (O_650,N_13966,N_13916);
nor UO_651 (O_651,N_13882,N_14381);
and UO_652 (O_652,N_14432,N_13654);
xor UO_653 (O_653,N_13521,N_14102);
and UO_654 (O_654,N_14572,N_14896);
nand UO_655 (O_655,N_14968,N_13537);
and UO_656 (O_656,N_14873,N_14997);
nor UO_657 (O_657,N_14556,N_14042);
xnor UO_658 (O_658,N_14631,N_14200);
nand UO_659 (O_659,N_14185,N_14250);
or UO_660 (O_660,N_13768,N_13930);
nor UO_661 (O_661,N_14141,N_14664);
and UO_662 (O_662,N_14264,N_13997);
nor UO_663 (O_663,N_14907,N_14491);
nor UO_664 (O_664,N_14034,N_13602);
xnor UO_665 (O_665,N_13868,N_14563);
nor UO_666 (O_666,N_14902,N_13658);
nand UO_667 (O_667,N_14984,N_14798);
xor UO_668 (O_668,N_13749,N_13645);
xor UO_669 (O_669,N_14795,N_14449);
nand UO_670 (O_670,N_13830,N_13810);
nand UO_671 (O_671,N_14983,N_14028);
or UO_672 (O_672,N_14339,N_14560);
nor UO_673 (O_673,N_14644,N_13719);
xnor UO_674 (O_674,N_13549,N_13608);
nor UO_675 (O_675,N_14331,N_14640);
nor UO_676 (O_676,N_13794,N_14980);
nand UO_677 (O_677,N_13993,N_13929);
and UO_678 (O_678,N_13688,N_13581);
and UO_679 (O_679,N_14365,N_14855);
xnor UO_680 (O_680,N_14181,N_14821);
or UO_681 (O_681,N_14852,N_14777);
xnor UO_682 (O_682,N_13650,N_14022);
nand UO_683 (O_683,N_14689,N_13973);
nand UO_684 (O_684,N_13919,N_14612);
or UO_685 (O_685,N_13612,N_14627);
nor UO_686 (O_686,N_14771,N_13850);
xor UO_687 (O_687,N_13784,N_13955);
nand UO_688 (O_688,N_14505,N_13681);
xor UO_689 (O_689,N_14753,N_13543);
nor UO_690 (O_690,N_14145,N_14005);
nor UO_691 (O_691,N_14880,N_13613);
and UO_692 (O_692,N_14422,N_14918);
and UO_693 (O_693,N_14916,N_14586);
and UO_694 (O_694,N_14908,N_14389);
nand UO_695 (O_695,N_13892,N_13556);
nor UO_696 (O_696,N_14506,N_13746);
xnor UO_697 (O_697,N_14347,N_14656);
nand UO_698 (O_698,N_13706,N_14641);
and UO_699 (O_699,N_14392,N_13564);
or UO_700 (O_700,N_13754,N_13846);
xor UO_701 (O_701,N_14544,N_13995);
xor UO_702 (O_702,N_13983,N_14667);
and UO_703 (O_703,N_14054,N_14885);
or UO_704 (O_704,N_13710,N_14335);
and UO_705 (O_705,N_13642,N_13914);
nor UO_706 (O_706,N_13873,N_14485);
or UO_707 (O_707,N_14866,N_13670);
nor UO_708 (O_708,N_14097,N_14747);
xnor UO_709 (O_709,N_14536,N_14178);
and UO_710 (O_710,N_14020,N_13663);
nand UO_711 (O_711,N_14334,N_14294);
or UO_712 (O_712,N_14361,N_14227);
and UO_713 (O_713,N_14940,N_14154);
or UO_714 (O_714,N_13510,N_13624);
and UO_715 (O_715,N_14116,N_14869);
nor UO_716 (O_716,N_14085,N_14708);
nand UO_717 (O_717,N_13702,N_13815);
or UO_718 (O_718,N_14288,N_14095);
xnor UO_719 (O_719,N_14297,N_14836);
or UO_720 (O_720,N_14194,N_13977);
and UO_721 (O_721,N_14788,N_13956);
xor UO_722 (O_722,N_14791,N_14404);
and UO_723 (O_723,N_13888,N_13851);
or UO_724 (O_724,N_14421,N_14203);
nor UO_725 (O_725,N_14262,N_14497);
and UO_726 (O_726,N_14735,N_14810);
xnor UO_727 (O_727,N_13978,N_14995);
xor UO_728 (O_728,N_14785,N_13547);
and UO_729 (O_729,N_14981,N_13819);
and UO_730 (O_730,N_14622,N_14436);
nor UO_731 (O_731,N_14579,N_14199);
and UO_732 (O_732,N_14025,N_14605);
or UO_733 (O_733,N_14012,N_13716);
or UO_734 (O_734,N_13635,N_14967);
and UO_735 (O_735,N_13555,N_14684);
nand UO_736 (O_736,N_14867,N_13540);
xnor UO_737 (O_737,N_14229,N_13600);
and UO_738 (O_738,N_13852,N_13769);
nand UO_739 (O_739,N_14120,N_14091);
and UO_740 (O_740,N_13856,N_14802);
nand UO_741 (O_741,N_13592,N_14801);
nor UO_742 (O_742,N_13771,N_14910);
nor UO_743 (O_743,N_14413,N_14370);
nand UO_744 (O_744,N_14522,N_14678);
nand UO_745 (O_745,N_14978,N_14829);
nand UO_746 (O_746,N_13946,N_14247);
and UO_747 (O_747,N_13813,N_14551);
and UO_748 (O_748,N_14140,N_13885);
or UO_749 (O_749,N_13826,N_14441);
or UO_750 (O_750,N_14490,N_14656);
or UO_751 (O_751,N_13621,N_13908);
xnor UO_752 (O_752,N_13948,N_13594);
or UO_753 (O_753,N_13900,N_14588);
nand UO_754 (O_754,N_13551,N_14538);
nand UO_755 (O_755,N_14752,N_14343);
and UO_756 (O_756,N_13979,N_14911);
nor UO_757 (O_757,N_14140,N_14427);
or UO_758 (O_758,N_14428,N_14830);
or UO_759 (O_759,N_13910,N_14785);
and UO_760 (O_760,N_14393,N_14415);
nor UO_761 (O_761,N_14384,N_14345);
xor UO_762 (O_762,N_14451,N_13946);
xnor UO_763 (O_763,N_14677,N_14432);
and UO_764 (O_764,N_14471,N_14078);
nand UO_765 (O_765,N_14415,N_14768);
and UO_766 (O_766,N_14275,N_14497);
nand UO_767 (O_767,N_14814,N_14802);
and UO_768 (O_768,N_14164,N_14955);
xor UO_769 (O_769,N_14069,N_13574);
or UO_770 (O_770,N_14362,N_13995);
nor UO_771 (O_771,N_14433,N_13935);
nor UO_772 (O_772,N_14067,N_13629);
and UO_773 (O_773,N_14457,N_14627);
or UO_774 (O_774,N_13824,N_14432);
xnor UO_775 (O_775,N_14916,N_14056);
xor UO_776 (O_776,N_13608,N_14883);
or UO_777 (O_777,N_14705,N_14183);
nand UO_778 (O_778,N_14795,N_14289);
nor UO_779 (O_779,N_13997,N_13875);
and UO_780 (O_780,N_13810,N_14896);
and UO_781 (O_781,N_14758,N_14978);
and UO_782 (O_782,N_14008,N_14164);
nor UO_783 (O_783,N_13781,N_14137);
xor UO_784 (O_784,N_14417,N_14080);
nor UO_785 (O_785,N_13572,N_14837);
nor UO_786 (O_786,N_13705,N_14200);
xnor UO_787 (O_787,N_14096,N_14847);
and UO_788 (O_788,N_14126,N_14563);
and UO_789 (O_789,N_14224,N_14433);
or UO_790 (O_790,N_14792,N_14294);
xor UO_791 (O_791,N_14404,N_13760);
xor UO_792 (O_792,N_13580,N_14216);
nor UO_793 (O_793,N_14998,N_14964);
xnor UO_794 (O_794,N_13949,N_14280);
and UO_795 (O_795,N_13914,N_13867);
or UO_796 (O_796,N_14206,N_14069);
xnor UO_797 (O_797,N_14933,N_14166);
nor UO_798 (O_798,N_13523,N_14342);
nor UO_799 (O_799,N_13858,N_14207);
and UO_800 (O_800,N_13921,N_13985);
or UO_801 (O_801,N_14807,N_14753);
xor UO_802 (O_802,N_14394,N_14526);
nand UO_803 (O_803,N_13789,N_14940);
or UO_804 (O_804,N_13667,N_14211);
nor UO_805 (O_805,N_14987,N_14999);
and UO_806 (O_806,N_14327,N_14968);
nand UO_807 (O_807,N_14227,N_13933);
nor UO_808 (O_808,N_13944,N_14355);
and UO_809 (O_809,N_14202,N_14972);
nand UO_810 (O_810,N_13744,N_13670);
or UO_811 (O_811,N_14728,N_13802);
or UO_812 (O_812,N_14500,N_14319);
nand UO_813 (O_813,N_14569,N_14648);
nand UO_814 (O_814,N_14546,N_14130);
xnor UO_815 (O_815,N_13570,N_14594);
nor UO_816 (O_816,N_14119,N_14470);
nor UO_817 (O_817,N_13991,N_13621);
and UO_818 (O_818,N_14465,N_14592);
xor UO_819 (O_819,N_14228,N_13850);
or UO_820 (O_820,N_14389,N_14813);
nor UO_821 (O_821,N_14517,N_14231);
xnor UO_822 (O_822,N_14611,N_14637);
or UO_823 (O_823,N_14846,N_14404);
or UO_824 (O_824,N_14113,N_14338);
and UO_825 (O_825,N_14501,N_14091);
or UO_826 (O_826,N_14726,N_13701);
nand UO_827 (O_827,N_14525,N_14632);
nand UO_828 (O_828,N_14973,N_13749);
nand UO_829 (O_829,N_14484,N_14561);
and UO_830 (O_830,N_14107,N_14269);
and UO_831 (O_831,N_14349,N_14804);
nand UO_832 (O_832,N_14685,N_14814);
nor UO_833 (O_833,N_13945,N_13769);
xnor UO_834 (O_834,N_14187,N_14726);
or UO_835 (O_835,N_14160,N_14215);
nand UO_836 (O_836,N_14143,N_14669);
and UO_837 (O_837,N_14718,N_13909);
nand UO_838 (O_838,N_14012,N_14133);
and UO_839 (O_839,N_14684,N_13824);
or UO_840 (O_840,N_13582,N_14843);
xor UO_841 (O_841,N_14406,N_14620);
xor UO_842 (O_842,N_14908,N_14926);
xor UO_843 (O_843,N_13508,N_13637);
nand UO_844 (O_844,N_14997,N_14345);
or UO_845 (O_845,N_14073,N_14084);
or UO_846 (O_846,N_14195,N_14639);
nor UO_847 (O_847,N_13936,N_14970);
nor UO_848 (O_848,N_14243,N_14213);
and UO_849 (O_849,N_14991,N_14945);
and UO_850 (O_850,N_14347,N_13678);
xor UO_851 (O_851,N_14867,N_13959);
xnor UO_852 (O_852,N_14627,N_14027);
nor UO_853 (O_853,N_14626,N_13826);
or UO_854 (O_854,N_13780,N_14596);
nand UO_855 (O_855,N_14076,N_13739);
or UO_856 (O_856,N_13530,N_14734);
and UO_857 (O_857,N_14102,N_14186);
or UO_858 (O_858,N_13784,N_14272);
or UO_859 (O_859,N_13788,N_13925);
and UO_860 (O_860,N_14139,N_14541);
nor UO_861 (O_861,N_14279,N_13918);
nor UO_862 (O_862,N_13729,N_14772);
xor UO_863 (O_863,N_14752,N_14859);
xor UO_864 (O_864,N_14110,N_14381);
xor UO_865 (O_865,N_13877,N_14862);
nand UO_866 (O_866,N_13988,N_14087);
or UO_867 (O_867,N_14246,N_14867);
xnor UO_868 (O_868,N_14286,N_14025);
nor UO_869 (O_869,N_14461,N_14910);
xnor UO_870 (O_870,N_14785,N_14128);
or UO_871 (O_871,N_14707,N_14587);
or UO_872 (O_872,N_13845,N_14892);
and UO_873 (O_873,N_14709,N_14297);
nor UO_874 (O_874,N_14537,N_13783);
nand UO_875 (O_875,N_14868,N_14177);
or UO_876 (O_876,N_14338,N_14106);
nand UO_877 (O_877,N_14935,N_13556);
xnor UO_878 (O_878,N_13502,N_14147);
nand UO_879 (O_879,N_14643,N_13639);
nand UO_880 (O_880,N_14908,N_14408);
nor UO_881 (O_881,N_14892,N_14602);
xnor UO_882 (O_882,N_14780,N_14662);
xor UO_883 (O_883,N_14186,N_13763);
nor UO_884 (O_884,N_13507,N_13987);
nand UO_885 (O_885,N_14946,N_13618);
nor UO_886 (O_886,N_13740,N_14842);
nand UO_887 (O_887,N_14911,N_13603);
nand UO_888 (O_888,N_14493,N_13751);
xor UO_889 (O_889,N_14256,N_14870);
nor UO_890 (O_890,N_14941,N_14570);
xnor UO_891 (O_891,N_13942,N_13992);
and UO_892 (O_892,N_14221,N_13992);
or UO_893 (O_893,N_13618,N_14835);
xnor UO_894 (O_894,N_14316,N_13981);
and UO_895 (O_895,N_14035,N_14009);
nand UO_896 (O_896,N_14978,N_13740);
nand UO_897 (O_897,N_13878,N_14273);
nor UO_898 (O_898,N_13686,N_13627);
nand UO_899 (O_899,N_14479,N_14316);
or UO_900 (O_900,N_14290,N_13878);
nand UO_901 (O_901,N_13894,N_13995);
or UO_902 (O_902,N_13967,N_14396);
xnor UO_903 (O_903,N_14012,N_14648);
xnor UO_904 (O_904,N_14340,N_13993);
and UO_905 (O_905,N_13855,N_14210);
and UO_906 (O_906,N_14728,N_13713);
or UO_907 (O_907,N_13818,N_14516);
or UO_908 (O_908,N_13853,N_13989);
nor UO_909 (O_909,N_13751,N_13916);
nor UO_910 (O_910,N_13588,N_14526);
nor UO_911 (O_911,N_14217,N_14657);
and UO_912 (O_912,N_13686,N_13866);
nor UO_913 (O_913,N_14898,N_14423);
nor UO_914 (O_914,N_14915,N_13523);
or UO_915 (O_915,N_14984,N_14526);
nor UO_916 (O_916,N_14828,N_14502);
xnor UO_917 (O_917,N_14236,N_13836);
nor UO_918 (O_918,N_14876,N_14018);
and UO_919 (O_919,N_14671,N_14257);
or UO_920 (O_920,N_14058,N_14241);
or UO_921 (O_921,N_14240,N_14455);
and UO_922 (O_922,N_13775,N_13538);
xor UO_923 (O_923,N_13516,N_13613);
xor UO_924 (O_924,N_14999,N_14819);
xor UO_925 (O_925,N_14418,N_14984);
and UO_926 (O_926,N_14782,N_13504);
or UO_927 (O_927,N_14907,N_14786);
and UO_928 (O_928,N_13681,N_14102);
or UO_929 (O_929,N_13624,N_14983);
nand UO_930 (O_930,N_13888,N_14644);
nor UO_931 (O_931,N_14473,N_14088);
xor UO_932 (O_932,N_14610,N_13602);
xnor UO_933 (O_933,N_14564,N_14409);
nor UO_934 (O_934,N_13514,N_14490);
and UO_935 (O_935,N_14984,N_13626);
and UO_936 (O_936,N_14079,N_14705);
nand UO_937 (O_937,N_14292,N_14229);
or UO_938 (O_938,N_13969,N_14831);
and UO_939 (O_939,N_13801,N_14874);
nor UO_940 (O_940,N_13533,N_13797);
nor UO_941 (O_941,N_13980,N_13707);
xnor UO_942 (O_942,N_14888,N_13633);
or UO_943 (O_943,N_14971,N_14092);
and UO_944 (O_944,N_14991,N_13623);
nor UO_945 (O_945,N_13819,N_13923);
nor UO_946 (O_946,N_14016,N_13615);
and UO_947 (O_947,N_14870,N_14623);
and UO_948 (O_948,N_14224,N_14351);
xor UO_949 (O_949,N_14661,N_14383);
xnor UO_950 (O_950,N_14707,N_13980);
and UO_951 (O_951,N_13716,N_14907);
or UO_952 (O_952,N_14917,N_13996);
nand UO_953 (O_953,N_14924,N_14032);
xor UO_954 (O_954,N_14510,N_14880);
nand UO_955 (O_955,N_14105,N_14050);
or UO_956 (O_956,N_13828,N_14574);
or UO_957 (O_957,N_14711,N_14461);
xnor UO_958 (O_958,N_13779,N_14990);
or UO_959 (O_959,N_13578,N_14233);
and UO_960 (O_960,N_14867,N_14750);
nand UO_961 (O_961,N_13607,N_14996);
or UO_962 (O_962,N_13958,N_13678);
or UO_963 (O_963,N_14731,N_14161);
xor UO_964 (O_964,N_14104,N_14952);
xnor UO_965 (O_965,N_14927,N_13638);
xnor UO_966 (O_966,N_14140,N_14262);
nor UO_967 (O_967,N_14853,N_14883);
nand UO_968 (O_968,N_14605,N_14451);
nand UO_969 (O_969,N_14642,N_13851);
and UO_970 (O_970,N_13561,N_13987);
or UO_971 (O_971,N_13802,N_14376);
and UO_972 (O_972,N_13860,N_14151);
and UO_973 (O_973,N_14204,N_14234);
and UO_974 (O_974,N_13686,N_14886);
nand UO_975 (O_975,N_13750,N_13597);
and UO_976 (O_976,N_13505,N_13631);
xor UO_977 (O_977,N_14310,N_14695);
nand UO_978 (O_978,N_14544,N_14493);
and UO_979 (O_979,N_14754,N_14724);
xor UO_980 (O_980,N_14593,N_13788);
nor UO_981 (O_981,N_14667,N_13920);
xnor UO_982 (O_982,N_14457,N_13823);
nand UO_983 (O_983,N_13608,N_14897);
xor UO_984 (O_984,N_13527,N_13711);
or UO_985 (O_985,N_14879,N_13702);
nand UO_986 (O_986,N_14211,N_14742);
or UO_987 (O_987,N_14130,N_14998);
or UO_988 (O_988,N_13737,N_14801);
nand UO_989 (O_989,N_14361,N_14994);
xor UO_990 (O_990,N_14145,N_13857);
nand UO_991 (O_991,N_14201,N_13732);
and UO_992 (O_992,N_14159,N_14969);
nand UO_993 (O_993,N_13811,N_13726);
nor UO_994 (O_994,N_14137,N_14231);
xor UO_995 (O_995,N_13590,N_14891);
xnor UO_996 (O_996,N_14013,N_14028);
or UO_997 (O_997,N_13761,N_14489);
xor UO_998 (O_998,N_14943,N_14304);
nor UO_999 (O_999,N_13892,N_14688);
nor UO_1000 (O_1000,N_14209,N_14073);
xnor UO_1001 (O_1001,N_14037,N_13803);
nor UO_1002 (O_1002,N_14358,N_14684);
xnor UO_1003 (O_1003,N_13729,N_14994);
xor UO_1004 (O_1004,N_13673,N_13873);
xor UO_1005 (O_1005,N_14967,N_13889);
xnor UO_1006 (O_1006,N_14687,N_13789);
nor UO_1007 (O_1007,N_14854,N_14875);
nand UO_1008 (O_1008,N_14413,N_14396);
xor UO_1009 (O_1009,N_14537,N_14602);
nand UO_1010 (O_1010,N_13980,N_13990);
xor UO_1011 (O_1011,N_13523,N_14090);
or UO_1012 (O_1012,N_14323,N_14381);
and UO_1013 (O_1013,N_14542,N_14134);
and UO_1014 (O_1014,N_13773,N_14662);
or UO_1015 (O_1015,N_13810,N_14249);
and UO_1016 (O_1016,N_14620,N_13887);
or UO_1017 (O_1017,N_14061,N_13676);
or UO_1018 (O_1018,N_14570,N_14730);
or UO_1019 (O_1019,N_13677,N_14616);
nor UO_1020 (O_1020,N_14199,N_13633);
xnor UO_1021 (O_1021,N_14235,N_13680);
nor UO_1022 (O_1022,N_14323,N_14453);
xor UO_1023 (O_1023,N_14415,N_14180);
or UO_1024 (O_1024,N_14668,N_14936);
nand UO_1025 (O_1025,N_14744,N_14245);
and UO_1026 (O_1026,N_13799,N_14190);
and UO_1027 (O_1027,N_14362,N_14876);
nor UO_1028 (O_1028,N_13870,N_13678);
nand UO_1029 (O_1029,N_14427,N_13536);
nand UO_1030 (O_1030,N_13598,N_14419);
xor UO_1031 (O_1031,N_14360,N_14833);
nor UO_1032 (O_1032,N_14763,N_13874);
nor UO_1033 (O_1033,N_14413,N_14218);
or UO_1034 (O_1034,N_14007,N_14016);
nand UO_1035 (O_1035,N_14018,N_13664);
xor UO_1036 (O_1036,N_14210,N_13747);
nor UO_1037 (O_1037,N_13526,N_13656);
nor UO_1038 (O_1038,N_14502,N_13790);
or UO_1039 (O_1039,N_14447,N_14819);
or UO_1040 (O_1040,N_14212,N_13766);
nand UO_1041 (O_1041,N_13914,N_14541);
xnor UO_1042 (O_1042,N_14956,N_13982);
nand UO_1043 (O_1043,N_14970,N_14168);
nand UO_1044 (O_1044,N_14089,N_13824);
and UO_1045 (O_1045,N_14494,N_14896);
or UO_1046 (O_1046,N_14324,N_14338);
xnor UO_1047 (O_1047,N_13607,N_14231);
and UO_1048 (O_1048,N_13524,N_13802);
or UO_1049 (O_1049,N_14814,N_14884);
nor UO_1050 (O_1050,N_14105,N_13604);
xor UO_1051 (O_1051,N_13701,N_13952);
xnor UO_1052 (O_1052,N_14766,N_13696);
xor UO_1053 (O_1053,N_14634,N_14423);
nor UO_1054 (O_1054,N_14142,N_13778);
nor UO_1055 (O_1055,N_14109,N_13649);
nand UO_1056 (O_1056,N_14638,N_13535);
nor UO_1057 (O_1057,N_14853,N_14274);
xnor UO_1058 (O_1058,N_14526,N_14976);
nand UO_1059 (O_1059,N_14997,N_14077);
or UO_1060 (O_1060,N_14388,N_14990);
nand UO_1061 (O_1061,N_14797,N_14569);
nand UO_1062 (O_1062,N_14412,N_14735);
and UO_1063 (O_1063,N_14683,N_14399);
or UO_1064 (O_1064,N_14353,N_14304);
nor UO_1065 (O_1065,N_14629,N_14455);
or UO_1066 (O_1066,N_14860,N_13659);
nor UO_1067 (O_1067,N_13579,N_14312);
and UO_1068 (O_1068,N_13823,N_14134);
nand UO_1069 (O_1069,N_14503,N_13880);
and UO_1070 (O_1070,N_14062,N_13902);
and UO_1071 (O_1071,N_13813,N_13745);
or UO_1072 (O_1072,N_14600,N_14734);
nor UO_1073 (O_1073,N_14857,N_14121);
or UO_1074 (O_1074,N_14698,N_14937);
and UO_1075 (O_1075,N_14516,N_13693);
or UO_1076 (O_1076,N_13714,N_14275);
nand UO_1077 (O_1077,N_14061,N_14376);
nand UO_1078 (O_1078,N_13760,N_14195);
and UO_1079 (O_1079,N_14424,N_14075);
or UO_1080 (O_1080,N_13662,N_14571);
nor UO_1081 (O_1081,N_13599,N_13762);
nor UO_1082 (O_1082,N_13949,N_13782);
xnor UO_1083 (O_1083,N_13584,N_13855);
nor UO_1084 (O_1084,N_14880,N_13625);
nand UO_1085 (O_1085,N_14570,N_13508);
nand UO_1086 (O_1086,N_14491,N_14349);
nand UO_1087 (O_1087,N_13575,N_13542);
nand UO_1088 (O_1088,N_13501,N_14272);
nor UO_1089 (O_1089,N_14292,N_14193);
xnor UO_1090 (O_1090,N_14746,N_13668);
or UO_1091 (O_1091,N_14916,N_14919);
or UO_1092 (O_1092,N_14860,N_14202);
nor UO_1093 (O_1093,N_14545,N_14509);
and UO_1094 (O_1094,N_13502,N_14024);
xnor UO_1095 (O_1095,N_13714,N_14261);
and UO_1096 (O_1096,N_14841,N_13570);
xnor UO_1097 (O_1097,N_13985,N_14360);
nand UO_1098 (O_1098,N_14691,N_14278);
nor UO_1099 (O_1099,N_13952,N_14425);
nand UO_1100 (O_1100,N_14932,N_13984);
xnor UO_1101 (O_1101,N_14663,N_14695);
nor UO_1102 (O_1102,N_14956,N_14869);
or UO_1103 (O_1103,N_14747,N_13952);
and UO_1104 (O_1104,N_14616,N_14911);
nor UO_1105 (O_1105,N_13984,N_14655);
nand UO_1106 (O_1106,N_14510,N_14910);
nor UO_1107 (O_1107,N_14338,N_14423);
nand UO_1108 (O_1108,N_14293,N_14361);
xnor UO_1109 (O_1109,N_13886,N_14233);
xnor UO_1110 (O_1110,N_13892,N_13561);
nand UO_1111 (O_1111,N_13634,N_14918);
xor UO_1112 (O_1112,N_14688,N_13788);
or UO_1113 (O_1113,N_14591,N_14530);
nor UO_1114 (O_1114,N_13806,N_13567);
nor UO_1115 (O_1115,N_13578,N_14185);
or UO_1116 (O_1116,N_14789,N_13778);
or UO_1117 (O_1117,N_14228,N_14775);
xnor UO_1118 (O_1118,N_13961,N_14920);
nor UO_1119 (O_1119,N_13750,N_14064);
and UO_1120 (O_1120,N_14661,N_14646);
nand UO_1121 (O_1121,N_14292,N_14230);
and UO_1122 (O_1122,N_13700,N_14931);
nand UO_1123 (O_1123,N_13989,N_14391);
nand UO_1124 (O_1124,N_13576,N_14055);
xor UO_1125 (O_1125,N_14292,N_13843);
xnor UO_1126 (O_1126,N_14831,N_13574);
nand UO_1127 (O_1127,N_14314,N_13756);
xnor UO_1128 (O_1128,N_13755,N_14778);
nor UO_1129 (O_1129,N_13974,N_14474);
and UO_1130 (O_1130,N_14527,N_14034);
or UO_1131 (O_1131,N_14665,N_13548);
xnor UO_1132 (O_1132,N_14978,N_14774);
xnor UO_1133 (O_1133,N_14649,N_14154);
xnor UO_1134 (O_1134,N_14175,N_13701);
and UO_1135 (O_1135,N_14040,N_14135);
xnor UO_1136 (O_1136,N_13567,N_14796);
and UO_1137 (O_1137,N_13762,N_13867);
xnor UO_1138 (O_1138,N_13558,N_13944);
nor UO_1139 (O_1139,N_14950,N_14031);
nand UO_1140 (O_1140,N_14499,N_13992);
nor UO_1141 (O_1141,N_14784,N_14936);
nor UO_1142 (O_1142,N_14558,N_14103);
and UO_1143 (O_1143,N_13885,N_14798);
nand UO_1144 (O_1144,N_14228,N_13500);
or UO_1145 (O_1145,N_13534,N_14877);
xor UO_1146 (O_1146,N_14889,N_13723);
xnor UO_1147 (O_1147,N_13778,N_13813);
nor UO_1148 (O_1148,N_14715,N_14859);
nand UO_1149 (O_1149,N_14837,N_14429);
nand UO_1150 (O_1150,N_13778,N_13868);
xnor UO_1151 (O_1151,N_14291,N_14031);
and UO_1152 (O_1152,N_13934,N_13955);
nand UO_1153 (O_1153,N_13622,N_14330);
xnor UO_1154 (O_1154,N_14618,N_13572);
nor UO_1155 (O_1155,N_14874,N_14231);
nor UO_1156 (O_1156,N_14131,N_14586);
and UO_1157 (O_1157,N_14456,N_13725);
and UO_1158 (O_1158,N_14211,N_13703);
and UO_1159 (O_1159,N_13724,N_14328);
nand UO_1160 (O_1160,N_13652,N_14840);
nor UO_1161 (O_1161,N_14299,N_13772);
xnor UO_1162 (O_1162,N_14409,N_14823);
nand UO_1163 (O_1163,N_14734,N_13931);
nand UO_1164 (O_1164,N_13752,N_13771);
nor UO_1165 (O_1165,N_14390,N_14356);
or UO_1166 (O_1166,N_13564,N_14230);
xnor UO_1167 (O_1167,N_14883,N_13668);
xnor UO_1168 (O_1168,N_14860,N_14264);
nand UO_1169 (O_1169,N_13810,N_14912);
xor UO_1170 (O_1170,N_13672,N_14479);
and UO_1171 (O_1171,N_14807,N_14125);
nand UO_1172 (O_1172,N_14844,N_13706);
and UO_1173 (O_1173,N_14597,N_13582);
nand UO_1174 (O_1174,N_14274,N_13590);
xnor UO_1175 (O_1175,N_14692,N_14979);
nand UO_1176 (O_1176,N_13587,N_14843);
nand UO_1177 (O_1177,N_13974,N_13950);
xor UO_1178 (O_1178,N_14119,N_14050);
and UO_1179 (O_1179,N_14340,N_14710);
xnor UO_1180 (O_1180,N_14529,N_14175);
nand UO_1181 (O_1181,N_14013,N_14292);
nor UO_1182 (O_1182,N_13503,N_14055);
xnor UO_1183 (O_1183,N_14615,N_13723);
xor UO_1184 (O_1184,N_14292,N_13782);
and UO_1185 (O_1185,N_14764,N_14895);
nor UO_1186 (O_1186,N_14023,N_14415);
xor UO_1187 (O_1187,N_14779,N_14768);
xor UO_1188 (O_1188,N_14148,N_14442);
and UO_1189 (O_1189,N_14971,N_14423);
nand UO_1190 (O_1190,N_13526,N_13893);
or UO_1191 (O_1191,N_13568,N_14467);
and UO_1192 (O_1192,N_14697,N_14599);
or UO_1193 (O_1193,N_13732,N_14363);
nor UO_1194 (O_1194,N_13807,N_13778);
nand UO_1195 (O_1195,N_13500,N_13794);
xor UO_1196 (O_1196,N_14120,N_14677);
xor UO_1197 (O_1197,N_14663,N_14048);
xnor UO_1198 (O_1198,N_14956,N_14880);
nor UO_1199 (O_1199,N_14373,N_14202);
nand UO_1200 (O_1200,N_14331,N_13909);
or UO_1201 (O_1201,N_13798,N_13922);
and UO_1202 (O_1202,N_13674,N_13732);
nor UO_1203 (O_1203,N_13675,N_13574);
nand UO_1204 (O_1204,N_14344,N_14815);
and UO_1205 (O_1205,N_13746,N_14972);
nor UO_1206 (O_1206,N_14231,N_14861);
or UO_1207 (O_1207,N_13751,N_14205);
and UO_1208 (O_1208,N_13819,N_14457);
or UO_1209 (O_1209,N_13953,N_14964);
xor UO_1210 (O_1210,N_14745,N_14330);
or UO_1211 (O_1211,N_14246,N_14905);
nand UO_1212 (O_1212,N_13528,N_13648);
nand UO_1213 (O_1213,N_14139,N_13547);
nand UO_1214 (O_1214,N_14582,N_14802);
and UO_1215 (O_1215,N_14934,N_14583);
nand UO_1216 (O_1216,N_14200,N_14064);
and UO_1217 (O_1217,N_14838,N_14527);
nor UO_1218 (O_1218,N_14548,N_14949);
and UO_1219 (O_1219,N_14789,N_14949);
nor UO_1220 (O_1220,N_14085,N_14453);
xor UO_1221 (O_1221,N_14148,N_14514);
nand UO_1222 (O_1222,N_14680,N_14568);
xor UO_1223 (O_1223,N_14553,N_13941);
xnor UO_1224 (O_1224,N_14340,N_13523);
nand UO_1225 (O_1225,N_14392,N_14506);
or UO_1226 (O_1226,N_13840,N_13704);
or UO_1227 (O_1227,N_14952,N_14012);
nor UO_1228 (O_1228,N_13952,N_14843);
nor UO_1229 (O_1229,N_14255,N_14589);
nand UO_1230 (O_1230,N_14659,N_14976);
xnor UO_1231 (O_1231,N_14042,N_14692);
or UO_1232 (O_1232,N_14912,N_14589);
nor UO_1233 (O_1233,N_13926,N_14949);
or UO_1234 (O_1234,N_14373,N_14779);
and UO_1235 (O_1235,N_14811,N_14203);
nand UO_1236 (O_1236,N_14128,N_13564);
nand UO_1237 (O_1237,N_13641,N_13854);
or UO_1238 (O_1238,N_14529,N_14667);
nor UO_1239 (O_1239,N_14163,N_14088);
and UO_1240 (O_1240,N_14830,N_14800);
nand UO_1241 (O_1241,N_14934,N_14654);
nor UO_1242 (O_1242,N_13859,N_14013);
xnor UO_1243 (O_1243,N_14142,N_14245);
or UO_1244 (O_1244,N_14956,N_13612);
xor UO_1245 (O_1245,N_14148,N_14902);
or UO_1246 (O_1246,N_13543,N_13868);
or UO_1247 (O_1247,N_14939,N_13907);
nand UO_1248 (O_1248,N_14708,N_13708);
xor UO_1249 (O_1249,N_14764,N_14122);
or UO_1250 (O_1250,N_13681,N_13711);
and UO_1251 (O_1251,N_13653,N_14129);
xnor UO_1252 (O_1252,N_13717,N_13914);
nor UO_1253 (O_1253,N_14819,N_14704);
nor UO_1254 (O_1254,N_13740,N_14640);
xor UO_1255 (O_1255,N_14771,N_14077);
or UO_1256 (O_1256,N_14453,N_14667);
nor UO_1257 (O_1257,N_13747,N_13852);
nor UO_1258 (O_1258,N_13649,N_14330);
nand UO_1259 (O_1259,N_13574,N_13577);
or UO_1260 (O_1260,N_14586,N_13928);
and UO_1261 (O_1261,N_14225,N_14859);
or UO_1262 (O_1262,N_13731,N_14937);
and UO_1263 (O_1263,N_14112,N_14487);
and UO_1264 (O_1264,N_13746,N_14441);
or UO_1265 (O_1265,N_14396,N_14927);
and UO_1266 (O_1266,N_14062,N_14561);
or UO_1267 (O_1267,N_13843,N_14778);
or UO_1268 (O_1268,N_14278,N_14676);
nor UO_1269 (O_1269,N_14421,N_13512);
nor UO_1270 (O_1270,N_14672,N_14184);
or UO_1271 (O_1271,N_13643,N_14664);
nand UO_1272 (O_1272,N_14948,N_14018);
or UO_1273 (O_1273,N_14145,N_13640);
and UO_1274 (O_1274,N_14499,N_14745);
and UO_1275 (O_1275,N_14125,N_14518);
xnor UO_1276 (O_1276,N_14627,N_14592);
nor UO_1277 (O_1277,N_14174,N_14800);
nand UO_1278 (O_1278,N_14062,N_13779);
nor UO_1279 (O_1279,N_14238,N_14953);
xnor UO_1280 (O_1280,N_14814,N_14902);
and UO_1281 (O_1281,N_14352,N_13837);
nor UO_1282 (O_1282,N_13866,N_14382);
and UO_1283 (O_1283,N_13802,N_14099);
and UO_1284 (O_1284,N_14577,N_14385);
xnor UO_1285 (O_1285,N_14155,N_13792);
and UO_1286 (O_1286,N_14135,N_13524);
nand UO_1287 (O_1287,N_14602,N_14497);
or UO_1288 (O_1288,N_14311,N_13728);
nor UO_1289 (O_1289,N_14011,N_14085);
or UO_1290 (O_1290,N_13520,N_14192);
and UO_1291 (O_1291,N_13840,N_13755);
nor UO_1292 (O_1292,N_14496,N_14609);
nor UO_1293 (O_1293,N_13909,N_14610);
or UO_1294 (O_1294,N_13615,N_13639);
nand UO_1295 (O_1295,N_14153,N_14372);
xor UO_1296 (O_1296,N_13664,N_14438);
and UO_1297 (O_1297,N_14082,N_14839);
xnor UO_1298 (O_1298,N_14282,N_13570);
xor UO_1299 (O_1299,N_13625,N_14175);
and UO_1300 (O_1300,N_14185,N_14107);
nor UO_1301 (O_1301,N_14723,N_14907);
or UO_1302 (O_1302,N_13783,N_14092);
and UO_1303 (O_1303,N_14138,N_14029);
nor UO_1304 (O_1304,N_13878,N_14939);
or UO_1305 (O_1305,N_14571,N_13915);
xnor UO_1306 (O_1306,N_14643,N_13721);
and UO_1307 (O_1307,N_13866,N_14170);
nand UO_1308 (O_1308,N_14354,N_14894);
nor UO_1309 (O_1309,N_13625,N_14024);
and UO_1310 (O_1310,N_14924,N_13502);
nand UO_1311 (O_1311,N_14247,N_14777);
nand UO_1312 (O_1312,N_13550,N_13812);
xnor UO_1313 (O_1313,N_14712,N_14803);
nor UO_1314 (O_1314,N_14517,N_13639);
and UO_1315 (O_1315,N_14891,N_14421);
nor UO_1316 (O_1316,N_13559,N_13617);
xor UO_1317 (O_1317,N_14861,N_13724);
xor UO_1318 (O_1318,N_14951,N_14771);
xor UO_1319 (O_1319,N_13925,N_14487);
xor UO_1320 (O_1320,N_14452,N_13925);
nand UO_1321 (O_1321,N_14425,N_13545);
or UO_1322 (O_1322,N_14475,N_13560);
nor UO_1323 (O_1323,N_14646,N_14653);
nand UO_1324 (O_1324,N_14828,N_14884);
and UO_1325 (O_1325,N_14575,N_14053);
nor UO_1326 (O_1326,N_13793,N_13765);
xnor UO_1327 (O_1327,N_14630,N_14762);
nor UO_1328 (O_1328,N_14832,N_14327);
nand UO_1329 (O_1329,N_13530,N_14912);
xnor UO_1330 (O_1330,N_13789,N_14171);
nand UO_1331 (O_1331,N_14154,N_13555);
or UO_1332 (O_1332,N_14163,N_13500);
nor UO_1333 (O_1333,N_14355,N_14506);
and UO_1334 (O_1334,N_14320,N_14459);
xnor UO_1335 (O_1335,N_13647,N_14976);
xor UO_1336 (O_1336,N_14018,N_14572);
or UO_1337 (O_1337,N_14118,N_13767);
or UO_1338 (O_1338,N_13947,N_13517);
nor UO_1339 (O_1339,N_13877,N_14390);
nor UO_1340 (O_1340,N_14405,N_14261);
nor UO_1341 (O_1341,N_13557,N_13949);
xor UO_1342 (O_1342,N_14428,N_14401);
xor UO_1343 (O_1343,N_14759,N_14175);
nor UO_1344 (O_1344,N_13836,N_13989);
nand UO_1345 (O_1345,N_14606,N_14328);
and UO_1346 (O_1346,N_14463,N_14130);
nor UO_1347 (O_1347,N_13716,N_13845);
or UO_1348 (O_1348,N_14649,N_13666);
nor UO_1349 (O_1349,N_14715,N_14245);
nor UO_1350 (O_1350,N_14699,N_14772);
xnor UO_1351 (O_1351,N_13788,N_14372);
or UO_1352 (O_1352,N_14515,N_14517);
and UO_1353 (O_1353,N_14969,N_14544);
and UO_1354 (O_1354,N_14933,N_14397);
or UO_1355 (O_1355,N_14519,N_14963);
xnor UO_1356 (O_1356,N_14011,N_14953);
nor UO_1357 (O_1357,N_14436,N_14053);
xor UO_1358 (O_1358,N_14768,N_14594);
xnor UO_1359 (O_1359,N_13905,N_14569);
and UO_1360 (O_1360,N_14380,N_14346);
nor UO_1361 (O_1361,N_14801,N_13967);
nand UO_1362 (O_1362,N_14260,N_13624);
nand UO_1363 (O_1363,N_14738,N_13575);
nor UO_1364 (O_1364,N_14662,N_14999);
nand UO_1365 (O_1365,N_14213,N_14582);
xor UO_1366 (O_1366,N_14201,N_13529);
or UO_1367 (O_1367,N_14612,N_13868);
nand UO_1368 (O_1368,N_13795,N_14373);
and UO_1369 (O_1369,N_13941,N_13730);
nor UO_1370 (O_1370,N_13919,N_13512);
nor UO_1371 (O_1371,N_14904,N_14834);
nor UO_1372 (O_1372,N_14873,N_14070);
and UO_1373 (O_1373,N_13584,N_14998);
nor UO_1374 (O_1374,N_13784,N_14972);
nor UO_1375 (O_1375,N_13664,N_14356);
nor UO_1376 (O_1376,N_14836,N_14875);
xnor UO_1377 (O_1377,N_14783,N_13774);
or UO_1378 (O_1378,N_14357,N_14480);
nor UO_1379 (O_1379,N_14000,N_14504);
nor UO_1380 (O_1380,N_14065,N_13638);
and UO_1381 (O_1381,N_14272,N_14192);
nand UO_1382 (O_1382,N_14427,N_14396);
nor UO_1383 (O_1383,N_14080,N_13625);
nand UO_1384 (O_1384,N_14538,N_14849);
xnor UO_1385 (O_1385,N_14686,N_14704);
xor UO_1386 (O_1386,N_14462,N_13652);
xor UO_1387 (O_1387,N_14285,N_13897);
xnor UO_1388 (O_1388,N_14441,N_13901);
and UO_1389 (O_1389,N_14712,N_14742);
or UO_1390 (O_1390,N_13885,N_13993);
nor UO_1391 (O_1391,N_14109,N_13689);
nand UO_1392 (O_1392,N_14373,N_13987);
or UO_1393 (O_1393,N_13982,N_14742);
nor UO_1394 (O_1394,N_14247,N_14505);
nor UO_1395 (O_1395,N_13528,N_14167);
and UO_1396 (O_1396,N_13534,N_14420);
or UO_1397 (O_1397,N_13818,N_14913);
nand UO_1398 (O_1398,N_14773,N_14806);
and UO_1399 (O_1399,N_13683,N_14187);
and UO_1400 (O_1400,N_13835,N_13548);
and UO_1401 (O_1401,N_14774,N_14198);
xor UO_1402 (O_1402,N_14984,N_14699);
nor UO_1403 (O_1403,N_14865,N_13665);
and UO_1404 (O_1404,N_14273,N_14058);
nand UO_1405 (O_1405,N_14867,N_13583);
nand UO_1406 (O_1406,N_13979,N_13820);
nand UO_1407 (O_1407,N_14323,N_13811);
nor UO_1408 (O_1408,N_14233,N_14222);
or UO_1409 (O_1409,N_14149,N_13844);
nor UO_1410 (O_1410,N_14312,N_14230);
or UO_1411 (O_1411,N_14060,N_13975);
xor UO_1412 (O_1412,N_14392,N_14013);
xor UO_1413 (O_1413,N_13866,N_14985);
or UO_1414 (O_1414,N_13743,N_13930);
nand UO_1415 (O_1415,N_14038,N_13944);
and UO_1416 (O_1416,N_13861,N_13971);
nand UO_1417 (O_1417,N_14180,N_13744);
nor UO_1418 (O_1418,N_14285,N_14572);
or UO_1419 (O_1419,N_13519,N_14171);
or UO_1420 (O_1420,N_14042,N_14377);
nand UO_1421 (O_1421,N_13950,N_13930);
nor UO_1422 (O_1422,N_14735,N_14282);
nor UO_1423 (O_1423,N_14501,N_14301);
nor UO_1424 (O_1424,N_14120,N_13680);
xnor UO_1425 (O_1425,N_14929,N_14772);
xnor UO_1426 (O_1426,N_13885,N_14997);
or UO_1427 (O_1427,N_13578,N_14600);
xnor UO_1428 (O_1428,N_14682,N_14376);
nor UO_1429 (O_1429,N_13507,N_13830);
nor UO_1430 (O_1430,N_14921,N_13642);
nor UO_1431 (O_1431,N_13961,N_14832);
or UO_1432 (O_1432,N_14554,N_13986);
or UO_1433 (O_1433,N_14940,N_14067);
nand UO_1434 (O_1434,N_13547,N_13645);
and UO_1435 (O_1435,N_13582,N_13530);
nand UO_1436 (O_1436,N_14152,N_14600);
or UO_1437 (O_1437,N_14140,N_13566);
or UO_1438 (O_1438,N_14164,N_13518);
and UO_1439 (O_1439,N_13644,N_14458);
xnor UO_1440 (O_1440,N_14010,N_13626);
and UO_1441 (O_1441,N_14435,N_13676);
nor UO_1442 (O_1442,N_13934,N_14013);
or UO_1443 (O_1443,N_13987,N_14703);
or UO_1444 (O_1444,N_13622,N_14683);
nand UO_1445 (O_1445,N_14127,N_13823);
or UO_1446 (O_1446,N_14500,N_14444);
xnor UO_1447 (O_1447,N_14262,N_13858);
nand UO_1448 (O_1448,N_14300,N_13592);
or UO_1449 (O_1449,N_14423,N_14978);
and UO_1450 (O_1450,N_14910,N_14505);
and UO_1451 (O_1451,N_13503,N_13614);
nor UO_1452 (O_1452,N_14210,N_14030);
or UO_1453 (O_1453,N_14060,N_14965);
or UO_1454 (O_1454,N_13712,N_14038);
nor UO_1455 (O_1455,N_14667,N_14991);
nand UO_1456 (O_1456,N_13972,N_13864);
and UO_1457 (O_1457,N_13814,N_14820);
and UO_1458 (O_1458,N_13576,N_14619);
and UO_1459 (O_1459,N_14372,N_13937);
nand UO_1460 (O_1460,N_13810,N_14784);
or UO_1461 (O_1461,N_14393,N_14380);
nand UO_1462 (O_1462,N_14835,N_14715);
nand UO_1463 (O_1463,N_14484,N_14517);
xnor UO_1464 (O_1464,N_13668,N_14535);
nand UO_1465 (O_1465,N_14857,N_13745);
and UO_1466 (O_1466,N_13659,N_14701);
nor UO_1467 (O_1467,N_13958,N_14818);
xor UO_1468 (O_1468,N_14610,N_14557);
or UO_1469 (O_1469,N_14400,N_14499);
or UO_1470 (O_1470,N_14720,N_14176);
nand UO_1471 (O_1471,N_13798,N_13752);
and UO_1472 (O_1472,N_13646,N_14561);
or UO_1473 (O_1473,N_13924,N_13735);
and UO_1474 (O_1474,N_14512,N_14643);
nand UO_1475 (O_1475,N_14369,N_13699);
nand UO_1476 (O_1476,N_14425,N_13523);
and UO_1477 (O_1477,N_14435,N_14167);
or UO_1478 (O_1478,N_14435,N_14128);
and UO_1479 (O_1479,N_13751,N_14906);
nand UO_1480 (O_1480,N_14944,N_14297);
nor UO_1481 (O_1481,N_14003,N_13542);
nor UO_1482 (O_1482,N_14703,N_14570);
and UO_1483 (O_1483,N_13743,N_13558);
and UO_1484 (O_1484,N_14384,N_14057);
nor UO_1485 (O_1485,N_14913,N_14967);
or UO_1486 (O_1486,N_14880,N_13805);
and UO_1487 (O_1487,N_14050,N_14301);
xor UO_1488 (O_1488,N_13728,N_14646);
or UO_1489 (O_1489,N_13545,N_14013);
nor UO_1490 (O_1490,N_14553,N_14067);
nor UO_1491 (O_1491,N_14447,N_14318);
nor UO_1492 (O_1492,N_14155,N_13881);
nand UO_1493 (O_1493,N_14312,N_14930);
and UO_1494 (O_1494,N_14586,N_14812);
xnor UO_1495 (O_1495,N_13699,N_13959);
nand UO_1496 (O_1496,N_14162,N_14653);
nand UO_1497 (O_1497,N_14044,N_14434);
nand UO_1498 (O_1498,N_14105,N_14540);
nor UO_1499 (O_1499,N_13683,N_14468);
and UO_1500 (O_1500,N_13897,N_14154);
nor UO_1501 (O_1501,N_14138,N_13658);
nor UO_1502 (O_1502,N_14608,N_13770);
nor UO_1503 (O_1503,N_13699,N_14769);
nor UO_1504 (O_1504,N_14133,N_13755);
nand UO_1505 (O_1505,N_13634,N_13835);
xor UO_1506 (O_1506,N_14693,N_13909);
or UO_1507 (O_1507,N_13787,N_14481);
or UO_1508 (O_1508,N_14216,N_13825);
or UO_1509 (O_1509,N_14148,N_14679);
nand UO_1510 (O_1510,N_13810,N_14873);
or UO_1511 (O_1511,N_13828,N_14953);
nor UO_1512 (O_1512,N_14799,N_14315);
nand UO_1513 (O_1513,N_14301,N_14300);
nand UO_1514 (O_1514,N_14930,N_14591);
nor UO_1515 (O_1515,N_14090,N_14081);
xnor UO_1516 (O_1516,N_14927,N_14700);
xor UO_1517 (O_1517,N_13730,N_13819);
xnor UO_1518 (O_1518,N_13949,N_14452);
and UO_1519 (O_1519,N_14273,N_14001);
and UO_1520 (O_1520,N_14380,N_14449);
nand UO_1521 (O_1521,N_13882,N_14447);
or UO_1522 (O_1522,N_14329,N_14102);
or UO_1523 (O_1523,N_14238,N_13684);
nand UO_1524 (O_1524,N_14686,N_14625);
nor UO_1525 (O_1525,N_13958,N_14540);
nor UO_1526 (O_1526,N_13888,N_14845);
nand UO_1527 (O_1527,N_14798,N_14221);
nor UO_1528 (O_1528,N_14118,N_13632);
or UO_1529 (O_1529,N_14169,N_14949);
and UO_1530 (O_1530,N_14258,N_13752);
xor UO_1531 (O_1531,N_14568,N_14400);
xor UO_1532 (O_1532,N_14168,N_14750);
or UO_1533 (O_1533,N_14295,N_14299);
nand UO_1534 (O_1534,N_14143,N_14963);
nor UO_1535 (O_1535,N_14836,N_13686);
nor UO_1536 (O_1536,N_14235,N_14411);
and UO_1537 (O_1537,N_14886,N_13838);
and UO_1538 (O_1538,N_14487,N_13789);
xor UO_1539 (O_1539,N_13662,N_14273);
and UO_1540 (O_1540,N_14660,N_13504);
or UO_1541 (O_1541,N_13740,N_14566);
nand UO_1542 (O_1542,N_13887,N_14948);
or UO_1543 (O_1543,N_13892,N_14005);
nand UO_1544 (O_1544,N_14883,N_14226);
xor UO_1545 (O_1545,N_13899,N_14192);
nand UO_1546 (O_1546,N_14774,N_14484);
and UO_1547 (O_1547,N_14054,N_13962);
nand UO_1548 (O_1548,N_13710,N_13696);
nand UO_1549 (O_1549,N_14330,N_14804);
and UO_1550 (O_1550,N_14446,N_14453);
or UO_1551 (O_1551,N_13960,N_14737);
or UO_1552 (O_1552,N_14256,N_13741);
or UO_1553 (O_1553,N_14982,N_13991);
or UO_1554 (O_1554,N_14847,N_14154);
nor UO_1555 (O_1555,N_14839,N_14093);
xor UO_1556 (O_1556,N_13604,N_13733);
nand UO_1557 (O_1557,N_14807,N_13648);
nor UO_1558 (O_1558,N_14735,N_14724);
nand UO_1559 (O_1559,N_14074,N_14753);
nor UO_1560 (O_1560,N_14783,N_13589);
nand UO_1561 (O_1561,N_14822,N_13865);
and UO_1562 (O_1562,N_14511,N_14838);
or UO_1563 (O_1563,N_13883,N_14694);
nor UO_1564 (O_1564,N_14453,N_14208);
xor UO_1565 (O_1565,N_14440,N_14005);
nor UO_1566 (O_1566,N_14929,N_13586);
nand UO_1567 (O_1567,N_13771,N_13794);
nor UO_1568 (O_1568,N_14115,N_14305);
nand UO_1569 (O_1569,N_14717,N_14564);
nand UO_1570 (O_1570,N_13934,N_13783);
nand UO_1571 (O_1571,N_13542,N_14082);
or UO_1572 (O_1572,N_14385,N_14831);
and UO_1573 (O_1573,N_14382,N_13624);
or UO_1574 (O_1574,N_14522,N_14320);
or UO_1575 (O_1575,N_14399,N_14203);
and UO_1576 (O_1576,N_14248,N_13905);
and UO_1577 (O_1577,N_14009,N_14582);
or UO_1578 (O_1578,N_14146,N_14391);
xor UO_1579 (O_1579,N_14746,N_14496);
or UO_1580 (O_1580,N_14477,N_14203);
xor UO_1581 (O_1581,N_13751,N_13647);
xor UO_1582 (O_1582,N_14740,N_14632);
or UO_1583 (O_1583,N_14561,N_14980);
nor UO_1584 (O_1584,N_14201,N_14370);
nor UO_1585 (O_1585,N_14191,N_14125);
and UO_1586 (O_1586,N_14891,N_14085);
or UO_1587 (O_1587,N_14521,N_14037);
nand UO_1588 (O_1588,N_14483,N_14719);
nor UO_1589 (O_1589,N_13594,N_14811);
and UO_1590 (O_1590,N_13595,N_14138);
nand UO_1591 (O_1591,N_13669,N_14272);
nor UO_1592 (O_1592,N_14549,N_13759);
nand UO_1593 (O_1593,N_14435,N_14192);
nor UO_1594 (O_1594,N_14275,N_13649);
xnor UO_1595 (O_1595,N_14671,N_14927);
or UO_1596 (O_1596,N_14408,N_13993);
and UO_1597 (O_1597,N_13621,N_14550);
or UO_1598 (O_1598,N_14152,N_14015);
or UO_1599 (O_1599,N_13694,N_14026);
and UO_1600 (O_1600,N_14212,N_13803);
xnor UO_1601 (O_1601,N_13580,N_14220);
nor UO_1602 (O_1602,N_14757,N_14211);
nand UO_1603 (O_1603,N_14301,N_14350);
nand UO_1604 (O_1604,N_14331,N_13803);
and UO_1605 (O_1605,N_13897,N_14218);
nand UO_1606 (O_1606,N_14137,N_14594);
nor UO_1607 (O_1607,N_14247,N_14731);
or UO_1608 (O_1608,N_13575,N_14211);
or UO_1609 (O_1609,N_14485,N_14397);
nand UO_1610 (O_1610,N_14764,N_14110);
or UO_1611 (O_1611,N_13892,N_14234);
or UO_1612 (O_1612,N_14437,N_14811);
nor UO_1613 (O_1613,N_13743,N_14671);
xor UO_1614 (O_1614,N_14355,N_14007);
nor UO_1615 (O_1615,N_13582,N_13777);
nor UO_1616 (O_1616,N_14140,N_14680);
and UO_1617 (O_1617,N_14633,N_13782);
xnor UO_1618 (O_1618,N_13542,N_14504);
or UO_1619 (O_1619,N_14919,N_13564);
nor UO_1620 (O_1620,N_14894,N_13568);
nor UO_1621 (O_1621,N_14949,N_13596);
or UO_1622 (O_1622,N_13783,N_13742);
or UO_1623 (O_1623,N_13707,N_14814);
xnor UO_1624 (O_1624,N_13529,N_14934);
nand UO_1625 (O_1625,N_13723,N_14593);
xor UO_1626 (O_1626,N_14587,N_13557);
and UO_1627 (O_1627,N_13581,N_13799);
xnor UO_1628 (O_1628,N_14046,N_14408);
nand UO_1629 (O_1629,N_13659,N_13948);
xnor UO_1630 (O_1630,N_13848,N_13742);
and UO_1631 (O_1631,N_14091,N_13550);
or UO_1632 (O_1632,N_13516,N_14978);
and UO_1633 (O_1633,N_14482,N_13731);
xnor UO_1634 (O_1634,N_14758,N_14543);
nor UO_1635 (O_1635,N_13540,N_14338);
or UO_1636 (O_1636,N_13584,N_14243);
or UO_1637 (O_1637,N_14233,N_14442);
nor UO_1638 (O_1638,N_14810,N_14162);
nand UO_1639 (O_1639,N_14532,N_14973);
or UO_1640 (O_1640,N_13678,N_14471);
and UO_1641 (O_1641,N_14426,N_14129);
and UO_1642 (O_1642,N_14876,N_13584);
and UO_1643 (O_1643,N_14668,N_14476);
xnor UO_1644 (O_1644,N_14810,N_13834);
and UO_1645 (O_1645,N_14651,N_14847);
and UO_1646 (O_1646,N_13955,N_13705);
nand UO_1647 (O_1647,N_13643,N_14024);
xnor UO_1648 (O_1648,N_14065,N_13670);
and UO_1649 (O_1649,N_14300,N_13870);
and UO_1650 (O_1650,N_14267,N_13574);
and UO_1651 (O_1651,N_13707,N_13877);
xor UO_1652 (O_1652,N_13759,N_14492);
nor UO_1653 (O_1653,N_14442,N_13599);
xnor UO_1654 (O_1654,N_13653,N_14833);
or UO_1655 (O_1655,N_14739,N_14357);
xnor UO_1656 (O_1656,N_13542,N_14718);
or UO_1657 (O_1657,N_14337,N_14757);
and UO_1658 (O_1658,N_14566,N_13972);
nor UO_1659 (O_1659,N_14861,N_14552);
nor UO_1660 (O_1660,N_13718,N_14480);
xor UO_1661 (O_1661,N_14249,N_13990);
and UO_1662 (O_1662,N_14105,N_14534);
and UO_1663 (O_1663,N_14644,N_14121);
nand UO_1664 (O_1664,N_14839,N_13842);
nand UO_1665 (O_1665,N_13910,N_14769);
xor UO_1666 (O_1666,N_13653,N_13769);
nand UO_1667 (O_1667,N_13716,N_13755);
nor UO_1668 (O_1668,N_13582,N_14051);
xnor UO_1669 (O_1669,N_14513,N_14466);
nand UO_1670 (O_1670,N_14889,N_13668);
xnor UO_1671 (O_1671,N_14606,N_13841);
xor UO_1672 (O_1672,N_14169,N_14316);
nand UO_1673 (O_1673,N_13726,N_14417);
nand UO_1674 (O_1674,N_14916,N_14400);
nand UO_1675 (O_1675,N_14270,N_14505);
and UO_1676 (O_1676,N_14761,N_14063);
nand UO_1677 (O_1677,N_13862,N_14168);
or UO_1678 (O_1678,N_14411,N_14052);
xnor UO_1679 (O_1679,N_14473,N_14065);
xnor UO_1680 (O_1680,N_14990,N_13550);
or UO_1681 (O_1681,N_14581,N_14906);
or UO_1682 (O_1682,N_14023,N_13847);
nand UO_1683 (O_1683,N_14301,N_14170);
or UO_1684 (O_1684,N_14742,N_13846);
nand UO_1685 (O_1685,N_13654,N_14186);
nand UO_1686 (O_1686,N_14096,N_14162);
nand UO_1687 (O_1687,N_13917,N_13720);
xor UO_1688 (O_1688,N_14486,N_14721);
or UO_1689 (O_1689,N_14814,N_14362);
nand UO_1690 (O_1690,N_14000,N_14352);
nor UO_1691 (O_1691,N_14330,N_13851);
xor UO_1692 (O_1692,N_14309,N_13723);
nand UO_1693 (O_1693,N_13917,N_13831);
nor UO_1694 (O_1694,N_14894,N_14384);
or UO_1695 (O_1695,N_13866,N_14061);
nand UO_1696 (O_1696,N_14090,N_13694);
or UO_1697 (O_1697,N_13799,N_14273);
and UO_1698 (O_1698,N_13693,N_14005);
xnor UO_1699 (O_1699,N_13732,N_14508);
nand UO_1700 (O_1700,N_14412,N_14816);
nor UO_1701 (O_1701,N_14262,N_14526);
xor UO_1702 (O_1702,N_14644,N_14616);
and UO_1703 (O_1703,N_13595,N_13644);
or UO_1704 (O_1704,N_14098,N_14937);
xnor UO_1705 (O_1705,N_14488,N_14172);
nor UO_1706 (O_1706,N_14679,N_14775);
or UO_1707 (O_1707,N_14375,N_14522);
or UO_1708 (O_1708,N_13750,N_13572);
or UO_1709 (O_1709,N_14278,N_14807);
and UO_1710 (O_1710,N_14798,N_13652);
xnor UO_1711 (O_1711,N_14500,N_13646);
xor UO_1712 (O_1712,N_13592,N_14624);
nand UO_1713 (O_1713,N_14083,N_13643);
and UO_1714 (O_1714,N_13939,N_14098);
nand UO_1715 (O_1715,N_14974,N_14224);
and UO_1716 (O_1716,N_13887,N_14589);
xnor UO_1717 (O_1717,N_14970,N_14127);
and UO_1718 (O_1718,N_13653,N_13538);
nor UO_1719 (O_1719,N_14710,N_14364);
or UO_1720 (O_1720,N_14165,N_14299);
or UO_1721 (O_1721,N_14379,N_14686);
nand UO_1722 (O_1722,N_14378,N_13661);
or UO_1723 (O_1723,N_14233,N_14303);
xor UO_1724 (O_1724,N_13606,N_14188);
nor UO_1725 (O_1725,N_14438,N_14450);
and UO_1726 (O_1726,N_14046,N_14023);
xnor UO_1727 (O_1727,N_14970,N_14683);
or UO_1728 (O_1728,N_14447,N_14984);
and UO_1729 (O_1729,N_13904,N_14756);
nor UO_1730 (O_1730,N_14438,N_13575);
nor UO_1731 (O_1731,N_13801,N_14560);
and UO_1732 (O_1732,N_14780,N_13702);
nor UO_1733 (O_1733,N_13561,N_13545);
or UO_1734 (O_1734,N_13753,N_14010);
xor UO_1735 (O_1735,N_14561,N_13745);
xor UO_1736 (O_1736,N_14365,N_14014);
or UO_1737 (O_1737,N_14721,N_13985);
nor UO_1738 (O_1738,N_13688,N_14439);
nand UO_1739 (O_1739,N_14998,N_13898);
or UO_1740 (O_1740,N_13553,N_14220);
nor UO_1741 (O_1741,N_13859,N_14831);
and UO_1742 (O_1742,N_14789,N_13552);
nor UO_1743 (O_1743,N_14752,N_13555);
xor UO_1744 (O_1744,N_14265,N_14018);
or UO_1745 (O_1745,N_14549,N_14249);
or UO_1746 (O_1746,N_14295,N_13666);
and UO_1747 (O_1747,N_13730,N_13747);
xnor UO_1748 (O_1748,N_14364,N_13769);
nand UO_1749 (O_1749,N_13758,N_14459);
or UO_1750 (O_1750,N_13609,N_13770);
and UO_1751 (O_1751,N_14462,N_14564);
and UO_1752 (O_1752,N_14525,N_14140);
nand UO_1753 (O_1753,N_14157,N_14729);
nand UO_1754 (O_1754,N_14681,N_13535);
nor UO_1755 (O_1755,N_13681,N_14906);
or UO_1756 (O_1756,N_14327,N_14167);
xnor UO_1757 (O_1757,N_14012,N_14512);
xnor UO_1758 (O_1758,N_14088,N_14917);
nor UO_1759 (O_1759,N_13909,N_14496);
or UO_1760 (O_1760,N_14448,N_14221);
and UO_1761 (O_1761,N_14508,N_14209);
xnor UO_1762 (O_1762,N_14106,N_14932);
xor UO_1763 (O_1763,N_13794,N_13636);
nor UO_1764 (O_1764,N_13682,N_14403);
or UO_1765 (O_1765,N_14950,N_14195);
and UO_1766 (O_1766,N_14203,N_14193);
and UO_1767 (O_1767,N_13828,N_14758);
xnor UO_1768 (O_1768,N_14415,N_14595);
or UO_1769 (O_1769,N_14702,N_14482);
and UO_1770 (O_1770,N_13559,N_14625);
nand UO_1771 (O_1771,N_14618,N_14522);
or UO_1772 (O_1772,N_14453,N_14882);
xnor UO_1773 (O_1773,N_14292,N_14882);
xor UO_1774 (O_1774,N_13841,N_14920);
nor UO_1775 (O_1775,N_13517,N_14978);
nor UO_1776 (O_1776,N_13730,N_13592);
nor UO_1777 (O_1777,N_14781,N_14586);
and UO_1778 (O_1778,N_14565,N_14668);
nand UO_1779 (O_1779,N_14130,N_14986);
nand UO_1780 (O_1780,N_14549,N_14052);
xor UO_1781 (O_1781,N_14348,N_13587);
nand UO_1782 (O_1782,N_13573,N_14237);
nor UO_1783 (O_1783,N_13574,N_14328);
nand UO_1784 (O_1784,N_14930,N_13585);
nand UO_1785 (O_1785,N_14819,N_14579);
nor UO_1786 (O_1786,N_14139,N_14690);
xor UO_1787 (O_1787,N_13508,N_14242);
and UO_1788 (O_1788,N_14501,N_14042);
or UO_1789 (O_1789,N_13733,N_14658);
and UO_1790 (O_1790,N_13982,N_14052);
nand UO_1791 (O_1791,N_13789,N_13704);
or UO_1792 (O_1792,N_13819,N_14263);
nand UO_1793 (O_1793,N_14207,N_14506);
nor UO_1794 (O_1794,N_13753,N_14060);
and UO_1795 (O_1795,N_14716,N_13948);
nor UO_1796 (O_1796,N_14563,N_14396);
and UO_1797 (O_1797,N_13873,N_14604);
and UO_1798 (O_1798,N_14700,N_13784);
or UO_1799 (O_1799,N_14196,N_14286);
or UO_1800 (O_1800,N_13706,N_14402);
and UO_1801 (O_1801,N_14221,N_14976);
and UO_1802 (O_1802,N_14374,N_14101);
or UO_1803 (O_1803,N_14150,N_14419);
and UO_1804 (O_1804,N_13963,N_14131);
or UO_1805 (O_1805,N_14262,N_14920);
nand UO_1806 (O_1806,N_14130,N_14301);
nand UO_1807 (O_1807,N_13757,N_13857);
nor UO_1808 (O_1808,N_14731,N_13595);
nand UO_1809 (O_1809,N_14520,N_14866);
nand UO_1810 (O_1810,N_13532,N_14837);
xnor UO_1811 (O_1811,N_14631,N_14690);
xnor UO_1812 (O_1812,N_14847,N_13523);
or UO_1813 (O_1813,N_13996,N_14015);
or UO_1814 (O_1814,N_13526,N_14249);
or UO_1815 (O_1815,N_14565,N_14468);
nand UO_1816 (O_1816,N_14173,N_13635);
xor UO_1817 (O_1817,N_13633,N_14028);
nand UO_1818 (O_1818,N_14540,N_14131);
xor UO_1819 (O_1819,N_14824,N_14548);
nand UO_1820 (O_1820,N_14272,N_13994);
or UO_1821 (O_1821,N_14231,N_14320);
or UO_1822 (O_1822,N_14829,N_14030);
nor UO_1823 (O_1823,N_14974,N_14707);
nor UO_1824 (O_1824,N_14864,N_14453);
nand UO_1825 (O_1825,N_14964,N_14704);
and UO_1826 (O_1826,N_14254,N_13726);
xor UO_1827 (O_1827,N_14698,N_14773);
and UO_1828 (O_1828,N_14598,N_14974);
and UO_1829 (O_1829,N_14646,N_14816);
xor UO_1830 (O_1830,N_13524,N_14957);
and UO_1831 (O_1831,N_14030,N_13972);
xnor UO_1832 (O_1832,N_14710,N_14333);
nor UO_1833 (O_1833,N_13510,N_14796);
and UO_1834 (O_1834,N_14413,N_14533);
nand UO_1835 (O_1835,N_14197,N_14418);
nor UO_1836 (O_1836,N_14157,N_13585);
xnor UO_1837 (O_1837,N_14247,N_14102);
xor UO_1838 (O_1838,N_14906,N_14058);
and UO_1839 (O_1839,N_14750,N_14039);
nand UO_1840 (O_1840,N_13910,N_13775);
xnor UO_1841 (O_1841,N_13764,N_14901);
nor UO_1842 (O_1842,N_14883,N_14304);
nor UO_1843 (O_1843,N_13558,N_14551);
xnor UO_1844 (O_1844,N_14502,N_13663);
nor UO_1845 (O_1845,N_13662,N_13740);
xor UO_1846 (O_1846,N_13716,N_14649);
and UO_1847 (O_1847,N_13901,N_14574);
or UO_1848 (O_1848,N_14682,N_14543);
nand UO_1849 (O_1849,N_14307,N_14356);
xnor UO_1850 (O_1850,N_14745,N_13848);
and UO_1851 (O_1851,N_14137,N_14019);
or UO_1852 (O_1852,N_13869,N_13585);
nor UO_1853 (O_1853,N_13559,N_14101);
xnor UO_1854 (O_1854,N_13807,N_13595);
nor UO_1855 (O_1855,N_14369,N_13591);
xnor UO_1856 (O_1856,N_14762,N_14907);
or UO_1857 (O_1857,N_14116,N_13510);
nand UO_1858 (O_1858,N_14809,N_13559);
or UO_1859 (O_1859,N_14458,N_14465);
nor UO_1860 (O_1860,N_13569,N_14095);
xor UO_1861 (O_1861,N_13966,N_13673);
xor UO_1862 (O_1862,N_14820,N_14445);
and UO_1863 (O_1863,N_13668,N_14331);
nor UO_1864 (O_1864,N_13584,N_14772);
or UO_1865 (O_1865,N_14115,N_14296);
nand UO_1866 (O_1866,N_14777,N_14767);
or UO_1867 (O_1867,N_14938,N_14088);
or UO_1868 (O_1868,N_14782,N_14218);
nand UO_1869 (O_1869,N_13777,N_13537);
or UO_1870 (O_1870,N_14092,N_14428);
or UO_1871 (O_1871,N_14618,N_13907);
xor UO_1872 (O_1872,N_14276,N_14489);
nor UO_1873 (O_1873,N_14280,N_14658);
and UO_1874 (O_1874,N_14118,N_14361);
or UO_1875 (O_1875,N_14831,N_14009);
nand UO_1876 (O_1876,N_13747,N_14804);
xnor UO_1877 (O_1877,N_13547,N_14436);
xor UO_1878 (O_1878,N_14936,N_14787);
and UO_1879 (O_1879,N_14133,N_14595);
nor UO_1880 (O_1880,N_14761,N_14335);
nor UO_1881 (O_1881,N_13775,N_14026);
and UO_1882 (O_1882,N_13551,N_14539);
nand UO_1883 (O_1883,N_14818,N_14971);
nor UO_1884 (O_1884,N_13679,N_14244);
xor UO_1885 (O_1885,N_14913,N_13965);
and UO_1886 (O_1886,N_13802,N_14608);
and UO_1887 (O_1887,N_13712,N_14162);
nand UO_1888 (O_1888,N_14573,N_13901);
or UO_1889 (O_1889,N_14672,N_14275);
nand UO_1890 (O_1890,N_14669,N_13559);
or UO_1891 (O_1891,N_14433,N_14988);
nor UO_1892 (O_1892,N_13834,N_14483);
and UO_1893 (O_1893,N_14150,N_14602);
or UO_1894 (O_1894,N_14761,N_13602);
and UO_1895 (O_1895,N_13619,N_14636);
xor UO_1896 (O_1896,N_14266,N_14170);
nor UO_1897 (O_1897,N_14740,N_13698);
nor UO_1898 (O_1898,N_13793,N_13532);
nand UO_1899 (O_1899,N_14663,N_13626);
nor UO_1900 (O_1900,N_14878,N_14395);
xor UO_1901 (O_1901,N_14281,N_14956);
nor UO_1902 (O_1902,N_14954,N_14544);
xnor UO_1903 (O_1903,N_14314,N_14985);
and UO_1904 (O_1904,N_13735,N_14452);
nor UO_1905 (O_1905,N_13533,N_14451);
xnor UO_1906 (O_1906,N_14202,N_13731);
xnor UO_1907 (O_1907,N_14721,N_14258);
and UO_1908 (O_1908,N_13899,N_13796);
nor UO_1909 (O_1909,N_13575,N_14838);
and UO_1910 (O_1910,N_13702,N_14889);
nand UO_1911 (O_1911,N_14685,N_14498);
xor UO_1912 (O_1912,N_13806,N_14150);
and UO_1913 (O_1913,N_14203,N_14669);
nor UO_1914 (O_1914,N_14736,N_14332);
and UO_1915 (O_1915,N_14496,N_14819);
or UO_1916 (O_1916,N_13626,N_14967);
or UO_1917 (O_1917,N_14676,N_14393);
nor UO_1918 (O_1918,N_13540,N_14274);
and UO_1919 (O_1919,N_14856,N_14131);
nor UO_1920 (O_1920,N_14997,N_14028);
and UO_1921 (O_1921,N_14488,N_14124);
xnor UO_1922 (O_1922,N_14406,N_14565);
or UO_1923 (O_1923,N_14210,N_14326);
nand UO_1924 (O_1924,N_14425,N_14078);
nand UO_1925 (O_1925,N_14650,N_13960);
nand UO_1926 (O_1926,N_14664,N_14035);
xnor UO_1927 (O_1927,N_14905,N_13563);
or UO_1928 (O_1928,N_14725,N_14380);
and UO_1929 (O_1929,N_13804,N_14554);
nand UO_1930 (O_1930,N_13906,N_13599);
nand UO_1931 (O_1931,N_14182,N_14082);
or UO_1932 (O_1932,N_14898,N_14298);
xor UO_1933 (O_1933,N_14646,N_14064);
nand UO_1934 (O_1934,N_14035,N_13758);
and UO_1935 (O_1935,N_14576,N_14088);
or UO_1936 (O_1936,N_14154,N_13989);
and UO_1937 (O_1937,N_14482,N_14806);
or UO_1938 (O_1938,N_14390,N_14146);
xnor UO_1939 (O_1939,N_14667,N_13654);
and UO_1940 (O_1940,N_14456,N_14244);
and UO_1941 (O_1941,N_14193,N_13832);
nand UO_1942 (O_1942,N_14986,N_14738);
or UO_1943 (O_1943,N_13843,N_13682);
xnor UO_1944 (O_1944,N_14612,N_14270);
xnor UO_1945 (O_1945,N_14082,N_14757);
xnor UO_1946 (O_1946,N_14473,N_13770);
or UO_1947 (O_1947,N_13746,N_13876);
and UO_1948 (O_1948,N_13890,N_14466);
or UO_1949 (O_1949,N_14810,N_13687);
xor UO_1950 (O_1950,N_14419,N_14757);
nor UO_1951 (O_1951,N_13572,N_13997);
and UO_1952 (O_1952,N_14809,N_13916);
nor UO_1953 (O_1953,N_14706,N_14225);
or UO_1954 (O_1954,N_14032,N_14195);
xnor UO_1955 (O_1955,N_14876,N_14418);
nand UO_1956 (O_1956,N_14404,N_14017);
nand UO_1957 (O_1957,N_13773,N_14253);
and UO_1958 (O_1958,N_14938,N_13614);
xnor UO_1959 (O_1959,N_14507,N_14424);
and UO_1960 (O_1960,N_13813,N_14772);
nor UO_1961 (O_1961,N_13940,N_14033);
nand UO_1962 (O_1962,N_13868,N_14073);
nor UO_1963 (O_1963,N_14434,N_14229);
and UO_1964 (O_1964,N_13594,N_14990);
nand UO_1965 (O_1965,N_14789,N_13573);
nand UO_1966 (O_1966,N_14951,N_13683);
nor UO_1967 (O_1967,N_14785,N_13843);
xor UO_1968 (O_1968,N_14579,N_13833);
nor UO_1969 (O_1969,N_14263,N_14065);
and UO_1970 (O_1970,N_14028,N_13705);
and UO_1971 (O_1971,N_14461,N_14522);
and UO_1972 (O_1972,N_14539,N_14220);
and UO_1973 (O_1973,N_13853,N_14240);
nand UO_1974 (O_1974,N_14639,N_14156);
nor UO_1975 (O_1975,N_14079,N_14015);
and UO_1976 (O_1976,N_14228,N_14140);
or UO_1977 (O_1977,N_14532,N_13567);
nand UO_1978 (O_1978,N_14976,N_14102);
and UO_1979 (O_1979,N_14126,N_14037);
xnor UO_1980 (O_1980,N_13869,N_13702);
nor UO_1981 (O_1981,N_14618,N_14591);
and UO_1982 (O_1982,N_13632,N_13928);
nor UO_1983 (O_1983,N_14905,N_14129);
and UO_1984 (O_1984,N_13667,N_14097);
nor UO_1985 (O_1985,N_13895,N_14893);
and UO_1986 (O_1986,N_14593,N_14072);
and UO_1987 (O_1987,N_14698,N_14753);
nand UO_1988 (O_1988,N_13856,N_14662);
or UO_1989 (O_1989,N_13971,N_14557);
xnor UO_1990 (O_1990,N_14292,N_14922);
and UO_1991 (O_1991,N_13525,N_13621);
nand UO_1992 (O_1992,N_14499,N_13907);
nand UO_1993 (O_1993,N_14656,N_13885);
xnor UO_1994 (O_1994,N_14465,N_14961);
nand UO_1995 (O_1995,N_13624,N_13749);
nor UO_1996 (O_1996,N_13681,N_13656);
nand UO_1997 (O_1997,N_13806,N_13853);
and UO_1998 (O_1998,N_13694,N_14326);
nand UO_1999 (O_1999,N_14847,N_14742);
endmodule