module basic_500_3000_500_50_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_333,In_458);
nor U1 (N_1,In_268,In_129);
or U2 (N_2,In_19,In_317);
or U3 (N_3,In_322,In_81);
nand U4 (N_4,In_424,In_140);
nand U5 (N_5,In_489,In_3);
or U6 (N_6,In_395,In_242);
or U7 (N_7,In_83,In_113);
xor U8 (N_8,In_102,In_125);
and U9 (N_9,In_288,In_35);
or U10 (N_10,In_319,In_362);
or U11 (N_11,In_97,In_176);
or U12 (N_12,In_192,In_130);
nand U13 (N_13,In_169,In_407);
and U14 (N_14,In_492,In_289);
nor U15 (N_15,In_269,In_165);
or U16 (N_16,In_20,In_281);
or U17 (N_17,In_300,In_25);
and U18 (N_18,In_157,In_109);
nand U19 (N_19,In_227,In_496);
nor U20 (N_20,In_141,In_441);
nand U21 (N_21,In_89,In_405);
and U22 (N_22,In_431,In_161);
xor U23 (N_23,In_43,In_200);
or U24 (N_24,In_133,In_206);
or U25 (N_25,In_122,In_173);
nor U26 (N_26,In_400,In_79);
nand U27 (N_27,In_7,In_360);
nor U28 (N_28,In_344,In_142);
nand U29 (N_29,In_33,In_264);
or U30 (N_30,In_175,In_308);
nor U31 (N_31,In_382,In_37);
and U32 (N_32,In_296,In_427);
nor U33 (N_33,In_0,In_442);
nor U34 (N_34,In_450,In_364);
and U35 (N_35,In_486,In_294);
and U36 (N_36,In_180,In_104);
nor U37 (N_37,In_318,In_485);
and U38 (N_38,In_218,In_316);
nor U39 (N_39,In_376,In_454);
and U40 (N_40,In_430,In_291);
or U41 (N_41,In_466,In_249);
and U42 (N_42,In_85,In_399);
and U43 (N_43,In_61,In_283);
nor U44 (N_44,In_66,In_132);
nand U45 (N_45,In_178,In_325);
nand U46 (N_46,In_114,In_260);
or U47 (N_47,In_383,In_44);
or U48 (N_48,In_42,In_480);
and U49 (N_49,In_315,In_267);
or U50 (N_50,In_82,In_396);
or U51 (N_51,In_185,In_251);
nand U52 (N_52,In_208,In_380);
or U53 (N_53,In_62,In_198);
and U54 (N_54,In_57,In_397);
or U55 (N_55,In_354,In_16);
nor U56 (N_56,In_170,In_247);
and U57 (N_57,In_95,In_499);
nand U58 (N_58,In_334,In_80);
and U59 (N_59,In_272,In_168);
nor U60 (N_60,In_301,In_93);
and U61 (N_61,In_307,In_409);
and U62 (N_62,In_460,In_342);
and U63 (N_63,In_92,In_416);
and U64 (N_64,In_10,In_50);
nand U65 (N_65,In_337,In_154);
nor U66 (N_66,In_422,N_38);
or U67 (N_67,In_320,In_94);
nand U68 (N_68,N_19,In_369);
nor U69 (N_69,In_265,In_151);
or U70 (N_70,In_49,In_131);
nand U71 (N_71,In_63,In_284);
and U72 (N_72,In_26,In_209);
or U73 (N_73,In_412,In_327);
nor U74 (N_74,In_236,N_4);
nand U75 (N_75,In_225,In_38);
nor U76 (N_76,In_363,In_415);
nand U77 (N_77,In_230,In_116);
nor U78 (N_78,In_343,In_495);
nor U79 (N_79,In_40,N_20);
or U80 (N_80,In_324,In_401);
and U81 (N_81,In_56,In_494);
or U82 (N_82,In_100,In_429);
or U83 (N_83,In_439,In_410);
nor U84 (N_84,N_40,In_403);
and U85 (N_85,In_381,In_243);
nor U86 (N_86,In_463,In_217);
or U87 (N_87,In_336,In_41);
or U88 (N_88,N_5,In_445);
nand U89 (N_89,N_33,In_457);
and U90 (N_90,In_271,In_348);
nor U91 (N_91,In_45,In_426);
and U92 (N_92,In_418,In_254);
nor U93 (N_93,In_475,In_367);
and U94 (N_94,In_34,In_448);
or U95 (N_95,In_196,In_358);
nand U96 (N_96,In_223,In_136);
nor U97 (N_97,In_446,In_275);
or U98 (N_98,In_118,In_237);
nand U99 (N_99,In_58,In_203);
or U100 (N_100,N_49,N_27);
or U101 (N_101,In_245,In_123);
nand U102 (N_102,In_436,In_77);
nor U103 (N_103,In_323,In_329);
and U104 (N_104,In_330,In_425);
nand U105 (N_105,In_166,In_210);
nand U106 (N_106,In_326,In_195);
nor U107 (N_107,In_224,In_359);
and U108 (N_108,In_191,In_314);
or U109 (N_109,In_404,In_179);
and U110 (N_110,In_366,In_444);
and U111 (N_111,In_304,N_44);
nand U112 (N_112,In_103,In_357);
nand U113 (N_113,In_467,In_321);
or U114 (N_114,In_378,In_392);
nor U115 (N_115,In_212,In_65);
nor U116 (N_116,N_23,In_69);
nor U117 (N_117,In_164,In_88);
or U118 (N_118,In_120,In_146);
nand U119 (N_119,In_101,In_110);
nor U120 (N_120,In_371,In_328);
nor U121 (N_121,In_465,N_59);
nand U122 (N_122,In_302,N_2);
and U123 (N_123,In_338,In_263);
and U124 (N_124,N_9,N_68);
or U125 (N_125,In_470,N_14);
nand U126 (N_126,In_350,In_440);
or U127 (N_127,In_473,In_258);
and U128 (N_128,In_469,In_32);
nand U129 (N_129,N_58,N_42);
nand U130 (N_130,In_280,In_287);
and U131 (N_131,N_88,In_174);
or U132 (N_132,N_78,N_6);
or U133 (N_133,N_26,In_127);
and U134 (N_134,In_435,N_30);
or U135 (N_135,In_64,In_353);
nand U136 (N_136,In_197,In_117);
nor U137 (N_137,In_148,N_45);
nand U138 (N_138,In_193,In_384);
and U139 (N_139,In_5,N_66);
or U140 (N_140,In_331,In_310);
nand U141 (N_141,In_414,In_278);
and U142 (N_142,In_163,In_241);
nor U143 (N_143,In_68,N_73);
nand U144 (N_144,In_262,In_75);
nand U145 (N_145,In_239,In_377);
nand U146 (N_146,N_35,In_172);
nor U147 (N_147,In_107,N_39);
and U148 (N_148,In_214,In_1);
nor U149 (N_149,In_55,In_472);
or U150 (N_150,N_119,In_213);
or U151 (N_151,In_189,N_62);
or U152 (N_152,N_117,In_452);
nand U153 (N_153,N_53,In_411);
nand U154 (N_154,In_459,In_462);
nand U155 (N_155,In_413,N_97);
and U156 (N_156,In_13,In_15);
nor U157 (N_157,In_158,N_65);
and U158 (N_158,N_93,In_71);
nor U159 (N_159,N_28,N_101);
nor U160 (N_160,N_43,N_87);
nand U161 (N_161,In_194,In_273);
xor U162 (N_162,In_87,N_3);
nand U163 (N_163,In_156,N_115);
and U164 (N_164,N_22,In_27);
or U165 (N_165,In_149,In_277);
or U166 (N_166,In_78,In_167);
nor U167 (N_167,In_276,In_250);
nand U168 (N_168,In_211,In_60);
nor U169 (N_169,In_143,In_220);
or U170 (N_170,N_71,N_75);
nand U171 (N_171,In_286,In_39);
nand U172 (N_172,In_370,N_111);
nor U173 (N_173,N_79,In_352);
and U174 (N_174,In_23,In_229);
nor U175 (N_175,N_8,In_244);
nor U176 (N_176,In_488,In_346);
nand U177 (N_177,In_135,N_96);
or U178 (N_178,In_390,N_34);
nand U179 (N_179,In_379,In_128);
or U180 (N_180,In_86,N_0);
or U181 (N_181,In_4,In_238);
or U182 (N_182,N_170,In_76);
nor U183 (N_183,N_64,In_279);
and U184 (N_184,In_160,N_146);
nor U185 (N_185,In_138,In_438);
nor U186 (N_186,In_368,N_54);
nor U187 (N_187,In_248,In_144);
and U188 (N_188,In_234,In_150);
xor U189 (N_189,In_171,In_456);
nor U190 (N_190,N_150,N_105);
nor U191 (N_191,N_140,N_152);
nand U192 (N_192,In_115,N_107);
nor U193 (N_193,In_256,In_186);
nand U194 (N_194,N_84,N_98);
or U195 (N_195,N_143,In_14);
or U196 (N_196,In_391,In_385);
nor U197 (N_197,In_52,In_389);
nor U198 (N_198,N_46,In_290);
and U199 (N_199,In_36,In_482);
xnor U200 (N_200,N_112,In_204);
or U201 (N_201,In_187,In_491);
nand U202 (N_202,N_144,In_6);
nor U203 (N_203,In_240,In_222);
or U204 (N_204,In_365,In_309);
nand U205 (N_205,In_282,In_285);
or U206 (N_206,In_434,N_156);
and U207 (N_207,In_408,N_167);
nor U208 (N_208,In_199,N_165);
nand U209 (N_209,In_112,In_487);
nor U210 (N_210,N_48,N_116);
nor U211 (N_211,In_266,N_128);
and U212 (N_212,In_339,N_157);
and U213 (N_213,N_109,N_120);
and U214 (N_214,N_164,N_174);
and U215 (N_215,In_183,N_7);
nand U216 (N_216,In_29,In_388);
nand U217 (N_217,In_124,In_184);
or U218 (N_218,In_443,In_257);
or U219 (N_219,In_349,In_181);
and U220 (N_220,N_85,N_83);
and U221 (N_221,N_137,N_100);
nand U222 (N_222,In_299,In_216);
or U223 (N_223,In_474,In_84);
and U224 (N_224,In_471,In_98);
nor U225 (N_225,In_493,In_259);
nor U226 (N_226,In_54,In_202);
nand U227 (N_227,N_57,In_31);
and U228 (N_228,N_21,In_46);
nor U229 (N_229,In_453,In_498);
and U230 (N_230,In_159,In_48);
or U231 (N_231,In_219,In_11);
and U232 (N_232,In_455,In_226);
and U233 (N_233,In_406,N_41);
or U234 (N_234,N_132,N_108);
nor U235 (N_235,N_148,In_67);
nand U236 (N_236,In_417,N_166);
or U237 (N_237,In_478,In_312);
and U238 (N_238,N_24,N_70);
or U239 (N_239,N_163,N_36);
nand U240 (N_240,In_228,In_137);
nor U241 (N_241,N_131,In_235);
and U242 (N_242,In_215,In_394);
nand U243 (N_243,In_207,In_232);
nand U244 (N_244,N_90,N_236);
or U245 (N_245,N_77,N_199);
nand U246 (N_246,In_437,N_212);
nand U247 (N_247,In_106,N_127);
or U248 (N_248,In_479,In_372);
or U249 (N_249,In_47,N_202);
nor U250 (N_250,In_205,N_63);
nand U251 (N_251,N_125,In_461);
nor U252 (N_252,In_332,N_192);
nand U253 (N_253,N_215,N_113);
nand U254 (N_254,N_145,In_91);
and U255 (N_255,In_177,In_433);
and U256 (N_256,N_16,In_423);
or U257 (N_257,In_451,In_2);
nor U258 (N_258,In_447,N_190);
and U259 (N_259,N_197,N_168);
nand U260 (N_260,In_96,N_13);
and U261 (N_261,N_110,N_179);
and U262 (N_262,N_89,N_126);
and U263 (N_263,N_86,In_155);
nand U264 (N_264,N_95,N_217);
nand U265 (N_265,N_92,In_72);
nand U266 (N_266,In_12,In_421);
and U267 (N_267,In_24,N_158);
or U268 (N_268,N_103,N_134);
and U269 (N_269,In_99,N_175);
or U270 (N_270,N_169,In_311);
or U271 (N_271,N_177,In_476);
or U272 (N_272,In_297,In_53);
nand U273 (N_273,N_61,In_373);
or U274 (N_274,N_106,N_12);
xor U275 (N_275,N_102,N_180);
or U276 (N_276,N_55,In_119);
nor U277 (N_277,N_204,In_108);
and U278 (N_278,N_29,N_155);
nand U279 (N_279,N_198,N_122);
nand U280 (N_280,In_419,In_387);
and U281 (N_281,In_246,N_124);
nor U282 (N_282,N_31,N_221);
or U283 (N_283,N_67,N_216);
or U284 (N_284,In_261,N_219);
and U285 (N_285,In_70,N_32);
or U286 (N_286,N_208,N_209);
nand U287 (N_287,N_205,N_191);
and U288 (N_288,N_118,N_193);
nor U289 (N_289,N_226,In_22);
nand U290 (N_290,In_361,In_111);
nor U291 (N_291,N_206,N_210);
and U292 (N_292,In_484,In_306);
and U293 (N_293,N_182,In_298);
and U294 (N_294,N_238,N_25);
or U295 (N_295,In_90,In_18);
nor U296 (N_296,N_227,N_232);
or U297 (N_297,N_229,N_173);
nand U298 (N_298,In_340,N_200);
or U299 (N_299,N_136,N_186);
nor U300 (N_300,N_207,N_283);
nor U301 (N_301,N_296,In_468);
nand U302 (N_302,In_59,In_375);
nor U303 (N_303,In_231,N_56);
nand U304 (N_304,N_214,N_181);
and U305 (N_305,N_82,N_187);
nand U306 (N_306,N_278,N_289);
nor U307 (N_307,N_203,N_268);
nand U308 (N_308,N_272,N_185);
and U309 (N_309,In_356,In_190);
or U310 (N_310,In_303,In_145);
nand U311 (N_311,N_255,N_287);
nor U312 (N_312,N_142,In_386);
and U313 (N_313,N_183,In_8);
nand U314 (N_314,N_243,N_270);
nand U315 (N_315,In_30,In_17);
or U316 (N_316,N_244,N_51);
nand U317 (N_317,N_263,N_121);
nand U318 (N_318,N_298,N_141);
nand U319 (N_319,N_247,N_235);
nor U320 (N_320,N_242,N_104);
and U321 (N_321,In_121,N_250);
nand U322 (N_322,In_420,N_276);
or U323 (N_323,N_114,N_50);
nand U324 (N_324,N_290,N_159);
nand U325 (N_325,N_195,In_73);
nand U326 (N_326,N_37,N_251);
and U327 (N_327,N_264,N_291);
nand U328 (N_328,In_252,N_176);
nand U329 (N_329,N_297,In_341);
nand U330 (N_330,N_249,In_295);
nand U331 (N_331,N_246,N_241);
or U332 (N_332,N_288,N_123);
or U333 (N_333,N_138,N_162);
and U334 (N_334,N_282,In_490);
or U335 (N_335,N_147,In_126);
and U336 (N_336,N_196,N_201);
nor U337 (N_337,N_60,N_171);
nand U338 (N_338,N_189,In_105);
nor U339 (N_339,N_153,N_252);
or U340 (N_340,N_80,N_172);
and U341 (N_341,In_428,N_224);
nor U342 (N_342,N_91,In_274);
or U343 (N_343,In_147,In_182);
or U344 (N_344,N_18,N_271);
or U345 (N_345,N_230,N_262);
nor U346 (N_346,N_253,In_233);
nand U347 (N_347,In_393,N_293);
nand U348 (N_348,N_260,N_257);
nor U349 (N_349,In_355,N_258);
and U350 (N_350,In_152,In_313);
and U351 (N_351,N_286,In_293);
and U352 (N_352,N_178,N_213);
or U353 (N_353,In_270,In_139);
nor U354 (N_354,In_402,N_237);
or U355 (N_355,N_130,In_292);
nand U356 (N_356,N_139,N_292);
nor U357 (N_357,N_256,In_477);
nand U358 (N_358,N_299,In_201);
and U359 (N_359,In_497,N_99);
or U360 (N_360,N_135,N_277);
nor U361 (N_361,N_331,In_335);
nor U362 (N_362,N_314,N_218);
or U363 (N_363,N_326,N_359);
nor U364 (N_364,N_302,N_325);
nor U365 (N_365,N_154,N_348);
or U366 (N_366,N_259,N_339);
and U367 (N_367,N_344,N_346);
and U368 (N_368,N_318,N_349);
and U369 (N_369,N_308,N_343);
nor U370 (N_370,N_341,N_222);
or U371 (N_371,N_231,N_347);
or U372 (N_372,N_307,N_194);
and U373 (N_373,In_253,In_483);
or U374 (N_374,In_464,In_153);
or U375 (N_375,N_254,N_327);
nand U376 (N_376,N_322,N_69);
nand U377 (N_377,N_300,In_221);
or U378 (N_378,N_315,N_338);
and U379 (N_379,N_358,In_398);
and U380 (N_380,N_225,N_320);
or U381 (N_381,N_310,N_1);
or U382 (N_382,In_51,N_311);
nor U383 (N_383,N_316,N_15);
or U384 (N_384,N_305,N_306);
nand U385 (N_385,N_345,In_374);
nor U386 (N_386,N_335,N_281);
nand U387 (N_387,N_319,In_449);
and U388 (N_388,N_261,N_266);
nand U389 (N_389,N_324,N_355);
nand U390 (N_390,N_357,In_351);
or U391 (N_391,In_162,In_9);
nor U392 (N_392,N_211,N_352);
or U393 (N_393,N_267,N_220);
nor U394 (N_394,N_285,N_265);
nor U395 (N_395,N_11,N_228);
nand U396 (N_396,N_340,N_334);
nor U397 (N_397,N_350,In_74);
and U398 (N_398,In_255,N_223);
and U399 (N_399,N_184,In_481);
nor U400 (N_400,N_337,N_94);
nand U401 (N_401,In_188,N_81);
or U402 (N_402,N_313,N_269);
nor U403 (N_403,N_356,N_149);
or U404 (N_404,N_336,In_28);
and U405 (N_405,N_151,N_74);
nor U406 (N_406,N_295,N_329);
and U407 (N_407,N_240,N_328);
nand U408 (N_408,In_21,N_351);
nor U409 (N_409,N_10,N_273);
nor U410 (N_410,In_305,N_160);
and U411 (N_411,In_345,N_323);
or U412 (N_412,N_188,N_301);
nand U413 (N_413,N_303,In_432);
or U414 (N_414,N_280,N_342);
and U415 (N_415,N_304,N_76);
nor U416 (N_416,N_279,N_72);
nor U417 (N_417,N_354,In_134);
nand U418 (N_418,N_233,N_248);
nand U419 (N_419,N_321,N_133);
xor U420 (N_420,N_401,N_384);
and U421 (N_421,N_17,N_129);
and U422 (N_422,N_369,N_383);
nor U423 (N_423,N_398,N_407);
nor U424 (N_424,N_368,N_378);
or U425 (N_425,N_396,N_239);
nand U426 (N_426,N_415,N_413);
nor U427 (N_427,N_400,N_385);
nor U428 (N_428,N_361,N_284);
nor U429 (N_429,N_394,N_379);
nand U430 (N_430,N_382,N_234);
nand U431 (N_431,In_347,N_363);
and U432 (N_432,N_371,N_402);
and U433 (N_433,N_412,N_416);
and U434 (N_434,N_408,N_370);
or U435 (N_435,N_387,N_409);
or U436 (N_436,N_245,N_373);
nor U437 (N_437,N_294,N_406);
nand U438 (N_438,N_390,N_380);
nor U439 (N_439,N_410,N_391);
nor U440 (N_440,N_386,N_161);
nor U441 (N_441,N_397,N_405);
nor U442 (N_442,N_417,N_333);
nor U443 (N_443,N_366,N_372);
or U444 (N_444,N_364,N_317);
nor U445 (N_445,N_52,N_388);
or U446 (N_446,N_389,N_403);
or U447 (N_447,N_404,N_360);
nor U448 (N_448,N_274,N_365);
or U449 (N_449,N_419,N_374);
nand U450 (N_450,N_399,N_381);
nand U451 (N_451,N_47,N_330);
or U452 (N_452,N_275,N_395);
nand U453 (N_453,N_414,N_411);
and U454 (N_454,N_376,N_393);
or U455 (N_455,N_362,N_418);
nand U456 (N_456,N_309,N_332);
and U457 (N_457,N_353,N_375);
and U458 (N_458,N_377,N_367);
or U459 (N_459,N_312,N_392);
and U460 (N_460,N_367,N_387);
nand U461 (N_461,N_17,N_365);
and U462 (N_462,N_416,N_391);
or U463 (N_463,N_370,N_409);
or U464 (N_464,N_366,N_360);
and U465 (N_465,N_394,N_386);
or U466 (N_466,N_364,N_373);
or U467 (N_467,N_52,N_413);
nand U468 (N_468,N_401,N_380);
nand U469 (N_469,N_367,N_412);
nand U470 (N_470,N_384,N_364);
and U471 (N_471,N_371,N_406);
and U472 (N_472,N_365,N_410);
and U473 (N_473,N_47,N_385);
nor U474 (N_474,N_362,N_312);
nand U475 (N_475,N_374,N_370);
and U476 (N_476,N_400,N_374);
nor U477 (N_477,N_161,N_234);
nand U478 (N_478,N_376,N_402);
nand U479 (N_479,N_364,N_416);
nand U480 (N_480,N_471,N_423);
and U481 (N_481,N_442,N_432);
nand U482 (N_482,N_433,N_454);
nand U483 (N_483,N_445,N_472);
nor U484 (N_484,N_461,N_456);
and U485 (N_485,N_421,N_470);
nor U486 (N_486,N_451,N_420);
nand U487 (N_487,N_431,N_436);
nor U488 (N_488,N_435,N_452);
nor U489 (N_489,N_434,N_466);
nor U490 (N_490,N_439,N_448);
nor U491 (N_491,N_460,N_449);
and U492 (N_492,N_440,N_457);
and U493 (N_493,N_459,N_468);
and U494 (N_494,N_426,N_474);
nor U495 (N_495,N_467,N_443);
nor U496 (N_496,N_430,N_444);
or U497 (N_497,N_478,N_458);
or U498 (N_498,N_429,N_476);
or U499 (N_499,N_463,N_424);
nand U500 (N_500,N_465,N_428);
or U501 (N_501,N_477,N_447);
and U502 (N_502,N_438,N_479);
nand U503 (N_503,N_469,N_450);
and U504 (N_504,N_473,N_441);
nand U505 (N_505,N_475,N_464);
nand U506 (N_506,N_425,N_462);
nor U507 (N_507,N_453,N_446);
or U508 (N_508,N_437,N_422);
nand U509 (N_509,N_427,N_455);
nand U510 (N_510,N_474,N_445);
and U511 (N_511,N_421,N_452);
and U512 (N_512,N_452,N_458);
nand U513 (N_513,N_479,N_458);
nor U514 (N_514,N_436,N_463);
nor U515 (N_515,N_437,N_451);
and U516 (N_516,N_438,N_421);
nand U517 (N_517,N_470,N_427);
and U518 (N_518,N_438,N_439);
and U519 (N_519,N_454,N_432);
nor U520 (N_520,N_452,N_440);
nand U521 (N_521,N_463,N_422);
nand U522 (N_522,N_452,N_455);
and U523 (N_523,N_478,N_423);
and U524 (N_524,N_472,N_454);
nand U525 (N_525,N_448,N_427);
or U526 (N_526,N_453,N_472);
and U527 (N_527,N_476,N_455);
or U528 (N_528,N_469,N_446);
or U529 (N_529,N_436,N_438);
nand U530 (N_530,N_422,N_454);
and U531 (N_531,N_443,N_463);
and U532 (N_532,N_452,N_431);
or U533 (N_533,N_474,N_468);
and U534 (N_534,N_424,N_470);
nand U535 (N_535,N_440,N_432);
nor U536 (N_536,N_437,N_431);
nand U537 (N_537,N_465,N_445);
nand U538 (N_538,N_479,N_431);
nor U539 (N_539,N_450,N_456);
and U540 (N_540,N_487,N_485);
and U541 (N_541,N_482,N_533);
and U542 (N_542,N_509,N_523);
and U543 (N_543,N_481,N_537);
nand U544 (N_544,N_489,N_522);
xor U545 (N_545,N_539,N_493);
nor U546 (N_546,N_515,N_517);
nor U547 (N_547,N_524,N_526);
nor U548 (N_548,N_505,N_507);
or U549 (N_549,N_530,N_480);
nor U550 (N_550,N_513,N_512);
nand U551 (N_551,N_501,N_492);
nor U552 (N_552,N_483,N_497);
or U553 (N_553,N_514,N_502);
or U554 (N_554,N_486,N_508);
or U555 (N_555,N_536,N_494);
nand U556 (N_556,N_511,N_519);
or U557 (N_557,N_534,N_490);
nor U558 (N_558,N_500,N_495);
nor U559 (N_559,N_520,N_503);
or U560 (N_560,N_529,N_518);
nor U561 (N_561,N_510,N_498);
nand U562 (N_562,N_528,N_499);
or U563 (N_563,N_521,N_516);
or U564 (N_564,N_496,N_525);
and U565 (N_565,N_506,N_491);
or U566 (N_566,N_527,N_532);
and U567 (N_567,N_488,N_535);
or U568 (N_568,N_504,N_484);
nor U569 (N_569,N_531,N_538);
nor U570 (N_570,N_500,N_514);
or U571 (N_571,N_516,N_497);
nand U572 (N_572,N_512,N_529);
and U573 (N_573,N_530,N_500);
or U574 (N_574,N_515,N_491);
or U575 (N_575,N_501,N_498);
nand U576 (N_576,N_515,N_489);
or U577 (N_577,N_517,N_481);
and U578 (N_578,N_489,N_492);
nand U579 (N_579,N_529,N_525);
nor U580 (N_580,N_538,N_500);
nor U581 (N_581,N_530,N_490);
and U582 (N_582,N_519,N_521);
and U583 (N_583,N_511,N_516);
or U584 (N_584,N_491,N_520);
nor U585 (N_585,N_522,N_521);
nor U586 (N_586,N_525,N_521);
nor U587 (N_587,N_535,N_505);
nand U588 (N_588,N_527,N_490);
nor U589 (N_589,N_485,N_493);
and U590 (N_590,N_522,N_523);
or U591 (N_591,N_531,N_530);
or U592 (N_592,N_518,N_522);
nand U593 (N_593,N_494,N_508);
nand U594 (N_594,N_497,N_496);
and U595 (N_595,N_506,N_527);
and U596 (N_596,N_523,N_485);
or U597 (N_597,N_498,N_500);
nand U598 (N_598,N_532,N_491);
and U599 (N_599,N_515,N_538);
nor U600 (N_600,N_572,N_570);
or U601 (N_601,N_599,N_553);
nor U602 (N_602,N_567,N_549);
nand U603 (N_603,N_544,N_598);
or U604 (N_604,N_550,N_573);
or U605 (N_605,N_583,N_593);
or U606 (N_606,N_565,N_551);
or U607 (N_607,N_552,N_554);
or U608 (N_608,N_596,N_548);
or U609 (N_609,N_558,N_546);
nor U610 (N_610,N_541,N_592);
and U611 (N_611,N_547,N_580);
and U612 (N_612,N_581,N_542);
nand U613 (N_613,N_556,N_575);
nor U614 (N_614,N_579,N_597);
and U615 (N_615,N_590,N_540);
or U616 (N_616,N_557,N_594);
nand U617 (N_617,N_568,N_574);
or U618 (N_618,N_577,N_571);
or U619 (N_619,N_588,N_589);
nand U620 (N_620,N_569,N_591);
and U621 (N_621,N_559,N_563);
and U622 (N_622,N_543,N_578);
or U623 (N_623,N_562,N_576);
and U624 (N_624,N_545,N_595);
nor U625 (N_625,N_582,N_585);
or U626 (N_626,N_560,N_561);
or U627 (N_627,N_555,N_587);
nor U628 (N_628,N_566,N_586);
or U629 (N_629,N_584,N_564);
or U630 (N_630,N_589,N_573);
or U631 (N_631,N_569,N_557);
nor U632 (N_632,N_599,N_578);
or U633 (N_633,N_551,N_588);
nor U634 (N_634,N_572,N_573);
and U635 (N_635,N_562,N_597);
and U636 (N_636,N_562,N_587);
nand U637 (N_637,N_580,N_565);
and U638 (N_638,N_587,N_568);
nand U639 (N_639,N_551,N_562);
nor U640 (N_640,N_561,N_593);
and U641 (N_641,N_575,N_561);
nor U642 (N_642,N_545,N_584);
or U643 (N_643,N_587,N_557);
nor U644 (N_644,N_568,N_559);
or U645 (N_645,N_553,N_588);
nand U646 (N_646,N_555,N_548);
and U647 (N_647,N_559,N_564);
and U648 (N_648,N_562,N_586);
xor U649 (N_649,N_597,N_574);
and U650 (N_650,N_592,N_544);
nor U651 (N_651,N_583,N_575);
nand U652 (N_652,N_569,N_585);
and U653 (N_653,N_592,N_579);
nand U654 (N_654,N_546,N_572);
or U655 (N_655,N_591,N_582);
or U656 (N_656,N_559,N_554);
or U657 (N_657,N_597,N_549);
or U658 (N_658,N_541,N_557);
nor U659 (N_659,N_547,N_578);
and U660 (N_660,N_616,N_617);
nor U661 (N_661,N_648,N_646);
xnor U662 (N_662,N_606,N_641);
or U663 (N_663,N_614,N_633);
nor U664 (N_664,N_627,N_612);
or U665 (N_665,N_649,N_621);
nor U666 (N_666,N_630,N_619);
and U667 (N_667,N_636,N_631);
nand U668 (N_668,N_622,N_659);
nand U669 (N_669,N_618,N_615);
nor U670 (N_670,N_653,N_637);
nand U671 (N_671,N_620,N_623);
nand U672 (N_672,N_647,N_654);
nor U673 (N_673,N_656,N_642);
and U674 (N_674,N_639,N_632);
or U675 (N_675,N_651,N_608);
and U676 (N_676,N_643,N_604);
nand U677 (N_677,N_640,N_628);
nand U678 (N_678,N_607,N_605);
nor U679 (N_679,N_655,N_613);
nand U680 (N_680,N_625,N_629);
nor U681 (N_681,N_650,N_602);
and U682 (N_682,N_645,N_634);
nor U683 (N_683,N_609,N_611);
and U684 (N_684,N_610,N_635);
or U685 (N_685,N_624,N_638);
nor U686 (N_686,N_657,N_644);
or U687 (N_687,N_601,N_603);
or U688 (N_688,N_652,N_626);
and U689 (N_689,N_600,N_658);
and U690 (N_690,N_637,N_624);
nor U691 (N_691,N_656,N_606);
nor U692 (N_692,N_600,N_623);
nor U693 (N_693,N_610,N_650);
and U694 (N_694,N_635,N_614);
or U695 (N_695,N_623,N_656);
or U696 (N_696,N_646,N_625);
nand U697 (N_697,N_650,N_623);
or U698 (N_698,N_648,N_629);
nand U699 (N_699,N_621,N_628);
nand U700 (N_700,N_644,N_619);
or U701 (N_701,N_603,N_616);
nor U702 (N_702,N_652,N_641);
nand U703 (N_703,N_644,N_612);
nor U704 (N_704,N_638,N_635);
and U705 (N_705,N_656,N_618);
nor U706 (N_706,N_628,N_616);
nand U707 (N_707,N_645,N_647);
nand U708 (N_708,N_626,N_633);
or U709 (N_709,N_652,N_614);
nand U710 (N_710,N_614,N_619);
and U711 (N_711,N_649,N_654);
or U712 (N_712,N_638,N_614);
nand U713 (N_713,N_642,N_658);
nor U714 (N_714,N_659,N_657);
nor U715 (N_715,N_600,N_652);
nor U716 (N_716,N_639,N_646);
nor U717 (N_717,N_658,N_641);
nor U718 (N_718,N_635,N_659);
nand U719 (N_719,N_607,N_639);
nand U720 (N_720,N_661,N_680);
nor U721 (N_721,N_688,N_682);
nor U722 (N_722,N_685,N_703);
nor U723 (N_723,N_667,N_702);
and U724 (N_724,N_676,N_719);
and U725 (N_725,N_662,N_698);
nor U726 (N_726,N_660,N_706);
nand U727 (N_727,N_677,N_673);
nor U728 (N_728,N_670,N_679);
nand U729 (N_729,N_705,N_665);
and U730 (N_730,N_697,N_674);
or U731 (N_731,N_712,N_687);
nand U732 (N_732,N_704,N_686);
and U733 (N_733,N_710,N_691);
nand U734 (N_734,N_707,N_663);
and U735 (N_735,N_684,N_681);
nand U736 (N_736,N_700,N_664);
and U737 (N_737,N_690,N_671);
nor U738 (N_738,N_717,N_714);
and U739 (N_739,N_668,N_695);
or U740 (N_740,N_699,N_716);
xnor U741 (N_741,N_693,N_672);
nand U742 (N_742,N_701,N_683);
xor U743 (N_743,N_669,N_692);
or U744 (N_744,N_696,N_711);
or U745 (N_745,N_694,N_678);
and U746 (N_746,N_715,N_666);
and U747 (N_747,N_708,N_718);
nand U748 (N_748,N_689,N_713);
nand U749 (N_749,N_675,N_709);
and U750 (N_750,N_671,N_675);
nor U751 (N_751,N_680,N_719);
and U752 (N_752,N_677,N_693);
or U753 (N_753,N_696,N_680);
nor U754 (N_754,N_719,N_708);
nand U755 (N_755,N_684,N_668);
and U756 (N_756,N_713,N_709);
or U757 (N_757,N_661,N_690);
nand U758 (N_758,N_699,N_673);
nand U759 (N_759,N_709,N_703);
nand U760 (N_760,N_695,N_675);
nand U761 (N_761,N_679,N_695);
nor U762 (N_762,N_712,N_669);
nor U763 (N_763,N_678,N_667);
and U764 (N_764,N_691,N_706);
and U765 (N_765,N_715,N_709);
xor U766 (N_766,N_691,N_699);
or U767 (N_767,N_709,N_671);
and U768 (N_768,N_690,N_717);
or U769 (N_769,N_682,N_671);
or U770 (N_770,N_680,N_717);
and U771 (N_771,N_670,N_683);
or U772 (N_772,N_710,N_662);
and U773 (N_773,N_670,N_685);
nor U774 (N_774,N_715,N_703);
or U775 (N_775,N_691,N_714);
and U776 (N_776,N_718,N_681);
and U777 (N_777,N_709,N_687);
and U778 (N_778,N_689,N_712);
nor U779 (N_779,N_707,N_719);
nand U780 (N_780,N_721,N_739);
or U781 (N_781,N_765,N_777);
nor U782 (N_782,N_748,N_746);
or U783 (N_783,N_747,N_763);
nand U784 (N_784,N_776,N_743);
or U785 (N_785,N_768,N_762);
and U786 (N_786,N_772,N_769);
or U787 (N_787,N_730,N_779);
or U788 (N_788,N_771,N_745);
nand U789 (N_789,N_727,N_756);
and U790 (N_790,N_770,N_761);
nor U791 (N_791,N_735,N_774);
and U792 (N_792,N_755,N_731);
and U793 (N_793,N_732,N_741);
and U794 (N_794,N_737,N_773);
nor U795 (N_795,N_754,N_728);
or U796 (N_796,N_723,N_742);
nor U797 (N_797,N_778,N_767);
and U798 (N_798,N_757,N_733);
nor U799 (N_799,N_740,N_738);
nor U800 (N_800,N_734,N_753);
nand U801 (N_801,N_736,N_729);
nand U802 (N_802,N_775,N_726);
and U803 (N_803,N_725,N_752);
or U804 (N_804,N_751,N_722);
nand U805 (N_805,N_749,N_760);
nand U806 (N_806,N_724,N_759);
and U807 (N_807,N_766,N_750);
and U808 (N_808,N_720,N_744);
and U809 (N_809,N_764,N_758);
or U810 (N_810,N_772,N_763);
nor U811 (N_811,N_729,N_763);
or U812 (N_812,N_753,N_727);
and U813 (N_813,N_778,N_774);
nor U814 (N_814,N_735,N_754);
or U815 (N_815,N_774,N_746);
and U816 (N_816,N_757,N_722);
nand U817 (N_817,N_726,N_770);
nor U818 (N_818,N_776,N_754);
and U819 (N_819,N_749,N_720);
nand U820 (N_820,N_754,N_751);
and U821 (N_821,N_765,N_752);
xnor U822 (N_822,N_760,N_753);
nor U823 (N_823,N_731,N_749);
and U824 (N_824,N_755,N_762);
and U825 (N_825,N_770,N_720);
nor U826 (N_826,N_750,N_775);
and U827 (N_827,N_770,N_747);
and U828 (N_828,N_754,N_777);
or U829 (N_829,N_734,N_771);
nor U830 (N_830,N_732,N_760);
nand U831 (N_831,N_763,N_750);
nand U832 (N_832,N_776,N_752);
nor U833 (N_833,N_736,N_720);
and U834 (N_834,N_722,N_730);
nor U835 (N_835,N_751,N_743);
and U836 (N_836,N_771,N_757);
or U837 (N_837,N_766,N_736);
and U838 (N_838,N_721,N_751);
nor U839 (N_839,N_746,N_728);
or U840 (N_840,N_799,N_803);
nand U841 (N_841,N_824,N_800);
nor U842 (N_842,N_780,N_788);
nand U843 (N_843,N_837,N_795);
nand U844 (N_844,N_789,N_825);
nor U845 (N_845,N_791,N_817);
nand U846 (N_846,N_797,N_782);
or U847 (N_847,N_828,N_781);
nor U848 (N_848,N_793,N_832);
xnor U849 (N_849,N_822,N_823);
nand U850 (N_850,N_812,N_818);
or U851 (N_851,N_819,N_783);
nor U852 (N_852,N_811,N_784);
or U853 (N_853,N_805,N_798);
nand U854 (N_854,N_831,N_792);
and U855 (N_855,N_826,N_786);
or U856 (N_856,N_801,N_813);
nor U857 (N_857,N_836,N_834);
and U858 (N_858,N_829,N_802);
nor U859 (N_859,N_830,N_814);
or U860 (N_860,N_809,N_833);
nor U861 (N_861,N_835,N_804);
nor U862 (N_862,N_796,N_808);
or U863 (N_863,N_785,N_806);
nor U864 (N_864,N_838,N_807);
nor U865 (N_865,N_816,N_787);
nor U866 (N_866,N_821,N_815);
nor U867 (N_867,N_790,N_794);
nor U868 (N_868,N_810,N_839);
and U869 (N_869,N_820,N_827);
nand U870 (N_870,N_837,N_807);
nand U871 (N_871,N_818,N_836);
nor U872 (N_872,N_818,N_790);
nand U873 (N_873,N_799,N_800);
or U874 (N_874,N_823,N_811);
and U875 (N_875,N_814,N_801);
and U876 (N_876,N_806,N_814);
and U877 (N_877,N_781,N_812);
nand U878 (N_878,N_786,N_791);
and U879 (N_879,N_782,N_802);
and U880 (N_880,N_812,N_837);
or U881 (N_881,N_837,N_822);
nand U882 (N_882,N_821,N_797);
or U883 (N_883,N_794,N_803);
or U884 (N_884,N_820,N_819);
or U885 (N_885,N_781,N_787);
and U886 (N_886,N_839,N_822);
nand U887 (N_887,N_827,N_791);
and U888 (N_888,N_830,N_803);
nand U889 (N_889,N_805,N_789);
nor U890 (N_890,N_838,N_834);
nand U891 (N_891,N_827,N_800);
nand U892 (N_892,N_789,N_792);
nand U893 (N_893,N_839,N_780);
or U894 (N_894,N_793,N_791);
nand U895 (N_895,N_802,N_799);
and U896 (N_896,N_819,N_807);
nand U897 (N_897,N_837,N_820);
and U898 (N_898,N_792,N_783);
and U899 (N_899,N_809,N_838);
and U900 (N_900,N_878,N_842);
nor U901 (N_901,N_855,N_858);
and U902 (N_902,N_861,N_898);
and U903 (N_903,N_856,N_844);
and U904 (N_904,N_868,N_896);
nor U905 (N_905,N_866,N_873);
nor U906 (N_906,N_899,N_877);
nor U907 (N_907,N_840,N_870);
and U908 (N_908,N_867,N_848);
and U909 (N_909,N_854,N_846);
or U910 (N_910,N_895,N_893);
nand U911 (N_911,N_845,N_871);
nand U912 (N_912,N_894,N_887);
and U913 (N_913,N_852,N_869);
nor U914 (N_914,N_892,N_843);
and U915 (N_915,N_888,N_881);
nor U916 (N_916,N_841,N_884);
nand U917 (N_917,N_885,N_863);
and U918 (N_918,N_859,N_891);
nor U919 (N_919,N_886,N_876);
nand U920 (N_920,N_860,N_890);
and U921 (N_921,N_889,N_880);
nor U922 (N_922,N_850,N_857);
nor U923 (N_923,N_882,N_879);
nor U924 (N_924,N_849,N_872);
nand U925 (N_925,N_853,N_883);
and U926 (N_926,N_874,N_847);
or U927 (N_927,N_875,N_862);
or U928 (N_928,N_897,N_851);
or U929 (N_929,N_864,N_865);
nor U930 (N_930,N_871,N_858);
nand U931 (N_931,N_874,N_855);
and U932 (N_932,N_842,N_879);
and U933 (N_933,N_895,N_881);
and U934 (N_934,N_870,N_867);
nor U935 (N_935,N_844,N_879);
and U936 (N_936,N_882,N_878);
nor U937 (N_937,N_851,N_858);
nor U938 (N_938,N_858,N_863);
or U939 (N_939,N_882,N_894);
nand U940 (N_940,N_878,N_846);
or U941 (N_941,N_899,N_876);
nand U942 (N_942,N_892,N_861);
or U943 (N_943,N_879,N_891);
nor U944 (N_944,N_861,N_878);
or U945 (N_945,N_885,N_840);
or U946 (N_946,N_856,N_892);
nand U947 (N_947,N_880,N_887);
nor U948 (N_948,N_877,N_862);
or U949 (N_949,N_896,N_841);
nand U950 (N_950,N_843,N_870);
nand U951 (N_951,N_896,N_880);
nand U952 (N_952,N_852,N_893);
nor U953 (N_953,N_876,N_853);
and U954 (N_954,N_875,N_842);
nand U955 (N_955,N_881,N_843);
and U956 (N_956,N_874,N_883);
nand U957 (N_957,N_896,N_881);
or U958 (N_958,N_850,N_896);
and U959 (N_959,N_877,N_855);
or U960 (N_960,N_948,N_922);
nor U961 (N_961,N_935,N_943);
nand U962 (N_962,N_908,N_942);
nor U963 (N_963,N_906,N_924);
nor U964 (N_964,N_911,N_950);
or U965 (N_965,N_959,N_954);
nor U966 (N_966,N_921,N_953);
nand U967 (N_967,N_917,N_947);
and U968 (N_968,N_904,N_903);
or U969 (N_969,N_956,N_910);
nand U970 (N_970,N_952,N_901);
nand U971 (N_971,N_909,N_958);
nor U972 (N_972,N_933,N_913);
or U973 (N_973,N_915,N_905);
or U974 (N_974,N_945,N_918);
nor U975 (N_975,N_929,N_944);
nor U976 (N_976,N_920,N_951);
nor U977 (N_977,N_941,N_957);
or U978 (N_978,N_923,N_900);
or U979 (N_979,N_919,N_926);
and U980 (N_980,N_912,N_946);
nor U981 (N_981,N_955,N_936);
nor U982 (N_982,N_938,N_914);
nor U983 (N_983,N_931,N_930);
and U984 (N_984,N_927,N_949);
and U985 (N_985,N_940,N_934);
nor U986 (N_986,N_932,N_939);
xnor U987 (N_987,N_902,N_925);
or U988 (N_988,N_907,N_916);
and U989 (N_989,N_937,N_928);
and U990 (N_990,N_959,N_906);
nor U991 (N_991,N_945,N_923);
nor U992 (N_992,N_901,N_928);
or U993 (N_993,N_920,N_936);
or U994 (N_994,N_929,N_901);
nand U995 (N_995,N_904,N_910);
nor U996 (N_996,N_935,N_947);
and U997 (N_997,N_939,N_951);
nor U998 (N_998,N_918,N_900);
or U999 (N_999,N_920,N_954);
and U1000 (N_1000,N_935,N_954);
nor U1001 (N_1001,N_948,N_906);
nand U1002 (N_1002,N_927,N_941);
or U1003 (N_1003,N_953,N_909);
and U1004 (N_1004,N_925,N_957);
nor U1005 (N_1005,N_945,N_907);
and U1006 (N_1006,N_953,N_912);
and U1007 (N_1007,N_900,N_916);
nor U1008 (N_1008,N_951,N_914);
or U1009 (N_1009,N_912,N_911);
or U1010 (N_1010,N_912,N_918);
nor U1011 (N_1011,N_937,N_900);
nor U1012 (N_1012,N_926,N_949);
nand U1013 (N_1013,N_938,N_924);
or U1014 (N_1014,N_915,N_916);
nand U1015 (N_1015,N_925,N_934);
and U1016 (N_1016,N_903,N_933);
or U1017 (N_1017,N_942,N_900);
and U1018 (N_1018,N_905,N_904);
nand U1019 (N_1019,N_926,N_932);
nor U1020 (N_1020,N_1013,N_981);
or U1021 (N_1021,N_969,N_992);
xor U1022 (N_1022,N_997,N_1012);
nor U1023 (N_1023,N_1018,N_1014);
nor U1024 (N_1024,N_964,N_984);
or U1025 (N_1025,N_1006,N_995);
or U1026 (N_1026,N_966,N_1005);
nor U1027 (N_1027,N_998,N_976);
nor U1028 (N_1028,N_993,N_1015);
nand U1029 (N_1029,N_987,N_973);
and U1030 (N_1030,N_965,N_961);
and U1031 (N_1031,N_968,N_974);
nand U1032 (N_1032,N_1004,N_977);
nor U1033 (N_1033,N_971,N_988);
nand U1034 (N_1034,N_985,N_1011);
or U1035 (N_1035,N_1016,N_1008);
nor U1036 (N_1036,N_994,N_982);
nor U1037 (N_1037,N_1003,N_991);
or U1038 (N_1038,N_960,N_996);
or U1039 (N_1039,N_1019,N_963);
nand U1040 (N_1040,N_1017,N_990);
nand U1041 (N_1041,N_967,N_979);
or U1042 (N_1042,N_989,N_1009);
or U1043 (N_1043,N_986,N_962);
and U1044 (N_1044,N_970,N_978);
or U1045 (N_1045,N_1010,N_980);
or U1046 (N_1046,N_1001,N_975);
nand U1047 (N_1047,N_983,N_999);
or U1048 (N_1048,N_972,N_1002);
nand U1049 (N_1049,N_1007,N_1000);
or U1050 (N_1050,N_969,N_1007);
xnor U1051 (N_1051,N_998,N_979);
and U1052 (N_1052,N_1016,N_990);
nand U1053 (N_1053,N_963,N_982);
or U1054 (N_1054,N_1002,N_992);
nor U1055 (N_1055,N_975,N_1007);
nor U1056 (N_1056,N_991,N_1005);
or U1057 (N_1057,N_999,N_1010);
and U1058 (N_1058,N_992,N_1005);
and U1059 (N_1059,N_963,N_993);
and U1060 (N_1060,N_1007,N_989);
nand U1061 (N_1061,N_984,N_979);
or U1062 (N_1062,N_982,N_981);
nand U1063 (N_1063,N_997,N_1001);
nand U1064 (N_1064,N_1013,N_969);
nand U1065 (N_1065,N_1015,N_975);
and U1066 (N_1066,N_1013,N_980);
or U1067 (N_1067,N_982,N_972);
nand U1068 (N_1068,N_986,N_999);
nand U1069 (N_1069,N_967,N_1011);
nor U1070 (N_1070,N_987,N_1015);
nor U1071 (N_1071,N_994,N_1004);
nor U1072 (N_1072,N_1000,N_985);
or U1073 (N_1073,N_971,N_1015);
or U1074 (N_1074,N_966,N_1014);
nand U1075 (N_1075,N_986,N_1003);
and U1076 (N_1076,N_1018,N_997);
and U1077 (N_1077,N_969,N_985);
or U1078 (N_1078,N_1011,N_1006);
or U1079 (N_1079,N_968,N_988);
nor U1080 (N_1080,N_1046,N_1048);
and U1081 (N_1081,N_1031,N_1077);
nand U1082 (N_1082,N_1020,N_1028);
nor U1083 (N_1083,N_1044,N_1034);
nor U1084 (N_1084,N_1026,N_1041);
and U1085 (N_1085,N_1067,N_1023);
nor U1086 (N_1086,N_1036,N_1058);
nand U1087 (N_1087,N_1055,N_1079);
nand U1088 (N_1088,N_1061,N_1065);
or U1089 (N_1089,N_1073,N_1056);
or U1090 (N_1090,N_1030,N_1039);
nor U1091 (N_1091,N_1043,N_1060);
and U1092 (N_1092,N_1064,N_1054);
nand U1093 (N_1093,N_1040,N_1024);
or U1094 (N_1094,N_1069,N_1038);
and U1095 (N_1095,N_1021,N_1042);
nor U1096 (N_1096,N_1047,N_1066);
or U1097 (N_1097,N_1052,N_1057);
and U1098 (N_1098,N_1027,N_1068);
and U1099 (N_1099,N_1076,N_1037);
and U1100 (N_1100,N_1045,N_1071);
nor U1101 (N_1101,N_1075,N_1035);
and U1102 (N_1102,N_1062,N_1070);
nand U1103 (N_1103,N_1051,N_1022);
or U1104 (N_1104,N_1032,N_1033);
nand U1105 (N_1105,N_1078,N_1025);
nor U1106 (N_1106,N_1029,N_1059);
and U1107 (N_1107,N_1074,N_1050);
and U1108 (N_1108,N_1053,N_1063);
or U1109 (N_1109,N_1049,N_1072);
nand U1110 (N_1110,N_1063,N_1025);
and U1111 (N_1111,N_1073,N_1058);
nand U1112 (N_1112,N_1046,N_1028);
nand U1113 (N_1113,N_1044,N_1078);
nor U1114 (N_1114,N_1078,N_1055);
or U1115 (N_1115,N_1024,N_1025);
and U1116 (N_1116,N_1053,N_1066);
nand U1117 (N_1117,N_1051,N_1021);
or U1118 (N_1118,N_1047,N_1022);
nand U1119 (N_1119,N_1044,N_1070);
and U1120 (N_1120,N_1059,N_1020);
nand U1121 (N_1121,N_1075,N_1070);
nand U1122 (N_1122,N_1060,N_1075);
nand U1123 (N_1123,N_1066,N_1049);
nor U1124 (N_1124,N_1058,N_1053);
nor U1125 (N_1125,N_1072,N_1023);
and U1126 (N_1126,N_1054,N_1069);
or U1127 (N_1127,N_1057,N_1040);
nand U1128 (N_1128,N_1042,N_1034);
nor U1129 (N_1129,N_1062,N_1033);
or U1130 (N_1130,N_1021,N_1044);
nor U1131 (N_1131,N_1033,N_1031);
nand U1132 (N_1132,N_1078,N_1036);
nor U1133 (N_1133,N_1075,N_1054);
nand U1134 (N_1134,N_1022,N_1062);
and U1135 (N_1135,N_1023,N_1020);
nor U1136 (N_1136,N_1044,N_1074);
and U1137 (N_1137,N_1066,N_1069);
and U1138 (N_1138,N_1078,N_1026);
nand U1139 (N_1139,N_1042,N_1043);
nand U1140 (N_1140,N_1080,N_1087);
or U1141 (N_1141,N_1083,N_1085);
and U1142 (N_1142,N_1084,N_1111);
or U1143 (N_1143,N_1088,N_1102);
and U1144 (N_1144,N_1138,N_1136);
or U1145 (N_1145,N_1125,N_1101);
nand U1146 (N_1146,N_1130,N_1115);
or U1147 (N_1147,N_1119,N_1126);
nor U1148 (N_1148,N_1127,N_1114);
or U1149 (N_1149,N_1135,N_1095);
nor U1150 (N_1150,N_1131,N_1137);
or U1151 (N_1151,N_1089,N_1090);
nor U1152 (N_1152,N_1099,N_1094);
or U1153 (N_1153,N_1105,N_1092);
or U1154 (N_1154,N_1129,N_1100);
nor U1155 (N_1155,N_1093,N_1134);
nand U1156 (N_1156,N_1123,N_1081);
or U1157 (N_1157,N_1097,N_1106);
or U1158 (N_1158,N_1116,N_1124);
or U1159 (N_1159,N_1109,N_1108);
nand U1160 (N_1160,N_1096,N_1120);
nand U1161 (N_1161,N_1113,N_1086);
or U1162 (N_1162,N_1107,N_1110);
nand U1163 (N_1163,N_1112,N_1132);
nor U1164 (N_1164,N_1091,N_1121);
or U1165 (N_1165,N_1139,N_1133);
and U1166 (N_1166,N_1104,N_1117);
nor U1167 (N_1167,N_1098,N_1122);
and U1168 (N_1168,N_1128,N_1082);
nor U1169 (N_1169,N_1118,N_1103);
and U1170 (N_1170,N_1122,N_1095);
nand U1171 (N_1171,N_1134,N_1135);
and U1172 (N_1172,N_1104,N_1135);
nor U1173 (N_1173,N_1128,N_1080);
and U1174 (N_1174,N_1108,N_1126);
nor U1175 (N_1175,N_1124,N_1114);
and U1176 (N_1176,N_1082,N_1111);
or U1177 (N_1177,N_1135,N_1107);
or U1178 (N_1178,N_1099,N_1091);
or U1179 (N_1179,N_1121,N_1133);
or U1180 (N_1180,N_1081,N_1130);
nand U1181 (N_1181,N_1090,N_1098);
nor U1182 (N_1182,N_1110,N_1136);
nand U1183 (N_1183,N_1087,N_1088);
nand U1184 (N_1184,N_1122,N_1107);
nor U1185 (N_1185,N_1124,N_1137);
or U1186 (N_1186,N_1095,N_1088);
nor U1187 (N_1187,N_1132,N_1134);
nand U1188 (N_1188,N_1119,N_1120);
nor U1189 (N_1189,N_1128,N_1098);
nor U1190 (N_1190,N_1127,N_1116);
or U1191 (N_1191,N_1138,N_1120);
or U1192 (N_1192,N_1135,N_1124);
nand U1193 (N_1193,N_1103,N_1096);
nand U1194 (N_1194,N_1125,N_1122);
nor U1195 (N_1195,N_1120,N_1128);
nand U1196 (N_1196,N_1103,N_1094);
nand U1197 (N_1197,N_1093,N_1131);
nand U1198 (N_1198,N_1109,N_1107);
and U1199 (N_1199,N_1118,N_1127);
xor U1200 (N_1200,N_1190,N_1199);
nor U1201 (N_1201,N_1168,N_1192);
or U1202 (N_1202,N_1194,N_1153);
nor U1203 (N_1203,N_1144,N_1177);
nor U1204 (N_1204,N_1175,N_1141);
and U1205 (N_1205,N_1165,N_1174);
and U1206 (N_1206,N_1156,N_1154);
nor U1207 (N_1207,N_1161,N_1181);
nand U1208 (N_1208,N_1148,N_1163);
or U1209 (N_1209,N_1158,N_1195);
or U1210 (N_1210,N_1167,N_1159);
nor U1211 (N_1211,N_1147,N_1160);
nor U1212 (N_1212,N_1185,N_1191);
nand U1213 (N_1213,N_1146,N_1157);
or U1214 (N_1214,N_1184,N_1178);
or U1215 (N_1215,N_1152,N_1172);
or U1216 (N_1216,N_1169,N_1189);
nor U1217 (N_1217,N_1182,N_1196);
or U1218 (N_1218,N_1193,N_1151);
or U1219 (N_1219,N_1179,N_1149);
nor U1220 (N_1220,N_1173,N_1143);
and U1221 (N_1221,N_1188,N_1171);
or U1222 (N_1222,N_1180,N_1197);
or U1223 (N_1223,N_1187,N_1164);
nor U1224 (N_1224,N_1170,N_1142);
and U1225 (N_1225,N_1183,N_1162);
and U1226 (N_1226,N_1198,N_1140);
or U1227 (N_1227,N_1186,N_1176);
nand U1228 (N_1228,N_1166,N_1150);
or U1229 (N_1229,N_1155,N_1145);
nand U1230 (N_1230,N_1176,N_1178);
and U1231 (N_1231,N_1165,N_1157);
nand U1232 (N_1232,N_1189,N_1196);
and U1233 (N_1233,N_1198,N_1196);
and U1234 (N_1234,N_1188,N_1146);
and U1235 (N_1235,N_1177,N_1181);
nor U1236 (N_1236,N_1154,N_1174);
nor U1237 (N_1237,N_1185,N_1184);
or U1238 (N_1238,N_1166,N_1183);
nand U1239 (N_1239,N_1184,N_1181);
nand U1240 (N_1240,N_1162,N_1168);
nand U1241 (N_1241,N_1196,N_1194);
nand U1242 (N_1242,N_1146,N_1166);
nand U1243 (N_1243,N_1147,N_1140);
nor U1244 (N_1244,N_1168,N_1145);
nor U1245 (N_1245,N_1149,N_1174);
nor U1246 (N_1246,N_1175,N_1176);
nand U1247 (N_1247,N_1192,N_1151);
and U1248 (N_1248,N_1161,N_1185);
or U1249 (N_1249,N_1193,N_1158);
or U1250 (N_1250,N_1171,N_1184);
nor U1251 (N_1251,N_1151,N_1164);
and U1252 (N_1252,N_1144,N_1150);
nand U1253 (N_1253,N_1152,N_1151);
and U1254 (N_1254,N_1141,N_1151);
nand U1255 (N_1255,N_1175,N_1143);
nor U1256 (N_1256,N_1168,N_1193);
and U1257 (N_1257,N_1187,N_1195);
or U1258 (N_1258,N_1160,N_1167);
xor U1259 (N_1259,N_1157,N_1156);
nor U1260 (N_1260,N_1251,N_1221);
and U1261 (N_1261,N_1246,N_1235);
nor U1262 (N_1262,N_1208,N_1209);
nand U1263 (N_1263,N_1258,N_1256);
or U1264 (N_1264,N_1249,N_1201);
or U1265 (N_1265,N_1237,N_1259);
nor U1266 (N_1266,N_1229,N_1206);
nand U1267 (N_1267,N_1217,N_1213);
nor U1268 (N_1268,N_1212,N_1211);
nor U1269 (N_1269,N_1216,N_1226);
nor U1270 (N_1270,N_1245,N_1253);
and U1271 (N_1271,N_1215,N_1203);
or U1272 (N_1272,N_1204,N_1244);
nand U1273 (N_1273,N_1202,N_1205);
or U1274 (N_1274,N_1233,N_1223);
nor U1275 (N_1275,N_1222,N_1231);
nand U1276 (N_1276,N_1230,N_1254);
nor U1277 (N_1277,N_1224,N_1214);
nor U1278 (N_1278,N_1234,N_1238);
nand U1279 (N_1279,N_1257,N_1248);
or U1280 (N_1280,N_1247,N_1236);
or U1281 (N_1281,N_1243,N_1250);
nand U1282 (N_1282,N_1255,N_1252);
or U1283 (N_1283,N_1218,N_1241);
nand U1284 (N_1284,N_1240,N_1227);
nor U1285 (N_1285,N_1219,N_1232);
nand U1286 (N_1286,N_1225,N_1220);
nor U1287 (N_1287,N_1228,N_1207);
nor U1288 (N_1288,N_1239,N_1210);
or U1289 (N_1289,N_1200,N_1242);
nor U1290 (N_1290,N_1229,N_1257);
and U1291 (N_1291,N_1235,N_1217);
and U1292 (N_1292,N_1213,N_1222);
xor U1293 (N_1293,N_1206,N_1235);
nand U1294 (N_1294,N_1230,N_1229);
nand U1295 (N_1295,N_1237,N_1226);
or U1296 (N_1296,N_1246,N_1220);
or U1297 (N_1297,N_1250,N_1206);
xnor U1298 (N_1298,N_1202,N_1247);
nor U1299 (N_1299,N_1248,N_1223);
or U1300 (N_1300,N_1252,N_1237);
nor U1301 (N_1301,N_1213,N_1203);
and U1302 (N_1302,N_1255,N_1205);
and U1303 (N_1303,N_1229,N_1204);
and U1304 (N_1304,N_1204,N_1237);
or U1305 (N_1305,N_1233,N_1239);
nor U1306 (N_1306,N_1208,N_1207);
nor U1307 (N_1307,N_1234,N_1229);
nor U1308 (N_1308,N_1242,N_1248);
and U1309 (N_1309,N_1238,N_1246);
nor U1310 (N_1310,N_1222,N_1201);
xor U1311 (N_1311,N_1247,N_1204);
or U1312 (N_1312,N_1256,N_1221);
and U1313 (N_1313,N_1238,N_1218);
or U1314 (N_1314,N_1255,N_1208);
and U1315 (N_1315,N_1258,N_1220);
nand U1316 (N_1316,N_1226,N_1204);
or U1317 (N_1317,N_1245,N_1203);
and U1318 (N_1318,N_1202,N_1242);
nand U1319 (N_1319,N_1226,N_1234);
nor U1320 (N_1320,N_1268,N_1294);
nor U1321 (N_1321,N_1278,N_1272);
or U1322 (N_1322,N_1312,N_1270);
or U1323 (N_1323,N_1296,N_1288);
and U1324 (N_1324,N_1262,N_1297);
and U1325 (N_1325,N_1314,N_1260);
or U1326 (N_1326,N_1275,N_1265);
and U1327 (N_1327,N_1307,N_1295);
xor U1328 (N_1328,N_1281,N_1290);
nor U1329 (N_1329,N_1309,N_1292);
or U1330 (N_1330,N_1313,N_1264);
or U1331 (N_1331,N_1277,N_1293);
nand U1332 (N_1332,N_1305,N_1274);
or U1333 (N_1333,N_1315,N_1283);
or U1334 (N_1334,N_1300,N_1291);
nor U1335 (N_1335,N_1303,N_1289);
nand U1336 (N_1336,N_1282,N_1304);
nor U1337 (N_1337,N_1298,N_1311);
or U1338 (N_1338,N_1269,N_1261);
nor U1339 (N_1339,N_1310,N_1308);
nor U1340 (N_1340,N_1271,N_1273);
and U1341 (N_1341,N_1266,N_1263);
or U1342 (N_1342,N_1299,N_1276);
and U1343 (N_1343,N_1284,N_1267);
nor U1344 (N_1344,N_1318,N_1285);
or U1345 (N_1345,N_1286,N_1302);
nor U1346 (N_1346,N_1301,N_1317);
nand U1347 (N_1347,N_1280,N_1306);
nor U1348 (N_1348,N_1279,N_1316);
and U1349 (N_1349,N_1287,N_1319);
and U1350 (N_1350,N_1306,N_1301);
or U1351 (N_1351,N_1298,N_1260);
nand U1352 (N_1352,N_1283,N_1313);
nor U1353 (N_1353,N_1268,N_1301);
nand U1354 (N_1354,N_1316,N_1277);
or U1355 (N_1355,N_1277,N_1296);
or U1356 (N_1356,N_1266,N_1270);
nand U1357 (N_1357,N_1299,N_1262);
or U1358 (N_1358,N_1304,N_1313);
or U1359 (N_1359,N_1300,N_1282);
nor U1360 (N_1360,N_1295,N_1281);
nor U1361 (N_1361,N_1305,N_1262);
or U1362 (N_1362,N_1291,N_1269);
nand U1363 (N_1363,N_1276,N_1271);
nand U1364 (N_1364,N_1278,N_1292);
and U1365 (N_1365,N_1312,N_1316);
nor U1366 (N_1366,N_1277,N_1297);
or U1367 (N_1367,N_1309,N_1269);
nor U1368 (N_1368,N_1307,N_1318);
nand U1369 (N_1369,N_1266,N_1302);
nor U1370 (N_1370,N_1284,N_1302);
xnor U1371 (N_1371,N_1287,N_1286);
or U1372 (N_1372,N_1272,N_1291);
nor U1373 (N_1373,N_1287,N_1263);
nor U1374 (N_1374,N_1289,N_1279);
nand U1375 (N_1375,N_1281,N_1287);
and U1376 (N_1376,N_1275,N_1309);
nand U1377 (N_1377,N_1311,N_1306);
or U1378 (N_1378,N_1281,N_1271);
nor U1379 (N_1379,N_1293,N_1313);
or U1380 (N_1380,N_1326,N_1345);
and U1381 (N_1381,N_1371,N_1372);
nor U1382 (N_1382,N_1349,N_1357);
xor U1383 (N_1383,N_1330,N_1377);
nor U1384 (N_1384,N_1351,N_1361);
nand U1385 (N_1385,N_1346,N_1344);
nand U1386 (N_1386,N_1343,N_1334);
nor U1387 (N_1387,N_1329,N_1374);
nand U1388 (N_1388,N_1375,N_1337);
nand U1389 (N_1389,N_1333,N_1358);
nor U1390 (N_1390,N_1379,N_1339);
and U1391 (N_1391,N_1367,N_1323);
nand U1392 (N_1392,N_1340,N_1360);
nor U1393 (N_1393,N_1369,N_1321);
or U1394 (N_1394,N_1370,N_1368);
nor U1395 (N_1395,N_1362,N_1354);
nor U1396 (N_1396,N_1327,N_1335);
and U1397 (N_1397,N_1365,N_1363);
or U1398 (N_1398,N_1325,N_1366);
nand U1399 (N_1399,N_1324,N_1338);
and U1400 (N_1400,N_1320,N_1373);
or U1401 (N_1401,N_1347,N_1350);
and U1402 (N_1402,N_1332,N_1352);
nand U1403 (N_1403,N_1355,N_1341);
nor U1404 (N_1404,N_1322,N_1348);
or U1405 (N_1405,N_1376,N_1359);
or U1406 (N_1406,N_1331,N_1353);
or U1407 (N_1407,N_1356,N_1336);
and U1408 (N_1408,N_1364,N_1342);
nand U1409 (N_1409,N_1328,N_1378);
nand U1410 (N_1410,N_1321,N_1324);
nor U1411 (N_1411,N_1369,N_1350);
or U1412 (N_1412,N_1321,N_1371);
and U1413 (N_1413,N_1356,N_1370);
nor U1414 (N_1414,N_1321,N_1358);
and U1415 (N_1415,N_1362,N_1359);
nor U1416 (N_1416,N_1320,N_1330);
nor U1417 (N_1417,N_1370,N_1353);
or U1418 (N_1418,N_1373,N_1330);
and U1419 (N_1419,N_1343,N_1369);
and U1420 (N_1420,N_1326,N_1346);
nand U1421 (N_1421,N_1370,N_1326);
or U1422 (N_1422,N_1363,N_1354);
xnor U1423 (N_1423,N_1320,N_1351);
nor U1424 (N_1424,N_1328,N_1372);
nor U1425 (N_1425,N_1356,N_1369);
and U1426 (N_1426,N_1354,N_1346);
nor U1427 (N_1427,N_1357,N_1370);
nor U1428 (N_1428,N_1323,N_1329);
nand U1429 (N_1429,N_1350,N_1341);
nor U1430 (N_1430,N_1325,N_1373);
and U1431 (N_1431,N_1347,N_1320);
nand U1432 (N_1432,N_1330,N_1364);
or U1433 (N_1433,N_1329,N_1350);
or U1434 (N_1434,N_1344,N_1329);
nand U1435 (N_1435,N_1358,N_1376);
nor U1436 (N_1436,N_1327,N_1338);
or U1437 (N_1437,N_1371,N_1320);
nand U1438 (N_1438,N_1359,N_1332);
or U1439 (N_1439,N_1339,N_1373);
or U1440 (N_1440,N_1429,N_1418);
and U1441 (N_1441,N_1411,N_1438);
nand U1442 (N_1442,N_1414,N_1409);
and U1443 (N_1443,N_1401,N_1435);
nor U1444 (N_1444,N_1400,N_1384);
nor U1445 (N_1445,N_1382,N_1419);
nand U1446 (N_1446,N_1393,N_1433);
or U1447 (N_1447,N_1437,N_1416);
or U1448 (N_1448,N_1407,N_1391);
or U1449 (N_1449,N_1422,N_1389);
nor U1450 (N_1450,N_1420,N_1388);
or U1451 (N_1451,N_1417,N_1415);
or U1452 (N_1452,N_1404,N_1402);
nand U1453 (N_1453,N_1430,N_1408);
and U1454 (N_1454,N_1403,N_1381);
and U1455 (N_1455,N_1392,N_1439);
and U1456 (N_1456,N_1398,N_1412);
and U1457 (N_1457,N_1406,N_1386);
nor U1458 (N_1458,N_1399,N_1413);
or U1459 (N_1459,N_1396,N_1383);
or U1460 (N_1460,N_1436,N_1432);
nand U1461 (N_1461,N_1427,N_1410);
or U1462 (N_1462,N_1387,N_1431);
or U1463 (N_1463,N_1434,N_1421);
and U1464 (N_1464,N_1397,N_1394);
nor U1465 (N_1465,N_1428,N_1423);
nor U1466 (N_1466,N_1385,N_1426);
or U1467 (N_1467,N_1395,N_1405);
or U1468 (N_1468,N_1380,N_1425);
nor U1469 (N_1469,N_1390,N_1424);
or U1470 (N_1470,N_1390,N_1386);
or U1471 (N_1471,N_1391,N_1439);
and U1472 (N_1472,N_1398,N_1402);
nand U1473 (N_1473,N_1389,N_1384);
and U1474 (N_1474,N_1424,N_1433);
or U1475 (N_1475,N_1396,N_1431);
nand U1476 (N_1476,N_1418,N_1423);
or U1477 (N_1477,N_1407,N_1386);
xnor U1478 (N_1478,N_1381,N_1436);
or U1479 (N_1479,N_1405,N_1424);
nand U1480 (N_1480,N_1390,N_1380);
nand U1481 (N_1481,N_1409,N_1426);
nor U1482 (N_1482,N_1435,N_1402);
or U1483 (N_1483,N_1413,N_1402);
nand U1484 (N_1484,N_1404,N_1406);
nand U1485 (N_1485,N_1424,N_1381);
or U1486 (N_1486,N_1384,N_1383);
or U1487 (N_1487,N_1435,N_1392);
nor U1488 (N_1488,N_1433,N_1434);
nand U1489 (N_1489,N_1394,N_1393);
nand U1490 (N_1490,N_1428,N_1397);
nand U1491 (N_1491,N_1393,N_1384);
or U1492 (N_1492,N_1397,N_1396);
and U1493 (N_1493,N_1406,N_1423);
or U1494 (N_1494,N_1398,N_1432);
and U1495 (N_1495,N_1407,N_1412);
and U1496 (N_1496,N_1406,N_1405);
nor U1497 (N_1497,N_1380,N_1398);
or U1498 (N_1498,N_1403,N_1397);
or U1499 (N_1499,N_1381,N_1409);
and U1500 (N_1500,N_1495,N_1499);
or U1501 (N_1501,N_1452,N_1465);
and U1502 (N_1502,N_1448,N_1444);
nand U1503 (N_1503,N_1443,N_1455);
nand U1504 (N_1504,N_1459,N_1476);
and U1505 (N_1505,N_1450,N_1486);
xnor U1506 (N_1506,N_1487,N_1471);
nand U1507 (N_1507,N_1496,N_1470);
and U1508 (N_1508,N_1480,N_1493);
and U1509 (N_1509,N_1447,N_1457);
and U1510 (N_1510,N_1492,N_1474);
and U1511 (N_1511,N_1484,N_1466);
and U1512 (N_1512,N_1485,N_1478);
or U1513 (N_1513,N_1491,N_1445);
and U1514 (N_1514,N_1473,N_1441);
or U1515 (N_1515,N_1482,N_1475);
nand U1516 (N_1516,N_1467,N_1458);
and U1517 (N_1517,N_1481,N_1464);
or U1518 (N_1518,N_1456,N_1461);
nor U1519 (N_1519,N_1454,N_1483);
nor U1520 (N_1520,N_1469,N_1490);
nor U1521 (N_1521,N_1489,N_1462);
or U1522 (N_1522,N_1479,N_1463);
or U1523 (N_1523,N_1442,N_1472);
and U1524 (N_1524,N_1453,N_1468);
nand U1525 (N_1525,N_1497,N_1446);
nand U1526 (N_1526,N_1449,N_1477);
nand U1527 (N_1527,N_1451,N_1498);
or U1528 (N_1528,N_1494,N_1460);
or U1529 (N_1529,N_1440,N_1488);
or U1530 (N_1530,N_1444,N_1450);
nor U1531 (N_1531,N_1452,N_1476);
nor U1532 (N_1532,N_1446,N_1499);
nor U1533 (N_1533,N_1468,N_1491);
nor U1534 (N_1534,N_1486,N_1481);
or U1535 (N_1535,N_1486,N_1482);
nand U1536 (N_1536,N_1492,N_1457);
or U1537 (N_1537,N_1498,N_1450);
nor U1538 (N_1538,N_1443,N_1487);
nand U1539 (N_1539,N_1444,N_1479);
or U1540 (N_1540,N_1491,N_1462);
and U1541 (N_1541,N_1463,N_1466);
or U1542 (N_1542,N_1498,N_1460);
nor U1543 (N_1543,N_1464,N_1448);
nor U1544 (N_1544,N_1467,N_1453);
or U1545 (N_1545,N_1441,N_1468);
nand U1546 (N_1546,N_1483,N_1456);
nand U1547 (N_1547,N_1448,N_1473);
and U1548 (N_1548,N_1484,N_1447);
nor U1549 (N_1549,N_1480,N_1460);
nor U1550 (N_1550,N_1471,N_1494);
nor U1551 (N_1551,N_1491,N_1495);
or U1552 (N_1552,N_1483,N_1498);
nand U1553 (N_1553,N_1489,N_1484);
nand U1554 (N_1554,N_1446,N_1493);
or U1555 (N_1555,N_1453,N_1464);
or U1556 (N_1556,N_1455,N_1483);
nor U1557 (N_1557,N_1487,N_1473);
nand U1558 (N_1558,N_1464,N_1463);
nor U1559 (N_1559,N_1488,N_1441);
nor U1560 (N_1560,N_1512,N_1524);
and U1561 (N_1561,N_1542,N_1523);
nand U1562 (N_1562,N_1549,N_1553);
or U1563 (N_1563,N_1547,N_1551);
and U1564 (N_1564,N_1529,N_1509);
or U1565 (N_1565,N_1508,N_1535);
and U1566 (N_1566,N_1504,N_1552);
nand U1567 (N_1567,N_1503,N_1555);
and U1568 (N_1568,N_1525,N_1505);
and U1569 (N_1569,N_1528,N_1516);
nor U1570 (N_1570,N_1536,N_1537);
nor U1571 (N_1571,N_1514,N_1500);
nand U1572 (N_1572,N_1550,N_1545);
nor U1573 (N_1573,N_1520,N_1518);
nand U1574 (N_1574,N_1515,N_1519);
or U1575 (N_1575,N_1539,N_1513);
xnor U1576 (N_1576,N_1527,N_1538);
nand U1577 (N_1577,N_1506,N_1511);
nand U1578 (N_1578,N_1559,N_1501);
nor U1579 (N_1579,N_1532,N_1534);
and U1580 (N_1580,N_1530,N_1546);
nand U1581 (N_1581,N_1557,N_1517);
nor U1582 (N_1582,N_1543,N_1558);
nand U1583 (N_1583,N_1521,N_1507);
or U1584 (N_1584,N_1502,N_1554);
nand U1585 (N_1585,N_1531,N_1533);
or U1586 (N_1586,N_1541,N_1510);
nor U1587 (N_1587,N_1522,N_1526);
nor U1588 (N_1588,N_1544,N_1540);
nor U1589 (N_1589,N_1548,N_1556);
nand U1590 (N_1590,N_1505,N_1507);
and U1591 (N_1591,N_1544,N_1541);
and U1592 (N_1592,N_1534,N_1526);
nand U1593 (N_1593,N_1510,N_1548);
and U1594 (N_1594,N_1559,N_1505);
or U1595 (N_1595,N_1551,N_1505);
nand U1596 (N_1596,N_1508,N_1556);
nor U1597 (N_1597,N_1539,N_1554);
nand U1598 (N_1598,N_1515,N_1508);
nor U1599 (N_1599,N_1533,N_1512);
nand U1600 (N_1600,N_1535,N_1521);
nor U1601 (N_1601,N_1519,N_1511);
nand U1602 (N_1602,N_1510,N_1558);
or U1603 (N_1603,N_1549,N_1547);
nand U1604 (N_1604,N_1501,N_1557);
or U1605 (N_1605,N_1553,N_1513);
nor U1606 (N_1606,N_1539,N_1544);
nor U1607 (N_1607,N_1531,N_1520);
nor U1608 (N_1608,N_1554,N_1543);
nand U1609 (N_1609,N_1543,N_1516);
nand U1610 (N_1610,N_1536,N_1510);
nand U1611 (N_1611,N_1525,N_1535);
and U1612 (N_1612,N_1523,N_1530);
or U1613 (N_1613,N_1547,N_1507);
nand U1614 (N_1614,N_1552,N_1553);
nand U1615 (N_1615,N_1509,N_1536);
nor U1616 (N_1616,N_1509,N_1518);
and U1617 (N_1617,N_1523,N_1532);
nand U1618 (N_1618,N_1502,N_1551);
nor U1619 (N_1619,N_1515,N_1523);
and U1620 (N_1620,N_1574,N_1608);
nand U1621 (N_1621,N_1606,N_1616);
nor U1622 (N_1622,N_1577,N_1570);
nand U1623 (N_1623,N_1578,N_1593);
nor U1624 (N_1624,N_1618,N_1605);
nor U1625 (N_1625,N_1564,N_1568);
and U1626 (N_1626,N_1612,N_1599);
nor U1627 (N_1627,N_1600,N_1586);
or U1628 (N_1628,N_1596,N_1585);
or U1629 (N_1629,N_1573,N_1607);
nor U1630 (N_1630,N_1604,N_1571);
nand U1631 (N_1631,N_1584,N_1610);
nand U1632 (N_1632,N_1566,N_1562);
or U1633 (N_1633,N_1576,N_1592);
and U1634 (N_1634,N_1595,N_1619);
nand U1635 (N_1635,N_1565,N_1583);
nor U1636 (N_1636,N_1582,N_1589);
and U1637 (N_1637,N_1598,N_1617);
nand U1638 (N_1638,N_1560,N_1597);
nand U1639 (N_1639,N_1572,N_1613);
or U1640 (N_1640,N_1561,N_1594);
and U1641 (N_1641,N_1563,N_1614);
nor U1642 (N_1642,N_1579,N_1581);
xnor U1643 (N_1643,N_1609,N_1588);
nor U1644 (N_1644,N_1615,N_1580);
nand U1645 (N_1645,N_1569,N_1590);
nor U1646 (N_1646,N_1611,N_1601);
or U1647 (N_1647,N_1603,N_1567);
and U1648 (N_1648,N_1587,N_1575);
nor U1649 (N_1649,N_1602,N_1591);
or U1650 (N_1650,N_1610,N_1598);
or U1651 (N_1651,N_1570,N_1600);
nor U1652 (N_1652,N_1570,N_1599);
and U1653 (N_1653,N_1574,N_1587);
and U1654 (N_1654,N_1592,N_1608);
and U1655 (N_1655,N_1581,N_1588);
or U1656 (N_1656,N_1581,N_1595);
and U1657 (N_1657,N_1585,N_1586);
or U1658 (N_1658,N_1585,N_1612);
nand U1659 (N_1659,N_1568,N_1562);
or U1660 (N_1660,N_1569,N_1587);
nand U1661 (N_1661,N_1616,N_1599);
nor U1662 (N_1662,N_1615,N_1599);
and U1663 (N_1663,N_1574,N_1616);
or U1664 (N_1664,N_1573,N_1569);
nand U1665 (N_1665,N_1565,N_1603);
or U1666 (N_1666,N_1562,N_1603);
nor U1667 (N_1667,N_1585,N_1563);
or U1668 (N_1668,N_1582,N_1596);
and U1669 (N_1669,N_1575,N_1562);
and U1670 (N_1670,N_1590,N_1601);
and U1671 (N_1671,N_1593,N_1610);
and U1672 (N_1672,N_1568,N_1579);
or U1673 (N_1673,N_1604,N_1602);
nand U1674 (N_1674,N_1571,N_1564);
and U1675 (N_1675,N_1608,N_1601);
nand U1676 (N_1676,N_1578,N_1572);
nor U1677 (N_1677,N_1577,N_1584);
nor U1678 (N_1678,N_1612,N_1575);
and U1679 (N_1679,N_1598,N_1602);
nor U1680 (N_1680,N_1654,N_1660);
nand U1681 (N_1681,N_1649,N_1626);
nor U1682 (N_1682,N_1663,N_1635);
or U1683 (N_1683,N_1627,N_1664);
and U1684 (N_1684,N_1653,N_1668);
and U1685 (N_1685,N_1655,N_1644);
nor U1686 (N_1686,N_1623,N_1670);
nand U1687 (N_1687,N_1677,N_1630);
and U1688 (N_1688,N_1628,N_1639);
or U1689 (N_1689,N_1666,N_1632);
nand U1690 (N_1690,N_1641,N_1678);
or U1691 (N_1691,N_1650,N_1661);
nor U1692 (N_1692,N_1624,N_1642);
nor U1693 (N_1693,N_1636,N_1667);
and U1694 (N_1694,N_1659,N_1629);
nand U1695 (N_1695,N_1648,N_1676);
and U1696 (N_1696,N_1662,N_1675);
or U1697 (N_1697,N_1631,N_1679);
or U1698 (N_1698,N_1634,N_1625);
xor U1699 (N_1699,N_1640,N_1637);
nor U1700 (N_1700,N_1671,N_1621);
nor U1701 (N_1701,N_1665,N_1622);
nand U1702 (N_1702,N_1651,N_1645);
nor U1703 (N_1703,N_1647,N_1633);
or U1704 (N_1704,N_1657,N_1643);
nor U1705 (N_1705,N_1673,N_1652);
nand U1706 (N_1706,N_1672,N_1620);
nor U1707 (N_1707,N_1674,N_1656);
and U1708 (N_1708,N_1638,N_1658);
nor U1709 (N_1709,N_1646,N_1669);
or U1710 (N_1710,N_1659,N_1654);
nand U1711 (N_1711,N_1633,N_1663);
or U1712 (N_1712,N_1622,N_1644);
nand U1713 (N_1713,N_1637,N_1648);
nor U1714 (N_1714,N_1658,N_1657);
or U1715 (N_1715,N_1666,N_1674);
and U1716 (N_1716,N_1632,N_1631);
and U1717 (N_1717,N_1623,N_1638);
and U1718 (N_1718,N_1661,N_1633);
nand U1719 (N_1719,N_1631,N_1647);
and U1720 (N_1720,N_1643,N_1677);
nand U1721 (N_1721,N_1649,N_1648);
nor U1722 (N_1722,N_1638,N_1629);
or U1723 (N_1723,N_1653,N_1624);
nor U1724 (N_1724,N_1657,N_1647);
nand U1725 (N_1725,N_1622,N_1675);
or U1726 (N_1726,N_1657,N_1638);
nand U1727 (N_1727,N_1649,N_1670);
and U1728 (N_1728,N_1652,N_1629);
and U1729 (N_1729,N_1632,N_1670);
and U1730 (N_1730,N_1674,N_1649);
and U1731 (N_1731,N_1621,N_1644);
nor U1732 (N_1732,N_1678,N_1655);
or U1733 (N_1733,N_1677,N_1648);
nand U1734 (N_1734,N_1624,N_1673);
nand U1735 (N_1735,N_1640,N_1666);
nor U1736 (N_1736,N_1650,N_1628);
and U1737 (N_1737,N_1664,N_1628);
or U1738 (N_1738,N_1635,N_1623);
or U1739 (N_1739,N_1642,N_1666);
and U1740 (N_1740,N_1681,N_1697);
and U1741 (N_1741,N_1729,N_1682);
nand U1742 (N_1742,N_1716,N_1734);
or U1743 (N_1743,N_1703,N_1705);
or U1744 (N_1744,N_1684,N_1689);
and U1745 (N_1745,N_1690,N_1724);
or U1746 (N_1746,N_1718,N_1738);
nor U1747 (N_1747,N_1727,N_1687);
nor U1748 (N_1748,N_1706,N_1691);
nor U1749 (N_1749,N_1728,N_1685);
and U1750 (N_1750,N_1707,N_1715);
nor U1751 (N_1751,N_1726,N_1704);
or U1752 (N_1752,N_1702,N_1725);
and U1753 (N_1753,N_1710,N_1711);
and U1754 (N_1754,N_1719,N_1721);
nand U1755 (N_1755,N_1730,N_1722);
or U1756 (N_1756,N_1680,N_1709);
nor U1757 (N_1757,N_1739,N_1737);
and U1758 (N_1758,N_1701,N_1712);
and U1759 (N_1759,N_1694,N_1735);
and U1760 (N_1760,N_1700,N_1732);
nor U1761 (N_1761,N_1736,N_1699);
nor U1762 (N_1762,N_1692,N_1695);
nand U1763 (N_1763,N_1688,N_1713);
nor U1764 (N_1764,N_1717,N_1683);
nor U1765 (N_1765,N_1696,N_1714);
nand U1766 (N_1766,N_1733,N_1686);
nor U1767 (N_1767,N_1723,N_1731);
and U1768 (N_1768,N_1693,N_1698);
or U1769 (N_1769,N_1720,N_1708);
nand U1770 (N_1770,N_1730,N_1694);
and U1771 (N_1771,N_1711,N_1704);
nor U1772 (N_1772,N_1680,N_1717);
and U1773 (N_1773,N_1697,N_1703);
nand U1774 (N_1774,N_1700,N_1713);
nor U1775 (N_1775,N_1719,N_1686);
nor U1776 (N_1776,N_1739,N_1716);
and U1777 (N_1777,N_1723,N_1725);
or U1778 (N_1778,N_1688,N_1705);
nand U1779 (N_1779,N_1715,N_1696);
nor U1780 (N_1780,N_1694,N_1727);
or U1781 (N_1781,N_1720,N_1681);
and U1782 (N_1782,N_1685,N_1719);
nor U1783 (N_1783,N_1702,N_1684);
and U1784 (N_1784,N_1686,N_1699);
nor U1785 (N_1785,N_1716,N_1685);
or U1786 (N_1786,N_1684,N_1728);
and U1787 (N_1787,N_1731,N_1681);
and U1788 (N_1788,N_1692,N_1717);
nand U1789 (N_1789,N_1704,N_1732);
xor U1790 (N_1790,N_1689,N_1681);
nand U1791 (N_1791,N_1688,N_1715);
or U1792 (N_1792,N_1694,N_1681);
and U1793 (N_1793,N_1732,N_1696);
nor U1794 (N_1794,N_1684,N_1695);
nor U1795 (N_1795,N_1700,N_1719);
or U1796 (N_1796,N_1709,N_1714);
and U1797 (N_1797,N_1696,N_1730);
nand U1798 (N_1798,N_1688,N_1700);
and U1799 (N_1799,N_1713,N_1684);
nor U1800 (N_1800,N_1799,N_1793);
and U1801 (N_1801,N_1777,N_1740);
and U1802 (N_1802,N_1765,N_1798);
nand U1803 (N_1803,N_1773,N_1779);
nand U1804 (N_1804,N_1762,N_1778);
and U1805 (N_1805,N_1797,N_1788);
or U1806 (N_1806,N_1783,N_1792);
nor U1807 (N_1807,N_1780,N_1770);
nor U1808 (N_1808,N_1744,N_1787);
and U1809 (N_1809,N_1761,N_1766);
and U1810 (N_1810,N_1791,N_1742);
and U1811 (N_1811,N_1747,N_1784);
nand U1812 (N_1812,N_1782,N_1767);
or U1813 (N_1813,N_1794,N_1785);
or U1814 (N_1814,N_1781,N_1790);
nor U1815 (N_1815,N_1789,N_1776);
or U1816 (N_1816,N_1764,N_1772);
nand U1817 (N_1817,N_1755,N_1749);
and U1818 (N_1818,N_1754,N_1753);
xnor U1819 (N_1819,N_1775,N_1795);
nand U1820 (N_1820,N_1786,N_1746);
or U1821 (N_1821,N_1751,N_1745);
and U1822 (N_1822,N_1741,N_1748);
nor U1823 (N_1823,N_1774,N_1763);
or U1824 (N_1824,N_1768,N_1760);
or U1825 (N_1825,N_1771,N_1757);
or U1826 (N_1826,N_1796,N_1756);
nor U1827 (N_1827,N_1752,N_1758);
or U1828 (N_1828,N_1759,N_1743);
and U1829 (N_1829,N_1769,N_1750);
or U1830 (N_1830,N_1758,N_1794);
nor U1831 (N_1831,N_1788,N_1751);
nor U1832 (N_1832,N_1751,N_1758);
nand U1833 (N_1833,N_1752,N_1745);
and U1834 (N_1834,N_1791,N_1789);
nor U1835 (N_1835,N_1765,N_1764);
nand U1836 (N_1836,N_1767,N_1771);
and U1837 (N_1837,N_1753,N_1798);
and U1838 (N_1838,N_1754,N_1750);
nor U1839 (N_1839,N_1759,N_1790);
and U1840 (N_1840,N_1766,N_1774);
and U1841 (N_1841,N_1799,N_1757);
nor U1842 (N_1842,N_1745,N_1778);
nor U1843 (N_1843,N_1756,N_1743);
and U1844 (N_1844,N_1771,N_1752);
nand U1845 (N_1845,N_1753,N_1770);
and U1846 (N_1846,N_1795,N_1766);
nor U1847 (N_1847,N_1756,N_1761);
nand U1848 (N_1848,N_1770,N_1745);
and U1849 (N_1849,N_1780,N_1787);
nor U1850 (N_1850,N_1789,N_1795);
nand U1851 (N_1851,N_1782,N_1783);
nor U1852 (N_1852,N_1784,N_1742);
nand U1853 (N_1853,N_1777,N_1754);
or U1854 (N_1854,N_1748,N_1764);
nand U1855 (N_1855,N_1750,N_1742);
nand U1856 (N_1856,N_1798,N_1785);
and U1857 (N_1857,N_1770,N_1776);
or U1858 (N_1858,N_1790,N_1750);
or U1859 (N_1859,N_1760,N_1755);
nand U1860 (N_1860,N_1851,N_1823);
and U1861 (N_1861,N_1857,N_1846);
or U1862 (N_1862,N_1824,N_1819);
nand U1863 (N_1863,N_1812,N_1808);
and U1864 (N_1864,N_1835,N_1833);
nor U1865 (N_1865,N_1806,N_1845);
nand U1866 (N_1866,N_1814,N_1829);
nor U1867 (N_1867,N_1815,N_1848);
and U1868 (N_1868,N_1800,N_1804);
nand U1869 (N_1869,N_1810,N_1856);
or U1870 (N_1870,N_1831,N_1817);
or U1871 (N_1871,N_1837,N_1802);
and U1872 (N_1872,N_1811,N_1832);
nand U1873 (N_1873,N_1826,N_1841);
nand U1874 (N_1874,N_1840,N_1809);
nor U1875 (N_1875,N_1805,N_1813);
and U1876 (N_1876,N_1842,N_1820);
and U1877 (N_1877,N_1854,N_1839);
and U1878 (N_1878,N_1822,N_1852);
nor U1879 (N_1879,N_1847,N_1836);
and U1880 (N_1880,N_1801,N_1858);
nand U1881 (N_1881,N_1830,N_1850);
or U1882 (N_1882,N_1853,N_1816);
nor U1883 (N_1883,N_1844,N_1855);
or U1884 (N_1884,N_1859,N_1838);
nand U1885 (N_1885,N_1807,N_1821);
and U1886 (N_1886,N_1827,N_1828);
or U1887 (N_1887,N_1818,N_1825);
and U1888 (N_1888,N_1803,N_1843);
and U1889 (N_1889,N_1849,N_1834);
nand U1890 (N_1890,N_1848,N_1844);
nor U1891 (N_1891,N_1836,N_1845);
and U1892 (N_1892,N_1841,N_1844);
nor U1893 (N_1893,N_1843,N_1800);
and U1894 (N_1894,N_1807,N_1844);
or U1895 (N_1895,N_1809,N_1822);
xnor U1896 (N_1896,N_1838,N_1819);
and U1897 (N_1897,N_1843,N_1812);
or U1898 (N_1898,N_1837,N_1813);
nand U1899 (N_1899,N_1833,N_1821);
nor U1900 (N_1900,N_1858,N_1834);
or U1901 (N_1901,N_1841,N_1823);
or U1902 (N_1902,N_1823,N_1858);
or U1903 (N_1903,N_1806,N_1817);
and U1904 (N_1904,N_1833,N_1856);
nand U1905 (N_1905,N_1856,N_1800);
and U1906 (N_1906,N_1818,N_1833);
or U1907 (N_1907,N_1839,N_1825);
nand U1908 (N_1908,N_1816,N_1857);
nand U1909 (N_1909,N_1831,N_1852);
nand U1910 (N_1910,N_1825,N_1824);
and U1911 (N_1911,N_1821,N_1801);
nor U1912 (N_1912,N_1857,N_1820);
nand U1913 (N_1913,N_1857,N_1852);
or U1914 (N_1914,N_1842,N_1806);
and U1915 (N_1915,N_1826,N_1814);
and U1916 (N_1916,N_1808,N_1814);
or U1917 (N_1917,N_1836,N_1812);
and U1918 (N_1918,N_1834,N_1812);
and U1919 (N_1919,N_1806,N_1850);
or U1920 (N_1920,N_1911,N_1891);
nand U1921 (N_1921,N_1904,N_1917);
or U1922 (N_1922,N_1909,N_1885);
nor U1923 (N_1923,N_1899,N_1892);
and U1924 (N_1924,N_1878,N_1915);
and U1925 (N_1925,N_1865,N_1919);
nor U1926 (N_1926,N_1887,N_1903);
nor U1927 (N_1927,N_1861,N_1916);
or U1928 (N_1928,N_1918,N_1876);
and U1929 (N_1929,N_1862,N_1912);
or U1930 (N_1930,N_1890,N_1872);
and U1931 (N_1931,N_1863,N_1893);
and U1932 (N_1932,N_1860,N_1902);
or U1933 (N_1933,N_1873,N_1906);
and U1934 (N_1934,N_1888,N_1868);
nor U1935 (N_1935,N_1883,N_1898);
nor U1936 (N_1936,N_1870,N_1871);
nand U1937 (N_1937,N_1880,N_1894);
and U1938 (N_1938,N_1907,N_1866);
or U1939 (N_1939,N_1908,N_1895);
nor U1940 (N_1940,N_1910,N_1869);
and U1941 (N_1941,N_1881,N_1884);
or U1942 (N_1942,N_1896,N_1864);
and U1943 (N_1943,N_1886,N_1897);
nor U1944 (N_1944,N_1867,N_1879);
nor U1945 (N_1945,N_1882,N_1905);
or U1946 (N_1946,N_1875,N_1889);
and U1947 (N_1947,N_1913,N_1877);
and U1948 (N_1948,N_1901,N_1874);
nor U1949 (N_1949,N_1914,N_1900);
and U1950 (N_1950,N_1866,N_1861);
nand U1951 (N_1951,N_1891,N_1896);
nor U1952 (N_1952,N_1916,N_1881);
and U1953 (N_1953,N_1909,N_1898);
nor U1954 (N_1954,N_1866,N_1895);
nand U1955 (N_1955,N_1869,N_1871);
or U1956 (N_1956,N_1886,N_1893);
and U1957 (N_1957,N_1916,N_1873);
and U1958 (N_1958,N_1897,N_1863);
nand U1959 (N_1959,N_1875,N_1873);
or U1960 (N_1960,N_1878,N_1894);
or U1961 (N_1961,N_1897,N_1875);
or U1962 (N_1962,N_1912,N_1913);
nand U1963 (N_1963,N_1919,N_1897);
nor U1964 (N_1964,N_1872,N_1919);
nand U1965 (N_1965,N_1870,N_1895);
or U1966 (N_1966,N_1873,N_1868);
nand U1967 (N_1967,N_1897,N_1896);
and U1968 (N_1968,N_1893,N_1915);
and U1969 (N_1969,N_1883,N_1903);
nand U1970 (N_1970,N_1880,N_1862);
and U1971 (N_1971,N_1888,N_1875);
nor U1972 (N_1972,N_1861,N_1874);
xnor U1973 (N_1973,N_1862,N_1878);
nor U1974 (N_1974,N_1892,N_1876);
nor U1975 (N_1975,N_1880,N_1915);
nand U1976 (N_1976,N_1864,N_1899);
or U1977 (N_1977,N_1910,N_1876);
nand U1978 (N_1978,N_1870,N_1878);
and U1979 (N_1979,N_1886,N_1867);
or U1980 (N_1980,N_1972,N_1941);
nor U1981 (N_1981,N_1942,N_1934);
nor U1982 (N_1982,N_1926,N_1933);
nand U1983 (N_1983,N_1944,N_1959);
nor U1984 (N_1984,N_1940,N_1955);
nand U1985 (N_1985,N_1931,N_1976);
nor U1986 (N_1986,N_1960,N_1954);
and U1987 (N_1987,N_1961,N_1943);
nor U1988 (N_1988,N_1964,N_1922);
or U1989 (N_1989,N_1974,N_1973);
nand U1990 (N_1990,N_1945,N_1953);
nand U1991 (N_1991,N_1920,N_1949);
and U1992 (N_1992,N_1929,N_1930);
or U1993 (N_1993,N_1963,N_1932);
or U1994 (N_1994,N_1946,N_1966);
nand U1995 (N_1995,N_1969,N_1939);
or U1996 (N_1996,N_1979,N_1938);
and U1997 (N_1997,N_1936,N_1928);
nand U1998 (N_1998,N_1975,N_1924);
and U1999 (N_1999,N_1956,N_1923);
and U2000 (N_2000,N_1971,N_1958);
nand U2001 (N_2001,N_1947,N_1951);
and U2002 (N_2002,N_1952,N_1962);
or U2003 (N_2003,N_1935,N_1965);
or U2004 (N_2004,N_1921,N_1978);
nand U2005 (N_2005,N_1937,N_1967);
nor U2006 (N_2006,N_1925,N_1950);
nor U2007 (N_2007,N_1970,N_1968);
nor U2008 (N_2008,N_1977,N_1957);
and U2009 (N_2009,N_1948,N_1927);
nor U2010 (N_2010,N_1926,N_1962);
and U2011 (N_2011,N_1976,N_1962);
nand U2012 (N_2012,N_1969,N_1973);
or U2013 (N_2013,N_1920,N_1957);
and U2014 (N_2014,N_1971,N_1933);
nand U2015 (N_2015,N_1969,N_1937);
nand U2016 (N_2016,N_1967,N_1949);
nand U2017 (N_2017,N_1961,N_1920);
nand U2018 (N_2018,N_1978,N_1975);
and U2019 (N_2019,N_1945,N_1933);
or U2020 (N_2020,N_1934,N_1972);
and U2021 (N_2021,N_1941,N_1971);
nand U2022 (N_2022,N_1946,N_1959);
nand U2023 (N_2023,N_1928,N_1938);
nor U2024 (N_2024,N_1961,N_1928);
nand U2025 (N_2025,N_1949,N_1923);
nand U2026 (N_2026,N_1926,N_1936);
nand U2027 (N_2027,N_1933,N_1960);
and U2028 (N_2028,N_1926,N_1960);
nand U2029 (N_2029,N_1974,N_1947);
and U2030 (N_2030,N_1956,N_1960);
or U2031 (N_2031,N_1970,N_1929);
nand U2032 (N_2032,N_1958,N_1965);
nor U2033 (N_2033,N_1976,N_1934);
and U2034 (N_2034,N_1976,N_1928);
nand U2035 (N_2035,N_1972,N_1975);
and U2036 (N_2036,N_1927,N_1969);
or U2037 (N_2037,N_1942,N_1923);
or U2038 (N_2038,N_1922,N_1958);
or U2039 (N_2039,N_1966,N_1963);
nand U2040 (N_2040,N_2023,N_2029);
and U2041 (N_2041,N_2035,N_2037);
or U2042 (N_2042,N_2015,N_2039);
and U2043 (N_2043,N_2011,N_2024);
or U2044 (N_2044,N_2014,N_2038);
or U2045 (N_2045,N_2034,N_2016);
and U2046 (N_2046,N_2012,N_2020);
nand U2047 (N_2047,N_1987,N_2003);
nand U2048 (N_2048,N_1990,N_1982);
nor U2049 (N_2049,N_2028,N_1993);
or U2050 (N_2050,N_1995,N_2006);
nand U2051 (N_2051,N_2008,N_2021);
and U2052 (N_2052,N_2031,N_1981);
nand U2053 (N_2053,N_1980,N_1998);
nor U2054 (N_2054,N_2005,N_2018);
or U2055 (N_2055,N_2017,N_1996);
or U2056 (N_2056,N_1997,N_2000);
or U2057 (N_2057,N_2033,N_2027);
nor U2058 (N_2058,N_2022,N_2019);
nor U2059 (N_2059,N_1988,N_1985);
nor U2060 (N_2060,N_1986,N_1983);
and U2061 (N_2061,N_2001,N_2013);
nand U2062 (N_2062,N_2032,N_2007);
and U2063 (N_2063,N_2009,N_1992);
nor U2064 (N_2064,N_1984,N_1989);
and U2065 (N_2065,N_2025,N_1999);
nor U2066 (N_2066,N_1994,N_2036);
and U2067 (N_2067,N_2030,N_2004);
nor U2068 (N_2068,N_2002,N_2026);
nor U2069 (N_2069,N_2010,N_1991);
nor U2070 (N_2070,N_2039,N_1991);
or U2071 (N_2071,N_1987,N_2008);
nor U2072 (N_2072,N_2016,N_2018);
xor U2073 (N_2073,N_2034,N_1992);
and U2074 (N_2074,N_2035,N_1996);
or U2075 (N_2075,N_1988,N_2017);
nor U2076 (N_2076,N_1988,N_2038);
nor U2077 (N_2077,N_2009,N_1988);
nand U2078 (N_2078,N_1987,N_2018);
nor U2079 (N_2079,N_2019,N_2005);
nand U2080 (N_2080,N_1980,N_2016);
nand U2081 (N_2081,N_2032,N_2024);
or U2082 (N_2082,N_1996,N_2009);
nand U2083 (N_2083,N_2030,N_2005);
nor U2084 (N_2084,N_2033,N_2031);
nor U2085 (N_2085,N_2017,N_2012);
nor U2086 (N_2086,N_1995,N_2025);
or U2087 (N_2087,N_2009,N_2036);
nand U2088 (N_2088,N_2035,N_2008);
and U2089 (N_2089,N_2027,N_1989);
and U2090 (N_2090,N_2019,N_1983);
nor U2091 (N_2091,N_2034,N_2032);
or U2092 (N_2092,N_1997,N_2009);
nor U2093 (N_2093,N_2010,N_2002);
nand U2094 (N_2094,N_2020,N_2008);
and U2095 (N_2095,N_1994,N_2000);
and U2096 (N_2096,N_2022,N_2026);
and U2097 (N_2097,N_1995,N_2013);
xor U2098 (N_2098,N_2027,N_2014);
or U2099 (N_2099,N_2031,N_2002);
or U2100 (N_2100,N_2087,N_2096);
nor U2101 (N_2101,N_2066,N_2081);
or U2102 (N_2102,N_2092,N_2048);
nand U2103 (N_2103,N_2064,N_2094);
or U2104 (N_2104,N_2083,N_2054);
nor U2105 (N_2105,N_2044,N_2070);
or U2106 (N_2106,N_2065,N_2056);
and U2107 (N_2107,N_2057,N_2041);
nor U2108 (N_2108,N_2052,N_2047);
or U2109 (N_2109,N_2071,N_2062);
nor U2110 (N_2110,N_2042,N_2063);
nor U2111 (N_2111,N_2088,N_2055);
nand U2112 (N_2112,N_2099,N_2082);
or U2113 (N_2113,N_2095,N_2045);
nand U2114 (N_2114,N_2080,N_2076);
nor U2115 (N_2115,N_2077,N_2046);
or U2116 (N_2116,N_2050,N_2075);
nor U2117 (N_2117,N_2051,N_2043);
and U2118 (N_2118,N_2084,N_2097);
or U2119 (N_2119,N_2067,N_2098);
and U2120 (N_2120,N_2040,N_2085);
nand U2121 (N_2121,N_2069,N_2078);
and U2122 (N_2122,N_2058,N_2049);
nand U2123 (N_2123,N_2079,N_2073);
and U2124 (N_2124,N_2068,N_2059);
or U2125 (N_2125,N_2053,N_2060);
nor U2126 (N_2126,N_2089,N_2091);
and U2127 (N_2127,N_2093,N_2086);
and U2128 (N_2128,N_2072,N_2061);
or U2129 (N_2129,N_2074,N_2090);
nor U2130 (N_2130,N_2088,N_2063);
or U2131 (N_2131,N_2049,N_2054);
nor U2132 (N_2132,N_2057,N_2048);
and U2133 (N_2133,N_2041,N_2067);
nand U2134 (N_2134,N_2089,N_2066);
and U2135 (N_2135,N_2051,N_2077);
or U2136 (N_2136,N_2096,N_2043);
and U2137 (N_2137,N_2095,N_2073);
or U2138 (N_2138,N_2082,N_2070);
nor U2139 (N_2139,N_2052,N_2073);
and U2140 (N_2140,N_2062,N_2045);
and U2141 (N_2141,N_2076,N_2048);
or U2142 (N_2142,N_2094,N_2062);
nor U2143 (N_2143,N_2073,N_2086);
or U2144 (N_2144,N_2044,N_2091);
nor U2145 (N_2145,N_2044,N_2076);
and U2146 (N_2146,N_2074,N_2081);
nand U2147 (N_2147,N_2078,N_2066);
nor U2148 (N_2148,N_2045,N_2063);
or U2149 (N_2149,N_2061,N_2049);
nor U2150 (N_2150,N_2067,N_2050);
nor U2151 (N_2151,N_2050,N_2093);
or U2152 (N_2152,N_2097,N_2069);
nand U2153 (N_2153,N_2086,N_2041);
nand U2154 (N_2154,N_2058,N_2075);
or U2155 (N_2155,N_2041,N_2079);
nor U2156 (N_2156,N_2046,N_2085);
nand U2157 (N_2157,N_2082,N_2049);
nor U2158 (N_2158,N_2063,N_2079);
nand U2159 (N_2159,N_2044,N_2065);
nand U2160 (N_2160,N_2145,N_2141);
and U2161 (N_2161,N_2148,N_2111);
and U2162 (N_2162,N_2123,N_2117);
nand U2163 (N_2163,N_2112,N_2118);
and U2164 (N_2164,N_2104,N_2122);
nand U2165 (N_2165,N_2130,N_2106);
and U2166 (N_2166,N_2153,N_2100);
nor U2167 (N_2167,N_2159,N_2132);
and U2168 (N_2168,N_2138,N_2124);
nor U2169 (N_2169,N_2146,N_2108);
nor U2170 (N_2170,N_2102,N_2155);
or U2171 (N_2171,N_2147,N_2121);
nor U2172 (N_2172,N_2140,N_2115);
nor U2173 (N_2173,N_2137,N_2149);
nand U2174 (N_2174,N_2142,N_2143);
or U2175 (N_2175,N_2151,N_2128);
and U2176 (N_2176,N_2127,N_2116);
or U2177 (N_2177,N_2125,N_2119);
and U2178 (N_2178,N_2157,N_2150);
nor U2179 (N_2179,N_2152,N_2154);
or U2180 (N_2180,N_2134,N_2144);
nand U2181 (N_2181,N_2135,N_2101);
nand U2182 (N_2182,N_2113,N_2131);
nor U2183 (N_2183,N_2105,N_2133);
nor U2184 (N_2184,N_2103,N_2126);
or U2185 (N_2185,N_2107,N_2120);
and U2186 (N_2186,N_2110,N_2114);
and U2187 (N_2187,N_2158,N_2136);
nand U2188 (N_2188,N_2156,N_2139);
nor U2189 (N_2189,N_2129,N_2109);
and U2190 (N_2190,N_2104,N_2121);
and U2191 (N_2191,N_2139,N_2126);
or U2192 (N_2192,N_2122,N_2143);
and U2193 (N_2193,N_2123,N_2155);
nor U2194 (N_2194,N_2129,N_2104);
or U2195 (N_2195,N_2152,N_2139);
and U2196 (N_2196,N_2156,N_2111);
or U2197 (N_2197,N_2113,N_2133);
or U2198 (N_2198,N_2152,N_2123);
nor U2199 (N_2199,N_2116,N_2135);
or U2200 (N_2200,N_2131,N_2108);
or U2201 (N_2201,N_2118,N_2123);
nor U2202 (N_2202,N_2127,N_2158);
or U2203 (N_2203,N_2127,N_2149);
and U2204 (N_2204,N_2123,N_2119);
nor U2205 (N_2205,N_2125,N_2128);
nor U2206 (N_2206,N_2155,N_2151);
nor U2207 (N_2207,N_2113,N_2129);
nor U2208 (N_2208,N_2147,N_2124);
or U2209 (N_2209,N_2151,N_2120);
nor U2210 (N_2210,N_2121,N_2131);
nor U2211 (N_2211,N_2142,N_2158);
xnor U2212 (N_2212,N_2136,N_2152);
nor U2213 (N_2213,N_2100,N_2128);
xnor U2214 (N_2214,N_2100,N_2116);
nor U2215 (N_2215,N_2149,N_2154);
or U2216 (N_2216,N_2108,N_2122);
and U2217 (N_2217,N_2109,N_2156);
or U2218 (N_2218,N_2158,N_2152);
and U2219 (N_2219,N_2134,N_2121);
nand U2220 (N_2220,N_2209,N_2168);
nor U2221 (N_2221,N_2198,N_2218);
and U2222 (N_2222,N_2214,N_2212);
nand U2223 (N_2223,N_2169,N_2208);
or U2224 (N_2224,N_2176,N_2206);
and U2225 (N_2225,N_2191,N_2184);
and U2226 (N_2226,N_2193,N_2183);
nor U2227 (N_2227,N_2170,N_2172);
nand U2228 (N_2228,N_2160,N_2217);
or U2229 (N_2229,N_2205,N_2207);
or U2230 (N_2230,N_2175,N_2216);
and U2231 (N_2231,N_2203,N_2204);
or U2232 (N_2232,N_2200,N_2181);
and U2233 (N_2233,N_2196,N_2190);
nor U2234 (N_2234,N_2189,N_2177);
nand U2235 (N_2235,N_2201,N_2213);
nand U2236 (N_2236,N_2202,N_2173);
nor U2237 (N_2237,N_2161,N_2174);
nand U2238 (N_2238,N_2171,N_2210);
and U2239 (N_2239,N_2163,N_2180);
nor U2240 (N_2240,N_2166,N_2188);
or U2241 (N_2241,N_2182,N_2185);
or U2242 (N_2242,N_2195,N_2192);
or U2243 (N_2243,N_2187,N_2219);
nand U2244 (N_2244,N_2162,N_2211);
or U2245 (N_2245,N_2186,N_2165);
nand U2246 (N_2246,N_2164,N_2179);
nand U2247 (N_2247,N_2178,N_2194);
nor U2248 (N_2248,N_2197,N_2167);
nand U2249 (N_2249,N_2215,N_2199);
or U2250 (N_2250,N_2174,N_2200);
nand U2251 (N_2251,N_2211,N_2179);
or U2252 (N_2252,N_2189,N_2166);
and U2253 (N_2253,N_2197,N_2208);
nor U2254 (N_2254,N_2165,N_2198);
and U2255 (N_2255,N_2204,N_2161);
nand U2256 (N_2256,N_2194,N_2208);
nor U2257 (N_2257,N_2190,N_2184);
nor U2258 (N_2258,N_2175,N_2170);
or U2259 (N_2259,N_2186,N_2176);
nor U2260 (N_2260,N_2219,N_2214);
nand U2261 (N_2261,N_2213,N_2170);
nor U2262 (N_2262,N_2170,N_2179);
nor U2263 (N_2263,N_2219,N_2162);
nand U2264 (N_2264,N_2213,N_2191);
nand U2265 (N_2265,N_2199,N_2217);
or U2266 (N_2266,N_2186,N_2215);
nand U2267 (N_2267,N_2176,N_2205);
or U2268 (N_2268,N_2191,N_2189);
nand U2269 (N_2269,N_2182,N_2166);
or U2270 (N_2270,N_2184,N_2175);
nor U2271 (N_2271,N_2187,N_2202);
nand U2272 (N_2272,N_2204,N_2178);
nand U2273 (N_2273,N_2198,N_2193);
nor U2274 (N_2274,N_2170,N_2199);
nor U2275 (N_2275,N_2180,N_2186);
nor U2276 (N_2276,N_2184,N_2168);
or U2277 (N_2277,N_2172,N_2183);
xnor U2278 (N_2278,N_2216,N_2186);
nand U2279 (N_2279,N_2202,N_2207);
nor U2280 (N_2280,N_2259,N_2247);
nand U2281 (N_2281,N_2278,N_2252);
and U2282 (N_2282,N_2272,N_2239);
nor U2283 (N_2283,N_2228,N_2279);
nor U2284 (N_2284,N_2270,N_2224);
and U2285 (N_2285,N_2260,N_2266);
xnor U2286 (N_2286,N_2220,N_2276);
and U2287 (N_2287,N_2248,N_2223);
or U2288 (N_2288,N_2232,N_2243);
or U2289 (N_2289,N_2256,N_2251);
and U2290 (N_2290,N_2262,N_2246);
nor U2291 (N_2291,N_2277,N_2275);
nor U2292 (N_2292,N_2237,N_2273);
nor U2293 (N_2293,N_2240,N_2254);
and U2294 (N_2294,N_2222,N_2235);
nand U2295 (N_2295,N_2221,N_2264);
nand U2296 (N_2296,N_2227,N_2241);
nand U2297 (N_2297,N_2238,N_2233);
and U2298 (N_2298,N_2271,N_2236);
nand U2299 (N_2299,N_2249,N_2265);
or U2300 (N_2300,N_2231,N_2268);
or U2301 (N_2301,N_2261,N_2269);
or U2302 (N_2302,N_2257,N_2250);
nand U2303 (N_2303,N_2244,N_2245);
nand U2304 (N_2304,N_2230,N_2225);
and U2305 (N_2305,N_2234,N_2258);
and U2306 (N_2306,N_2255,N_2226);
nand U2307 (N_2307,N_2263,N_2229);
nand U2308 (N_2308,N_2253,N_2274);
nand U2309 (N_2309,N_2242,N_2267);
or U2310 (N_2310,N_2230,N_2253);
nand U2311 (N_2311,N_2242,N_2247);
nand U2312 (N_2312,N_2238,N_2244);
and U2313 (N_2313,N_2238,N_2243);
or U2314 (N_2314,N_2244,N_2248);
or U2315 (N_2315,N_2226,N_2259);
nor U2316 (N_2316,N_2256,N_2224);
and U2317 (N_2317,N_2273,N_2227);
nor U2318 (N_2318,N_2276,N_2227);
or U2319 (N_2319,N_2257,N_2236);
or U2320 (N_2320,N_2271,N_2226);
and U2321 (N_2321,N_2239,N_2238);
nand U2322 (N_2322,N_2265,N_2241);
or U2323 (N_2323,N_2225,N_2257);
nor U2324 (N_2324,N_2254,N_2246);
nand U2325 (N_2325,N_2226,N_2265);
nor U2326 (N_2326,N_2269,N_2257);
nor U2327 (N_2327,N_2226,N_2253);
and U2328 (N_2328,N_2276,N_2225);
or U2329 (N_2329,N_2276,N_2259);
or U2330 (N_2330,N_2233,N_2230);
or U2331 (N_2331,N_2232,N_2227);
or U2332 (N_2332,N_2266,N_2273);
and U2333 (N_2333,N_2268,N_2243);
nor U2334 (N_2334,N_2275,N_2228);
and U2335 (N_2335,N_2264,N_2244);
nand U2336 (N_2336,N_2241,N_2243);
nand U2337 (N_2337,N_2242,N_2268);
or U2338 (N_2338,N_2268,N_2250);
and U2339 (N_2339,N_2237,N_2231);
or U2340 (N_2340,N_2286,N_2309);
or U2341 (N_2341,N_2288,N_2302);
nand U2342 (N_2342,N_2335,N_2326);
nor U2343 (N_2343,N_2316,N_2322);
nor U2344 (N_2344,N_2299,N_2285);
nor U2345 (N_2345,N_2329,N_2311);
nor U2346 (N_2346,N_2305,N_2304);
or U2347 (N_2347,N_2331,N_2297);
or U2348 (N_2348,N_2318,N_2296);
nand U2349 (N_2349,N_2289,N_2303);
xor U2350 (N_2350,N_2310,N_2314);
nor U2351 (N_2351,N_2283,N_2320);
or U2352 (N_2352,N_2328,N_2338);
nor U2353 (N_2353,N_2295,N_2294);
nor U2354 (N_2354,N_2319,N_2301);
or U2355 (N_2355,N_2323,N_2315);
nand U2356 (N_2356,N_2290,N_2337);
nand U2357 (N_2357,N_2308,N_2321);
and U2358 (N_2358,N_2287,N_2339);
or U2359 (N_2359,N_2332,N_2281);
nand U2360 (N_2360,N_2300,N_2334);
and U2361 (N_2361,N_2336,N_2291);
or U2362 (N_2362,N_2313,N_2312);
and U2363 (N_2363,N_2317,N_2324);
nand U2364 (N_2364,N_2306,N_2282);
and U2365 (N_2365,N_2330,N_2325);
nand U2366 (N_2366,N_2333,N_2327);
and U2367 (N_2367,N_2292,N_2280);
or U2368 (N_2368,N_2293,N_2307);
or U2369 (N_2369,N_2284,N_2298);
or U2370 (N_2370,N_2316,N_2284);
and U2371 (N_2371,N_2320,N_2305);
and U2372 (N_2372,N_2335,N_2325);
and U2373 (N_2373,N_2303,N_2320);
and U2374 (N_2374,N_2332,N_2323);
nor U2375 (N_2375,N_2310,N_2312);
or U2376 (N_2376,N_2304,N_2318);
nand U2377 (N_2377,N_2281,N_2296);
nand U2378 (N_2378,N_2300,N_2321);
and U2379 (N_2379,N_2318,N_2333);
or U2380 (N_2380,N_2290,N_2333);
nand U2381 (N_2381,N_2312,N_2287);
nor U2382 (N_2382,N_2296,N_2333);
and U2383 (N_2383,N_2282,N_2320);
nand U2384 (N_2384,N_2299,N_2288);
and U2385 (N_2385,N_2313,N_2290);
nand U2386 (N_2386,N_2324,N_2288);
and U2387 (N_2387,N_2292,N_2335);
nand U2388 (N_2388,N_2331,N_2318);
nor U2389 (N_2389,N_2304,N_2301);
and U2390 (N_2390,N_2310,N_2332);
nand U2391 (N_2391,N_2281,N_2327);
and U2392 (N_2392,N_2314,N_2284);
or U2393 (N_2393,N_2334,N_2326);
or U2394 (N_2394,N_2304,N_2288);
and U2395 (N_2395,N_2302,N_2306);
nor U2396 (N_2396,N_2299,N_2301);
and U2397 (N_2397,N_2309,N_2307);
nor U2398 (N_2398,N_2325,N_2306);
nor U2399 (N_2399,N_2312,N_2293);
and U2400 (N_2400,N_2393,N_2374);
or U2401 (N_2401,N_2352,N_2367);
or U2402 (N_2402,N_2397,N_2379);
nor U2403 (N_2403,N_2376,N_2396);
nand U2404 (N_2404,N_2350,N_2346);
and U2405 (N_2405,N_2364,N_2343);
or U2406 (N_2406,N_2357,N_2390);
or U2407 (N_2407,N_2377,N_2340);
or U2408 (N_2408,N_2392,N_2359);
or U2409 (N_2409,N_2349,N_2387);
nand U2410 (N_2410,N_2371,N_2354);
and U2411 (N_2411,N_2368,N_2382);
nand U2412 (N_2412,N_2385,N_2394);
or U2413 (N_2413,N_2360,N_2381);
nor U2414 (N_2414,N_2361,N_2345);
nor U2415 (N_2415,N_2348,N_2362);
or U2416 (N_2416,N_2369,N_2344);
or U2417 (N_2417,N_2358,N_2355);
nor U2418 (N_2418,N_2380,N_2399);
nor U2419 (N_2419,N_2363,N_2388);
or U2420 (N_2420,N_2341,N_2391);
or U2421 (N_2421,N_2373,N_2386);
nor U2422 (N_2422,N_2383,N_2342);
or U2423 (N_2423,N_2378,N_2398);
nand U2424 (N_2424,N_2375,N_2384);
and U2425 (N_2425,N_2389,N_2353);
nor U2426 (N_2426,N_2356,N_2370);
or U2427 (N_2427,N_2366,N_2351);
nand U2428 (N_2428,N_2347,N_2372);
and U2429 (N_2429,N_2395,N_2365);
or U2430 (N_2430,N_2387,N_2380);
nand U2431 (N_2431,N_2353,N_2340);
and U2432 (N_2432,N_2356,N_2346);
nand U2433 (N_2433,N_2391,N_2343);
or U2434 (N_2434,N_2353,N_2342);
nand U2435 (N_2435,N_2392,N_2366);
nand U2436 (N_2436,N_2397,N_2363);
or U2437 (N_2437,N_2350,N_2369);
or U2438 (N_2438,N_2376,N_2345);
nor U2439 (N_2439,N_2344,N_2365);
nor U2440 (N_2440,N_2397,N_2366);
or U2441 (N_2441,N_2366,N_2389);
or U2442 (N_2442,N_2372,N_2363);
and U2443 (N_2443,N_2343,N_2369);
nand U2444 (N_2444,N_2349,N_2345);
nor U2445 (N_2445,N_2376,N_2392);
and U2446 (N_2446,N_2366,N_2399);
nor U2447 (N_2447,N_2360,N_2399);
nand U2448 (N_2448,N_2366,N_2374);
nor U2449 (N_2449,N_2361,N_2343);
and U2450 (N_2450,N_2392,N_2399);
nor U2451 (N_2451,N_2369,N_2395);
nand U2452 (N_2452,N_2390,N_2399);
xnor U2453 (N_2453,N_2346,N_2385);
or U2454 (N_2454,N_2386,N_2366);
nor U2455 (N_2455,N_2384,N_2386);
and U2456 (N_2456,N_2342,N_2366);
nor U2457 (N_2457,N_2347,N_2342);
and U2458 (N_2458,N_2383,N_2341);
nor U2459 (N_2459,N_2360,N_2356);
and U2460 (N_2460,N_2442,N_2437);
and U2461 (N_2461,N_2406,N_2403);
and U2462 (N_2462,N_2451,N_2414);
and U2463 (N_2463,N_2445,N_2401);
nor U2464 (N_2464,N_2447,N_2400);
and U2465 (N_2465,N_2419,N_2422);
or U2466 (N_2466,N_2420,N_2450);
or U2467 (N_2467,N_2415,N_2431);
and U2468 (N_2468,N_2423,N_2424);
nand U2469 (N_2469,N_2446,N_2449);
and U2470 (N_2470,N_2421,N_2458);
and U2471 (N_2471,N_2418,N_2444);
nor U2472 (N_2472,N_2411,N_2454);
or U2473 (N_2473,N_2452,N_2435);
nor U2474 (N_2474,N_2409,N_2408);
nor U2475 (N_2475,N_2426,N_2436);
nor U2476 (N_2476,N_2434,N_2402);
nor U2477 (N_2477,N_2432,N_2425);
or U2478 (N_2478,N_2417,N_2429);
nand U2479 (N_2479,N_2448,N_2456);
or U2480 (N_2480,N_2413,N_2427);
nor U2481 (N_2481,N_2428,N_2416);
or U2482 (N_2482,N_2453,N_2443);
or U2483 (N_2483,N_2404,N_2412);
or U2484 (N_2484,N_2433,N_2407);
nand U2485 (N_2485,N_2441,N_2439);
nand U2486 (N_2486,N_2410,N_2459);
and U2487 (N_2487,N_2455,N_2440);
or U2488 (N_2488,N_2438,N_2405);
nor U2489 (N_2489,N_2430,N_2457);
nand U2490 (N_2490,N_2401,N_2443);
nor U2491 (N_2491,N_2430,N_2423);
xnor U2492 (N_2492,N_2452,N_2440);
or U2493 (N_2493,N_2458,N_2404);
and U2494 (N_2494,N_2442,N_2415);
nand U2495 (N_2495,N_2422,N_2401);
and U2496 (N_2496,N_2423,N_2410);
nor U2497 (N_2497,N_2422,N_2435);
or U2498 (N_2498,N_2432,N_2421);
nand U2499 (N_2499,N_2411,N_2436);
xor U2500 (N_2500,N_2444,N_2425);
or U2501 (N_2501,N_2400,N_2416);
nor U2502 (N_2502,N_2436,N_2424);
or U2503 (N_2503,N_2423,N_2450);
and U2504 (N_2504,N_2443,N_2442);
and U2505 (N_2505,N_2426,N_2408);
or U2506 (N_2506,N_2431,N_2409);
or U2507 (N_2507,N_2447,N_2431);
or U2508 (N_2508,N_2436,N_2422);
or U2509 (N_2509,N_2456,N_2411);
and U2510 (N_2510,N_2423,N_2418);
xnor U2511 (N_2511,N_2448,N_2405);
or U2512 (N_2512,N_2426,N_2440);
xor U2513 (N_2513,N_2435,N_2419);
nor U2514 (N_2514,N_2455,N_2447);
and U2515 (N_2515,N_2404,N_2448);
and U2516 (N_2516,N_2424,N_2440);
or U2517 (N_2517,N_2429,N_2448);
nand U2518 (N_2518,N_2446,N_2430);
or U2519 (N_2519,N_2418,N_2438);
nand U2520 (N_2520,N_2488,N_2515);
and U2521 (N_2521,N_2518,N_2489);
or U2522 (N_2522,N_2514,N_2503);
or U2523 (N_2523,N_2493,N_2476);
nand U2524 (N_2524,N_2509,N_2519);
or U2525 (N_2525,N_2464,N_2516);
nand U2526 (N_2526,N_2487,N_2490);
nand U2527 (N_2527,N_2485,N_2478);
or U2528 (N_2528,N_2468,N_2504);
and U2529 (N_2529,N_2505,N_2508);
or U2530 (N_2530,N_2486,N_2492);
or U2531 (N_2531,N_2495,N_2460);
and U2532 (N_2532,N_2465,N_2501);
nand U2533 (N_2533,N_2463,N_2491);
or U2534 (N_2534,N_2473,N_2466);
nand U2535 (N_2535,N_2512,N_2499);
nor U2536 (N_2536,N_2513,N_2517);
and U2537 (N_2537,N_2496,N_2474);
nand U2538 (N_2538,N_2482,N_2470);
nor U2539 (N_2539,N_2469,N_2467);
nor U2540 (N_2540,N_2484,N_2497);
and U2541 (N_2541,N_2506,N_2494);
or U2542 (N_2542,N_2461,N_2507);
nor U2543 (N_2543,N_2500,N_2480);
nand U2544 (N_2544,N_2475,N_2510);
and U2545 (N_2545,N_2477,N_2483);
nand U2546 (N_2546,N_2462,N_2479);
and U2547 (N_2547,N_2471,N_2472);
nand U2548 (N_2548,N_2498,N_2511);
or U2549 (N_2549,N_2481,N_2502);
nand U2550 (N_2550,N_2498,N_2484);
nor U2551 (N_2551,N_2490,N_2513);
or U2552 (N_2552,N_2510,N_2507);
nor U2553 (N_2553,N_2497,N_2506);
or U2554 (N_2554,N_2471,N_2491);
nor U2555 (N_2555,N_2504,N_2503);
or U2556 (N_2556,N_2503,N_2486);
and U2557 (N_2557,N_2469,N_2483);
or U2558 (N_2558,N_2506,N_2460);
nand U2559 (N_2559,N_2480,N_2505);
or U2560 (N_2560,N_2518,N_2492);
nand U2561 (N_2561,N_2482,N_2508);
nand U2562 (N_2562,N_2464,N_2466);
and U2563 (N_2563,N_2513,N_2489);
or U2564 (N_2564,N_2501,N_2495);
or U2565 (N_2565,N_2496,N_2476);
and U2566 (N_2566,N_2511,N_2503);
and U2567 (N_2567,N_2484,N_2505);
and U2568 (N_2568,N_2512,N_2474);
or U2569 (N_2569,N_2477,N_2465);
nand U2570 (N_2570,N_2496,N_2483);
and U2571 (N_2571,N_2462,N_2503);
nand U2572 (N_2572,N_2477,N_2494);
and U2573 (N_2573,N_2497,N_2461);
or U2574 (N_2574,N_2501,N_2467);
nor U2575 (N_2575,N_2480,N_2482);
and U2576 (N_2576,N_2468,N_2510);
nand U2577 (N_2577,N_2516,N_2512);
nor U2578 (N_2578,N_2502,N_2467);
nor U2579 (N_2579,N_2493,N_2470);
nor U2580 (N_2580,N_2534,N_2559);
nor U2581 (N_2581,N_2520,N_2574);
nor U2582 (N_2582,N_2547,N_2555);
nor U2583 (N_2583,N_2532,N_2571);
and U2584 (N_2584,N_2577,N_2546);
nand U2585 (N_2585,N_2550,N_2542);
or U2586 (N_2586,N_2539,N_2524);
and U2587 (N_2587,N_2568,N_2579);
xor U2588 (N_2588,N_2545,N_2557);
or U2589 (N_2589,N_2554,N_2530);
nand U2590 (N_2590,N_2572,N_2535);
and U2591 (N_2591,N_2576,N_2538);
nand U2592 (N_2592,N_2526,N_2558);
and U2593 (N_2593,N_2560,N_2541);
nor U2594 (N_2594,N_2567,N_2561);
nor U2595 (N_2595,N_2531,N_2552);
nand U2596 (N_2596,N_2528,N_2578);
or U2597 (N_2597,N_2564,N_2544);
nor U2598 (N_2598,N_2529,N_2553);
or U2599 (N_2599,N_2523,N_2551);
or U2600 (N_2600,N_2573,N_2522);
and U2601 (N_2601,N_2562,N_2566);
nor U2602 (N_2602,N_2536,N_2543);
and U2603 (N_2603,N_2525,N_2533);
or U2604 (N_2604,N_2548,N_2521);
nor U2605 (N_2605,N_2569,N_2556);
or U2606 (N_2606,N_2537,N_2565);
nor U2607 (N_2607,N_2540,N_2549);
and U2608 (N_2608,N_2575,N_2527);
nand U2609 (N_2609,N_2570,N_2563);
nor U2610 (N_2610,N_2521,N_2571);
or U2611 (N_2611,N_2545,N_2573);
and U2612 (N_2612,N_2554,N_2550);
or U2613 (N_2613,N_2571,N_2551);
and U2614 (N_2614,N_2560,N_2563);
or U2615 (N_2615,N_2548,N_2534);
xor U2616 (N_2616,N_2564,N_2527);
nand U2617 (N_2617,N_2536,N_2538);
nand U2618 (N_2618,N_2550,N_2537);
or U2619 (N_2619,N_2542,N_2537);
nand U2620 (N_2620,N_2574,N_2532);
nand U2621 (N_2621,N_2570,N_2538);
and U2622 (N_2622,N_2521,N_2567);
nand U2623 (N_2623,N_2525,N_2540);
and U2624 (N_2624,N_2568,N_2569);
nand U2625 (N_2625,N_2573,N_2574);
nor U2626 (N_2626,N_2534,N_2531);
nor U2627 (N_2627,N_2574,N_2561);
nor U2628 (N_2628,N_2536,N_2572);
nor U2629 (N_2629,N_2555,N_2567);
nand U2630 (N_2630,N_2526,N_2542);
nor U2631 (N_2631,N_2555,N_2526);
or U2632 (N_2632,N_2579,N_2529);
nand U2633 (N_2633,N_2555,N_2562);
and U2634 (N_2634,N_2541,N_2548);
nor U2635 (N_2635,N_2550,N_2563);
nor U2636 (N_2636,N_2548,N_2573);
or U2637 (N_2637,N_2545,N_2566);
or U2638 (N_2638,N_2563,N_2577);
or U2639 (N_2639,N_2531,N_2551);
or U2640 (N_2640,N_2591,N_2589);
and U2641 (N_2641,N_2632,N_2588);
xor U2642 (N_2642,N_2603,N_2609);
or U2643 (N_2643,N_2631,N_2613);
nor U2644 (N_2644,N_2628,N_2604);
and U2645 (N_2645,N_2621,N_2617);
or U2646 (N_2646,N_2614,N_2595);
nor U2647 (N_2647,N_2618,N_2612);
nand U2648 (N_2648,N_2622,N_2633);
nor U2649 (N_2649,N_2610,N_2615);
and U2650 (N_2650,N_2585,N_2598);
or U2651 (N_2651,N_2616,N_2580);
nand U2652 (N_2652,N_2624,N_2581);
nand U2653 (N_2653,N_2597,N_2601);
nand U2654 (N_2654,N_2600,N_2629);
or U2655 (N_2655,N_2623,N_2625);
nand U2656 (N_2656,N_2626,N_2619);
nor U2657 (N_2657,N_2605,N_2608);
and U2658 (N_2658,N_2583,N_2630);
nand U2659 (N_2659,N_2611,N_2638);
and U2660 (N_2660,N_2635,N_2636);
or U2661 (N_2661,N_2606,N_2607);
nor U2662 (N_2662,N_2586,N_2627);
nand U2663 (N_2663,N_2582,N_2587);
or U2664 (N_2664,N_2634,N_2620);
and U2665 (N_2665,N_2596,N_2599);
or U2666 (N_2666,N_2584,N_2592);
or U2667 (N_2667,N_2637,N_2594);
nand U2668 (N_2668,N_2639,N_2593);
nand U2669 (N_2669,N_2590,N_2602);
nor U2670 (N_2670,N_2603,N_2608);
and U2671 (N_2671,N_2591,N_2629);
nor U2672 (N_2672,N_2588,N_2601);
nand U2673 (N_2673,N_2620,N_2614);
nand U2674 (N_2674,N_2631,N_2606);
or U2675 (N_2675,N_2609,N_2615);
or U2676 (N_2676,N_2607,N_2603);
or U2677 (N_2677,N_2618,N_2606);
or U2678 (N_2678,N_2592,N_2613);
and U2679 (N_2679,N_2595,N_2613);
nor U2680 (N_2680,N_2634,N_2619);
nor U2681 (N_2681,N_2595,N_2628);
or U2682 (N_2682,N_2615,N_2590);
nand U2683 (N_2683,N_2622,N_2632);
or U2684 (N_2684,N_2584,N_2626);
nand U2685 (N_2685,N_2632,N_2630);
or U2686 (N_2686,N_2592,N_2628);
or U2687 (N_2687,N_2596,N_2633);
or U2688 (N_2688,N_2581,N_2633);
xor U2689 (N_2689,N_2600,N_2614);
nor U2690 (N_2690,N_2627,N_2618);
nand U2691 (N_2691,N_2602,N_2612);
nand U2692 (N_2692,N_2586,N_2607);
or U2693 (N_2693,N_2617,N_2635);
or U2694 (N_2694,N_2601,N_2606);
nor U2695 (N_2695,N_2625,N_2611);
and U2696 (N_2696,N_2612,N_2605);
and U2697 (N_2697,N_2592,N_2638);
or U2698 (N_2698,N_2639,N_2626);
and U2699 (N_2699,N_2585,N_2609);
or U2700 (N_2700,N_2657,N_2678);
nor U2701 (N_2701,N_2668,N_2693);
and U2702 (N_2702,N_2677,N_2650);
nand U2703 (N_2703,N_2695,N_2653);
or U2704 (N_2704,N_2660,N_2643);
or U2705 (N_2705,N_2682,N_2674);
xor U2706 (N_2706,N_2648,N_2672);
nor U2707 (N_2707,N_2673,N_2691);
or U2708 (N_2708,N_2664,N_2681);
nand U2709 (N_2709,N_2662,N_2696);
nand U2710 (N_2710,N_2679,N_2641);
nor U2711 (N_2711,N_2652,N_2685);
nand U2712 (N_2712,N_2688,N_2690);
and U2713 (N_2713,N_2684,N_2683);
nor U2714 (N_2714,N_2646,N_2687);
and U2715 (N_2715,N_2692,N_2663);
and U2716 (N_2716,N_2676,N_2697);
nor U2717 (N_2717,N_2671,N_2647);
or U2718 (N_2718,N_2666,N_2659);
nor U2719 (N_2719,N_2644,N_2699);
nor U2720 (N_2720,N_2642,N_2649);
nand U2721 (N_2721,N_2655,N_2680);
or U2722 (N_2722,N_2689,N_2654);
or U2723 (N_2723,N_2640,N_2656);
nor U2724 (N_2724,N_2645,N_2698);
nand U2725 (N_2725,N_2661,N_2651);
and U2726 (N_2726,N_2665,N_2667);
and U2727 (N_2727,N_2686,N_2675);
nor U2728 (N_2728,N_2669,N_2694);
nand U2729 (N_2729,N_2658,N_2670);
nor U2730 (N_2730,N_2689,N_2657);
and U2731 (N_2731,N_2655,N_2683);
nand U2732 (N_2732,N_2682,N_2648);
and U2733 (N_2733,N_2647,N_2645);
or U2734 (N_2734,N_2677,N_2689);
nand U2735 (N_2735,N_2653,N_2666);
or U2736 (N_2736,N_2651,N_2641);
nor U2737 (N_2737,N_2643,N_2687);
nand U2738 (N_2738,N_2662,N_2668);
nand U2739 (N_2739,N_2694,N_2697);
nand U2740 (N_2740,N_2680,N_2690);
or U2741 (N_2741,N_2673,N_2684);
nor U2742 (N_2742,N_2663,N_2681);
nand U2743 (N_2743,N_2691,N_2675);
nor U2744 (N_2744,N_2686,N_2648);
xor U2745 (N_2745,N_2661,N_2692);
xor U2746 (N_2746,N_2651,N_2679);
nand U2747 (N_2747,N_2686,N_2676);
nor U2748 (N_2748,N_2644,N_2681);
and U2749 (N_2749,N_2677,N_2653);
nor U2750 (N_2750,N_2684,N_2693);
nand U2751 (N_2751,N_2664,N_2685);
nand U2752 (N_2752,N_2661,N_2645);
or U2753 (N_2753,N_2666,N_2688);
nor U2754 (N_2754,N_2686,N_2672);
nor U2755 (N_2755,N_2683,N_2644);
nor U2756 (N_2756,N_2674,N_2687);
and U2757 (N_2757,N_2688,N_2654);
nor U2758 (N_2758,N_2653,N_2657);
or U2759 (N_2759,N_2699,N_2645);
or U2760 (N_2760,N_2739,N_2718);
and U2761 (N_2761,N_2758,N_2742);
or U2762 (N_2762,N_2731,N_2755);
or U2763 (N_2763,N_2757,N_2722);
nor U2764 (N_2764,N_2707,N_2708);
nand U2765 (N_2765,N_2712,N_2705);
nor U2766 (N_2766,N_2749,N_2738);
or U2767 (N_2767,N_2743,N_2720);
and U2768 (N_2768,N_2726,N_2741);
or U2769 (N_2769,N_2700,N_2734);
nand U2770 (N_2770,N_2729,N_2746);
nand U2771 (N_2771,N_2719,N_2752);
and U2772 (N_2772,N_2714,N_2710);
and U2773 (N_2773,N_2730,N_2723);
nor U2774 (N_2774,N_2702,N_2754);
or U2775 (N_2775,N_2744,N_2753);
and U2776 (N_2776,N_2751,N_2706);
and U2777 (N_2777,N_2735,N_2732);
and U2778 (N_2778,N_2716,N_2703);
nor U2779 (N_2779,N_2725,N_2715);
and U2780 (N_2780,N_2756,N_2728);
or U2781 (N_2781,N_2759,N_2713);
nor U2782 (N_2782,N_2736,N_2727);
or U2783 (N_2783,N_2724,N_2748);
or U2784 (N_2784,N_2721,N_2740);
nand U2785 (N_2785,N_2733,N_2747);
and U2786 (N_2786,N_2717,N_2711);
or U2787 (N_2787,N_2750,N_2704);
nor U2788 (N_2788,N_2701,N_2737);
or U2789 (N_2789,N_2745,N_2709);
and U2790 (N_2790,N_2714,N_2751);
nand U2791 (N_2791,N_2723,N_2759);
and U2792 (N_2792,N_2718,N_2733);
and U2793 (N_2793,N_2713,N_2709);
nor U2794 (N_2794,N_2702,N_2731);
or U2795 (N_2795,N_2701,N_2750);
and U2796 (N_2796,N_2740,N_2759);
and U2797 (N_2797,N_2756,N_2722);
nand U2798 (N_2798,N_2717,N_2756);
or U2799 (N_2799,N_2707,N_2740);
nor U2800 (N_2800,N_2712,N_2721);
nand U2801 (N_2801,N_2721,N_2731);
nor U2802 (N_2802,N_2701,N_2728);
nor U2803 (N_2803,N_2755,N_2754);
or U2804 (N_2804,N_2757,N_2711);
or U2805 (N_2805,N_2759,N_2753);
and U2806 (N_2806,N_2706,N_2701);
or U2807 (N_2807,N_2724,N_2711);
nor U2808 (N_2808,N_2726,N_2736);
and U2809 (N_2809,N_2759,N_2743);
and U2810 (N_2810,N_2701,N_2722);
nand U2811 (N_2811,N_2708,N_2758);
nand U2812 (N_2812,N_2754,N_2707);
nor U2813 (N_2813,N_2754,N_2725);
nand U2814 (N_2814,N_2737,N_2735);
nand U2815 (N_2815,N_2737,N_2731);
or U2816 (N_2816,N_2705,N_2715);
nand U2817 (N_2817,N_2701,N_2735);
and U2818 (N_2818,N_2716,N_2753);
nor U2819 (N_2819,N_2722,N_2745);
and U2820 (N_2820,N_2800,N_2768);
or U2821 (N_2821,N_2769,N_2792);
nor U2822 (N_2822,N_2808,N_2796);
or U2823 (N_2823,N_2818,N_2794);
and U2824 (N_2824,N_2773,N_2787);
and U2825 (N_2825,N_2781,N_2811);
and U2826 (N_2826,N_2783,N_2778);
or U2827 (N_2827,N_2790,N_2819);
and U2828 (N_2828,N_2804,N_2793);
nor U2829 (N_2829,N_2772,N_2761);
nor U2830 (N_2830,N_2767,N_2766);
or U2831 (N_2831,N_2812,N_2788);
or U2832 (N_2832,N_2791,N_2813);
nor U2833 (N_2833,N_2776,N_2770);
nand U2834 (N_2834,N_2816,N_2763);
or U2835 (N_2835,N_2784,N_2780);
nor U2836 (N_2836,N_2765,N_2801);
nand U2837 (N_2837,N_2785,N_2815);
or U2838 (N_2838,N_2807,N_2797);
nand U2839 (N_2839,N_2809,N_2775);
or U2840 (N_2840,N_2762,N_2814);
nor U2841 (N_2841,N_2802,N_2771);
and U2842 (N_2842,N_2789,N_2774);
nand U2843 (N_2843,N_2777,N_2806);
or U2844 (N_2844,N_2786,N_2760);
nand U2845 (N_2845,N_2805,N_2810);
or U2846 (N_2846,N_2803,N_2817);
or U2847 (N_2847,N_2782,N_2799);
nand U2848 (N_2848,N_2764,N_2779);
or U2849 (N_2849,N_2798,N_2795);
or U2850 (N_2850,N_2779,N_2785);
nor U2851 (N_2851,N_2806,N_2795);
or U2852 (N_2852,N_2785,N_2799);
and U2853 (N_2853,N_2768,N_2806);
and U2854 (N_2854,N_2783,N_2794);
and U2855 (N_2855,N_2766,N_2782);
nand U2856 (N_2856,N_2795,N_2818);
and U2857 (N_2857,N_2816,N_2817);
and U2858 (N_2858,N_2817,N_2776);
or U2859 (N_2859,N_2805,N_2816);
or U2860 (N_2860,N_2769,N_2780);
and U2861 (N_2861,N_2770,N_2795);
nor U2862 (N_2862,N_2815,N_2766);
or U2863 (N_2863,N_2784,N_2786);
and U2864 (N_2864,N_2779,N_2762);
or U2865 (N_2865,N_2785,N_2767);
nor U2866 (N_2866,N_2818,N_2792);
or U2867 (N_2867,N_2770,N_2785);
nor U2868 (N_2868,N_2774,N_2782);
or U2869 (N_2869,N_2816,N_2814);
nor U2870 (N_2870,N_2801,N_2760);
nand U2871 (N_2871,N_2772,N_2774);
nor U2872 (N_2872,N_2765,N_2780);
nand U2873 (N_2873,N_2808,N_2775);
or U2874 (N_2874,N_2808,N_2810);
nand U2875 (N_2875,N_2779,N_2777);
nor U2876 (N_2876,N_2767,N_2818);
or U2877 (N_2877,N_2794,N_2789);
or U2878 (N_2878,N_2772,N_2766);
and U2879 (N_2879,N_2765,N_2816);
nand U2880 (N_2880,N_2848,N_2833);
and U2881 (N_2881,N_2820,N_2849);
and U2882 (N_2882,N_2874,N_2831);
nor U2883 (N_2883,N_2865,N_2862);
or U2884 (N_2884,N_2827,N_2875);
or U2885 (N_2885,N_2836,N_2829);
or U2886 (N_2886,N_2841,N_2856);
nor U2887 (N_2887,N_2867,N_2845);
nor U2888 (N_2888,N_2852,N_2878);
nand U2889 (N_2889,N_2832,N_2876);
nor U2890 (N_2890,N_2830,N_2853);
nand U2891 (N_2891,N_2858,N_2872);
nand U2892 (N_2892,N_2855,N_2823);
nor U2893 (N_2893,N_2826,N_2879);
or U2894 (N_2894,N_2835,N_2850);
and U2895 (N_2895,N_2834,N_2843);
nand U2896 (N_2896,N_2871,N_2822);
nand U2897 (N_2897,N_2864,N_2854);
and U2898 (N_2898,N_2863,N_2869);
nor U2899 (N_2899,N_2847,N_2866);
nor U2900 (N_2900,N_2839,N_2821);
and U2901 (N_2901,N_2824,N_2840);
nand U2902 (N_2902,N_2828,N_2873);
or U2903 (N_2903,N_2857,N_2837);
nor U2904 (N_2904,N_2868,N_2870);
nor U2905 (N_2905,N_2844,N_2860);
or U2906 (N_2906,N_2825,N_2842);
or U2907 (N_2907,N_2846,N_2859);
and U2908 (N_2908,N_2877,N_2861);
or U2909 (N_2909,N_2838,N_2851);
nand U2910 (N_2910,N_2868,N_2878);
or U2911 (N_2911,N_2870,N_2822);
and U2912 (N_2912,N_2870,N_2852);
and U2913 (N_2913,N_2824,N_2838);
and U2914 (N_2914,N_2849,N_2840);
and U2915 (N_2915,N_2834,N_2825);
and U2916 (N_2916,N_2878,N_2859);
or U2917 (N_2917,N_2871,N_2872);
nand U2918 (N_2918,N_2867,N_2861);
nor U2919 (N_2919,N_2866,N_2857);
nor U2920 (N_2920,N_2823,N_2869);
nand U2921 (N_2921,N_2821,N_2846);
and U2922 (N_2922,N_2830,N_2865);
nor U2923 (N_2923,N_2863,N_2878);
and U2924 (N_2924,N_2837,N_2847);
and U2925 (N_2925,N_2831,N_2852);
nand U2926 (N_2926,N_2843,N_2879);
nand U2927 (N_2927,N_2827,N_2869);
nand U2928 (N_2928,N_2874,N_2828);
nand U2929 (N_2929,N_2876,N_2870);
and U2930 (N_2930,N_2833,N_2826);
nor U2931 (N_2931,N_2834,N_2860);
and U2932 (N_2932,N_2855,N_2822);
and U2933 (N_2933,N_2826,N_2842);
and U2934 (N_2934,N_2846,N_2874);
nand U2935 (N_2935,N_2866,N_2852);
or U2936 (N_2936,N_2835,N_2851);
or U2937 (N_2937,N_2825,N_2838);
and U2938 (N_2938,N_2841,N_2834);
nor U2939 (N_2939,N_2853,N_2866);
nor U2940 (N_2940,N_2927,N_2900);
and U2941 (N_2941,N_2906,N_2909);
and U2942 (N_2942,N_2901,N_2923);
and U2943 (N_2943,N_2889,N_2894);
or U2944 (N_2944,N_2890,N_2912);
nand U2945 (N_2945,N_2905,N_2915);
and U2946 (N_2946,N_2922,N_2917);
and U2947 (N_2947,N_2891,N_2897);
nor U2948 (N_2948,N_2887,N_2895);
or U2949 (N_2949,N_2930,N_2902);
and U2950 (N_2950,N_2918,N_2884);
nand U2951 (N_2951,N_2937,N_2883);
nand U2952 (N_2952,N_2921,N_2924);
and U2953 (N_2953,N_2903,N_2907);
and U2954 (N_2954,N_2911,N_2925);
nor U2955 (N_2955,N_2908,N_2919);
or U2956 (N_2956,N_2939,N_2896);
nor U2957 (N_2957,N_2914,N_2892);
or U2958 (N_2958,N_2932,N_2926);
or U2959 (N_2959,N_2938,N_2886);
or U2960 (N_2960,N_2935,N_2904);
and U2961 (N_2961,N_2882,N_2899);
or U2962 (N_2962,N_2928,N_2885);
or U2963 (N_2963,N_2931,N_2913);
and U2964 (N_2964,N_2916,N_2910);
nand U2965 (N_2965,N_2880,N_2929);
and U2966 (N_2966,N_2898,N_2934);
or U2967 (N_2967,N_2920,N_2893);
xor U2968 (N_2968,N_2936,N_2881);
or U2969 (N_2969,N_2888,N_2933);
and U2970 (N_2970,N_2893,N_2892);
nor U2971 (N_2971,N_2901,N_2893);
nor U2972 (N_2972,N_2931,N_2894);
and U2973 (N_2973,N_2934,N_2913);
and U2974 (N_2974,N_2925,N_2898);
nor U2975 (N_2975,N_2917,N_2891);
nor U2976 (N_2976,N_2906,N_2887);
nand U2977 (N_2977,N_2907,N_2900);
or U2978 (N_2978,N_2905,N_2933);
nand U2979 (N_2979,N_2935,N_2908);
nand U2980 (N_2980,N_2913,N_2881);
and U2981 (N_2981,N_2899,N_2907);
and U2982 (N_2982,N_2889,N_2913);
nor U2983 (N_2983,N_2904,N_2895);
or U2984 (N_2984,N_2935,N_2897);
or U2985 (N_2985,N_2935,N_2928);
or U2986 (N_2986,N_2929,N_2936);
or U2987 (N_2987,N_2894,N_2891);
and U2988 (N_2988,N_2896,N_2927);
or U2989 (N_2989,N_2896,N_2900);
nand U2990 (N_2990,N_2925,N_2936);
and U2991 (N_2991,N_2903,N_2932);
xor U2992 (N_2992,N_2927,N_2934);
or U2993 (N_2993,N_2915,N_2918);
or U2994 (N_2994,N_2880,N_2915);
nor U2995 (N_2995,N_2937,N_2935);
nor U2996 (N_2996,N_2900,N_2934);
or U2997 (N_2997,N_2887,N_2907);
nand U2998 (N_2998,N_2910,N_2886);
nor U2999 (N_2999,N_2904,N_2924);
nor UO_0 (O_0,N_2957,N_2969);
or UO_1 (O_1,N_2959,N_2955);
or UO_2 (O_2,N_2943,N_2954);
nand UO_3 (O_3,N_2987,N_2971);
nor UO_4 (O_4,N_2970,N_2972);
nand UO_5 (O_5,N_2974,N_2941);
nand UO_6 (O_6,N_2944,N_2952);
xnor UO_7 (O_7,N_2982,N_2956);
or UO_8 (O_8,N_2949,N_2967);
nand UO_9 (O_9,N_2977,N_2948);
nor UO_10 (O_10,N_2991,N_2947);
and UO_11 (O_11,N_2950,N_2973);
nor UO_12 (O_12,N_2985,N_2995);
and UO_13 (O_13,N_2979,N_2992);
and UO_14 (O_14,N_2946,N_2965);
xor UO_15 (O_15,N_2966,N_2964);
nand UO_16 (O_16,N_2998,N_2968);
nand UO_17 (O_17,N_2953,N_2990);
nand UO_18 (O_18,N_2942,N_2961);
or UO_19 (O_19,N_2993,N_2981);
and UO_20 (O_20,N_2976,N_2983);
and UO_21 (O_21,N_2984,N_2975);
or UO_22 (O_22,N_2986,N_2999);
and UO_23 (O_23,N_2960,N_2989);
nor UO_24 (O_24,N_2945,N_2958);
nand UO_25 (O_25,N_2978,N_2980);
and UO_26 (O_26,N_2940,N_2996);
or UO_27 (O_27,N_2997,N_2994);
and UO_28 (O_28,N_2951,N_2962);
nand UO_29 (O_29,N_2963,N_2988);
or UO_30 (O_30,N_2995,N_2988);
nand UO_31 (O_31,N_2960,N_2947);
nand UO_32 (O_32,N_2953,N_2970);
and UO_33 (O_33,N_2992,N_2983);
or UO_34 (O_34,N_2943,N_2965);
or UO_35 (O_35,N_2973,N_2941);
xnor UO_36 (O_36,N_2994,N_2983);
and UO_37 (O_37,N_2951,N_2968);
nand UO_38 (O_38,N_2954,N_2972);
or UO_39 (O_39,N_2990,N_2942);
nor UO_40 (O_40,N_2955,N_2965);
and UO_41 (O_41,N_2953,N_2963);
and UO_42 (O_42,N_2968,N_2978);
or UO_43 (O_43,N_2941,N_2991);
nand UO_44 (O_44,N_2990,N_2970);
nand UO_45 (O_45,N_2991,N_2995);
and UO_46 (O_46,N_2957,N_2967);
and UO_47 (O_47,N_2962,N_2954);
and UO_48 (O_48,N_2998,N_2978);
or UO_49 (O_49,N_2968,N_2986);
and UO_50 (O_50,N_2953,N_2977);
or UO_51 (O_51,N_2954,N_2963);
and UO_52 (O_52,N_2975,N_2986);
nor UO_53 (O_53,N_2980,N_2995);
nand UO_54 (O_54,N_2987,N_2943);
nor UO_55 (O_55,N_2964,N_2975);
nand UO_56 (O_56,N_2963,N_2946);
nor UO_57 (O_57,N_2989,N_2966);
nand UO_58 (O_58,N_2968,N_2960);
or UO_59 (O_59,N_2990,N_2984);
and UO_60 (O_60,N_2966,N_2992);
nand UO_61 (O_61,N_2963,N_2984);
nand UO_62 (O_62,N_2988,N_2979);
or UO_63 (O_63,N_2947,N_2957);
or UO_64 (O_64,N_2984,N_2947);
nand UO_65 (O_65,N_2991,N_2960);
nand UO_66 (O_66,N_2964,N_2946);
nand UO_67 (O_67,N_2955,N_2966);
nand UO_68 (O_68,N_2991,N_2967);
and UO_69 (O_69,N_2952,N_2990);
nand UO_70 (O_70,N_2987,N_2979);
and UO_71 (O_71,N_2950,N_2967);
nor UO_72 (O_72,N_2983,N_2962);
and UO_73 (O_73,N_2948,N_2942);
nor UO_74 (O_74,N_2979,N_2960);
or UO_75 (O_75,N_2963,N_2957);
nor UO_76 (O_76,N_2981,N_2982);
nand UO_77 (O_77,N_2976,N_2971);
and UO_78 (O_78,N_2945,N_2978);
nand UO_79 (O_79,N_2998,N_2941);
nor UO_80 (O_80,N_2985,N_2958);
nor UO_81 (O_81,N_2978,N_2997);
nor UO_82 (O_82,N_2949,N_2948);
or UO_83 (O_83,N_2942,N_2963);
or UO_84 (O_84,N_2982,N_2969);
nand UO_85 (O_85,N_2944,N_2956);
and UO_86 (O_86,N_2990,N_2973);
nor UO_87 (O_87,N_2990,N_2994);
and UO_88 (O_88,N_2994,N_2964);
or UO_89 (O_89,N_2978,N_2970);
or UO_90 (O_90,N_2981,N_2956);
nor UO_91 (O_91,N_2970,N_2998);
and UO_92 (O_92,N_2956,N_2997);
nand UO_93 (O_93,N_2988,N_2980);
nand UO_94 (O_94,N_2965,N_2987);
nor UO_95 (O_95,N_2999,N_2985);
or UO_96 (O_96,N_2998,N_2983);
nand UO_97 (O_97,N_2987,N_2998);
nand UO_98 (O_98,N_2940,N_2993);
or UO_99 (O_99,N_2983,N_2955);
and UO_100 (O_100,N_2941,N_2982);
and UO_101 (O_101,N_2986,N_2979);
and UO_102 (O_102,N_2988,N_2957);
and UO_103 (O_103,N_2988,N_2960);
nand UO_104 (O_104,N_2947,N_2998);
nand UO_105 (O_105,N_2969,N_2960);
or UO_106 (O_106,N_2993,N_2965);
or UO_107 (O_107,N_2993,N_2986);
and UO_108 (O_108,N_2956,N_2968);
nand UO_109 (O_109,N_2966,N_2993);
nand UO_110 (O_110,N_2994,N_2977);
nor UO_111 (O_111,N_2942,N_2992);
nor UO_112 (O_112,N_2947,N_2958);
and UO_113 (O_113,N_2973,N_2982);
or UO_114 (O_114,N_2989,N_2973);
nor UO_115 (O_115,N_2992,N_2989);
and UO_116 (O_116,N_2969,N_2977);
nor UO_117 (O_117,N_2966,N_2942);
nor UO_118 (O_118,N_2992,N_2952);
nor UO_119 (O_119,N_2981,N_2970);
and UO_120 (O_120,N_2943,N_2967);
nand UO_121 (O_121,N_2969,N_2968);
nand UO_122 (O_122,N_2974,N_2952);
nor UO_123 (O_123,N_2940,N_2960);
and UO_124 (O_124,N_2979,N_2971);
or UO_125 (O_125,N_2995,N_2963);
and UO_126 (O_126,N_2979,N_2995);
or UO_127 (O_127,N_2950,N_2992);
nor UO_128 (O_128,N_2957,N_2991);
nor UO_129 (O_129,N_2974,N_2962);
or UO_130 (O_130,N_2950,N_2986);
and UO_131 (O_131,N_2976,N_2955);
or UO_132 (O_132,N_2949,N_2955);
and UO_133 (O_133,N_2954,N_2958);
and UO_134 (O_134,N_2951,N_2997);
or UO_135 (O_135,N_2959,N_2949);
nor UO_136 (O_136,N_2959,N_2947);
or UO_137 (O_137,N_2993,N_2971);
or UO_138 (O_138,N_2944,N_2957);
or UO_139 (O_139,N_2984,N_2958);
nor UO_140 (O_140,N_2945,N_2990);
and UO_141 (O_141,N_2965,N_2957);
nand UO_142 (O_142,N_2992,N_2958);
nand UO_143 (O_143,N_2955,N_2957);
or UO_144 (O_144,N_2950,N_2945);
and UO_145 (O_145,N_2969,N_2996);
nand UO_146 (O_146,N_2987,N_2956);
nand UO_147 (O_147,N_2994,N_2973);
nor UO_148 (O_148,N_2945,N_2960);
and UO_149 (O_149,N_2998,N_2980);
or UO_150 (O_150,N_2987,N_2977);
nand UO_151 (O_151,N_2964,N_2978);
nand UO_152 (O_152,N_2967,N_2951);
nor UO_153 (O_153,N_2978,N_2951);
or UO_154 (O_154,N_2989,N_2946);
or UO_155 (O_155,N_2954,N_2992);
nand UO_156 (O_156,N_2972,N_2952);
nor UO_157 (O_157,N_2985,N_2951);
or UO_158 (O_158,N_2957,N_2942);
or UO_159 (O_159,N_2988,N_2976);
nor UO_160 (O_160,N_2969,N_2941);
nand UO_161 (O_161,N_2968,N_2975);
nor UO_162 (O_162,N_2960,N_2946);
and UO_163 (O_163,N_2975,N_2987);
nor UO_164 (O_164,N_2956,N_2966);
nor UO_165 (O_165,N_2994,N_2957);
nor UO_166 (O_166,N_2942,N_2995);
and UO_167 (O_167,N_2990,N_2951);
nand UO_168 (O_168,N_2969,N_2993);
or UO_169 (O_169,N_2948,N_2960);
and UO_170 (O_170,N_2988,N_2962);
nand UO_171 (O_171,N_2983,N_2961);
nand UO_172 (O_172,N_2956,N_2989);
or UO_173 (O_173,N_2981,N_2984);
or UO_174 (O_174,N_2990,N_2996);
nor UO_175 (O_175,N_2982,N_2993);
or UO_176 (O_176,N_2955,N_2995);
and UO_177 (O_177,N_2973,N_2958);
nor UO_178 (O_178,N_2945,N_2970);
and UO_179 (O_179,N_2987,N_2963);
xnor UO_180 (O_180,N_2961,N_2979);
or UO_181 (O_181,N_2992,N_2975);
or UO_182 (O_182,N_2966,N_2948);
nand UO_183 (O_183,N_2945,N_2966);
and UO_184 (O_184,N_2949,N_2991);
or UO_185 (O_185,N_2985,N_2987);
or UO_186 (O_186,N_2995,N_2954);
or UO_187 (O_187,N_2946,N_2966);
nand UO_188 (O_188,N_2991,N_2972);
or UO_189 (O_189,N_2960,N_2973);
or UO_190 (O_190,N_2999,N_2969);
and UO_191 (O_191,N_2975,N_2949);
nand UO_192 (O_192,N_2992,N_2940);
nor UO_193 (O_193,N_2947,N_2973);
or UO_194 (O_194,N_2963,N_2969);
nor UO_195 (O_195,N_2988,N_2971);
nor UO_196 (O_196,N_2968,N_2944);
and UO_197 (O_197,N_2997,N_2970);
nor UO_198 (O_198,N_2972,N_2994);
nand UO_199 (O_199,N_2993,N_2951);
nor UO_200 (O_200,N_2961,N_2958);
and UO_201 (O_201,N_2997,N_2966);
and UO_202 (O_202,N_2982,N_2950);
nor UO_203 (O_203,N_2985,N_2975);
and UO_204 (O_204,N_2970,N_2994);
nor UO_205 (O_205,N_2969,N_2949);
nor UO_206 (O_206,N_2970,N_2974);
and UO_207 (O_207,N_2975,N_2947);
nor UO_208 (O_208,N_2968,N_2980);
or UO_209 (O_209,N_2942,N_2979);
and UO_210 (O_210,N_2950,N_2955);
and UO_211 (O_211,N_2970,N_2955);
or UO_212 (O_212,N_2972,N_2956);
nand UO_213 (O_213,N_2993,N_2994);
or UO_214 (O_214,N_2971,N_2963);
nor UO_215 (O_215,N_2971,N_2974);
or UO_216 (O_216,N_2965,N_2990);
nand UO_217 (O_217,N_2962,N_2969);
nand UO_218 (O_218,N_2960,N_2980);
or UO_219 (O_219,N_2988,N_2984);
nand UO_220 (O_220,N_2973,N_2998);
nand UO_221 (O_221,N_2971,N_2994);
nor UO_222 (O_222,N_2972,N_2969);
or UO_223 (O_223,N_2995,N_2947);
nand UO_224 (O_224,N_2997,N_2961);
nand UO_225 (O_225,N_2980,N_2977);
nor UO_226 (O_226,N_2969,N_2989);
nand UO_227 (O_227,N_2964,N_2969);
or UO_228 (O_228,N_2990,N_2978);
nand UO_229 (O_229,N_2991,N_2968);
and UO_230 (O_230,N_2952,N_2976);
nand UO_231 (O_231,N_2974,N_2993);
nor UO_232 (O_232,N_2967,N_2953);
nor UO_233 (O_233,N_2941,N_2952);
nor UO_234 (O_234,N_2973,N_2949);
and UO_235 (O_235,N_2983,N_2949);
and UO_236 (O_236,N_2968,N_2958);
nor UO_237 (O_237,N_2957,N_2997);
or UO_238 (O_238,N_2987,N_2941);
nor UO_239 (O_239,N_2980,N_2983);
nor UO_240 (O_240,N_2959,N_2977);
nand UO_241 (O_241,N_2950,N_2941);
nand UO_242 (O_242,N_2996,N_2980);
or UO_243 (O_243,N_2953,N_2983);
or UO_244 (O_244,N_2996,N_2962);
and UO_245 (O_245,N_2940,N_2988);
or UO_246 (O_246,N_2974,N_2949);
nor UO_247 (O_247,N_2992,N_2948);
and UO_248 (O_248,N_2995,N_2940);
and UO_249 (O_249,N_2972,N_2962);
nand UO_250 (O_250,N_2983,N_2971);
nor UO_251 (O_251,N_2966,N_2986);
nand UO_252 (O_252,N_2949,N_2992);
and UO_253 (O_253,N_2987,N_2997);
nor UO_254 (O_254,N_2956,N_2962);
or UO_255 (O_255,N_2973,N_2956);
or UO_256 (O_256,N_2952,N_2947);
nand UO_257 (O_257,N_2965,N_2988);
or UO_258 (O_258,N_2941,N_2968);
or UO_259 (O_259,N_2972,N_2964);
nand UO_260 (O_260,N_2953,N_2966);
and UO_261 (O_261,N_2952,N_2983);
and UO_262 (O_262,N_2974,N_2943);
or UO_263 (O_263,N_2948,N_2959);
nor UO_264 (O_264,N_2985,N_2976);
nor UO_265 (O_265,N_2982,N_2992);
nor UO_266 (O_266,N_2946,N_2959);
nor UO_267 (O_267,N_2950,N_2987);
and UO_268 (O_268,N_2977,N_2944);
nand UO_269 (O_269,N_2944,N_2969);
nor UO_270 (O_270,N_2941,N_2957);
nor UO_271 (O_271,N_2963,N_2947);
nor UO_272 (O_272,N_2962,N_2994);
or UO_273 (O_273,N_2960,N_2958);
or UO_274 (O_274,N_2972,N_2990);
nand UO_275 (O_275,N_2962,N_2977);
nor UO_276 (O_276,N_2942,N_2973);
or UO_277 (O_277,N_2982,N_2961);
and UO_278 (O_278,N_2963,N_2948);
and UO_279 (O_279,N_2991,N_2965);
or UO_280 (O_280,N_2944,N_2974);
nor UO_281 (O_281,N_2946,N_2955);
and UO_282 (O_282,N_2980,N_2945);
nand UO_283 (O_283,N_2966,N_2981);
nand UO_284 (O_284,N_2966,N_2940);
or UO_285 (O_285,N_2988,N_2956);
nor UO_286 (O_286,N_2960,N_2995);
nand UO_287 (O_287,N_2950,N_2951);
nor UO_288 (O_288,N_2987,N_2986);
nor UO_289 (O_289,N_2943,N_2999);
nand UO_290 (O_290,N_2999,N_2945);
nand UO_291 (O_291,N_2956,N_2961);
nand UO_292 (O_292,N_2981,N_2942);
nor UO_293 (O_293,N_2984,N_2942);
or UO_294 (O_294,N_2975,N_2959);
or UO_295 (O_295,N_2984,N_2987);
nand UO_296 (O_296,N_2950,N_2980);
or UO_297 (O_297,N_2980,N_2952);
nor UO_298 (O_298,N_2963,N_2952);
and UO_299 (O_299,N_2956,N_2942);
and UO_300 (O_300,N_2959,N_2990);
and UO_301 (O_301,N_2955,N_2981);
and UO_302 (O_302,N_2946,N_2997);
nand UO_303 (O_303,N_2998,N_2962);
nor UO_304 (O_304,N_2959,N_2976);
nor UO_305 (O_305,N_2995,N_2972);
or UO_306 (O_306,N_2997,N_2955);
or UO_307 (O_307,N_2952,N_2940);
nand UO_308 (O_308,N_2986,N_2997);
nor UO_309 (O_309,N_2971,N_2954);
or UO_310 (O_310,N_2993,N_2948);
and UO_311 (O_311,N_2951,N_2971);
nor UO_312 (O_312,N_2976,N_2995);
or UO_313 (O_313,N_2996,N_2987);
nor UO_314 (O_314,N_2995,N_2981);
or UO_315 (O_315,N_2987,N_2980);
nand UO_316 (O_316,N_2997,N_2960);
nor UO_317 (O_317,N_2963,N_2958);
nand UO_318 (O_318,N_2949,N_2968);
and UO_319 (O_319,N_2966,N_2970);
nor UO_320 (O_320,N_2995,N_2967);
or UO_321 (O_321,N_2994,N_2982);
nand UO_322 (O_322,N_2987,N_2945);
or UO_323 (O_323,N_2950,N_2940);
or UO_324 (O_324,N_2985,N_2963);
and UO_325 (O_325,N_2989,N_2958);
and UO_326 (O_326,N_2983,N_2970);
nor UO_327 (O_327,N_2979,N_2946);
nor UO_328 (O_328,N_2943,N_2941);
and UO_329 (O_329,N_2971,N_2978);
and UO_330 (O_330,N_2993,N_2996);
and UO_331 (O_331,N_2983,N_2989);
nor UO_332 (O_332,N_2953,N_2961);
or UO_333 (O_333,N_2941,N_2955);
nor UO_334 (O_334,N_2967,N_2942);
or UO_335 (O_335,N_2997,N_2995);
nor UO_336 (O_336,N_2988,N_2955);
or UO_337 (O_337,N_2969,N_2947);
or UO_338 (O_338,N_2996,N_2954);
nand UO_339 (O_339,N_2985,N_2968);
nand UO_340 (O_340,N_2971,N_2970);
and UO_341 (O_341,N_2987,N_2988);
nand UO_342 (O_342,N_2953,N_2948);
nor UO_343 (O_343,N_2959,N_2981);
and UO_344 (O_344,N_2950,N_2946);
nor UO_345 (O_345,N_2969,N_2961);
nand UO_346 (O_346,N_2957,N_2982);
and UO_347 (O_347,N_2949,N_2940);
nor UO_348 (O_348,N_2943,N_2946);
nor UO_349 (O_349,N_2994,N_2989);
and UO_350 (O_350,N_2975,N_2958);
and UO_351 (O_351,N_2996,N_2975);
nand UO_352 (O_352,N_2972,N_2960);
nor UO_353 (O_353,N_2950,N_2943);
or UO_354 (O_354,N_2947,N_2988);
or UO_355 (O_355,N_2967,N_2978);
nand UO_356 (O_356,N_2981,N_2963);
and UO_357 (O_357,N_2989,N_2952);
and UO_358 (O_358,N_2963,N_2956);
and UO_359 (O_359,N_2978,N_2981);
nor UO_360 (O_360,N_2984,N_2991);
nand UO_361 (O_361,N_2979,N_2989);
nand UO_362 (O_362,N_2988,N_2967);
and UO_363 (O_363,N_2980,N_2986);
and UO_364 (O_364,N_2983,N_2967);
nand UO_365 (O_365,N_2974,N_2954);
nor UO_366 (O_366,N_2961,N_2949);
or UO_367 (O_367,N_2994,N_2995);
nand UO_368 (O_368,N_2995,N_2945);
or UO_369 (O_369,N_2981,N_2964);
and UO_370 (O_370,N_2948,N_2952);
and UO_371 (O_371,N_2947,N_2941);
and UO_372 (O_372,N_2948,N_2975);
or UO_373 (O_373,N_2981,N_2997);
nor UO_374 (O_374,N_2994,N_2966);
nand UO_375 (O_375,N_2959,N_2987);
and UO_376 (O_376,N_2957,N_2951);
nand UO_377 (O_377,N_2971,N_2984);
and UO_378 (O_378,N_2954,N_2987);
nor UO_379 (O_379,N_2976,N_2951);
nand UO_380 (O_380,N_2993,N_2949);
and UO_381 (O_381,N_2999,N_2965);
or UO_382 (O_382,N_2945,N_2959);
nand UO_383 (O_383,N_2948,N_2974);
and UO_384 (O_384,N_2984,N_2964);
nor UO_385 (O_385,N_2965,N_2996);
nand UO_386 (O_386,N_2951,N_2989);
nand UO_387 (O_387,N_2959,N_2951);
or UO_388 (O_388,N_2987,N_2992);
nand UO_389 (O_389,N_2984,N_2976);
nand UO_390 (O_390,N_2980,N_2958);
and UO_391 (O_391,N_2949,N_2990);
or UO_392 (O_392,N_2970,N_2943);
nand UO_393 (O_393,N_2991,N_2971);
nor UO_394 (O_394,N_2941,N_2959);
nand UO_395 (O_395,N_2977,N_2986);
nand UO_396 (O_396,N_2966,N_2969);
nand UO_397 (O_397,N_2993,N_2973);
and UO_398 (O_398,N_2951,N_2944);
and UO_399 (O_399,N_2970,N_2964);
or UO_400 (O_400,N_2999,N_2987);
nand UO_401 (O_401,N_2982,N_2985);
and UO_402 (O_402,N_2978,N_2953);
and UO_403 (O_403,N_2940,N_2973);
and UO_404 (O_404,N_2999,N_2977);
nand UO_405 (O_405,N_2964,N_2988);
nand UO_406 (O_406,N_2976,N_2942);
nand UO_407 (O_407,N_2975,N_2967);
or UO_408 (O_408,N_2998,N_2993);
xor UO_409 (O_409,N_2988,N_2998);
and UO_410 (O_410,N_2981,N_2965);
nor UO_411 (O_411,N_2992,N_2971);
nand UO_412 (O_412,N_2964,N_2968);
nor UO_413 (O_413,N_2987,N_2968);
and UO_414 (O_414,N_2961,N_2964);
and UO_415 (O_415,N_2953,N_2998);
or UO_416 (O_416,N_2948,N_2951);
and UO_417 (O_417,N_2992,N_2997);
nand UO_418 (O_418,N_2978,N_2969);
nor UO_419 (O_419,N_2941,N_2996);
nor UO_420 (O_420,N_2999,N_2964);
nand UO_421 (O_421,N_2985,N_2980);
nor UO_422 (O_422,N_2946,N_2977);
nor UO_423 (O_423,N_2981,N_2985);
nand UO_424 (O_424,N_2961,N_2941);
or UO_425 (O_425,N_2978,N_2940);
nor UO_426 (O_426,N_2998,N_2961);
or UO_427 (O_427,N_2954,N_2984);
and UO_428 (O_428,N_2960,N_2999);
nand UO_429 (O_429,N_2982,N_2978);
or UO_430 (O_430,N_2999,N_2976);
and UO_431 (O_431,N_2976,N_2996);
or UO_432 (O_432,N_2970,N_2942);
nor UO_433 (O_433,N_2960,N_2956);
and UO_434 (O_434,N_2955,N_2967);
or UO_435 (O_435,N_2992,N_2986);
or UO_436 (O_436,N_2968,N_2993);
and UO_437 (O_437,N_2951,N_2952);
nor UO_438 (O_438,N_2942,N_2958);
nor UO_439 (O_439,N_2988,N_2985);
and UO_440 (O_440,N_2952,N_2945);
and UO_441 (O_441,N_2942,N_2953);
nor UO_442 (O_442,N_2961,N_2943);
nand UO_443 (O_443,N_2973,N_2970);
nor UO_444 (O_444,N_2948,N_2955);
or UO_445 (O_445,N_2970,N_2969);
or UO_446 (O_446,N_2985,N_2948);
or UO_447 (O_447,N_2960,N_2950);
nand UO_448 (O_448,N_2946,N_2970);
or UO_449 (O_449,N_2993,N_2964);
and UO_450 (O_450,N_2940,N_2947);
or UO_451 (O_451,N_2951,N_2996);
nor UO_452 (O_452,N_2984,N_2973);
nor UO_453 (O_453,N_2959,N_2952);
nor UO_454 (O_454,N_2977,N_2961);
or UO_455 (O_455,N_2969,N_2986);
or UO_456 (O_456,N_2973,N_2944);
nand UO_457 (O_457,N_2988,N_2953);
or UO_458 (O_458,N_2964,N_2948);
nor UO_459 (O_459,N_2990,N_2962);
nand UO_460 (O_460,N_2965,N_2967);
or UO_461 (O_461,N_2996,N_2956);
or UO_462 (O_462,N_2989,N_2942);
or UO_463 (O_463,N_2983,N_2982);
or UO_464 (O_464,N_2948,N_2976);
nor UO_465 (O_465,N_2941,N_2948);
or UO_466 (O_466,N_2962,N_2949);
nand UO_467 (O_467,N_2956,N_2946);
or UO_468 (O_468,N_2993,N_2988);
or UO_469 (O_469,N_2991,N_2993);
nor UO_470 (O_470,N_2975,N_2978);
and UO_471 (O_471,N_2963,N_2989);
nor UO_472 (O_472,N_2996,N_2946);
nand UO_473 (O_473,N_2972,N_2980);
or UO_474 (O_474,N_2971,N_2965);
and UO_475 (O_475,N_2941,N_2997);
and UO_476 (O_476,N_2966,N_2987);
or UO_477 (O_477,N_2994,N_2967);
and UO_478 (O_478,N_2989,N_2967);
nor UO_479 (O_479,N_2974,N_2994);
or UO_480 (O_480,N_2945,N_2989);
nor UO_481 (O_481,N_2972,N_2967);
nand UO_482 (O_482,N_2945,N_2951);
or UO_483 (O_483,N_2999,N_2978);
and UO_484 (O_484,N_2966,N_2980);
nand UO_485 (O_485,N_2994,N_2955);
and UO_486 (O_486,N_2959,N_2982);
or UO_487 (O_487,N_2986,N_2948);
nor UO_488 (O_488,N_2965,N_2956);
nand UO_489 (O_489,N_2962,N_2965);
nor UO_490 (O_490,N_2981,N_2986);
or UO_491 (O_491,N_2944,N_2965);
and UO_492 (O_492,N_2981,N_2996);
nor UO_493 (O_493,N_2947,N_2970);
nor UO_494 (O_494,N_2943,N_2992);
nor UO_495 (O_495,N_2996,N_2972);
and UO_496 (O_496,N_2948,N_2968);
or UO_497 (O_497,N_2995,N_2973);
and UO_498 (O_498,N_2994,N_2944);
or UO_499 (O_499,N_2958,N_2995);
endmodule