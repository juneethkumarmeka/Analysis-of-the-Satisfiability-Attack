module basic_750_5000_1000_25_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_376,In_312);
nand U1 (N_1,In_11,In_443);
or U2 (N_2,In_322,In_703);
nor U3 (N_3,In_553,In_237);
nor U4 (N_4,In_184,In_699);
nand U5 (N_5,In_556,In_676);
nor U6 (N_6,In_387,In_537);
and U7 (N_7,In_209,In_632);
and U8 (N_8,In_68,In_300);
and U9 (N_9,In_23,In_308);
or U10 (N_10,In_539,In_18);
and U11 (N_11,In_151,In_395);
or U12 (N_12,In_232,In_79);
and U13 (N_13,In_313,In_275);
or U14 (N_14,In_270,In_586);
nand U15 (N_15,In_114,In_630);
nand U16 (N_16,In_32,In_233);
nor U17 (N_17,In_574,In_545);
and U18 (N_18,In_656,In_616);
or U19 (N_19,In_50,In_37);
nor U20 (N_20,In_249,In_123);
and U21 (N_21,In_567,In_364);
nor U22 (N_22,In_548,In_621);
and U23 (N_23,In_712,In_116);
or U24 (N_24,In_602,In_399);
and U25 (N_25,In_347,In_671);
nand U26 (N_26,In_659,In_730);
nor U27 (N_27,In_409,In_558);
and U28 (N_28,In_670,In_277);
and U29 (N_29,In_113,In_133);
nor U30 (N_30,In_278,In_637);
nor U31 (N_31,In_49,In_696);
and U32 (N_32,In_500,In_138);
nor U33 (N_33,In_326,In_431);
nor U34 (N_34,In_693,In_361);
nor U35 (N_35,In_413,In_101);
nand U36 (N_36,In_236,In_441);
or U37 (N_37,In_69,In_746);
or U38 (N_38,In_723,In_144);
and U39 (N_39,In_107,In_108);
nor U40 (N_40,In_664,In_105);
nor U41 (N_41,In_36,In_421);
and U42 (N_42,In_345,In_6);
or U43 (N_43,In_305,In_285);
and U44 (N_44,In_515,In_747);
nand U45 (N_45,In_672,In_43);
and U46 (N_46,In_17,In_77);
and U47 (N_47,In_620,In_562);
nor U48 (N_48,In_212,In_555);
nand U49 (N_49,In_743,In_609);
nor U50 (N_50,In_241,In_647);
and U51 (N_51,In_150,In_328);
nand U52 (N_52,In_367,In_135);
or U53 (N_53,In_454,In_463);
nand U54 (N_54,In_452,In_280);
nor U55 (N_55,In_502,In_360);
or U56 (N_56,In_461,In_149);
or U57 (N_57,In_47,In_682);
nor U58 (N_58,In_170,In_388);
nor U59 (N_59,In_97,In_412);
nand U60 (N_60,In_286,In_271);
nor U61 (N_61,In_717,In_284);
xnor U62 (N_62,In_343,In_62);
and U63 (N_63,In_119,In_147);
nor U64 (N_64,In_171,In_531);
and U65 (N_65,In_614,In_464);
nand U66 (N_66,In_336,In_268);
and U67 (N_67,In_686,In_642);
or U68 (N_68,In_509,In_530);
or U69 (N_69,In_91,In_125);
and U70 (N_70,In_207,In_707);
nor U71 (N_71,In_60,In_87);
or U72 (N_72,In_456,In_424);
nand U73 (N_73,In_403,In_708);
nor U74 (N_74,In_635,In_475);
nor U75 (N_75,In_155,In_660);
nor U76 (N_76,In_64,In_302);
nor U77 (N_77,In_615,In_414);
nor U78 (N_78,In_710,In_472);
nand U79 (N_79,In_134,In_401);
nor U80 (N_80,In_473,In_365);
nor U81 (N_81,In_396,In_73);
and U82 (N_82,In_353,In_75);
and U83 (N_83,In_422,In_356);
or U84 (N_84,In_53,In_222);
and U85 (N_85,In_481,In_718);
nand U86 (N_86,In_220,In_593);
and U87 (N_87,In_380,In_583);
and U88 (N_88,In_433,In_645);
nor U89 (N_89,In_164,In_569);
nor U90 (N_90,In_375,In_89);
nand U91 (N_91,In_181,In_327);
nand U92 (N_92,In_226,In_467);
nand U93 (N_93,In_216,In_8);
nand U94 (N_94,In_366,In_82);
nor U95 (N_95,In_315,In_223);
and U96 (N_96,In_253,In_294);
nand U97 (N_97,In_261,In_72);
nand U98 (N_98,In_158,In_288);
and U99 (N_99,In_483,In_4);
nor U100 (N_100,In_404,In_344);
nor U101 (N_101,In_435,In_38);
and U102 (N_102,In_355,In_596);
nand U103 (N_103,In_160,In_229);
or U104 (N_104,In_332,In_653);
and U105 (N_105,In_319,In_157);
or U106 (N_106,In_126,In_678);
nor U107 (N_107,In_745,In_522);
nor U108 (N_108,In_691,In_242);
and U109 (N_109,In_316,In_254);
and U110 (N_110,In_67,In_384);
and U111 (N_111,In_186,In_304);
nand U112 (N_112,In_398,In_694);
or U113 (N_113,In_425,In_243);
and U114 (N_114,In_208,In_100);
nor U115 (N_115,In_440,In_546);
and U116 (N_116,In_202,In_183);
and U117 (N_117,In_489,In_71);
and U118 (N_118,In_26,In_371);
and U119 (N_119,In_31,In_564);
or U120 (N_120,In_258,In_468);
nand U121 (N_121,In_27,In_448);
nand U122 (N_122,In_102,In_78);
nand U123 (N_123,In_514,In_10);
nor U124 (N_124,In_57,In_311);
nor U125 (N_125,In_307,In_737);
nand U126 (N_126,In_634,In_290);
nor U127 (N_127,In_504,In_111);
and U128 (N_128,In_442,In_650);
nor U129 (N_129,In_195,In_188);
and U130 (N_130,In_550,In_154);
nand U131 (N_131,In_20,In_695);
nand U132 (N_132,In_638,In_698);
nor U133 (N_133,In_495,In_684);
nand U134 (N_134,In_210,In_118);
nor U135 (N_135,In_219,In_667);
and U136 (N_136,In_370,In_628);
and U137 (N_137,In_320,In_196);
nand U138 (N_138,In_636,In_655);
nand U139 (N_139,In_559,In_449);
or U140 (N_140,In_629,In_225);
or U141 (N_141,In_625,In_30);
nor U142 (N_142,In_103,In_543);
and U143 (N_143,In_257,In_16);
or U144 (N_144,In_457,In_681);
nand U145 (N_145,In_402,In_604);
nor U146 (N_146,In_148,In_458);
nand U147 (N_147,In_534,In_644);
or U148 (N_148,In_520,In_488);
or U149 (N_149,In_14,In_675);
nor U150 (N_150,In_211,In_3);
nor U151 (N_151,In_45,In_266);
or U152 (N_152,In_214,In_643);
nor U153 (N_153,In_189,In_131);
or U154 (N_154,In_466,In_627);
nor U155 (N_155,In_446,In_329);
nor U156 (N_156,In_600,In_436);
and U157 (N_157,In_339,In_714);
nor U158 (N_158,In_680,In_601);
or U159 (N_159,In_540,In_617);
nand U160 (N_160,In_581,In_174);
nand U161 (N_161,In_267,In_706);
nand U162 (N_162,In_649,In_206);
nor U163 (N_163,In_631,In_83);
nand U164 (N_164,In_21,In_362);
and U165 (N_165,In_470,In_231);
or U166 (N_166,In_727,In_416);
nand U167 (N_167,In_679,In_462);
nand U168 (N_168,In_74,In_608);
or U169 (N_169,In_245,In_56);
nor U170 (N_170,In_142,In_692);
or U171 (N_171,In_39,In_527);
nor U172 (N_172,In_390,In_611);
nor U173 (N_173,In_51,In_244);
nand U174 (N_174,In_544,In_44);
and U175 (N_175,In_169,In_197);
or U176 (N_176,In_263,In_742);
and U177 (N_177,In_22,In_391);
and U178 (N_178,In_256,In_265);
nand U179 (N_179,In_292,In_494);
nor U180 (N_180,In_552,In_110);
and U181 (N_181,In_283,In_333);
nor U182 (N_182,In_260,In_287);
or U183 (N_183,In_410,In_598);
or U184 (N_184,In_106,In_240);
nor U185 (N_185,In_591,In_640);
and U186 (N_186,In_704,In_505);
nand U187 (N_187,In_733,In_182);
nand U188 (N_188,In_112,In_748);
nor U189 (N_189,In_507,In_377);
xnor U190 (N_190,In_324,In_81);
or U191 (N_191,In_687,In_622);
nand U192 (N_192,In_354,In_274);
nand U193 (N_193,In_716,In_582);
nor U194 (N_194,In_536,In_584);
nor U195 (N_195,In_291,In_549);
or U196 (N_196,In_340,In_603);
nand U197 (N_197,In_426,In_688);
nand U198 (N_198,In_535,In_476);
nand U199 (N_199,In_646,In_34);
nor U200 (N_200,In_25,In_94);
or U201 (N_201,In_683,N_56);
or U202 (N_202,In_29,N_118);
nor U203 (N_203,N_148,In_690);
or U204 (N_204,N_182,In_2);
nor U205 (N_205,In_289,In_215);
nor U206 (N_206,N_175,N_146);
nand U207 (N_207,In_378,N_60);
nor U208 (N_208,In_415,N_188);
and U209 (N_209,N_168,In_173);
and U210 (N_210,In_735,In_613);
or U211 (N_211,N_120,N_173);
nor U212 (N_212,N_165,N_104);
nor U213 (N_213,In_374,In_651);
nor U214 (N_214,N_147,In_33);
nand U215 (N_215,In_120,N_59);
nand U216 (N_216,N_68,In_230);
and U217 (N_217,In_477,In_610);
or U218 (N_218,In_262,N_199);
or U219 (N_219,N_99,In_565);
or U220 (N_220,In_12,In_547);
or U221 (N_221,N_55,N_44);
and U222 (N_222,N_110,In_619);
nand U223 (N_223,In_512,In_529);
and U224 (N_224,In_542,In_92);
nand U225 (N_225,N_142,In_41);
or U226 (N_226,N_181,In_363);
nand U227 (N_227,In_314,N_162);
or U228 (N_228,In_573,In_238);
nand U229 (N_229,In_255,In_204);
and U230 (N_230,In_162,N_139);
and U231 (N_231,In_523,N_155);
nor U232 (N_232,N_54,In_471);
or U233 (N_233,In_342,In_579);
nor U234 (N_234,In_568,N_1);
nand U235 (N_235,In_427,In_297);
or U236 (N_236,In_439,In_348);
and U237 (N_237,N_167,N_82);
or U238 (N_238,In_589,In_503);
or U239 (N_239,N_169,N_96);
nand U240 (N_240,N_171,In_0);
nand U241 (N_241,N_40,In_729);
or U242 (N_242,N_183,In_478);
or U243 (N_243,N_77,In_459);
or U244 (N_244,In_1,N_144);
nor U245 (N_245,In_161,In_259);
nand U246 (N_246,N_16,In_55);
and U247 (N_247,In_666,In_741);
nor U248 (N_248,In_251,N_8);
and U249 (N_249,In_84,In_423);
or U250 (N_250,In_334,In_654);
nand U251 (N_251,In_176,N_97);
nor U252 (N_252,N_117,In_63);
and U253 (N_253,N_29,In_234);
and U254 (N_254,In_217,In_331);
nor U255 (N_255,N_137,In_595);
or U256 (N_256,In_299,In_563);
nor U257 (N_257,N_47,In_557);
nor U258 (N_258,In_734,In_357);
nor U259 (N_259,In_213,In_321);
xnor U260 (N_260,In_194,N_161);
and U261 (N_261,N_86,In_411);
or U262 (N_262,In_434,In_715);
or U263 (N_263,N_37,N_102);
xor U264 (N_264,In_175,N_71);
and U265 (N_265,In_590,N_46);
or U266 (N_266,N_191,In_479);
nor U267 (N_267,In_137,N_128);
and U268 (N_268,N_95,N_195);
or U269 (N_269,In_430,In_235);
or U270 (N_270,In_740,In_95);
nor U271 (N_271,In_199,In_187);
or U272 (N_272,In_652,In_533);
nor U273 (N_273,N_185,In_351);
and U274 (N_274,N_19,In_524);
nand U275 (N_275,In_246,In_618);
nor U276 (N_276,In_393,N_126);
or U277 (N_277,N_35,In_517);
or U278 (N_278,In_372,In_571);
nor U279 (N_279,In_382,In_228);
or U280 (N_280,In_224,N_66);
and U281 (N_281,In_469,In_480);
or U282 (N_282,N_52,N_23);
or U283 (N_283,In_658,N_27);
nor U284 (N_284,In_205,In_521);
or U285 (N_285,In_491,In_685);
nor U286 (N_286,In_657,In_335);
nand U287 (N_287,In_191,In_561);
nor U288 (N_288,N_133,In_541);
nand U289 (N_289,In_420,In_177);
and U290 (N_290,In_178,N_41);
or U291 (N_291,In_48,In_310);
and U292 (N_292,In_484,In_373);
and U293 (N_293,N_134,N_65);
nor U294 (N_294,In_725,In_368);
nor U295 (N_295,In_570,N_93);
nand U296 (N_296,In_510,In_247);
or U297 (N_297,N_62,In_381);
nor U298 (N_298,In_624,In_295);
nor U299 (N_299,In_732,In_519);
and U300 (N_300,N_88,In_665);
and U301 (N_301,N_58,N_151);
nor U302 (N_302,N_170,In_709);
nand U303 (N_303,In_701,N_73);
xor U304 (N_304,N_176,N_198);
nor U305 (N_305,In_296,N_160);
nor U306 (N_306,N_94,In_282);
or U307 (N_307,In_386,In_606);
nor U308 (N_308,N_12,In_566);
nor U309 (N_309,In_428,In_337);
and U310 (N_310,N_87,N_70);
and U311 (N_311,N_13,In_490);
nor U312 (N_312,N_34,N_100);
or U313 (N_313,In_13,In_451);
or U314 (N_314,In_88,In_576);
or U315 (N_315,N_138,N_129);
nand U316 (N_316,In_744,N_21);
nor U317 (N_317,In_90,N_83);
or U318 (N_318,In_513,In_407);
nand U319 (N_319,In_721,N_125);
nor U320 (N_320,N_79,In_346);
nor U321 (N_321,N_136,In_104);
nand U322 (N_322,In_293,In_156);
nor U323 (N_323,N_192,In_98);
nor U324 (N_324,In_493,In_577);
nor U325 (N_325,In_739,In_722);
and U326 (N_326,In_159,N_6);
nor U327 (N_327,In_318,N_92);
nand U328 (N_328,In_516,In_61);
nand U329 (N_329,N_172,N_89);
nand U330 (N_330,N_193,In_487);
or U331 (N_331,In_724,N_42);
nand U332 (N_332,In_417,In_24);
nand U333 (N_333,In_532,N_84);
or U334 (N_334,In_528,N_124);
nor U335 (N_335,N_158,In_506);
and U336 (N_336,In_117,In_677);
and U337 (N_337,N_2,In_641);
nand U338 (N_338,N_5,In_65);
nor U339 (N_339,N_15,N_61);
and U340 (N_340,N_197,N_69);
and U341 (N_341,N_74,In_736);
and U342 (N_342,N_143,In_662);
and U343 (N_343,N_3,In_444);
nor U344 (N_344,In_124,In_705);
or U345 (N_345,In_554,In_406);
or U346 (N_346,In_59,In_418);
nor U347 (N_347,In_359,In_306);
and U348 (N_348,In_498,N_112);
and U349 (N_349,In_383,In_673);
or U350 (N_350,In_58,In_668);
or U351 (N_351,In_585,N_33);
or U352 (N_352,In_9,In_394);
nand U353 (N_353,In_330,N_153);
nor U354 (N_354,In_221,N_0);
nand U355 (N_355,N_78,In_501);
nor U356 (N_356,N_10,In_146);
or U357 (N_357,In_269,In_453);
or U358 (N_358,In_728,In_281);
nor U359 (N_359,In_499,In_180);
nand U360 (N_360,In_465,In_607);
nand U361 (N_361,In_248,In_445);
nor U362 (N_362,In_99,In_85);
and U363 (N_363,N_130,N_26);
or U364 (N_364,In_437,In_96);
and U365 (N_365,In_485,N_9);
nand U366 (N_366,In_203,N_7);
and U367 (N_367,N_145,In_389);
nand U368 (N_368,In_70,N_109);
and U369 (N_369,In_127,N_121);
nand U370 (N_370,In_7,In_711);
and U371 (N_371,In_28,In_15);
nor U372 (N_372,N_48,In_719);
and U373 (N_373,N_184,In_369);
and U374 (N_374,In_508,In_447);
nor U375 (N_375,In_40,In_526);
or U376 (N_376,N_116,In_168);
xnor U377 (N_377,N_156,N_187);
or U378 (N_378,In_626,N_31);
and U379 (N_379,N_123,In_309);
or U380 (N_380,N_90,In_397);
or U381 (N_381,N_103,In_648);
nor U382 (N_382,N_107,N_111);
nor U383 (N_383,In_700,In_538);
or U384 (N_384,In_450,In_227);
nor U385 (N_385,In_518,In_511);
nand U386 (N_386,In_419,N_177);
nor U387 (N_387,N_152,N_140);
or U388 (N_388,In_192,In_460);
nor U389 (N_389,N_39,In_438);
nor U390 (N_390,N_196,In_145);
and U391 (N_391,N_115,In_726);
nor U392 (N_392,In_5,In_35);
nand U393 (N_393,In_578,N_98);
nand U394 (N_394,In_166,N_194);
nor U395 (N_395,In_201,In_279);
nor U396 (N_396,In_486,In_674);
nand U397 (N_397,In_19,In_128);
and U398 (N_398,N_45,N_43);
and U399 (N_399,N_114,In_588);
and U400 (N_400,N_236,In_185);
nand U401 (N_401,N_330,N_290);
nor U402 (N_402,N_303,N_242);
and U403 (N_403,In_76,N_85);
nand U404 (N_404,N_150,N_296);
and U405 (N_405,N_333,N_212);
nand U406 (N_406,N_350,N_36);
and U407 (N_407,In_301,N_317);
or U408 (N_408,N_387,N_274);
or U409 (N_409,In_385,N_241);
nand U410 (N_410,N_294,N_268);
or U411 (N_411,In_167,In_352);
nand U412 (N_412,N_373,N_253);
nand U413 (N_413,In_338,N_270);
nand U414 (N_414,N_249,In_455);
or U415 (N_415,N_154,In_713);
nand U416 (N_416,In_303,N_244);
and U417 (N_417,N_319,N_131);
nand U418 (N_418,N_336,N_298);
and U419 (N_419,N_375,In_432);
nand U420 (N_420,N_366,N_291);
nand U421 (N_421,N_306,N_246);
and U422 (N_422,In_633,N_222);
nor U423 (N_423,N_75,In_139);
and U424 (N_424,N_157,In_560);
nor U425 (N_425,N_390,N_232);
or U426 (N_426,N_382,In_323);
nand U427 (N_427,In_689,N_262);
or U428 (N_428,In_264,N_230);
nor U429 (N_429,N_214,In_497);
or U430 (N_430,In_136,In_198);
nor U431 (N_431,N_349,N_81);
and U432 (N_432,N_149,N_210);
nand U433 (N_433,In_525,N_248);
xnor U434 (N_434,N_269,In_612);
nand U435 (N_435,N_346,N_331);
or U436 (N_436,N_313,In_153);
nand U437 (N_437,In_663,N_367);
nand U438 (N_438,N_135,N_50);
nor U439 (N_439,N_280,In_429);
or U440 (N_440,N_240,N_254);
and U441 (N_441,N_328,N_14);
xor U442 (N_442,In_350,N_163);
and U443 (N_443,N_368,N_216);
nand U444 (N_444,N_166,N_80);
and U445 (N_445,In_392,N_233);
nand U446 (N_446,N_28,In_669);
and U447 (N_447,N_231,In_551);
nor U448 (N_448,In_218,N_206);
and U449 (N_449,N_378,In_52);
or U450 (N_450,N_318,In_623);
nor U451 (N_451,N_320,N_361);
nand U452 (N_452,N_219,N_392);
nand U453 (N_453,In_580,N_341);
nand U454 (N_454,In_172,In_54);
xnor U455 (N_455,N_22,In_405);
nand U456 (N_456,In_86,In_200);
and U457 (N_457,N_76,N_372);
nor U458 (N_458,N_394,In_597);
nor U459 (N_459,N_203,N_220);
nand U460 (N_460,N_63,In_749);
nor U461 (N_461,N_374,N_327);
and U462 (N_462,N_243,N_257);
or U463 (N_463,In_46,N_363);
or U464 (N_464,In_193,N_381);
or U465 (N_465,N_369,In_702);
nand U466 (N_466,N_189,N_324);
and U467 (N_467,N_273,In_121);
and U468 (N_468,N_279,N_263);
and U469 (N_469,In_115,In_152);
or U470 (N_470,N_379,N_57);
nor U471 (N_471,In_80,In_697);
nor U472 (N_472,N_395,N_218);
and U473 (N_473,N_179,N_340);
or U474 (N_474,N_229,N_261);
or U475 (N_475,N_302,N_234);
nand U476 (N_476,N_223,In_141);
nor U477 (N_477,In_239,In_731);
nor U478 (N_478,N_310,N_332);
nor U479 (N_479,N_164,N_282);
nor U480 (N_480,In_273,In_587);
nand U481 (N_481,N_278,N_380);
xnor U482 (N_482,In_132,N_4);
nand U483 (N_483,N_384,N_342);
xor U484 (N_484,N_284,N_245);
and U485 (N_485,N_299,N_347);
nor U486 (N_486,In_379,In_592);
nand U487 (N_487,N_383,N_202);
or U488 (N_488,In_109,N_386);
nor U489 (N_489,N_101,N_49);
nor U490 (N_490,N_24,In_599);
nor U491 (N_491,N_370,N_204);
nand U492 (N_492,N_224,N_295);
xnor U493 (N_493,N_51,In_250);
and U494 (N_494,N_235,N_67);
nor U495 (N_495,N_283,N_276);
nor U496 (N_496,N_275,In_575);
nor U497 (N_497,In_143,N_64);
or U498 (N_498,N_399,N_205);
or U499 (N_499,N_272,N_334);
nand U500 (N_500,N_285,In_720);
and U501 (N_501,N_264,In_400);
or U502 (N_502,In_140,N_72);
and U503 (N_503,N_377,N_127);
nor U504 (N_504,N_326,N_364);
nor U505 (N_505,In_661,In_272);
nor U506 (N_506,N_389,In_252);
and U507 (N_507,N_18,N_25);
or U508 (N_508,In_474,In_408);
nor U509 (N_509,N_316,N_260);
nor U510 (N_510,N_180,N_238);
or U511 (N_511,N_356,N_348);
or U512 (N_512,N_255,N_337);
xor U513 (N_513,In_276,N_397);
or U514 (N_514,N_208,N_201);
and U515 (N_515,N_388,N_267);
or U516 (N_516,N_371,N_105);
or U517 (N_517,N_314,In_130);
and U518 (N_518,N_225,In_605);
and U519 (N_519,N_178,In_492);
nand U520 (N_520,In_163,N_343);
nor U521 (N_521,N_271,N_281);
or U522 (N_522,In_298,N_174);
nand U523 (N_523,In_165,N_385);
nand U524 (N_524,In_482,N_288);
nand U525 (N_525,N_239,N_250);
nand U526 (N_526,N_353,N_358);
nor U527 (N_527,N_221,N_122);
or U528 (N_528,N_265,N_300);
and U529 (N_529,N_323,N_292);
or U530 (N_530,N_362,N_396);
and U531 (N_531,N_322,N_247);
nand U532 (N_532,N_258,N_53);
nand U533 (N_533,N_141,N_308);
nand U534 (N_534,N_365,N_312);
nor U535 (N_535,In_639,N_211);
nor U536 (N_536,N_91,N_311);
nand U537 (N_537,N_251,In_122);
and U538 (N_538,In_341,In_179);
nand U539 (N_539,N_315,In_66);
nand U540 (N_540,N_309,N_106);
nor U541 (N_541,In_42,N_297);
and U542 (N_542,N_391,N_289);
and U543 (N_543,N_321,N_354);
and U544 (N_544,N_32,N_325);
and U545 (N_545,In_738,N_228);
or U546 (N_546,N_213,N_252);
and U547 (N_547,N_355,N_339);
nand U548 (N_548,N_256,N_30);
and U549 (N_549,N_335,In_349);
and U550 (N_550,In_317,N_307);
nor U551 (N_551,N_113,N_217);
nor U552 (N_552,N_352,N_186);
nor U553 (N_553,N_259,N_237);
and U554 (N_554,N_338,N_301);
nand U555 (N_555,In_325,N_304);
nor U556 (N_556,N_376,N_344);
or U557 (N_557,N_11,N_393);
or U558 (N_558,N_20,In_358);
and U559 (N_559,N_359,In_190);
nand U560 (N_560,N_398,In_129);
or U561 (N_561,N_108,In_572);
and U562 (N_562,N_227,N_200);
xor U563 (N_563,N_329,In_496);
and U564 (N_564,N_357,N_345);
nand U565 (N_565,N_209,N_305);
or U566 (N_566,N_351,N_17);
or U567 (N_567,N_132,N_286);
nand U568 (N_568,N_287,N_277);
nand U569 (N_569,In_93,N_119);
nand U570 (N_570,N_190,N_293);
nor U571 (N_571,In_594,N_266);
or U572 (N_572,N_159,N_38);
nor U573 (N_573,N_360,N_207);
and U574 (N_574,N_226,N_215);
nand U575 (N_575,In_597,N_72);
nor U576 (N_576,N_324,In_352);
and U577 (N_577,N_272,N_222);
or U578 (N_578,N_282,N_302);
nand U579 (N_579,In_200,N_359);
or U580 (N_580,N_326,N_294);
nand U581 (N_581,In_663,N_223);
nor U582 (N_582,N_127,N_219);
and U583 (N_583,N_246,N_239);
and U584 (N_584,In_140,N_76);
nor U585 (N_585,In_76,In_93);
nor U586 (N_586,N_331,N_297);
nand U587 (N_587,N_233,In_633);
and U588 (N_588,N_127,N_201);
nand U589 (N_589,In_385,N_32);
or U590 (N_590,In_109,N_255);
nand U591 (N_591,N_289,N_248);
or U592 (N_592,In_153,N_201);
or U593 (N_593,N_351,N_32);
or U594 (N_594,N_30,N_235);
or U595 (N_595,N_245,N_349);
nor U596 (N_596,N_127,N_352);
or U597 (N_597,N_245,N_274);
nor U598 (N_598,N_204,In_551);
nor U599 (N_599,In_633,In_301);
nor U600 (N_600,N_492,N_595);
nor U601 (N_601,N_583,N_593);
nor U602 (N_602,N_424,N_457);
nand U603 (N_603,N_517,N_568);
nand U604 (N_604,N_502,N_431);
and U605 (N_605,N_495,N_529);
and U606 (N_606,N_499,N_464);
and U607 (N_607,N_539,N_591);
and U608 (N_608,N_441,N_423);
or U609 (N_609,N_460,N_475);
nand U610 (N_610,N_404,N_552);
and U611 (N_611,N_479,N_514);
and U612 (N_612,N_481,N_439);
nor U613 (N_613,N_581,N_544);
nand U614 (N_614,N_503,N_512);
and U615 (N_615,N_509,N_508);
or U616 (N_616,N_419,N_445);
nor U617 (N_617,N_594,N_532);
nor U618 (N_618,N_426,N_561);
nor U619 (N_619,N_483,N_435);
and U620 (N_620,N_578,N_537);
or U621 (N_621,N_418,N_449);
nor U622 (N_622,N_430,N_577);
and U623 (N_623,N_564,N_559);
or U624 (N_624,N_500,N_478);
and U625 (N_625,N_513,N_553);
nor U626 (N_626,N_573,N_429);
or U627 (N_627,N_543,N_451);
nor U628 (N_628,N_538,N_540);
nor U629 (N_629,N_473,N_422);
nand U630 (N_630,N_554,N_472);
nand U631 (N_631,N_549,N_470);
nand U632 (N_632,N_516,N_410);
or U633 (N_633,N_491,N_582);
nand U634 (N_634,N_504,N_597);
and U635 (N_635,N_528,N_530);
and U636 (N_636,N_574,N_586);
or U637 (N_637,N_520,N_412);
and U638 (N_638,N_444,N_531);
nor U639 (N_639,N_471,N_468);
and U640 (N_640,N_456,N_527);
nand U641 (N_641,N_521,N_407);
or U642 (N_642,N_488,N_400);
nor U643 (N_643,N_534,N_421);
nor U644 (N_644,N_555,N_585);
nor U645 (N_645,N_415,N_526);
and U646 (N_646,N_482,N_570);
nor U647 (N_647,N_571,N_416);
and U648 (N_648,N_519,N_566);
nand U649 (N_649,N_589,N_401);
and U650 (N_650,N_598,N_545);
nor U651 (N_651,N_427,N_515);
nor U652 (N_652,N_498,N_408);
nand U653 (N_653,N_434,N_556);
nor U654 (N_654,N_563,N_494);
nor U655 (N_655,N_487,N_425);
nand U656 (N_656,N_465,N_541);
and U657 (N_657,N_480,N_442);
nand U658 (N_658,N_546,N_522);
nand U659 (N_659,N_402,N_575);
nor U660 (N_660,N_560,N_474);
xor U661 (N_661,N_413,N_428);
xor U662 (N_662,N_588,N_524);
and U663 (N_663,N_443,N_458);
or U664 (N_664,N_459,N_551);
and U665 (N_665,N_525,N_596);
nand U666 (N_666,N_463,N_414);
nand U667 (N_667,N_490,N_505);
or U668 (N_668,N_448,N_572);
and U669 (N_669,N_417,N_511);
nand U670 (N_670,N_587,N_432);
and U671 (N_671,N_462,N_405);
nand U672 (N_672,N_550,N_523);
and U673 (N_673,N_501,N_453);
and U674 (N_674,N_562,N_454);
nand U675 (N_675,N_599,N_584);
nand U676 (N_676,N_510,N_455);
and U677 (N_677,N_438,N_558);
nor U678 (N_678,N_469,N_446);
nor U679 (N_679,N_411,N_440);
xor U680 (N_680,N_485,N_518);
nor U681 (N_681,N_437,N_409);
or U682 (N_682,N_576,N_420);
nand U683 (N_683,N_497,N_542);
and U684 (N_684,N_436,N_580);
nand U685 (N_685,N_447,N_493);
and U686 (N_686,N_496,N_567);
nand U687 (N_687,N_507,N_403);
nor U688 (N_688,N_450,N_579);
nor U689 (N_689,N_476,N_533);
nor U690 (N_690,N_557,N_467);
nand U691 (N_691,N_565,N_484);
nor U692 (N_692,N_406,N_535);
and U693 (N_693,N_592,N_466);
nand U694 (N_694,N_461,N_452);
nand U695 (N_695,N_548,N_569);
nand U696 (N_696,N_536,N_506);
nand U697 (N_697,N_590,N_486);
or U698 (N_698,N_477,N_547);
or U699 (N_699,N_433,N_489);
and U700 (N_700,N_584,N_506);
and U701 (N_701,N_518,N_455);
nor U702 (N_702,N_562,N_456);
nand U703 (N_703,N_595,N_457);
or U704 (N_704,N_442,N_593);
and U705 (N_705,N_427,N_497);
nand U706 (N_706,N_437,N_572);
nor U707 (N_707,N_579,N_433);
nor U708 (N_708,N_563,N_545);
nand U709 (N_709,N_593,N_490);
and U710 (N_710,N_421,N_452);
or U711 (N_711,N_580,N_505);
and U712 (N_712,N_522,N_467);
nand U713 (N_713,N_473,N_543);
nor U714 (N_714,N_585,N_441);
or U715 (N_715,N_401,N_414);
nand U716 (N_716,N_408,N_447);
nor U717 (N_717,N_575,N_595);
and U718 (N_718,N_405,N_568);
or U719 (N_719,N_471,N_532);
and U720 (N_720,N_527,N_403);
and U721 (N_721,N_454,N_574);
nand U722 (N_722,N_451,N_500);
and U723 (N_723,N_570,N_558);
nor U724 (N_724,N_449,N_551);
and U725 (N_725,N_504,N_513);
nor U726 (N_726,N_432,N_522);
nor U727 (N_727,N_464,N_420);
or U728 (N_728,N_596,N_412);
and U729 (N_729,N_487,N_585);
and U730 (N_730,N_430,N_457);
nor U731 (N_731,N_406,N_426);
nor U732 (N_732,N_424,N_578);
nand U733 (N_733,N_441,N_430);
or U734 (N_734,N_443,N_459);
and U735 (N_735,N_411,N_425);
xor U736 (N_736,N_573,N_419);
nor U737 (N_737,N_526,N_523);
and U738 (N_738,N_591,N_445);
and U739 (N_739,N_589,N_538);
nor U740 (N_740,N_499,N_506);
nor U741 (N_741,N_402,N_435);
or U742 (N_742,N_598,N_463);
and U743 (N_743,N_438,N_429);
or U744 (N_744,N_582,N_408);
nand U745 (N_745,N_453,N_597);
nand U746 (N_746,N_432,N_553);
or U747 (N_747,N_564,N_558);
or U748 (N_748,N_498,N_467);
nand U749 (N_749,N_459,N_540);
and U750 (N_750,N_543,N_502);
nand U751 (N_751,N_499,N_587);
nor U752 (N_752,N_424,N_413);
nand U753 (N_753,N_413,N_544);
nor U754 (N_754,N_557,N_410);
and U755 (N_755,N_442,N_521);
and U756 (N_756,N_486,N_457);
nand U757 (N_757,N_554,N_412);
nand U758 (N_758,N_541,N_451);
nand U759 (N_759,N_565,N_594);
nor U760 (N_760,N_406,N_448);
or U761 (N_761,N_551,N_405);
and U762 (N_762,N_547,N_418);
or U763 (N_763,N_557,N_480);
nor U764 (N_764,N_442,N_580);
nor U765 (N_765,N_535,N_598);
or U766 (N_766,N_438,N_539);
nor U767 (N_767,N_468,N_486);
nor U768 (N_768,N_574,N_542);
nor U769 (N_769,N_492,N_501);
or U770 (N_770,N_557,N_594);
and U771 (N_771,N_547,N_567);
nand U772 (N_772,N_578,N_493);
nand U773 (N_773,N_523,N_558);
or U774 (N_774,N_503,N_539);
nor U775 (N_775,N_476,N_420);
nand U776 (N_776,N_488,N_462);
and U777 (N_777,N_489,N_450);
nor U778 (N_778,N_474,N_545);
and U779 (N_779,N_425,N_453);
nor U780 (N_780,N_472,N_423);
nor U781 (N_781,N_431,N_467);
nor U782 (N_782,N_573,N_538);
nand U783 (N_783,N_497,N_441);
and U784 (N_784,N_549,N_533);
nand U785 (N_785,N_566,N_584);
nor U786 (N_786,N_457,N_518);
nor U787 (N_787,N_588,N_502);
and U788 (N_788,N_565,N_530);
nand U789 (N_789,N_490,N_521);
or U790 (N_790,N_497,N_540);
nor U791 (N_791,N_593,N_559);
and U792 (N_792,N_497,N_400);
and U793 (N_793,N_561,N_568);
and U794 (N_794,N_528,N_428);
and U795 (N_795,N_444,N_450);
nand U796 (N_796,N_576,N_464);
nand U797 (N_797,N_545,N_498);
and U798 (N_798,N_558,N_559);
nor U799 (N_799,N_580,N_445);
xnor U800 (N_800,N_689,N_766);
nor U801 (N_801,N_710,N_738);
nand U802 (N_802,N_761,N_757);
nor U803 (N_803,N_643,N_702);
nor U804 (N_804,N_603,N_637);
or U805 (N_805,N_795,N_722);
or U806 (N_806,N_748,N_638);
or U807 (N_807,N_786,N_790);
nor U808 (N_808,N_633,N_762);
and U809 (N_809,N_657,N_724);
and U810 (N_810,N_734,N_779);
or U811 (N_811,N_628,N_687);
nor U812 (N_812,N_613,N_784);
nand U813 (N_813,N_769,N_707);
or U814 (N_814,N_640,N_673);
nand U815 (N_815,N_614,N_726);
and U816 (N_816,N_659,N_601);
nand U817 (N_817,N_745,N_768);
and U818 (N_818,N_703,N_732);
and U819 (N_819,N_743,N_654);
nor U820 (N_820,N_604,N_605);
nor U821 (N_821,N_616,N_792);
nand U822 (N_822,N_778,N_629);
nor U823 (N_823,N_789,N_758);
nand U824 (N_824,N_671,N_693);
nand U825 (N_825,N_797,N_642);
and U826 (N_826,N_684,N_680);
nand U827 (N_827,N_735,N_721);
and U828 (N_828,N_696,N_699);
or U829 (N_829,N_728,N_796);
nor U830 (N_830,N_641,N_647);
nand U831 (N_831,N_685,N_754);
nand U832 (N_832,N_669,N_717);
nand U833 (N_833,N_697,N_660);
or U834 (N_834,N_747,N_715);
or U835 (N_835,N_645,N_737);
nor U836 (N_836,N_794,N_709);
nor U837 (N_837,N_764,N_644);
or U838 (N_838,N_705,N_617);
nor U839 (N_839,N_700,N_675);
nand U840 (N_840,N_690,N_706);
or U841 (N_841,N_608,N_676);
nand U842 (N_842,N_656,N_625);
and U843 (N_843,N_630,N_719);
nor U844 (N_844,N_623,N_772);
and U845 (N_845,N_632,N_677);
or U846 (N_846,N_730,N_672);
nand U847 (N_847,N_631,N_782);
nor U848 (N_848,N_612,N_752);
nor U849 (N_849,N_636,N_740);
nor U850 (N_850,N_718,N_733);
or U851 (N_851,N_799,N_686);
nand U852 (N_852,N_650,N_666);
and U853 (N_853,N_777,N_716);
or U854 (N_854,N_714,N_727);
nand U855 (N_855,N_793,N_746);
nor U856 (N_856,N_661,N_663);
nand U857 (N_857,N_635,N_621);
and U858 (N_858,N_664,N_736);
and U859 (N_859,N_634,N_725);
nand U860 (N_860,N_607,N_620);
or U861 (N_861,N_627,N_610);
xnor U862 (N_862,N_655,N_711);
and U863 (N_863,N_611,N_651);
and U864 (N_864,N_708,N_723);
nand U865 (N_865,N_798,N_759);
nand U866 (N_866,N_649,N_704);
or U867 (N_867,N_668,N_618);
xor U868 (N_868,N_713,N_701);
nor U869 (N_869,N_776,N_658);
nand U870 (N_870,N_788,N_750);
nor U871 (N_871,N_683,N_744);
or U872 (N_872,N_681,N_760);
and U873 (N_873,N_780,N_646);
nand U874 (N_874,N_694,N_606);
or U875 (N_875,N_662,N_648);
and U876 (N_876,N_787,N_753);
or U877 (N_877,N_691,N_653);
and U878 (N_878,N_609,N_791);
or U879 (N_879,N_674,N_729);
nand U880 (N_880,N_742,N_783);
or U881 (N_881,N_781,N_755);
and U882 (N_882,N_767,N_667);
nand U883 (N_883,N_698,N_773);
or U884 (N_884,N_626,N_775);
nand U885 (N_885,N_652,N_749);
xor U886 (N_886,N_756,N_751);
nor U887 (N_887,N_771,N_619);
nand U888 (N_888,N_739,N_731);
nand U889 (N_889,N_765,N_602);
and U890 (N_890,N_639,N_682);
or U891 (N_891,N_678,N_670);
or U892 (N_892,N_665,N_785);
and U893 (N_893,N_741,N_615);
and U894 (N_894,N_695,N_712);
or U895 (N_895,N_774,N_720);
or U896 (N_896,N_600,N_692);
and U897 (N_897,N_679,N_763);
nor U898 (N_898,N_624,N_688);
nand U899 (N_899,N_770,N_622);
xnor U900 (N_900,N_687,N_618);
nand U901 (N_901,N_666,N_667);
and U902 (N_902,N_615,N_705);
and U903 (N_903,N_751,N_608);
nand U904 (N_904,N_708,N_668);
and U905 (N_905,N_603,N_616);
and U906 (N_906,N_761,N_600);
nand U907 (N_907,N_792,N_692);
and U908 (N_908,N_639,N_754);
nand U909 (N_909,N_756,N_606);
and U910 (N_910,N_612,N_736);
nand U911 (N_911,N_747,N_721);
or U912 (N_912,N_693,N_603);
or U913 (N_913,N_744,N_696);
nand U914 (N_914,N_624,N_623);
nor U915 (N_915,N_666,N_790);
nor U916 (N_916,N_710,N_697);
nand U917 (N_917,N_624,N_714);
nor U918 (N_918,N_691,N_629);
nor U919 (N_919,N_748,N_790);
nand U920 (N_920,N_717,N_657);
nor U921 (N_921,N_619,N_683);
or U922 (N_922,N_622,N_612);
nand U923 (N_923,N_619,N_754);
and U924 (N_924,N_705,N_612);
nand U925 (N_925,N_742,N_745);
nand U926 (N_926,N_756,N_665);
or U927 (N_927,N_707,N_798);
or U928 (N_928,N_658,N_687);
nor U929 (N_929,N_705,N_704);
or U930 (N_930,N_697,N_617);
and U931 (N_931,N_786,N_739);
nor U932 (N_932,N_753,N_783);
and U933 (N_933,N_712,N_699);
and U934 (N_934,N_687,N_728);
xnor U935 (N_935,N_783,N_709);
nand U936 (N_936,N_758,N_750);
nor U937 (N_937,N_604,N_732);
nand U938 (N_938,N_794,N_643);
and U939 (N_939,N_708,N_612);
and U940 (N_940,N_615,N_787);
nor U941 (N_941,N_626,N_728);
nand U942 (N_942,N_674,N_642);
nor U943 (N_943,N_707,N_607);
nor U944 (N_944,N_610,N_799);
nor U945 (N_945,N_789,N_648);
nor U946 (N_946,N_601,N_751);
or U947 (N_947,N_741,N_799);
nor U948 (N_948,N_644,N_602);
and U949 (N_949,N_737,N_655);
or U950 (N_950,N_744,N_707);
nand U951 (N_951,N_704,N_647);
nor U952 (N_952,N_685,N_708);
nor U953 (N_953,N_785,N_681);
and U954 (N_954,N_799,N_771);
nand U955 (N_955,N_713,N_602);
nand U956 (N_956,N_726,N_626);
nand U957 (N_957,N_747,N_668);
or U958 (N_958,N_674,N_797);
and U959 (N_959,N_788,N_714);
and U960 (N_960,N_601,N_607);
and U961 (N_961,N_650,N_762);
nor U962 (N_962,N_761,N_639);
nand U963 (N_963,N_705,N_752);
and U964 (N_964,N_662,N_799);
or U965 (N_965,N_609,N_634);
or U966 (N_966,N_653,N_742);
or U967 (N_967,N_610,N_743);
or U968 (N_968,N_790,N_632);
or U969 (N_969,N_680,N_739);
nor U970 (N_970,N_625,N_781);
or U971 (N_971,N_789,N_615);
nor U972 (N_972,N_703,N_625);
nor U973 (N_973,N_610,N_722);
and U974 (N_974,N_687,N_644);
nor U975 (N_975,N_645,N_695);
nand U976 (N_976,N_644,N_709);
nor U977 (N_977,N_613,N_789);
or U978 (N_978,N_739,N_665);
nand U979 (N_979,N_645,N_697);
or U980 (N_980,N_660,N_699);
xor U981 (N_981,N_784,N_696);
or U982 (N_982,N_679,N_768);
nor U983 (N_983,N_775,N_799);
nor U984 (N_984,N_672,N_652);
nand U985 (N_985,N_703,N_609);
or U986 (N_986,N_771,N_774);
and U987 (N_987,N_717,N_645);
nor U988 (N_988,N_628,N_736);
or U989 (N_989,N_733,N_767);
and U990 (N_990,N_638,N_774);
or U991 (N_991,N_749,N_708);
or U992 (N_992,N_602,N_637);
or U993 (N_993,N_715,N_798);
or U994 (N_994,N_672,N_760);
nor U995 (N_995,N_679,N_747);
nor U996 (N_996,N_687,N_748);
nor U997 (N_997,N_657,N_629);
or U998 (N_998,N_666,N_700);
nand U999 (N_999,N_796,N_676);
and U1000 (N_1000,N_892,N_970);
or U1001 (N_1001,N_925,N_999);
nand U1002 (N_1002,N_957,N_898);
and U1003 (N_1003,N_845,N_886);
nand U1004 (N_1004,N_917,N_848);
nand U1005 (N_1005,N_894,N_987);
nand U1006 (N_1006,N_828,N_947);
nand U1007 (N_1007,N_988,N_901);
xnor U1008 (N_1008,N_928,N_882);
or U1009 (N_1009,N_971,N_893);
and U1010 (N_1010,N_939,N_823);
or U1011 (N_1011,N_962,N_857);
nand U1012 (N_1012,N_909,N_833);
nand U1013 (N_1013,N_883,N_844);
nand U1014 (N_1014,N_896,N_940);
or U1015 (N_1015,N_946,N_801);
and U1016 (N_1016,N_881,N_887);
nor U1017 (N_1017,N_888,N_919);
or U1018 (N_1018,N_908,N_968);
or U1019 (N_1019,N_934,N_854);
and U1020 (N_1020,N_842,N_983);
and U1021 (N_1021,N_964,N_984);
or U1022 (N_1022,N_953,N_829);
nor U1023 (N_1023,N_834,N_976);
or U1024 (N_1024,N_849,N_921);
or U1025 (N_1025,N_932,N_808);
nor U1026 (N_1026,N_821,N_958);
nor U1027 (N_1027,N_814,N_811);
nor U1028 (N_1028,N_944,N_911);
nor U1029 (N_1029,N_914,N_998);
nor U1030 (N_1030,N_897,N_993);
nor U1031 (N_1031,N_884,N_871);
nor U1032 (N_1032,N_920,N_948);
or U1033 (N_1033,N_954,N_870);
and U1034 (N_1034,N_863,N_855);
nand U1035 (N_1035,N_975,N_858);
or U1036 (N_1036,N_942,N_803);
nand U1037 (N_1037,N_860,N_843);
and U1038 (N_1038,N_874,N_837);
nor U1039 (N_1039,N_873,N_906);
nand U1040 (N_1040,N_869,N_916);
nand U1041 (N_1041,N_952,N_885);
and U1042 (N_1042,N_889,N_856);
or U1043 (N_1043,N_997,N_903);
nand U1044 (N_1044,N_972,N_912);
nand U1045 (N_1045,N_937,N_991);
nor U1046 (N_1046,N_876,N_836);
or U1047 (N_1047,N_847,N_959);
nor U1048 (N_1048,N_986,N_977);
nand U1049 (N_1049,N_899,N_929);
nor U1050 (N_1050,N_852,N_840);
nor U1051 (N_1051,N_965,N_868);
and U1052 (N_1052,N_864,N_985);
and U1053 (N_1053,N_802,N_902);
nor U1054 (N_1054,N_861,N_825);
xnor U1055 (N_1055,N_973,N_807);
and U1056 (N_1056,N_865,N_996);
or U1057 (N_1057,N_880,N_877);
and U1058 (N_1058,N_812,N_831);
nor U1059 (N_1059,N_878,N_820);
or U1060 (N_1060,N_879,N_941);
or U1061 (N_1061,N_804,N_931);
nor U1062 (N_1062,N_950,N_980);
or U1063 (N_1063,N_978,N_872);
nor U1064 (N_1064,N_859,N_936);
nor U1065 (N_1065,N_918,N_943);
and U1066 (N_1066,N_891,N_815);
or U1067 (N_1067,N_813,N_994);
nor U1068 (N_1068,N_810,N_955);
and U1069 (N_1069,N_851,N_819);
nand U1070 (N_1070,N_995,N_966);
and U1071 (N_1071,N_949,N_830);
nand U1072 (N_1072,N_924,N_905);
or U1073 (N_1073,N_930,N_963);
and U1074 (N_1074,N_956,N_907);
nor U1075 (N_1075,N_800,N_895);
nor U1076 (N_1076,N_826,N_816);
and U1077 (N_1077,N_989,N_926);
and U1078 (N_1078,N_822,N_866);
or U1079 (N_1079,N_846,N_945);
and U1080 (N_1080,N_967,N_990);
or U1081 (N_1081,N_951,N_969);
nand U1082 (N_1082,N_862,N_805);
or U1083 (N_1083,N_961,N_817);
nand U1084 (N_1084,N_850,N_938);
and U1085 (N_1085,N_933,N_981);
or U1086 (N_1086,N_979,N_853);
or U1087 (N_1087,N_935,N_904);
or U1088 (N_1088,N_922,N_835);
nor U1089 (N_1089,N_910,N_839);
xor U1090 (N_1090,N_832,N_992);
nor U1091 (N_1091,N_827,N_982);
or U1092 (N_1092,N_875,N_809);
or U1093 (N_1093,N_824,N_900);
or U1094 (N_1094,N_867,N_841);
nand U1095 (N_1095,N_818,N_915);
and U1096 (N_1096,N_838,N_806);
and U1097 (N_1097,N_960,N_890);
and U1098 (N_1098,N_923,N_913);
or U1099 (N_1099,N_974,N_927);
or U1100 (N_1100,N_880,N_967);
nand U1101 (N_1101,N_939,N_875);
or U1102 (N_1102,N_916,N_934);
nand U1103 (N_1103,N_920,N_999);
nor U1104 (N_1104,N_997,N_973);
nor U1105 (N_1105,N_952,N_881);
nand U1106 (N_1106,N_869,N_832);
nand U1107 (N_1107,N_963,N_995);
nor U1108 (N_1108,N_929,N_907);
nand U1109 (N_1109,N_941,N_957);
nand U1110 (N_1110,N_810,N_801);
or U1111 (N_1111,N_861,N_800);
nor U1112 (N_1112,N_822,N_975);
or U1113 (N_1113,N_897,N_821);
nand U1114 (N_1114,N_803,N_825);
and U1115 (N_1115,N_802,N_812);
or U1116 (N_1116,N_995,N_815);
nand U1117 (N_1117,N_984,N_847);
nor U1118 (N_1118,N_955,N_990);
or U1119 (N_1119,N_878,N_945);
nor U1120 (N_1120,N_867,N_921);
and U1121 (N_1121,N_853,N_873);
or U1122 (N_1122,N_978,N_992);
and U1123 (N_1123,N_995,N_867);
nor U1124 (N_1124,N_898,N_986);
nor U1125 (N_1125,N_881,N_843);
nor U1126 (N_1126,N_847,N_857);
or U1127 (N_1127,N_857,N_939);
xor U1128 (N_1128,N_963,N_928);
nor U1129 (N_1129,N_885,N_850);
nand U1130 (N_1130,N_874,N_961);
nand U1131 (N_1131,N_807,N_848);
nor U1132 (N_1132,N_886,N_873);
and U1133 (N_1133,N_862,N_807);
nand U1134 (N_1134,N_918,N_939);
nand U1135 (N_1135,N_838,N_970);
and U1136 (N_1136,N_966,N_821);
and U1137 (N_1137,N_849,N_876);
nand U1138 (N_1138,N_914,N_992);
nor U1139 (N_1139,N_807,N_880);
nand U1140 (N_1140,N_890,N_874);
or U1141 (N_1141,N_917,N_888);
nand U1142 (N_1142,N_941,N_835);
and U1143 (N_1143,N_937,N_958);
nor U1144 (N_1144,N_908,N_860);
or U1145 (N_1145,N_810,N_808);
and U1146 (N_1146,N_838,N_974);
and U1147 (N_1147,N_802,N_928);
nor U1148 (N_1148,N_888,N_867);
nor U1149 (N_1149,N_883,N_965);
or U1150 (N_1150,N_888,N_845);
or U1151 (N_1151,N_970,N_853);
nand U1152 (N_1152,N_861,N_889);
nor U1153 (N_1153,N_871,N_802);
and U1154 (N_1154,N_880,N_879);
and U1155 (N_1155,N_950,N_959);
and U1156 (N_1156,N_957,N_944);
nand U1157 (N_1157,N_966,N_864);
nor U1158 (N_1158,N_855,N_985);
nand U1159 (N_1159,N_807,N_967);
nor U1160 (N_1160,N_883,N_986);
nand U1161 (N_1161,N_861,N_826);
nor U1162 (N_1162,N_950,N_832);
or U1163 (N_1163,N_896,N_866);
or U1164 (N_1164,N_989,N_879);
or U1165 (N_1165,N_929,N_833);
and U1166 (N_1166,N_839,N_925);
nand U1167 (N_1167,N_836,N_955);
nand U1168 (N_1168,N_890,N_893);
nand U1169 (N_1169,N_873,N_863);
nand U1170 (N_1170,N_961,N_958);
and U1171 (N_1171,N_921,N_941);
or U1172 (N_1172,N_954,N_833);
or U1173 (N_1173,N_936,N_943);
and U1174 (N_1174,N_927,N_934);
or U1175 (N_1175,N_870,N_914);
nand U1176 (N_1176,N_811,N_836);
or U1177 (N_1177,N_949,N_960);
or U1178 (N_1178,N_850,N_918);
nor U1179 (N_1179,N_834,N_993);
nand U1180 (N_1180,N_838,N_915);
nand U1181 (N_1181,N_849,N_856);
and U1182 (N_1182,N_989,N_901);
nor U1183 (N_1183,N_902,N_931);
nand U1184 (N_1184,N_801,N_816);
nand U1185 (N_1185,N_939,N_909);
nor U1186 (N_1186,N_829,N_885);
nand U1187 (N_1187,N_931,N_965);
and U1188 (N_1188,N_856,N_949);
or U1189 (N_1189,N_882,N_814);
nand U1190 (N_1190,N_935,N_970);
nand U1191 (N_1191,N_840,N_835);
and U1192 (N_1192,N_940,N_802);
or U1193 (N_1193,N_928,N_835);
nor U1194 (N_1194,N_805,N_959);
or U1195 (N_1195,N_880,N_919);
nand U1196 (N_1196,N_811,N_937);
nor U1197 (N_1197,N_901,N_818);
and U1198 (N_1198,N_928,N_908);
nor U1199 (N_1199,N_943,N_990);
nand U1200 (N_1200,N_1066,N_1093);
and U1201 (N_1201,N_1046,N_1025);
and U1202 (N_1202,N_1043,N_1016);
and U1203 (N_1203,N_1050,N_1071);
and U1204 (N_1204,N_1088,N_1157);
or U1205 (N_1205,N_1196,N_1040);
nand U1206 (N_1206,N_1119,N_1121);
and U1207 (N_1207,N_1104,N_1031);
nand U1208 (N_1208,N_1154,N_1173);
nand U1209 (N_1209,N_1064,N_1117);
nor U1210 (N_1210,N_1092,N_1059);
nor U1211 (N_1211,N_1091,N_1185);
nor U1212 (N_1212,N_1168,N_1027);
nand U1213 (N_1213,N_1160,N_1035);
or U1214 (N_1214,N_1177,N_1130);
and U1215 (N_1215,N_1165,N_1105);
or U1216 (N_1216,N_1118,N_1017);
nand U1217 (N_1217,N_1137,N_1174);
nor U1218 (N_1218,N_1026,N_1183);
nand U1219 (N_1219,N_1187,N_1170);
or U1220 (N_1220,N_1002,N_1044);
and U1221 (N_1221,N_1139,N_1065);
and U1222 (N_1222,N_1129,N_1111);
nand U1223 (N_1223,N_1100,N_1024);
and U1224 (N_1224,N_1041,N_1166);
nand U1225 (N_1225,N_1193,N_1136);
and U1226 (N_1226,N_1133,N_1009);
and U1227 (N_1227,N_1152,N_1135);
nor U1228 (N_1228,N_1124,N_1120);
nor U1229 (N_1229,N_1055,N_1158);
and U1230 (N_1230,N_1029,N_1097);
and U1231 (N_1231,N_1192,N_1090);
nand U1232 (N_1232,N_1075,N_1030);
and U1233 (N_1233,N_1003,N_1047);
or U1234 (N_1234,N_1038,N_1186);
xnor U1235 (N_1235,N_1179,N_1072);
nand U1236 (N_1236,N_1085,N_1132);
and U1237 (N_1237,N_1079,N_1062);
nor U1238 (N_1238,N_1051,N_1042);
or U1239 (N_1239,N_1109,N_1014);
or U1240 (N_1240,N_1069,N_1045);
nor U1241 (N_1241,N_1018,N_1161);
or U1242 (N_1242,N_1061,N_1167);
or U1243 (N_1243,N_1163,N_1140);
and U1244 (N_1244,N_1034,N_1149);
nor U1245 (N_1245,N_1015,N_1068);
nor U1246 (N_1246,N_1058,N_1028);
and U1247 (N_1247,N_1176,N_1073);
or U1248 (N_1248,N_1110,N_1067);
or U1249 (N_1249,N_1122,N_1115);
or U1250 (N_1250,N_1142,N_1178);
nand U1251 (N_1251,N_1123,N_1021);
nand U1252 (N_1252,N_1172,N_1011);
nor U1253 (N_1253,N_1189,N_1008);
nor U1254 (N_1254,N_1083,N_1150);
nand U1255 (N_1255,N_1020,N_1127);
nand U1256 (N_1256,N_1169,N_1007);
nand U1257 (N_1257,N_1039,N_1155);
nand U1258 (N_1258,N_1175,N_1099);
or U1259 (N_1259,N_1087,N_1146);
nor U1260 (N_1260,N_1147,N_1005);
nand U1261 (N_1261,N_1125,N_1191);
or U1262 (N_1262,N_1080,N_1076);
nor U1263 (N_1263,N_1126,N_1103);
nand U1264 (N_1264,N_1096,N_1144);
and U1265 (N_1265,N_1153,N_1048);
nand U1266 (N_1266,N_1112,N_1106);
nor U1267 (N_1267,N_1114,N_1084);
and U1268 (N_1268,N_1060,N_1164);
or U1269 (N_1269,N_1162,N_1010);
and U1270 (N_1270,N_1134,N_1098);
and U1271 (N_1271,N_1023,N_1052);
nand U1272 (N_1272,N_1116,N_1077);
or U1273 (N_1273,N_1082,N_1081);
nor U1274 (N_1274,N_1156,N_1053);
nand U1275 (N_1275,N_1188,N_1180);
and U1276 (N_1276,N_1190,N_1128);
and U1277 (N_1277,N_1004,N_1145);
and U1278 (N_1278,N_1006,N_1022);
nor U1279 (N_1279,N_1151,N_1102);
or U1280 (N_1280,N_1032,N_1199);
nor U1281 (N_1281,N_1001,N_1108);
and U1282 (N_1282,N_1113,N_1074);
or U1283 (N_1283,N_1036,N_1181);
and U1284 (N_1284,N_1197,N_1107);
or U1285 (N_1285,N_1141,N_1019);
nand U1286 (N_1286,N_1138,N_1159);
nand U1287 (N_1287,N_1194,N_1131);
nor U1288 (N_1288,N_1063,N_1049);
nor U1289 (N_1289,N_1184,N_1195);
or U1290 (N_1290,N_1089,N_1143);
nand U1291 (N_1291,N_1056,N_1054);
nand U1292 (N_1292,N_1033,N_1070);
or U1293 (N_1293,N_1094,N_1000);
and U1294 (N_1294,N_1198,N_1182);
nor U1295 (N_1295,N_1086,N_1037);
and U1296 (N_1296,N_1012,N_1078);
and U1297 (N_1297,N_1095,N_1171);
nand U1298 (N_1298,N_1013,N_1057);
nand U1299 (N_1299,N_1148,N_1101);
nand U1300 (N_1300,N_1171,N_1083);
or U1301 (N_1301,N_1114,N_1000);
nor U1302 (N_1302,N_1059,N_1115);
xnor U1303 (N_1303,N_1156,N_1173);
nor U1304 (N_1304,N_1185,N_1067);
nor U1305 (N_1305,N_1001,N_1098);
or U1306 (N_1306,N_1012,N_1079);
or U1307 (N_1307,N_1153,N_1131);
nand U1308 (N_1308,N_1138,N_1069);
nand U1309 (N_1309,N_1134,N_1132);
nand U1310 (N_1310,N_1126,N_1052);
or U1311 (N_1311,N_1054,N_1147);
nor U1312 (N_1312,N_1071,N_1162);
or U1313 (N_1313,N_1051,N_1029);
nand U1314 (N_1314,N_1178,N_1038);
and U1315 (N_1315,N_1119,N_1067);
nand U1316 (N_1316,N_1156,N_1120);
and U1317 (N_1317,N_1114,N_1111);
nor U1318 (N_1318,N_1050,N_1195);
nand U1319 (N_1319,N_1042,N_1108);
or U1320 (N_1320,N_1120,N_1017);
or U1321 (N_1321,N_1070,N_1035);
nor U1322 (N_1322,N_1029,N_1012);
and U1323 (N_1323,N_1007,N_1080);
and U1324 (N_1324,N_1148,N_1011);
nand U1325 (N_1325,N_1160,N_1097);
or U1326 (N_1326,N_1089,N_1134);
or U1327 (N_1327,N_1130,N_1174);
or U1328 (N_1328,N_1121,N_1048);
nor U1329 (N_1329,N_1131,N_1008);
nand U1330 (N_1330,N_1081,N_1027);
and U1331 (N_1331,N_1108,N_1031);
or U1332 (N_1332,N_1130,N_1027);
nand U1333 (N_1333,N_1074,N_1079);
and U1334 (N_1334,N_1194,N_1152);
and U1335 (N_1335,N_1102,N_1176);
or U1336 (N_1336,N_1192,N_1124);
or U1337 (N_1337,N_1121,N_1020);
or U1338 (N_1338,N_1110,N_1098);
nor U1339 (N_1339,N_1012,N_1184);
and U1340 (N_1340,N_1031,N_1036);
nand U1341 (N_1341,N_1068,N_1170);
nor U1342 (N_1342,N_1159,N_1121);
nor U1343 (N_1343,N_1037,N_1032);
xnor U1344 (N_1344,N_1027,N_1073);
and U1345 (N_1345,N_1196,N_1096);
and U1346 (N_1346,N_1187,N_1086);
nand U1347 (N_1347,N_1001,N_1051);
and U1348 (N_1348,N_1178,N_1186);
nand U1349 (N_1349,N_1087,N_1033);
nor U1350 (N_1350,N_1080,N_1022);
and U1351 (N_1351,N_1148,N_1136);
xor U1352 (N_1352,N_1033,N_1103);
nor U1353 (N_1353,N_1078,N_1018);
nor U1354 (N_1354,N_1086,N_1100);
nand U1355 (N_1355,N_1034,N_1179);
nor U1356 (N_1356,N_1066,N_1082);
and U1357 (N_1357,N_1014,N_1064);
or U1358 (N_1358,N_1120,N_1123);
and U1359 (N_1359,N_1014,N_1152);
nand U1360 (N_1360,N_1193,N_1051);
nand U1361 (N_1361,N_1154,N_1132);
nand U1362 (N_1362,N_1123,N_1083);
or U1363 (N_1363,N_1002,N_1069);
nor U1364 (N_1364,N_1197,N_1177);
or U1365 (N_1365,N_1158,N_1183);
and U1366 (N_1366,N_1102,N_1069);
nor U1367 (N_1367,N_1158,N_1021);
or U1368 (N_1368,N_1000,N_1059);
nor U1369 (N_1369,N_1086,N_1077);
nand U1370 (N_1370,N_1015,N_1052);
nand U1371 (N_1371,N_1183,N_1028);
or U1372 (N_1372,N_1096,N_1126);
and U1373 (N_1373,N_1189,N_1124);
nand U1374 (N_1374,N_1042,N_1064);
nor U1375 (N_1375,N_1086,N_1113);
or U1376 (N_1376,N_1129,N_1125);
nand U1377 (N_1377,N_1024,N_1022);
nor U1378 (N_1378,N_1029,N_1112);
and U1379 (N_1379,N_1048,N_1134);
or U1380 (N_1380,N_1036,N_1196);
nor U1381 (N_1381,N_1198,N_1119);
nand U1382 (N_1382,N_1069,N_1091);
and U1383 (N_1383,N_1180,N_1035);
and U1384 (N_1384,N_1124,N_1180);
or U1385 (N_1385,N_1118,N_1195);
or U1386 (N_1386,N_1128,N_1110);
nor U1387 (N_1387,N_1086,N_1180);
nor U1388 (N_1388,N_1136,N_1090);
and U1389 (N_1389,N_1150,N_1044);
or U1390 (N_1390,N_1003,N_1058);
nand U1391 (N_1391,N_1155,N_1088);
nand U1392 (N_1392,N_1103,N_1089);
nand U1393 (N_1393,N_1075,N_1162);
and U1394 (N_1394,N_1140,N_1022);
nand U1395 (N_1395,N_1182,N_1184);
or U1396 (N_1396,N_1084,N_1005);
nand U1397 (N_1397,N_1136,N_1174);
and U1398 (N_1398,N_1011,N_1187);
nand U1399 (N_1399,N_1039,N_1031);
nand U1400 (N_1400,N_1270,N_1226);
nand U1401 (N_1401,N_1319,N_1364);
and U1402 (N_1402,N_1325,N_1398);
or U1403 (N_1403,N_1278,N_1333);
nor U1404 (N_1404,N_1281,N_1315);
or U1405 (N_1405,N_1310,N_1258);
nand U1406 (N_1406,N_1371,N_1245);
or U1407 (N_1407,N_1248,N_1240);
nand U1408 (N_1408,N_1362,N_1316);
and U1409 (N_1409,N_1323,N_1296);
or U1410 (N_1410,N_1377,N_1369);
nand U1411 (N_1411,N_1290,N_1211);
nand U1412 (N_1412,N_1229,N_1206);
nor U1413 (N_1413,N_1274,N_1263);
and U1414 (N_1414,N_1228,N_1349);
xor U1415 (N_1415,N_1291,N_1380);
nor U1416 (N_1416,N_1300,N_1356);
xor U1417 (N_1417,N_1336,N_1328);
or U1418 (N_1418,N_1210,N_1326);
and U1419 (N_1419,N_1313,N_1312);
and U1420 (N_1420,N_1350,N_1268);
or U1421 (N_1421,N_1282,N_1277);
nand U1422 (N_1422,N_1217,N_1232);
or U1423 (N_1423,N_1353,N_1280);
and U1424 (N_1424,N_1394,N_1273);
and U1425 (N_1425,N_1203,N_1223);
nand U1426 (N_1426,N_1392,N_1256);
nand U1427 (N_1427,N_1236,N_1244);
nand U1428 (N_1428,N_1269,N_1321);
or U1429 (N_1429,N_1387,N_1322);
and U1430 (N_1430,N_1383,N_1209);
nand U1431 (N_1431,N_1287,N_1347);
and U1432 (N_1432,N_1397,N_1327);
nand U1433 (N_1433,N_1242,N_1324);
or U1434 (N_1434,N_1262,N_1395);
and U1435 (N_1435,N_1344,N_1303);
or U1436 (N_1436,N_1225,N_1332);
nand U1437 (N_1437,N_1218,N_1253);
or U1438 (N_1438,N_1304,N_1293);
nor U1439 (N_1439,N_1348,N_1261);
nor U1440 (N_1440,N_1202,N_1257);
xnor U1441 (N_1441,N_1250,N_1376);
and U1442 (N_1442,N_1288,N_1330);
or U1443 (N_1443,N_1289,N_1241);
nand U1444 (N_1444,N_1339,N_1255);
nand U1445 (N_1445,N_1351,N_1302);
and U1446 (N_1446,N_1357,N_1360);
nor U1447 (N_1447,N_1301,N_1345);
nor U1448 (N_1448,N_1393,N_1317);
xor U1449 (N_1449,N_1213,N_1286);
and U1450 (N_1450,N_1243,N_1222);
and U1451 (N_1451,N_1205,N_1352);
and U1452 (N_1452,N_1237,N_1389);
nand U1453 (N_1453,N_1285,N_1238);
and U1454 (N_1454,N_1335,N_1254);
and U1455 (N_1455,N_1386,N_1361);
nand U1456 (N_1456,N_1391,N_1234);
nor U1457 (N_1457,N_1382,N_1396);
and U1458 (N_1458,N_1329,N_1271);
nand U1459 (N_1459,N_1272,N_1221);
and U1460 (N_1460,N_1311,N_1385);
and U1461 (N_1461,N_1299,N_1201);
and U1462 (N_1462,N_1341,N_1233);
nor U1463 (N_1463,N_1267,N_1375);
nand U1464 (N_1464,N_1388,N_1283);
and U1465 (N_1465,N_1252,N_1359);
or U1466 (N_1466,N_1340,N_1370);
nand U1467 (N_1467,N_1390,N_1338);
and U1468 (N_1468,N_1305,N_1227);
nand U1469 (N_1469,N_1294,N_1320);
nor U1470 (N_1470,N_1284,N_1378);
nand U1471 (N_1471,N_1247,N_1220);
nand U1472 (N_1472,N_1342,N_1231);
nand U1473 (N_1473,N_1314,N_1251);
or U1474 (N_1474,N_1307,N_1373);
or U1475 (N_1475,N_1260,N_1354);
or U1476 (N_1476,N_1384,N_1214);
nand U1477 (N_1477,N_1239,N_1297);
and U1478 (N_1478,N_1246,N_1358);
nand U1479 (N_1479,N_1346,N_1276);
and U1480 (N_1480,N_1399,N_1230);
and U1481 (N_1481,N_1308,N_1365);
nor U1482 (N_1482,N_1355,N_1331);
nor U1483 (N_1483,N_1363,N_1367);
nor U1484 (N_1484,N_1215,N_1295);
nor U1485 (N_1485,N_1212,N_1368);
nor U1486 (N_1486,N_1334,N_1318);
nor U1487 (N_1487,N_1204,N_1266);
and U1488 (N_1488,N_1235,N_1381);
nand U1489 (N_1489,N_1249,N_1275);
xnor U1490 (N_1490,N_1219,N_1374);
nand U1491 (N_1491,N_1208,N_1216);
or U1492 (N_1492,N_1224,N_1207);
and U1493 (N_1493,N_1306,N_1200);
or U1494 (N_1494,N_1265,N_1337);
or U1495 (N_1495,N_1379,N_1264);
and U1496 (N_1496,N_1343,N_1366);
or U1497 (N_1497,N_1298,N_1279);
and U1498 (N_1498,N_1292,N_1259);
nor U1499 (N_1499,N_1372,N_1309);
nand U1500 (N_1500,N_1211,N_1294);
nand U1501 (N_1501,N_1208,N_1321);
nor U1502 (N_1502,N_1253,N_1259);
nor U1503 (N_1503,N_1289,N_1269);
nor U1504 (N_1504,N_1346,N_1286);
nand U1505 (N_1505,N_1356,N_1399);
nand U1506 (N_1506,N_1301,N_1235);
or U1507 (N_1507,N_1372,N_1290);
nand U1508 (N_1508,N_1306,N_1227);
or U1509 (N_1509,N_1226,N_1325);
nor U1510 (N_1510,N_1330,N_1313);
and U1511 (N_1511,N_1243,N_1387);
nand U1512 (N_1512,N_1352,N_1215);
nand U1513 (N_1513,N_1226,N_1285);
and U1514 (N_1514,N_1246,N_1290);
and U1515 (N_1515,N_1222,N_1274);
nor U1516 (N_1516,N_1378,N_1257);
nand U1517 (N_1517,N_1272,N_1399);
and U1518 (N_1518,N_1396,N_1280);
and U1519 (N_1519,N_1227,N_1268);
and U1520 (N_1520,N_1389,N_1219);
or U1521 (N_1521,N_1399,N_1359);
or U1522 (N_1522,N_1273,N_1280);
nand U1523 (N_1523,N_1229,N_1224);
nand U1524 (N_1524,N_1320,N_1332);
and U1525 (N_1525,N_1293,N_1264);
nor U1526 (N_1526,N_1341,N_1243);
and U1527 (N_1527,N_1259,N_1288);
nor U1528 (N_1528,N_1277,N_1320);
nor U1529 (N_1529,N_1230,N_1336);
or U1530 (N_1530,N_1371,N_1277);
or U1531 (N_1531,N_1370,N_1327);
nand U1532 (N_1532,N_1341,N_1203);
nand U1533 (N_1533,N_1339,N_1240);
nor U1534 (N_1534,N_1315,N_1248);
nor U1535 (N_1535,N_1241,N_1305);
nor U1536 (N_1536,N_1375,N_1369);
nand U1537 (N_1537,N_1318,N_1293);
and U1538 (N_1538,N_1368,N_1302);
nand U1539 (N_1539,N_1360,N_1210);
or U1540 (N_1540,N_1392,N_1370);
nand U1541 (N_1541,N_1205,N_1202);
and U1542 (N_1542,N_1327,N_1354);
and U1543 (N_1543,N_1228,N_1328);
and U1544 (N_1544,N_1243,N_1318);
nor U1545 (N_1545,N_1352,N_1338);
and U1546 (N_1546,N_1345,N_1218);
nor U1547 (N_1547,N_1344,N_1294);
or U1548 (N_1548,N_1284,N_1201);
nand U1549 (N_1549,N_1241,N_1209);
and U1550 (N_1550,N_1323,N_1389);
nor U1551 (N_1551,N_1293,N_1250);
nand U1552 (N_1552,N_1391,N_1208);
nand U1553 (N_1553,N_1364,N_1285);
nor U1554 (N_1554,N_1279,N_1244);
xor U1555 (N_1555,N_1321,N_1346);
nor U1556 (N_1556,N_1367,N_1327);
or U1557 (N_1557,N_1303,N_1381);
nand U1558 (N_1558,N_1341,N_1332);
nand U1559 (N_1559,N_1282,N_1306);
nor U1560 (N_1560,N_1386,N_1384);
nand U1561 (N_1561,N_1254,N_1330);
or U1562 (N_1562,N_1205,N_1262);
or U1563 (N_1563,N_1295,N_1369);
nand U1564 (N_1564,N_1257,N_1342);
or U1565 (N_1565,N_1263,N_1243);
nor U1566 (N_1566,N_1325,N_1234);
or U1567 (N_1567,N_1215,N_1228);
nand U1568 (N_1568,N_1324,N_1262);
nor U1569 (N_1569,N_1341,N_1336);
and U1570 (N_1570,N_1297,N_1396);
and U1571 (N_1571,N_1332,N_1200);
and U1572 (N_1572,N_1290,N_1320);
and U1573 (N_1573,N_1232,N_1363);
or U1574 (N_1574,N_1335,N_1384);
nand U1575 (N_1575,N_1375,N_1235);
or U1576 (N_1576,N_1252,N_1336);
nor U1577 (N_1577,N_1382,N_1294);
and U1578 (N_1578,N_1394,N_1380);
nor U1579 (N_1579,N_1381,N_1323);
and U1580 (N_1580,N_1302,N_1339);
or U1581 (N_1581,N_1340,N_1267);
or U1582 (N_1582,N_1350,N_1395);
xor U1583 (N_1583,N_1295,N_1296);
nand U1584 (N_1584,N_1396,N_1253);
nor U1585 (N_1585,N_1382,N_1218);
or U1586 (N_1586,N_1359,N_1303);
nor U1587 (N_1587,N_1377,N_1360);
or U1588 (N_1588,N_1294,N_1317);
or U1589 (N_1589,N_1256,N_1279);
nor U1590 (N_1590,N_1388,N_1262);
nor U1591 (N_1591,N_1348,N_1253);
nand U1592 (N_1592,N_1354,N_1318);
nor U1593 (N_1593,N_1388,N_1334);
and U1594 (N_1594,N_1374,N_1213);
nor U1595 (N_1595,N_1303,N_1313);
nor U1596 (N_1596,N_1314,N_1201);
or U1597 (N_1597,N_1385,N_1273);
and U1598 (N_1598,N_1344,N_1311);
nand U1599 (N_1599,N_1393,N_1295);
and U1600 (N_1600,N_1576,N_1517);
or U1601 (N_1601,N_1522,N_1482);
nand U1602 (N_1602,N_1414,N_1594);
nor U1603 (N_1603,N_1416,N_1543);
nor U1604 (N_1604,N_1512,N_1508);
or U1605 (N_1605,N_1525,N_1528);
nor U1606 (N_1606,N_1431,N_1488);
and U1607 (N_1607,N_1439,N_1511);
nor U1608 (N_1608,N_1462,N_1577);
nor U1609 (N_1609,N_1432,N_1474);
nand U1610 (N_1610,N_1570,N_1535);
nor U1611 (N_1611,N_1583,N_1533);
or U1612 (N_1612,N_1481,N_1446);
or U1613 (N_1613,N_1538,N_1557);
or U1614 (N_1614,N_1598,N_1530);
and U1615 (N_1615,N_1447,N_1449);
and U1616 (N_1616,N_1561,N_1441);
nand U1617 (N_1617,N_1514,N_1501);
and U1618 (N_1618,N_1551,N_1458);
and U1619 (N_1619,N_1451,N_1578);
and U1620 (N_1620,N_1539,N_1411);
or U1621 (N_1621,N_1491,N_1548);
nand U1622 (N_1622,N_1541,N_1540);
nor U1623 (N_1623,N_1579,N_1567);
nor U1624 (N_1624,N_1554,N_1503);
and U1625 (N_1625,N_1582,N_1587);
nor U1626 (N_1626,N_1562,N_1599);
nand U1627 (N_1627,N_1590,N_1572);
and U1628 (N_1628,N_1592,N_1495);
nand U1629 (N_1629,N_1448,N_1526);
or U1630 (N_1630,N_1549,N_1407);
and U1631 (N_1631,N_1523,N_1473);
nand U1632 (N_1632,N_1454,N_1437);
or U1633 (N_1633,N_1415,N_1468);
or U1634 (N_1634,N_1597,N_1430);
and U1635 (N_1635,N_1521,N_1585);
and U1636 (N_1636,N_1450,N_1435);
nor U1637 (N_1637,N_1479,N_1445);
nand U1638 (N_1638,N_1575,N_1493);
or U1639 (N_1639,N_1403,N_1565);
and U1640 (N_1640,N_1589,N_1586);
and U1641 (N_1641,N_1553,N_1552);
nor U1642 (N_1642,N_1515,N_1485);
or U1643 (N_1643,N_1534,N_1452);
and U1644 (N_1644,N_1519,N_1404);
nor U1645 (N_1645,N_1467,N_1444);
or U1646 (N_1646,N_1555,N_1588);
and U1647 (N_1647,N_1424,N_1584);
nand U1648 (N_1648,N_1593,N_1571);
or U1649 (N_1649,N_1433,N_1580);
or U1650 (N_1650,N_1560,N_1470);
nor U1651 (N_1651,N_1504,N_1544);
and U1652 (N_1652,N_1478,N_1400);
or U1653 (N_1653,N_1486,N_1496);
or U1654 (N_1654,N_1546,N_1475);
nand U1655 (N_1655,N_1509,N_1505);
nor U1656 (N_1656,N_1401,N_1559);
and U1657 (N_1657,N_1426,N_1547);
nor U1658 (N_1658,N_1428,N_1492);
or U1659 (N_1659,N_1516,N_1455);
nand U1660 (N_1660,N_1410,N_1408);
and U1661 (N_1661,N_1440,N_1418);
nand U1662 (N_1662,N_1550,N_1513);
and U1663 (N_1663,N_1510,N_1558);
and U1664 (N_1664,N_1569,N_1499);
or U1665 (N_1665,N_1484,N_1596);
or U1666 (N_1666,N_1419,N_1436);
or U1667 (N_1667,N_1472,N_1461);
xnor U1668 (N_1668,N_1480,N_1469);
nand U1669 (N_1669,N_1425,N_1497);
or U1670 (N_1670,N_1456,N_1542);
or U1671 (N_1671,N_1420,N_1409);
nand U1672 (N_1672,N_1532,N_1556);
and U1673 (N_1673,N_1581,N_1498);
nand U1674 (N_1674,N_1563,N_1490);
or U1675 (N_1675,N_1412,N_1477);
nor U1676 (N_1676,N_1423,N_1413);
nand U1677 (N_1677,N_1465,N_1489);
nand U1678 (N_1678,N_1564,N_1457);
nand U1679 (N_1679,N_1545,N_1402);
or U1680 (N_1680,N_1417,N_1591);
nand U1681 (N_1681,N_1422,N_1453);
nor U1682 (N_1682,N_1438,N_1500);
nand U1683 (N_1683,N_1427,N_1476);
nor U1684 (N_1684,N_1494,N_1443);
nand U1685 (N_1685,N_1460,N_1531);
and U1686 (N_1686,N_1459,N_1464);
or U1687 (N_1687,N_1527,N_1529);
nor U1688 (N_1688,N_1434,N_1566);
nand U1689 (N_1689,N_1524,N_1507);
nand U1690 (N_1690,N_1406,N_1573);
nor U1691 (N_1691,N_1502,N_1466);
and U1692 (N_1692,N_1405,N_1483);
or U1693 (N_1693,N_1471,N_1421);
nand U1694 (N_1694,N_1487,N_1595);
nor U1695 (N_1695,N_1506,N_1568);
or U1696 (N_1696,N_1536,N_1463);
or U1697 (N_1697,N_1429,N_1574);
nand U1698 (N_1698,N_1520,N_1442);
and U1699 (N_1699,N_1537,N_1518);
or U1700 (N_1700,N_1538,N_1406);
nor U1701 (N_1701,N_1406,N_1509);
and U1702 (N_1702,N_1588,N_1457);
nand U1703 (N_1703,N_1435,N_1532);
and U1704 (N_1704,N_1500,N_1593);
nor U1705 (N_1705,N_1547,N_1566);
and U1706 (N_1706,N_1505,N_1407);
nor U1707 (N_1707,N_1513,N_1490);
xnor U1708 (N_1708,N_1477,N_1525);
nand U1709 (N_1709,N_1564,N_1559);
nand U1710 (N_1710,N_1587,N_1562);
or U1711 (N_1711,N_1509,N_1526);
and U1712 (N_1712,N_1439,N_1539);
or U1713 (N_1713,N_1473,N_1403);
nand U1714 (N_1714,N_1492,N_1541);
nand U1715 (N_1715,N_1514,N_1519);
nand U1716 (N_1716,N_1528,N_1574);
or U1717 (N_1717,N_1414,N_1466);
nand U1718 (N_1718,N_1410,N_1541);
and U1719 (N_1719,N_1422,N_1510);
or U1720 (N_1720,N_1478,N_1446);
or U1721 (N_1721,N_1508,N_1410);
or U1722 (N_1722,N_1485,N_1578);
and U1723 (N_1723,N_1504,N_1445);
nand U1724 (N_1724,N_1529,N_1564);
nand U1725 (N_1725,N_1482,N_1489);
xnor U1726 (N_1726,N_1481,N_1406);
or U1727 (N_1727,N_1442,N_1430);
and U1728 (N_1728,N_1436,N_1467);
and U1729 (N_1729,N_1569,N_1503);
or U1730 (N_1730,N_1428,N_1467);
and U1731 (N_1731,N_1436,N_1543);
nand U1732 (N_1732,N_1534,N_1573);
nand U1733 (N_1733,N_1494,N_1581);
nor U1734 (N_1734,N_1506,N_1521);
nand U1735 (N_1735,N_1527,N_1494);
and U1736 (N_1736,N_1480,N_1594);
and U1737 (N_1737,N_1577,N_1565);
and U1738 (N_1738,N_1468,N_1426);
nand U1739 (N_1739,N_1455,N_1552);
and U1740 (N_1740,N_1566,N_1544);
and U1741 (N_1741,N_1528,N_1480);
and U1742 (N_1742,N_1408,N_1451);
nor U1743 (N_1743,N_1516,N_1533);
and U1744 (N_1744,N_1468,N_1480);
nand U1745 (N_1745,N_1443,N_1490);
and U1746 (N_1746,N_1464,N_1531);
nor U1747 (N_1747,N_1400,N_1405);
and U1748 (N_1748,N_1592,N_1586);
nor U1749 (N_1749,N_1588,N_1564);
nand U1750 (N_1750,N_1531,N_1478);
nand U1751 (N_1751,N_1488,N_1521);
nand U1752 (N_1752,N_1444,N_1483);
nand U1753 (N_1753,N_1440,N_1565);
or U1754 (N_1754,N_1596,N_1568);
or U1755 (N_1755,N_1485,N_1525);
or U1756 (N_1756,N_1425,N_1427);
nand U1757 (N_1757,N_1513,N_1578);
and U1758 (N_1758,N_1515,N_1572);
and U1759 (N_1759,N_1557,N_1473);
or U1760 (N_1760,N_1456,N_1450);
nand U1761 (N_1761,N_1478,N_1564);
and U1762 (N_1762,N_1464,N_1451);
or U1763 (N_1763,N_1467,N_1430);
nand U1764 (N_1764,N_1528,N_1592);
nand U1765 (N_1765,N_1596,N_1438);
nor U1766 (N_1766,N_1592,N_1599);
nor U1767 (N_1767,N_1441,N_1469);
nand U1768 (N_1768,N_1583,N_1516);
nor U1769 (N_1769,N_1512,N_1445);
and U1770 (N_1770,N_1528,N_1582);
nand U1771 (N_1771,N_1414,N_1412);
nor U1772 (N_1772,N_1469,N_1593);
and U1773 (N_1773,N_1508,N_1548);
and U1774 (N_1774,N_1519,N_1405);
or U1775 (N_1775,N_1557,N_1549);
or U1776 (N_1776,N_1438,N_1514);
nand U1777 (N_1777,N_1498,N_1406);
or U1778 (N_1778,N_1494,N_1418);
nor U1779 (N_1779,N_1421,N_1534);
nand U1780 (N_1780,N_1438,N_1508);
nor U1781 (N_1781,N_1463,N_1483);
or U1782 (N_1782,N_1492,N_1534);
or U1783 (N_1783,N_1525,N_1545);
nand U1784 (N_1784,N_1486,N_1577);
nand U1785 (N_1785,N_1598,N_1553);
or U1786 (N_1786,N_1515,N_1567);
or U1787 (N_1787,N_1400,N_1562);
nand U1788 (N_1788,N_1540,N_1408);
or U1789 (N_1789,N_1578,N_1595);
or U1790 (N_1790,N_1524,N_1488);
or U1791 (N_1791,N_1538,N_1563);
and U1792 (N_1792,N_1460,N_1506);
nor U1793 (N_1793,N_1481,N_1488);
and U1794 (N_1794,N_1454,N_1572);
or U1795 (N_1795,N_1513,N_1478);
and U1796 (N_1796,N_1534,N_1473);
nor U1797 (N_1797,N_1447,N_1555);
nand U1798 (N_1798,N_1569,N_1516);
or U1799 (N_1799,N_1473,N_1563);
nand U1800 (N_1800,N_1795,N_1770);
or U1801 (N_1801,N_1749,N_1635);
or U1802 (N_1802,N_1641,N_1728);
nor U1803 (N_1803,N_1600,N_1636);
or U1804 (N_1804,N_1796,N_1703);
or U1805 (N_1805,N_1702,N_1697);
or U1806 (N_1806,N_1760,N_1689);
nand U1807 (N_1807,N_1683,N_1738);
nand U1808 (N_1808,N_1656,N_1691);
nand U1809 (N_1809,N_1752,N_1696);
nand U1810 (N_1810,N_1693,N_1648);
and U1811 (N_1811,N_1637,N_1632);
and U1812 (N_1812,N_1616,N_1649);
or U1813 (N_1813,N_1720,N_1774);
and U1814 (N_1814,N_1751,N_1747);
nor U1815 (N_1815,N_1629,N_1737);
or U1816 (N_1816,N_1646,N_1617);
or U1817 (N_1817,N_1706,N_1692);
or U1818 (N_1818,N_1647,N_1654);
nor U1819 (N_1819,N_1726,N_1682);
or U1820 (N_1820,N_1677,N_1766);
and U1821 (N_1821,N_1783,N_1773);
or U1822 (N_1822,N_1622,N_1750);
or U1823 (N_1823,N_1605,N_1763);
nor U1824 (N_1824,N_1761,N_1615);
nor U1825 (N_1825,N_1607,N_1765);
or U1826 (N_1826,N_1601,N_1700);
nand U1827 (N_1827,N_1671,N_1608);
or U1828 (N_1828,N_1757,N_1781);
or U1829 (N_1829,N_1694,N_1735);
nor U1830 (N_1830,N_1707,N_1665);
nor U1831 (N_1831,N_1606,N_1745);
nor U1832 (N_1832,N_1681,N_1744);
and U1833 (N_1833,N_1715,N_1621);
and U1834 (N_1834,N_1734,N_1784);
and U1835 (N_1835,N_1624,N_1713);
nor U1836 (N_1836,N_1643,N_1674);
or U1837 (N_1837,N_1759,N_1709);
nand U1838 (N_1838,N_1631,N_1791);
nor U1839 (N_1839,N_1739,N_1613);
nand U1840 (N_1840,N_1730,N_1618);
or U1841 (N_1841,N_1782,N_1764);
nand U1842 (N_1842,N_1663,N_1772);
nand U1843 (N_1843,N_1667,N_1655);
nor U1844 (N_1844,N_1708,N_1630);
nor U1845 (N_1845,N_1602,N_1793);
or U1846 (N_1846,N_1776,N_1639);
and U1847 (N_1847,N_1798,N_1625);
nand U1848 (N_1848,N_1695,N_1657);
and U1849 (N_1849,N_1789,N_1741);
and U1850 (N_1850,N_1660,N_1669);
and U1851 (N_1851,N_1699,N_1668);
or U1852 (N_1852,N_1628,N_1797);
nor U1853 (N_1853,N_1725,N_1661);
or U1854 (N_1854,N_1690,N_1620);
or U1855 (N_1855,N_1729,N_1685);
nor U1856 (N_1856,N_1609,N_1673);
nand U1857 (N_1857,N_1788,N_1792);
nand U1858 (N_1858,N_1701,N_1645);
and U1859 (N_1859,N_1658,N_1704);
and U1860 (N_1860,N_1780,N_1698);
nor U1861 (N_1861,N_1659,N_1653);
nor U1862 (N_1862,N_1705,N_1724);
nand U1863 (N_1863,N_1771,N_1650);
nand U1864 (N_1864,N_1614,N_1619);
or U1865 (N_1865,N_1758,N_1678);
or U1866 (N_1866,N_1640,N_1686);
or U1867 (N_1867,N_1768,N_1718);
nor U1868 (N_1868,N_1779,N_1664);
or U1869 (N_1869,N_1627,N_1633);
nor U1870 (N_1870,N_1722,N_1799);
nor U1871 (N_1871,N_1767,N_1688);
nor U1872 (N_1872,N_1604,N_1762);
and U1873 (N_1873,N_1710,N_1743);
or U1874 (N_1874,N_1623,N_1756);
xor U1875 (N_1875,N_1714,N_1626);
nand U1876 (N_1876,N_1716,N_1740);
xnor U1877 (N_1877,N_1727,N_1610);
nand U1878 (N_1878,N_1638,N_1755);
or U1879 (N_1879,N_1721,N_1642);
or U1880 (N_1880,N_1687,N_1679);
nor U1881 (N_1881,N_1711,N_1712);
nor U1882 (N_1882,N_1675,N_1670);
nor U1883 (N_1883,N_1754,N_1736);
or U1884 (N_1884,N_1603,N_1634);
nand U1885 (N_1885,N_1732,N_1786);
or U1886 (N_1886,N_1794,N_1723);
and U1887 (N_1887,N_1651,N_1666);
nor U1888 (N_1888,N_1787,N_1790);
nand U1889 (N_1889,N_1733,N_1785);
and U1890 (N_1890,N_1611,N_1672);
nor U1891 (N_1891,N_1746,N_1612);
nor U1892 (N_1892,N_1680,N_1719);
and U1893 (N_1893,N_1769,N_1731);
nor U1894 (N_1894,N_1775,N_1684);
or U1895 (N_1895,N_1748,N_1778);
and U1896 (N_1896,N_1777,N_1652);
and U1897 (N_1897,N_1753,N_1644);
or U1898 (N_1898,N_1742,N_1676);
and U1899 (N_1899,N_1717,N_1662);
xnor U1900 (N_1900,N_1740,N_1713);
nand U1901 (N_1901,N_1772,N_1757);
nand U1902 (N_1902,N_1784,N_1799);
and U1903 (N_1903,N_1709,N_1622);
nor U1904 (N_1904,N_1779,N_1660);
nor U1905 (N_1905,N_1655,N_1775);
nor U1906 (N_1906,N_1735,N_1645);
and U1907 (N_1907,N_1753,N_1637);
nand U1908 (N_1908,N_1742,N_1660);
or U1909 (N_1909,N_1682,N_1674);
or U1910 (N_1910,N_1758,N_1680);
nor U1911 (N_1911,N_1707,N_1649);
or U1912 (N_1912,N_1719,N_1764);
and U1913 (N_1913,N_1645,N_1673);
or U1914 (N_1914,N_1631,N_1749);
nand U1915 (N_1915,N_1775,N_1648);
nand U1916 (N_1916,N_1611,N_1747);
or U1917 (N_1917,N_1771,N_1658);
nor U1918 (N_1918,N_1699,N_1778);
xnor U1919 (N_1919,N_1725,N_1765);
nor U1920 (N_1920,N_1648,N_1633);
nor U1921 (N_1921,N_1740,N_1719);
or U1922 (N_1922,N_1640,N_1618);
nor U1923 (N_1923,N_1607,N_1645);
and U1924 (N_1924,N_1787,N_1726);
and U1925 (N_1925,N_1714,N_1718);
nand U1926 (N_1926,N_1733,N_1754);
nand U1927 (N_1927,N_1714,N_1756);
nand U1928 (N_1928,N_1640,N_1739);
nand U1929 (N_1929,N_1719,N_1683);
or U1930 (N_1930,N_1634,N_1686);
and U1931 (N_1931,N_1738,N_1766);
nor U1932 (N_1932,N_1608,N_1632);
nand U1933 (N_1933,N_1671,N_1722);
and U1934 (N_1934,N_1667,N_1657);
and U1935 (N_1935,N_1761,N_1709);
nor U1936 (N_1936,N_1735,N_1756);
and U1937 (N_1937,N_1690,N_1625);
nor U1938 (N_1938,N_1767,N_1634);
nand U1939 (N_1939,N_1792,N_1761);
nor U1940 (N_1940,N_1636,N_1620);
nand U1941 (N_1941,N_1665,N_1771);
nor U1942 (N_1942,N_1753,N_1649);
and U1943 (N_1943,N_1733,N_1702);
or U1944 (N_1944,N_1730,N_1711);
or U1945 (N_1945,N_1663,N_1758);
and U1946 (N_1946,N_1656,N_1600);
or U1947 (N_1947,N_1718,N_1797);
or U1948 (N_1948,N_1659,N_1641);
and U1949 (N_1949,N_1672,N_1667);
nand U1950 (N_1950,N_1604,N_1668);
or U1951 (N_1951,N_1648,N_1736);
or U1952 (N_1952,N_1747,N_1713);
or U1953 (N_1953,N_1738,N_1732);
and U1954 (N_1954,N_1787,N_1740);
nor U1955 (N_1955,N_1778,N_1609);
nand U1956 (N_1956,N_1759,N_1634);
and U1957 (N_1957,N_1663,N_1675);
nand U1958 (N_1958,N_1767,N_1671);
nor U1959 (N_1959,N_1672,N_1702);
nand U1960 (N_1960,N_1634,N_1619);
nor U1961 (N_1961,N_1753,N_1692);
nand U1962 (N_1962,N_1647,N_1770);
nor U1963 (N_1963,N_1676,N_1756);
or U1964 (N_1964,N_1673,N_1730);
and U1965 (N_1965,N_1601,N_1678);
and U1966 (N_1966,N_1667,N_1716);
and U1967 (N_1967,N_1766,N_1683);
or U1968 (N_1968,N_1662,N_1753);
nor U1969 (N_1969,N_1773,N_1758);
or U1970 (N_1970,N_1651,N_1702);
and U1971 (N_1971,N_1615,N_1710);
and U1972 (N_1972,N_1727,N_1604);
and U1973 (N_1973,N_1673,N_1763);
and U1974 (N_1974,N_1767,N_1694);
nor U1975 (N_1975,N_1686,N_1734);
and U1976 (N_1976,N_1788,N_1795);
nor U1977 (N_1977,N_1643,N_1759);
and U1978 (N_1978,N_1727,N_1726);
nand U1979 (N_1979,N_1711,N_1682);
and U1980 (N_1980,N_1667,N_1786);
nor U1981 (N_1981,N_1784,N_1713);
or U1982 (N_1982,N_1646,N_1677);
and U1983 (N_1983,N_1772,N_1730);
nor U1984 (N_1984,N_1715,N_1651);
or U1985 (N_1985,N_1754,N_1761);
or U1986 (N_1986,N_1673,N_1643);
and U1987 (N_1987,N_1699,N_1638);
nand U1988 (N_1988,N_1603,N_1632);
nand U1989 (N_1989,N_1685,N_1782);
and U1990 (N_1990,N_1625,N_1621);
or U1991 (N_1991,N_1680,N_1631);
nand U1992 (N_1992,N_1618,N_1663);
or U1993 (N_1993,N_1612,N_1736);
and U1994 (N_1994,N_1627,N_1737);
or U1995 (N_1995,N_1784,N_1685);
or U1996 (N_1996,N_1668,N_1732);
or U1997 (N_1997,N_1710,N_1622);
nand U1998 (N_1998,N_1630,N_1738);
or U1999 (N_1999,N_1767,N_1689);
or U2000 (N_2000,N_1949,N_1801);
nand U2001 (N_2001,N_1978,N_1937);
nor U2002 (N_2002,N_1811,N_1824);
or U2003 (N_2003,N_1928,N_1874);
and U2004 (N_2004,N_1871,N_1815);
or U2005 (N_2005,N_1860,N_1907);
nand U2006 (N_2006,N_1851,N_1955);
nand U2007 (N_2007,N_1879,N_1971);
and U2008 (N_2008,N_1926,N_1935);
or U2009 (N_2009,N_1808,N_1803);
nand U2010 (N_2010,N_1876,N_1950);
or U2011 (N_2011,N_1837,N_1968);
nand U2012 (N_2012,N_1983,N_1957);
and U2013 (N_2013,N_1966,N_1880);
nor U2014 (N_2014,N_1891,N_1838);
nand U2015 (N_2015,N_1840,N_1980);
and U2016 (N_2016,N_1910,N_1868);
or U2017 (N_2017,N_1967,N_1912);
nor U2018 (N_2018,N_1946,N_1836);
nand U2019 (N_2019,N_1988,N_1858);
nor U2020 (N_2020,N_1855,N_1816);
nand U2021 (N_2021,N_1959,N_1960);
or U2022 (N_2022,N_1850,N_1927);
nor U2023 (N_2023,N_1929,N_1911);
nor U2024 (N_2024,N_1873,N_1847);
and U2025 (N_2025,N_1898,N_1941);
or U2026 (N_2026,N_1992,N_1843);
and U2027 (N_2027,N_1896,N_1886);
and U2028 (N_2028,N_1982,N_1881);
nor U2029 (N_2029,N_1922,N_1953);
and U2030 (N_2030,N_1997,N_1807);
nand U2031 (N_2031,N_1852,N_1999);
or U2032 (N_2032,N_1817,N_1956);
nor U2033 (N_2033,N_1825,N_1913);
or U2034 (N_2034,N_1828,N_1904);
nor U2035 (N_2035,N_1854,N_1962);
nand U2036 (N_2036,N_1899,N_1931);
nand U2037 (N_2037,N_1882,N_1853);
nand U2038 (N_2038,N_1819,N_1975);
or U2039 (N_2039,N_1839,N_1844);
or U2040 (N_2040,N_1893,N_1859);
nand U2041 (N_2041,N_1892,N_1945);
or U2042 (N_2042,N_1933,N_1930);
nand U2043 (N_2043,N_1890,N_1921);
xor U2044 (N_2044,N_1845,N_1832);
or U2045 (N_2045,N_1924,N_1821);
nor U2046 (N_2046,N_1963,N_1936);
and U2047 (N_2047,N_1800,N_1866);
or U2048 (N_2048,N_1917,N_1867);
nand U2049 (N_2049,N_1834,N_1900);
nor U2050 (N_2050,N_1823,N_1806);
nor U2051 (N_2051,N_1835,N_1994);
or U2052 (N_2052,N_1932,N_1878);
nor U2053 (N_2053,N_1961,N_1986);
nand U2054 (N_2054,N_1830,N_1894);
or U2055 (N_2055,N_1903,N_1885);
nand U2056 (N_2056,N_1831,N_1901);
or U2057 (N_2057,N_1925,N_1862);
or U2058 (N_2058,N_1857,N_1954);
or U2059 (N_2059,N_1883,N_1849);
nand U2060 (N_2060,N_1914,N_1906);
nor U2061 (N_2061,N_1991,N_1948);
and U2062 (N_2062,N_1870,N_1947);
nor U2063 (N_2063,N_1919,N_1827);
nor U2064 (N_2064,N_1942,N_1993);
nor U2065 (N_2065,N_1820,N_1958);
and U2066 (N_2066,N_1923,N_1841);
nand U2067 (N_2067,N_1872,N_1969);
nand U2068 (N_2068,N_1984,N_1965);
nand U2069 (N_2069,N_1805,N_1829);
and U2070 (N_2070,N_1943,N_1809);
nor U2071 (N_2071,N_1875,N_1905);
nand U2072 (N_2072,N_1918,N_1814);
nand U2073 (N_2073,N_1856,N_1848);
or U2074 (N_2074,N_1822,N_1812);
and U2075 (N_2075,N_1915,N_1951);
or U2076 (N_2076,N_1884,N_1940);
nor U2077 (N_2077,N_1908,N_1833);
and U2078 (N_2078,N_1864,N_1861);
nor U2079 (N_2079,N_1964,N_1877);
nor U2080 (N_2080,N_1869,N_1863);
nand U2081 (N_2081,N_1985,N_1998);
nor U2082 (N_2082,N_1818,N_1916);
and U2083 (N_2083,N_1939,N_1887);
or U2084 (N_2084,N_1989,N_1976);
or U2085 (N_2085,N_1974,N_1804);
and U2086 (N_2086,N_1895,N_1909);
or U2087 (N_2087,N_1826,N_1987);
and U2088 (N_2088,N_1977,N_1952);
nor U2089 (N_2089,N_1995,N_1889);
or U2090 (N_2090,N_1902,N_1996);
or U2091 (N_2091,N_1979,N_1810);
and U2092 (N_2092,N_1981,N_1972);
nand U2093 (N_2093,N_1944,N_1920);
or U2094 (N_2094,N_1897,N_1865);
and U2095 (N_2095,N_1990,N_1802);
nor U2096 (N_2096,N_1934,N_1813);
nor U2097 (N_2097,N_1888,N_1973);
nand U2098 (N_2098,N_1846,N_1938);
nand U2099 (N_2099,N_1842,N_1970);
and U2100 (N_2100,N_1940,N_1948);
and U2101 (N_2101,N_1875,N_1974);
and U2102 (N_2102,N_1855,N_1802);
or U2103 (N_2103,N_1831,N_1984);
or U2104 (N_2104,N_1875,N_1958);
nand U2105 (N_2105,N_1941,N_1993);
nor U2106 (N_2106,N_1809,N_1989);
and U2107 (N_2107,N_1947,N_1904);
nand U2108 (N_2108,N_1982,N_1906);
or U2109 (N_2109,N_1994,N_1952);
nand U2110 (N_2110,N_1953,N_1968);
and U2111 (N_2111,N_1839,N_1827);
and U2112 (N_2112,N_1938,N_1876);
or U2113 (N_2113,N_1895,N_1806);
and U2114 (N_2114,N_1963,N_1973);
or U2115 (N_2115,N_1986,N_1982);
nor U2116 (N_2116,N_1926,N_1844);
nand U2117 (N_2117,N_1963,N_1804);
or U2118 (N_2118,N_1921,N_1816);
or U2119 (N_2119,N_1826,N_1974);
nand U2120 (N_2120,N_1945,N_1851);
nor U2121 (N_2121,N_1954,N_1852);
or U2122 (N_2122,N_1897,N_1871);
xnor U2123 (N_2123,N_1820,N_1934);
or U2124 (N_2124,N_1840,N_1806);
or U2125 (N_2125,N_1872,N_1811);
or U2126 (N_2126,N_1803,N_1942);
nor U2127 (N_2127,N_1806,N_1930);
or U2128 (N_2128,N_1867,N_1902);
and U2129 (N_2129,N_1830,N_1959);
and U2130 (N_2130,N_1809,N_1851);
nand U2131 (N_2131,N_1946,N_1975);
and U2132 (N_2132,N_1821,N_1888);
or U2133 (N_2133,N_1968,N_1993);
nor U2134 (N_2134,N_1971,N_1870);
nor U2135 (N_2135,N_1925,N_1900);
and U2136 (N_2136,N_1817,N_1849);
and U2137 (N_2137,N_1959,N_1995);
or U2138 (N_2138,N_1968,N_1864);
or U2139 (N_2139,N_1976,N_1851);
or U2140 (N_2140,N_1992,N_1808);
and U2141 (N_2141,N_1875,N_1944);
and U2142 (N_2142,N_1894,N_1987);
or U2143 (N_2143,N_1927,N_1901);
or U2144 (N_2144,N_1878,N_1987);
and U2145 (N_2145,N_1844,N_1913);
and U2146 (N_2146,N_1924,N_1975);
nor U2147 (N_2147,N_1891,N_1873);
nand U2148 (N_2148,N_1832,N_1800);
and U2149 (N_2149,N_1943,N_1939);
nor U2150 (N_2150,N_1974,N_1913);
nor U2151 (N_2151,N_1933,N_1897);
or U2152 (N_2152,N_1801,N_1881);
and U2153 (N_2153,N_1871,N_1981);
nand U2154 (N_2154,N_1979,N_1827);
and U2155 (N_2155,N_1998,N_1883);
nand U2156 (N_2156,N_1918,N_1961);
nand U2157 (N_2157,N_1861,N_1987);
and U2158 (N_2158,N_1876,N_1937);
and U2159 (N_2159,N_1820,N_1878);
and U2160 (N_2160,N_1809,N_1853);
and U2161 (N_2161,N_1900,N_1983);
and U2162 (N_2162,N_1878,N_1971);
or U2163 (N_2163,N_1920,N_1868);
and U2164 (N_2164,N_1974,N_1948);
nand U2165 (N_2165,N_1832,N_1809);
or U2166 (N_2166,N_1918,N_1811);
nand U2167 (N_2167,N_1848,N_1841);
nor U2168 (N_2168,N_1895,N_1948);
and U2169 (N_2169,N_1903,N_1834);
and U2170 (N_2170,N_1834,N_1879);
and U2171 (N_2171,N_1841,N_1958);
xor U2172 (N_2172,N_1871,N_1907);
nor U2173 (N_2173,N_1802,N_1809);
and U2174 (N_2174,N_1977,N_1862);
and U2175 (N_2175,N_1962,N_1816);
nor U2176 (N_2176,N_1867,N_1879);
or U2177 (N_2177,N_1947,N_1910);
nand U2178 (N_2178,N_1822,N_1959);
and U2179 (N_2179,N_1847,N_1853);
and U2180 (N_2180,N_1869,N_1871);
nand U2181 (N_2181,N_1825,N_1929);
or U2182 (N_2182,N_1812,N_1928);
and U2183 (N_2183,N_1991,N_1994);
and U2184 (N_2184,N_1867,N_1884);
and U2185 (N_2185,N_1856,N_1887);
nand U2186 (N_2186,N_1997,N_1856);
or U2187 (N_2187,N_1988,N_1916);
nand U2188 (N_2188,N_1841,N_1856);
nand U2189 (N_2189,N_1921,N_1853);
and U2190 (N_2190,N_1911,N_1949);
nor U2191 (N_2191,N_1993,N_1980);
nand U2192 (N_2192,N_1991,N_1813);
or U2193 (N_2193,N_1883,N_1921);
and U2194 (N_2194,N_1950,N_1813);
nor U2195 (N_2195,N_1862,N_1839);
nor U2196 (N_2196,N_1876,N_1839);
and U2197 (N_2197,N_1921,N_1848);
nand U2198 (N_2198,N_1964,N_1807);
or U2199 (N_2199,N_1878,N_1918);
nand U2200 (N_2200,N_2148,N_2161);
nand U2201 (N_2201,N_2063,N_2039);
nor U2202 (N_2202,N_2061,N_2015);
or U2203 (N_2203,N_2132,N_2195);
or U2204 (N_2204,N_2027,N_2090);
nand U2205 (N_2205,N_2141,N_2186);
nor U2206 (N_2206,N_2126,N_2182);
or U2207 (N_2207,N_2146,N_2175);
nor U2208 (N_2208,N_2120,N_2026);
nand U2209 (N_2209,N_2150,N_2049);
and U2210 (N_2210,N_2180,N_2054);
or U2211 (N_2211,N_2002,N_2174);
or U2212 (N_2212,N_2199,N_2038);
nand U2213 (N_2213,N_2151,N_2080);
and U2214 (N_2214,N_2031,N_2152);
nand U2215 (N_2215,N_2050,N_2144);
nand U2216 (N_2216,N_2022,N_2106);
nor U2217 (N_2217,N_2127,N_2094);
nor U2218 (N_2218,N_2165,N_2024);
nand U2219 (N_2219,N_2045,N_2133);
or U2220 (N_2220,N_2108,N_2083);
nor U2221 (N_2221,N_2000,N_2060);
or U2222 (N_2222,N_2142,N_2135);
or U2223 (N_2223,N_2157,N_2035);
nor U2224 (N_2224,N_2190,N_2008);
or U2225 (N_2225,N_2053,N_2105);
and U2226 (N_2226,N_2025,N_2103);
nand U2227 (N_2227,N_2170,N_2143);
xnor U2228 (N_2228,N_2079,N_2003);
and U2229 (N_2229,N_2128,N_2107);
and U2230 (N_2230,N_2011,N_2006);
and U2231 (N_2231,N_2189,N_2185);
nor U2232 (N_2232,N_2131,N_2168);
or U2233 (N_2233,N_2081,N_2092);
nand U2234 (N_2234,N_2001,N_2183);
or U2235 (N_2235,N_2198,N_2159);
or U2236 (N_2236,N_2057,N_2058);
or U2237 (N_2237,N_2172,N_2123);
nor U2238 (N_2238,N_2030,N_2005);
and U2239 (N_2239,N_2163,N_2016);
nand U2240 (N_2240,N_2072,N_2178);
nand U2241 (N_2241,N_2154,N_2064);
or U2242 (N_2242,N_2147,N_2089);
or U2243 (N_2243,N_2076,N_2114);
nor U2244 (N_2244,N_2084,N_2129);
nor U2245 (N_2245,N_2096,N_2149);
or U2246 (N_2246,N_2125,N_2034);
nand U2247 (N_2247,N_2071,N_2075);
or U2248 (N_2248,N_2051,N_2121);
and U2249 (N_2249,N_2077,N_2110);
nor U2250 (N_2250,N_2193,N_2100);
nand U2251 (N_2251,N_2137,N_2047);
or U2252 (N_2252,N_2017,N_2088);
and U2253 (N_2253,N_2082,N_2028);
and U2254 (N_2254,N_2164,N_2041);
or U2255 (N_2255,N_2020,N_2007);
nand U2256 (N_2256,N_2104,N_2169);
nand U2257 (N_2257,N_2134,N_2059);
nand U2258 (N_2258,N_2037,N_2098);
and U2259 (N_2259,N_2162,N_2192);
and U2260 (N_2260,N_2176,N_2187);
nand U2261 (N_2261,N_2069,N_2109);
nand U2262 (N_2262,N_2099,N_2145);
and U2263 (N_2263,N_2130,N_2197);
nor U2264 (N_2264,N_2062,N_2046);
and U2265 (N_2265,N_2171,N_2097);
nand U2266 (N_2266,N_2018,N_2010);
nand U2267 (N_2267,N_2067,N_2184);
nand U2268 (N_2268,N_2138,N_2117);
and U2269 (N_2269,N_2055,N_2085);
or U2270 (N_2270,N_2042,N_2066);
or U2271 (N_2271,N_2153,N_2086);
or U2272 (N_2272,N_2116,N_2068);
or U2273 (N_2273,N_2124,N_2023);
and U2274 (N_2274,N_2115,N_2009);
or U2275 (N_2275,N_2056,N_2074);
nand U2276 (N_2276,N_2118,N_2158);
nand U2277 (N_2277,N_2113,N_2188);
nand U2278 (N_2278,N_2112,N_2044);
or U2279 (N_2279,N_2029,N_2087);
nand U2280 (N_2280,N_2102,N_2093);
and U2281 (N_2281,N_2177,N_2160);
and U2282 (N_2282,N_2052,N_2156);
nor U2283 (N_2283,N_2070,N_2019);
nand U2284 (N_2284,N_2014,N_2048);
and U2285 (N_2285,N_2065,N_2013);
or U2286 (N_2286,N_2111,N_2040);
nor U2287 (N_2287,N_2139,N_2095);
nand U2288 (N_2288,N_2181,N_2032);
or U2289 (N_2289,N_2122,N_2073);
or U2290 (N_2290,N_2166,N_2012);
nand U2291 (N_2291,N_2167,N_2194);
nor U2292 (N_2292,N_2155,N_2196);
and U2293 (N_2293,N_2036,N_2179);
and U2294 (N_2294,N_2043,N_2119);
or U2295 (N_2295,N_2004,N_2078);
nor U2296 (N_2296,N_2091,N_2021);
nand U2297 (N_2297,N_2173,N_2136);
or U2298 (N_2298,N_2033,N_2191);
nand U2299 (N_2299,N_2101,N_2140);
nor U2300 (N_2300,N_2191,N_2048);
nor U2301 (N_2301,N_2150,N_2056);
nand U2302 (N_2302,N_2027,N_2196);
nand U2303 (N_2303,N_2002,N_2008);
nor U2304 (N_2304,N_2146,N_2099);
nor U2305 (N_2305,N_2026,N_2117);
and U2306 (N_2306,N_2093,N_2169);
nor U2307 (N_2307,N_2177,N_2016);
nand U2308 (N_2308,N_2145,N_2078);
and U2309 (N_2309,N_2129,N_2181);
nand U2310 (N_2310,N_2109,N_2180);
nor U2311 (N_2311,N_2176,N_2191);
or U2312 (N_2312,N_2033,N_2024);
or U2313 (N_2313,N_2055,N_2128);
and U2314 (N_2314,N_2176,N_2030);
nand U2315 (N_2315,N_2017,N_2127);
nor U2316 (N_2316,N_2149,N_2025);
xor U2317 (N_2317,N_2051,N_2068);
or U2318 (N_2318,N_2127,N_2168);
nor U2319 (N_2319,N_2008,N_2035);
and U2320 (N_2320,N_2083,N_2119);
nand U2321 (N_2321,N_2180,N_2158);
or U2322 (N_2322,N_2192,N_2117);
nand U2323 (N_2323,N_2106,N_2070);
or U2324 (N_2324,N_2062,N_2112);
and U2325 (N_2325,N_2036,N_2040);
nand U2326 (N_2326,N_2089,N_2042);
nand U2327 (N_2327,N_2032,N_2034);
and U2328 (N_2328,N_2148,N_2017);
and U2329 (N_2329,N_2181,N_2012);
nor U2330 (N_2330,N_2099,N_2161);
or U2331 (N_2331,N_2062,N_2174);
or U2332 (N_2332,N_2001,N_2161);
nand U2333 (N_2333,N_2174,N_2042);
and U2334 (N_2334,N_2092,N_2096);
nand U2335 (N_2335,N_2027,N_2011);
nor U2336 (N_2336,N_2159,N_2174);
nor U2337 (N_2337,N_2133,N_2164);
and U2338 (N_2338,N_2018,N_2068);
and U2339 (N_2339,N_2171,N_2052);
or U2340 (N_2340,N_2109,N_2199);
nor U2341 (N_2341,N_2142,N_2079);
nand U2342 (N_2342,N_2168,N_2154);
and U2343 (N_2343,N_2167,N_2081);
or U2344 (N_2344,N_2148,N_2174);
and U2345 (N_2345,N_2192,N_2035);
and U2346 (N_2346,N_2181,N_2146);
nor U2347 (N_2347,N_2019,N_2057);
nand U2348 (N_2348,N_2136,N_2122);
nor U2349 (N_2349,N_2032,N_2068);
or U2350 (N_2350,N_2071,N_2022);
xnor U2351 (N_2351,N_2134,N_2136);
nand U2352 (N_2352,N_2086,N_2081);
or U2353 (N_2353,N_2182,N_2066);
nand U2354 (N_2354,N_2020,N_2169);
and U2355 (N_2355,N_2102,N_2052);
nand U2356 (N_2356,N_2115,N_2100);
or U2357 (N_2357,N_2067,N_2003);
nor U2358 (N_2358,N_2062,N_2142);
or U2359 (N_2359,N_2035,N_2177);
or U2360 (N_2360,N_2118,N_2030);
nor U2361 (N_2361,N_2177,N_2168);
nor U2362 (N_2362,N_2093,N_2149);
nand U2363 (N_2363,N_2003,N_2037);
nor U2364 (N_2364,N_2095,N_2015);
or U2365 (N_2365,N_2031,N_2036);
nand U2366 (N_2366,N_2146,N_2190);
nand U2367 (N_2367,N_2072,N_2108);
or U2368 (N_2368,N_2182,N_2167);
nor U2369 (N_2369,N_2156,N_2007);
and U2370 (N_2370,N_2190,N_2029);
nand U2371 (N_2371,N_2113,N_2069);
and U2372 (N_2372,N_2171,N_2176);
nand U2373 (N_2373,N_2059,N_2072);
nor U2374 (N_2374,N_2193,N_2123);
and U2375 (N_2375,N_2095,N_2118);
and U2376 (N_2376,N_2038,N_2177);
nand U2377 (N_2377,N_2023,N_2169);
nand U2378 (N_2378,N_2007,N_2063);
nor U2379 (N_2379,N_2148,N_2061);
nand U2380 (N_2380,N_2018,N_2066);
nor U2381 (N_2381,N_2154,N_2029);
nor U2382 (N_2382,N_2166,N_2141);
nor U2383 (N_2383,N_2195,N_2121);
nor U2384 (N_2384,N_2095,N_2129);
or U2385 (N_2385,N_2151,N_2096);
and U2386 (N_2386,N_2094,N_2095);
and U2387 (N_2387,N_2170,N_2129);
nor U2388 (N_2388,N_2174,N_2137);
nor U2389 (N_2389,N_2084,N_2067);
nor U2390 (N_2390,N_2147,N_2183);
and U2391 (N_2391,N_2036,N_2028);
nor U2392 (N_2392,N_2176,N_2072);
nand U2393 (N_2393,N_2160,N_2039);
and U2394 (N_2394,N_2024,N_2063);
nor U2395 (N_2395,N_2049,N_2014);
nand U2396 (N_2396,N_2044,N_2098);
nand U2397 (N_2397,N_2148,N_2175);
nand U2398 (N_2398,N_2180,N_2048);
nor U2399 (N_2399,N_2084,N_2190);
and U2400 (N_2400,N_2324,N_2234);
and U2401 (N_2401,N_2210,N_2290);
xor U2402 (N_2402,N_2345,N_2275);
and U2403 (N_2403,N_2328,N_2327);
nand U2404 (N_2404,N_2280,N_2362);
and U2405 (N_2405,N_2294,N_2288);
and U2406 (N_2406,N_2395,N_2273);
and U2407 (N_2407,N_2396,N_2201);
nand U2408 (N_2408,N_2238,N_2223);
or U2409 (N_2409,N_2245,N_2263);
or U2410 (N_2410,N_2231,N_2279);
nor U2411 (N_2411,N_2262,N_2265);
and U2412 (N_2412,N_2269,N_2207);
nor U2413 (N_2413,N_2364,N_2353);
or U2414 (N_2414,N_2386,N_2319);
and U2415 (N_2415,N_2249,N_2251);
and U2416 (N_2416,N_2323,N_2213);
and U2417 (N_2417,N_2233,N_2237);
and U2418 (N_2418,N_2241,N_2232);
and U2419 (N_2419,N_2369,N_2310);
nor U2420 (N_2420,N_2256,N_2217);
and U2421 (N_2421,N_2359,N_2260);
and U2422 (N_2422,N_2379,N_2295);
or U2423 (N_2423,N_2302,N_2293);
or U2424 (N_2424,N_2242,N_2202);
or U2425 (N_2425,N_2229,N_2289);
or U2426 (N_2426,N_2296,N_2322);
nand U2427 (N_2427,N_2321,N_2399);
xnor U2428 (N_2428,N_2236,N_2352);
nand U2429 (N_2429,N_2307,N_2381);
and U2430 (N_2430,N_2230,N_2305);
and U2431 (N_2431,N_2339,N_2252);
nor U2432 (N_2432,N_2246,N_2346);
nand U2433 (N_2433,N_2258,N_2375);
nor U2434 (N_2434,N_2349,N_2311);
nand U2435 (N_2435,N_2240,N_2221);
or U2436 (N_2436,N_2350,N_2378);
xnor U2437 (N_2437,N_2270,N_2373);
nand U2438 (N_2438,N_2341,N_2309);
and U2439 (N_2439,N_2392,N_2286);
or U2440 (N_2440,N_2203,N_2224);
nor U2441 (N_2441,N_2285,N_2243);
or U2442 (N_2442,N_2325,N_2371);
nand U2443 (N_2443,N_2361,N_2266);
and U2444 (N_2444,N_2344,N_2215);
nand U2445 (N_2445,N_2316,N_2209);
and U2446 (N_2446,N_2351,N_2365);
nand U2447 (N_2447,N_2254,N_2332);
and U2448 (N_2448,N_2297,N_2397);
nand U2449 (N_2449,N_2264,N_2267);
or U2450 (N_2450,N_2355,N_2383);
nand U2451 (N_2451,N_2342,N_2301);
or U2452 (N_2452,N_2206,N_2326);
nand U2453 (N_2453,N_2214,N_2387);
and U2454 (N_2454,N_2281,N_2366);
nand U2455 (N_2455,N_2368,N_2382);
nor U2456 (N_2456,N_2216,N_2261);
and U2457 (N_2457,N_2391,N_2313);
nand U2458 (N_2458,N_2314,N_2398);
or U2459 (N_2459,N_2259,N_2204);
and U2460 (N_2460,N_2300,N_2219);
or U2461 (N_2461,N_2304,N_2337);
nand U2462 (N_2462,N_2250,N_2340);
and U2463 (N_2463,N_2389,N_2222);
or U2464 (N_2464,N_2357,N_2200);
or U2465 (N_2465,N_2334,N_2348);
or U2466 (N_2466,N_2315,N_2338);
or U2467 (N_2467,N_2329,N_2211);
nand U2468 (N_2468,N_2218,N_2306);
or U2469 (N_2469,N_2303,N_2388);
and U2470 (N_2470,N_2372,N_2276);
nand U2471 (N_2471,N_2283,N_2374);
nor U2472 (N_2472,N_2298,N_2244);
nand U2473 (N_2473,N_2287,N_2292);
nor U2474 (N_2474,N_2271,N_2385);
or U2475 (N_2475,N_2308,N_2354);
and U2476 (N_2476,N_2394,N_2312);
or U2477 (N_2477,N_2335,N_2225);
or U2478 (N_2478,N_2268,N_2226);
or U2479 (N_2479,N_2277,N_2212);
or U2480 (N_2480,N_2291,N_2255);
and U2481 (N_2481,N_2333,N_2336);
and U2482 (N_2482,N_2390,N_2208);
and U2483 (N_2483,N_2393,N_2367);
nor U2484 (N_2484,N_2253,N_2228);
nand U2485 (N_2485,N_2377,N_2299);
nor U2486 (N_2486,N_2247,N_2358);
and U2487 (N_2487,N_2272,N_2257);
or U2488 (N_2488,N_2248,N_2278);
nor U2489 (N_2489,N_2360,N_2205);
nor U2490 (N_2490,N_2284,N_2384);
and U2491 (N_2491,N_2282,N_2370);
and U2492 (N_2492,N_2330,N_2318);
nor U2493 (N_2493,N_2331,N_2376);
nor U2494 (N_2494,N_2320,N_2274);
nand U2495 (N_2495,N_2220,N_2363);
or U2496 (N_2496,N_2239,N_2227);
nand U2497 (N_2497,N_2235,N_2317);
xor U2498 (N_2498,N_2343,N_2380);
nand U2499 (N_2499,N_2356,N_2347);
and U2500 (N_2500,N_2307,N_2275);
or U2501 (N_2501,N_2232,N_2251);
or U2502 (N_2502,N_2254,N_2358);
and U2503 (N_2503,N_2283,N_2345);
and U2504 (N_2504,N_2219,N_2381);
nand U2505 (N_2505,N_2284,N_2233);
or U2506 (N_2506,N_2323,N_2352);
nand U2507 (N_2507,N_2386,N_2232);
nor U2508 (N_2508,N_2265,N_2310);
or U2509 (N_2509,N_2329,N_2366);
or U2510 (N_2510,N_2237,N_2229);
nand U2511 (N_2511,N_2327,N_2366);
and U2512 (N_2512,N_2330,N_2259);
or U2513 (N_2513,N_2399,N_2330);
and U2514 (N_2514,N_2228,N_2393);
nand U2515 (N_2515,N_2200,N_2372);
or U2516 (N_2516,N_2388,N_2336);
nor U2517 (N_2517,N_2234,N_2327);
nor U2518 (N_2518,N_2322,N_2278);
nor U2519 (N_2519,N_2298,N_2275);
and U2520 (N_2520,N_2268,N_2329);
nand U2521 (N_2521,N_2267,N_2221);
nor U2522 (N_2522,N_2261,N_2218);
nand U2523 (N_2523,N_2209,N_2308);
nor U2524 (N_2524,N_2232,N_2237);
and U2525 (N_2525,N_2348,N_2277);
nand U2526 (N_2526,N_2214,N_2264);
and U2527 (N_2527,N_2348,N_2378);
nand U2528 (N_2528,N_2388,N_2276);
and U2529 (N_2529,N_2375,N_2272);
or U2530 (N_2530,N_2383,N_2309);
and U2531 (N_2531,N_2277,N_2268);
nor U2532 (N_2532,N_2315,N_2248);
nor U2533 (N_2533,N_2355,N_2215);
nand U2534 (N_2534,N_2358,N_2375);
nand U2535 (N_2535,N_2202,N_2259);
and U2536 (N_2536,N_2368,N_2206);
and U2537 (N_2537,N_2368,N_2251);
and U2538 (N_2538,N_2346,N_2226);
or U2539 (N_2539,N_2336,N_2233);
and U2540 (N_2540,N_2272,N_2254);
nand U2541 (N_2541,N_2385,N_2359);
or U2542 (N_2542,N_2389,N_2379);
nor U2543 (N_2543,N_2377,N_2290);
and U2544 (N_2544,N_2245,N_2200);
and U2545 (N_2545,N_2259,N_2205);
and U2546 (N_2546,N_2367,N_2279);
nand U2547 (N_2547,N_2379,N_2267);
xor U2548 (N_2548,N_2395,N_2366);
nand U2549 (N_2549,N_2297,N_2237);
nand U2550 (N_2550,N_2248,N_2394);
and U2551 (N_2551,N_2274,N_2386);
or U2552 (N_2552,N_2248,N_2204);
or U2553 (N_2553,N_2278,N_2330);
or U2554 (N_2554,N_2384,N_2355);
nor U2555 (N_2555,N_2240,N_2332);
nand U2556 (N_2556,N_2352,N_2376);
and U2557 (N_2557,N_2378,N_2233);
or U2558 (N_2558,N_2365,N_2332);
nor U2559 (N_2559,N_2342,N_2362);
nand U2560 (N_2560,N_2328,N_2248);
nand U2561 (N_2561,N_2385,N_2365);
and U2562 (N_2562,N_2260,N_2223);
nand U2563 (N_2563,N_2207,N_2302);
nor U2564 (N_2564,N_2328,N_2307);
or U2565 (N_2565,N_2314,N_2274);
or U2566 (N_2566,N_2341,N_2262);
nor U2567 (N_2567,N_2287,N_2371);
nand U2568 (N_2568,N_2299,N_2396);
and U2569 (N_2569,N_2244,N_2247);
nand U2570 (N_2570,N_2230,N_2326);
or U2571 (N_2571,N_2220,N_2261);
nand U2572 (N_2572,N_2310,N_2256);
and U2573 (N_2573,N_2202,N_2296);
and U2574 (N_2574,N_2341,N_2300);
or U2575 (N_2575,N_2254,N_2383);
nand U2576 (N_2576,N_2216,N_2369);
or U2577 (N_2577,N_2304,N_2294);
and U2578 (N_2578,N_2209,N_2312);
nand U2579 (N_2579,N_2378,N_2284);
or U2580 (N_2580,N_2331,N_2287);
nand U2581 (N_2581,N_2244,N_2213);
and U2582 (N_2582,N_2340,N_2350);
or U2583 (N_2583,N_2395,N_2334);
and U2584 (N_2584,N_2378,N_2326);
and U2585 (N_2585,N_2276,N_2259);
or U2586 (N_2586,N_2371,N_2395);
or U2587 (N_2587,N_2236,N_2237);
and U2588 (N_2588,N_2299,N_2204);
xnor U2589 (N_2589,N_2209,N_2260);
nand U2590 (N_2590,N_2246,N_2283);
nor U2591 (N_2591,N_2286,N_2395);
nor U2592 (N_2592,N_2249,N_2372);
or U2593 (N_2593,N_2325,N_2379);
or U2594 (N_2594,N_2296,N_2301);
nand U2595 (N_2595,N_2313,N_2283);
nor U2596 (N_2596,N_2214,N_2272);
nor U2597 (N_2597,N_2261,N_2341);
or U2598 (N_2598,N_2343,N_2201);
and U2599 (N_2599,N_2269,N_2245);
nand U2600 (N_2600,N_2531,N_2413);
and U2601 (N_2601,N_2458,N_2461);
nand U2602 (N_2602,N_2479,N_2598);
and U2603 (N_2603,N_2572,N_2450);
nor U2604 (N_2604,N_2564,N_2555);
nand U2605 (N_2605,N_2596,N_2520);
and U2606 (N_2606,N_2421,N_2501);
or U2607 (N_2607,N_2467,N_2484);
and U2608 (N_2608,N_2430,N_2474);
or U2609 (N_2609,N_2448,N_2457);
and U2610 (N_2610,N_2595,N_2575);
nor U2611 (N_2611,N_2422,N_2464);
nand U2612 (N_2612,N_2489,N_2497);
nand U2613 (N_2613,N_2434,N_2540);
or U2614 (N_2614,N_2488,N_2469);
and U2615 (N_2615,N_2560,N_2447);
and U2616 (N_2616,N_2411,N_2512);
or U2617 (N_2617,N_2557,N_2569);
or U2618 (N_2618,N_2437,N_2582);
nor U2619 (N_2619,N_2403,N_2427);
or U2620 (N_2620,N_2528,N_2571);
and U2621 (N_2621,N_2420,N_2452);
or U2622 (N_2622,N_2505,N_2473);
and U2623 (N_2623,N_2532,N_2435);
and U2624 (N_2624,N_2521,N_2502);
nand U2625 (N_2625,N_2405,N_2547);
xor U2626 (N_2626,N_2466,N_2591);
and U2627 (N_2627,N_2406,N_2481);
nor U2628 (N_2628,N_2593,N_2523);
xnor U2629 (N_2629,N_2424,N_2537);
nor U2630 (N_2630,N_2415,N_2476);
or U2631 (N_2631,N_2419,N_2409);
nand U2632 (N_2632,N_2412,N_2443);
and U2633 (N_2633,N_2556,N_2562);
or U2634 (N_2634,N_2518,N_2599);
or U2635 (N_2635,N_2465,N_2519);
nor U2636 (N_2636,N_2579,N_2586);
and U2637 (N_2637,N_2529,N_2553);
nand U2638 (N_2638,N_2533,N_2515);
and U2639 (N_2639,N_2574,N_2590);
or U2640 (N_2640,N_2468,N_2576);
and U2641 (N_2641,N_2485,N_2459);
and U2642 (N_2642,N_2456,N_2548);
nor U2643 (N_2643,N_2490,N_2581);
or U2644 (N_2644,N_2508,N_2472);
nor U2645 (N_2645,N_2417,N_2538);
or U2646 (N_2646,N_2402,N_2425);
or U2647 (N_2647,N_2525,N_2580);
and U2648 (N_2648,N_2462,N_2517);
nor U2649 (N_2649,N_2433,N_2597);
and U2650 (N_2650,N_2463,N_2573);
or U2651 (N_2651,N_2535,N_2483);
nand U2652 (N_2652,N_2480,N_2565);
or U2653 (N_2653,N_2426,N_2583);
nor U2654 (N_2654,N_2549,N_2500);
nor U2655 (N_2655,N_2559,N_2416);
nand U2656 (N_2656,N_2563,N_2527);
or U2657 (N_2657,N_2453,N_2509);
and U2658 (N_2658,N_2552,N_2478);
nand U2659 (N_2659,N_2541,N_2514);
or U2660 (N_2660,N_2445,N_2455);
nand U2661 (N_2661,N_2460,N_2585);
and U2662 (N_2662,N_2539,N_2431);
nor U2663 (N_2663,N_2534,N_2516);
and U2664 (N_2664,N_2470,N_2438);
nand U2665 (N_2665,N_2471,N_2545);
and U2666 (N_2666,N_2584,N_2400);
and U2667 (N_2667,N_2594,N_2546);
nand U2668 (N_2668,N_2578,N_2446);
or U2669 (N_2669,N_2410,N_2414);
or U2670 (N_2670,N_2404,N_2429);
and U2671 (N_2671,N_2522,N_2492);
or U2672 (N_2672,N_2401,N_2442);
xor U2673 (N_2673,N_2499,N_2524);
nand U2674 (N_2674,N_2566,N_2588);
and U2675 (N_2675,N_2526,N_2506);
or U2676 (N_2676,N_2589,N_2475);
or U2677 (N_2677,N_2408,N_2592);
nor U2678 (N_2678,N_2454,N_2543);
and U2679 (N_2679,N_2551,N_2503);
and U2680 (N_2680,N_2495,N_2504);
nor U2681 (N_2681,N_2407,N_2428);
or U2682 (N_2682,N_2439,N_2510);
nor U2683 (N_2683,N_2494,N_2570);
or U2684 (N_2684,N_2513,N_2491);
nand U2685 (N_2685,N_2558,N_2567);
or U2686 (N_2686,N_2493,N_2440);
nor U2687 (N_2687,N_2441,N_2561);
nor U2688 (N_2688,N_2542,N_2577);
and U2689 (N_2689,N_2550,N_2496);
nand U2690 (N_2690,N_2487,N_2449);
nor U2691 (N_2691,N_2436,N_2423);
nand U2692 (N_2692,N_2418,N_2477);
or U2693 (N_2693,N_2486,N_2544);
nor U2694 (N_2694,N_2587,N_2482);
nor U2695 (N_2695,N_2511,N_2451);
and U2696 (N_2696,N_2568,N_2507);
nor U2697 (N_2697,N_2554,N_2536);
or U2698 (N_2698,N_2498,N_2432);
nand U2699 (N_2699,N_2530,N_2444);
nand U2700 (N_2700,N_2407,N_2409);
nor U2701 (N_2701,N_2512,N_2518);
nor U2702 (N_2702,N_2509,N_2589);
nand U2703 (N_2703,N_2434,N_2534);
and U2704 (N_2704,N_2503,N_2580);
nor U2705 (N_2705,N_2567,N_2446);
nand U2706 (N_2706,N_2450,N_2499);
nor U2707 (N_2707,N_2405,N_2470);
and U2708 (N_2708,N_2413,N_2475);
or U2709 (N_2709,N_2532,N_2459);
nor U2710 (N_2710,N_2586,N_2581);
and U2711 (N_2711,N_2485,N_2598);
nor U2712 (N_2712,N_2526,N_2580);
and U2713 (N_2713,N_2522,N_2578);
and U2714 (N_2714,N_2451,N_2464);
or U2715 (N_2715,N_2482,N_2409);
nand U2716 (N_2716,N_2400,N_2563);
nand U2717 (N_2717,N_2522,N_2403);
nor U2718 (N_2718,N_2523,N_2518);
xor U2719 (N_2719,N_2546,N_2579);
and U2720 (N_2720,N_2457,N_2492);
nand U2721 (N_2721,N_2445,N_2518);
nor U2722 (N_2722,N_2447,N_2481);
nand U2723 (N_2723,N_2457,N_2580);
nand U2724 (N_2724,N_2487,N_2521);
nor U2725 (N_2725,N_2570,N_2451);
or U2726 (N_2726,N_2552,N_2446);
nand U2727 (N_2727,N_2473,N_2403);
nand U2728 (N_2728,N_2573,N_2445);
nor U2729 (N_2729,N_2596,N_2563);
or U2730 (N_2730,N_2571,N_2578);
or U2731 (N_2731,N_2440,N_2425);
and U2732 (N_2732,N_2443,N_2599);
or U2733 (N_2733,N_2520,N_2527);
or U2734 (N_2734,N_2565,N_2580);
and U2735 (N_2735,N_2501,N_2579);
nor U2736 (N_2736,N_2592,N_2407);
and U2737 (N_2737,N_2485,N_2458);
and U2738 (N_2738,N_2409,N_2527);
nand U2739 (N_2739,N_2518,N_2544);
nor U2740 (N_2740,N_2412,N_2521);
and U2741 (N_2741,N_2453,N_2431);
or U2742 (N_2742,N_2419,N_2581);
nand U2743 (N_2743,N_2551,N_2432);
nor U2744 (N_2744,N_2435,N_2414);
nor U2745 (N_2745,N_2537,N_2538);
or U2746 (N_2746,N_2547,N_2482);
nor U2747 (N_2747,N_2453,N_2430);
and U2748 (N_2748,N_2551,N_2508);
nor U2749 (N_2749,N_2450,N_2466);
nand U2750 (N_2750,N_2485,N_2515);
nand U2751 (N_2751,N_2433,N_2468);
and U2752 (N_2752,N_2527,N_2464);
and U2753 (N_2753,N_2432,N_2452);
nand U2754 (N_2754,N_2414,N_2594);
and U2755 (N_2755,N_2503,N_2418);
or U2756 (N_2756,N_2499,N_2573);
and U2757 (N_2757,N_2597,N_2437);
nor U2758 (N_2758,N_2540,N_2415);
nor U2759 (N_2759,N_2597,N_2444);
or U2760 (N_2760,N_2594,N_2576);
and U2761 (N_2761,N_2560,N_2490);
or U2762 (N_2762,N_2449,N_2454);
and U2763 (N_2763,N_2419,N_2445);
or U2764 (N_2764,N_2402,N_2405);
and U2765 (N_2765,N_2543,N_2513);
and U2766 (N_2766,N_2583,N_2455);
and U2767 (N_2767,N_2442,N_2592);
or U2768 (N_2768,N_2428,N_2531);
nor U2769 (N_2769,N_2540,N_2559);
and U2770 (N_2770,N_2475,N_2545);
or U2771 (N_2771,N_2530,N_2503);
xnor U2772 (N_2772,N_2458,N_2430);
nor U2773 (N_2773,N_2463,N_2539);
xnor U2774 (N_2774,N_2467,N_2518);
and U2775 (N_2775,N_2594,N_2577);
and U2776 (N_2776,N_2551,N_2402);
nor U2777 (N_2777,N_2580,N_2559);
or U2778 (N_2778,N_2597,N_2473);
or U2779 (N_2779,N_2484,N_2571);
nand U2780 (N_2780,N_2513,N_2507);
or U2781 (N_2781,N_2469,N_2443);
and U2782 (N_2782,N_2447,N_2599);
nor U2783 (N_2783,N_2474,N_2426);
nand U2784 (N_2784,N_2446,N_2599);
and U2785 (N_2785,N_2520,N_2588);
or U2786 (N_2786,N_2544,N_2422);
nand U2787 (N_2787,N_2532,N_2450);
or U2788 (N_2788,N_2426,N_2499);
nand U2789 (N_2789,N_2459,N_2594);
or U2790 (N_2790,N_2523,N_2528);
and U2791 (N_2791,N_2417,N_2435);
nor U2792 (N_2792,N_2493,N_2513);
nand U2793 (N_2793,N_2518,N_2462);
nor U2794 (N_2794,N_2520,N_2503);
and U2795 (N_2795,N_2448,N_2523);
nor U2796 (N_2796,N_2551,N_2524);
nand U2797 (N_2797,N_2470,N_2532);
nand U2798 (N_2798,N_2413,N_2577);
nand U2799 (N_2799,N_2430,N_2426);
nand U2800 (N_2800,N_2629,N_2795);
and U2801 (N_2801,N_2641,N_2672);
or U2802 (N_2802,N_2745,N_2627);
and U2803 (N_2803,N_2716,N_2642);
nand U2804 (N_2804,N_2690,N_2653);
or U2805 (N_2805,N_2602,N_2604);
nor U2806 (N_2806,N_2778,N_2770);
or U2807 (N_2807,N_2717,N_2676);
nand U2808 (N_2808,N_2726,N_2668);
or U2809 (N_2809,N_2677,N_2622);
and U2810 (N_2810,N_2774,N_2789);
and U2811 (N_2811,N_2709,N_2648);
nor U2812 (N_2812,N_2740,N_2634);
and U2813 (N_2813,N_2727,N_2760);
and U2814 (N_2814,N_2744,N_2776);
and U2815 (N_2815,N_2759,N_2763);
and U2816 (N_2816,N_2714,N_2682);
and U2817 (N_2817,N_2781,N_2688);
or U2818 (N_2818,N_2769,N_2616);
and U2819 (N_2819,N_2601,N_2669);
or U2820 (N_2820,N_2683,N_2638);
and U2821 (N_2821,N_2606,N_2700);
nand U2822 (N_2822,N_2633,N_2645);
nand U2823 (N_2823,N_2733,N_2628);
nand U2824 (N_2824,N_2703,N_2773);
and U2825 (N_2825,N_2617,N_2724);
nand U2826 (N_2826,N_2687,N_2783);
or U2827 (N_2827,N_2710,N_2663);
nor U2828 (N_2828,N_2654,N_2610);
nor U2829 (N_2829,N_2649,N_2799);
or U2830 (N_2830,N_2766,N_2785);
and U2831 (N_2831,N_2751,N_2664);
nand U2832 (N_2832,N_2779,N_2630);
xnor U2833 (N_2833,N_2608,N_2678);
nand U2834 (N_2834,N_2704,N_2739);
or U2835 (N_2835,N_2637,N_2711);
nor U2836 (N_2836,N_2666,N_2758);
and U2837 (N_2837,N_2671,N_2775);
nor U2838 (N_2838,N_2721,N_2761);
nand U2839 (N_2839,N_2656,N_2743);
and U2840 (N_2840,N_2600,N_2796);
nand U2841 (N_2841,N_2715,N_2749);
or U2842 (N_2842,N_2702,N_2732);
nor U2843 (N_2843,N_2765,N_2662);
or U2844 (N_2844,N_2680,N_2786);
nor U2845 (N_2845,N_2691,N_2772);
and U2846 (N_2846,N_2698,N_2718);
nand U2847 (N_2847,N_2607,N_2706);
or U2848 (N_2848,N_2791,N_2712);
and U2849 (N_2849,N_2767,N_2603);
or U2850 (N_2850,N_2699,N_2614);
nand U2851 (N_2851,N_2755,N_2665);
or U2852 (N_2852,N_2696,N_2675);
nand U2853 (N_2853,N_2756,N_2693);
or U2854 (N_2854,N_2753,N_2626);
and U2855 (N_2855,N_2750,N_2788);
and U2856 (N_2856,N_2613,N_2636);
and U2857 (N_2857,N_2742,N_2764);
nor U2858 (N_2858,N_2708,N_2689);
or U2859 (N_2859,N_2797,N_2748);
and U2860 (N_2860,N_2635,N_2639);
or U2861 (N_2861,N_2787,N_2620);
and U2862 (N_2862,N_2728,N_2734);
nand U2863 (N_2863,N_2762,N_2657);
nand U2864 (N_2864,N_2771,N_2793);
and U2865 (N_2865,N_2650,N_2659);
nand U2866 (N_2866,N_2674,N_2652);
nand U2867 (N_2867,N_2679,N_2757);
and U2868 (N_2868,N_2692,N_2735);
or U2869 (N_2869,N_2655,N_2660);
and U2870 (N_2870,N_2782,N_2720);
or U2871 (N_2871,N_2752,N_2792);
nand U2872 (N_2872,N_2612,N_2694);
and U2873 (N_2873,N_2673,N_2661);
and U2874 (N_2874,N_2798,N_2605);
and U2875 (N_2875,N_2777,N_2646);
and U2876 (N_2876,N_2618,N_2651);
and U2877 (N_2877,N_2707,N_2701);
nor U2878 (N_2878,N_2737,N_2609);
and U2879 (N_2879,N_2621,N_2623);
nor U2880 (N_2880,N_2611,N_2624);
nand U2881 (N_2881,N_2725,N_2731);
nor U2882 (N_2882,N_2615,N_2741);
nand U2883 (N_2883,N_2730,N_2729);
nor U2884 (N_2884,N_2768,N_2738);
and U2885 (N_2885,N_2670,N_2794);
nand U2886 (N_2886,N_2705,N_2647);
and U2887 (N_2887,N_2685,N_2658);
nor U2888 (N_2888,N_2643,N_2722);
and U2889 (N_2889,N_2681,N_2625);
nand U2890 (N_2890,N_2695,N_2747);
nand U2891 (N_2891,N_2644,N_2640);
or U2892 (N_2892,N_2736,N_2619);
and U2893 (N_2893,N_2780,N_2684);
nor U2894 (N_2894,N_2686,N_2790);
nand U2895 (N_2895,N_2746,N_2723);
nand U2896 (N_2896,N_2784,N_2719);
or U2897 (N_2897,N_2667,N_2697);
and U2898 (N_2898,N_2754,N_2713);
and U2899 (N_2899,N_2631,N_2632);
nand U2900 (N_2900,N_2795,N_2646);
and U2901 (N_2901,N_2786,N_2647);
nand U2902 (N_2902,N_2751,N_2790);
nand U2903 (N_2903,N_2728,N_2660);
nand U2904 (N_2904,N_2705,N_2648);
nor U2905 (N_2905,N_2678,N_2626);
nor U2906 (N_2906,N_2624,N_2643);
nor U2907 (N_2907,N_2679,N_2776);
or U2908 (N_2908,N_2785,N_2670);
nand U2909 (N_2909,N_2621,N_2729);
or U2910 (N_2910,N_2646,N_2782);
and U2911 (N_2911,N_2637,N_2792);
nand U2912 (N_2912,N_2778,N_2668);
and U2913 (N_2913,N_2742,N_2605);
or U2914 (N_2914,N_2774,N_2706);
or U2915 (N_2915,N_2753,N_2670);
or U2916 (N_2916,N_2783,N_2727);
and U2917 (N_2917,N_2688,N_2701);
nand U2918 (N_2918,N_2769,N_2632);
and U2919 (N_2919,N_2736,N_2704);
nor U2920 (N_2920,N_2735,N_2717);
or U2921 (N_2921,N_2639,N_2720);
nand U2922 (N_2922,N_2628,N_2763);
or U2923 (N_2923,N_2718,N_2760);
nor U2924 (N_2924,N_2736,N_2728);
nand U2925 (N_2925,N_2648,N_2638);
nand U2926 (N_2926,N_2636,N_2687);
nor U2927 (N_2927,N_2682,N_2789);
nand U2928 (N_2928,N_2610,N_2639);
nand U2929 (N_2929,N_2608,N_2793);
nand U2930 (N_2930,N_2756,N_2677);
nor U2931 (N_2931,N_2793,N_2798);
nor U2932 (N_2932,N_2799,N_2680);
nand U2933 (N_2933,N_2630,N_2601);
nand U2934 (N_2934,N_2758,N_2724);
and U2935 (N_2935,N_2662,N_2631);
nand U2936 (N_2936,N_2637,N_2744);
nor U2937 (N_2937,N_2718,N_2659);
nor U2938 (N_2938,N_2758,N_2675);
nand U2939 (N_2939,N_2789,N_2686);
nor U2940 (N_2940,N_2771,N_2644);
nand U2941 (N_2941,N_2724,N_2629);
nand U2942 (N_2942,N_2763,N_2743);
nor U2943 (N_2943,N_2781,N_2699);
nor U2944 (N_2944,N_2697,N_2712);
or U2945 (N_2945,N_2640,N_2698);
nor U2946 (N_2946,N_2705,N_2738);
or U2947 (N_2947,N_2610,N_2700);
or U2948 (N_2948,N_2709,N_2743);
and U2949 (N_2949,N_2751,N_2665);
nor U2950 (N_2950,N_2719,N_2736);
nor U2951 (N_2951,N_2778,N_2764);
or U2952 (N_2952,N_2636,N_2609);
and U2953 (N_2953,N_2629,N_2641);
or U2954 (N_2954,N_2780,N_2735);
and U2955 (N_2955,N_2675,N_2630);
nand U2956 (N_2956,N_2705,N_2788);
nand U2957 (N_2957,N_2644,N_2739);
nand U2958 (N_2958,N_2602,N_2645);
and U2959 (N_2959,N_2765,N_2633);
nor U2960 (N_2960,N_2745,N_2769);
nand U2961 (N_2961,N_2725,N_2746);
nor U2962 (N_2962,N_2734,N_2721);
nor U2963 (N_2963,N_2688,N_2783);
nor U2964 (N_2964,N_2629,N_2706);
and U2965 (N_2965,N_2700,N_2618);
and U2966 (N_2966,N_2756,N_2772);
or U2967 (N_2967,N_2705,N_2704);
and U2968 (N_2968,N_2689,N_2784);
nor U2969 (N_2969,N_2755,N_2606);
nand U2970 (N_2970,N_2630,N_2609);
nor U2971 (N_2971,N_2713,N_2680);
nand U2972 (N_2972,N_2662,N_2720);
and U2973 (N_2973,N_2635,N_2630);
nor U2974 (N_2974,N_2722,N_2617);
nor U2975 (N_2975,N_2769,N_2799);
and U2976 (N_2976,N_2690,N_2677);
or U2977 (N_2977,N_2636,N_2657);
nand U2978 (N_2978,N_2710,N_2771);
or U2979 (N_2979,N_2667,N_2636);
or U2980 (N_2980,N_2795,N_2710);
nand U2981 (N_2981,N_2644,N_2687);
nand U2982 (N_2982,N_2680,N_2774);
and U2983 (N_2983,N_2762,N_2724);
nand U2984 (N_2984,N_2732,N_2673);
nor U2985 (N_2985,N_2722,N_2759);
or U2986 (N_2986,N_2660,N_2760);
nand U2987 (N_2987,N_2786,N_2727);
nor U2988 (N_2988,N_2604,N_2792);
nand U2989 (N_2989,N_2680,N_2691);
and U2990 (N_2990,N_2682,N_2683);
nor U2991 (N_2991,N_2764,N_2684);
nand U2992 (N_2992,N_2696,N_2635);
nor U2993 (N_2993,N_2686,N_2717);
or U2994 (N_2994,N_2754,N_2785);
and U2995 (N_2995,N_2768,N_2625);
or U2996 (N_2996,N_2662,N_2725);
or U2997 (N_2997,N_2762,N_2743);
or U2998 (N_2998,N_2647,N_2728);
and U2999 (N_2999,N_2760,N_2652);
nor U3000 (N_3000,N_2942,N_2850);
or U3001 (N_3001,N_2933,N_2853);
and U3002 (N_3002,N_2924,N_2967);
nand U3003 (N_3003,N_2875,N_2886);
and U3004 (N_3004,N_2815,N_2894);
nand U3005 (N_3005,N_2876,N_2839);
nor U3006 (N_3006,N_2874,N_2871);
nand U3007 (N_3007,N_2873,N_2964);
nor U3008 (N_3008,N_2938,N_2981);
nor U3009 (N_3009,N_2996,N_2891);
or U3010 (N_3010,N_2945,N_2818);
nand U3011 (N_3011,N_2977,N_2954);
and U3012 (N_3012,N_2937,N_2855);
or U3013 (N_3013,N_2805,N_2892);
or U3014 (N_3014,N_2987,N_2923);
nand U3015 (N_3015,N_2903,N_2939);
nand U3016 (N_3016,N_2951,N_2819);
nor U3017 (N_3017,N_2866,N_2861);
or U3018 (N_3018,N_2847,N_2989);
and U3019 (N_3019,N_2864,N_2829);
and U3020 (N_3020,N_2925,N_2856);
nand U3021 (N_3021,N_2956,N_2965);
nand U3022 (N_3022,N_2851,N_2978);
and U3023 (N_3023,N_2960,N_2994);
and U3024 (N_3024,N_2830,N_2804);
or U3025 (N_3025,N_2880,N_2838);
xor U3026 (N_3026,N_2801,N_2976);
nand U3027 (N_3027,N_2911,N_2917);
nor U3028 (N_3028,N_2859,N_2950);
nor U3029 (N_3029,N_2966,N_2803);
and U3030 (N_3030,N_2953,N_2835);
or U3031 (N_3031,N_2910,N_2958);
nand U3032 (N_3032,N_2833,N_2800);
nor U3033 (N_3033,N_2992,N_2814);
or U3034 (N_3034,N_2932,N_2905);
or U3035 (N_3035,N_2808,N_2899);
and U3036 (N_3036,N_2837,N_2869);
or U3037 (N_3037,N_2972,N_2918);
or U3038 (N_3038,N_2935,N_2936);
nor U3039 (N_3039,N_2995,N_2900);
and U3040 (N_3040,N_2840,N_2926);
or U3041 (N_3041,N_2922,N_2811);
or U3042 (N_3042,N_2947,N_2946);
nor U3043 (N_3043,N_2895,N_2969);
or U3044 (N_3044,N_2963,N_2844);
or U3045 (N_3045,N_2944,N_2898);
nand U3046 (N_3046,N_2821,N_2885);
nand U3047 (N_3047,N_2893,N_2842);
nand U3048 (N_3048,N_2998,N_2883);
or U3049 (N_3049,N_2881,N_2948);
and U3050 (N_3050,N_2985,N_2897);
nor U3051 (N_3051,N_2809,N_2862);
nor U3052 (N_3052,N_2857,N_2968);
nor U3053 (N_3053,N_2984,N_2979);
nand U3054 (N_3054,N_2882,N_2986);
or U3055 (N_3055,N_2826,N_2955);
and U3056 (N_3056,N_2878,N_2823);
nand U3057 (N_3057,N_2832,N_2999);
or U3058 (N_3058,N_2971,N_2975);
nor U3059 (N_3059,N_2993,N_2970);
nor U3060 (N_3060,N_2887,N_2959);
and U3061 (N_3061,N_2843,N_2820);
nor U3062 (N_3062,N_2879,N_2921);
nor U3063 (N_3063,N_2845,N_2863);
nand U3064 (N_3064,N_2848,N_2824);
and U3065 (N_3065,N_2904,N_2908);
nor U3066 (N_3066,N_2974,N_2827);
nand U3067 (N_3067,N_2816,N_2867);
nand U3068 (N_3068,N_2930,N_2907);
and U3069 (N_3069,N_2961,N_2884);
or U3070 (N_3070,N_2822,N_2929);
and U3071 (N_3071,N_2849,N_2983);
nor U3072 (N_3072,N_2872,N_2825);
or U3073 (N_3073,N_2877,N_2828);
nand U3074 (N_3074,N_2901,N_2906);
and U3075 (N_3075,N_2988,N_2860);
and U3076 (N_3076,N_2991,N_2831);
nor U3077 (N_3077,N_2914,N_2817);
nand U3078 (N_3078,N_2806,N_2865);
nand U3079 (N_3079,N_2949,N_2802);
or U3080 (N_3080,N_2957,N_2931);
nand U3081 (N_3081,N_2927,N_2813);
xor U3082 (N_3082,N_2896,N_2997);
nand U3083 (N_3083,N_2812,N_2928);
and U3084 (N_3084,N_2919,N_2952);
and U3085 (N_3085,N_2807,N_2890);
or U3086 (N_3086,N_2934,N_2889);
or U3087 (N_3087,N_2912,N_2870);
and U3088 (N_3088,N_2973,N_2915);
nor U3089 (N_3089,N_2810,N_2888);
nor U3090 (N_3090,N_2980,N_2920);
and U3091 (N_3091,N_2834,N_2990);
and U3092 (N_3092,N_2841,N_2846);
or U3093 (N_3093,N_2852,N_2940);
nand U3094 (N_3094,N_2836,N_2909);
or U3095 (N_3095,N_2854,N_2943);
or U3096 (N_3096,N_2941,N_2868);
or U3097 (N_3097,N_2913,N_2902);
and U3098 (N_3098,N_2982,N_2916);
nand U3099 (N_3099,N_2858,N_2962);
or U3100 (N_3100,N_2983,N_2808);
nor U3101 (N_3101,N_2822,N_2983);
and U3102 (N_3102,N_2862,N_2868);
or U3103 (N_3103,N_2963,N_2981);
or U3104 (N_3104,N_2924,N_2972);
nand U3105 (N_3105,N_2886,N_2808);
and U3106 (N_3106,N_2922,N_2936);
nor U3107 (N_3107,N_2869,N_2895);
or U3108 (N_3108,N_2926,N_2910);
nand U3109 (N_3109,N_2840,N_2850);
nand U3110 (N_3110,N_2870,N_2839);
or U3111 (N_3111,N_2875,N_2896);
nor U3112 (N_3112,N_2861,N_2857);
nor U3113 (N_3113,N_2925,N_2931);
nor U3114 (N_3114,N_2938,N_2952);
nand U3115 (N_3115,N_2803,N_2837);
and U3116 (N_3116,N_2812,N_2951);
and U3117 (N_3117,N_2914,N_2836);
nor U3118 (N_3118,N_2836,N_2882);
or U3119 (N_3119,N_2838,N_2834);
or U3120 (N_3120,N_2937,N_2966);
or U3121 (N_3121,N_2826,N_2802);
nand U3122 (N_3122,N_2804,N_2979);
or U3123 (N_3123,N_2845,N_2826);
nand U3124 (N_3124,N_2999,N_2968);
nor U3125 (N_3125,N_2889,N_2875);
nand U3126 (N_3126,N_2874,N_2999);
nand U3127 (N_3127,N_2848,N_2822);
or U3128 (N_3128,N_2981,N_2831);
and U3129 (N_3129,N_2935,N_2854);
nor U3130 (N_3130,N_2997,N_2880);
or U3131 (N_3131,N_2993,N_2998);
or U3132 (N_3132,N_2880,N_2968);
nor U3133 (N_3133,N_2974,N_2825);
or U3134 (N_3134,N_2922,N_2941);
nor U3135 (N_3135,N_2969,N_2880);
or U3136 (N_3136,N_2972,N_2937);
nand U3137 (N_3137,N_2875,N_2806);
or U3138 (N_3138,N_2881,N_2854);
nand U3139 (N_3139,N_2902,N_2820);
and U3140 (N_3140,N_2948,N_2987);
and U3141 (N_3141,N_2992,N_2869);
nand U3142 (N_3142,N_2898,N_2899);
nand U3143 (N_3143,N_2863,N_2987);
xnor U3144 (N_3144,N_2991,N_2826);
and U3145 (N_3145,N_2968,N_2817);
nand U3146 (N_3146,N_2965,N_2864);
nor U3147 (N_3147,N_2993,N_2802);
nand U3148 (N_3148,N_2902,N_2993);
and U3149 (N_3149,N_2924,N_2946);
nor U3150 (N_3150,N_2819,N_2846);
and U3151 (N_3151,N_2800,N_2952);
and U3152 (N_3152,N_2991,N_2861);
or U3153 (N_3153,N_2806,N_2828);
nand U3154 (N_3154,N_2986,N_2959);
nand U3155 (N_3155,N_2870,N_2935);
or U3156 (N_3156,N_2838,N_2905);
nand U3157 (N_3157,N_2882,N_2895);
and U3158 (N_3158,N_2818,N_2990);
and U3159 (N_3159,N_2962,N_2837);
or U3160 (N_3160,N_2887,N_2873);
nor U3161 (N_3161,N_2860,N_2836);
and U3162 (N_3162,N_2951,N_2867);
and U3163 (N_3163,N_2998,N_2882);
and U3164 (N_3164,N_2810,N_2900);
or U3165 (N_3165,N_2973,N_2855);
or U3166 (N_3166,N_2904,N_2944);
nand U3167 (N_3167,N_2841,N_2946);
and U3168 (N_3168,N_2815,N_2976);
nand U3169 (N_3169,N_2833,N_2847);
nand U3170 (N_3170,N_2910,N_2825);
nand U3171 (N_3171,N_2875,N_2853);
nor U3172 (N_3172,N_2826,N_2911);
or U3173 (N_3173,N_2828,N_2916);
or U3174 (N_3174,N_2803,N_2990);
and U3175 (N_3175,N_2880,N_2892);
nor U3176 (N_3176,N_2813,N_2856);
or U3177 (N_3177,N_2901,N_2885);
xor U3178 (N_3178,N_2910,N_2896);
nor U3179 (N_3179,N_2950,N_2984);
or U3180 (N_3180,N_2863,N_2800);
nand U3181 (N_3181,N_2810,N_2884);
nor U3182 (N_3182,N_2984,N_2976);
and U3183 (N_3183,N_2805,N_2918);
or U3184 (N_3184,N_2856,N_2844);
and U3185 (N_3185,N_2896,N_2906);
and U3186 (N_3186,N_2893,N_2895);
or U3187 (N_3187,N_2830,N_2896);
or U3188 (N_3188,N_2932,N_2859);
and U3189 (N_3189,N_2863,N_2911);
nor U3190 (N_3190,N_2980,N_2921);
and U3191 (N_3191,N_2817,N_2967);
nor U3192 (N_3192,N_2904,N_2838);
nand U3193 (N_3193,N_2849,N_2876);
and U3194 (N_3194,N_2948,N_2914);
nand U3195 (N_3195,N_2971,N_2925);
and U3196 (N_3196,N_2859,N_2968);
and U3197 (N_3197,N_2931,N_2860);
nand U3198 (N_3198,N_2975,N_2848);
nand U3199 (N_3199,N_2884,N_2990);
nor U3200 (N_3200,N_3094,N_3058);
nand U3201 (N_3201,N_3142,N_3073);
nor U3202 (N_3202,N_3081,N_3011);
or U3203 (N_3203,N_3032,N_3159);
or U3204 (N_3204,N_3119,N_3050);
nor U3205 (N_3205,N_3164,N_3095);
or U3206 (N_3206,N_3184,N_3116);
or U3207 (N_3207,N_3083,N_3173);
and U3208 (N_3208,N_3088,N_3014);
or U3209 (N_3209,N_3111,N_3177);
nor U3210 (N_3210,N_3158,N_3188);
and U3211 (N_3211,N_3074,N_3194);
nand U3212 (N_3212,N_3080,N_3037);
and U3213 (N_3213,N_3135,N_3153);
nand U3214 (N_3214,N_3065,N_3017);
nor U3215 (N_3215,N_3165,N_3055);
and U3216 (N_3216,N_3009,N_3108);
or U3217 (N_3217,N_3072,N_3033);
and U3218 (N_3218,N_3199,N_3028);
nand U3219 (N_3219,N_3040,N_3048);
nor U3220 (N_3220,N_3183,N_3043);
or U3221 (N_3221,N_3086,N_3059);
and U3222 (N_3222,N_3117,N_3105);
or U3223 (N_3223,N_3109,N_3123);
nor U3224 (N_3224,N_3044,N_3106);
and U3225 (N_3225,N_3075,N_3092);
nor U3226 (N_3226,N_3112,N_3064);
nand U3227 (N_3227,N_3013,N_3030);
or U3228 (N_3228,N_3178,N_3035);
nand U3229 (N_3229,N_3138,N_3019);
nor U3230 (N_3230,N_3039,N_3099);
and U3231 (N_3231,N_3176,N_3069);
nor U3232 (N_3232,N_3193,N_3150);
nand U3233 (N_3233,N_3031,N_3162);
or U3234 (N_3234,N_3101,N_3042);
and U3235 (N_3235,N_3053,N_3102);
and U3236 (N_3236,N_3051,N_3062);
nor U3237 (N_3237,N_3133,N_3128);
nand U3238 (N_3238,N_3190,N_3026);
nand U3239 (N_3239,N_3181,N_3169);
nand U3240 (N_3240,N_3085,N_3110);
or U3241 (N_3241,N_3021,N_3047);
nor U3242 (N_3242,N_3168,N_3146);
and U3243 (N_3243,N_3163,N_3100);
nand U3244 (N_3244,N_3152,N_3170);
nor U3245 (N_3245,N_3126,N_3096);
nand U3246 (N_3246,N_3174,N_3179);
and U3247 (N_3247,N_3036,N_3157);
and U3248 (N_3248,N_3041,N_3134);
or U3249 (N_3249,N_3196,N_3071);
and U3250 (N_3250,N_3161,N_3003);
nor U3251 (N_3251,N_3077,N_3187);
or U3252 (N_3252,N_3137,N_3001);
nor U3253 (N_3253,N_3038,N_3066);
and U3254 (N_3254,N_3049,N_3104);
or U3255 (N_3255,N_3167,N_3082);
or U3256 (N_3256,N_3129,N_3034);
nand U3257 (N_3257,N_3007,N_3068);
nor U3258 (N_3258,N_3045,N_3186);
and U3259 (N_3259,N_3022,N_3078);
and U3260 (N_3260,N_3124,N_3097);
nand U3261 (N_3261,N_3182,N_3046);
nor U3262 (N_3262,N_3018,N_3079);
and U3263 (N_3263,N_3145,N_3107);
and U3264 (N_3264,N_3144,N_3127);
or U3265 (N_3265,N_3012,N_3185);
and U3266 (N_3266,N_3091,N_3004);
or U3267 (N_3267,N_3000,N_3067);
nand U3268 (N_3268,N_3103,N_3180);
nor U3269 (N_3269,N_3155,N_3131);
nand U3270 (N_3270,N_3197,N_3115);
nand U3271 (N_3271,N_3029,N_3160);
nand U3272 (N_3272,N_3070,N_3132);
nor U3273 (N_3273,N_3052,N_3060);
nor U3274 (N_3274,N_3166,N_3192);
or U3275 (N_3275,N_3143,N_3057);
or U3276 (N_3276,N_3076,N_3139);
nand U3277 (N_3277,N_3008,N_3151);
or U3278 (N_3278,N_3148,N_3063);
or U3279 (N_3279,N_3016,N_3130);
or U3280 (N_3280,N_3084,N_3114);
or U3281 (N_3281,N_3195,N_3120);
nand U3282 (N_3282,N_3122,N_3020);
and U3283 (N_3283,N_3141,N_3113);
nand U3284 (N_3284,N_3136,N_3191);
nand U3285 (N_3285,N_3054,N_3010);
and U3286 (N_3286,N_3093,N_3140);
and U3287 (N_3287,N_3089,N_3147);
nand U3288 (N_3288,N_3121,N_3090);
or U3289 (N_3289,N_3198,N_3175);
or U3290 (N_3290,N_3024,N_3087);
nor U3291 (N_3291,N_3156,N_3002);
nand U3292 (N_3292,N_3118,N_3027);
nand U3293 (N_3293,N_3189,N_3171);
or U3294 (N_3294,N_3061,N_3005);
nor U3295 (N_3295,N_3006,N_3098);
nand U3296 (N_3296,N_3015,N_3149);
and U3297 (N_3297,N_3154,N_3023);
or U3298 (N_3298,N_3172,N_3056);
nand U3299 (N_3299,N_3125,N_3025);
or U3300 (N_3300,N_3198,N_3144);
nand U3301 (N_3301,N_3070,N_3166);
xnor U3302 (N_3302,N_3040,N_3150);
nand U3303 (N_3303,N_3082,N_3194);
nand U3304 (N_3304,N_3023,N_3014);
and U3305 (N_3305,N_3032,N_3053);
and U3306 (N_3306,N_3100,N_3055);
nand U3307 (N_3307,N_3122,N_3021);
or U3308 (N_3308,N_3027,N_3037);
and U3309 (N_3309,N_3010,N_3066);
nand U3310 (N_3310,N_3086,N_3165);
nor U3311 (N_3311,N_3093,N_3130);
nand U3312 (N_3312,N_3083,N_3080);
nand U3313 (N_3313,N_3000,N_3175);
nor U3314 (N_3314,N_3088,N_3160);
and U3315 (N_3315,N_3036,N_3071);
nand U3316 (N_3316,N_3180,N_3079);
and U3317 (N_3317,N_3183,N_3086);
nand U3318 (N_3318,N_3154,N_3065);
or U3319 (N_3319,N_3132,N_3154);
nand U3320 (N_3320,N_3149,N_3108);
nand U3321 (N_3321,N_3190,N_3104);
and U3322 (N_3322,N_3139,N_3089);
nor U3323 (N_3323,N_3187,N_3192);
and U3324 (N_3324,N_3175,N_3147);
nor U3325 (N_3325,N_3170,N_3144);
nor U3326 (N_3326,N_3101,N_3092);
or U3327 (N_3327,N_3098,N_3077);
or U3328 (N_3328,N_3040,N_3010);
and U3329 (N_3329,N_3128,N_3110);
or U3330 (N_3330,N_3075,N_3133);
or U3331 (N_3331,N_3049,N_3135);
and U3332 (N_3332,N_3168,N_3071);
or U3333 (N_3333,N_3062,N_3109);
and U3334 (N_3334,N_3006,N_3102);
or U3335 (N_3335,N_3053,N_3131);
nor U3336 (N_3336,N_3006,N_3112);
nor U3337 (N_3337,N_3099,N_3046);
nor U3338 (N_3338,N_3122,N_3117);
or U3339 (N_3339,N_3178,N_3153);
or U3340 (N_3340,N_3065,N_3196);
and U3341 (N_3341,N_3050,N_3003);
or U3342 (N_3342,N_3108,N_3052);
nor U3343 (N_3343,N_3051,N_3158);
or U3344 (N_3344,N_3072,N_3100);
and U3345 (N_3345,N_3158,N_3187);
nand U3346 (N_3346,N_3015,N_3099);
nor U3347 (N_3347,N_3036,N_3177);
and U3348 (N_3348,N_3021,N_3091);
and U3349 (N_3349,N_3069,N_3184);
and U3350 (N_3350,N_3154,N_3019);
and U3351 (N_3351,N_3166,N_3191);
nand U3352 (N_3352,N_3182,N_3161);
nand U3353 (N_3353,N_3119,N_3159);
nand U3354 (N_3354,N_3149,N_3091);
or U3355 (N_3355,N_3173,N_3124);
nand U3356 (N_3356,N_3110,N_3158);
nand U3357 (N_3357,N_3065,N_3067);
nand U3358 (N_3358,N_3135,N_3107);
nand U3359 (N_3359,N_3173,N_3053);
or U3360 (N_3360,N_3007,N_3190);
nand U3361 (N_3361,N_3165,N_3163);
and U3362 (N_3362,N_3129,N_3086);
or U3363 (N_3363,N_3153,N_3005);
and U3364 (N_3364,N_3045,N_3077);
or U3365 (N_3365,N_3033,N_3115);
and U3366 (N_3366,N_3182,N_3156);
nand U3367 (N_3367,N_3024,N_3188);
nor U3368 (N_3368,N_3123,N_3045);
and U3369 (N_3369,N_3081,N_3199);
and U3370 (N_3370,N_3037,N_3108);
or U3371 (N_3371,N_3144,N_3071);
nor U3372 (N_3372,N_3135,N_3088);
nand U3373 (N_3373,N_3123,N_3154);
nand U3374 (N_3374,N_3117,N_3138);
nand U3375 (N_3375,N_3042,N_3050);
nand U3376 (N_3376,N_3156,N_3168);
nand U3377 (N_3377,N_3034,N_3145);
or U3378 (N_3378,N_3017,N_3085);
or U3379 (N_3379,N_3177,N_3133);
or U3380 (N_3380,N_3042,N_3116);
and U3381 (N_3381,N_3082,N_3170);
nand U3382 (N_3382,N_3095,N_3105);
or U3383 (N_3383,N_3061,N_3008);
nor U3384 (N_3384,N_3179,N_3096);
nand U3385 (N_3385,N_3077,N_3159);
nand U3386 (N_3386,N_3168,N_3018);
nand U3387 (N_3387,N_3019,N_3054);
or U3388 (N_3388,N_3117,N_3135);
or U3389 (N_3389,N_3001,N_3012);
nor U3390 (N_3390,N_3021,N_3014);
and U3391 (N_3391,N_3110,N_3177);
and U3392 (N_3392,N_3100,N_3134);
nor U3393 (N_3393,N_3109,N_3128);
nor U3394 (N_3394,N_3193,N_3011);
and U3395 (N_3395,N_3120,N_3154);
nor U3396 (N_3396,N_3163,N_3130);
and U3397 (N_3397,N_3111,N_3197);
nand U3398 (N_3398,N_3159,N_3064);
and U3399 (N_3399,N_3031,N_3151);
nor U3400 (N_3400,N_3319,N_3306);
nand U3401 (N_3401,N_3211,N_3256);
nor U3402 (N_3402,N_3329,N_3212);
nand U3403 (N_3403,N_3268,N_3367);
or U3404 (N_3404,N_3361,N_3371);
and U3405 (N_3405,N_3237,N_3308);
or U3406 (N_3406,N_3249,N_3258);
and U3407 (N_3407,N_3229,N_3206);
and U3408 (N_3408,N_3382,N_3250);
and U3409 (N_3409,N_3265,N_3251);
nand U3410 (N_3410,N_3354,N_3242);
or U3411 (N_3411,N_3398,N_3321);
nor U3412 (N_3412,N_3219,N_3289);
nor U3413 (N_3413,N_3243,N_3307);
or U3414 (N_3414,N_3340,N_3297);
or U3415 (N_3415,N_3356,N_3370);
nand U3416 (N_3416,N_3223,N_3246);
nor U3417 (N_3417,N_3344,N_3314);
nor U3418 (N_3418,N_3368,N_3225);
nor U3419 (N_3419,N_3385,N_3337);
nand U3420 (N_3420,N_3362,N_3294);
nor U3421 (N_3421,N_3279,N_3214);
and U3422 (N_3422,N_3240,N_3208);
or U3423 (N_3423,N_3204,N_3280);
nand U3424 (N_3424,N_3347,N_3332);
or U3425 (N_3425,N_3239,N_3357);
nand U3426 (N_3426,N_3313,N_3376);
nand U3427 (N_3427,N_3252,N_3301);
nand U3428 (N_3428,N_3277,N_3262);
nor U3429 (N_3429,N_3325,N_3389);
nand U3430 (N_3430,N_3349,N_3202);
nand U3431 (N_3431,N_3236,N_3261);
nand U3432 (N_3432,N_3311,N_3284);
nand U3433 (N_3433,N_3318,N_3230);
or U3434 (N_3434,N_3273,N_3335);
or U3435 (N_3435,N_3247,N_3386);
xnor U3436 (N_3436,N_3355,N_3302);
nand U3437 (N_3437,N_3215,N_3231);
and U3438 (N_3438,N_3263,N_3383);
or U3439 (N_3439,N_3336,N_3377);
nor U3440 (N_3440,N_3373,N_3283);
or U3441 (N_3441,N_3266,N_3345);
and U3442 (N_3442,N_3217,N_3288);
nand U3443 (N_3443,N_3227,N_3264);
nor U3444 (N_3444,N_3369,N_3360);
nand U3445 (N_3445,N_3248,N_3365);
or U3446 (N_3446,N_3276,N_3228);
nand U3447 (N_3447,N_3224,N_3269);
nor U3448 (N_3448,N_3222,N_3327);
nand U3449 (N_3449,N_3339,N_3282);
or U3450 (N_3450,N_3320,N_3375);
nor U3451 (N_3451,N_3312,N_3203);
xnor U3452 (N_3452,N_3293,N_3226);
or U3453 (N_3453,N_3274,N_3275);
or U3454 (N_3454,N_3399,N_3333);
nand U3455 (N_3455,N_3235,N_3343);
and U3456 (N_3456,N_3322,N_3272);
nor U3457 (N_3457,N_3346,N_3392);
and U3458 (N_3458,N_3374,N_3270);
and U3459 (N_3459,N_3304,N_3380);
or U3460 (N_3460,N_3213,N_3326);
nor U3461 (N_3461,N_3358,N_3384);
and U3462 (N_3462,N_3232,N_3395);
and U3463 (N_3463,N_3364,N_3210);
or U3464 (N_3464,N_3216,N_3207);
nand U3465 (N_3465,N_3300,N_3396);
and U3466 (N_3466,N_3342,N_3220);
nand U3467 (N_3467,N_3387,N_3330);
and U3468 (N_3468,N_3244,N_3281);
xor U3469 (N_3469,N_3287,N_3218);
nor U3470 (N_3470,N_3315,N_3241);
nand U3471 (N_3471,N_3201,N_3391);
nor U3472 (N_3472,N_3394,N_3298);
nand U3473 (N_3473,N_3317,N_3352);
or U3474 (N_3474,N_3310,N_3200);
nand U3475 (N_3475,N_3234,N_3253);
nand U3476 (N_3476,N_3350,N_3233);
and U3477 (N_3477,N_3379,N_3255);
nor U3478 (N_3478,N_3397,N_3245);
nand U3479 (N_3479,N_3290,N_3324);
and U3480 (N_3480,N_3351,N_3295);
nor U3481 (N_3481,N_3388,N_3323);
nor U3482 (N_3482,N_3381,N_3285);
nor U3483 (N_3483,N_3299,N_3334);
nor U3484 (N_3484,N_3221,N_3292);
nand U3485 (N_3485,N_3359,N_3205);
nand U3486 (N_3486,N_3348,N_3291);
and U3487 (N_3487,N_3372,N_3254);
nand U3488 (N_3488,N_3209,N_3338);
nand U3489 (N_3489,N_3260,N_3309);
nand U3490 (N_3490,N_3238,N_3259);
nor U3491 (N_3491,N_3393,N_3378);
and U3492 (N_3492,N_3296,N_3353);
nor U3493 (N_3493,N_3390,N_3271);
and U3494 (N_3494,N_3303,N_3341);
or U3495 (N_3495,N_3363,N_3278);
nor U3496 (N_3496,N_3305,N_3366);
nand U3497 (N_3497,N_3257,N_3331);
nand U3498 (N_3498,N_3267,N_3328);
nor U3499 (N_3499,N_3316,N_3286);
and U3500 (N_3500,N_3320,N_3334);
and U3501 (N_3501,N_3368,N_3251);
and U3502 (N_3502,N_3349,N_3281);
or U3503 (N_3503,N_3379,N_3344);
or U3504 (N_3504,N_3389,N_3230);
nand U3505 (N_3505,N_3370,N_3357);
nand U3506 (N_3506,N_3281,N_3250);
nor U3507 (N_3507,N_3357,N_3244);
and U3508 (N_3508,N_3261,N_3243);
and U3509 (N_3509,N_3279,N_3364);
or U3510 (N_3510,N_3376,N_3319);
nor U3511 (N_3511,N_3366,N_3363);
nand U3512 (N_3512,N_3363,N_3303);
nand U3513 (N_3513,N_3366,N_3246);
or U3514 (N_3514,N_3338,N_3329);
or U3515 (N_3515,N_3285,N_3228);
or U3516 (N_3516,N_3289,N_3325);
nor U3517 (N_3517,N_3295,N_3378);
nand U3518 (N_3518,N_3245,N_3211);
nor U3519 (N_3519,N_3205,N_3312);
and U3520 (N_3520,N_3303,N_3287);
nor U3521 (N_3521,N_3221,N_3270);
nor U3522 (N_3522,N_3263,N_3221);
nand U3523 (N_3523,N_3360,N_3390);
and U3524 (N_3524,N_3347,N_3315);
and U3525 (N_3525,N_3368,N_3284);
xor U3526 (N_3526,N_3378,N_3256);
and U3527 (N_3527,N_3264,N_3369);
or U3528 (N_3528,N_3211,N_3397);
nor U3529 (N_3529,N_3324,N_3332);
nand U3530 (N_3530,N_3245,N_3322);
nand U3531 (N_3531,N_3229,N_3216);
or U3532 (N_3532,N_3399,N_3304);
nand U3533 (N_3533,N_3355,N_3305);
or U3534 (N_3534,N_3229,N_3285);
or U3535 (N_3535,N_3288,N_3282);
or U3536 (N_3536,N_3207,N_3325);
or U3537 (N_3537,N_3318,N_3287);
nand U3538 (N_3538,N_3367,N_3251);
nand U3539 (N_3539,N_3221,N_3372);
or U3540 (N_3540,N_3329,N_3213);
nor U3541 (N_3541,N_3345,N_3280);
nand U3542 (N_3542,N_3306,N_3388);
and U3543 (N_3543,N_3337,N_3322);
nand U3544 (N_3544,N_3337,N_3276);
or U3545 (N_3545,N_3226,N_3335);
and U3546 (N_3546,N_3233,N_3261);
nand U3547 (N_3547,N_3251,N_3364);
nand U3548 (N_3548,N_3296,N_3262);
nand U3549 (N_3549,N_3339,N_3280);
nand U3550 (N_3550,N_3209,N_3373);
and U3551 (N_3551,N_3333,N_3272);
nand U3552 (N_3552,N_3282,N_3251);
nor U3553 (N_3553,N_3384,N_3348);
or U3554 (N_3554,N_3276,N_3261);
nor U3555 (N_3555,N_3271,N_3384);
or U3556 (N_3556,N_3398,N_3258);
and U3557 (N_3557,N_3363,N_3393);
nand U3558 (N_3558,N_3297,N_3348);
and U3559 (N_3559,N_3312,N_3391);
and U3560 (N_3560,N_3342,N_3294);
and U3561 (N_3561,N_3330,N_3239);
and U3562 (N_3562,N_3378,N_3398);
and U3563 (N_3563,N_3259,N_3278);
nor U3564 (N_3564,N_3386,N_3384);
or U3565 (N_3565,N_3382,N_3314);
or U3566 (N_3566,N_3230,N_3258);
or U3567 (N_3567,N_3357,N_3259);
nand U3568 (N_3568,N_3363,N_3269);
nor U3569 (N_3569,N_3385,N_3227);
or U3570 (N_3570,N_3294,N_3239);
or U3571 (N_3571,N_3377,N_3359);
nand U3572 (N_3572,N_3227,N_3338);
or U3573 (N_3573,N_3285,N_3396);
nand U3574 (N_3574,N_3230,N_3365);
and U3575 (N_3575,N_3281,N_3227);
nand U3576 (N_3576,N_3305,N_3384);
nor U3577 (N_3577,N_3230,N_3310);
nor U3578 (N_3578,N_3379,N_3257);
nand U3579 (N_3579,N_3269,N_3229);
and U3580 (N_3580,N_3251,N_3296);
and U3581 (N_3581,N_3254,N_3332);
nor U3582 (N_3582,N_3337,N_3369);
nor U3583 (N_3583,N_3216,N_3260);
and U3584 (N_3584,N_3258,N_3312);
and U3585 (N_3585,N_3272,N_3394);
or U3586 (N_3586,N_3296,N_3286);
or U3587 (N_3587,N_3237,N_3389);
and U3588 (N_3588,N_3260,N_3322);
and U3589 (N_3589,N_3207,N_3300);
and U3590 (N_3590,N_3340,N_3370);
nor U3591 (N_3591,N_3345,N_3379);
or U3592 (N_3592,N_3247,N_3276);
nor U3593 (N_3593,N_3250,N_3319);
nor U3594 (N_3594,N_3359,N_3346);
or U3595 (N_3595,N_3369,N_3395);
nor U3596 (N_3596,N_3304,N_3393);
or U3597 (N_3597,N_3285,N_3220);
nand U3598 (N_3598,N_3296,N_3372);
nor U3599 (N_3599,N_3362,N_3385);
nand U3600 (N_3600,N_3505,N_3525);
nor U3601 (N_3601,N_3424,N_3415);
and U3602 (N_3602,N_3537,N_3554);
or U3603 (N_3603,N_3440,N_3592);
nor U3604 (N_3604,N_3421,N_3543);
nand U3605 (N_3605,N_3426,N_3545);
nor U3606 (N_3606,N_3599,N_3457);
or U3607 (N_3607,N_3491,N_3450);
or U3608 (N_3608,N_3578,N_3502);
nor U3609 (N_3609,N_3506,N_3559);
nor U3610 (N_3610,N_3584,N_3404);
nor U3611 (N_3611,N_3403,N_3596);
or U3612 (N_3612,N_3581,N_3494);
nand U3613 (N_3613,N_3573,N_3446);
nor U3614 (N_3614,N_3425,N_3515);
and U3615 (N_3615,N_3423,N_3516);
or U3616 (N_3616,N_3501,N_3433);
nand U3617 (N_3617,N_3513,N_3416);
and U3618 (N_3618,N_3548,N_3409);
nand U3619 (N_3619,N_3411,N_3412);
or U3620 (N_3620,N_3597,N_3406);
or U3621 (N_3621,N_3474,N_3527);
nor U3622 (N_3622,N_3488,N_3585);
nand U3623 (N_3623,N_3577,N_3514);
or U3624 (N_3624,N_3435,N_3448);
and U3625 (N_3625,N_3436,N_3495);
nor U3626 (N_3626,N_3442,N_3452);
and U3627 (N_3627,N_3571,N_3539);
and U3628 (N_3628,N_3492,N_3588);
or U3629 (N_3629,N_3430,N_3538);
and U3630 (N_3630,N_3528,N_3498);
nor U3631 (N_3631,N_3402,N_3493);
nor U3632 (N_3632,N_3487,N_3428);
nor U3633 (N_3633,N_3590,N_3437);
and U3634 (N_3634,N_3497,N_3504);
nand U3635 (N_3635,N_3458,N_3532);
nand U3636 (N_3636,N_3541,N_3467);
nand U3637 (N_3637,N_3459,N_3558);
nor U3638 (N_3638,N_3510,N_3526);
or U3639 (N_3639,N_3553,N_3564);
nor U3640 (N_3640,N_3427,N_3536);
nor U3641 (N_3641,N_3561,N_3560);
nand U3642 (N_3642,N_3464,N_3480);
nor U3643 (N_3643,N_3531,N_3562);
nor U3644 (N_3644,N_3439,N_3575);
or U3645 (N_3645,N_3441,N_3586);
nand U3646 (N_3646,N_3593,N_3552);
and U3647 (N_3647,N_3456,N_3598);
nand U3648 (N_3648,N_3566,N_3434);
nand U3649 (N_3649,N_3455,N_3414);
nor U3650 (N_3650,N_3482,N_3460);
or U3651 (N_3651,N_3582,N_3509);
and U3652 (N_3652,N_3410,N_3484);
and U3653 (N_3653,N_3529,N_3544);
and U3654 (N_3654,N_3591,N_3533);
and U3655 (N_3655,N_3438,N_3471);
and U3656 (N_3656,N_3530,N_3481);
or U3657 (N_3657,N_3469,N_3546);
and U3658 (N_3658,N_3419,N_3449);
nand U3659 (N_3659,N_3507,N_3508);
and U3660 (N_3660,N_3476,N_3549);
or U3661 (N_3661,N_3583,N_3444);
and U3662 (N_3662,N_3589,N_3555);
nand U3663 (N_3663,N_3521,N_3475);
nand U3664 (N_3664,N_3518,N_3557);
or U3665 (N_3665,N_3500,N_3477);
nand U3666 (N_3666,N_3454,N_3429);
or U3667 (N_3667,N_3468,N_3574);
nand U3668 (N_3668,N_3567,N_3473);
nor U3669 (N_3669,N_3556,N_3451);
nand U3670 (N_3670,N_3535,N_3496);
nand U3671 (N_3671,N_3453,N_3579);
nor U3672 (N_3672,N_3517,N_3540);
and U3673 (N_3673,N_3490,N_3405);
and U3674 (N_3674,N_3551,N_3580);
or U3675 (N_3675,N_3466,N_3565);
and U3676 (N_3676,N_3524,N_3511);
or U3677 (N_3677,N_3595,N_3483);
or U3678 (N_3678,N_3523,N_3443);
nor U3679 (N_3679,N_3408,N_3470);
or U3680 (N_3680,N_3568,N_3520);
nand U3681 (N_3681,N_3576,N_3570);
nor U3682 (N_3682,N_3418,N_3401);
and U3683 (N_3683,N_3542,N_3461);
nand U3684 (N_3684,N_3445,N_3547);
or U3685 (N_3685,N_3479,N_3550);
or U3686 (N_3686,N_3489,N_3465);
or U3687 (N_3687,N_3417,N_3431);
and U3688 (N_3688,N_3485,N_3400);
and U3689 (N_3689,N_3407,N_3422);
or U3690 (N_3690,N_3519,N_3594);
and U3691 (N_3691,N_3478,N_3447);
and U3692 (N_3692,N_3486,N_3499);
nand U3693 (N_3693,N_3463,N_3432);
or U3694 (N_3694,N_3472,N_3503);
nor U3695 (N_3695,N_3512,N_3563);
nor U3696 (N_3696,N_3462,N_3522);
nor U3697 (N_3697,N_3534,N_3569);
or U3698 (N_3698,N_3572,N_3587);
or U3699 (N_3699,N_3413,N_3420);
and U3700 (N_3700,N_3522,N_3548);
or U3701 (N_3701,N_3498,N_3412);
or U3702 (N_3702,N_3514,N_3427);
nor U3703 (N_3703,N_3410,N_3418);
or U3704 (N_3704,N_3458,N_3559);
or U3705 (N_3705,N_3592,N_3478);
or U3706 (N_3706,N_3515,N_3500);
nor U3707 (N_3707,N_3406,N_3551);
nand U3708 (N_3708,N_3542,N_3419);
nand U3709 (N_3709,N_3413,N_3492);
nor U3710 (N_3710,N_3581,N_3444);
nor U3711 (N_3711,N_3429,N_3406);
nand U3712 (N_3712,N_3413,N_3456);
nand U3713 (N_3713,N_3519,N_3445);
nor U3714 (N_3714,N_3544,N_3509);
nand U3715 (N_3715,N_3578,N_3539);
and U3716 (N_3716,N_3568,N_3460);
nor U3717 (N_3717,N_3566,N_3509);
or U3718 (N_3718,N_3553,N_3528);
nor U3719 (N_3719,N_3577,N_3515);
and U3720 (N_3720,N_3590,N_3498);
nand U3721 (N_3721,N_3549,N_3517);
nor U3722 (N_3722,N_3402,N_3458);
or U3723 (N_3723,N_3549,N_3587);
and U3724 (N_3724,N_3505,N_3587);
nand U3725 (N_3725,N_3552,N_3529);
and U3726 (N_3726,N_3411,N_3518);
nand U3727 (N_3727,N_3412,N_3501);
nand U3728 (N_3728,N_3573,N_3419);
or U3729 (N_3729,N_3502,N_3473);
nor U3730 (N_3730,N_3508,N_3554);
nand U3731 (N_3731,N_3525,N_3511);
and U3732 (N_3732,N_3509,N_3545);
and U3733 (N_3733,N_3439,N_3419);
or U3734 (N_3734,N_3540,N_3489);
nand U3735 (N_3735,N_3436,N_3500);
nand U3736 (N_3736,N_3491,N_3587);
or U3737 (N_3737,N_3493,N_3543);
nor U3738 (N_3738,N_3462,N_3484);
nor U3739 (N_3739,N_3545,N_3560);
and U3740 (N_3740,N_3492,N_3428);
or U3741 (N_3741,N_3447,N_3407);
or U3742 (N_3742,N_3508,N_3555);
nor U3743 (N_3743,N_3596,N_3495);
nor U3744 (N_3744,N_3598,N_3586);
and U3745 (N_3745,N_3493,N_3439);
and U3746 (N_3746,N_3581,N_3592);
and U3747 (N_3747,N_3462,N_3460);
nor U3748 (N_3748,N_3467,N_3446);
nand U3749 (N_3749,N_3433,N_3463);
or U3750 (N_3750,N_3507,N_3524);
nor U3751 (N_3751,N_3569,N_3422);
nor U3752 (N_3752,N_3481,N_3419);
nand U3753 (N_3753,N_3459,N_3556);
xor U3754 (N_3754,N_3410,N_3535);
or U3755 (N_3755,N_3541,N_3586);
nand U3756 (N_3756,N_3438,N_3460);
or U3757 (N_3757,N_3446,N_3531);
nand U3758 (N_3758,N_3520,N_3463);
and U3759 (N_3759,N_3489,N_3428);
or U3760 (N_3760,N_3538,N_3452);
and U3761 (N_3761,N_3593,N_3547);
or U3762 (N_3762,N_3589,N_3492);
or U3763 (N_3763,N_3573,N_3435);
nand U3764 (N_3764,N_3533,N_3599);
and U3765 (N_3765,N_3424,N_3490);
nor U3766 (N_3766,N_3506,N_3489);
nand U3767 (N_3767,N_3538,N_3457);
or U3768 (N_3768,N_3547,N_3468);
or U3769 (N_3769,N_3452,N_3533);
or U3770 (N_3770,N_3400,N_3566);
and U3771 (N_3771,N_3400,N_3456);
or U3772 (N_3772,N_3488,N_3443);
or U3773 (N_3773,N_3457,N_3519);
nand U3774 (N_3774,N_3562,N_3532);
or U3775 (N_3775,N_3512,N_3492);
nand U3776 (N_3776,N_3477,N_3595);
or U3777 (N_3777,N_3441,N_3446);
nor U3778 (N_3778,N_3566,N_3525);
or U3779 (N_3779,N_3574,N_3540);
nand U3780 (N_3780,N_3421,N_3506);
nor U3781 (N_3781,N_3437,N_3582);
or U3782 (N_3782,N_3400,N_3573);
and U3783 (N_3783,N_3521,N_3547);
nor U3784 (N_3784,N_3564,N_3485);
nor U3785 (N_3785,N_3596,N_3579);
nor U3786 (N_3786,N_3527,N_3558);
and U3787 (N_3787,N_3541,N_3453);
and U3788 (N_3788,N_3552,N_3433);
or U3789 (N_3789,N_3525,N_3503);
nor U3790 (N_3790,N_3426,N_3439);
nand U3791 (N_3791,N_3400,N_3538);
nor U3792 (N_3792,N_3460,N_3504);
nand U3793 (N_3793,N_3438,N_3467);
or U3794 (N_3794,N_3536,N_3437);
nor U3795 (N_3795,N_3413,N_3529);
or U3796 (N_3796,N_3553,N_3448);
nand U3797 (N_3797,N_3577,N_3457);
nand U3798 (N_3798,N_3529,N_3531);
and U3799 (N_3799,N_3542,N_3533);
nor U3800 (N_3800,N_3709,N_3736);
and U3801 (N_3801,N_3676,N_3753);
and U3802 (N_3802,N_3735,N_3724);
or U3803 (N_3803,N_3672,N_3717);
or U3804 (N_3804,N_3739,N_3690);
nand U3805 (N_3805,N_3796,N_3760);
and U3806 (N_3806,N_3726,N_3623);
nor U3807 (N_3807,N_3620,N_3614);
or U3808 (N_3808,N_3763,N_3636);
or U3809 (N_3809,N_3751,N_3689);
or U3810 (N_3810,N_3624,N_3775);
or U3811 (N_3811,N_3792,N_3698);
and U3812 (N_3812,N_3765,N_3741);
nand U3813 (N_3813,N_3706,N_3646);
nor U3814 (N_3814,N_3693,N_3779);
nand U3815 (N_3815,N_3714,N_3604);
or U3816 (N_3816,N_3766,N_3642);
nand U3817 (N_3817,N_3686,N_3795);
nand U3818 (N_3818,N_3746,N_3626);
or U3819 (N_3819,N_3794,N_3648);
nand U3820 (N_3820,N_3713,N_3667);
nand U3821 (N_3821,N_3639,N_3619);
and U3822 (N_3822,N_3680,N_3643);
or U3823 (N_3823,N_3668,N_3694);
nand U3824 (N_3824,N_3789,N_3634);
and U3825 (N_3825,N_3611,N_3749);
and U3826 (N_3826,N_3647,N_3748);
nand U3827 (N_3827,N_3652,N_3788);
or U3828 (N_3828,N_3710,N_3691);
or U3829 (N_3829,N_3768,N_3613);
or U3830 (N_3830,N_3600,N_3712);
or U3831 (N_3831,N_3752,N_3756);
nand U3832 (N_3832,N_3678,N_3778);
nand U3833 (N_3833,N_3612,N_3754);
and U3834 (N_3834,N_3675,N_3635);
nor U3835 (N_3835,N_3708,N_3727);
and U3836 (N_3836,N_3773,N_3610);
xnor U3837 (N_3837,N_3790,N_3660);
nor U3838 (N_3838,N_3637,N_3670);
nand U3839 (N_3839,N_3621,N_3605);
nand U3840 (N_3840,N_3615,N_3704);
nand U3841 (N_3841,N_3638,N_3662);
and U3842 (N_3842,N_3664,N_3697);
nand U3843 (N_3843,N_3733,N_3774);
nor U3844 (N_3844,N_3750,N_3658);
nand U3845 (N_3845,N_3742,N_3687);
nand U3846 (N_3846,N_3780,N_3718);
and U3847 (N_3847,N_3701,N_3650);
and U3848 (N_3848,N_3762,N_3761);
nand U3849 (N_3849,N_3716,N_3757);
nor U3850 (N_3850,N_3622,N_3793);
nor U3851 (N_3851,N_3719,N_3609);
and U3852 (N_3852,N_3783,N_3711);
nand U3853 (N_3853,N_3731,N_3734);
and U3854 (N_3854,N_3781,N_3633);
nand U3855 (N_3855,N_3758,N_3617);
nand U3856 (N_3856,N_3606,N_3671);
nand U3857 (N_3857,N_3674,N_3673);
or U3858 (N_3858,N_3723,N_3649);
nand U3859 (N_3859,N_3759,N_3745);
and U3860 (N_3860,N_3702,N_3641);
nor U3861 (N_3861,N_3707,N_3772);
nor U3862 (N_3862,N_3737,N_3721);
nand U3863 (N_3863,N_3669,N_3755);
or U3864 (N_3864,N_3703,N_3679);
and U3865 (N_3865,N_3651,N_3782);
and U3866 (N_3866,N_3628,N_3629);
nor U3867 (N_3867,N_3616,N_3644);
or U3868 (N_3868,N_3603,N_3767);
and U3869 (N_3869,N_3738,N_3784);
nor U3870 (N_3870,N_3684,N_3663);
nand U3871 (N_3871,N_3655,N_3627);
or U3872 (N_3872,N_3720,N_3744);
or U3873 (N_3873,N_3728,N_3677);
nor U3874 (N_3874,N_3657,N_3631);
nand U3875 (N_3875,N_3791,N_3787);
and U3876 (N_3876,N_3699,N_3799);
nor U3877 (N_3877,N_3654,N_3666);
nor U3878 (N_3878,N_3681,N_3786);
or U3879 (N_3879,N_3771,N_3770);
nor U3880 (N_3880,N_3625,N_3705);
and U3881 (N_3881,N_3640,N_3601);
and U3882 (N_3882,N_3682,N_3743);
nor U3883 (N_3883,N_3777,N_3722);
nor U3884 (N_3884,N_3607,N_3688);
or U3885 (N_3885,N_3618,N_3729);
nor U3886 (N_3886,N_3797,N_3764);
nand U3887 (N_3887,N_3659,N_3776);
nor U3888 (N_3888,N_3769,N_3730);
or U3889 (N_3889,N_3696,N_3732);
nor U3890 (N_3890,N_3747,N_3715);
or U3891 (N_3891,N_3695,N_3645);
and U3892 (N_3892,N_3683,N_3740);
and U3893 (N_3893,N_3785,N_3632);
or U3894 (N_3894,N_3661,N_3656);
and U3895 (N_3895,N_3798,N_3602);
nor U3896 (N_3896,N_3692,N_3725);
and U3897 (N_3897,N_3630,N_3700);
and U3898 (N_3898,N_3665,N_3685);
nand U3899 (N_3899,N_3653,N_3608);
nor U3900 (N_3900,N_3754,N_3698);
and U3901 (N_3901,N_3766,N_3644);
nand U3902 (N_3902,N_3792,N_3786);
or U3903 (N_3903,N_3776,N_3633);
or U3904 (N_3904,N_3719,N_3718);
or U3905 (N_3905,N_3722,N_3729);
and U3906 (N_3906,N_3656,N_3715);
nor U3907 (N_3907,N_3615,N_3675);
and U3908 (N_3908,N_3776,N_3781);
or U3909 (N_3909,N_3679,N_3687);
and U3910 (N_3910,N_3744,N_3670);
nor U3911 (N_3911,N_3701,N_3715);
nand U3912 (N_3912,N_3705,N_3743);
nor U3913 (N_3913,N_3739,N_3681);
nor U3914 (N_3914,N_3621,N_3614);
and U3915 (N_3915,N_3643,N_3687);
nand U3916 (N_3916,N_3775,N_3778);
nand U3917 (N_3917,N_3668,N_3601);
or U3918 (N_3918,N_3660,N_3611);
and U3919 (N_3919,N_3709,N_3638);
nand U3920 (N_3920,N_3755,N_3788);
xnor U3921 (N_3921,N_3710,N_3687);
nand U3922 (N_3922,N_3718,N_3798);
nor U3923 (N_3923,N_3777,N_3641);
nand U3924 (N_3924,N_3749,N_3693);
nand U3925 (N_3925,N_3716,N_3688);
or U3926 (N_3926,N_3660,N_3722);
or U3927 (N_3927,N_3749,N_3615);
nor U3928 (N_3928,N_3724,N_3734);
and U3929 (N_3929,N_3627,N_3668);
nand U3930 (N_3930,N_3632,N_3684);
nor U3931 (N_3931,N_3727,N_3684);
nor U3932 (N_3932,N_3621,N_3664);
or U3933 (N_3933,N_3730,N_3721);
xor U3934 (N_3934,N_3603,N_3694);
and U3935 (N_3935,N_3631,N_3632);
nand U3936 (N_3936,N_3764,N_3774);
nand U3937 (N_3937,N_3700,N_3603);
nand U3938 (N_3938,N_3746,N_3659);
nand U3939 (N_3939,N_3678,N_3611);
nor U3940 (N_3940,N_3711,N_3679);
and U3941 (N_3941,N_3736,N_3762);
and U3942 (N_3942,N_3735,N_3730);
nor U3943 (N_3943,N_3748,N_3657);
nor U3944 (N_3944,N_3629,N_3722);
or U3945 (N_3945,N_3725,N_3606);
nor U3946 (N_3946,N_3634,N_3633);
and U3947 (N_3947,N_3720,N_3742);
nand U3948 (N_3948,N_3757,N_3613);
and U3949 (N_3949,N_3693,N_3697);
and U3950 (N_3950,N_3634,N_3761);
and U3951 (N_3951,N_3775,N_3796);
nand U3952 (N_3952,N_3681,N_3776);
and U3953 (N_3953,N_3761,N_3605);
and U3954 (N_3954,N_3627,N_3730);
nor U3955 (N_3955,N_3698,N_3668);
and U3956 (N_3956,N_3684,N_3644);
and U3957 (N_3957,N_3620,N_3792);
nor U3958 (N_3958,N_3789,N_3738);
nor U3959 (N_3959,N_3667,N_3660);
nor U3960 (N_3960,N_3729,N_3602);
or U3961 (N_3961,N_3751,N_3613);
or U3962 (N_3962,N_3690,N_3723);
and U3963 (N_3963,N_3797,N_3701);
and U3964 (N_3964,N_3642,N_3791);
nor U3965 (N_3965,N_3615,N_3702);
or U3966 (N_3966,N_3693,N_3641);
or U3967 (N_3967,N_3794,N_3713);
or U3968 (N_3968,N_3686,N_3637);
and U3969 (N_3969,N_3610,N_3640);
and U3970 (N_3970,N_3788,N_3639);
nand U3971 (N_3971,N_3768,N_3743);
or U3972 (N_3972,N_3798,N_3758);
or U3973 (N_3973,N_3690,N_3671);
nand U3974 (N_3974,N_3644,N_3794);
nor U3975 (N_3975,N_3602,N_3683);
nand U3976 (N_3976,N_3775,N_3767);
and U3977 (N_3977,N_3650,N_3639);
or U3978 (N_3978,N_3679,N_3786);
nand U3979 (N_3979,N_3615,N_3677);
xor U3980 (N_3980,N_3790,N_3779);
nand U3981 (N_3981,N_3650,N_3749);
and U3982 (N_3982,N_3665,N_3700);
or U3983 (N_3983,N_3601,N_3713);
and U3984 (N_3984,N_3693,N_3681);
or U3985 (N_3985,N_3683,N_3796);
nor U3986 (N_3986,N_3748,N_3792);
or U3987 (N_3987,N_3741,N_3634);
or U3988 (N_3988,N_3656,N_3756);
or U3989 (N_3989,N_3641,N_3766);
nor U3990 (N_3990,N_3701,N_3770);
or U3991 (N_3991,N_3743,N_3621);
nor U3992 (N_3992,N_3791,N_3640);
nand U3993 (N_3993,N_3708,N_3684);
or U3994 (N_3994,N_3715,N_3621);
or U3995 (N_3995,N_3742,N_3688);
nor U3996 (N_3996,N_3622,N_3790);
or U3997 (N_3997,N_3767,N_3725);
nor U3998 (N_3998,N_3601,N_3704);
or U3999 (N_3999,N_3664,N_3647);
and U4000 (N_4000,N_3854,N_3846);
nand U4001 (N_4001,N_3801,N_3962);
nand U4002 (N_4002,N_3885,N_3910);
or U4003 (N_4003,N_3866,N_3900);
nor U4004 (N_4004,N_3805,N_3889);
or U4005 (N_4005,N_3983,N_3850);
and U4006 (N_4006,N_3862,N_3902);
nand U4007 (N_4007,N_3883,N_3894);
nor U4008 (N_4008,N_3965,N_3852);
or U4009 (N_4009,N_3917,N_3817);
nor U4010 (N_4010,N_3870,N_3928);
and U4011 (N_4011,N_3923,N_3864);
and U4012 (N_4012,N_3899,N_3958);
nor U4013 (N_4013,N_3897,N_3924);
nand U4014 (N_4014,N_3851,N_3814);
or U4015 (N_4015,N_3811,N_3944);
nor U4016 (N_4016,N_3874,N_3806);
nor U4017 (N_4017,N_3825,N_3886);
nand U4018 (N_4018,N_3990,N_3830);
and U4019 (N_4019,N_3999,N_3873);
nor U4020 (N_4020,N_3991,N_3833);
nor U4021 (N_4021,N_3935,N_3929);
nor U4022 (N_4022,N_3884,N_3842);
nor U4023 (N_4023,N_3980,N_3994);
and U4024 (N_4024,N_3967,N_3845);
and U4025 (N_4025,N_3841,N_3822);
or U4026 (N_4026,N_3998,N_3997);
and U4027 (N_4027,N_3986,N_3926);
nor U4028 (N_4028,N_3802,N_3875);
nor U4029 (N_4029,N_3911,N_3871);
and U4030 (N_4030,N_3966,N_3819);
or U4031 (N_4031,N_3843,N_3880);
nand U4032 (N_4032,N_3920,N_3823);
or U4033 (N_4033,N_3934,N_3878);
and U4034 (N_4034,N_3907,N_3933);
nor U4035 (N_4035,N_3867,N_3963);
nand U4036 (N_4036,N_3856,N_3804);
or U4037 (N_4037,N_3898,N_3930);
nor U4038 (N_4038,N_3912,N_3977);
nand U4039 (N_4039,N_3839,N_3987);
xor U4040 (N_4040,N_3890,N_3913);
nand U4041 (N_4041,N_3813,N_3946);
nand U4042 (N_4042,N_3887,N_3820);
and U4043 (N_4043,N_3893,N_3824);
nand U4044 (N_4044,N_3948,N_3868);
nand U4045 (N_4045,N_3859,N_3931);
nor U4046 (N_4046,N_3952,N_3838);
and U4047 (N_4047,N_3937,N_3895);
and U4048 (N_4048,N_3949,N_3849);
and U4049 (N_4049,N_3916,N_3959);
nor U4050 (N_4050,N_3972,N_3800);
nor U4051 (N_4051,N_3834,N_3985);
nand U4052 (N_4052,N_3975,N_3858);
nand U4053 (N_4053,N_3982,N_3844);
or U4054 (N_4054,N_3812,N_3888);
and U4055 (N_4055,N_3973,N_3943);
nand U4056 (N_4056,N_3938,N_3992);
nor U4057 (N_4057,N_3969,N_3974);
and U4058 (N_4058,N_3891,N_3970);
nand U4059 (N_4059,N_3951,N_3932);
or U4060 (N_4060,N_3837,N_3840);
or U4061 (N_4061,N_3908,N_3978);
and U4062 (N_4062,N_3818,N_3836);
or U4063 (N_4063,N_3989,N_3984);
and U4064 (N_4064,N_3879,N_3921);
and U4065 (N_4065,N_3956,N_3855);
nand U4066 (N_4066,N_3809,N_3955);
nor U4067 (N_4067,N_3872,N_3810);
nor U4068 (N_4068,N_3828,N_3922);
and U4069 (N_4069,N_3953,N_3863);
or U4070 (N_4070,N_3815,N_3803);
or U4071 (N_4071,N_3904,N_3925);
nand U4072 (N_4072,N_3941,N_3892);
nor U4073 (N_4073,N_3979,N_3865);
nand U4074 (N_4074,N_3832,N_3847);
or U4075 (N_4075,N_3876,N_3860);
nor U4076 (N_4076,N_3957,N_3816);
nor U4077 (N_4077,N_3993,N_3915);
or U4078 (N_4078,N_3882,N_3881);
nor U4079 (N_4079,N_3936,N_3954);
nand U4080 (N_4080,N_3961,N_3960);
nand U4081 (N_4081,N_3914,N_3848);
or U4082 (N_4082,N_3968,N_3976);
or U4083 (N_4083,N_3821,N_3861);
and U4084 (N_4084,N_3901,N_3877);
or U4085 (N_4085,N_3835,N_3853);
nand U4086 (N_4086,N_3831,N_3995);
nand U4087 (N_4087,N_3939,N_3950);
or U4088 (N_4088,N_3896,N_3827);
and U4089 (N_4089,N_3981,N_3808);
or U4090 (N_4090,N_3996,N_3906);
nor U4091 (N_4091,N_3829,N_3988);
nand U4092 (N_4092,N_3971,N_3857);
nor U4093 (N_4093,N_3940,N_3903);
and U4094 (N_4094,N_3919,N_3909);
nand U4095 (N_4095,N_3947,N_3905);
nor U4096 (N_4096,N_3826,N_3807);
nor U4097 (N_4097,N_3942,N_3918);
or U4098 (N_4098,N_3869,N_3945);
nor U4099 (N_4099,N_3964,N_3927);
and U4100 (N_4100,N_3867,N_3845);
nor U4101 (N_4101,N_3886,N_3987);
nand U4102 (N_4102,N_3946,N_3908);
nor U4103 (N_4103,N_3938,N_3804);
nor U4104 (N_4104,N_3901,N_3998);
and U4105 (N_4105,N_3982,N_3895);
and U4106 (N_4106,N_3932,N_3976);
and U4107 (N_4107,N_3998,N_3992);
or U4108 (N_4108,N_3924,N_3965);
and U4109 (N_4109,N_3958,N_3956);
and U4110 (N_4110,N_3854,N_3948);
and U4111 (N_4111,N_3963,N_3869);
and U4112 (N_4112,N_3958,N_3974);
nor U4113 (N_4113,N_3907,N_3871);
and U4114 (N_4114,N_3967,N_3828);
or U4115 (N_4115,N_3983,N_3806);
nand U4116 (N_4116,N_3882,N_3818);
and U4117 (N_4117,N_3958,N_3911);
and U4118 (N_4118,N_3830,N_3962);
and U4119 (N_4119,N_3875,N_3854);
nand U4120 (N_4120,N_3803,N_3836);
nand U4121 (N_4121,N_3881,N_3873);
nor U4122 (N_4122,N_3910,N_3831);
nand U4123 (N_4123,N_3986,N_3947);
nand U4124 (N_4124,N_3845,N_3907);
nor U4125 (N_4125,N_3857,N_3981);
and U4126 (N_4126,N_3950,N_3816);
or U4127 (N_4127,N_3869,N_3993);
and U4128 (N_4128,N_3867,N_3900);
and U4129 (N_4129,N_3896,N_3858);
and U4130 (N_4130,N_3824,N_3919);
or U4131 (N_4131,N_3940,N_3848);
nor U4132 (N_4132,N_3821,N_3974);
nor U4133 (N_4133,N_3922,N_3995);
and U4134 (N_4134,N_3803,N_3968);
nand U4135 (N_4135,N_3847,N_3828);
and U4136 (N_4136,N_3871,N_3921);
nand U4137 (N_4137,N_3912,N_3938);
and U4138 (N_4138,N_3887,N_3916);
or U4139 (N_4139,N_3930,N_3936);
nand U4140 (N_4140,N_3961,N_3872);
nor U4141 (N_4141,N_3918,N_3833);
nor U4142 (N_4142,N_3950,N_3858);
nor U4143 (N_4143,N_3974,N_3948);
nand U4144 (N_4144,N_3994,N_3919);
or U4145 (N_4145,N_3850,N_3838);
nor U4146 (N_4146,N_3916,N_3926);
nand U4147 (N_4147,N_3808,N_3826);
or U4148 (N_4148,N_3937,N_3964);
or U4149 (N_4149,N_3975,N_3980);
or U4150 (N_4150,N_3922,N_3893);
and U4151 (N_4151,N_3921,N_3873);
or U4152 (N_4152,N_3932,N_3831);
or U4153 (N_4153,N_3953,N_3855);
and U4154 (N_4154,N_3855,N_3827);
nand U4155 (N_4155,N_3999,N_3850);
nor U4156 (N_4156,N_3927,N_3828);
nor U4157 (N_4157,N_3942,N_3857);
or U4158 (N_4158,N_3940,N_3993);
nor U4159 (N_4159,N_3919,N_3803);
and U4160 (N_4160,N_3998,N_3965);
or U4161 (N_4161,N_3879,N_3969);
and U4162 (N_4162,N_3861,N_3964);
or U4163 (N_4163,N_3966,N_3910);
or U4164 (N_4164,N_3933,N_3878);
nand U4165 (N_4165,N_3988,N_3998);
xor U4166 (N_4166,N_3995,N_3814);
and U4167 (N_4167,N_3912,N_3871);
or U4168 (N_4168,N_3889,N_3935);
nor U4169 (N_4169,N_3999,N_3921);
or U4170 (N_4170,N_3922,N_3830);
nor U4171 (N_4171,N_3891,N_3928);
nand U4172 (N_4172,N_3893,N_3801);
and U4173 (N_4173,N_3894,N_3990);
or U4174 (N_4174,N_3990,N_3976);
and U4175 (N_4175,N_3909,N_3929);
nand U4176 (N_4176,N_3848,N_3971);
nand U4177 (N_4177,N_3977,N_3966);
nand U4178 (N_4178,N_3928,N_3994);
nor U4179 (N_4179,N_3824,N_3899);
nand U4180 (N_4180,N_3879,N_3839);
nor U4181 (N_4181,N_3998,N_3860);
and U4182 (N_4182,N_3826,N_3938);
or U4183 (N_4183,N_3950,N_3800);
nand U4184 (N_4184,N_3934,N_3868);
or U4185 (N_4185,N_3880,N_3983);
nor U4186 (N_4186,N_3840,N_3991);
nand U4187 (N_4187,N_3958,N_3811);
nand U4188 (N_4188,N_3991,N_3974);
or U4189 (N_4189,N_3875,N_3939);
nand U4190 (N_4190,N_3820,N_3976);
or U4191 (N_4191,N_3847,N_3845);
nor U4192 (N_4192,N_3889,N_3915);
and U4193 (N_4193,N_3858,N_3805);
and U4194 (N_4194,N_3817,N_3860);
nand U4195 (N_4195,N_3916,N_3832);
nor U4196 (N_4196,N_3946,N_3951);
nor U4197 (N_4197,N_3806,N_3880);
nor U4198 (N_4198,N_3982,N_3840);
nor U4199 (N_4199,N_3876,N_3980);
nor U4200 (N_4200,N_4017,N_4164);
nor U4201 (N_4201,N_4167,N_4171);
or U4202 (N_4202,N_4198,N_4073);
nor U4203 (N_4203,N_4033,N_4157);
or U4204 (N_4204,N_4173,N_4008);
nor U4205 (N_4205,N_4006,N_4098);
nor U4206 (N_4206,N_4087,N_4183);
and U4207 (N_4207,N_4194,N_4131);
nand U4208 (N_4208,N_4094,N_4185);
nand U4209 (N_4209,N_4177,N_4020);
nand U4210 (N_4210,N_4090,N_4019);
nor U4211 (N_4211,N_4065,N_4132);
nand U4212 (N_4212,N_4123,N_4011);
and U4213 (N_4213,N_4158,N_4076);
or U4214 (N_4214,N_4053,N_4142);
or U4215 (N_4215,N_4089,N_4088);
or U4216 (N_4216,N_4086,N_4047);
nor U4217 (N_4217,N_4037,N_4122);
nor U4218 (N_4218,N_4139,N_4030);
nor U4219 (N_4219,N_4068,N_4039);
or U4220 (N_4220,N_4197,N_4057);
or U4221 (N_4221,N_4191,N_4182);
nand U4222 (N_4222,N_4100,N_4025);
and U4223 (N_4223,N_4199,N_4118);
or U4224 (N_4224,N_4134,N_4113);
nand U4225 (N_4225,N_4045,N_4140);
or U4226 (N_4226,N_4052,N_4166);
nor U4227 (N_4227,N_4162,N_4061);
nand U4228 (N_4228,N_4168,N_4032);
or U4229 (N_4229,N_4069,N_4156);
nand U4230 (N_4230,N_4049,N_4135);
nor U4231 (N_4231,N_4026,N_4038);
nand U4232 (N_4232,N_4048,N_4040);
and U4233 (N_4233,N_4070,N_4195);
xor U4234 (N_4234,N_4097,N_4112);
or U4235 (N_4235,N_4064,N_4138);
nor U4236 (N_4236,N_4169,N_4159);
or U4237 (N_4237,N_4192,N_4063);
and U4238 (N_4238,N_4075,N_4143);
nor U4239 (N_4239,N_4092,N_4083);
or U4240 (N_4240,N_4161,N_4196);
or U4241 (N_4241,N_4145,N_4129);
or U4242 (N_4242,N_4104,N_4080);
and U4243 (N_4243,N_4108,N_4190);
or U4244 (N_4244,N_4015,N_4103);
and U4245 (N_4245,N_4029,N_4095);
nand U4246 (N_4246,N_4188,N_4114);
and U4247 (N_4247,N_4154,N_4148);
or U4248 (N_4248,N_4165,N_4137);
nand U4249 (N_4249,N_4124,N_4160);
nand U4250 (N_4250,N_4181,N_4189);
and U4251 (N_4251,N_4041,N_4078);
nand U4252 (N_4252,N_4013,N_4119);
nor U4253 (N_4253,N_4060,N_4042);
or U4254 (N_4254,N_4051,N_4043);
nand U4255 (N_4255,N_4133,N_4186);
or U4256 (N_4256,N_4116,N_4022);
nand U4257 (N_4257,N_4151,N_4121);
or U4258 (N_4258,N_4127,N_4102);
and U4259 (N_4259,N_4152,N_4021);
and U4260 (N_4260,N_4193,N_4144);
or U4261 (N_4261,N_4099,N_4105);
nor U4262 (N_4262,N_4009,N_4031);
nand U4263 (N_4263,N_4176,N_4110);
nand U4264 (N_4264,N_4172,N_4128);
nand U4265 (N_4265,N_4077,N_4179);
and U4266 (N_4266,N_4184,N_4111);
nand U4267 (N_4267,N_4027,N_4072);
nand U4268 (N_4268,N_4175,N_4056);
or U4269 (N_4269,N_4091,N_4126);
nand U4270 (N_4270,N_4012,N_4106);
and U4271 (N_4271,N_4004,N_4001);
and U4272 (N_4272,N_4000,N_4059);
and U4273 (N_4273,N_4034,N_4010);
nand U4274 (N_4274,N_4085,N_4005);
and U4275 (N_4275,N_4007,N_4180);
and U4276 (N_4276,N_4046,N_4093);
and U4277 (N_4277,N_4082,N_4035);
nor U4278 (N_4278,N_4147,N_4146);
nor U4279 (N_4279,N_4044,N_4081);
or U4280 (N_4280,N_4066,N_4117);
or U4281 (N_4281,N_4071,N_4141);
or U4282 (N_4282,N_4058,N_4187);
nor U4283 (N_4283,N_4120,N_4050);
nor U4284 (N_4284,N_4136,N_4014);
nand U4285 (N_4285,N_4036,N_4163);
nor U4286 (N_4286,N_4079,N_4024);
or U4287 (N_4287,N_4174,N_4074);
and U4288 (N_4288,N_4149,N_4018);
or U4289 (N_4289,N_4096,N_4130);
or U4290 (N_4290,N_4016,N_4101);
and U4291 (N_4291,N_4028,N_4054);
nand U4292 (N_4292,N_4003,N_4155);
or U4293 (N_4293,N_4084,N_4125);
nand U4294 (N_4294,N_4109,N_4002);
or U4295 (N_4295,N_4178,N_4055);
nor U4296 (N_4296,N_4170,N_4150);
nand U4297 (N_4297,N_4023,N_4062);
nand U4298 (N_4298,N_4115,N_4107);
and U4299 (N_4299,N_4067,N_4153);
nand U4300 (N_4300,N_4098,N_4080);
and U4301 (N_4301,N_4151,N_4149);
nand U4302 (N_4302,N_4196,N_4137);
and U4303 (N_4303,N_4106,N_4119);
or U4304 (N_4304,N_4127,N_4159);
nor U4305 (N_4305,N_4173,N_4097);
xor U4306 (N_4306,N_4120,N_4150);
and U4307 (N_4307,N_4022,N_4064);
or U4308 (N_4308,N_4074,N_4007);
and U4309 (N_4309,N_4123,N_4034);
and U4310 (N_4310,N_4102,N_4153);
or U4311 (N_4311,N_4089,N_4143);
nand U4312 (N_4312,N_4111,N_4006);
or U4313 (N_4313,N_4084,N_4102);
or U4314 (N_4314,N_4166,N_4016);
or U4315 (N_4315,N_4134,N_4111);
nor U4316 (N_4316,N_4092,N_4161);
and U4317 (N_4317,N_4179,N_4188);
nor U4318 (N_4318,N_4197,N_4145);
nor U4319 (N_4319,N_4062,N_4005);
nand U4320 (N_4320,N_4065,N_4182);
or U4321 (N_4321,N_4109,N_4003);
nand U4322 (N_4322,N_4078,N_4038);
or U4323 (N_4323,N_4009,N_4054);
nor U4324 (N_4324,N_4093,N_4174);
nor U4325 (N_4325,N_4107,N_4074);
nor U4326 (N_4326,N_4080,N_4181);
nand U4327 (N_4327,N_4170,N_4047);
nand U4328 (N_4328,N_4131,N_4120);
or U4329 (N_4329,N_4194,N_4048);
nor U4330 (N_4330,N_4071,N_4188);
and U4331 (N_4331,N_4121,N_4075);
nor U4332 (N_4332,N_4159,N_4186);
or U4333 (N_4333,N_4131,N_4153);
and U4334 (N_4334,N_4195,N_4083);
and U4335 (N_4335,N_4023,N_4065);
and U4336 (N_4336,N_4102,N_4037);
and U4337 (N_4337,N_4157,N_4190);
or U4338 (N_4338,N_4092,N_4097);
nor U4339 (N_4339,N_4103,N_4192);
or U4340 (N_4340,N_4099,N_4193);
nor U4341 (N_4341,N_4070,N_4026);
nand U4342 (N_4342,N_4033,N_4083);
nand U4343 (N_4343,N_4030,N_4007);
and U4344 (N_4344,N_4152,N_4167);
or U4345 (N_4345,N_4077,N_4008);
or U4346 (N_4346,N_4086,N_4041);
or U4347 (N_4347,N_4190,N_4166);
and U4348 (N_4348,N_4090,N_4023);
or U4349 (N_4349,N_4162,N_4129);
nor U4350 (N_4350,N_4132,N_4069);
nand U4351 (N_4351,N_4069,N_4065);
or U4352 (N_4352,N_4110,N_4162);
nand U4353 (N_4353,N_4108,N_4126);
and U4354 (N_4354,N_4077,N_4146);
and U4355 (N_4355,N_4135,N_4154);
and U4356 (N_4356,N_4141,N_4105);
and U4357 (N_4357,N_4010,N_4163);
nor U4358 (N_4358,N_4109,N_4013);
nor U4359 (N_4359,N_4120,N_4065);
nand U4360 (N_4360,N_4199,N_4053);
nand U4361 (N_4361,N_4160,N_4151);
nor U4362 (N_4362,N_4021,N_4167);
or U4363 (N_4363,N_4109,N_4153);
and U4364 (N_4364,N_4016,N_4065);
nor U4365 (N_4365,N_4106,N_4073);
or U4366 (N_4366,N_4057,N_4098);
nand U4367 (N_4367,N_4044,N_4059);
nor U4368 (N_4368,N_4082,N_4160);
or U4369 (N_4369,N_4000,N_4061);
nand U4370 (N_4370,N_4137,N_4162);
and U4371 (N_4371,N_4119,N_4132);
nor U4372 (N_4372,N_4181,N_4100);
or U4373 (N_4373,N_4172,N_4025);
nor U4374 (N_4374,N_4057,N_4158);
nor U4375 (N_4375,N_4143,N_4156);
and U4376 (N_4376,N_4064,N_4184);
or U4377 (N_4377,N_4138,N_4028);
nor U4378 (N_4378,N_4103,N_4180);
and U4379 (N_4379,N_4140,N_4028);
nor U4380 (N_4380,N_4024,N_4096);
nor U4381 (N_4381,N_4000,N_4154);
nor U4382 (N_4382,N_4140,N_4004);
nor U4383 (N_4383,N_4091,N_4160);
nor U4384 (N_4384,N_4103,N_4061);
or U4385 (N_4385,N_4048,N_4028);
nand U4386 (N_4386,N_4082,N_4104);
nor U4387 (N_4387,N_4132,N_4177);
nor U4388 (N_4388,N_4162,N_4034);
or U4389 (N_4389,N_4198,N_4172);
or U4390 (N_4390,N_4053,N_4123);
nor U4391 (N_4391,N_4112,N_4137);
and U4392 (N_4392,N_4193,N_4102);
or U4393 (N_4393,N_4096,N_4103);
and U4394 (N_4394,N_4116,N_4189);
and U4395 (N_4395,N_4155,N_4074);
nor U4396 (N_4396,N_4108,N_4196);
nand U4397 (N_4397,N_4143,N_4000);
nor U4398 (N_4398,N_4105,N_4001);
nor U4399 (N_4399,N_4166,N_4098);
and U4400 (N_4400,N_4289,N_4386);
nand U4401 (N_4401,N_4215,N_4260);
nand U4402 (N_4402,N_4268,N_4334);
nor U4403 (N_4403,N_4281,N_4351);
or U4404 (N_4404,N_4229,N_4329);
and U4405 (N_4405,N_4220,N_4364);
nor U4406 (N_4406,N_4237,N_4291);
nor U4407 (N_4407,N_4280,N_4217);
nand U4408 (N_4408,N_4342,N_4208);
and U4409 (N_4409,N_4224,N_4321);
or U4410 (N_4410,N_4396,N_4264);
or U4411 (N_4411,N_4286,N_4212);
or U4412 (N_4412,N_4344,N_4262);
and U4413 (N_4413,N_4335,N_4257);
or U4414 (N_4414,N_4241,N_4200);
and U4415 (N_4415,N_4216,N_4387);
and U4416 (N_4416,N_4375,N_4211);
and U4417 (N_4417,N_4361,N_4383);
nand U4418 (N_4418,N_4398,N_4290);
and U4419 (N_4419,N_4206,N_4274);
and U4420 (N_4420,N_4338,N_4205);
and U4421 (N_4421,N_4303,N_4359);
nor U4422 (N_4422,N_4341,N_4323);
or U4423 (N_4423,N_4372,N_4324);
or U4424 (N_4424,N_4249,N_4306);
nand U4425 (N_4425,N_4201,N_4267);
or U4426 (N_4426,N_4265,N_4242);
nor U4427 (N_4427,N_4231,N_4270);
nor U4428 (N_4428,N_4238,N_4261);
xor U4429 (N_4429,N_4331,N_4311);
nor U4430 (N_4430,N_4292,N_4307);
and U4431 (N_4431,N_4388,N_4239);
nand U4432 (N_4432,N_4340,N_4374);
nor U4433 (N_4433,N_4373,N_4279);
nor U4434 (N_4434,N_4310,N_4380);
or U4435 (N_4435,N_4272,N_4235);
nor U4436 (N_4436,N_4254,N_4395);
nor U4437 (N_4437,N_4252,N_4271);
or U4438 (N_4438,N_4213,N_4382);
and U4439 (N_4439,N_4230,N_4283);
or U4440 (N_4440,N_4243,N_4333);
nand U4441 (N_4441,N_4357,N_4317);
nor U4442 (N_4442,N_4297,N_4332);
or U4443 (N_4443,N_4240,N_4360);
and U4444 (N_4444,N_4245,N_4392);
nand U4445 (N_4445,N_4207,N_4325);
nor U4446 (N_4446,N_4393,N_4326);
nor U4447 (N_4447,N_4223,N_4219);
xor U4448 (N_4448,N_4348,N_4247);
xor U4449 (N_4449,N_4222,N_4336);
and U4450 (N_4450,N_4355,N_4378);
nand U4451 (N_4451,N_4248,N_4371);
nand U4452 (N_4452,N_4285,N_4236);
nand U4453 (N_4453,N_4397,N_4308);
nand U4454 (N_4454,N_4256,N_4246);
nand U4455 (N_4455,N_4379,N_4314);
nor U4456 (N_4456,N_4255,N_4287);
nor U4457 (N_4457,N_4391,N_4278);
and U4458 (N_4458,N_4253,N_4221);
nand U4459 (N_4459,N_4273,N_4366);
and U4460 (N_4460,N_4353,N_4367);
or U4461 (N_4461,N_4202,N_4269);
or U4462 (N_4462,N_4210,N_4302);
and U4463 (N_4463,N_4365,N_4250);
nand U4464 (N_4464,N_4381,N_4214);
nand U4465 (N_4465,N_4244,N_4316);
nor U4466 (N_4466,N_4251,N_4209);
or U4467 (N_4467,N_4259,N_4218);
nor U4468 (N_4468,N_4295,N_4370);
and U4469 (N_4469,N_4343,N_4347);
or U4470 (N_4470,N_4377,N_4376);
nand U4471 (N_4471,N_4266,N_4389);
nand U4472 (N_4472,N_4305,N_4309);
nand U4473 (N_4473,N_4349,N_4350);
nor U4474 (N_4474,N_4358,N_4282);
or U4475 (N_4475,N_4363,N_4277);
nor U4476 (N_4476,N_4339,N_4368);
or U4477 (N_4477,N_4327,N_4293);
nand U4478 (N_4478,N_4225,N_4232);
nand U4479 (N_4479,N_4330,N_4233);
or U4480 (N_4480,N_4258,N_4318);
and U4481 (N_4481,N_4313,N_4298);
and U4482 (N_4482,N_4346,N_4362);
nand U4483 (N_4483,N_4328,N_4284);
nand U4484 (N_4484,N_4322,N_4354);
or U4485 (N_4485,N_4204,N_4369);
nor U4486 (N_4486,N_4228,N_4263);
nor U4487 (N_4487,N_4352,N_4394);
nand U4488 (N_4488,N_4399,N_4304);
and U4489 (N_4489,N_4315,N_4319);
nand U4490 (N_4490,N_4345,N_4390);
nand U4491 (N_4491,N_4356,N_4234);
or U4492 (N_4492,N_4275,N_4312);
nand U4493 (N_4493,N_4203,N_4300);
and U4494 (N_4494,N_4384,N_4301);
nand U4495 (N_4495,N_4296,N_4288);
or U4496 (N_4496,N_4337,N_4227);
or U4497 (N_4497,N_4320,N_4299);
nand U4498 (N_4498,N_4276,N_4226);
nor U4499 (N_4499,N_4385,N_4294);
nor U4500 (N_4500,N_4357,N_4364);
and U4501 (N_4501,N_4399,N_4312);
or U4502 (N_4502,N_4336,N_4259);
and U4503 (N_4503,N_4388,N_4363);
or U4504 (N_4504,N_4306,N_4315);
or U4505 (N_4505,N_4343,N_4270);
nor U4506 (N_4506,N_4374,N_4380);
nor U4507 (N_4507,N_4311,N_4324);
and U4508 (N_4508,N_4325,N_4393);
or U4509 (N_4509,N_4258,N_4319);
nand U4510 (N_4510,N_4236,N_4229);
nor U4511 (N_4511,N_4360,N_4210);
nor U4512 (N_4512,N_4319,N_4366);
or U4513 (N_4513,N_4368,N_4323);
and U4514 (N_4514,N_4284,N_4268);
nor U4515 (N_4515,N_4284,N_4226);
and U4516 (N_4516,N_4376,N_4266);
nand U4517 (N_4517,N_4381,N_4331);
nor U4518 (N_4518,N_4397,N_4260);
and U4519 (N_4519,N_4319,N_4317);
nor U4520 (N_4520,N_4306,N_4345);
nor U4521 (N_4521,N_4293,N_4390);
or U4522 (N_4522,N_4311,N_4262);
nand U4523 (N_4523,N_4383,N_4381);
and U4524 (N_4524,N_4278,N_4367);
nand U4525 (N_4525,N_4339,N_4221);
nor U4526 (N_4526,N_4389,N_4221);
nor U4527 (N_4527,N_4370,N_4214);
nand U4528 (N_4528,N_4327,N_4307);
nand U4529 (N_4529,N_4372,N_4291);
or U4530 (N_4530,N_4323,N_4284);
nand U4531 (N_4531,N_4329,N_4293);
nor U4532 (N_4532,N_4382,N_4348);
nor U4533 (N_4533,N_4339,N_4216);
and U4534 (N_4534,N_4226,N_4343);
nor U4535 (N_4535,N_4243,N_4242);
or U4536 (N_4536,N_4231,N_4336);
nand U4537 (N_4537,N_4292,N_4323);
and U4538 (N_4538,N_4220,N_4361);
or U4539 (N_4539,N_4208,N_4266);
nor U4540 (N_4540,N_4359,N_4353);
or U4541 (N_4541,N_4310,N_4211);
nand U4542 (N_4542,N_4324,N_4338);
nor U4543 (N_4543,N_4271,N_4285);
nand U4544 (N_4544,N_4299,N_4201);
nor U4545 (N_4545,N_4299,N_4333);
and U4546 (N_4546,N_4296,N_4395);
nand U4547 (N_4547,N_4204,N_4292);
and U4548 (N_4548,N_4384,N_4228);
nand U4549 (N_4549,N_4294,N_4341);
or U4550 (N_4550,N_4335,N_4212);
nand U4551 (N_4551,N_4318,N_4279);
and U4552 (N_4552,N_4260,N_4333);
and U4553 (N_4553,N_4297,N_4356);
nor U4554 (N_4554,N_4225,N_4218);
nand U4555 (N_4555,N_4326,N_4292);
nand U4556 (N_4556,N_4337,N_4282);
and U4557 (N_4557,N_4291,N_4355);
nand U4558 (N_4558,N_4235,N_4302);
nor U4559 (N_4559,N_4231,N_4221);
and U4560 (N_4560,N_4249,N_4346);
and U4561 (N_4561,N_4226,N_4330);
or U4562 (N_4562,N_4250,N_4313);
nand U4563 (N_4563,N_4351,N_4231);
nor U4564 (N_4564,N_4312,N_4331);
nor U4565 (N_4565,N_4346,N_4268);
and U4566 (N_4566,N_4328,N_4341);
nand U4567 (N_4567,N_4298,N_4297);
nor U4568 (N_4568,N_4354,N_4215);
nor U4569 (N_4569,N_4229,N_4247);
or U4570 (N_4570,N_4287,N_4371);
and U4571 (N_4571,N_4362,N_4224);
and U4572 (N_4572,N_4268,N_4376);
and U4573 (N_4573,N_4336,N_4212);
nor U4574 (N_4574,N_4394,N_4368);
or U4575 (N_4575,N_4370,N_4280);
nand U4576 (N_4576,N_4274,N_4229);
nor U4577 (N_4577,N_4385,N_4368);
nand U4578 (N_4578,N_4203,N_4275);
or U4579 (N_4579,N_4302,N_4321);
or U4580 (N_4580,N_4397,N_4384);
or U4581 (N_4581,N_4254,N_4219);
or U4582 (N_4582,N_4396,N_4303);
nand U4583 (N_4583,N_4258,N_4300);
nand U4584 (N_4584,N_4234,N_4240);
nor U4585 (N_4585,N_4320,N_4342);
nor U4586 (N_4586,N_4257,N_4253);
nor U4587 (N_4587,N_4349,N_4315);
or U4588 (N_4588,N_4269,N_4388);
or U4589 (N_4589,N_4377,N_4373);
nor U4590 (N_4590,N_4381,N_4291);
and U4591 (N_4591,N_4285,N_4245);
or U4592 (N_4592,N_4305,N_4370);
nand U4593 (N_4593,N_4347,N_4207);
and U4594 (N_4594,N_4253,N_4220);
nor U4595 (N_4595,N_4264,N_4257);
nor U4596 (N_4596,N_4321,N_4367);
and U4597 (N_4597,N_4358,N_4308);
nand U4598 (N_4598,N_4310,N_4364);
nor U4599 (N_4599,N_4246,N_4343);
nor U4600 (N_4600,N_4486,N_4493);
or U4601 (N_4601,N_4533,N_4444);
nand U4602 (N_4602,N_4580,N_4404);
nand U4603 (N_4603,N_4438,N_4521);
or U4604 (N_4604,N_4453,N_4432);
and U4605 (N_4605,N_4416,N_4531);
or U4606 (N_4606,N_4482,N_4490);
and U4607 (N_4607,N_4562,N_4400);
nand U4608 (N_4608,N_4410,N_4544);
nand U4609 (N_4609,N_4460,N_4512);
nand U4610 (N_4610,N_4534,N_4450);
and U4611 (N_4611,N_4518,N_4478);
nor U4612 (N_4612,N_4553,N_4592);
nor U4613 (N_4613,N_4506,N_4436);
nor U4614 (N_4614,N_4520,N_4441);
nand U4615 (N_4615,N_4408,N_4567);
or U4616 (N_4616,N_4437,N_4421);
or U4617 (N_4617,N_4401,N_4536);
and U4618 (N_4618,N_4523,N_4557);
and U4619 (N_4619,N_4476,N_4428);
nand U4620 (N_4620,N_4508,N_4491);
nand U4621 (N_4621,N_4528,N_4429);
nand U4622 (N_4622,N_4412,N_4530);
and U4623 (N_4623,N_4470,N_4403);
nand U4624 (N_4624,N_4517,N_4575);
nand U4625 (N_4625,N_4524,N_4417);
or U4626 (N_4626,N_4415,N_4431);
nand U4627 (N_4627,N_4496,N_4465);
and U4628 (N_4628,N_4402,N_4502);
or U4629 (N_4629,N_4595,N_4519);
xor U4630 (N_4630,N_4591,N_4419);
or U4631 (N_4631,N_4598,N_4448);
nand U4632 (N_4632,N_4549,N_4462);
nand U4633 (N_4633,N_4498,N_4464);
nor U4634 (N_4634,N_4452,N_4563);
nor U4635 (N_4635,N_4568,N_4426);
nor U4636 (N_4636,N_4588,N_4573);
and U4637 (N_4637,N_4546,N_4541);
nor U4638 (N_4638,N_4420,N_4487);
or U4639 (N_4639,N_4561,N_4550);
nand U4640 (N_4640,N_4593,N_4494);
nor U4641 (N_4641,N_4527,N_4529);
nand U4642 (N_4642,N_4499,N_4578);
nand U4643 (N_4643,N_4433,N_4525);
nand U4644 (N_4644,N_4405,N_4547);
nand U4645 (N_4645,N_4511,N_4583);
and U4646 (N_4646,N_4514,N_4463);
and U4647 (N_4647,N_4477,N_4467);
and U4648 (N_4648,N_4451,N_4579);
and U4649 (N_4649,N_4570,N_4459);
xor U4650 (N_4650,N_4474,N_4440);
and U4651 (N_4651,N_4468,N_4409);
nand U4652 (N_4652,N_4425,N_4590);
nand U4653 (N_4653,N_4475,N_4449);
and U4654 (N_4654,N_4522,N_4571);
or U4655 (N_4655,N_4473,N_4542);
nor U4656 (N_4656,N_4548,N_4430);
nor U4657 (N_4657,N_4551,N_4565);
nor U4658 (N_4658,N_4545,N_4532);
or U4659 (N_4659,N_4479,N_4501);
nand U4660 (N_4660,N_4585,N_4576);
or U4661 (N_4661,N_4543,N_4407);
or U4662 (N_4662,N_4504,N_4439);
or U4663 (N_4663,N_4503,N_4446);
nand U4664 (N_4664,N_4596,N_4454);
or U4665 (N_4665,N_4569,N_4558);
nor U4666 (N_4666,N_4427,N_4485);
nor U4667 (N_4667,N_4555,N_4535);
nand U4668 (N_4668,N_4566,N_4552);
nand U4669 (N_4669,N_4577,N_4564);
nor U4670 (N_4670,N_4472,N_4414);
and U4671 (N_4671,N_4586,N_4418);
and U4672 (N_4672,N_4554,N_4599);
nand U4673 (N_4673,N_4574,N_4471);
or U4674 (N_4674,N_4589,N_4516);
nor U4675 (N_4675,N_4484,N_4424);
nand U4676 (N_4676,N_4456,N_4495);
and U4677 (N_4677,N_4513,N_4556);
and U4678 (N_4678,N_4537,N_4507);
and U4679 (N_4679,N_4455,N_4413);
nor U4680 (N_4680,N_4435,N_4434);
or U4681 (N_4681,N_4560,N_4510);
nand U4682 (N_4682,N_4497,N_4466);
nor U4683 (N_4683,N_4481,N_4445);
nand U4684 (N_4684,N_4480,N_4488);
or U4685 (N_4685,N_4447,N_4442);
nand U4686 (N_4686,N_4587,N_4500);
and U4687 (N_4687,N_4594,N_4509);
and U4688 (N_4688,N_4411,N_4443);
or U4689 (N_4689,N_4539,N_4559);
nand U4690 (N_4690,N_4461,N_4458);
nand U4691 (N_4691,N_4526,N_4406);
or U4692 (N_4692,N_4483,N_4597);
nand U4693 (N_4693,N_4572,N_4540);
nor U4694 (N_4694,N_4422,N_4469);
or U4695 (N_4695,N_4581,N_4538);
and U4696 (N_4696,N_4423,N_4582);
nor U4697 (N_4697,N_4584,N_4489);
nor U4698 (N_4698,N_4505,N_4515);
nand U4699 (N_4699,N_4457,N_4492);
or U4700 (N_4700,N_4578,N_4441);
nand U4701 (N_4701,N_4549,N_4465);
and U4702 (N_4702,N_4533,N_4475);
and U4703 (N_4703,N_4531,N_4458);
or U4704 (N_4704,N_4502,N_4546);
and U4705 (N_4705,N_4462,N_4519);
and U4706 (N_4706,N_4597,N_4548);
nand U4707 (N_4707,N_4524,N_4452);
nand U4708 (N_4708,N_4542,N_4567);
or U4709 (N_4709,N_4592,N_4561);
nand U4710 (N_4710,N_4548,N_4552);
nor U4711 (N_4711,N_4468,N_4426);
nor U4712 (N_4712,N_4499,N_4576);
and U4713 (N_4713,N_4506,N_4437);
nand U4714 (N_4714,N_4542,N_4479);
nor U4715 (N_4715,N_4597,N_4547);
and U4716 (N_4716,N_4459,N_4515);
nor U4717 (N_4717,N_4537,N_4453);
nor U4718 (N_4718,N_4492,N_4516);
nor U4719 (N_4719,N_4481,N_4448);
nor U4720 (N_4720,N_4538,N_4474);
nor U4721 (N_4721,N_4415,N_4411);
nor U4722 (N_4722,N_4587,N_4432);
nand U4723 (N_4723,N_4572,N_4583);
nor U4724 (N_4724,N_4553,N_4460);
nand U4725 (N_4725,N_4523,N_4479);
and U4726 (N_4726,N_4444,N_4432);
nor U4727 (N_4727,N_4593,N_4419);
and U4728 (N_4728,N_4596,N_4552);
or U4729 (N_4729,N_4435,N_4588);
or U4730 (N_4730,N_4591,N_4501);
or U4731 (N_4731,N_4458,N_4444);
and U4732 (N_4732,N_4595,N_4547);
or U4733 (N_4733,N_4570,N_4517);
or U4734 (N_4734,N_4467,N_4491);
and U4735 (N_4735,N_4526,N_4401);
nor U4736 (N_4736,N_4405,N_4535);
and U4737 (N_4737,N_4425,N_4447);
nor U4738 (N_4738,N_4410,N_4515);
nor U4739 (N_4739,N_4499,N_4460);
nand U4740 (N_4740,N_4587,N_4446);
and U4741 (N_4741,N_4513,N_4481);
nor U4742 (N_4742,N_4540,N_4476);
nand U4743 (N_4743,N_4585,N_4566);
or U4744 (N_4744,N_4473,N_4444);
xnor U4745 (N_4745,N_4412,N_4507);
and U4746 (N_4746,N_4450,N_4413);
nor U4747 (N_4747,N_4404,N_4540);
and U4748 (N_4748,N_4499,N_4583);
or U4749 (N_4749,N_4514,N_4418);
nand U4750 (N_4750,N_4483,N_4547);
nor U4751 (N_4751,N_4455,N_4564);
nor U4752 (N_4752,N_4564,N_4426);
nor U4753 (N_4753,N_4586,N_4508);
or U4754 (N_4754,N_4489,N_4537);
nor U4755 (N_4755,N_4421,N_4493);
xor U4756 (N_4756,N_4524,N_4517);
and U4757 (N_4757,N_4465,N_4595);
nor U4758 (N_4758,N_4577,N_4582);
nand U4759 (N_4759,N_4554,N_4589);
or U4760 (N_4760,N_4497,N_4403);
and U4761 (N_4761,N_4468,N_4517);
nor U4762 (N_4762,N_4544,N_4461);
nand U4763 (N_4763,N_4550,N_4548);
nand U4764 (N_4764,N_4575,N_4500);
nand U4765 (N_4765,N_4520,N_4462);
nor U4766 (N_4766,N_4551,N_4406);
or U4767 (N_4767,N_4533,N_4405);
or U4768 (N_4768,N_4467,N_4432);
and U4769 (N_4769,N_4412,N_4521);
nor U4770 (N_4770,N_4599,N_4543);
and U4771 (N_4771,N_4493,N_4418);
nor U4772 (N_4772,N_4553,N_4501);
nand U4773 (N_4773,N_4571,N_4583);
nand U4774 (N_4774,N_4474,N_4401);
or U4775 (N_4775,N_4417,N_4440);
and U4776 (N_4776,N_4519,N_4439);
xor U4777 (N_4777,N_4426,N_4549);
and U4778 (N_4778,N_4539,N_4497);
xnor U4779 (N_4779,N_4559,N_4424);
or U4780 (N_4780,N_4540,N_4430);
and U4781 (N_4781,N_4478,N_4483);
nand U4782 (N_4782,N_4427,N_4489);
or U4783 (N_4783,N_4403,N_4445);
and U4784 (N_4784,N_4444,N_4423);
xor U4785 (N_4785,N_4510,N_4541);
nor U4786 (N_4786,N_4433,N_4405);
nor U4787 (N_4787,N_4431,N_4435);
and U4788 (N_4788,N_4500,N_4407);
or U4789 (N_4789,N_4431,N_4595);
and U4790 (N_4790,N_4533,N_4563);
or U4791 (N_4791,N_4563,N_4592);
nand U4792 (N_4792,N_4432,N_4456);
or U4793 (N_4793,N_4528,N_4586);
nor U4794 (N_4794,N_4542,N_4482);
nor U4795 (N_4795,N_4497,N_4577);
nor U4796 (N_4796,N_4568,N_4550);
nand U4797 (N_4797,N_4588,N_4567);
and U4798 (N_4798,N_4585,N_4598);
nand U4799 (N_4799,N_4460,N_4426);
nand U4800 (N_4800,N_4773,N_4711);
and U4801 (N_4801,N_4732,N_4605);
nor U4802 (N_4802,N_4672,N_4717);
or U4803 (N_4803,N_4639,N_4739);
and U4804 (N_4804,N_4626,N_4693);
nand U4805 (N_4805,N_4680,N_4759);
or U4806 (N_4806,N_4785,N_4766);
or U4807 (N_4807,N_4757,N_4608);
or U4808 (N_4808,N_4613,N_4687);
nand U4809 (N_4809,N_4784,N_4606);
or U4810 (N_4810,N_4673,N_4601);
nand U4811 (N_4811,N_4659,N_4665);
nor U4812 (N_4812,N_4628,N_4780);
or U4813 (N_4813,N_4789,N_4707);
or U4814 (N_4814,N_4640,N_4612);
nor U4815 (N_4815,N_4741,N_4703);
nand U4816 (N_4816,N_4768,N_4798);
or U4817 (N_4817,N_4704,N_4735);
nor U4818 (N_4818,N_4736,N_4682);
nor U4819 (N_4819,N_4622,N_4633);
nor U4820 (N_4820,N_4635,N_4714);
nor U4821 (N_4821,N_4775,N_4660);
and U4822 (N_4822,N_4716,N_4718);
or U4823 (N_4823,N_4638,N_4676);
nor U4824 (N_4824,N_4730,N_4697);
nor U4825 (N_4825,N_4740,N_4647);
nor U4826 (N_4826,N_4708,N_4683);
nor U4827 (N_4827,N_4685,N_4765);
and U4828 (N_4828,N_4669,N_4778);
and U4829 (N_4829,N_4652,N_4603);
or U4830 (N_4830,N_4701,N_4787);
and U4831 (N_4831,N_4607,N_4793);
or U4832 (N_4832,N_4706,N_4772);
nand U4833 (N_4833,N_4667,N_4634);
and U4834 (N_4834,N_4769,N_4637);
and U4835 (N_4835,N_4630,N_4783);
and U4836 (N_4836,N_4642,N_4770);
and U4837 (N_4837,N_4602,N_4752);
or U4838 (N_4838,N_4729,N_4650);
nor U4839 (N_4839,N_4699,N_4748);
nor U4840 (N_4840,N_4725,N_4636);
nor U4841 (N_4841,N_4745,N_4742);
xnor U4842 (N_4842,N_4782,N_4743);
nor U4843 (N_4843,N_4781,N_4698);
or U4844 (N_4844,N_4670,N_4727);
nand U4845 (N_4845,N_4734,N_4648);
nand U4846 (N_4846,N_4651,N_4666);
nand U4847 (N_4847,N_4604,N_4649);
nand U4848 (N_4848,N_4689,N_4653);
and U4849 (N_4849,N_4702,N_4654);
or U4850 (N_4850,N_4746,N_4617);
and U4851 (N_4851,N_4720,N_4762);
and U4852 (N_4852,N_4629,N_4758);
and U4853 (N_4853,N_4696,N_4795);
or U4854 (N_4854,N_4750,N_4709);
and U4855 (N_4855,N_4763,N_4663);
nor U4856 (N_4856,N_4712,N_4799);
or U4857 (N_4857,N_4662,N_4722);
nand U4858 (N_4858,N_4645,N_4779);
nand U4859 (N_4859,N_4747,N_4731);
and U4860 (N_4860,N_4668,N_4797);
nor U4861 (N_4861,N_4688,N_4710);
nand U4862 (N_4862,N_4794,N_4691);
nor U4863 (N_4863,N_4726,N_4627);
and U4864 (N_4864,N_4611,N_4671);
nand U4865 (N_4865,N_4675,N_4756);
and U4866 (N_4866,N_4771,N_4681);
and U4867 (N_4867,N_4641,N_4791);
or U4868 (N_4868,N_4620,N_4615);
and U4869 (N_4869,N_4621,N_4624);
nor U4870 (N_4870,N_4788,N_4658);
nand U4871 (N_4871,N_4677,N_4690);
nand U4872 (N_4872,N_4796,N_4625);
and U4873 (N_4873,N_4655,N_4656);
or U4874 (N_4874,N_4737,N_4723);
and U4875 (N_4875,N_4679,N_4644);
nand U4876 (N_4876,N_4761,N_4616);
nand U4877 (N_4877,N_4774,N_4678);
and U4878 (N_4878,N_4610,N_4755);
or U4879 (N_4879,N_4753,N_4764);
or U4880 (N_4880,N_4674,N_4600);
and U4881 (N_4881,N_4684,N_4694);
and U4882 (N_4882,N_4754,N_4749);
and U4883 (N_4883,N_4614,N_4777);
or U4884 (N_4884,N_4724,N_4618);
or U4885 (N_4885,N_4776,N_4713);
or U4886 (N_4886,N_4631,N_4751);
and U4887 (N_4887,N_4661,N_4705);
nand U4888 (N_4888,N_4632,N_4664);
or U4889 (N_4889,N_4646,N_4686);
nand U4890 (N_4890,N_4767,N_4792);
nor U4891 (N_4891,N_4619,N_4643);
and U4892 (N_4892,N_4715,N_4738);
nor U4893 (N_4893,N_4609,N_4695);
nand U4894 (N_4894,N_4790,N_4760);
nand U4895 (N_4895,N_4692,N_4721);
nand U4896 (N_4896,N_4623,N_4728);
nor U4897 (N_4897,N_4657,N_4744);
or U4898 (N_4898,N_4786,N_4700);
nor U4899 (N_4899,N_4719,N_4733);
nand U4900 (N_4900,N_4745,N_4764);
nor U4901 (N_4901,N_4721,N_4618);
or U4902 (N_4902,N_4685,N_4748);
xnor U4903 (N_4903,N_4755,N_4781);
or U4904 (N_4904,N_4610,N_4684);
or U4905 (N_4905,N_4711,N_4694);
nor U4906 (N_4906,N_4755,N_4680);
or U4907 (N_4907,N_4773,N_4744);
nand U4908 (N_4908,N_4741,N_4723);
nand U4909 (N_4909,N_4655,N_4734);
nor U4910 (N_4910,N_4745,N_4600);
or U4911 (N_4911,N_4693,N_4718);
nand U4912 (N_4912,N_4799,N_4766);
or U4913 (N_4913,N_4657,N_4772);
or U4914 (N_4914,N_4794,N_4638);
nor U4915 (N_4915,N_4673,N_4667);
nor U4916 (N_4916,N_4665,N_4728);
nand U4917 (N_4917,N_4742,N_4719);
nor U4918 (N_4918,N_4626,N_4765);
or U4919 (N_4919,N_4709,N_4767);
nand U4920 (N_4920,N_4750,N_4650);
nand U4921 (N_4921,N_4792,N_4714);
and U4922 (N_4922,N_4672,N_4707);
nand U4923 (N_4923,N_4777,N_4700);
and U4924 (N_4924,N_4753,N_4681);
nand U4925 (N_4925,N_4798,N_4653);
nor U4926 (N_4926,N_4759,N_4631);
and U4927 (N_4927,N_4745,N_4618);
and U4928 (N_4928,N_4780,N_4686);
or U4929 (N_4929,N_4650,N_4620);
or U4930 (N_4930,N_4602,N_4616);
and U4931 (N_4931,N_4699,N_4743);
or U4932 (N_4932,N_4738,N_4739);
nand U4933 (N_4933,N_4648,N_4612);
or U4934 (N_4934,N_4619,N_4725);
nand U4935 (N_4935,N_4629,N_4717);
nand U4936 (N_4936,N_4634,N_4616);
or U4937 (N_4937,N_4749,N_4718);
and U4938 (N_4938,N_4790,N_4786);
nand U4939 (N_4939,N_4628,N_4668);
and U4940 (N_4940,N_4675,N_4639);
xor U4941 (N_4941,N_4724,N_4655);
nand U4942 (N_4942,N_4752,N_4634);
nor U4943 (N_4943,N_4699,N_4668);
nor U4944 (N_4944,N_4751,N_4746);
or U4945 (N_4945,N_4686,N_4653);
and U4946 (N_4946,N_4726,N_4771);
nor U4947 (N_4947,N_4666,N_4679);
or U4948 (N_4948,N_4689,N_4615);
nand U4949 (N_4949,N_4627,N_4608);
and U4950 (N_4950,N_4736,N_4782);
nand U4951 (N_4951,N_4787,N_4665);
nand U4952 (N_4952,N_4601,N_4733);
or U4953 (N_4953,N_4692,N_4739);
and U4954 (N_4954,N_4749,N_4604);
nand U4955 (N_4955,N_4693,N_4665);
or U4956 (N_4956,N_4690,N_4611);
or U4957 (N_4957,N_4619,N_4713);
or U4958 (N_4958,N_4761,N_4777);
nor U4959 (N_4959,N_4793,N_4614);
or U4960 (N_4960,N_4749,N_4685);
xnor U4961 (N_4961,N_4768,N_4673);
and U4962 (N_4962,N_4776,N_4653);
nor U4963 (N_4963,N_4764,N_4680);
and U4964 (N_4964,N_4700,N_4690);
nand U4965 (N_4965,N_4636,N_4779);
and U4966 (N_4966,N_4641,N_4655);
nor U4967 (N_4967,N_4746,N_4769);
or U4968 (N_4968,N_4708,N_4697);
nor U4969 (N_4969,N_4670,N_4750);
nand U4970 (N_4970,N_4706,N_4720);
nand U4971 (N_4971,N_4645,N_4783);
nand U4972 (N_4972,N_4772,N_4640);
nand U4973 (N_4973,N_4653,N_4691);
and U4974 (N_4974,N_4669,N_4635);
and U4975 (N_4975,N_4628,N_4610);
nand U4976 (N_4976,N_4743,N_4744);
and U4977 (N_4977,N_4731,N_4627);
nor U4978 (N_4978,N_4738,N_4601);
and U4979 (N_4979,N_4665,N_4790);
nand U4980 (N_4980,N_4615,N_4693);
nor U4981 (N_4981,N_4783,N_4660);
or U4982 (N_4982,N_4675,N_4648);
nor U4983 (N_4983,N_4694,N_4784);
or U4984 (N_4984,N_4747,N_4660);
and U4985 (N_4985,N_4643,N_4668);
nand U4986 (N_4986,N_4743,N_4609);
or U4987 (N_4987,N_4670,N_4720);
nor U4988 (N_4988,N_4674,N_4733);
or U4989 (N_4989,N_4671,N_4666);
nand U4990 (N_4990,N_4719,N_4716);
and U4991 (N_4991,N_4769,N_4602);
nor U4992 (N_4992,N_4641,N_4688);
or U4993 (N_4993,N_4747,N_4799);
nand U4994 (N_4994,N_4677,N_4704);
nand U4995 (N_4995,N_4740,N_4765);
and U4996 (N_4996,N_4709,N_4755);
nor U4997 (N_4997,N_4738,N_4609);
nor U4998 (N_4998,N_4676,N_4723);
nand U4999 (N_4999,N_4698,N_4742);
nor UO_0 (O_0,N_4913,N_4961);
or UO_1 (O_1,N_4868,N_4859);
nand UO_2 (O_2,N_4890,N_4878);
nand UO_3 (O_3,N_4843,N_4911);
or UO_4 (O_4,N_4864,N_4821);
nand UO_5 (O_5,N_4965,N_4819);
nor UO_6 (O_6,N_4930,N_4809);
or UO_7 (O_7,N_4866,N_4900);
and UO_8 (O_8,N_4826,N_4899);
or UO_9 (O_9,N_4943,N_4835);
and UO_10 (O_10,N_4901,N_4855);
nor UO_11 (O_11,N_4974,N_4823);
nand UO_12 (O_12,N_4937,N_4877);
nand UO_13 (O_13,N_4895,N_4801);
or UO_14 (O_14,N_4882,N_4828);
or UO_15 (O_15,N_4825,N_4894);
or UO_16 (O_16,N_4947,N_4881);
and UO_17 (O_17,N_4939,N_4910);
or UO_18 (O_18,N_4898,N_4906);
or UO_19 (O_19,N_4852,N_4812);
nor UO_20 (O_20,N_4970,N_4936);
nor UO_21 (O_21,N_4805,N_4872);
nand UO_22 (O_22,N_4811,N_4917);
and UO_23 (O_23,N_4827,N_4952);
or UO_24 (O_24,N_4922,N_4946);
or UO_25 (O_25,N_4967,N_4973);
nor UO_26 (O_26,N_4863,N_4953);
nand UO_27 (O_27,N_4839,N_4888);
and UO_28 (O_28,N_4975,N_4954);
and UO_29 (O_29,N_4813,N_4912);
nand UO_30 (O_30,N_4807,N_4822);
and UO_31 (O_31,N_4981,N_4892);
and UO_32 (O_32,N_4842,N_4870);
nand UO_33 (O_33,N_4982,N_4902);
or UO_34 (O_34,N_4833,N_4932);
or UO_35 (O_35,N_4847,N_4924);
nand UO_36 (O_36,N_4921,N_4829);
and UO_37 (O_37,N_4925,N_4968);
or UO_38 (O_38,N_4830,N_4996);
or UO_39 (O_39,N_4966,N_4986);
or UO_40 (O_40,N_4923,N_4824);
nand UO_41 (O_41,N_4960,N_4927);
and UO_42 (O_42,N_4950,N_4958);
and UO_43 (O_43,N_4942,N_4959);
or UO_44 (O_44,N_4837,N_4919);
or UO_45 (O_45,N_4834,N_4831);
xnor UO_46 (O_46,N_4934,N_4893);
or UO_47 (O_47,N_4991,N_4955);
nand UO_48 (O_48,N_4978,N_4860);
nor UO_49 (O_49,N_4818,N_4886);
nor UO_50 (O_50,N_4814,N_4815);
and UO_51 (O_51,N_4940,N_4997);
nor UO_52 (O_52,N_4883,N_4979);
and UO_53 (O_53,N_4887,N_4989);
xor UO_54 (O_54,N_4964,N_4915);
nand UO_55 (O_55,N_4841,N_4856);
nor UO_56 (O_56,N_4914,N_4971);
nand UO_57 (O_57,N_4916,N_4990);
nand UO_58 (O_58,N_4820,N_4846);
and UO_59 (O_59,N_4988,N_4869);
nor UO_60 (O_60,N_4963,N_4817);
or UO_61 (O_61,N_4929,N_4832);
nor UO_62 (O_62,N_4999,N_4836);
and UO_63 (O_63,N_4951,N_4897);
nor UO_64 (O_64,N_4962,N_4920);
or UO_65 (O_65,N_4987,N_4972);
nor UO_66 (O_66,N_4994,N_4861);
nand UO_67 (O_67,N_4876,N_4858);
nor UO_68 (O_68,N_4851,N_4867);
or UO_69 (O_69,N_4875,N_4945);
nand UO_70 (O_70,N_4984,N_4879);
nor UO_71 (O_71,N_4905,N_4896);
nor UO_72 (O_72,N_4845,N_4992);
nand UO_73 (O_73,N_4800,N_4880);
and UO_74 (O_74,N_4926,N_4844);
or UO_75 (O_75,N_4816,N_4865);
and UO_76 (O_76,N_4884,N_4810);
nor UO_77 (O_77,N_4849,N_4903);
nand UO_78 (O_78,N_4909,N_4993);
or UO_79 (O_79,N_4980,N_4804);
and UO_80 (O_80,N_4969,N_4806);
and UO_81 (O_81,N_4857,N_4891);
nor UO_82 (O_82,N_4853,N_4854);
or UO_83 (O_83,N_4941,N_4977);
nand UO_84 (O_84,N_4983,N_4848);
and UO_85 (O_85,N_4948,N_4873);
or UO_86 (O_86,N_4956,N_4957);
nor UO_87 (O_87,N_4933,N_4802);
nand UO_88 (O_88,N_4907,N_4998);
nand UO_89 (O_89,N_4976,N_4904);
nor UO_90 (O_90,N_4944,N_4808);
or UO_91 (O_91,N_4949,N_4874);
nand UO_92 (O_92,N_4871,N_4803);
nor UO_93 (O_93,N_4931,N_4935);
and UO_94 (O_94,N_4885,N_4862);
or UO_95 (O_95,N_4995,N_4928);
or UO_96 (O_96,N_4938,N_4838);
or UO_97 (O_97,N_4889,N_4918);
and UO_98 (O_98,N_4908,N_4840);
nand UO_99 (O_99,N_4985,N_4850);
or UO_100 (O_100,N_4966,N_4917);
and UO_101 (O_101,N_4881,N_4844);
or UO_102 (O_102,N_4919,N_4911);
nor UO_103 (O_103,N_4968,N_4804);
nand UO_104 (O_104,N_4925,N_4833);
nand UO_105 (O_105,N_4804,N_4967);
and UO_106 (O_106,N_4869,N_4920);
and UO_107 (O_107,N_4901,N_4909);
nand UO_108 (O_108,N_4884,N_4973);
or UO_109 (O_109,N_4833,N_4810);
nand UO_110 (O_110,N_4930,N_4812);
and UO_111 (O_111,N_4821,N_4934);
nand UO_112 (O_112,N_4805,N_4913);
nor UO_113 (O_113,N_4885,N_4898);
nand UO_114 (O_114,N_4983,N_4994);
nand UO_115 (O_115,N_4895,N_4823);
nor UO_116 (O_116,N_4938,N_4880);
nor UO_117 (O_117,N_4935,N_4855);
nor UO_118 (O_118,N_4826,N_4932);
or UO_119 (O_119,N_4967,N_4837);
or UO_120 (O_120,N_4921,N_4981);
nor UO_121 (O_121,N_4939,N_4898);
nand UO_122 (O_122,N_4873,N_4884);
and UO_123 (O_123,N_4923,N_4819);
nand UO_124 (O_124,N_4822,N_4937);
and UO_125 (O_125,N_4900,N_4927);
or UO_126 (O_126,N_4846,N_4960);
nor UO_127 (O_127,N_4912,N_4929);
and UO_128 (O_128,N_4883,N_4983);
nor UO_129 (O_129,N_4962,N_4812);
and UO_130 (O_130,N_4893,N_4949);
and UO_131 (O_131,N_4861,N_4920);
nor UO_132 (O_132,N_4908,N_4842);
nand UO_133 (O_133,N_4929,N_4954);
and UO_134 (O_134,N_4886,N_4893);
nand UO_135 (O_135,N_4888,N_4960);
or UO_136 (O_136,N_4802,N_4973);
nor UO_137 (O_137,N_4956,N_4968);
nor UO_138 (O_138,N_4885,N_4901);
and UO_139 (O_139,N_4877,N_4872);
or UO_140 (O_140,N_4813,N_4933);
nor UO_141 (O_141,N_4817,N_4927);
and UO_142 (O_142,N_4991,N_4849);
nor UO_143 (O_143,N_4861,N_4961);
and UO_144 (O_144,N_4920,N_4955);
nor UO_145 (O_145,N_4966,N_4894);
nor UO_146 (O_146,N_4870,N_4844);
and UO_147 (O_147,N_4959,N_4957);
nand UO_148 (O_148,N_4857,N_4991);
and UO_149 (O_149,N_4976,N_4833);
nor UO_150 (O_150,N_4944,N_4904);
and UO_151 (O_151,N_4863,N_4989);
xnor UO_152 (O_152,N_4979,N_4900);
nand UO_153 (O_153,N_4988,N_4829);
and UO_154 (O_154,N_4878,N_4853);
and UO_155 (O_155,N_4801,N_4833);
nor UO_156 (O_156,N_4922,N_4836);
nand UO_157 (O_157,N_4850,N_4825);
or UO_158 (O_158,N_4839,N_4970);
nand UO_159 (O_159,N_4818,N_4989);
nand UO_160 (O_160,N_4914,N_4804);
nand UO_161 (O_161,N_4900,N_4913);
nand UO_162 (O_162,N_4848,N_4959);
or UO_163 (O_163,N_4967,N_4886);
or UO_164 (O_164,N_4937,N_4914);
or UO_165 (O_165,N_4979,N_4946);
nor UO_166 (O_166,N_4873,N_4823);
nor UO_167 (O_167,N_4828,N_4881);
nand UO_168 (O_168,N_4851,N_4854);
nand UO_169 (O_169,N_4845,N_4871);
and UO_170 (O_170,N_4874,N_4969);
nor UO_171 (O_171,N_4934,N_4857);
and UO_172 (O_172,N_4892,N_4952);
nor UO_173 (O_173,N_4817,N_4979);
and UO_174 (O_174,N_4917,N_4853);
xnor UO_175 (O_175,N_4940,N_4812);
nand UO_176 (O_176,N_4944,N_4984);
or UO_177 (O_177,N_4985,N_4963);
and UO_178 (O_178,N_4809,N_4813);
nand UO_179 (O_179,N_4897,N_4809);
xor UO_180 (O_180,N_4970,N_4931);
nand UO_181 (O_181,N_4854,N_4806);
and UO_182 (O_182,N_4867,N_4874);
nand UO_183 (O_183,N_4802,N_4875);
nor UO_184 (O_184,N_4836,N_4918);
nand UO_185 (O_185,N_4953,N_4900);
nor UO_186 (O_186,N_4938,N_4829);
nor UO_187 (O_187,N_4829,N_4962);
or UO_188 (O_188,N_4842,N_4983);
or UO_189 (O_189,N_4963,N_4881);
nand UO_190 (O_190,N_4820,N_4823);
or UO_191 (O_191,N_4972,N_4965);
and UO_192 (O_192,N_4922,N_4980);
nand UO_193 (O_193,N_4814,N_4962);
and UO_194 (O_194,N_4901,N_4978);
or UO_195 (O_195,N_4976,N_4827);
nand UO_196 (O_196,N_4977,N_4908);
or UO_197 (O_197,N_4954,N_4825);
nand UO_198 (O_198,N_4887,N_4843);
nand UO_199 (O_199,N_4959,N_4812);
nand UO_200 (O_200,N_4975,N_4869);
nor UO_201 (O_201,N_4872,N_4854);
nor UO_202 (O_202,N_4809,N_4893);
nor UO_203 (O_203,N_4897,N_4928);
or UO_204 (O_204,N_4976,N_4855);
nor UO_205 (O_205,N_4903,N_4973);
and UO_206 (O_206,N_4924,N_4898);
nand UO_207 (O_207,N_4870,N_4943);
and UO_208 (O_208,N_4933,N_4885);
or UO_209 (O_209,N_4833,N_4959);
nand UO_210 (O_210,N_4898,N_4963);
nor UO_211 (O_211,N_4802,N_4948);
and UO_212 (O_212,N_4840,N_4809);
or UO_213 (O_213,N_4994,N_4933);
nand UO_214 (O_214,N_4857,N_4815);
nand UO_215 (O_215,N_4910,N_4820);
or UO_216 (O_216,N_4909,N_4900);
nor UO_217 (O_217,N_4994,N_4970);
nand UO_218 (O_218,N_4810,N_4866);
nor UO_219 (O_219,N_4929,N_4934);
and UO_220 (O_220,N_4815,N_4825);
nand UO_221 (O_221,N_4959,N_4949);
nand UO_222 (O_222,N_4841,N_4951);
nand UO_223 (O_223,N_4937,N_4845);
and UO_224 (O_224,N_4939,N_4938);
or UO_225 (O_225,N_4930,N_4974);
or UO_226 (O_226,N_4962,N_4838);
or UO_227 (O_227,N_4910,N_4875);
and UO_228 (O_228,N_4994,N_4880);
nand UO_229 (O_229,N_4809,N_4802);
nand UO_230 (O_230,N_4887,N_4851);
and UO_231 (O_231,N_4940,N_4875);
and UO_232 (O_232,N_4911,N_4996);
or UO_233 (O_233,N_4867,N_4806);
and UO_234 (O_234,N_4934,N_4870);
or UO_235 (O_235,N_4998,N_4801);
or UO_236 (O_236,N_4814,N_4836);
nor UO_237 (O_237,N_4808,N_4875);
nor UO_238 (O_238,N_4865,N_4891);
nand UO_239 (O_239,N_4953,N_4956);
or UO_240 (O_240,N_4982,N_4950);
or UO_241 (O_241,N_4927,N_4929);
and UO_242 (O_242,N_4977,N_4810);
nor UO_243 (O_243,N_4848,N_4908);
and UO_244 (O_244,N_4878,N_4842);
nor UO_245 (O_245,N_4894,N_4900);
nor UO_246 (O_246,N_4873,N_4822);
or UO_247 (O_247,N_4987,N_4958);
nor UO_248 (O_248,N_4889,N_4949);
or UO_249 (O_249,N_4921,N_4832);
and UO_250 (O_250,N_4952,N_4841);
nand UO_251 (O_251,N_4946,N_4859);
and UO_252 (O_252,N_4847,N_4852);
nor UO_253 (O_253,N_4983,N_4966);
and UO_254 (O_254,N_4801,N_4887);
and UO_255 (O_255,N_4821,N_4982);
or UO_256 (O_256,N_4971,N_4906);
nand UO_257 (O_257,N_4870,N_4929);
nor UO_258 (O_258,N_4951,N_4974);
nand UO_259 (O_259,N_4945,N_4998);
nor UO_260 (O_260,N_4846,N_4863);
nor UO_261 (O_261,N_4989,N_4990);
nor UO_262 (O_262,N_4895,N_4887);
nor UO_263 (O_263,N_4812,N_4894);
or UO_264 (O_264,N_4866,N_4825);
xor UO_265 (O_265,N_4928,N_4841);
nand UO_266 (O_266,N_4805,N_4961);
and UO_267 (O_267,N_4823,N_4835);
nor UO_268 (O_268,N_4918,N_4890);
nand UO_269 (O_269,N_4966,N_4961);
nand UO_270 (O_270,N_4866,N_4886);
nand UO_271 (O_271,N_4928,N_4989);
nand UO_272 (O_272,N_4833,N_4977);
or UO_273 (O_273,N_4802,N_4986);
nand UO_274 (O_274,N_4863,N_4958);
nand UO_275 (O_275,N_4915,N_4836);
nor UO_276 (O_276,N_4909,N_4946);
xnor UO_277 (O_277,N_4821,N_4834);
or UO_278 (O_278,N_4919,N_4913);
or UO_279 (O_279,N_4841,N_4983);
nand UO_280 (O_280,N_4948,N_4919);
nor UO_281 (O_281,N_4820,N_4960);
nand UO_282 (O_282,N_4930,N_4999);
and UO_283 (O_283,N_4924,N_4841);
nand UO_284 (O_284,N_4825,N_4953);
and UO_285 (O_285,N_4815,N_4949);
or UO_286 (O_286,N_4986,N_4885);
nor UO_287 (O_287,N_4990,N_4828);
and UO_288 (O_288,N_4818,N_4861);
and UO_289 (O_289,N_4986,N_4923);
or UO_290 (O_290,N_4881,N_4926);
nor UO_291 (O_291,N_4960,N_4976);
and UO_292 (O_292,N_4979,N_4836);
nor UO_293 (O_293,N_4924,N_4915);
and UO_294 (O_294,N_4838,N_4877);
and UO_295 (O_295,N_4982,N_4852);
and UO_296 (O_296,N_4806,N_4970);
and UO_297 (O_297,N_4928,N_4843);
and UO_298 (O_298,N_4808,N_4984);
nor UO_299 (O_299,N_4805,N_4948);
nor UO_300 (O_300,N_4885,N_4883);
and UO_301 (O_301,N_4819,N_4908);
or UO_302 (O_302,N_4807,N_4873);
or UO_303 (O_303,N_4816,N_4852);
or UO_304 (O_304,N_4883,N_4887);
nand UO_305 (O_305,N_4996,N_4840);
nand UO_306 (O_306,N_4800,N_4986);
xnor UO_307 (O_307,N_4935,N_4975);
nand UO_308 (O_308,N_4906,N_4998);
or UO_309 (O_309,N_4978,N_4918);
nor UO_310 (O_310,N_4821,N_4801);
or UO_311 (O_311,N_4842,N_4953);
or UO_312 (O_312,N_4871,N_4959);
nand UO_313 (O_313,N_4977,N_4824);
and UO_314 (O_314,N_4831,N_4995);
and UO_315 (O_315,N_4871,N_4973);
or UO_316 (O_316,N_4904,N_4895);
nand UO_317 (O_317,N_4845,N_4851);
or UO_318 (O_318,N_4932,N_4950);
nor UO_319 (O_319,N_4827,N_4807);
nand UO_320 (O_320,N_4941,N_4884);
nand UO_321 (O_321,N_4985,N_4890);
nor UO_322 (O_322,N_4803,N_4961);
or UO_323 (O_323,N_4874,N_4975);
nor UO_324 (O_324,N_4804,N_4806);
nand UO_325 (O_325,N_4895,N_4861);
or UO_326 (O_326,N_4800,N_4949);
nand UO_327 (O_327,N_4816,N_4994);
or UO_328 (O_328,N_4995,N_4983);
or UO_329 (O_329,N_4939,N_4897);
or UO_330 (O_330,N_4860,N_4834);
nor UO_331 (O_331,N_4883,N_4893);
nand UO_332 (O_332,N_4945,N_4836);
or UO_333 (O_333,N_4806,N_4966);
and UO_334 (O_334,N_4916,N_4991);
and UO_335 (O_335,N_4843,N_4858);
and UO_336 (O_336,N_4891,N_4970);
nand UO_337 (O_337,N_4932,N_4957);
and UO_338 (O_338,N_4986,N_4941);
xor UO_339 (O_339,N_4932,N_4831);
or UO_340 (O_340,N_4854,N_4979);
or UO_341 (O_341,N_4945,N_4974);
and UO_342 (O_342,N_4859,N_4816);
nand UO_343 (O_343,N_4857,N_4909);
nand UO_344 (O_344,N_4893,N_4954);
nand UO_345 (O_345,N_4991,N_4889);
nor UO_346 (O_346,N_4845,N_4861);
and UO_347 (O_347,N_4996,N_4820);
and UO_348 (O_348,N_4967,N_4937);
and UO_349 (O_349,N_4854,N_4819);
and UO_350 (O_350,N_4864,N_4932);
nand UO_351 (O_351,N_4811,N_4855);
or UO_352 (O_352,N_4984,N_4922);
and UO_353 (O_353,N_4821,N_4805);
nor UO_354 (O_354,N_4860,N_4821);
xor UO_355 (O_355,N_4885,N_4800);
nand UO_356 (O_356,N_4824,N_4806);
and UO_357 (O_357,N_4989,N_4808);
nand UO_358 (O_358,N_4985,N_4964);
or UO_359 (O_359,N_4849,N_4935);
nor UO_360 (O_360,N_4808,N_4927);
nand UO_361 (O_361,N_4985,N_4954);
nor UO_362 (O_362,N_4930,N_4806);
or UO_363 (O_363,N_4806,N_4990);
nand UO_364 (O_364,N_4874,N_4834);
nand UO_365 (O_365,N_4905,N_4832);
nand UO_366 (O_366,N_4892,N_4951);
or UO_367 (O_367,N_4839,N_4822);
nand UO_368 (O_368,N_4851,N_4902);
and UO_369 (O_369,N_4813,N_4903);
nand UO_370 (O_370,N_4875,N_4830);
or UO_371 (O_371,N_4811,N_4990);
nand UO_372 (O_372,N_4887,N_4978);
nor UO_373 (O_373,N_4835,N_4822);
or UO_374 (O_374,N_4859,N_4808);
or UO_375 (O_375,N_4833,N_4806);
and UO_376 (O_376,N_4899,N_4989);
nor UO_377 (O_377,N_4871,N_4833);
nor UO_378 (O_378,N_4893,N_4860);
and UO_379 (O_379,N_4864,N_4959);
and UO_380 (O_380,N_4998,N_4922);
or UO_381 (O_381,N_4807,N_4845);
and UO_382 (O_382,N_4990,N_4835);
nand UO_383 (O_383,N_4986,N_4921);
nand UO_384 (O_384,N_4850,N_4805);
nand UO_385 (O_385,N_4852,N_4825);
and UO_386 (O_386,N_4842,N_4885);
xor UO_387 (O_387,N_4889,N_4884);
nor UO_388 (O_388,N_4948,N_4803);
nor UO_389 (O_389,N_4829,N_4947);
or UO_390 (O_390,N_4891,N_4987);
nor UO_391 (O_391,N_4938,N_4946);
nor UO_392 (O_392,N_4992,N_4972);
nand UO_393 (O_393,N_4916,N_4954);
or UO_394 (O_394,N_4813,N_4857);
nor UO_395 (O_395,N_4925,N_4932);
or UO_396 (O_396,N_4883,N_4889);
nand UO_397 (O_397,N_4873,N_4918);
or UO_398 (O_398,N_4919,N_4997);
nand UO_399 (O_399,N_4819,N_4879);
nand UO_400 (O_400,N_4965,N_4954);
and UO_401 (O_401,N_4973,N_4855);
nor UO_402 (O_402,N_4885,N_4830);
and UO_403 (O_403,N_4807,N_4880);
nand UO_404 (O_404,N_4813,N_4925);
xor UO_405 (O_405,N_4929,N_4841);
nand UO_406 (O_406,N_4940,N_4986);
and UO_407 (O_407,N_4886,N_4907);
nor UO_408 (O_408,N_4908,N_4975);
and UO_409 (O_409,N_4968,N_4847);
or UO_410 (O_410,N_4802,N_4800);
nor UO_411 (O_411,N_4810,N_4995);
nor UO_412 (O_412,N_4941,N_4993);
or UO_413 (O_413,N_4932,N_4801);
nor UO_414 (O_414,N_4910,N_4816);
nor UO_415 (O_415,N_4904,N_4822);
nand UO_416 (O_416,N_4850,N_4896);
and UO_417 (O_417,N_4962,N_4897);
and UO_418 (O_418,N_4950,N_4979);
and UO_419 (O_419,N_4842,N_4859);
and UO_420 (O_420,N_4952,N_4888);
nor UO_421 (O_421,N_4946,N_4874);
and UO_422 (O_422,N_4859,N_4807);
and UO_423 (O_423,N_4991,N_4859);
nor UO_424 (O_424,N_4959,N_4991);
nand UO_425 (O_425,N_4853,N_4803);
and UO_426 (O_426,N_4992,N_4891);
nor UO_427 (O_427,N_4865,N_4923);
and UO_428 (O_428,N_4939,N_4927);
nor UO_429 (O_429,N_4964,N_4870);
and UO_430 (O_430,N_4800,N_4991);
or UO_431 (O_431,N_4978,N_4886);
nand UO_432 (O_432,N_4817,N_4860);
and UO_433 (O_433,N_4981,N_4849);
and UO_434 (O_434,N_4806,N_4918);
or UO_435 (O_435,N_4872,N_4880);
nand UO_436 (O_436,N_4887,N_4815);
or UO_437 (O_437,N_4906,N_4870);
and UO_438 (O_438,N_4966,N_4853);
and UO_439 (O_439,N_4960,N_4838);
nand UO_440 (O_440,N_4825,N_4831);
nand UO_441 (O_441,N_4872,N_4916);
or UO_442 (O_442,N_4801,N_4892);
nor UO_443 (O_443,N_4977,N_4930);
or UO_444 (O_444,N_4892,N_4988);
and UO_445 (O_445,N_4888,N_4967);
nor UO_446 (O_446,N_4847,N_4923);
and UO_447 (O_447,N_4942,N_4920);
nor UO_448 (O_448,N_4978,N_4991);
and UO_449 (O_449,N_4976,N_4928);
and UO_450 (O_450,N_4875,N_4951);
and UO_451 (O_451,N_4935,N_4912);
and UO_452 (O_452,N_4954,N_4805);
nand UO_453 (O_453,N_4824,N_4950);
or UO_454 (O_454,N_4968,N_4924);
nor UO_455 (O_455,N_4833,N_4875);
nor UO_456 (O_456,N_4857,N_4803);
nand UO_457 (O_457,N_4932,N_4897);
and UO_458 (O_458,N_4849,N_4887);
and UO_459 (O_459,N_4872,N_4853);
nand UO_460 (O_460,N_4896,N_4846);
or UO_461 (O_461,N_4861,N_4836);
nand UO_462 (O_462,N_4850,N_4816);
nand UO_463 (O_463,N_4872,N_4947);
or UO_464 (O_464,N_4972,N_4949);
or UO_465 (O_465,N_4916,N_4917);
nand UO_466 (O_466,N_4972,N_4874);
and UO_467 (O_467,N_4988,N_4902);
nor UO_468 (O_468,N_4856,N_4814);
and UO_469 (O_469,N_4889,N_4830);
and UO_470 (O_470,N_4861,N_4941);
nor UO_471 (O_471,N_4886,N_4995);
nand UO_472 (O_472,N_4805,N_4883);
and UO_473 (O_473,N_4963,N_4845);
nand UO_474 (O_474,N_4846,N_4881);
and UO_475 (O_475,N_4864,N_4869);
or UO_476 (O_476,N_4982,N_4891);
or UO_477 (O_477,N_4982,N_4849);
and UO_478 (O_478,N_4861,N_4919);
or UO_479 (O_479,N_4867,N_4907);
and UO_480 (O_480,N_4832,N_4954);
and UO_481 (O_481,N_4907,N_4972);
nand UO_482 (O_482,N_4804,N_4885);
and UO_483 (O_483,N_4832,N_4875);
nand UO_484 (O_484,N_4808,N_4979);
and UO_485 (O_485,N_4987,N_4955);
nand UO_486 (O_486,N_4897,N_4904);
or UO_487 (O_487,N_4806,N_4982);
nor UO_488 (O_488,N_4997,N_4910);
nor UO_489 (O_489,N_4901,N_4917);
or UO_490 (O_490,N_4918,N_4907);
nor UO_491 (O_491,N_4835,N_4986);
and UO_492 (O_492,N_4915,N_4916);
and UO_493 (O_493,N_4864,N_4975);
nand UO_494 (O_494,N_4904,N_4830);
nand UO_495 (O_495,N_4808,N_4946);
and UO_496 (O_496,N_4803,N_4841);
nand UO_497 (O_497,N_4974,N_4820);
nand UO_498 (O_498,N_4837,N_4920);
and UO_499 (O_499,N_4999,N_4885);
nor UO_500 (O_500,N_4817,N_4894);
and UO_501 (O_501,N_4904,N_4812);
and UO_502 (O_502,N_4951,N_4862);
nor UO_503 (O_503,N_4874,N_4928);
or UO_504 (O_504,N_4836,N_4816);
nand UO_505 (O_505,N_4998,N_4851);
nand UO_506 (O_506,N_4892,N_4923);
and UO_507 (O_507,N_4924,N_4812);
nand UO_508 (O_508,N_4911,N_4981);
nor UO_509 (O_509,N_4989,N_4910);
nor UO_510 (O_510,N_4913,N_4820);
nor UO_511 (O_511,N_4910,N_4894);
nand UO_512 (O_512,N_4959,N_4932);
or UO_513 (O_513,N_4981,N_4894);
nor UO_514 (O_514,N_4823,N_4838);
and UO_515 (O_515,N_4917,N_4860);
and UO_516 (O_516,N_4936,N_4821);
nor UO_517 (O_517,N_4978,N_4892);
or UO_518 (O_518,N_4953,N_4901);
nor UO_519 (O_519,N_4823,N_4854);
nand UO_520 (O_520,N_4900,N_4942);
and UO_521 (O_521,N_4954,N_4953);
or UO_522 (O_522,N_4845,N_4842);
nor UO_523 (O_523,N_4850,N_4845);
or UO_524 (O_524,N_4809,N_4860);
and UO_525 (O_525,N_4915,N_4878);
or UO_526 (O_526,N_4916,N_4993);
nand UO_527 (O_527,N_4807,N_4913);
nor UO_528 (O_528,N_4886,N_4872);
nor UO_529 (O_529,N_4836,N_4931);
or UO_530 (O_530,N_4868,N_4991);
nor UO_531 (O_531,N_4887,N_4878);
and UO_532 (O_532,N_4991,N_4829);
and UO_533 (O_533,N_4918,N_4815);
or UO_534 (O_534,N_4846,N_4823);
and UO_535 (O_535,N_4885,N_4926);
or UO_536 (O_536,N_4976,N_4822);
nor UO_537 (O_537,N_4820,N_4981);
and UO_538 (O_538,N_4875,N_4846);
nand UO_539 (O_539,N_4977,N_4881);
and UO_540 (O_540,N_4925,N_4907);
nor UO_541 (O_541,N_4925,N_4880);
and UO_542 (O_542,N_4955,N_4906);
and UO_543 (O_543,N_4834,N_4869);
and UO_544 (O_544,N_4896,N_4815);
nor UO_545 (O_545,N_4896,N_4904);
and UO_546 (O_546,N_4824,N_4994);
and UO_547 (O_547,N_4812,N_4955);
and UO_548 (O_548,N_4805,N_4863);
nor UO_549 (O_549,N_4885,N_4915);
nor UO_550 (O_550,N_4954,N_4874);
nor UO_551 (O_551,N_4846,N_4975);
and UO_552 (O_552,N_4882,N_4922);
or UO_553 (O_553,N_4835,N_4848);
or UO_554 (O_554,N_4835,N_4903);
and UO_555 (O_555,N_4981,N_4901);
nor UO_556 (O_556,N_4841,N_4974);
or UO_557 (O_557,N_4890,N_4828);
nor UO_558 (O_558,N_4917,N_4874);
nand UO_559 (O_559,N_4906,N_4949);
nor UO_560 (O_560,N_4864,N_4964);
nor UO_561 (O_561,N_4918,N_4830);
or UO_562 (O_562,N_4932,N_4935);
nand UO_563 (O_563,N_4946,N_4991);
or UO_564 (O_564,N_4926,N_4925);
or UO_565 (O_565,N_4891,N_4896);
nor UO_566 (O_566,N_4992,N_4955);
nand UO_567 (O_567,N_4955,N_4864);
nor UO_568 (O_568,N_4881,N_4819);
and UO_569 (O_569,N_4914,N_4934);
nand UO_570 (O_570,N_4909,N_4839);
nand UO_571 (O_571,N_4887,N_4901);
and UO_572 (O_572,N_4912,N_4905);
and UO_573 (O_573,N_4984,N_4856);
nor UO_574 (O_574,N_4961,N_4838);
or UO_575 (O_575,N_4888,N_4981);
nand UO_576 (O_576,N_4950,N_4973);
and UO_577 (O_577,N_4858,N_4900);
and UO_578 (O_578,N_4804,N_4970);
and UO_579 (O_579,N_4912,N_4848);
nand UO_580 (O_580,N_4876,N_4833);
and UO_581 (O_581,N_4814,N_4837);
and UO_582 (O_582,N_4811,N_4871);
nand UO_583 (O_583,N_4855,N_4909);
nor UO_584 (O_584,N_4963,N_4989);
nor UO_585 (O_585,N_4899,N_4805);
nor UO_586 (O_586,N_4827,N_4911);
nand UO_587 (O_587,N_4929,N_4931);
or UO_588 (O_588,N_4918,N_4863);
nand UO_589 (O_589,N_4892,N_4817);
nand UO_590 (O_590,N_4909,N_4808);
or UO_591 (O_591,N_4961,N_4833);
nor UO_592 (O_592,N_4889,N_4961);
nand UO_593 (O_593,N_4800,N_4904);
and UO_594 (O_594,N_4842,N_4806);
nor UO_595 (O_595,N_4854,N_4923);
nand UO_596 (O_596,N_4962,N_4956);
or UO_597 (O_597,N_4905,N_4986);
xnor UO_598 (O_598,N_4827,N_4894);
or UO_599 (O_599,N_4936,N_4955);
nor UO_600 (O_600,N_4922,N_4923);
and UO_601 (O_601,N_4830,N_4976);
or UO_602 (O_602,N_4876,N_4995);
or UO_603 (O_603,N_4846,N_4885);
nand UO_604 (O_604,N_4867,N_4810);
nand UO_605 (O_605,N_4882,N_4824);
nand UO_606 (O_606,N_4948,N_4927);
nor UO_607 (O_607,N_4947,N_4892);
or UO_608 (O_608,N_4842,N_4990);
and UO_609 (O_609,N_4892,N_4914);
and UO_610 (O_610,N_4810,N_4882);
and UO_611 (O_611,N_4867,N_4832);
nor UO_612 (O_612,N_4806,N_4950);
nand UO_613 (O_613,N_4838,N_4926);
or UO_614 (O_614,N_4997,N_4925);
or UO_615 (O_615,N_4926,N_4826);
nand UO_616 (O_616,N_4856,N_4857);
or UO_617 (O_617,N_4894,N_4830);
and UO_618 (O_618,N_4976,N_4942);
and UO_619 (O_619,N_4816,N_4987);
or UO_620 (O_620,N_4862,N_4910);
nor UO_621 (O_621,N_4952,N_4823);
nor UO_622 (O_622,N_4999,N_4955);
nand UO_623 (O_623,N_4849,N_4928);
and UO_624 (O_624,N_4848,N_4863);
or UO_625 (O_625,N_4961,N_4882);
and UO_626 (O_626,N_4897,N_4816);
nor UO_627 (O_627,N_4994,N_4979);
or UO_628 (O_628,N_4955,N_4840);
xor UO_629 (O_629,N_4957,N_4885);
and UO_630 (O_630,N_4996,N_4907);
nand UO_631 (O_631,N_4833,N_4849);
and UO_632 (O_632,N_4847,N_4917);
nor UO_633 (O_633,N_4807,N_4942);
or UO_634 (O_634,N_4961,N_4881);
and UO_635 (O_635,N_4920,N_4886);
and UO_636 (O_636,N_4934,N_4815);
and UO_637 (O_637,N_4926,N_4919);
nand UO_638 (O_638,N_4920,N_4944);
or UO_639 (O_639,N_4893,N_4835);
and UO_640 (O_640,N_4923,N_4811);
nor UO_641 (O_641,N_4836,N_4942);
nor UO_642 (O_642,N_4979,N_4976);
or UO_643 (O_643,N_4864,N_4844);
or UO_644 (O_644,N_4997,N_4952);
and UO_645 (O_645,N_4851,N_4883);
nor UO_646 (O_646,N_4814,N_4983);
nor UO_647 (O_647,N_4967,N_4958);
and UO_648 (O_648,N_4844,N_4804);
or UO_649 (O_649,N_4999,N_4851);
nand UO_650 (O_650,N_4898,N_4813);
and UO_651 (O_651,N_4827,N_4833);
or UO_652 (O_652,N_4919,N_4820);
nand UO_653 (O_653,N_4825,N_4941);
nand UO_654 (O_654,N_4974,N_4939);
or UO_655 (O_655,N_4936,N_4842);
and UO_656 (O_656,N_4983,N_4977);
nor UO_657 (O_657,N_4979,N_4834);
nor UO_658 (O_658,N_4827,N_4892);
or UO_659 (O_659,N_4804,N_4826);
and UO_660 (O_660,N_4883,N_4816);
and UO_661 (O_661,N_4880,N_4869);
nor UO_662 (O_662,N_4929,N_4849);
xor UO_663 (O_663,N_4978,N_4880);
and UO_664 (O_664,N_4995,N_4890);
or UO_665 (O_665,N_4928,N_4988);
and UO_666 (O_666,N_4913,N_4872);
nor UO_667 (O_667,N_4988,N_4824);
and UO_668 (O_668,N_4870,N_4873);
nor UO_669 (O_669,N_4953,N_4933);
and UO_670 (O_670,N_4804,N_4845);
nor UO_671 (O_671,N_4806,N_4926);
or UO_672 (O_672,N_4918,N_4971);
or UO_673 (O_673,N_4876,N_4986);
xor UO_674 (O_674,N_4856,N_4969);
and UO_675 (O_675,N_4925,N_4920);
and UO_676 (O_676,N_4800,N_4826);
nand UO_677 (O_677,N_4988,N_4887);
and UO_678 (O_678,N_4902,N_4821);
nor UO_679 (O_679,N_4857,N_4904);
or UO_680 (O_680,N_4912,N_4956);
or UO_681 (O_681,N_4803,N_4817);
nand UO_682 (O_682,N_4911,N_4871);
or UO_683 (O_683,N_4947,N_4993);
and UO_684 (O_684,N_4952,N_4873);
nand UO_685 (O_685,N_4974,N_4824);
nor UO_686 (O_686,N_4806,N_4846);
nand UO_687 (O_687,N_4869,N_4961);
nand UO_688 (O_688,N_4917,N_4899);
nor UO_689 (O_689,N_4906,N_4944);
nor UO_690 (O_690,N_4966,N_4946);
nor UO_691 (O_691,N_4829,N_4878);
or UO_692 (O_692,N_4867,N_4953);
nor UO_693 (O_693,N_4829,N_4979);
nor UO_694 (O_694,N_4918,N_4822);
and UO_695 (O_695,N_4858,N_4863);
nand UO_696 (O_696,N_4967,N_4999);
or UO_697 (O_697,N_4900,N_4872);
nand UO_698 (O_698,N_4875,N_4822);
and UO_699 (O_699,N_4889,N_4835);
or UO_700 (O_700,N_4965,N_4809);
nor UO_701 (O_701,N_4835,N_4809);
or UO_702 (O_702,N_4823,N_4824);
nand UO_703 (O_703,N_4984,N_4958);
nand UO_704 (O_704,N_4951,N_4979);
nand UO_705 (O_705,N_4835,N_4914);
or UO_706 (O_706,N_4845,N_4951);
nor UO_707 (O_707,N_4930,N_4970);
nor UO_708 (O_708,N_4912,N_4807);
nor UO_709 (O_709,N_4893,N_4952);
and UO_710 (O_710,N_4866,N_4809);
nor UO_711 (O_711,N_4812,N_4980);
nor UO_712 (O_712,N_4915,N_4830);
nor UO_713 (O_713,N_4947,N_4926);
nor UO_714 (O_714,N_4823,N_4926);
and UO_715 (O_715,N_4925,N_4893);
nor UO_716 (O_716,N_4866,N_4884);
nor UO_717 (O_717,N_4857,N_4959);
or UO_718 (O_718,N_4961,N_4830);
nor UO_719 (O_719,N_4961,N_4988);
nand UO_720 (O_720,N_4999,N_4979);
and UO_721 (O_721,N_4818,N_4954);
and UO_722 (O_722,N_4820,N_4887);
xor UO_723 (O_723,N_4939,N_4851);
and UO_724 (O_724,N_4807,N_4865);
nand UO_725 (O_725,N_4944,N_4954);
nor UO_726 (O_726,N_4830,N_4880);
nand UO_727 (O_727,N_4997,N_4969);
nor UO_728 (O_728,N_4807,N_4922);
or UO_729 (O_729,N_4853,N_4855);
nand UO_730 (O_730,N_4909,N_4934);
nand UO_731 (O_731,N_4905,N_4974);
nor UO_732 (O_732,N_4950,N_4885);
nor UO_733 (O_733,N_4852,N_4851);
and UO_734 (O_734,N_4940,N_4932);
nand UO_735 (O_735,N_4879,N_4955);
or UO_736 (O_736,N_4936,N_4882);
and UO_737 (O_737,N_4959,N_4860);
and UO_738 (O_738,N_4972,N_4879);
or UO_739 (O_739,N_4921,N_4924);
nor UO_740 (O_740,N_4949,N_4821);
and UO_741 (O_741,N_4966,N_4857);
or UO_742 (O_742,N_4916,N_4926);
or UO_743 (O_743,N_4829,N_4956);
or UO_744 (O_744,N_4833,N_4909);
nand UO_745 (O_745,N_4991,N_4818);
and UO_746 (O_746,N_4805,N_4857);
nor UO_747 (O_747,N_4900,N_4855);
or UO_748 (O_748,N_4995,N_4930);
and UO_749 (O_749,N_4939,N_4904);
nor UO_750 (O_750,N_4922,N_4909);
and UO_751 (O_751,N_4945,N_4947);
or UO_752 (O_752,N_4887,N_4864);
nor UO_753 (O_753,N_4996,N_4992);
or UO_754 (O_754,N_4948,N_4979);
nand UO_755 (O_755,N_4955,N_4907);
and UO_756 (O_756,N_4824,N_4860);
nand UO_757 (O_757,N_4977,N_4912);
or UO_758 (O_758,N_4918,N_4876);
or UO_759 (O_759,N_4838,N_4933);
and UO_760 (O_760,N_4836,N_4841);
or UO_761 (O_761,N_4812,N_4893);
nor UO_762 (O_762,N_4904,N_4890);
or UO_763 (O_763,N_4997,N_4889);
nor UO_764 (O_764,N_4961,N_4866);
nand UO_765 (O_765,N_4908,N_4923);
nand UO_766 (O_766,N_4974,N_4855);
or UO_767 (O_767,N_4984,N_4892);
or UO_768 (O_768,N_4820,N_4896);
or UO_769 (O_769,N_4911,N_4831);
or UO_770 (O_770,N_4896,N_4911);
and UO_771 (O_771,N_4936,N_4918);
nand UO_772 (O_772,N_4834,N_4858);
and UO_773 (O_773,N_4980,N_4972);
nand UO_774 (O_774,N_4863,N_4908);
or UO_775 (O_775,N_4967,N_4951);
nor UO_776 (O_776,N_4912,N_4845);
nor UO_777 (O_777,N_4940,N_4985);
nand UO_778 (O_778,N_4861,N_4834);
and UO_779 (O_779,N_4955,N_4924);
nand UO_780 (O_780,N_4998,N_4881);
or UO_781 (O_781,N_4858,N_4884);
nor UO_782 (O_782,N_4884,N_4948);
xnor UO_783 (O_783,N_4808,N_4815);
nand UO_784 (O_784,N_4953,N_4829);
nor UO_785 (O_785,N_4915,N_4902);
and UO_786 (O_786,N_4832,N_4804);
or UO_787 (O_787,N_4837,N_4936);
or UO_788 (O_788,N_4965,N_4881);
and UO_789 (O_789,N_4967,N_4823);
xnor UO_790 (O_790,N_4967,N_4847);
or UO_791 (O_791,N_4887,N_4830);
and UO_792 (O_792,N_4810,N_4845);
and UO_793 (O_793,N_4922,N_4901);
nand UO_794 (O_794,N_4892,N_4882);
nor UO_795 (O_795,N_4898,N_4981);
xnor UO_796 (O_796,N_4831,N_4960);
and UO_797 (O_797,N_4831,N_4871);
nor UO_798 (O_798,N_4869,N_4873);
nand UO_799 (O_799,N_4917,N_4878);
or UO_800 (O_800,N_4981,N_4827);
nor UO_801 (O_801,N_4873,N_4976);
nand UO_802 (O_802,N_4963,N_4919);
and UO_803 (O_803,N_4949,N_4905);
or UO_804 (O_804,N_4818,N_4812);
or UO_805 (O_805,N_4839,N_4976);
nor UO_806 (O_806,N_4984,N_4805);
and UO_807 (O_807,N_4803,N_4922);
and UO_808 (O_808,N_4976,N_4808);
or UO_809 (O_809,N_4812,N_4804);
and UO_810 (O_810,N_4929,N_4817);
or UO_811 (O_811,N_4918,N_4852);
or UO_812 (O_812,N_4895,N_4831);
nand UO_813 (O_813,N_4828,N_4910);
nor UO_814 (O_814,N_4813,N_4900);
or UO_815 (O_815,N_4945,N_4876);
nor UO_816 (O_816,N_4880,N_4951);
nor UO_817 (O_817,N_4938,N_4983);
or UO_818 (O_818,N_4989,N_4885);
and UO_819 (O_819,N_4821,N_4907);
nor UO_820 (O_820,N_4836,N_4960);
nand UO_821 (O_821,N_4838,N_4998);
nand UO_822 (O_822,N_4868,N_4835);
and UO_823 (O_823,N_4887,N_4881);
or UO_824 (O_824,N_4868,N_4988);
and UO_825 (O_825,N_4917,N_4887);
or UO_826 (O_826,N_4995,N_4891);
and UO_827 (O_827,N_4835,N_4821);
or UO_828 (O_828,N_4879,N_4866);
and UO_829 (O_829,N_4973,N_4824);
and UO_830 (O_830,N_4910,N_4935);
nand UO_831 (O_831,N_4992,N_4983);
and UO_832 (O_832,N_4939,N_4865);
nor UO_833 (O_833,N_4947,N_4924);
and UO_834 (O_834,N_4864,N_4881);
and UO_835 (O_835,N_4834,N_4960);
and UO_836 (O_836,N_4973,N_4954);
and UO_837 (O_837,N_4943,N_4920);
nand UO_838 (O_838,N_4824,N_4900);
xnor UO_839 (O_839,N_4839,N_4986);
nand UO_840 (O_840,N_4917,N_4820);
nor UO_841 (O_841,N_4801,N_4936);
or UO_842 (O_842,N_4935,N_4886);
or UO_843 (O_843,N_4925,N_4846);
nor UO_844 (O_844,N_4808,N_4967);
nand UO_845 (O_845,N_4881,N_4953);
xor UO_846 (O_846,N_4973,N_4897);
nand UO_847 (O_847,N_4988,N_4865);
and UO_848 (O_848,N_4894,N_4914);
nor UO_849 (O_849,N_4983,N_4993);
nor UO_850 (O_850,N_4915,N_4882);
nand UO_851 (O_851,N_4872,N_4924);
or UO_852 (O_852,N_4897,N_4848);
and UO_853 (O_853,N_4869,N_4960);
or UO_854 (O_854,N_4831,N_4963);
or UO_855 (O_855,N_4989,N_4801);
nand UO_856 (O_856,N_4813,N_4816);
nor UO_857 (O_857,N_4998,N_4804);
or UO_858 (O_858,N_4834,N_4823);
and UO_859 (O_859,N_4811,N_4926);
and UO_860 (O_860,N_4899,N_4949);
and UO_861 (O_861,N_4996,N_4822);
nor UO_862 (O_862,N_4898,N_4972);
and UO_863 (O_863,N_4901,N_4940);
nand UO_864 (O_864,N_4817,N_4851);
or UO_865 (O_865,N_4978,N_4916);
or UO_866 (O_866,N_4806,N_4877);
nand UO_867 (O_867,N_4815,N_4899);
or UO_868 (O_868,N_4800,N_4990);
or UO_869 (O_869,N_4878,N_4935);
nor UO_870 (O_870,N_4920,N_4887);
nor UO_871 (O_871,N_4868,N_4817);
nand UO_872 (O_872,N_4937,N_4959);
nand UO_873 (O_873,N_4971,N_4866);
or UO_874 (O_874,N_4916,N_4971);
and UO_875 (O_875,N_4880,N_4992);
or UO_876 (O_876,N_4914,N_4998);
nor UO_877 (O_877,N_4916,N_4999);
and UO_878 (O_878,N_4803,N_4966);
nor UO_879 (O_879,N_4805,N_4903);
xor UO_880 (O_880,N_4885,N_4927);
nor UO_881 (O_881,N_4933,N_4904);
nor UO_882 (O_882,N_4911,N_4986);
or UO_883 (O_883,N_4806,N_4998);
nor UO_884 (O_884,N_4929,N_4967);
nor UO_885 (O_885,N_4802,N_4810);
or UO_886 (O_886,N_4905,N_4836);
nor UO_887 (O_887,N_4814,N_4848);
nand UO_888 (O_888,N_4967,N_4940);
nand UO_889 (O_889,N_4904,N_4945);
nor UO_890 (O_890,N_4997,N_4907);
or UO_891 (O_891,N_4933,N_4897);
nand UO_892 (O_892,N_4876,N_4931);
nand UO_893 (O_893,N_4957,N_4940);
or UO_894 (O_894,N_4980,N_4881);
and UO_895 (O_895,N_4888,N_4805);
nor UO_896 (O_896,N_4819,N_4917);
nand UO_897 (O_897,N_4830,N_4981);
nor UO_898 (O_898,N_4891,N_4877);
nor UO_899 (O_899,N_4951,N_4970);
and UO_900 (O_900,N_4813,N_4815);
or UO_901 (O_901,N_4942,N_4989);
nand UO_902 (O_902,N_4858,N_4894);
nand UO_903 (O_903,N_4925,N_4984);
nand UO_904 (O_904,N_4933,N_4814);
nand UO_905 (O_905,N_4878,N_4990);
nand UO_906 (O_906,N_4969,N_4981);
or UO_907 (O_907,N_4940,N_4891);
or UO_908 (O_908,N_4949,N_4960);
or UO_909 (O_909,N_4940,N_4803);
nand UO_910 (O_910,N_4803,N_4900);
or UO_911 (O_911,N_4843,N_4857);
nor UO_912 (O_912,N_4820,N_4803);
nand UO_913 (O_913,N_4983,N_4964);
and UO_914 (O_914,N_4978,N_4838);
nor UO_915 (O_915,N_4998,N_4860);
nor UO_916 (O_916,N_4975,N_4889);
nand UO_917 (O_917,N_4914,N_4857);
and UO_918 (O_918,N_4887,N_4842);
nor UO_919 (O_919,N_4903,N_4800);
and UO_920 (O_920,N_4950,N_4821);
or UO_921 (O_921,N_4995,N_4822);
or UO_922 (O_922,N_4861,N_4829);
nor UO_923 (O_923,N_4899,N_4854);
nand UO_924 (O_924,N_4995,N_4997);
and UO_925 (O_925,N_4965,N_4814);
nand UO_926 (O_926,N_4999,N_4951);
nand UO_927 (O_927,N_4954,N_4861);
and UO_928 (O_928,N_4946,N_4960);
or UO_929 (O_929,N_4829,N_4823);
and UO_930 (O_930,N_4873,N_4895);
and UO_931 (O_931,N_4894,N_4861);
nand UO_932 (O_932,N_4849,N_4874);
or UO_933 (O_933,N_4978,N_4935);
or UO_934 (O_934,N_4877,N_4940);
and UO_935 (O_935,N_4886,N_4940);
or UO_936 (O_936,N_4815,N_4801);
nor UO_937 (O_937,N_4814,N_4951);
nor UO_938 (O_938,N_4941,N_4998);
or UO_939 (O_939,N_4885,N_4881);
nor UO_940 (O_940,N_4981,N_4907);
nor UO_941 (O_941,N_4917,N_4800);
nand UO_942 (O_942,N_4996,N_4857);
or UO_943 (O_943,N_4801,N_4993);
nand UO_944 (O_944,N_4876,N_4889);
or UO_945 (O_945,N_4903,N_4822);
nand UO_946 (O_946,N_4863,N_4822);
nor UO_947 (O_947,N_4821,N_4842);
nor UO_948 (O_948,N_4958,N_4973);
nor UO_949 (O_949,N_4906,N_4942);
or UO_950 (O_950,N_4925,N_4940);
or UO_951 (O_951,N_4942,N_4988);
and UO_952 (O_952,N_4929,N_4876);
nor UO_953 (O_953,N_4801,N_4891);
nand UO_954 (O_954,N_4839,N_4863);
nor UO_955 (O_955,N_4971,N_4853);
or UO_956 (O_956,N_4941,N_4965);
and UO_957 (O_957,N_4943,N_4853);
and UO_958 (O_958,N_4806,N_4894);
nor UO_959 (O_959,N_4992,N_4957);
nor UO_960 (O_960,N_4930,N_4821);
nor UO_961 (O_961,N_4858,N_4980);
or UO_962 (O_962,N_4857,N_4958);
and UO_963 (O_963,N_4890,N_4889);
nand UO_964 (O_964,N_4999,N_4960);
nand UO_965 (O_965,N_4951,N_4900);
nand UO_966 (O_966,N_4828,N_4895);
nand UO_967 (O_967,N_4814,N_4823);
nand UO_968 (O_968,N_4842,N_4949);
or UO_969 (O_969,N_4931,N_4947);
nor UO_970 (O_970,N_4868,N_4860);
nor UO_971 (O_971,N_4876,N_4818);
or UO_972 (O_972,N_4832,N_4893);
or UO_973 (O_973,N_4877,N_4822);
nand UO_974 (O_974,N_4810,N_4932);
nor UO_975 (O_975,N_4931,N_4844);
and UO_976 (O_976,N_4853,N_4958);
and UO_977 (O_977,N_4941,N_4838);
nand UO_978 (O_978,N_4862,N_4961);
nand UO_979 (O_979,N_4892,N_4826);
or UO_980 (O_980,N_4812,N_4827);
nor UO_981 (O_981,N_4906,N_4999);
nand UO_982 (O_982,N_4802,N_4887);
and UO_983 (O_983,N_4900,N_4804);
or UO_984 (O_984,N_4977,N_4950);
nor UO_985 (O_985,N_4836,N_4869);
nand UO_986 (O_986,N_4908,N_4834);
and UO_987 (O_987,N_4967,N_4944);
nand UO_988 (O_988,N_4929,N_4998);
or UO_989 (O_989,N_4886,N_4960);
nor UO_990 (O_990,N_4962,N_4887);
nor UO_991 (O_991,N_4820,N_4994);
or UO_992 (O_992,N_4938,N_4947);
and UO_993 (O_993,N_4871,N_4867);
or UO_994 (O_994,N_4829,N_4880);
nor UO_995 (O_995,N_4859,N_4942);
nor UO_996 (O_996,N_4915,N_4863);
nor UO_997 (O_997,N_4938,N_4870);
and UO_998 (O_998,N_4829,N_4905);
or UO_999 (O_999,N_4816,N_4999);
endmodule